name mem_ctrl
i pi0000
i pi0001
i pi0002
i pi0003
i pi0004
i pi0005
i pi0006
i pi0007
i pi0008
i pi0009
i pi0010
i pi0011
i pi0012
i pi0013
i pi0014
i pi0015
i pi0016
i pi0017
i pi0018
i pi0019
i pi0020
i pi0021
i pi0022
i pi0023
i pi0024
i pi0025
i pi0026
i pi0027
i pi0028
i pi0029
i pi0030
i pi0031
i pi0032
i pi0033
i pi0034
i pi0035
i pi0036
i pi0037
i pi0038
i pi0039
i pi0040
i pi0041
i pi0042
i pi0043
i pi0044
i pi0045
i pi0046
i pi0047
i pi0048
i pi0049
i pi0050
i pi0051
i pi0052
i pi0053
i pi0054
i pi0055
i pi0056
i pi0057
i pi0058
i pi0059
i pi0060
i pi0061
i pi0062
i pi0063
i pi0064
i pi0065
i pi0066
i pi0067
i pi0068
i pi0069
i pi0070
i pi0071
i pi0072
i pi0073
i pi0074
i pi0075
i pi0076
i pi0077
i pi0078
i pi0079
i pi0080
i pi0081
i pi0082
i pi0083
i pi0084
i pi0085
i pi0086
i pi0087
i pi0088
i pi0089
i pi0090
i pi0091
i pi0092
i pi0093
i pi0094
i pi0095
i pi0096
i pi0097
i pi0098
i pi0099
i pi0100
i pi0101
i pi0102
i pi0103
i pi0104
i pi0105
i pi0106
i pi0107
i pi0108
i pi0109
i pi0110
i pi0111
i pi0112
i pi0113
i pi0114
i pi0115
i pi0116
i pi0117
i pi0118
i pi0119
i pi0120
i pi0121
i pi0122
i pi0123
i pi0124
i pi0125
i pi0126
i pi0127
i pi0128
i pi0129
i pi0130
i pi0131
i pi0132
i pi0133
i pi0134
i pi0135
i pi0136
i pi0137
i pi0138
i pi0139
i pi0140
i pi0141
i pi0142
i pi0143
i pi0144
i pi0145
i pi0146
i pi0147
i pi0148
i pi0149
i pi0150
i pi0151
i pi0152
i pi0153
i pi0154
i pi0155
i pi0156
i pi0157
i pi0158
i pi0159
i pi0160
i pi0161
i pi0162
i pi0163
i pi0164
i pi0165
i pi0166
i pi0167
i pi0168
i pi0169
i pi0170
i pi0171
i pi0172
i pi0173
i pi0174
i pi0175
i pi0176
i pi0177
i pi0178
i pi0179
i pi0180
i pi0181
i pi0182
i pi0183
i pi0184
i pi0185
i pi0186
i pi0187
i pi0188
i pi0189
i pi0190
i pi0191
i pi0192
i pi0193
i pi0194
i pi0195
i pi0196
i pi0197
i pi0198
i pi0199
i pi0200
i pi0201
i pi0202
i pi0203
i pi0204
i pi0205
i pi0206
i pi0207
i pi0208
i pi0209
i pi0210
i pi0211
i pi0212
i pi0213
i pi0214
i pi0215
i pi0216
i pi0217
i pi0218
i pi0219
i pi0220
i pi0221
i pi0222
i pi0223
i pi0224
i pi0225
i pi0226
i pi0227
i pi0228
i pi0229
i pi0230
i pi0231
i pi0232
i pi0233
i pi0234
i pi0235
i pi0236
i pi0237
i pi0238
i pi0239
i pi0240
i pi0241
i pi0242
i pi0243
i pi0244
i pi0245
i pi0246
i pi0247
i pi0248
i pi0249
i pi0250
i pi0251
i pi0252
i pi0253
i pi0254
i pi0255
i pi0256
i pi0257
i pi0258
i pi0259
i pi0260
i pi0261
i pi0262
i pi0263
i pi0264
i pi0265
i pi0266
i pi0267
i pi0268
i pi0269
i pi0270
i pi0271
i pi0272
i pi0273
i pi0274
i pi0275
i pi0276
i pi0277
i pi0278
i pi0279
i pi0280
i pi0281
i pi0282
i pi0283
i pi0284
i pi0285
i pi0286
i pi0287
i pi0288
i pi0289
i pi0290
i pi0291
i pi0292
i pi0293
i pi0294
i pi0295
i pi0296
i pi0297
i pi0298
i pi0299
i pi0300
i pi0301
i pi0302
i pi0303
i pi0304
i pi0305
i pi0306
i pi0307
i pi0308
i pi0309
i pi0310
i pi0311
i pi0312
i pi0313
i pi0314
i pi0315
i pi0316
i pi0317
i pi0318
i pi0319
i pi0320
i pi0321
i pi0322
i pi0323
i pi0324
i pi0325
i pi0326
i pi0327
i pi0328
i pi0329
i pi0330
i pi0331
i pi0332
i pi0333
i pi0334
i pi0335
i pi0336
i pi0337
i pi0338
i pi0339
i pi0340
i pi0341
i pi0342
i pi0343
i pi0344
i pi0345
i pi0346
i pi0347
i pi0348
i pi0349
i pi0350
i pi0351
i pi0352
i pi0353
i pi0354
i pi0355
i pi0356
i pi0357
i pi0358
i pi0359
i pi0360
i pi0361
i pi0362
i pi0363
i pi0364
i pi0365
i pi0366
i pi0367
i pi0368
i pi0369
i pi0370
i pi0371
i pi0372
i pi0373
i pi0374
i pi0375
i pi0376
i pi0377
i pi0378
i pi0379
i pi0380
i pi0381
i pi0382
i pi0383
i pi0384
i pi0385
i pi0386
i pi0387
i pi0388
i pi0389
i pi0390
i pi0391
i pi0392
i pi0393
i pi0394
i pi0395
i pi0396
i pi0397
i pi0398
i pi0399
i pi0400
i pi0401
i pi0402
i pi0403
i pi0404
i pi0405
i pi0406
i pi0407
i pi0408
i pi0409
i pi0410
i pi0411
i pi0412
i pi0413
i pi0414
i pi0415
i pi0416
i pi0417
i pi0418
i pi0419
i pi0420
i pi0421
i pi0422
i pi0423
i pi0424
i pi0425
i pi0426
i pi0427
i pi0428
i pi0429
i pi0430
i pi0431
i pi0432
i pi0433
i pi0434
i pi0435
i pi0436
i pi0437
i pi0438
i pi0439
i pi0440
i pi0441
i pi0442
i pi0443
i pi0444
i pi0445
i pi0446
i pi0447
i pi0448
i pi0449
i pi0450
i pi0451
i pi0452
i pi0453
i pi0454
i pi0455
i pi0456
i pi0457
i pi0458
i pi0459
i pi0460
i pi0461
i pi0462
i pi0463
i pi0464
i pi0465
i pi0466
i pi0467
i pi0468
i pi0469
i pi0470
i pi0471
i pi0472
i pi0473
i pi0474
i pi0475
i pi0476
i pi0477
i pi0478
i pi0479
i pi0480
i pi0481
i pi0482
i pi0483
i pi0484
i pi0485
i pi0486
i pi0487
i pi0488
i pi0489
i pi0490
i pi0491
i pi0492
i pi0493
i pi0494
i pi0495
i pi0496
i pi0497
i pi0498
i pi0499
i pi0500
i pi0501
i pi0502
i pi0503
i pi0504
i pi0505
i pi0506
i pi0507
i pi0508
i pi0509
i pi0510
i pi0511
i pi0512
i pi0513
i pi0514
i pi0515
i pi0516
i pi0517
i pi0518
i pi0519
i pi0520
i pi0521
i pi0522
i pi0523
i pi0524
i pi0525
i pi0526
i pi0527
i pi0528
i pi0529
i pi0530
i pi0531
i pi0532
i pi0533
i pi0534
i pi0535
i pi0536
i pi0537
i pi0538
i pi0539
i pi0540
i pi0541
i pi0542
i pi0543
i pi0544
i pi0545
i pi0546
i pi0547
i pi0548
i pi0549
i pi0550
i pi0551
i pi0552
i pi0553
i pi0554
i pi0555
i pi0556
i pi0557
i pi0558
i pi0559
i pi0560
i pi0561
i pi0562
i pi0563
i pi0564
i pi0565
i pi0566
i pi0567
i pi0568
i pi0569
i pi0570
i pi0571
i pi0572
i pi0573
i pi0574
i pi0575
i pi0576
i pi0577
i pi0578
i pi0579
i pi0580
i pi0581
i pi0582
i pi0583
i pi0584
i pi0585
i pi0586
i pi0587
i pi0588
i pi0589
i pi0590
i pi0591
i pi0592
i pi0593
i pi0594
i pi0595
i pi0596
i pi0597
i pi0598
i pi0599
i pi0600
i pi0601
i pi0602
i pi0603
i pi0604
i pi0605
i pi0606
i pi0607
i pi0608
i pi0609
i pi0610
i pi0611
i pi0612
i pi0613
i pi0614
i pi0615
i pi0616
i pi0617
i pi0618
i pi0619
i pi0620
i pi0621
i pi0622
i pi0623
i pi0624
i pi0625
i pi0626
i pi0627
i pi0628
i pi0629
i pi0630
i pi0631
i pi0632
i pi0633
i pi0634
i pi0635
i pi0636
i pi0637
i pi0638
i pi0639
i pi0640
i pi0641
i pi0642
i pi0643
i pi0644
i pi0645
i pi0646
i pi0647
i pi0648
i pi0649
i pi0650
i pi0651
i pi0652
i pi0653
i pi0654
i pi0655
i pi0656
i pi0657
i pi0658
i pi0659
i pi0660
i pi0661
i pi0662
i pi0663
i pi0664
i pi0665
i pi0666
i pi0667
i pi0668
i pi0669
i pi0670
i pi0671
i pi0672
i pi0673
i pi0674
i pi0675
i pi0676
i pi0677
i pi0678
i pi0679
i pi0680
i pi0681
i pi0682
i pi0683
i pi0684
i pi0685
i pi0686
i pi0687
i pi0688
i pi0689
i pi0690
i pi0691
i pi0692
i pi0693
i pi0694
i pi0695
i pi0696
i pi0697
i pi0698
i pi0699
i pi0700
i pi0701
i pi0702
i pi0703
i pi0704
i pi0705
i pi0706
i pi0707
i pi0708
i pi0709
i pi0710
i pi0711
i pi0712
i pi0713
i pi0714
i pi0715
i pi0716
i pi0717
i pi0718
i pi0719
i pi0720
i pi0721
i pi0722
i pi0723
i pi0724
i pi0725
i pi0726
i pi0727
i pi0728
i pi0729
i pi0730
i pi0731
i pi0732
i pi0733
i pi0734
i pi0735
i pi0736
i pi0737
i pi0738
i pi0739
i pi0740
i pi0741
i pi0742
i pi0743
i pi0744
i pi0745
i pi0746
i pi0747
i pi0748
i pi0749
i pi0750
i pi0751
i pi0752
i pi0753
i pi0754
i pi0755
i pi0756
i pi0757
i pi0758
i pi0759
i pi0760
i pi0761
i pi0762
i pi0763
i pi0764
i pi0765
i pi0766
i pi0767
i pi0768
i pi0769
i pi0770
i pi0771
i pi0772
i pi0773
i pi0774
i pi0775
i pi0776
i pi0777
i pi0778
i pi0779
i pi0780
i pi0781
i pi0782
i pi0783
i pi0784
i pi0785
i pi0786
i pi0787
i pi0788
i pi0789
i pi0790
i pi0791
i pi0792
i pi0793
i pi0794
i pi0795
i pi0796
i pi0797
i pi0798
i pi0799
i pi0800
i pi0801
i pi0802
i pi0803
i pi0804
i pi0805
i pi0806
i pi0807
i pi0808
i pi0809
i pi0810
i pi0811
i pi0812
i pi0813
i pi0814
i pi0815
i pi0816
i pi0817
i pi0818
i pi0819
i pi0820
i pi0821
i pi0822
i pi0823
i pi0824
i pi0825
i pi0826
i pi0827
i pi0828
i pi0829
i pi0830
i pi0831
i pi0832
i pi0833
i pi0834
i pi0835
i pi0836
i pi0837
i pi0838
i pi0839
i pi0840
i pi0841
i pi0842
i pi0843
i pi0844
i pi0845
i pi0846
i pi0847
i pi0848
i pi0849
i pi0850
i pi0851
i pi0852
i pi0853
i pi0854
i pi0855
i pi0856
i pi0857
i pi0858
i pi0859
i pi0860
i pi0861
i pi0862
i pi0863
i pi0864
i pi0865
i pi0866
i pi0867
i pi0868
i pi0869
i pi0870
i pi0871
i pi0872
i pi0873
i pi0874
i pi0875
i pi0876
i pi0877
i pi0878
i pi0879
i pi0880
i pi0881
i pi0882
i pi0883
i pi0884
i pi0885
i pi0886
i pi0887
i pi0888
i pi0889
i pi0890
i pi0891
i pi0892
i pi0893
i pi0894
i pi0895
i pi0896
i pi0897
i pi0898
i pi0899
i pi0900
i pi0901
i pi0902
i pi0903
i pi0904
i pi0905
i pi0906
i pi0907
i pi0908
i pi0909
i pi0910
i pi0911
i pi0912
i pi0913
i pi0914
i pi0915
i pi0916
i pi0917
i pi0918
i pi0919
i pi0920
i pi0921
i pi0922
i pi0923
i pi0924
i pi0925
i pi0926
i pi0927
i pi0928
i pi0929
i pi0930
i pi0931
i pi0932
i pi0933
i pi0934
i pi0935
i pi0936
i pi0937
i pi0938
i pi0939
i pi0940
i pi0941
i pi0942
i pi0943
i pi0944
i pi0945
i pi0946
i pi0947
i pi0948
i pi0949
i pi0950
i pi0951
i pi0952
i pi0953
i pi0954
i pi0955
i pi0956
i pi0957
i pi0958
i pi0959
i pi0960
i pi0961
i pi0962
i pi0963
i pi0964
i pi0965
i pi0966
i pi0967
i pi0968
i pi0969
i pi0970
i pi0971
i pi0972
i pi0973
i pi0974
i pi0975
i pi0976
i pi0977
i pi0978
i pi0979
i pi0980
i pi0981
i pi0982
i pi0983
i pi0984
i pi0985
i pi0986
i pi0987
i pi0988
i pi0989
i pi0990
i pi0991
i pi0992
i pi0993
i pi0994
i pi0995
i pi0996
i pi0997
i pi0998
i pi0999
i pi1000
i pi1001
i pi1002
i pi1003
i pi1004
i pi1005
i pi1006
i pi1007
i pi1008
i pi1009
i pi1010
i pi1011
i pi1012
i pi1013
i pi1014
i pi1015
i pi1016
i pi1017
i pi1018
i pi1019
i pi1020
i pi1021
i pi1022
i pi1023
i pi1024
i pi1025
i pi1026
i pi1027
i pi1028
i pi1029
i pi1030
i pi1031
i pi1032
i pi1033
i pi1034
i pi1035
i pi1036
i pi1037
i pi1038
i pi1039
i pi1040
i pi1041
i pi1042
i pi1043
i pi1044
i pi1045
i pi1046
i pi1047
i pi1048
i pi1049
i pi1050
i pi1051
i pi1052
i pi1053
i pi1054
i pi1055
i pi1056
i pi1057
i pi1058
i pi1059
i pi1060
i pi1061
i pi1062
i pi1063
i pi1064
i pi1065
i pi1066
i pi1067
i pi1068
i pi1069
i pi1070
i pi1071
i pi1072
i pi1073
i pi1074
i pi1075
i pi1076
i pi1077
i pi1078
i pi1079
i pi1080
i pi1081
i pi1082
i pi1083
i pi1084
i pi1085
i pi1086
i pi1087
i pi1088
i pi1089
i pi1090
i pi1091
i pi1092
i pi1093
i pi1094
i pi1095
i pi1096
i pi1097
i pi1098
i pi1099
i pi1100
i pi1101
i pi1102
i pi1103
i pi1104
i pi1105
i pi1106
i pi1107
i pi1108
i pi1109
i pi1110
i pi1111
i pi1112
i pi1113
i pi1114
i pi1115
i pi1116
i pi1117
i pi1118
i pi1119
i pi1120
i pi1121
i pi1122
i pi1123
i pi1124
i pi1125
i pi1126
i pi1127
i pi1128
i pi1129
i pi1130
i pi1131
i pi1132
i pi1133
i pi1134
i pi1135
i pi1136
i pi1137
i pi1138
i pi1139
i pi1140
i pi1141
i pi1142
i pi1143
i pi1144
i pi1145
i pi1146
i pi1147
i pi1148
i pi1149
i pi1150
i pi1151
i pi1152
i pi1153
i pi1154
i pi1155
i pi1156
i pi1157
i pi1158
i pi1159
i pi1160
i pi1161
i pi1162
i pi1163
i pi1164
i pi1165
i pi1166
i pi1167
i pi1168
i pi1169
i pi1170
i pi1171
i pi1172
i pi1173
i pi1174
i pi1175
i pi1176
i pi1177
i pi1178
i pi1179
i pi1180
i pi1181
i pi1182
i pi1183
i pi1184
i pi1185
i pi1186
i pi1187
i pi1188
i pi1189
i pi1190
i pi1191
i pi1192
i pi1193
i pi1194
i pi1195
i pi1196
i pi1197
i pi1198
i pi1199
i pi1200
i pi1201
i pi1202
i pi1203

o po0000
o po0001
o po0002
o po0003
o po0004
o po0005
o po0006
o po0007
o po0008
o po0009
o po0010
o po0011
o po0012
o po0013
o po0014
o po0015
o po0016
o po0017
o po0018
o po0019
o po0020
o po0021
o po0022
o po0023
o po0024
o po0025
o po0026
o po0027
o po0028
o po0029
o po0030
o po0031
o po0032
o po0033
o po0034
o po0035
o po0036
o po0037
o po0038
o po0039
o po0040
o po0041
o po0042
o po0043
o po0044
o po0045
o po0046
o po0047
o po0048
o po0049
o po0050
o po0051
o po0052
o po0053
o po0054
o po0055
o po0056
o po0057
o po0058
o po0059
o po0060
o po0061
o po0062
o po0063
o po0064
o po0065
o po0066
o po0067
o po0068
o po0069
o po0070
o po0071
o po0072
o po0073
o po0074
o po0075
o po0076
o po0077
o po0078
o po0079
o po0080
o po0081
o po0082
o po0083
o po0084
o po0085
o po0086
o po0087
o po0088
o po0089
o po0090
o po0091
o po0092
o po0093
o po0094
o po0095
o po0096
o po0097
o po0098
o po0099
o po0100
o po0101
o po0102
o po0103
o po0104
o po0105
o po0106
o po0107
o po0108
o po0109
o po0110
o po0111
o po0112
o po0113
o po0114
o po0115
o po0116
o po0117
o po0118
o po0119
o po0120
o po0121
o po0122
o po0123
o po0124
o po0125
o po0126
o po0127
o po0128
o po0129
o po0130
o po0131
o po0132
o po0133
o po0134
o po0135
o po0136
o po0137
o po0138
o po0139
o po0140
o po0141
o po0142
o po0143
o po0144
o po0145
o po0146
o po0147
o po0148
o po0149
o po0150
o po0151
o po0152
o po0153
o po0154
o po0155
o po0156
o po0157
o po0158
o po0159
o po0160
o po0161
o po0162
o po0163
o po0164
o po0165
o po0166
o po0167
o po0168
o po0169
o po0170
o po0171
o po0172
o po0173
o po0174
o po0175
o po0176
o po0177
o po0178
o po0179
o po0180
o po0181
o po0182
o po0183
o po0184
o po0185
o po0186
o po0187
o po0188
o po0189
o po0190
o po0191
o po0192
o po0193
o po0194
o po0195
o po0196
o po0197
o po0198
o po0199
o po0200
o po0201
o po0202
o po0203
o po0204
o po0205
o po0206
o po0207
o po0208
o po0209
o po0210
o po0211
o po0212
o po0213
o po0214
o po0215
o po0216
o po0217
o po0218
o po0219
o po0220
o po0221
o po0222
o po0223
o po0224
o po0225
o po0226
o po0227
o po0228
o po0229
o po0230
o po0231
o po0232
o po0233
o po0234
o po0235
o po0236
o po0237
o po0238
o po0239
o po0240
o po0241
o po0242
o po0243
o po0244
o po0245
o po0246
o po0247
o po0248
o po0249
o po0250
o po0251
o po0252
o po0253
o po0254
o po0255
o po0256
o po0257
o po0258
o po0259
o po0260
o po0261
o po0262
o po0263
o po0264
o po0265
o po0266
o po0267
o po0268
o po0269
o po0270
o po0271
o po0272
o po0273
o po0274
o po0275
o po0276
o po0277
o po0278
o po0279
o po0280
o po0281
o po0282
o po0283
o po0284
o po0285
o po0286
o po0287
o po0288
o po0289
o po0290
o po0291
o po0292
o po0293
o po0294
o po0295
o po0296
o po0297
o po0298
o po0299
o po0300
o po0301
o po0302
o po0303
o po0304
o po0305
o po0306
o po0307
o po0308
o po0309
o po0310
o po0311
o po0312
o po0313
o po0314
o po0315
o po0316
o po0317
o po0318
o po0319
o po0320
o po0321
o po0322
o po0323
o po0324
o po0325
o po0326
o po0327
o po0328
o po0329
o po0330
o po0331
o po0332
o po0333
o po0334
o po0335
o po0336
o po0337
o po0338
o po0339
o po0340
o po0341
o po0342
o po0343
o po0344
o po0345
o po0346
o po0347
o po0348
o po0349
o po0350
o po0351
o po0352
o po0353
o po0354
o po0355
o po0356
o po0357
o po0358
o po0359
o po0360
o po0361
o po0362
o po0363
o po0364
o po0365
o po0366
o po0367
o po0368
o po0369
o po0370
o po0371
o po0372
o po0373
o po0374
o po0375
o po0376
o po0377
o po0378
o po0379
o po0380
o po0381
o po0382
o po0383
o po0384
o po0385
o po0386
o po0387
o po0388
o po0389
o po0390
o po0391
o po0392
o po0393
o po0394
o po0395
o po0396
o po0397
o po0398
o po0399
o po0400
o po0401
o po0402
o po0403
o po0404
o po0405
o po0406
o po0407
o po0408
o po0409
o po0410
o po0411
o po0412
o po0413
o po0414
o po0415
o po0416
o po0417
o po0418
o po0419
o po0420
o po0421
o po0422
o po0423
o po0424
o po0425
o po0426
o po0427
o po0428
o po0429
o po0430
o po0431
o po0432
o po0433
o po0434
o po0435
o po0436
o po0437
o po0438
o po0439
o po0440
o po0441
o po0442
o po0443
o po0444
o po0445
o po0446
o po0447
o po0448
o po0449
o po0450
o po0451
o po0452
o po0453
o po0454
o po0455
o po0456
o po0457
o po0458
o po0459
o po0460
o po0461
o po0462
o po0463
o po0464
o po0465
o po0466
o po0467
o po0468
o po0469
o po0470
o po0471
o po0472
o po0473
o po0474
o po0475
o po0476
o po0477
o po0478
o po0479
o po0480
o po0481
o po0482
o po0483
o po0484
o po0485
o po0486
o po0487
o po0488
o po0489
o po0490
o po0491
o po0492
o po0493
o po0494
o po0495
o po0496
o po0497
o po0498
o po0499
o po0500
o po0501
o po0502
o po0503
o po0504
o po0505
o po0506
o po0507
o po0508
o po0509
o po0510
o po0511
o po0512
o po0513
o po0514
o po0515
o po0516
o po0517
o po0518
o po0519
o po0520
o po0521
o po0522
o po0523
o po0524
o po0525
o po0526
o po0527
o po0528
o po0529
o po0530
o po0531
o po0532
o po0533
o po0534
o po0535
o po0536
o po0537
o po0538
o po0539
o po0540
o po0541
o po0542
o po0543
o po0544
o po0545
o po0546
o po0547
o po0548
o po0549
o po0550
o po0551
o po0552
o po0553
o po0554
o po0555
o po0556
o po0557
o po0558
o po0559
o po0560
o po0561
o po0562
o po0563
o po0564
o po0565
o po0566
o po0567
o po0568
o po0569
o po0570
o po0571
o po0572
o po0573
o po0574
o po0575
o po0576
o po0577
o po0578
o po0579
o po0580
o po0581
o po0582
o po0583
o po0584
o po0585
o po0586
o po0587
o po0588
o po0589
o po0590
o po0591
o po0592
o po0593
o po0594
o po0595
o po0596
o po0597
o po0598
o po0599
o po0600
o po0601
o po0602
o po0603
o po0604
o po0605
o po0606
o po0607
o po0608
o po0609
o po0610
o po0611
o po0612
o po0613
o po0614
o po0615
o po0616
o po0617
o po0618
o po0619
o po0620
o po0621
o po0622
o po0623
o po0624
o po0625
o po0626
o po0627
o po0628
o po0629
o po0630
o po0631
o po0632
o po0633
o po0634
o po0635
o po0636
o po0637
o po0638
o po0639
o po0640
o po0641
o po0642
o po0643
o po0644
o po0645
o po0646
o po0647
o po0648
o po0649
o po0650
o po0651
o po0652
o po0653
o po0654
o po0655
o po0656
o po0657
o po0658
o po0659
o po0660
o po0661
o po0662
o po0663
o po0664
o po0665
o po0666
o po0667
o po0668
o po0669
o po0670
o po0671
o po0672
o po0673
o po0674
o po0675
o po0676
o po0677
o po0678
o po0679
o po0680
o po0681
o po0682
o po0683
o po0684
o po0685
o po0686
o po0687
o po0688
o po0689
o po0690
o po0691
o po0692
o po0693
o po0694
o po0695
o po0696
o po0697
o po0698
o po0699
o po0700
o po0701
o po0702
o po0703
o po0704
o po0705
o po0706
o po0707
o po0708
o po0709
o po0710
o po0711
o po0712
o po0713
o po0714
o po0715
o po0716
o po0717
o po0718
o po0719
o po0720
o po0721
o po0722
o po0723
o po0724
o po0725
o po0726
o po0727
o po0728
o po0729
o po0730
o po0731
o po0732
o po0733
o po0734
o po0735
o po0736
o po0737
o po0738
o po0739
o po0740
o po0741
o po0742
o po0743
o po0744
o po0745
o po0746
o po0747
o po0748
o po0749
o po0750
o po0751
o po0752
o po0753
o po0754
o po0755
o po0756
o po0757
o po0758
o po0759
o po0760
o po0761
o po0762
o po0763
o po0764
o po0765
o po0766
o po0767
o po0768
o po0769
o po0770
o po0771
o po0772
o po0773
o po0774
o po0775
o po0776
o po0777
o po0778
o po0779
o po0780
o po0781
o po0782
o po0783
o po0784
o po0785
o po0786
o po0787
o po0788
o po0789
o po0790
o po0791
o po0792
o po0793
o po0794
o po0795
o po0796
o po0797
o po0798
o po0799
o po0800
o po0801
o po0802
o po0803
o po0804
o po0805
o po0806
o po0807
o po0808
o po0809
o po0810
o po0811
o po0812
o po0813
o po0814
o po0815
o po0816
o po0817
o po0818
o po0819
o po0820
o po0821
o po0822
o po0823
o po0824
o po0825
o po0826
o po0827
o po0828
o po0829
o po0830
o po0831
o po0832
o po0833
o po0834
o po0835
o po0836
o po0837
o po0838
o po0839
o po0840
o po0841
o po0842
o po0843
o po0844
o po0845
o po0846
o po0847
o po0848
o po0849
o po0850
o po0851
o po0852
o po0853
o po0854
o po0855
o po0856
o po0857
o po0858
o po0859
o po0860
o po0861
o po0862
o po0863
o po0864
o po0865
o po0866
o po0867
o po0868
o po0869
o po0870
o po0871
o po0872
o po0873
o po0874
o po0875
o po0876
o po0877
o po0878
o po0879
o po0880
o po0881
o po0882
o po0883
o po0884
o po0885
o po0886
o po0887
o po0888
o po0889
o po0890
o po0891
o po0892
o po0893
o po0894
o po0895
o po0896
o po0897
o po0898
o po0899
o po0900
o po0901
o po0902
o po0903
o po0904
o po0905
o po0906
o po0907
o po0908
o po0909
o po0910
o po0911
o po0912
o po0913
o po0914
o po0915
o po0916
o po0917
o po0918
o po0919
o po0920
o po0921
o po0922
o po0923
o po0924
o po0925
o po0926
o po0927
o po0928
o po0929
o po0930
o po0931
o po0932
o po0933
o po0934
o po0935
o po0936
o po0937
o po0938
o po0939
o po0940
o po0941
o po0942
o po0943
o po0944
o po0945
o po0946
o po0947
o po0948
o po0949
o po0950
o po0951
o po0952
o po0953
o po0954
o po0955
o po0956
o po0957
o po0958
o po0959
o po0960
o po0961
o po0962
o po0963
o po0964
o po0965
o po0966
o po0967
o po0968
o po0969
o po0970
o po0971
o po0972
o po0973
o po0974
o po0975
o po0976
o po0977
o po0978
o po0979
o po0980
o po0981
o po0982
o po0983
o po0984
o po0985
o po0986
o po0987
o po0988
o po0989
o po0990
o po0991
o po0992
o po0993
o po0994
o po0995
o po0996
o po0997
o po0998
o po0999
o po1000
o po1001
o po1002
o po1003
o po1004
o po1005
o po1006
o po1007
o po1008
o po1009
o po1010
o po1011
o po1012
o po1013
o po1014
o po1015
o po1016
o po1017
o po1018
o po1019
o po1020
o po1021
o po1022
o po1023
o po1024
o po1025
o po1026
o po1027
o po1028
o po1029
o po1030
o po1031
o po1032
o po1033
o po1034
o po1035
o po1036
o po1037
o po1038
o po1039
o po1040
o po1041
o po1042
o po1043
o po1044
o po1045
o po1046
o po1047
o po1048
o po1049
o po1050
o po1051
o po1052
o po1053
o po1054
o po1055
o po1056
o po1057
o po1058
o po1059
o po1060
o po1061
o po1062
o po1063
o po1064
o po1065
o po1066
o po1067
o po1068
o po1069
o po1070
o po1071
o po1072
o po1073
o po1074
o po1075
o po1076
o po1077
o po1078
o po1079
o po1080
o po1081
o po1082
o po1083
o po1084
o po1085
o po1086
o po1087
o po1088
o po1089
o po1090
o po1091
o po1092
o po1093
o po1094
o po1095
o po1096
o po1097
o po1098
o po1099
o po1100
o po1101
o po1102
o po1103
o po1104
o po1105
o po1106
o po1107
o po1108
o po1109
o po1110
o po1111
o po1112
o po1113
o po1114
o po1115
o po1116
o po1117
o po1118
o po1119
o po1120
o po1121
o po1122
o po1123
o po1124
o po1125
o po1126
o po1127
o po1128
o po1129
o po1130
o po1131
o po1132
o po1133
o po1134
o po1135
o po1136
o po1137
o po1138
o po1139
o po1140
o po1141
o po1142
o po1143
o po1144
o po1145
o po1146
o po1147
o po1148
o po1149
o po1150
o po1151
o po1152
o po1153
o po1154
o po1155
o po1156
o po1157
o po1158
o po1159
o po1160
o po1161
o po1162
o po1163
o po1164
o po1165
o po1166
o po1167
o po1168
o po1169
o po1170
o po1171
o po1172
o po1173
o po1174
o po1175
o po1176
o po1177
o po1178
o po1179
o po1180
o po1181
o po1182
o po1183
o po1184
o po1185
o po1186
o po1187
o po1188
o po1189
o po1190
o po1191
o po1192
o po1193
o po1194
o po1195
o po1196
o po1197
o po1198
o po1199
o po1200
o po1201
o po1202
o po1203
o po1204
o po1205
o po1206
o po1207
o po1208
o po1209
o po1210
o po1211
o po1212
o po1213
o po1214
o po1215
o po1216
o po1217
o po1218
o po1219
o po1220
o po1221
o po1222
o po1223
o po1224
o po1225
o po1226
o po1227
o po1228
o po1229
o po1230

g1 nor pi0332 pi1144 ; n2437
g2 and pi0215 n2437_not ; n2438
g3 and pi0265 pi0332_not ; n2439
g4 and pi0216 n2439_not ; n2440
g5 and pi0105 pi0228 ; n2441
g6 and pi0095 pi0479_not ; n2442
g7 and pi0234 n2442 ; n2443
g8 nor pi0332 n2443 ; n2444
g9 and n2441 n2444 ; n2445
g10 and pi0153 pi0332_not ; n2446
g11 and n2441_not n2446 ; n2447
g12 nor pi0216 n2447 ; n2448
g13 and n2445_not n2448 ; n2449
g14 nor n2440 n2449 ; n2450
g15 nor pi0221 n2450 ; n2451
g16 and pi0216_not pi0833 ; n2452
g17 and pi1144 n2452_not ; n2453
g18 and pi0929 n2452 ; n2454
g19 nor pi0332 n2453 ; n2455
g20 and n2454_not n2455 ; n2456
g21 and pi0221 n2456_not ; n2457
g22 nor n2451 n2457 ; n2458
g23 nor pi0215 n2458 ; n2459
g24 nor n2438 n2459 ; n2460
g25 nor pi0058 pi0090 ; n2461
g26 nor pi0088 pi0098 ; n2462
g27 and pi0077_not n2462 ; n2463
g28 and pi0050_not n2463 ; n2464
g29 and pi0102_not n2464 ; n2465
g30 nor pi0065 pi0071 ; n2466
g31 nor pi0083 pi0103 ; n2467
g32 nor pi0067 pi0069 ; n2468
g33 nor pi0066 pi0073 ; n2469
g34 nor pi0061 pi0076 ; n2470
g35 nor pi0085 pi0106 ; n2471
g36 and n2470 n2471 ; n2472
g37 and pi0048_not n2472 ; n2473
g38 and pi0089_not n2473 ; n2474
g39 and pi0049_not n2474 ; n2475
g40 and pi0104_not n2475 ; n2476
g41 and pi0045_not n2476 ; n2477
g42 nor pi0068 pi0084 ; n2478
g43 nor pi0082 pi0111 ; n2479
g44 and pi0036_not n2479 ; n2480
g45 and n2478 n2480 ; n2481
g46 and n2477 n2481 ; n2482
g47 and n2469 n2482 ; n2483
g48 and n2468 n2483 ; n2484
g49 and n2467 n2484 ; n2485
g50 and n2466 n2485 ; n2486
g51 nor pi0063 pi0107 ; n2487
g52 and n2486 n2487 ; n2488
g53 and pi0064_not n2488 ; n2489
g54 and pi0081_not n2489 ; n2490
g55 and n2465 n2490 ; n2491
g56 nor pi0047 pi0091 ; n2492
g57 nor pi0109 pi0110 ; n2493
g58 nor pi0053 pi0060 ; n2494
g59 and pi0086_not n2494 ; n2495
g60 nor pi0097 pi0108 ; n2496
g61 and pi0094_not n2496 ; n2497
g62 and pi0046_not n2495 ; n2498
g63 and n2497 n2498 ; n2499
g64 and n2493 n2499 ; n2500
g65 and n2492 n2500 ; n2501
g66 and n2491 n2501 ; n2502
g67 and n2461 n2502 ; n2503
g68 nor pi0035 pi0093 ; n2504
g69 and n2503 n2504 ; n2505
g70 nor pi0072 pi0096 ; n2506
g71 nor pi0051 pi0070 ; n2507
g72 and n2506 n2507 ; n2508
g73 and n2505 n2508 ; n2509
g74 nor pi0032 pi0040 ; n2510
g75 and n2509 n2510 ; n2511
g76 and pi0095_not n2511 ; n2512
g77 nor n2442 n2512 ; n2513
g78 and pi0234 n2513_not ; n2514
g79 and pi0070_not n2505 ; n2515
g80 nor pi0051 pi0096 ; n2516
g81 nor pi0040 pi0072 ; n2517
g82 nor pi0032 pi0095 ; n2518
g83 and n2517 n2518 ; n2519
g84 and n2516 n2519 ; n2520
g85 and n2515 n2520 ; n2521
g86 and pi0234_not n2521 ; n2522
g87 nor n2514 n2522 ; n2523
g88 and pi0137 n2523_not ; n2524
g89 and n2444 n2524_not ; n2525
g90 nor pi0215 pi0221 ; n2526
g91 and n2448 n2526 ; n2527
g92 and n2525_not n2527 ; n2528
g93 nor pi0056 pi0062 ; n2529
g94 nor pi0038 pi0039 ; n2530
g95 and pi0100_not n2530 ; n2531
g96 nor pi0054 pi0074 ; n2532
g97 nor pi0075 pi0087 ; n2533
g98 and pi0092_not n2533 ; n2534
g99 and n2532 n2534 ; n2535
g100 and pi0055_not n2535 ; n2536
g101 and n2531 n2536 ; n2537
g102 and n2529 n2537 ; n2538
g103 and n2528 n2538 ; n2539
g104 and pi0059 n2460 ; n2540
g105 and n2539_not n2540 ; n2541
g106 and n2460 n2537_not ; n2542
g107 nor pi0105 n2446 ; n2543
g108 and pi0105 n2525_not ; n2544
g109 nor n2543 n2544 ; n2545
g110 and pi0228 n2545_not ; n2546
g111 and pi0137 n2521 ; n2547
g112 and n2446 n2547_not ; n2548
g113 and pi0332_not n2512 ; n2549
g114 nor pi0137 pi0153 ; n2550
g115 and n2549 n2550 ; n2551
g116 nor pi0228 n2548 ; n2552
g117 and n2551_not n2552 ; n2553
g118 nor n2546 n2553 ; n2554
g119 nor pi0216 n2554 ; n2555
g120 nor n2440 n2555 ; n2556
g121 nor pi0221 n2556 ; n2557
g122 nor n2457 n2557 ; n2558
g123 nor pi0215 n2558 ; n2559
g124 nor n2438 n2559 ; n2560
g125 and n2537 n2560 ; n2561
g126 nor n2542 n2561 ; n2562
g127 nor pi0056 n2562 ; n2563
g128 and pi0056 n2460 ; n2564
g129 and pi0062 n2564_not ; n2565
g130 and n2563_not n2565 ; n2566
g131 and pi0056 n2562_not ; n2567
g132 nor pi0087 pi0100 ; n2568
g133 nor pi0075 pi0092 ; n2569
g134 and n2532 n2569 ; n2570
g135 and n2568 n2570 ; n2571
g136 and n2530 n2571 ; n2572
g137 and n2460 n2572_not ; n2573
g138 and pi0228 n2543_not ; n2574
g139 and pi0332_not n2523 ; n2575
g140 and pi0105 n2575_not ; n2576
g141 and n2574 n2576_not ; n2577
g142 and pi0228_not n2446 ; n2578
g143 and n2521_not n2578 ; n2579
g144 nor pi0216 n2579 ; n2580
g145 and n2577_not n2580 ; n2581
g146 nor n2440 n2581 ; n2582
g147 nor pi0221 n2582 ; n2583
g148 nor n2457 n2583 ; n2584
g149 nor pi0215 n2584 ; n2585
g150 and n2438_not n2572 ; n2586
g151 and n2585_not n2586 ; n2587
g152 and pi0055 n2573_not ; n2588
g153 and n2587_not n2588 ; n2589
g154 and pi0299 n2460 ; n2590
g155 and pi0224_not pi0833 ; n2591
g156 and pi0222 n2591_not ; n2592
g157 nor pi0223 n2592 ; n2593
g158 and n2437 n2593_not ; n2594
g159 and pi0224 n2439_not ; n2595
g160 nor pi0222 n2595 ; n2596
g161 nor pi0332 pi0929 ; n2597
g162 and n2591 n2597 ; n2598
g163 nor n2596 n2598 ; n2599
g164 nor pi0223 n2599 ; n2600
g165 nor n2594 n2600 ; n2601
g166 nor pi0299 n2601 ; n2602
g167 nor pi0222 pi0224 ; n2603
g168 and pi0223_not n2603 ; n2604
g169 and n2444_not n2604 ; n2605
g170 and n2602 n2605_not ; n2606
g171 nor n2590 n2606 ; n2607
g172 nor pi0038 pi0100 ; n2608
g173 nor pi0039 pi0087 ; n2609
g174 and n2608 n2609 ; n2610
g175 and n2569 n2610 ; n2611
g176 and n2607 n2611_not ; n2612
g177 and n2525_not n2604 ; n2613
g178 nor n2601 n2613 ; n2614
g179 nor pi0299 n2614 ; n2615
g180 and n2460 n2528_not ; n2616
g181 and pi0299 n2616_not ; n2617
g182 nor n2615 n2617 ; n2618
g183 nor pi0039 n2618 ; n2619
g184 and pi0038_not n2568 ; n2620
g185 and n2569 n2620 ; n2621
g186 and n2619 n2621 ; n2622
g187 nor n2612 n2622 ; n2623
g188 and pi0054 n2623 ; n2624
g189 and pi0039_not n2608 ; n2625
g190 nor n2607 n2625 ; n2626
g191 and pi0299 n2560_not ; n2627
g192 nor n2615 n2627 ; n2628
g193 and n2625 n2628 ; n2629
g194 nor n2626 n2629 ; n2630
g195 and n2533 n2630_not ; n2631
g196 nor n2533 n2607 ; n2632
g197 and pi0092 n2632_not ; n2633
g198 and n2631_not n2633 ; n2634
g199 and pi0087 n2630_not ; n2635
g200 nor n2530 n2607 ; n2636
g201 and pi0095 pi0234 ; n2637
g202 nor pi0152 pi0161 ; n2638
g203 and pi0166_not n2638 ; n2639
g204 nor pi0146 n2639 ; n2640
g205 nor pi0210 n2640 ; n2641
g206 nor pi0137 n2637 ; n2642
g207 and n2641_not n2642 ; n2643
g208 nor n2523 n2643 ; n2644
g209 nor pi0332 n2644 ; n2645
g210 and pi0105 n2645_not ; n2646
g211 and n2574 n2646_not ; n2647
g212 and n2547 n2640 ; n2648
g213 and pi0137_not pi0210 ; n2649
g214 nor pi0252 n2649 ; n2650
g215 and n2640_not n2650 ; n2651
g216 and n2549 n2651 ; n2652
g217 and n2446 n2648_not ; n2653
g218 and n2652_not n2653 ; n2654
g219 and pi0252 n2640_not ; n2655
g220 nor n2641 n2655 ; n2656
g221 and n2551 n2656 ; n2657
g222 nor n2654 n2657 ; n2658
g223 nor pi0228 n2658 ; n2659
g224 nor pi0216 n2659 ; n2660
g225 and n2647_not n2660 ; n2661
g226 nor n2440 n2661 ; n2662
g227 nor pi0221 n2662 ; n2663
g228 nor n2457 n2663 ; n2664
g229 nor pi0215 n2664 ; n2665
g230 nor n2438 n2665 ; n2666
g231 and pi0299 n2666_not ; n2667
g232 nor pi0144 pi0174 ; n2668
g233 and pi0189_not n2668 ; n2669
g234 nor pi0223 n2669 ; n2670
g235 and pi0142 pi0198_not ; n2671
g236 nor pi0137 n2671 ; n2672
g237 nor n2523 n2672 ; n2673
g238 and n2444 n2673_not ; n2674
g239 and n2670 n2674_not ; n2675
g240 nor pi0234 pi0332 ; n2676
g241 and pi0137_not pi0198 ; n2677
g242 and n2521 n2677_not ; n2678
g243 and n2676 n2678_not ; n2679
g244 and pi0223_not n2669 ; n2680
g245 and pi0234 pi0332_not ; n2681
g246 and pi0095_not n2677 ; n2682
g247 nor n2513 n2682 ; n2683
g248 and n2681 n2683_not ; n2684
g249 and n2679_not n2680 ; n2685
g250 and n2684_not n2685 ; n2686
g251 nor n2675 n2686 ; n2687
g252 and n2603 n2687_not ; n2688
g253 nor n2601 n2688 ; n2689
g254 nor pi0299 n2689 ; n2690
g255 and n2530 n2690_not ; n2691
g256 and n2667_not n2691 ; n2692
g257 and pi0100 n2636_not ; n2693
g258 and n2692_not n2693 ; n2694
g259 and pi0039 n2607 ; n2695
g260 and pi0038 n2695_not ; n2696
g261 and n2619_not n2696 ; n2697
g262 and pi0039 n2628_not ; n2698
g263 and n2491 n2499 ; n2699
g264 nor pi0058 pi0091 ; n2700
g265 and pi0047_not n2700 ; n2701
g266 and n2493 n2701 ; n2702
g267 and n2699 n2702 ; n2703
g268 nor pi0090 pi0093 ; n2704
g269 nor pi0070 pi0096 ; n2705
g270 nor pi0035 pi0051 ; n2706
g271 and n2705 n2706 ; n2707
g272 and n2704 n2707 ; n2708
g273 and n2703 n2708 ; n2709
g274 and n2517 n2709 ; n2710
g275 and pi0225 n2710 ; n2711
g276 and pi0032 n2711_not ; n2712
g277 nor pi0095 n2712 ; n2713
g278 and pi0046_not n2493 ; n2714
g279 and n2492 n2496 ; n2715
g280 and n2714 n2715 ; n2716
g281 and pi0058_not n2716 ; n2717
g282 and pi0060 n2491 ; n2718
g283 nor pi0053 n2718 ; n2719
g284 nor pi0086 pi0094 ; n2720
g285 and pi0060_not n2491 ; n2721
g286 and pi0053 n2721_not ; n2722
g287 and n2720 n2722_not ; n2723
g288 and n2719_not n2723 ; n2724
g289 and n2704 n2717 ; n2725
g290 and n2724 n2725 ; n2726
g291 nor pi0035 n2726 ; n2727
g292 and pi0093_not n2503 ; n2728
g293 and pi0035 n2728_not ; n2729
g294 and pi0035 n2728 ; n2730
g295 and pi0225_not n2730 ; n2731
g296 nor pi0070 n2731 ; n2732
g297 and pi0051_not n2732 ; n2733
g298 and n2729_not n2733 ; n2734
g299 and n2727_not n2734 ; n2735
g300 and pi0040_not n2506 ; n2736
g301 and n2735 n2736 ; n2737
g302 nor pi0032 n2737 ; n2738
g303 and n2713 n2738_not ; n2739
g304 nor pi0137 n2739 ; n2740
g305 and pi0095 n2511_not ; n2741
g306 nor n2442 n2741 ; n2742
g307 and pi0040 n2509 ; n2743
g308 nor pi0032 n2743 ; n2744
g309 and pi0072 n2709_not ; n2745
g310 nor pi0040 n2745 ; n2746
g311 and pi0051 n2515_not ; n2747
g312 nor pi0096 n2747 ; n2748
g313 and pi0051_not pi0070 ; n2749
g314 and n2748 n2749_not ; n2750
g315 nor n2729 n2731 ; n2751
g316 and pi0093 n2503 ; n2752
g317 nor pi0035 n2752 ; n2753
g318 and pi0047_not n2500 ; n2754
g319 and n2491 n2754 ; n2755
g320 and pi0091 n2755 ; n2756
g321 and n2461 n2756_not ; n2757
g322 and pi0109_not n2699 ; n2758
g323 and pi0110 n2758_not ; n2759
g324 and pi0047 n2491 ; n2760
g325 and n2500 n2760 ; n2761
g326 and pi0047 n2761_not ; n2762
g327 nor pi0091 n2762 ; n2763
g328 and n2759_not n2763 ; n2764
g329 nor pi0047 pi0110 ; n2765
g330 and pi0109 n2699_not ; n2766
g331 and pi0102_not n2490 ; n2767
g332 and n2462 n2767 ; n2768
g333 and pi0050_not n2494 ; n2769
g334 and pi0077_not n2769 ; n2770
g335 and n2720 n2770 ; n2771
g336 and n2768 n2771 ; n2772
g337 and pi0097_not n2772 ; n2773
g338 and pi0108 n2773_not ; n2774
g339 nor pi0046 n2774 ; n2775
g340 and pi0097 n2772_not ; n2776
g341 and n2463 n2767 ; n2777
g342 and n2769 n2777 ; n2778
g343 and pi0086_not pi0094 ; n2779
g344 and n2778 n2779 ; n2780
g345 nor pi0097 n2780 ; n2781
g346 and pi0086 n2778_not ; n2782
g347 nor pi0094 n2782 ; n2783
g348 and pi0077 n2768 ; n2784
g349 nor pi0050 n2784 ; n2785
g350 and pi0081 n2489_not ; n2786
g351 and pi0102 n2490_not ; n2787
g352 nor n2786 n2787 ; n2788
g353 and pi0064 n2488_not ; n2789
g354 and pi0071 n2485_not ; n2790
g355 nor pi0065 n2790 ; n2791
g356 and pi0067_not n2483 ; n2792
g357 and pi0069 n2792_not ; n2793
g358 and pi0083 n2484_not ; n2794
g359 nor pi0103 n2794 ; n2795
g360 and n2793_not n2795 ; n2796
g361 nor pi0069 pi0083 ; n2797
g362 and pi0067 n2483_not ; n2798
g363 and n2469 n2477 ; n2799
g364 and pi0084_not n2799 ; n2800
g365 and pi0068_not n2800 ; n2801
g366 and n2479 n2801 ; n2802
g367 and pi0036 n2802_not ; n2803
g368 nor pi0036 pi0067 ; n2804
g369 nor pi0068 pi0111 ; n2805
g370 and pi0082 n2805 ; n2806
g371 and n2800 n2806 ; n2807
g372 and pi0111 n2801_not ; n2808
g373 nor pi0082 n2808 ; n2809
g374 and pi0068 n2800_not ; n2810
g375 and pi0084 n2799_not ; n2811
g376 and pi0104 n2475_not ; n2812
g377 and pi0085 pi0106 ; n2813
g378 and n2470 n2813_not ; n2814
g379 and pi0061 pi0076 ; n2815
g380 and n2471 n2815_not ; n2816
g381 nor n2814 n2816 ; n2817
g382 nor pi0048 n2817 ; n2818
g383 nor n2472 n2818 ; n2819
g384 and pi0089 n2473_not ; n2820
g385 nor pi0049 n2820 ; n2821
g386 and n2819_not n2821 ; n2822
g387 nor n2474 n2822 ; n2823
g388 nor pi0045 n2812 ; n2824
g389 and n2823_not n2824 ; n2825
g390 nor n2476 n2825 ; n2826
g391 nor n2477 n2826 ; n2827
g392 and n2469 n2827_not ; n2828
g393 and pi0066 pi0073 ; n2829
g394 nor n2469 n2477 ; n2830
g395 nor n2829 n2830 ; n2831
g396 and n2828_not n2831 ; n2832
g397 nor pi0084 n2832 ; n2833
g398 nor n2811 n2833 ; n2834
g399 and n2805 n2834_not ; n2835
g400 and n2809 n2810_not ; n2836
g401 and n2835_not n2836 ; n2837
g402 and n2804 n2807_not ; n2838
g403 and n2837_not n2838 ; n2839
g404 nor n2798 n2803 ; n2840
g405 and n2839_not n2840 ; n2841
g406 and n2797 n2841_not ; n2842
g407 and n2796 n2842_not ; n2843
g408 and pi0103 n2797 ; n2844
g409 and n2792 n2844 ; n2845
g410 nor pi0071 n2845 ; n2846
g411 and n2843_not n2846 ; n2847
g412 and n2791 n2847_not ; n2848
g413 nor pi0107 n2848 ; n2849
g414 and pi0065 pi0071_not ; n2850
g415 and n2485 n2850 ; n2851
g416 and n2849 n2851_not ; n2852
g417 and pi0107 n2486_not ; n2853
g418 nor pi0063 n2853 ; n2854
g419 and n2852_not n2854 ; n2855
g420 nor pi0064 n2855 ; n2856
g421 nor n2789 n2856 ; n2857
g422 nor pi0081 pi0102 ; n2858
g423 and n2857_not n2858 ; n2859
g424 and n2849_not n2854 ; n2860
g425 and pi0063 pi0107_not ; n2861
g426 and n2486 n2861 ; n2862
g427 nor pi0064 n2862 ; n2863
g428 and n2860_not n2863 ; n2864
g429 nor n2789 n2864 ; n2865
g430 and n2859 n2865_not ; n2866
g431 and n2788 n2866_not ; n2867
g432 and n2462 n2867_not ; n2868
g433 and pi0098 n2767_not ; n2869
g434 and pi0098_not n2767 ; n2870
g435 and pi0088 n2870_not ; n2871
g436 nor pi0077 n2869 ; n2872
g437 and n2871_not n2872 ; n2873
g438 and n2868_not n2873 ; n2874
g439 and n2785 n2874_not ; n2875
g440 and pi0050 n2777_not ; n2876
g441 nor pi0060 n2876 ; n2877
g442 and n2875_not n2877 ; n2878
g443 and n2719 n2878_not ; n2879
g444 nor n2722 n2879 ; n2880
g445 nor pi0086 n2880 ; n2881
g446 and n2783 n2881_not ; n2882
g447 and n2781 n2882_not ; n2883
g448 nor n2776 n2883 ; n2884
g449 nor pi0108 n2884 ; n2885
g450 and n2775 n2885_not ; n2886
g451 and pi0046 n2496 ; n2887
g452 and n2772 n2887 ; n2888
g453 nor pi0109 n2888 ; n2889
g454 and n2886_not n2889 ; n2890
g455 nor n2766 n2890 ; n2891
g456 and n2765 n2891_not ; n2892
g457 and n2764 n2892_not ; n2893
g458 and n2757 n2893_not ; n2894
g459 and pi0058 n2502_not ; n2895
g460 and pi0090 n2703_not ; n2896
g461 nor pi0093 n2896 ; n2897
g462 and n2895_not n2897 ; n2898
g463 and n2894_not n2898 ; n2899
g464 and n2753 n2899_not ; n2900
g465 and n2751 n2900_not ; n2901
g466 nor pi0051 n2901 ; n2902
g467 and n2750 n2902_not ; n2903
g468 nor pi0072 n2903 ; n2904
g469 and n2746 n2904_not ; n2905
g470 and n2744 n2905_not ; n2906
g471 nor n2712 n2906 ; n2907
g472 nor pi0095 n2907 ; n2908
g473 and n2742 n2908_not ; n2909
g474 and pi0137 n2909_not ; n2910
g475 nor n2740 n2910 ; n2911
g476 and pi0210 n2911_not ; n2912
g477 nor pi0051 pi0072 ; n2913
g478 and pi0841 n2503 ; n2914
g479 and pi0093_not n2914 ; n2915
g480 and n2913 n2915 ; n2916
g481 nor pi0035 pi0040 ; n2917
g482 and pi0225 n2917 ; n2918
g483 and n2705 n2918 ; n2919
g484 and n2916 n2919 ; n2920
g485 and pi0032 n2920_not ; n2921
g486 nor pi0095 n2921 ; n2922
g487 and pi0833_not pi0957 ; n2923
g488 and pi1091 n2923_not ; n2924
g489 and pi0829 pi0950 ; n2925
g490 and pi1092 pi1093 ; n2926
g491 and n2925 n2926 ; n2927
g492 and n2924 n2927 ; n2928
g493 nor n2727 n2928 ; n2929
g494 and pi1091 pi1093 ; n2930
g495 and n2923_not n2930 ; n2931
g496 and pi0950 pi1092 ; n2932
g497 and pi0829 n2932 ; n2933
g498 nor pi0046 pi0109 ; n2934
g499 and n2492 n2934 ; n2935
g500 nor pi0108 n2776 ; n2936
g501 and pi0110_not n2936 ; n2937
g502 and pi0093_not n2461 ; n2938
g503 nor pi0097 n2724 ; n2939
g504 and n2935 n2938 ; n2940
g505 and n2937 n2940 ; n2941
g506 and n2939_not n2941 ; n2942
g507 nor pi0035 n2942 ; n2943
g508 and n2931 n2933 ; n2944
g509 and n2943_not n2944 ; n2945
g510 nor n2929 n2945 ; n2946
g511 and n2734 n2736 ; n2947
g512 and n2946_not n2947 ; n2948
g513 nor pi0032 n2948 ; n2949
g514 and n2922 n2949_not ; n2950
g515 nor pi0137 n2950 ; n2951
g516 nor n2906 n2921 ; n2952
g517 nor pi0095 n2952 ; n2953
g518 and n2742 n2953_not ; n2954
g519 and pi0137 n2954_not ; n2955
g520 nor n2951 n2955 ; n2956
g521 nor pi0210 n2956 ; n2957
g522 nor n2912 n2957 ; n2958
g523 and pi0234_not n2958 ; n2959
g524 nor pi0096 n2735 ; n2960
g525 nor pi0035 pi0070 ; n2961
g526 and pi0051_not n2961 ; n2962
g527 and pi0091_not n2938 ; n2963
g528 and n2962 n2963 ; n2964
g529 and n2755 n2964 ; n2965
g530 and pi0096 n2965_not ; n2966
g531 and n2517 n2966_not ; n2967
g532 and n2960_not n2967 ; n2968
g533 nor pi0032 n2968 ; n2969
g534 and n2713 n2969_not ; n2970
g535 nor n2442 n2970 ; n2971
g536 and pi0137_not n2971 ; n2972
g537 and pi0096 n2965 ; n2973
g538 and pi0040_not n2913 ; n2974
g539 and n2505 n2974 ; n2975
g540 and n2973 n2975 ; n2976
g541 and n2906 n2976_not ; n2977
g542 nor n2712 n2977 ; n2978
g543 nor pi0095 n2978 ; n2979
g544 and pi0479 n2741 ; n2980
g545 nor n2979 n2980 ; n2981
g546 and pi0137 n2981_not ; n2982
g547 nor n2972 n2982 ; n2983
g548 and pi0210 n2983_not ; n2984
g549 nor n2921 n2977 ; n2985
g550 nor pi0095 n2985 ; n2986
g551 nor n2980 n2986 ; n2987
g552 and pi0137 n2987_not ; n2988
g553 and pi0095 pi0479 ; n2989
g554 nor n2921 n2969 ; n2990
g555 nor pi0095 n2990 ; n2991
g556 nor n2989 n2991 ; n2992
g557 nor pi0137 n2992 ; n2993
g558 nor n2988 n2993 ; n2994
g559 and n2924_not n2994 ; n2995
g560 and n2734 n2943_not ; n2996
g561 nor pi0096 n2996 ; n2997
g562 and n2967 n2997_not ; n2998
g563 nor pi0032 n2998 ; n2999
g564 nor n2921 n2999 ; n3000
g565 nor pi0095 n3000 ; n3001
g566 and n2927 n2989_not ; n3002
g567 and n3001_not n3002 ; n3003
g568 and n2927_not n2992 ; n3004
g569 nor pi0137 n3003 ; n3005
g570 and n3004_not n3005 ; n3006
g571 and n2924 n3006_not ; n3007
g572 and n2988_not n3007 ; n3008
g573 nor n2995 n3008 ; n3009
g574 and pi0210_not n3009 ; n3010
g575 nor n2984 n3010 ; n3011
g576 and pi0234 n3011 ; n3012
g577 nor pi0332 n2959 ; n3013
g578 and n3012_not n3013 ; n3014
g579 and n2639 n3014_not ; n3015
g580 and pi0146 n3011 ; n3016
g581 nor pi0210 n2994 ; n3017
g582 nor pi0146 n2984 ; n3018
g583 and n3017_not n3018 ; n3019
g584 and n2681 n3019_not ; n3020
g585 and n3016_not n3020 ; n3021
g586 and pi0146 n2958 ; n3022
g587 and n2738_not n2922 ; n3023
g588 nor pi0137 n3023 ; n3024
g589 nor n2955 n3024 ; n3025
g590 nor pi0210 n3025 ; n3026
g591 nor pi0146 n2912 ; n3027
g592 and n3026_not n3027 ; n3028
g593 and n2676 n3022_not ; n3029
g594 and n3028_not n3029 ; n3030
g595 nor n2639 n3030 ; n3031
g596 and n3021_not n3031 ; n3032
g597 nor n3015 n3032 ; n3033
g598 and pi0105 n3033_not ; n3034
g599 nor n2543 n3034 ; n3035
g600 and pi0228 n3035_not ; n3036
g601 nor pi0109 n2886 ; n3037
g602 nor n2766 n3037 ; n3038
g603 and n2765 n3038_not ; n3039
g604 and n2764 n3039_not ; n3040
g605 and n2757 n3040_not ; n3041
g606 and n2898 n3041_not ; n3042
g607 and n2753 n3042_not ; n3043
g608 and n2751 n3043_not ; n3044
g609 nor pi0051 n3044 ; n3045
g610 and n2750 n3045_not ; n3046
g611 nor pi0072 n3046 ; n3047
g612 and n2746 n3047_not ; n3048
g613 and n2744 n3048_not ; n3049
g614 nor n2921 n3049 ; n3050
g615 nor pi0095 n3050 ; n3051
g616 and n2742 n3051_not ; n3052
g617 and pi0137 n3052_not ; n3053
g618 and n2640 n3024 ; n3054
g619 and n2640_not n2951 ; n3055
g620 nor pi0210 pi0234 ; n3056
g621 and n3054_not n3056 ; n3057
g622 and n3055_not n3057 ; n3058
g623 and n3053_not n3058 ; n3059
g624 nor n2712 n3049 ; n3060
g625 nor pi0095 n3060 ; n3061
g626 and n2742 n3061_not ; n3062
g627 and pi0137 n3062_not ; n3063
g628 and pi0210 n2740_not ; n3064
g629 and n3063_not n3064 ; n3065
g630 and n2976_not n3049 ; n3066
g631 nor n2921 n3066 ; n3067
g632 nor pi0095 n3067 ; n3068
g633 nor n2741 n3068 ; n3069
g634 and pi0137 n3069_not ; n3070
g635 and n2640_not n2924 ; n3071
g636 and n3004_not n3071 ; n3072
g637 and n2741_not n2992 ; n3073
g638 and n3072_not n3073 ; n3074
g639 and n2741_not n3071 ; n3075
g640 and n3003 n3075 ; n3076
g641 nor pi0137 n3076 ; n3077
g642 and n3074_not n3077 ; n3078
g643 nor n3070 n3078 ; n3079
g644 nor pi0210 n3079 ; n3080
g645 and pi0234 n3080_not ; n3081
g646 nor n3059 n3065 ; n3082
g647 and n3081_not n3082 ; n3083
g648 nor pi0137 n2741 ; n3084
g649 and n2971_not n3084 ; n3085
g650 nor n2712 n3066 ; n3086
g651 nor pi0095 n3086 ; n3087
g652 and pi0137 n2741_not ; n3088
g653 and n3087_not n3088 ; n3089
g654 and pi0210 pi0234 ; n3090
g655 and n3085_not n3090 ; n3091
g656 and n3089_not n3091 ; n3092
g657 nor n3083 n3092 ; n3093
g658 and n2446 n3093_not ; n3094
g659 and pi0225 pi0841 ; n3095
g660 and n2710 n3095_not ; n3096
g661 and pi0032 n3096_not ; n3097
g662 nor pi0095 n3097 ; n3098
g663 and pi0070 n2505_not ; n3099
g664 and n2516 n3099_not ; n3100
g665 and n2517 n3100 ; n3101
g666 and n2732_not n3101 ; n3102
g667 nor pi0032 n3102 ; n3103
g668 and n3098 n3103_not ; n3104
g669 and pi0137 n3104_not ; n3105
g670 and pi0093 n2503_not ; n3106
g671 nor pi0035 n3106 ; n3107
g672 nor n2895 n2896 ; n3108
g673 and pi0053_not n2878 ; n3109
g674 nor pi0086 n3109 ; n3110
g675 and n2783 n3110_not ; n3111
g676 and n2781 n3111_not ; n3112
g677 nor n2776 n3112 ; n3113
g678 nor pi0108 n3113 ; n3114
g679 and n2775 n3114_not ; n3115
g680 nor pi0109 n3115 ; n3116
g681 nor n2766 n3116 ; n3117
g682 and n2765 n3117_not ; n3118
g683 and n2764 n3118_not ; n3119
g684 and n2757 n3119_not ; n3120
g685 and n3108 n3120_not ; n3121
g686 nor pi0093 n3121 ; n3122
g687 and n3107 n3122_not ; n3123
g688 and n2733 n3123_not ; n3124
g689 and n2748 n3099_not ; n3125
g690 and n3124_not n3125 ; n3126
g691 nor pi0072 n3126 ; n3127
g692 and n2746 n3127_not ; n3128
g693 and n2744 n3128_not ; n3129
g694 and n2928_not n3129 ; n3130
g695 and n2744 n2928 ; n3131
g696 nor pi0097 n3112 ; n3132
g697 nor pi0108 n3132 ; n3133
g698 and n2775 n3133_not ; n3134
g699 nor pi0109 n3134 ; n3135
g700 nor n2766 n3135 ; n3136
g701 and n2765 n3136_not ; n3137
g702 and n2764 n3137_not ; n3138
g703 and n2757 n3138_not ; n3139
g704 and n3108 n3139_not ; n3140
g705 nor pi0093 n3140 ; n3141
g706 and n3107 n3141_not ; n3142
g707 and n2733 n3142_not ; n3143
g708 and n3125 n3143_not ; n3144
g709 nor pi0072 n3144 ; n3145
g710 and n2746 n3145_not ; n3146
g711 and n3131 n3146_not ; n3147
g712 nor n3097 n3147 ; n3148
g713 and n3130_not n3148 ; n3149
g714 nor pi0095 n3149 ; n3150
g715 and n2742 n3150_not ; n3151
g716 nor pi0137 n3151 ; n3152
g717 nor n3105 n3152 ; n3153
g718 nor pi0210 n3153 ; n3154
g719 and pi0225_not n2710 ; n3155
g720 and pi0032 n3155_not ; n3156
g721 nor pi0095 n3156 ; n3157
g722 and pi0137 n3157 ; n3158
g723 and n3103_not n3158 ; n3159
g724 nor n3129 n3156 ; n3160
g725 nor pi0095 n3160 ; n3161
g726 and pi0137_not n2742 ; n3162
g727 and n3161_not n3162 ; n3163
g728 and pi0210 n3159_not ; n3164
g729 and n3163_not n3164 ; n3165
g730 and n2681 n3165_not ; n3166
g731 and n3154_not n3166 ; n3167
g732 nor pi0072 n2973 ; n3168
g733 and n3126_not n3168 ; n3169
g734 and n2746 n3169_not ; n3170
g735 and n2744 n3170_not ; n3171
g736 and n2928_not n3171 ; n3172
g737 and n3144_not n3168 ; n3173
g738 and n2746 n3173_not ; n3174
g739 and n3131 n3174_not ; n3175
g740 nor n3097 n3175 ; n3176
g741 and n3172_not n3176 ; n3177
g742 nor pi0095 n3177 ; n3178
g743 nor n2741 n3178 ; n3179
g744 nor pi0137 n3179 ; n3180
g745 and n2442 n2511 ; n3181
g746 and pi0072_not n2510 ; n3182
g747 and n2973 n3182 ; n3183
g748 and n3103 n3183_not ; n3184
g749 and n3098 n3184_not ; n3185
g750 and pi0137 n3181_not ; n3186
g751 and n3185_not n3186 ; n3187
g752 nor n3180 n3187 ; n3188
g753 nor pi0210 n3188 ; n3189
g754 nor n3156 n3171 ; n3190
g755 nor pi0095 n3190 ; n3191
g756 and n3084 n3191_not ; n3192
g757 and n3157 n3184_not ; n3193
g758 nor n3181 n3193 ; n3194
g759 and pi0137 n3194_not ; n3195
g760 and pi0210 n3195_not ; n3196
g761 and n3192_not n3196 ; n3197
g762 and n2676 n3197_not ; n3198
g763 and n3189_not n3198 ; n3199
g764 and n2639 n3167_not ; n3200
g765 and n3199_not n3200 ; n3201
g766 and pi0146 n3189 ; n3202
g767 nor pi0146 pi0210 ; n3203
g768 nor n3097 n3171 ; n3204
g769 nor pi0095 n3204 ; n3205
g770 nor n2741 n3205 ; n3206
g771 nor pi0137 n3206 ; n3207
g772 nor n3187 n3207 ; n3208
g773 and n3203 n3208_not ; n3209
g774 and n3198 n3209_not ; n3210
g775 and n3202_not n3210 ; n3211
g776 nor n3097 n3129 ; n3212
g777 nor pi0095 n3212 ; n3213
g778 and n2742 n3213_not ; n3214
g779 nor pi0137 n3214 ; n3215
g780 nor n3105 n3215 ; n3216
g781 and n3203 n3216_not ; n3217
g782 and pi0146 n3154 ; n3218
g783 and n3166 n3217_not ; n3219
g784 and n3218_not n3219 ; n3220
g785 nor n2639 n3211 ; n3221
g786 and n3220_not n3221 ; n3222
g787 nor pi0153 n3201 ; n3223
g788 and n3222_not n3223 ; n3224
g789 nor pi0228 n3094 ; n3225
g790 and n3224_not n3225 ; n3226
g791 nor n3036 n3226 ; n3227
g792 nor pi0216 n3227 ; n3228
g793 nor n2440 n3228 ; n3229
g794 nor pi0221 n3229 ; n3230
g795 nor n2457 n3230 ; n3231
g796 nor pi0215 n3231 ; n3232
g797 and pi0299 n2438_not ; n3233
g798 and n3232_not n3233 ; n3234
g799 and pi0198 n2983_not ; n3235
g800 and pi0198_not n3009 ; n3236
g801 nor n3235 n3236 ; n3237
g802 and pi0142 n3237 ; n3238
g803 nor pi0198 n2994 ; n3239
g804 nor pi0142 n3235 ; n3240
g805 and n3239_not n3240 ; n3241
g806 and n2681 n3241_not ; n3242
g807 and n3238_not n3242 ; n3243
g808 and pi0198 n2911_not ; n3244
g809 nor pi0198 n2956 ; n3245
g810 nor n3244 n3245 ; n3246
g811 and pi0142 n3246 ; n3247
g812 nor pi0198 n3025 ; n3248
g813 nor pi0142 n3244 ; n3249
g814 and n3248_not n3249 ; n3250
g815 and n2676 n3247_not ; n3251
g816 and n3250_not n3251 ; n3252
g817 and n2670 n3252_not ; n3253
g818 and n3243_not n3253 ; n3254
g819 and pi0234_not n3246 ; n3255
g820 and pi0234 n3237 ; n3256
g821 nor pi0332 n3255 ; n3257
g822 and n3256_not n3257 ; n3258
g823 and n2680 n3258_not ; n3259
g824 nor n3254 n3259 ; n3260
g825 and n2603 n3260_not ; n3261
g826 and n2602 n3261_not ; n3262
g827 nor pi0039 n3262 ; n3263
g828 and n3234_not n3263 ; n3264
g829 nor pi0038 n2698 ; n3265
g830 and n3264_not n3265 ; n3266
g831 nor pi0100 n2697 ; n3267
g832 and n3266_not n3267 ; n3268
g833 nor pi0087 n2694 ; n3269
g834 and n3268_not n3269 ; n3270
g835 nor pi0075 n2635 ; n3271
g836 and n3270_not n3271 ; n3272
g837 nor n2607 n2610 ; n3273
g838 and n2448 n2647_not ; n3274
g839 nor n2440 n3274 ; n3275
g840 nor pi0221 n3275 ; n3276
g841 nor n2457 n3276 ; n3277
g842 nor pi0215 n3277 ; n3278
g843 nor n2438 n3278 ; n3279
g844 and pi0299 n3279_not ; n3280
g845 and n2610 n2690_not ; n3281
g846 and n3280_not n3281 ; n3282
g847 and pi0075 n3273_not ; n3283
g848 and n3282_not n3283 ; n3284
g849 nor n3272 n3284 ; n3285
g850 nor pi0092 n3285 ; n3286
g851 nor pi0054 n2634 ; n3287
g852 and n3286_not n3287 ; n3288
g853 nor pi0074 n2624 ; n3289
g854 and n3288_not n3289 ; n3290
g855 and pi0054 n2607_not ; n3291
g856 and pi0054_not n2623 ; n3292
g857 and pi0074 n3291_not ; n3293
g858 and n3292_not n3293 ; n3294
g859 nor n3290 n3294 ; n3295
g860 nor pi0055 n3295 ; n3296
g861 nor pi0056 n2589 ; n3297
g862 and n3296_not n3297 ; n3298
g863 nor pi0062 n2567 ; n3299
g864 and n3298_not n3299 ; n3300
g865 nor pi0059 n2566 ; n3301
g866 and n3300_not n3301 ; n3302
g867 nor pi0057 n2541 ; n3303
g868 and n3302_not n3303 ; n3304
g869 and pi0059_not n2539 ; n3305
g870 and n2460 n3305_not ; n3306
g871 and pi0057 n3306_not ; n3307
g872 or n3304 n3307 ; po0153
g873 and pi0215 pi1146 ; n3309
g874 and pi0216 pi0221_not ; n3310
g875 and pi0276 n3310 ; n3311
g876 nor pi1146 n2452 ; n3312
g877 and pi0939_not n2452 ; n3313
g878 and pi0221 n3312_not ; n3314
g879 and n3313_not n3314 ; n3315
g880 nor n3311 n3315 ; n3316
g881 nor pi0215 n3316 ; n3317
g882 nor n3309 n3317 ; n3318
g883 and pi0154 n3318_not ; n3319
g884 nor pi0216 n2441 ; n3320
g885 nor n3311 n3320 ; n3321
g886 nor pi0221 n3321 ; n3322
g887 nor n3315 n3322 ; n3323
g888 nor pi0215 n3323 ; n3324
g889 nor n3309 n3324 ; n3325
g890 nor pi0154 n3325 ; n3326
g891 nor n3319 n3326 ; n3327
g892 nor pi0057 pi0059 ; n3328
g893 and n3327 n3328_not ; n3329
g894 and pi0056_not n2536 ; n3330
g895 and n2531 n3330 ; n3331
g896 nor n3327 n3331 ; n3332
g897 and pi0055_not n2572 ; n3333
g898 nor n3309 n3315 ; n3334
g899 and pi0228_not n2521 ; n3335
g900 and pi0216_not n3335 ; n3336
g901 and n3334 n3336 ; n3337
g902 and n3319_not n3337 ; n3338
g903 and n3327_not n3333 ; n3339
g904 and n3338_not n3339 ; n3340
g905 nor n3332 n3340 ; n3341
g906 and pi0062 n3341_not ; n3342
g907 nor n2537 n3327 ; n3343
g908 and pi0056 n3343_not ; n3344
g909 and n3340_not n3344 ; n3345
g910 and n2572 n3338 ; n3346
g911 and pi0055 n3327_not ; n3347
g912 and n3346_not n3347 ; n3348
g913 and pi0299 n3327_not ; n3349
g914 and pi0223 pi1146_not ; n3350
g915 and pi0222_not pi0224 ; n3351
g916 and pi0276 n3351 ; n3352
g917 nor pi1146 n2591 ; n3353
g918 and pi0939_not n2591 ; n3354
g919 and pi0222 n3353_not ; n3355
g920 and n3354_not n3355 ; n3356
g921 nor pi0223 n3352 ; n3357
g922 and n3356_not n3357 ; n3358
g923 nor pi0299 n3350 ; n3359
g924 and n3358_not n3359 ; n3360
g925 nor n3349 n3360 ; n3361
g926 and n2532_not n3361 ; n3362
g927 and pi0299 n3318_not ; n3363
g928 nor n3360 n3363 ; n3364
g929 and pi0154 n3364_not ; n3365
g930 and pi0299 n3325_not ; n3366
g931 and n3337_not n3366 ; n3367
g932 nor n3360 n3367 ; n3368
g933 nor pi0154 n3368 ; n3369
g934 and n2625 n3365_not ; n3370
g935 and n3369_not n3370 ; n3371
g936 and n2533 n3371 ; n3372
g937 and n2531 n2533 ; n3373
g938 and n3361 n3373_not ; n3374
g939 and pi0092 n3374_not ; n3375
g940 and n3372_not n3375 ; n3376
g941 and pi0075 n3361 ; n3377
g942 and n2625_not n3361 ; n3378
g943 nor n3371 n3378 ; n3379
g944 and pi0087 n3379_not ; n3380
g945 nor pi0038 pi0216 ; n3381
g946 and pi0228_not n3381 ; n3382
g947 and pi0154_not pi0299 ; n3383
g948 nor pi0146 n2521 ; n3384
g949 and pi0252_not n2521 ; n3385
g950 and pi0146 n3385_not ; n3386
g951 nor n3384 n3386 ; n3387
g952 and pi0152 n3387_not ; n3388
g953 nor pi0161 pi0166 ; n3389
g954 and n3385 n3389 ; n3390
g955 and n3387 n3389_not ; n3391
g956 nor pi0152 n3390 ; n3392
g957 and n3391_not n3392 ; n3393
g958 nor n3388 n3393 ; n3394
g959 and pi0039_not n3383 ; n3395
g960 and n3382 n3395 ; n3396
g961 and n3334 n3396 ; n3397
g962 and n3394 n3397 ; n3398
g963 and pi0100 n3361_not ; n3399
g964 and n3398_not n3399 ; n3400
g965 and pi0038 n3361 ; n3401
g966 and pi0039 n2521_not ; n3402
g967 and pi0070_not n3043 ; n3403
g968 nor n2729 n3099 ; n3404
g969 and n3403_not n3404 ; n3405
g970 nor pi0051 n3405 ; n3406
g971 and n2748 n3406_not ; n3407
g972 and n3168 n3407_not ; n3408
g973 nor n2745 n3408 ; n3409
g974 and n2510 n3409_not ; n3410
g975 and pi0040 n2509_not ; n3411
g976 and pi0032 n2710_not ; n3412
g977 nor n3411 n3412 ; n3413
g978 and n3410_not n3413 ; n3414
g979 nor pi0095 n3414 ; n3415
g980 nor n2741 n3415 ; n3416
g981 nor pi0039 n3416 ; n3417
g982 nor n3402 n3417 ; n3418
g983 nor pi0216 pi0228 ; n3419
g984 and n3334 n3419 ; n3420
g985 and n3418 n3420 ; n3421
g986 and n3366 n3421_not ; n3422
g987 nor n3360 n3422 ; n3423
g988 nor pi0154 n3423 ; n3424
g989 nor pi0038 n3365 ; n3425
g990 and n3424_not n3425 ; n3426
g991 nor pi0100 n3401 ; n3427
g992 and n3426_not n3427 ; n3428
g993 nor pi0087 n3400 ; n3429
g994 and n3428_not n3429 ; n3430
g995 nor n3380 n3430 ; n3431
g996 nor pi0075 n3431 ; n3432
g997 nor pi0092 n3377 ; n3433
g998 and n3432_not n3433 ; n3434
g999 and n2532 n3376_not ; n3435
g1000 and n3434_not n3435 ; n3436
g1001 nor pi0055 n3362 ; n3437
g1002 and n3436_not n3437 ; n3438
g1003 nor pi0056 n3348 ; n3439
g1004 and n3438_not n3439 ; n3440
g1005 nor pi0062 n3345 ; n3441
g1006 and n3440_not n3441 ; n3442
g1007 and n3328 n3342_not ; n3443
g1008 and n3442_not n3443 ; n3444
g1009 nor pi0239 n3329 ; n3445
g1010 and n3444_not n3445 ; n3446
g1011 and n2441 n2442 ; n3447
g1012 nor pi0216 pi0221 ; n3448
g1013 and pi0215_not n3448 ; n3449
g1014 and n3447 n3449 ; n3450
g1015 and n3318 n3450_not ; n3451
g1016 nor pi0215 n3451 ; n3452
g1017 and pi0154 n3451_not ; n3453
g1018 nor n3326 n3452 ; n3454
g1019 and n3453_not n3454 ; n3455
g1020 and n3328_not n3455 ; n3456
g1021 nor n3331 n3455 ; n3457
g1022 and n3337 n3453_not ; n3458
g1023 nor n3455 n3458 ; n3459
g1024 and n3333 n3459 ; n3460
g1025 and pi0056_not n3460 ; n3461
g1026 nor n3457 n3461 ; n3462
g1027 and pi0062 n3462_not ; n3463
g1028 nor n2537 n3455 ; n3464
g1029 and pi0056 n3464_not ; n3465
g1030 and n3460_not n3465 ; n3466
g1031 and n2572 n3458 ; n3467
g1032 and pi0055 n3455_not ; n3468
g1033 and n3467_not n3468 ; n3469
g1034 nor pi0223 pi0299 ; n3470
g1035 and n2603 n3470 ; n3471
g1036 and n2442 n3471 ; n3472
g1037 and pi0299 n3455_not ; n3473
g1038 nor n3360 n3472 ; n3474
g1039 and n3473_not n3474 ; n3475
g1040 and n2532_not n3475 ; n3476
g1041 and pi0299 n3459_not ; n3477
g1042 and n3373 n3477 ; n3478
g1043 and pi0092 n3475_not ; n3479
g1044 and n3478_not n3479 ; n3480
g1045 and pi0075 n3475 ; n3481
g1046 and n2625 n3477 ; n3482
g1047 and pi0087 n3475_not ; n3483
g1048 and n3482_not n3483 ; n3484
g1049 nor n3475 n3477 ; n3485
g1050 and pi0039 n3485_not ; n3486
g1051 and n2519 n2973 ; n3487
g1052 nor n2442 n3487 ; n3488
g1053 and pi0224_not n3488 ; n3489
g1054 and pi0224 pi0276_not ; n3490
g1055 nor pi0222 n3490 ; n3491
g1056 and n3489_not n3491 ; n3492
g1057 nor pi0223 n3356 ; n3493
g1058 and n3492_not n3493 ; n3494
g1059 nor n3350 n3494 ; n3495
g1060 nor pi0299 n3495 ; n3496
g1061 and pi0105 n3488_not ; n3497
g1062 and pi0228 n3497_not ; n3498
g1063 nor n2741 n3488 ; n3499
g1064 nor pi0228 n3499 ; n3500
g1065 nor n3498 n3500 ; n3501
g1066 and pi0154 n3501_not ; n3502
g1067 nor pi0072 n3407 ; n3503
g1068 nor n2745 n3503 ; n3504
g1069 and n2510 n3504_not ; n3505
g1070 and n3413 n3505_not ; n3506
g1071 nor pi0095 n3506 ; n3507
g1072 and n2742 n3507_not ; n3508
g1073 and pi0228_not n3508 ; n3509
g1074 and n2441 n3488 ; n3510
g1075 nor n3509 n3510 ; n3511
g1076 nor pi0154 n3511 ; n3512
g1077 and n3449 n3502_not ; n3513
g1078 and n3512_not n3513 ; n3514
g1079 and pi0299 n3318 ; n3515
g1080 and n3514_not n3515 ; n3516
g1081 nor n3496 n3516 ; n3517
g1082 nor pi0039 n3517 ; n3518
g1083 and n2608 n3486_not ; n3519
g1084 and n3518_not n3519 ; n3520
g1085 and pi0100 n3398 ; n3521
g1086 nor n2608 n3475 ; n3522
g1087 and n3521_not n3522 ; n3523
g1088 nor n3520 n3523 ; n3524
g1089 nor pi0087 n3524 ; n3525
g1090 nor pi0075 n3484 ; n3526
g1091 and n3525_not n3526 ; n3527
g1092 nor pi0092 n3481 ; n3528
g1093 and n3527_not n3528 ; n3529
g1094 and n2532 n3480_not ; n3530
g1095 and n3529_not n3530 ; n3531
g1096 nor pi0055 n3476 ; n3532
g1097 and n3531_not n3532 ; n3533
g1098 nor pi0056 n3469 ; n3534
g1099 and n3533_not n3534 ; n3535
g1100 nor pi0062 n3466 ; n3536
g1101 and n3535_not n3536 ; n3537
g1102 and n3328 n3463_not ; n3538
g1103 and n3537_not n3538 ; n3539
g1104 and pi0239 n3456_not ; n3540
g1105 and n3539_not n3540 ; n3541
g1106 or n3446 n3541 ; po0154
g1107 and pi0215 pi1145 ; n3543
g1108 and pi0216 pi0274 ; n3544
g1109 nor pi0221 n3544 ; n3545
g1110 nor pi0151 n2441 ; n3546
g1111 nor pi0216 n3546 ; n3547
g1112 and n3545 n3547_not ; n3548
g1113 nor pi1145 n2452 ; n3549
g1114 and pi0927_not n2452 ; n3550
g1115 and pi0221 n3549_not ; n3551
g1116 and n3550_not n3551 ; n3552
g1117 nor n3548 n3552 ; n3553
g1118 nor pi0215 n3553 ; n3554
g1119 nor n3543 n3554 ; n3555
g1120 and n2526 n3447 ; n3556
g1121 and n3544_not n3556 ; n3557
g1122 and n3555 n3557_not ; n3558
g1123 and n3331_not n3558 ; n3559
g1124 nor n3447 n3546 ; n3560
g1125 and pi0151_not n3335 ; n3561
g1126 nor n3560 n3561 ; n3562
g1127 nor pi0216 n3562 ; n3563
g1128 and n3545 n3563_not ; n3564
g1129 nor n3552 n3564 ; n3565
g1130 nor pi0215 n3565 ; n3566
g1131 nor n3543 n3566 ; n3567
g1132 and n3331 n3567 ; n3568
g1133 and pi0062 n3559_not ; n3569
g1134 and n3568_not n3569 ; n3570
g1135 nor n2537 n3558 ; n3571
g1136 and n2537 n3567_not ; n3572
g1137 and pi0056 n3571_not ; n3573
g1138 and n3572_not n3573 ; n3574
g1139 and n2572_not n3558 ; n3575
g1140 and n2572 n3567 ; n3576
g1141 and pi0055 n3575_not ; n3577
g1142 and n3576_not n3577 ; n3578
g1143 and pi0223 pi1145 ; n3579
g1144 nor pi1145 n2591 ; n3580
g1145 and pi0927_not n2591 ; n3581
g1146 and pi0222 n3580_not ; n3582
g1147 and n3581_not n3582 ; n3583
g1148 and pi0224 pi0274 ; n3584
g1149 and n3351 n3584_not ; n3585
g1150 nor n3583 n3585 ; n3586
g1151 nor pi0223 n3586 ; n3587
g1152 nor n3579 n3587 ; n3588
g1153 nor pi0299 n3588 ; n3589
g1154 nor n3472 n3589 ; n3590
g1155 and pi0299 n3558_not ; n3591
g1156 and n3590 n3591_not ; n3592
g1157 and n2532_not n3592 ; n3593
g1158 and n2625_not n3592 ; n3594
g1159 and pi0299 n3567_not ; n3595
g1160 and n3590 n3595_not ; n3596
g1161 and n2625 n3596 ; n3597
g1162 nor n3594 n3597 ; n3598
g1163 and n2533 n3598_not ; n3599
g1164 and n2533_not n3592 ; n3600
g1165 and pi0092 n3600_not ; n3601
g1166 and n3599_not n3601 ; n3602
g1167 and pi0075 n3592 ; n3603
g1168 and pi0087 n3598 ; n3604
g1169 and pi0038 n3592 ; n3605
g1170 and pi0039 n3596_not ; n3606
g1171 nor pi0222 n3584 ; n3607
g1172 and n3489_not n3607 ; n3608
g1173 nor n3583 n3608 ; n3609
g1174 nor pi0223 n3609 ; n3610
g1175 nor pi0299 n3579 ; n3611
g1176 and n3610_not n3611 ; n3612
g1177 and pi0151_not n3511 ; n3613
g1178 and pi0151 n3501 ; n3614
g1179 nor pi0216 n3614 ; n3615
g1180 and n3613_not n3615 ; n3616
g1181 and n3545 n3616_not ; n3617
g1182 nor n3552 n3617 ; n3618
g1183 nor pi0215 n3618 ; n3619
g1184 and pi0299 n3543_not ; n3620
g1185 and n3619_not n3620 ; n3621
g1186 nor pi0039 n3612 ; n3622
g1187 and n3621_not n3622 ; n3623
g1188 nor pi0038 n3606 ; n3624
g1189 and n3623_not n3624 ; n3625
g1190 nor pi0100 n3605 ; n3626
g1191 and n3625_not n3626 ; n3627
g1192 and n2530_not n3592 ; n3628
g1193 and pi0228_not n3394 ; n3629
g1194 and n2441 n2442_not ; n3630
g1195 nor n3629 n3630 ; n3631
g1196 and pi0151_not n3631 ; n3632
g1197 and n3563 n3632_not ; n3633
g1198 and n3545 n3633_not ; n3634
g1199 nor n3552 n3634 ; n3635
g1200 nor pi0215 n3635 ; n3636
g1201 nor n3543 n3636 ; n3637
g1202 and pi0299 n3637_not ; n3638
g1203 and n2530 n3590 ; n3639
g1204 and n3638_not n3639 ; n3640
g1205 and pi0100 n3628_not ; n3641
g1206 and n3640_not n3641 ; n3642
g1207 nor n3627 n3642 ; n3643
g1208 nor pi0087 n3643 ; n3644
g1209 nor pi0075 n3604 ; n3645
g1210 and n3644_not n3645 ; n3646
g1211 nor pi0092 n3603 ; n3647
g1212 and n3646_not n3647 ; n3648
g1213 and n2532 n3602_not ; n3649
g1214 and n3648_not n3649 ; n3650
g1215 nor pi0055 n3593 ; n3651
g1216 and n3650_not n3651 ; n3652
g1217 nor pi0056 n3578 ; n3653
g1218 and n3652_not n3653 ; n3654
g1219 nor pi0062 n3574 ; n3655
g1220 and n3654_not n3655 ; n3656
g1221 and pi0235 n3328 ; n3657
g1222 and n3570_not n3657 ; n3658
g1223 and n3656_not n3658 ; n3659
g1224 nor n3543 n3552 ; n3660
g1225 and n3336 n3660 ; n3661
g1226 and n2537 n3661 ; n3662
g1227 and pi0056_not n3662 ; n3663
g1228 and pi0062 n3555_not ; n3664
g1229 and n3663_not n3664 ; n3665
g1230 nor n3555 n3662 ; n3666
g1231 and pi0056 n3666_not ; n3667
g1232 and n2572 n3661 ; n3668
g1233 and pi0055 n3555_not ; n3669
g1234 and n3668_not n3669 ; n3670
g1235 and pi0299 n3555_not ; n3671
g1236 nor n3589 n3671 ; n3672
g1237 and n2532_not n3672 ; n3673
g1238 and n3661_not n3671 ; n3674
g1239 and n2531 n3589_not ; n3675
g1240 and n3674_not n3675 ; n3676
g1241 and n2533 n3676 ; n3677
g1242 and n3373_not n3672 ; n3678
g1243 and pi0092 n3678_not ; n3679
g1244 and n3677_not n3679 ; n3680
g1245 and pi0075 n3672 ; n3681
g1246 and n2625_not n3672 ; n3682
g1247 nor n3676 n3682 ; n3683
g1248 and pi0087 n3683_not ; n3684
g1249 and pi0100_not n3418 ; n3685
g1250 and pi0039_not pi0100 ; n3686
g1251 and n3394 n3686 ; n3687
g1252 nor n3685 n3687 ; n3688
g1253 and n3382 n3660 ; n3689
g1254 and n3688_not n3689 ; n3690
g1255 and n3671 n3690_not ; n3691
g1256 nor pi0087 n3589 ; n3692
g1257 and n3691_not n3692 ; n3693
g1258 nor n3684 n3693 ; n3694
g1259 nor pi0075 n3694 ; n3695
g1260 nor pi0092 n3681 ; n3696
g1261 and n3695_not n3696 ; n3697
g1262 and n2532 n3680_not ; n3698
g1263 and n3697_not n3698 ; n3699
g1264 nor pi0055 n3673 ; n3700
g1265 and n3699_not n3700 ; n3701
g1266 nor pi0056 n3670 ; n3702
g1267 and n3701_not n3702 ; n3703
g1268 nor pi0062 n3667 ; n3704
g1269 and n3703_not n3704 ; n3705
g1270 and pi0235_not n3328 ; n3706
g1271 and n3665_not n3706 ; n3707
g1272 and n3705_not n3707 ; n3708
g1273 and pi0235 n3557 ; n3709
g1274 nor n3328 n3709 ; n3710
g1275 and n3555 n3710 ; n3711
g1276 nor n3708 n3711 ; n3712
g1277 and n3659_not n3712 ; po0155
g1278 and pi0215 pi1143 ; n3714
g1279 and pi0216 pi0264 ; n3715
g1280 nor pi0221 n3715 ; n3716
g1281 and pi0105_not pi0146 ; n3717
g1282 and pi0284 n2442_not ; n3718
g1283 and pi0105 n3718_not ; n3719
g1284 and pi0228 n3717_not ; n3720
g1285 and n3719_not n3720 ; n3721
g1286 nor n3447 n3721 ; n3722
g1287 nor pi0146 pi0228 ; n3723
g1288 and n3722 n3723_not ; n3724
g1289 nor pi0216 n3724 ; n3725
g1290 and n3716 n3725_not ; n3726
g1291 nor pi1143 n2452 ; n3727
g1292 and pi0944_not n2452 ; n3728
g1293 and pi0221 n3727_not ; n3729
g1294 and n3728_not n3729 ; n3730
g1295 nor n3726 n3730 ; n3731
g1296 nor pi0215 n3731 ; n3732
g1297 nor n3714 n3732 ; n3733
g1298 and n3331_not n3733 ; n3734
g1299 and pi0284 n2521 ; n3735
g1300 nor n3384 n3735 ; n3736
g1301 nor pi0228 n3736 ; n3737
g1302 and n3722 n3737_not ; n3738
g1303 nor pi0216 n3738 ; n3739
g1304 and n3716 n3739_not ; n3740
g1305 nor n3730 n3740 ; n3741
g1306 nor pi0215 n3741 ; n3742
g1307 nor n3714 n3742 ; n3743
g1308 and n3331 n3743 ; n3744
g1309 and pi0062 n3734_not ; n3745
g1310 and n3744_not n3745 ; n3746
g1311 nor n2537 n3733 ; n3747
g1312 and n2537 n3743_not ; n3748
g1313 and pi0056 n3747_not ; n3749
g1314 and n3748_not n3749 ; n3750
g1315 and n2572_not n3733 ; n3751
g1316 and n2572 n3743 ; n3752
g1317 and pi0055 n3751_not ; n3753
g1318 and n3752_not n3753 ; n3754
g1319 and n2442 n2604 ; n3755
g1320 and pi0223 pi1143 ; n3756
g1321 and pi0224 pi0264 ; n3757
g1322 nor pi0222 n3757 ; n3758
g1323 and pi0224_not n3718 ; n3759
g1324 and n3758 n3759_not ; n3760
g1325 nor pi1143 n2591 ; n3761
g1326 and pi0944_not n2591 ; n3762
g1327 and pi0222 n3761_not ; n3763
g1328 and n3762_not n3763 ; n3764
g1329 nor n3760 n3764 ; n3765
g1330 nor pi0223 n3765 ; n3766
g1331 nor n3756 n3766 ; n3767
g1332 nor pi0299 n3767 ; n3768
g1333 and n3755_not n3768 ; n3769
g1334 and pi0299 n3733_not ; n3770
g1335 nor n3769 n3770 ; n3771
g1336 and n2532_not n3771 ; n3772
g1337 and n2625_not n3771 ; n3773
g1338 and pi0299 n3743_not ; n3774
g1339 nor n3769 n3774 ; n3775
g1340 and n2625 n3775 ; n3776
g1341 nor n3773 n3776 ; n3777
g1342 and n2533 n3777_not ; n3778
g1343 and n2533_not n3771 ; n3779
g1344 and pi0092 n3779_not ; n3780
g1345 and n3778_not n3780 ; n3781
g1346 and pi0075 n3771 ; n3782
g1347 and pi0087 n3777 ; n3783
g1348 and pi0038 n3771 ; n3784
g1349 and pi0039 n3775_not ; n3785
g1350 nor pi0299 n3756 ; n3786
g1351 and pi0284_not n3488 ; n3787
g1352 nor pi0224 n3787 ; n3788
g1353 and n3758 n3788_not ; n3789
g1354 nor n3764 n3789 ; n3790
g1355 and n3786 n3790 ; n3791
g1356 and pi0299 n3714_not ; n3792
g1357 and n2441 n3488_not ; n3793
g1358 nor pi0146 n3508 ; n3794
g1359 and pi0146 n3499 ; n3795
g1360 nor pi0284 n3795 ; n3796
g1361 and pi0146 pi0284 ; n3797
g1362 and n3416_not n3797 ; n3798
g1363 nor n3796 n3798 ; n3799
g1364 nor n3794 n3799 ; n3800
g1365 nor pi0228 n3800 ; n3801
g1366 nor n3721 n3793 ; n3802
g1367 and n3801_not n3802 ; n3803
g1368 nor pi0216 n3803 ; n3804
g1369 and n3716 n3804_not ; n3805
g1370 nor n3730 n3805 ; n3806
g1371 nor pi0215 n3806 ; n3807
g1372 and n3792 n3807_not ; n3808
g1373 and n3488_not n3758 ; n3809
g1374 and n3790 n3809_not ; n3810
g1375 nor pi0223 n3810 ; n3811
g1376 and n3786 n3811_not ; n3812
g1377 nor pi0039 n3812 ; n3813
g1378 and n3791_not n3813 ; n3814
g1379 and n3808_not n3814 ; n3815
g1380 nor pi0038 n3785 ; n3816
g1381 and n3815_not n3816 ; n3817
g1382 nor pi0100 n3784 ; n3818
g1383 and n3817_not n3818 ; n3819
g1384 and n2530_not n3771 ; n3820
g1385 and pi0252 n2639 ; n3821
g1386 nor pi0284 n3821 ; n3822
g1387 and n2521 n3822 ; n3823
g1388 nor pi0228 n3823 ; n3824
g1389 and n3386_not n3824 ; n3825
g1390 and n3722 n3825_not ; n3826
g1391 nor pi0216 n3826 ; n3827
g1392 and n3716 n3827_not ; n3828
g1393 nor n3730 n3828 ; n3829
g1394 nor pi0215 n3829 ; n3830
g1395 nor n3714 n3830 ; n3831
g1396 and pi0299 n3831_not ; n3832
g1397 and n2530 n3769_not ; n3833
g1398 and n3832_not n3833 ; n3834
g1399 and pi0100 n3820_not ; n3835
g1400 and n3834_not n3835 ; n3836
g1401 nor n3819 n3836 ; n3837
g1402 nor pi0087 n3837 ; n3838
g1403 nor pi0075 n3783 ; n3839
g1404 and n3838_not n3839 ; n3840
g1405 nor pi0092 n3782 ; n3841
g1406 and n3840_not n3841 ; n3842
g1407 and n2532 n3781_not ; n3843
g1408 and n3842_not n3843 ; n3844
g1409 nor pi0055 n3772 ; n3845
g1410 and n3844_not n3845 ; n3846
g1411 nor pi0056 n3754 ; n3847
g1412 and n3846_not n3847 ; n3848
g1413 nor pi0062 n3750 ; n3849
g1414 and n3848_not n3849 ; n3850
g1415 and pi0238_not n3328 ; n3851
g1416 and n3746_not n3851 ; n3852
g1417 and n3850_not n3852 ; n3853
g1418 nor n3721 n3737 ; n3854
g1419 nor pi0216 n3854 ; n3855
g1420 and n3716 n3855_not ; n3856
g1421 nor n3730 n3856 ; n3857
g1422 nor pi0215 n3857 ; n3858
g1423 nor n3714 n3858 ; n3859
g1424 and n3331 n3859 ; n3860
g1425 and n3556 n3715_not ; n3861
g1426 and n3733 n3861_not ; n3862
g1427 and n3331_not n3862 ; n3863
g1428 and pi0062 n3863_not ; n3864
g1429 and n3860_not n3864 ; n3865
g1430 nor n2537 n3862 ; n3866
g1431 and n2537 n3859_not ; n3867
g1432 and pi0056 n3866_not ; n3868
g1433 and n3867_not n3868 ; n3869
g1434 and n2572 n3859 ; n3870
g1435 and n2572_not n3862 ; n3871
g1436 and pi0055 n3871_not ; n3872
g1437 and n3870_not n3872 ; n3873
g1438 and pi0299 n3862_not ; n3874
g1439 nor n3768 n3874 ; n3875
g1440 and n2532_not n3875 ; n3876
g1441 and n2625_not n3875 ; n3877
g1442 and pi0299 n3859_not ; n3878
g1443 nor n3768 n3878 ; n3879
g1444 and n2625 n3879 ; n3880
g1445 nor n3877 n3880 ; n3881
g1446 and n2533 n3881_not ; n3882
g1447 and n2533_not n3875 ; n3883
g1448 and pi0092 n3883_not ; n3884
g1449 and n3882_not n3884 ; n3885
g1450 and pi0075 n3875 ; n3886
g1451 and pi0087 n3881 ; n3887
g1452 and pi0038 n3875 ; n3888
g1453 and pi0039 n3879_not ; n3889
g1454 and n3497_not n3721 ; n3890
g1455 and pi0146_not n3499 ; n3891
g1456 and pi0146 n3508_not ; n3892
g1457 and pi0284 n3891_not ; n3893
g1458 and n3892_not n3893 ; n3894
g1459 nor pi0146 pi0284 ; n3895
g1460 and n3416_not n3895 ; n3896
g1461 nor n3894 n3896 ; n3897
g1462 nor pi0228 n3897 ; n3898
g1463 nor n3890 n3898 ; n3899
g1464 nor pi0216 n3899 ; n3900
g1465 and n3716 n3900_not ; n3901
g1466 nor n3730 n3901 ; n3902
g1467 nor pi0215 n3902 ; n3903
g1468 and n3792 n3903_not ; n3904
g1469 and n3813 n3904_not ; n3905
g1470 nor pi0038 n3889 ; n3906
g1471 and n3905_not n3906 ; n3907
g1472 nor pi0100 n3888 ; n3908
g1473 and n3907_not n3908 ; n3909
g1474 and n2530_not n3875 ; n3910
g1475 nor n3721 n3825 ; n3911
g1476 nor pi0216 n3911 ; n3912
g1477 and n3716 n3912_not ; n3913
g1478 nor n3730 n3913 ; n3914
g1479 nor pi0215 n3914 ; n3915
g1480 nor n3714 n3915 ; n3916
g1481 and pi0299 n3916_not ; n3917
g1482 and n2530 n3768_not ; n3918
g1483 and n3917_not n3918 ; n3919
g1484 and pi0100 n3910_not ; n3920
g1485 and n3919_not n3920 ; n3921
g1486 nor n3909 n3921 ; n3922
g1487 nor pi0087 n3922 ; n3923
g1488 nor pi0075 n3887 ; n3924
g1489 and n3923_not n3924 ; n3925
g1490 nor pi0092 n3886 ; n3926
g1491 and n3925_not n3926 ; n3927
g1492 and n2532 n3885_not ; n3928
g1493 and n3927_not n3928 ; n3929
g1494 nor pi0055 n3876 ; n3930
g1495 and n3929_not n3930 ; n3931
g1496 nor pi0056 n3873 ; n3932
g1497 and n3931_not n3932 ; n3933
g1498 nor pi0062 n3869 ; n3934
g1499 and n3933_not n3934 ; n3935
g1500 and pi0238 n3328 ; n3936
g1501 and n3865_not n3936 ; n3937
g1502 and n3935_not n3937 ; n3938
g1503 and pi0238 n3861 ; n3939
g1504 nor n3328 n3939 ; n3940
g1505 and n3733 n3940 ; n3941
g1506 nor n3853 n3941 ; n3942
g1507 and n3938_not n3942 ; po0156
g1508 and pi0215 pi1142 ; n3944
g1509 and pi0216 pi0277 ; n3945
g1510 nor pi0221 n3945 ; n3946
g1511 and pi0172 pi0228_not ; n3947
g1512 and pi0105_not pi0172 ; n3948
g1513 and pi0262 n2442_not ; n3949
g1514 and pi0105 n3949 ; n3950
g1515 nor n3948 n3950 ; n3951
g1516 and pi0228 n3951_not ; n3952
g1517 nor n3947 n3952 ; n3953
g1518 nor pi0216 n3953 ; n3954
g1519 and n3946 n3954_not ; n3955
g1520 nor pi1142 n2452 ; n3956
g1521 and pi0932_not n2452 ; n3957
g1522 and pi0221 n3956_not ; n3958
g1523 and n3957_not n3958 ; n3959
g1524 nor n3955 n3959 ; n3960
g1525 nor pi0215 n3960 ; n3961
g1526 nor n3944 n3961 ; n3962
g1527 nor n3450 n3962 ; n3963
g1528 nor n3328 n3963 ; n3964
g1529 nor n3331 n3963 ; n3965
g1530 and pi0262_not n2521 ; n3966
g1531 nor n3335 n3947 ; n3967
g1532 nor n3966 n3967 ; n3968
g1533 nor n3447 n3952 ; n3969
g1534 and n3968_not n3969 ; n3970
g1535 nor pi0216 n3970 ; n3971
g1536 and n3946 n3971_not ; n3972
g1537 nor n3959 n3972 ; n3973
g1538 nor pi0215 n3973 ; n3974
g1539 nor n3944 n3974 ; n3975
g1540 and n3331 n3975 ; n3976
g1541 and pi0062 n3965_not ; n3977
g1542 and n3976_not n3977 ; n3978
g1543 and n2537 n3975_not ; n3979
g1544 and n2537_not n3963 ; n3980
g1545 and pi0056 n3980_not ; n3981
g1546 and n3979_not n3981 ; n3982
g1547 nor n2572 n3963 ; n3983
g1548 and n2572 n3975 ; n3984
g1549 and pi0055 n3983_not ; n3985
g1550 and n3984_not n3985 ; n3986
g1551 and pi0223 pi1142 ; n3987
g1552 and pi0224 pi0277 ; n3988
g1553 nor pi0222 n3988 ; n3989
g1554 and pi0224_not n3949 ; n3990
g1555 and n3989 n3990_not ; n3991
g1556 nor pi1142 n2591 ; n3992
g1557 and pi0932_not n2591 ; n3993
g1558 and pi0222 n3992_not ; n3994
g1559 and n3993_not n3994 ; n3995
g1560 nor n3991 n3995 ; n3996
g1561 nor pi0223 n3996 ; n3997
g1562 nor n3987 n3997 ; n3998
g1563 nor pi0299 n3998 ; n3999
g1564 and n3755_not n3999 ; n4000
g1565 and pi0299 n3963 ; n4001
g1566 nor n4000 n4001 ; n4002
g1567 and n2532_not n4002 ; n4003
g1568 and n2625_not n4002 ; n4004
g1569 and pi0299 n3975_not ; n4005
g1570 nor n4000 n4005 ; n4006
g1571 and n2625 n4006 ; n4007
g1572 nor n4004 n4007 ; n4008
g1573 and n2533 n4008_not ; n4009
g1574 and n2533_not n4002 ; n4010
g1575 and pi0092 n4010_not ; n4011
g1576 and n4009_not n4011 ; n4012
g1577 and pi0075 n4002 ; n4013
g1578 and pi0087 n4008 ; n4014
g1579 and pi0038 n4002 ; n4015
g1580 and pi0039 n4006_not ; n4016
g1581 nor pi0299 n3987 ; n4017
g1582 and pi0262_not n3488 ; n4018
g1583 nor pi0224 n4018 ; n4019
g1584 and n3989 n4019_not ; n4020
g1585 nor n3995 n4020 ; n4021
g1586 and n4017 n4021 ; n4022
g1587 and pi0299 n3944_not ; n4023
g1588 and pi0262 n3416 ; n4024
g1589 and pi0262_not n3499 ; n4025
g1590 nor pi0172 n4025 ; n4026
g1591 and pi0172 pi0262_not ; n4027
g1592 and n3508 n4027 ; n4028
g1593 nor n4026 n4028 ; n4029
g1594 nor pi0228 n4024 ; n4030
g1595 and n4029_not n4030 ; n4031
g1596 and n3487_not n3950 ; n4032
g1597 and pi0228 n3948_not ; n4033
g1598 and n4032_not n4033 ; n4034
g1599 and n3497_not n4034 ; n4035
g1600 nor pi0216 n4035 ; n4036
g1601 and n4031_not n4036 ; n4037
g1602 and n3946 n4037_not ; n4038
g1603 nor n3959 n4038 ; n4039
g1604 nor pi0215 n4039 ; n4040
g1605 and n4023 n4040_not ; n4041
g1606 and n3488_not n3989 ; n4042
g1607 and n4021 n4042_not ; n4043
g1608 nor pi0223 n4043 ; n4044
g1609 and n4017 n4044_not ; n4045
g1610 nor pi0039 n4045 ; n4046
g1611 and n4022_not n4046 ; n4047
g1612 and n4041_not n4047 ; n4048
g1613 nor pi0038 n4016 ; n4049
g1614 and n4048_not n4049 ; n4050
g1615 nor pi0100 n4015 ; n4051
g1616 and n4050_not n4051 ; n4052
g1617 and n2530_not n4002 ; n4053
g1618 and pi0262_not n3394 ; n4054
g1619 nor n3629 n3947 ; n4055
g1620 nor n4054 n4055 ; n4056
g1621 and n3969 n4056_not ; n4057
g1622 nor pi0216 n4057 ; n4058
g1623 and n3946 n4058_not ; n4059
g1624 nor n3959 n4059 ; n4060
g1625 nor pi0215 n4060 ; n4061
g1626 nor n3944 n4061 ; n4062
g1627 and pi0299 n4062_not ; n4063
g1628 and n2530 n4000_not ; n4064
g1629 and n4063_not n4064 ; n4065
g1630 and pi0100 n4053_not ; n4066
g1631 and n4065_not n4066 ; n4067
g1632 nor n4052 n4067 ; n4068
g1633 nor pi0087 n4068 ; n4069
g1634 nor pi0075 n4014 ; n4070
g1635 and n4069_not n4070 ; n4071
g1636 nor pi0092 n4013 ; n4072
g1637 and n4071_not n4072 ; n4073
g1638 and n2532 n4012_not ; n4074
g1639 and n4073_not n4074 ; n4075
g1640 nor pi0055 n4003 ; n4076
g1641 and n4075_not n4076 ; n4077
g1642 nor pi0056 n3986 ; n4078
g1643 and n4077_not n4078 ; n4079
g1644 nor pi0062 n3982 ; n4080
g1645 and n4079_not n4080 ; n4081
g1646 and n3328 n3978_not ; n4082
g1647 and n4081_not n4082 ; n4083
g1648 nor pi0249 n3964 ; n4084
g1649 and n4083_not n4084 ; n4085
g1650 and n3328_not n3962 ; n4086
g1651 and n3331_not n3962 ; n4087
g1652 nor n3952 n3968 ; n4088
g1653 nor pi0216 n4088 ; n4089
g1654 and n3946 n4089_not ; n4090
g1655 nor n3959 n4090 ; n4091
g1656 nor pi0215 n4091 ; n4092
g1657 nor n3944 n4092 ; n4093
g1658 and n3331 n4093 ; n4094
g1659 and pi0062 n4087_not ; n4095
g1660 and n4094_not n4095 ; n4096
g1661 nor n2537 n3962 ; n4097
g1662 and n2537 n4093_not ; n4098
g1663 and pi0056 n4097_not ; n4099
g1664 and n4098_not n4099 ; n4100
g1665 and n2572_not n3962 ; n4101
g1666 and n2572 n4093 ; n4102
g1667 and pi0055 n4101_not ; n4103
g1668 and n4102_not n4103 ; n4104
g1669 and pi0299 n3962_not ; n4105
g1670 nor n3999 n4105 ; n4106
g1671 and n2532_not n4106 ; n4107
g1672 and n2625_not n4106 ; n4108
g1673 and pi0299 n4093_not ; n4109
g1674 nor n3999 n4109 ; n4110
g1675 and n2625 n4110 ; n4111
g1676 nor n4108 n4111 ; n4112
g1677 and n2533 n4112_not ; n4113
g1678 and n2533_not n4106 ; n4114
g1679 and pi0092 n4114_not ; n4115
g1680 and n4113_not n4115 ; n4116
g1681 and pi0075 n4106 ; n4117
g1682 and pi0087 n4112 ; n4118
g1683 and pi0038 n4106 ; n4119
g1684 and pi0039 n4110_not ; n4120
g1685 and pi0262 n3508 ; n4121
g1686 nor pi0172 n4121 ; n4122
g1687 and pi0262 n3499_not ; n4123
g1688 nor pi0262 n3416 ; n4124
g1689 and pi0172 n4123_not ; n4125
g1690 and n4124_not n4125 ; n4126
g1691 nor n4122 n4126 ; n4127
g1692 nor pi0228 n4127 ; n4128
g1693 nor pi0216 n4034 ; n4129
g1694 and n4128_not n4129 ; n4130
g1695 and n3946 n4130_not ; n4131
g1696 nor n3959 n4131 ; n4132
g1697 nor pi0215 n4132 ; n4133
g1698 and n4023 n4133_not ; n4134
g1699 and n4046 n4134_not ; n4135
g1700 nor pi0038 n4120 ; n4136
g1701 and n4135_not n4136 ; n4137
g1702 nor pi0100 n4119 ; n4138
g1703 and n4137_not n4138 ; n4139
g1704 and n2530_not n4106 ; n4140
g1705 nor n3952 n4056 ; n4141
g1706 nor pi0216 n4141 ; n4142
g1707 and n3946 n4142_not ; n4143
g1708 nor n3959 n4143 ; n4144
g1709 nor pi0215 n4144 ; n4145
g1710 nor n3944 n4145 ; n4146
g1711 and pi0299 n4146_not ; n4147
g1712 and n2530 n3999_not ; n4148
g1713 and n4147_not n4148 ; n4149
g1714 and pi0100 n4140_not ; n4150
g1715 and n4149_not n4150 ; n4151
g1716 nor n4139 n4151 ; n4152
g1717 nor pi0087 n4152 ; n4153
g1718 nor pi0075 n4118 ; n4154
g1719 and n4153_not n4154 ; n4155
g1720 nor pi0092 n4117 ; n4156
g1721 and n4155_not n4156 ; n4157
g1722 and n2532 n4116_not ; n4158
g1723 and n4157_not n4158 ; n4159
g1724 nor pi0055 n4107 ; n4160
g1725 and n4159_not n4160 ; n4161
g1726 nor pi0056 n4104 ; n4162
g1727 and n4161_not n4162 ; n4163
g1728 nor pi0062 n4100 ; n4164
g1729 and n4163_not n4164 ; n4165
g1730 and n3328 n4096_not ; n4166
g1731 and n4165_not n4166 ; n4167
g1732 and pi0249 n4086_not ; n4168
g1733 and n4167_not n4168 ; n4169
g1734 or n4085 n4169 ; po0157
g1735 and pi0215 pi1141 ; n4171
g1736 and pi0216 pi0270 ; n4172
g1737 nor pi0221 n4172 ; n4173
g1738 and pi0105_not pi0171 ; n4174
g1739 and pi0861 n2442_not ; n4175
g1740 and pi0105 n4175_not ; n4176
g1741 and pi0228 n4174_not ; n4177
g1742 and n4176_not n4177 ; n4178
g1743 nor pi0216 n4178 ; n4179
g1744 nor pi0171 pi0228 ; n4180
g1745 and n4179 n4180_not ; n4181
g1746 and n4173 n4181_not ; n4182
g1747 nor pi1141 n2452 ; n4183
g1748 and pi0935_not n2452 ; n4184
g1749 and pi0221 n4183_not ; n4185
g1750 and n4184_not n4185 ; n4186
g1751 nor n4182 n4186 ; n4187
g1752 nor pi0215 n4187 ; n4188
g1753 nor n4171 n4188 ; n4189
g1754 and n3331_not n4189 ; n4190
g1755 and pi0861_not n2521 ; n4191
g1756 and pi0171 n2521_not ; n4192
g1757 nor pi0228 n4191 ; n4193
g1758 and n4192_not n4193 ; n4194
g1759 and n4179 n4194_not ; n4195
g1760 and n4173 n4195_not ; n4196
g1761 nor n4186 n4196 ; n4197
g1762 nor pi0215 n4197 ; n4198
g1763 nor n4171 n4198 ; n4199
g1764 and n3331 n4199 ; n4200
g1765 and pi0062 n4190_not ; n4201
g1766 and n4200_not n4201 ; n4202
g1767 nor n2537 n4189 ; n4203
g1768 and n2537 n4199_not ; n4204
g1769 and pi0056 n4203_not ; n4205
g1770 and n4204_not n4205 ; n4206
g1771 and n2572_not n4189 ; n4207
g1772 and n2572 n4199 ; n4208
g1773 and pi0055 n4207_not ; n4209
g1774 and n4208_not n4209 ; n4210
g1775 and pi0223 pi1141 ; n4211
g1776 and pi0224 pi0270 ; n4212
g1777 nor pi0222 n4212 ; n4213
g1778 nor pi0224 n4175 ; n4214
g1779 and n4213 n4214_not ; n4215
g1780 nor pi1141 n2591 ; n4216
g1781 and pi0935_not n2591 ; n4217
g1782 and pi0222 n4216_not ; n4218
g1783 and n4217_not n4218 ; n4219
g1784 nor n4215 n4219 ; n4220
g1785 nor pi0223 n4220 ; n4221
g1786 nor n4211 n4221 ; n4222
g1787 nor pi0299 n4222 ; n4223
g1788 and pi0299 n4189_not ; n4224
g1789 nor n4223 n4224 ; n4225
g1790 and n2532_not n4225 ; n4226
g1791 and n2625_not n4225 ; n4227
g1792 and pi0299 n4199_not ; n4228
g1793 nor n4223 n4228 ; n4229
g1794 and n2625 n4229 ; n4230
g1795 nor n4227 n4230 ; n4231
g1796 and n2533 n4231_not ; n4232
g1797 and n2533_not n4225 ; n4233
g1798 and pi0092 n4233_not ; n4234
g1799 and n4232_not n4234 ; n4235
g1800 and pi0075 n4225 ; n4236
g1801 and pi0087 n4231 ; n4237
g1802 and pi0038 n4225 ; n4238
g1803 and pi0039 n4229_not ; n4239
g1804 nor pi0299 n4211 ; n4240
g1805 and pi0861 n3488 ; n4241
g1806 nor pi0224 n4241 ; n4242
g1807 and n4213 n4242_not ; n4243
g1808 nor n4219 n4243 ; n4244
g1809 and n4240 n4244 ; n4245
g1810 and pi0299 n4171_not ; n4246
g1811 and pi0861 n3499 ; n4247
g1812 nor pi0171 n4247 ; n4248
g1813 and pi0171 n3508 ; n4249
g1814 nor n4248 n4249 ; n4250
g1815 and pi0861 n4250_not ; n4251
g1816 and n3416_not n4248 ; n4252
g1817 nor n4251 n4252 ; n4253
g1818 nor pi0228 n4253 ; n4254
g1819 and n3497_not n4178 ; n4255
g1820 nor pi0216 n4255 ; n4256
g1821 and n4254_not n4256 ; n4257
g1822 and n4173 n4257_not ; n4258
g1823 nor n4186 n4258 ; n4259
g1824 nor pi0215 n4259 ; n4260
g1825 and n4246 n4260_not ; n4261
g1826 and n3488_not n4213 ; n4262
g1827 and n4244 n4262_not ; n4263
g1828 nor pi0223 n4263 ; n4264
g1829 and n4240 n4264_not ; n4265
g1830 nor pi0039 n4265 ; n4266
g1831 and n4245_not n4266 ; n4267
g1832 and n4261_not n4267 ; n4268
g1833 nor pi0038 n4239 ; n4269
g1834 and n4268_not n4269 ; n4270
g1835 nor pi0100 n4238 ; n4271
g1836 and n4270_not n4271 ; n4272
g1837 and n2530_not n4225 ; n4273
g1838 and pi0861_not n3394 ; n4274
g1839 and pi0171 n3394_not ; n4275
g1840 nor pi0228 n4274 ; n4276
g1841 and n4275_not n4276 ; n4277
g1842 and n4179 n4277_not ; n4278
g1843 and n4173 n4278_not ; n4279
g1844 nor n4186 n4279 ; n4280
g1845 nor pi0215 n4280 ; n4281
g1846 nor n4171 n4281 ; n4282
g1847 and pi0299 n4282_not ; n4283
g1848 and n2530 n4223_not ; n4284
g1849 and n4283_not n4284 ; n4285
g1850 and pi0100 n4273_not ; n4286
g1851 and n4285_not n4286 ; n4287
g1852 nor n4272 n4287 ; n4288
g1853 nor pi0087 n4288 ; n4289
g1854 nor pi0075 n4237 ; n4290
g1855 and n4289_not n4290 ; n4291
g1856 nor pi0092 n4236 ; n4292
g1857 and n4291_not n4292 ; n4293
g1858 and n2532 n4235_not ; n4294
g1859 and n4293_not n4294 ; n4295
g1860 nor pi0055 n4226 ; n4296
g1861 and n4295_not n4296 ; n4297
g1862 nor pi0056 n4210 ; n4298
g1863 and n4297_not n4298 ; n4299
g1864 nor pi0062 n4206 ; n4300
g1865 and n4299_not n4300 ; n4301
g1866 and pi0241_not n3328 ; n4302
g1867 and n4202_not n4302 ; n4303
g1868 and n4301_not n4303 ; n4304
g1869 and n3447_not n4179 ; n4305
g1870 and n4194_not n4305 ; n4306
g1871 and n4173 n4306_not ; n4307
g1872 nor n4186 n4307 ; n4308
g1873 nor pi0215 n4308 ; n4309
g1874 nor n4171 n4309 ; n4310
g1875 and n3331 n4310 ; n4311
g1876 and n3556 n4172_not ; n4312
g1877 and n4189 n4312_not ; n4313
g1878 and n3331_not n4313 ; n4314
g1879 and pi0062 n4314_not ; n4315
g1880 and n4311_not n4315 ; n4316
g1881 nor n2537 n4313 ; n4317
g1882 and n2537 n4310_not ; n4318
g1883 and pi0056 n4317_not ; n4319
g1884 and n4318_not n4319 ; n4320
g1885 and n2572 n4310 ; n4321
g1886 and n2572_not n4313 ; n4322
g1887 and pi0055 n4322_not ; n4323
g1888 and n4321_not n4323 ; n4324
g1889 nor n3472 n4223 ; n4325
g1890 and pi0299 n4313_not ; n4326
g1891 and n4325 n4326_not ; n4327
g1892 and n2532_not n4327 ; n4328
g1893 and n2625_not n4327 ; n4329
g1894 and pi0299 n4310_not ; n4330
g1895 and n4325 n4330_not ; n4331
g1896 and n2625 n4331 ; n4332
g1897 nor n4329 n4332 ; n4333
g1898 and n2533 n4333_not ; n4334
g1899 and n2533_not n4327 ; n4335
g1900 and pi0092 n4335_not ; n4336
g1901 and n4334_not n4336 ; n4337
g1902 and pi0075 n4327 ; n4338
g1903 and pi0087 n4333 ; n4339
g1904 and pi0038 n4327 ; n4340
g1905 and pi0039 n4331_not ; n4341
g1906 and pi0861_not n3508 ; n4342
g1907 nor pi0171 n4342 ; n4343
g1908 nor pi0861 n3499 ; n4344
g1909 and pi0861 n3416_not ; n4345
g1910 and pi0171 n4344_not ; n4346
g1911 and n4345_not n4346 ; n4347
g1912 nor n4343 n4347 ; n4348
g1913 nor pi0228 n4348 ; n4349
g1914 and n3793_not n4179 ; n4350
g1915 and n4349_not n4350 ; n4351
g1916 and n4173 n4351_not ; n4352
g1917 nor n4186 n4352 ; n4353
g1918 nor pi0215 n4353 ; n4354
g1919 and n4246 n4354_not ; n4355
g1920 and n4266 n4355_not ; n4356
g1921 nor pi0038 n4341 ; n4357
g1922 and n4356_not n4357 ; n4358
g1923 nor pi0100 n4340 ; n4359
g1924 and n4358_not n4359 ; n4360
g1925 and n2530_not n4327 ; n4361
g1926 and n4277_not n4305 ; n4362
g1927 and n4173 n4362_not ; n4363
g1928 nor n4186 n4363 ; n4364
g1929 nor pi0215 n4364 ; n4365
g1930 nor n4171 n4365 ; n4366
g1931 and pi0299 n4366_not ; n4367
g1932 and n2530 n4325 ; n4368
g1933 and n4367_not n4368 ; n4369
g1934 and pi0100 n4361_not ; n4370
g1935 and n4369_not n4370 ; n4371
g1936 nor n4360 n4371 ; n4372
g1937 nor pi0087 n4372 ; n4373
g1938 nor pi0075 n4339 ; n4374
g1939 and n4373_not n4374 ; n4375
g1940 nor pi0092 n4338 ; n4376
g1941 and n4375_not n4376 ; n4377
g1942 and n2532 n4337_not ; n4378
g1943 and n4377_not n4378 ; n4379
g1944 nor pi0055 n4328 ; n4380
g1945 and n4379_not n4380 ; n4381
g1946 nor pi0056 n4324 ; n4382
g1947 and n4381_not n4382 ; n4383
g1948 nor pi0062 n4320 ; n4384
g1949 and n4383_not n4384 ; n4385
g1950 and pi0241 n3328 ; n4386
g1951 and n4316_not n4386 ; n4387
g1952 and n4385_not n4387 ; n4388
g1953 and pi0241 n4312 ; n4389
g1954 nor n3328 n4389 ; n4390
g1955 and n4189 n4390 ; n4391
g1956 nor n4388 n4391 ; n4392
g1957 and n4304_not n4392 ; po0158
g1958 and pi0215 pi1140 ; n4394
g1959 and pi0216 pi0282 ; n4395
g1960 nor pi0221 n4395 ; n4396
g1961 and pi0105_not pi0170 ; n4397
g1962 and pi0869 n2442_not ; n4398
g1963 and pi0105 n4398_not ; n4399
g1964 and pi0228 n4397_not ; n4400
g1965 and n4399_not n4400 ; n4401
g1966 nor pi0216 n4401 ; n4402
g1967 nor pi0170 pi0228 ; n4403
g1968 and n4402 n4403_not ; n4404
g1969 and n4396 n4404_not ; n4405
g1970 nor pi1140 n2452 ; n4406
g1971 and pi0921_not n2452 ; n4407
g1972 and pi0221 n4406_not ; n4408
g1973 and n4407_not n4408 ; n4409
g1974 nor n4405 n4409 ; n4410
g1975 nor pi0215 n4410 ; n4411
g1976 nor n4394 n4411 ; n4412
g1977 and n3331_not n4412 ; n4413
g1978 and pi0869_not n2521 ; n4414
g1979 and pi0170 n2521_not ; n4415
g1980 nor pi0228 n4414 ; n4416
g1981 and n4415_not n4416 ; n4417
g1982 and n4402 n4417_not ; n4418
g1983 and n4396 n4418_not ; n4419
g1984 nor n4409 n4419 ; n4420
g1985 nor pi0215 n4420 ; n4421
g1986 nor n4394 n4421 ; n4422
g1987 and n3331 n4422 ; n4423
g1988 and pi0062 n4413_not ; n4424
g1989 and n4423_not n4424 ; n4425
g1990 nor n2537 n4412 ; n4426
g1991 and n2537 n4422_not ; n4427
g1992 and pi0056 n4426_not ; n4428
g1993 and n4427_not n4428 ; n4429
g1994 and n2572_not n4412 ; n4430
g1995 and n2572 n4422 ; n4431
g1996 and pi0055 n4430_not ; n4432
g1997 and n4431_not n4432 ; n4433
g1998 and pi0223 pi1140 ; n4434
g1999 and pi0224 pi0282 ; n4435
g2000 nor pi0222 n4435 ; n4436
g2001 nor pi0224 n4398 ; n4437
g2002 and n4436 n4437_not ; n4438
g2003 nor pi1140 n2591 ; n4439
g2004 and pi0921_not n2591 ; n4440
g2005 and pi0222 n4439_not ; n4441
g2006 and n4440_not n4441 ; n4442
g2007 nor n4438 n4442 ; n4443
g2008 nor pi0223 n4443 ; n4444
g2009 nor n4434 n4444 ; n4445
g2010 nor pi0299 n4445 ; n4446
g2011 and pi0299 n4412_not ; n4447
g2012 nor n4446 n4447 ; n4448
g2013 and n2532_not n4448 ; n4449
g2014 and n2625_not n4448 ; n4450
g2015 and pi0299 n4422_not ; n4451
g2016 nor n4446 n4451 ; n4452
g2017 and n2625 n4452 ; n4453
g2018 nor n4450 n4453 ; n4454
g2019 and n2533 n4454_not ; n4455
g2020 and n2533_not n4448 ; n4456
g2021 and pi0092 n4456_not ; n4457
g2022 and n4455_not n4457 ; n4458
g2023 and pi0075 n4448 ; n4459
g2024 and pi0087 n4454 ; n4460
g2025 and pi0038 n4448 ; n4461
g2026 and pi0039 n4452_not ; n4462
g2027 nor pi0299 n4434 ; n4463
g2028 and pi0869 n3488 ; n4464
g2029 nor pi0224 n4464 ; n4465
g2030 and n4436 n4465_not ; n4466
g2031 nor n4442 n4466 ; n4467
g2032 and n4463 n4467 ; n4468
g2033 and pi0299 n4394_not ; n4469
g2034 and pi0869 n3499 ; n4470
g2035 nor pi0170 n4470 ; n4471
g2036 and pi0170 n3508 ; n4472
g2037 nor n4471 n4472 ; n4473
g2038 and pi0869 n4473_not ; n4474
g2039 and n3416_not n4471 ; n4475
g2040 nor n4474 n4475 ; n4476
g2041 nor pi0228 n4476 ; n4477
g2042 and n3497_not n4401 ; n4478
g2043 nor pi0216 n4478 ; n4479
g2044 and n4477_not n4479 ; n4480
g2045 and n4396 n4480_not ; n4481
g2046 nor n4409 n4481 ; n4482
g2047 nor pi0215 n4482 ; n4483
g2048 and n4469 n4483_not ; n4484
g2049 and n3488_not n4436 ; n4485
g2050 and n4467 n4485_not ; n4486
g2051 nor pi0223 n4486 ; n4487
g2052 and n4463 n4487_not ; n4488
g2053 nor pi0039 n4488 ; n4489
g2054 and n4468_not n4489 ; n4490
g2055 and n4484_not n4490 ; n4491
g2056 nor pi0038 n4462 ; n4492
g2057 and n4491_not n4492 ; n4493
g2058 nor pi0100 n4461 ; n4494
g2059 and n4493_not n4494 ; n4495
g2060 and n2530_not n4448 ; n4496
g2061 and pi0869_not n3394 ; n4497
g2062 and pi0170 n3394_not ; n4498
g2063 nor pi0228 n4497 ; n4499
g2064 and n4498_not n4499 ; n4500
g2065 and n4402 n4500_not ; n4501
g2066 and n4396 n4501_not ; n4502
g2067 nor n4409 n4502 ; n4503
g2068 nor pi0215 n4503 ; n4504
g2069 nor n4394 n4504 ; n4505
g2070 and pi0299 n4505_not ; n4506
g2071 and n2530 n4446_not ; n4507
g2072 and n4506_not n4507 ; n4508
g2073 and pi0100 n4496_not ; n4509
g2074 and n4508_not n4509 ; n4510
g2075 nor n4495 n4510 ; n4511
g2076 nor pi0087 n4511 ; n4512
g2077 nor pi0075 n4460 ; n4513
g2078 and n4512_not n4513 ; n4514
g2079 nor pi0092 n4459 ; n4515
g2080 and n4514_not n4515 ; n4516
g2081 and n2532 n4458_not ; n4517
g2082 and n4516_not n4517 ; n4518
g2083 nor pi0055 n4449 ; n4519
g2084 and n4518_not n4519 ; n4520
g2085 nor pi0056 n4433 ; n4521
g2086 and n4520_not n4521 ; n4522
g2087 nor pi0062 n4429 ; n4523
g2088 and n4522_not n4523 ; n4524
g2089 and pi0248_not n3328 ; n4525
g2090 and n4425_not n4525 ; n4526
g2091 and n4524_not n4526 ; n4527
g2092 and n3447_not n4402 ; n4528
g2093 and n4417_not n4528 ; n4529
g2094 and n4396 n4529_not ; n4530
g2095 nor n4409 n4530 ; n4531
g2096 nor pi0215 n4531 ; n4532
g2097 nor n4394 n4532 ; n4533
g2098 and n3331 n4533 ; n4534
g2099 and n3556 n4395_not ; n4535
g2100 and n4412 n4535_not ; n4536
g2101 and n3331_not n4536 ; n4537
g2102 and pi0062 n4537_not ; n4538
g2103 and n4534_not n4538 ; n4539
g2104 nor n2537 n4536 ; n4540
g2105 and n2537 n4533_not ; n4541
g2106 and pi0056 n4540_not ; n4542
g2107 and n4541_not n4542 ; n4543
g2108 and n2572 n4533 ; n4544
g2109 and n2572_not n4536 ; n4545
g2110 and pi0055 n4545_not ; n4546
g2111 and n4544_not n4546 ; n4547
g2112 nor n3472 n4446 ; n4548
g2113 and pi0299 n4536_not ; n4549
g2114 and n4548 n4549_not ; n4550
g2115 and n2532_not n4550 ; n4551
g2116 and n2625_not n4550 ; n4552
g2117 and pi0299 n4533_not ; n4553
g2118 and n4548 n4553_not ; n4554
g2119 and n2625 n4554 ; n4555
g2120 nor n4552 n4555 ; n4556
g2121 and n2533 n4556_not ; n4557
g2122 and n2533_not n4550 ; n4558
g2123 and pi0092 n4558_not ; n4559
g2124 and n4557_not n4559 ; n4560
g2125 and pi0075 n4550 ; n4561
g2126 and pi0087 n4556 ; n4562
g2127 and pi0038 n4550 ; n4563
g2128 and pi0039 n4554_not ; n4564
g2129 and pi0869_not n3508 ; n4565
g2130 nor pi0170 n4565 ; n4566
g2131 nor pi0869 n3499 ; n4567
g2132 and pi0869 n3416_not ; n4568
g2133 and pi0170 n4567_not ; n4569
g2134 and n4568_not n4569 ; n4570
g2135 nor n4566 n4570 ; n4571
g2136 nor pi0228 n4571 ; n4572
g2137 and n3793_not n4402 ; n4573
g2138 and n4572_not n4573 ; n4574
g2139 and n4396 n4574_not ; n4575
g2140 nor n4409 n4575 ; n4576
g2141 nor pi0215 n4576 ; n4577
g2142 and n4469 n4577_not ; n4578
g2143 and n4489 n4578_not ; n4579
g2144 nor pi0038 n4564 ; n4580
g2145 and n4579_not n4580 ; n4581
g2146 nor pi0100 n4563 ; n4582
g2147 and n4581_not n4582 ; n4583
g2148 and n2530_not n4550 ; n4584
g2149 and n4500_not n4528 ; n4585
g2150 and n4396 n4585_not ; n4586
g2151 nor n4409 n4586 ; n4587
g2152 nor pi0215 n4587 ; n4588
g2153 nor n4394 n4588 ; n4589
g2154 and pi0299 n4589_not ; n4590
g2155 and n2530 n4548 ; n4591
g2156 and n4590_not n4591 ; n4592
g2157 and pi0100 n4584_not ; n4593
g2158 and n4592_not n4593 ; n4594
g2159 nor n4583 n4594 ; n4595
g2160 nor pi0087 n4595 ; n4596
g2161 nor pi0075 n4562 ; n4597
g2162 and n4596_not n4597 ; n4598
g2163 nor pi0092 n4561 ; n4599
g2164 and n4598_not n4599 ; n4600
g2165 and n2532 n4560_not ; n4601
g2166 and n4600_not n4601 ; n4602
g2167 nor pi0055 n4551 ; n4603
g2168 and n4602_not n4603 ; n4604
g2169 nor pi0056 n4547 ; n4605
g2170 and n4604_not n4605 ; n4606
g2171 nor pi0062 n4543 ; n4607
g2172 and n4606_not n4607 ; n4608
g2173 and pi0248 n3328 ; n4609
g2174 and n4539_not n4609 ; n4610
g2175 and n4608_not n4610 ; n4611
g2176 and pi0248 n4535 ; n4612
g2177 nor n3328 n4612 ; n4613
g2178 and n4412 n4613 ; n4614
g2179 nor n4611 n4614 ; n4615
g2180 and n4527_not n4615 ; po0159
g2181 and pi0215 pi1139 ; n4617
g2182 and pi0216 pi1139_not ; n4618
g2183 and pi0833 pi0920 ; n4619
g2184 and pi0833_not pi1139 ; n4620
g2185 nor pi0216 n4619 ; n4621
g2186 and n4620_not n4621 ; n4622
g2187 and pi0221 n4622_not ; n4623
g2188 and n4618_not n4623 ; n4624
g2189 and pi0216 pi0281 ; n4625
g2190 nor pi0221 n4625 ; n4626
g2191 nor pi0216 pi0862 ; n4627
g2192 and n3630 n4627 ; n4628
g2193 and n4626 n4628_not ; n4629
g2194 nor n4624 n4629 ; n4630
g2195 nor pi0216 n4623 ; n4631
g2196 and pi0148 n2441_not ; n4632
g2197 and n4631 n4632 ; n4633
g2198 nor pi0215 n4633 ; n4634
g2199 and n4630_not n4634 ; n4635
g2200 nor n4617 n4635 ; n4636
g2201 nor n3450 n4636 ; n4637
g2202 nor n3328 n4637 ; n4638
g2203 nor n3331 n4637 ; n4639
g2204 nor pi0148 pi0215 ; n4640
g2205 and pi0862 n3447_not ; n4641
g2206 nor n2441 n3335 ; n4642
g2207 nor pi0216 n4641 ; n4643
g2208 and n4642_not n4643 ; n4644
g2209 and n4626 n4644_not ; n4645
g2210 nor n4624 n4645 ; n4646
g2211 and n4640 n4646_not ; n4647
g2212 and pi0148 pi0215_not ; n4648
g2213 nor n3335 n3630 ; n4649
g2214 and n4627 n4649_not ; n4650
g2215 and n4626 n4650_not ; n4651
g2216 nor n4624 n4651 ; n4652
g2217 and n4631 n4649 ; n4653
g2218 and n4648 n4653_not ; n4654
g2219 and n4652_not n4654 ; n4655
g2220 nor n4617 n4655 ; n4656
g2221 and n4647_not n4656 ; n4657
g2222 and n3331 n4657 ; n4658
g2223 and pi0062 n4639_not ; n4659
g2224 and n4658_not n4659 ; n4660
g2225 and n2537 n4657_not ; n4661
g2226 and n2537_not n4637 ; n4662
g2227 and pi0056 n4662_not ; n4663
g2228 and n4661_not n4663 ; n4664
g2229 nor n2572 n4637 ; n4665
g2230 and n2572 n4657 ; n4666
g2231 and pi0055 n4665_not ; n4667
g2232 and n4666_not n4667 ; n4668
g2233 and pi0223 pi1139 ; n4669
g2234 nor pi1139 n2591 ; n4670
g2235 and pi0920_not n2591 ; n4671
g2236 and pi0222 n4670_not ; n4672
g2237 and n4671_not n4672 ; n4673
g2238 nor pi0224 n4669 ; n4674
g2239 and n4673_not n4674 ; n4675
g2240 and n2442 n4675 ; n4676
g2241 and pi0862_not n4675 ; n4677
g2242 and pi0224 pi0281 ; n4678
g2243 nor pi0222 n4678 ; n4679
g2244 nor n4673 n4679 ; n4680
g2245 nor pi0223 n4680 ; n4681
g2246 nor n4669 n4681 ; n4682
g2247 nor pi0299 n4682 ; n4683
g2248 and n4677_not n4683 ; n4684
g2249 and n4676_not n4684 ; n4685
g2250 and pi0299 n4637 ; n4686
g2251 nor n4685 n4686 ; n4687
g2252 and n2532_not n4687 ; n4688
g2253 and n2625_not n4687 ; n4689
g2254 and pi0299 n4657_not ; n4690
g2255 nor n4685 n4690 ; n4691
g2256 and n2625 n4691 ; n4692
g2257 nor n4689 n4692 ; n4693
g2258 and n2533 n4693_not ; n4694
g2259 and n2533_not n4687 ; n4695
g2260 and pi0092 n4695_not ; n4696
g2261 and n4694_not n4696 ; n4697
g2262 and pi0075 n4687 ; n4698
g2263 and pi0087 n4693 ; n4699
g2264 and n2530_not n4687 ; n4700
g2265 nor n2441 n3629 ; n4701
g2266 and n4626 n4701 ; n4702
g2267 and n4646 n4702_not ; n4703
g2268 and n4640 n4703_not ; n4704
g2269 and n3631 n4626 ; n4705
g2270 and n4652 n4705_not ; n4706
g2271 and n3631 n4631 ; n4707
g2272 and n4648 n4707_not ; n4708
g2273 and n4706_not n4708 ; n4709
g2274 nor n4617 n4704 ; n4710
g2275 and n4709_not n4710 ; n4711
g2276 and pi0299 n4711_not ; n4712
g2277 and n2530 n4685_not ; n4713
g2278 and n4712_not n4713 ; n4714
g2279 and pi0100 n4700_not ; n4715
g2280 and n4714_not n4715 ; n4716
g2281 and pi0038 n4687 ; n4717
g2282 and pi0039 n4691_not ; n4718
g2283 and n3488_not n4675 ; n4719
g2284 nor n4677 n4682 ; n4720
g2285 and n4719_not n4720 ; n4721
g2286 nor pi0299 n4721 ; n4722
g2287 and n3511_not n4627 ; n4723
g2288 and n4626 n4723_not ; n4724
g2289 nor n4624 n4724 ; n4725
g2290 and n3511 n4631 ; n4726
g2291 and n4648 n4726_not ; n4727
g2292 and n4725_not n4727 ; n4728
g2293 and pi0862 n3501_not ; n4729
g2294 and pi0228_not n3416 ; n4730
g2295 nor n2441 n4730 ; n4731
g2296 and pi0862_not n4731 ; n4732
g2297 nor pi0216 n4729 ; n4733
g2298 and n4732_not n4733 ; n4734
g2299 and n4626 n4734_not ; n4735
g2300 nor n4624 n4735 ; n4736
g2301 and n4640 n4736_not ; n4737
g2302 and pi0299 n4617_not ; n4738
g2303 and n4728_not n4738 ; n4739
g2304 and n4737_not n4739 ; n4740
g2305 nor pi0039 n4722 ; n4741
g2306 and n4740_not n4741 ; n4742
g2307 nor pi0038 n4718 ; n4743
g2308 and n4742_not n4743 ; n4744
g2309 nor pi0100 n4717 ; n4745
g2310 and n4744_not n4745 ; n4746
g2311 nor n4716 n4746 ; n4747
g2312 nor pi0087 n4747 ; n4748
g2313 nor pi0075 n4699 ; n4749
g2314 and n4748_not n4749 ; n4750
g2315 nor pi0092 n4698 ; n4751
g2316 and n4750_not n4751 ; n4752
g2317 and n2532 n4697_not ; n4753
g2318 and n4752_not n4753 ; n4754
g2319 nor pi0055 n4688 ; n4755
g2320 and n4754_not n4755 ; n4756
g2321 nor pi0056 n4668 ; n4757
g2322 and n4756_not n4757 ; n4758
g2323 nor pi0062 n4664 ; n4759
g2324 and n4758_not n4759 ; n4760
g2325 and n3328 n4660_not ; n4761
g2326 and n4760_not n4761 ; n4762
g2327 nor pi0247 n4638 ; n4763
g2328 and n4762_not n4763 ; n4764
g2329 and n3328_not n4636 ; n4765
g2330 and n3331_not n4636 ; n4766
g2331 and n4634 n4652_not ; n4767
g2332 and n4656 n4767_not ; n4768
g2333 and n3331 n4768 ; n4769
g2334 and pi0062 n4766_not ; n4770
g2335 and n4769_not n4770 ; n4771
g2336 nor n2537 n4636 ; n4772
g2337 and n2537 n4768_not ; n4773
g2338 and pi0056 n4772_not ; n4774
g2339 and n4773_not n4774 ; n4775
g2340 and n2572_not n4636 ; n4776
g2341 and n2572 n4768 ; n4777
g2342 and pi0055 n4776_not ; n4778
g2343 and n4777_not n4778 ; n4779
g2344 nor n3472 n4684 ; n4780
g2345 and pi0299 n4636_not ; n4781
g2346 and n4780 n4781_not ; n4782
g2347 and n2532_not n4782 ; n4783
g2348 and n2625_not n4782 ; n4784
g2349 and pi0299 n4768_not ; n4785
g2350 and n4780 n4785_not ; n4786
g2351 and n2625 n4786 ; n4787
g2352 nor n4784 n4787 ; n4788
g2353 and n2533 n4788_not ; n4789
g2354 and n2533_not n4782 ; n4790
g2355 and pi0092 n4790_not ; n4791
g2356 and n4789_not n4791 ; n4792
g2357 and pi0075 n4782 ; n4793
g2358 and pi0087 n4788 ; n4794
g2359 and n2530_not n4782 ; n4795
g2360 and n4640 n4706_not ; n4796
g2361 nor pi0216 n4624 ; n4797
g2362 and n4701 n4797 ; n4798
g2363 and n4648 n4652_not ; n4799
g2364 and n4798_not n4799 ; n4800
g2365 nor n4617 n4800 ; n4801
g2366 and n4796_not n4801 ; n4802
g2367 and pi0299 n4802_not ; n4803
g2368 and n2530 n4780 ; n4804
g2369 and n4803_not n4804 ; n4805
g2370 and pi0100 n4795_not ; n4806
g2371 and n4805_not n4806 ; n4807
g2372 and pi0038 n4782 ; n4808
g2373 and pi0039 n4786_not ; n4809
g2374 and n3488 n4677 ; n4810
g2375 and n4683 n4810_not ; n4811
g2376 and pi0862 n4731_not ; n4812
g2377 and pi0862_not n3501 ; n4813
g2378 nor pi0216 n4813 ; n4814
g2379 and n4812_not n4814 ; n4815
g2380 and n4626 n4815_not ; n4816
g2381 nor n4624 n4816 ; n4817
g2382 and n4648 n4817_not ; n4818
g2383 and n4640 n4725_not ; n4819
g2384 nor n4617 n4819 ; n4820
g2385 and n4818_not n4820 ; n4821
g2386 and pi0299 n4821_not ; n4822
g2387 nor n4811 n4822 ; n4823
g2388 nor pi0039 n4823 ; n4824
g2389 nor pi0038 n4809 ; n4825
g2390 and n4824_not n4825 ; n4826
g2391 nor pi0100 n4808 ; n4827
g2392 and n4826_not n4827 ; n4828
g2393 nor n4807 n4828 ; n4829
g2394 nor pi0087 n4829 ; n4830
g2395 nor pi0075 n4794 ; n4831
g2396 and n4830_not n4831 ; n4832
g2397 nor pi0092 n4793 ; n4833
g2398 and n4832_not n4833 ; n4834
g2399 and n2532 n4792_not ; n4835
g2400 and n4834_not n4835 ; n4836
g2401 nor pi0055 n4783 ; n4837
g2402 and n4836_not n4837 ; n4838
g2403 nor pi0056 n4779 ; n4839
g2404 and n4838_not n4839 ; n4840
g2405 nor pi0062 n4775 ; n4841
g2406 and n4840_not n4841 ; n4842
g2407 and n3328 n4771_not ; n4843
g2408 and n4842_not n4843 ; n4844
g2409 and pi0247 n4765_not ; n4845
g2410 and n4844_not n4845 ; n4846
g2411 or n4764 n4846 ; po0160
g2412 and pi0215 pi1138 ; n4848
g2413 and pi0216 pi0269 ; n4849
g2414 nor pi0221 n4849 ; n4850
g2415 and pi0105_not pi0169 ; n4851
g2416 and pi0877 n2442_not ; n4852
g2417 and pi0105 n4852_not ; n4853
g2418 and pi0228 n4851_not ; n4854
g2419 and n4853_not n4854 ; n4855
g2420 nor pi0216 n4855 ; n4856
g2421 nor pi0169 pi0228 ; n4857
g2422 and n4856 n4857_not ; n4858
g2423 and n4850 n4858_not ; n4859
g2424 nor pi1138 n2452 ; n4860
g2425 and pi0940_not n2452 ; n4861
g2426 and pi0221 n4860_not ; n4862
g2427 and n4861_not n4862 ; n4863
g2428 nor n4859 n4863 ; n4864
g2429 nor pi0215 n4864 ; n4865
g2430 nor n4848 n4865 ; n4866
g2431 and n3331_not n4866 ; n4867
g2432 and pi0877_not n2521 ; n4868
g2433 and pi0169 n2521_not ; n4869
g2434 nor pi0228 n4868 ; n4870
g2435 and n4869_not n4870 ; n4871
g2436 and n4856 n4871_not ; n4872
g2437 and n4850 n4872_not ; n4873
g2438 nor n4863 n4873 ; n4874
g2439 nor pi0215 n4874 ; n4875
g2440 nor n4848 n4875 ; n4876
g2441 and n3331 n4876 ; n4877
g2442 and pi0062 n4867_not ; n4878
g2443 and n4877_not n4878 ; n4879
g2444 nor n2537 n4866 ; n4880
g2445 and n2537 n4876_not ; n4881
g2446 and pi0056 n4880_not ; n4882
g2447 and n4881_not n4882 ; n4883
g2448 and n2572_not n4866 ; n4884
g2449 and n2572 n4876 ; n4885
g2450 and pi0055 n4884_not ; n4886
g2451 and n4885_not n4886 ; n4887
g2452 and pi0223 pi1138 ; n4888
g2453 and pi0224 pi0269 ; n4889
g2454 nor pi0222 n4889 ; n4890
g2455 nor pi0224 n4852 ; n4891
g2456 and n4890 n4891_not ; n4892
g2457 nor pi1138 n2591 ; n4893
g2458 and pi0940_not n2591 ; n4894
g2459 and pi0222 n4893_not ; n4895
g2460 and n4894_not n4895 ; n4896
g2461 nor n4892 n4896 ; n4897
g2462 nor pi0223 n4897 ; n4898
g2463 nor n4888 n4898 ; n4899
g2464 nor pi0299 n4899 ; n4900
g2465 and pi0299 n4866_not ; n4901
g2466 nor n4900 n4901 ; n4902
g2467 and n2532_not n4902 ; n4903
g2468 and n2625_not n4902 ; n4904
g2469 and pi0299 n4876_not ; n4905
g2470 nor n4900 n4905 ; n4906
g2471 and n2625 n4906 ; n4907
g2472 nor n4904 n4907 ; n4908
g2473 and n2533 n4908_not ; n4909
g2474 and n2533_not n4902 ; n4910
g2475 and pi0092 n4910_not ; n4911
g2476 and n4909_not n4911 ; n4912
g2477 and pi0075 n4902 ; n4913
g2478 and pi0087 n4908 ; n4914
g2479 and pi0038 n4902 ; n4915
g2480 and pi0039 n4906_not ; n4916
g2481 nor pi0299 n4888 ; n4917
g2482 and pi0877 n3488 ; n4918
g2483 nor pi0224 n4918 ; n4919
g2484 and n4890 n4919_not ; n4920
g2485 nor n4896 n4920 ; n4921
g2486 and n4917 n4921 ; n4922
g2487 and pi0299 n4848_not ; n4923
g2488 and pi0877 n3499 ; n4924
g2489 nor pi0169 n4924 ; n4925
g2490 and pi0169 n3508 ; n4926
g2491 nor n4925 n4926 ; n4927
g2492 and pi0877 n4927_not ; n4928
g2493 and n3416_not n4925 ; n4929
g2494 nor n4928 n4929 ; n4930
g2495 nor pi0228 n4930 ; n4931
g2496 and n3497_not n4855 ; n4932
g2497 nor pi0216 n4932 ; n4933
g2498 and n4931_not n4933 ; n4934
g2499 and n4850 n4934_not ; n4935
g2500 nor n4863 n4935 ; n4936
g2501 nor pi0215 n4936 ; n4937
g2502 and n4923 n4937_not ; n4938
g2503 and n3488_not n4890 ; n4939
g2504 and n4921 n4939_not ; n4940
g2505 nor pi0223 n4940 ; n4941
g2506 and n4917 n4941_not ; n4942
g2507 nor pi0039 n4942 ; n4943
g2508 and n4922_not n4943 ; n4944
g2509 and n4938_not n4944 ; n4945
g2510 nor pi0038 n4916 ; n4946
g2511 and n4945_not n4946 ; n4947
g2512 nor pi0100 n4915 ; n4948
g2513 and n4947_not n4948 ; n4949
g2514 and n2530_not n4902 ; n4950
g2515 and pi0877_not n3394 ; n4951
g2516 and pi0169 n3394_not ; n4952
g2517 nor pi0228 n4951 ; n4953
g2518 and n4952_not n4953 ; n4954
g2519 and n4856 n4954_not ; n4955
g2520 and n4850 n4955_not ; n4956
g2521 nor n4863 n4956 ; n4957
g2522 nor pi0215 n4957 ; n4958
g2523 nor n4848 n4958 ; n4959
g2524 and pi0299 n4959_not ; n4960
g2525 and n2530 n4900_not ; n4961
g2526 and n4960_not n4961 ; n4962
g2527 and pi0100 n4950_not ; n4963
g2528 and n4962_not n4963 ; n4964
g2529 nor n4949 n4964 ; n4965
g2530 nor pi0087 n4965 ; n4966
g2531 nor pi0075 n4914 ; n4967
g2532 and n4966_not n4967 ; n4968
g2533 nor pi0092 n4913 ; n4969
g2534 and n4968_not n4969 ; n4970
g2535 and n2532 n4912_not ; n4971
g2536 and n4970_not n4971 ; n4972
g2537 nor pi0055 n4903 ; n4973
g2538 and n4972_not n4973 ; n4974
g2539 nor pi0056 n4887 ; n4975
g2540 and n4974_not n4975 ; n4976
g2541 nor pi0062 n4883 ; n4977
g2542 and n4976_not n4977 ; n4978
g2543 and pi0246_not n3328 ; n4979
g2544 and n4879_not n4979 ; n4980
g2545 and n4978_not n4980 ; n4981
g2546 and n3447_not n4856 ; n4982
g2547 and n4871_not n4982 ; n4983
g2548 and n4850 n4983_not ; n4984
g2549 nor n4863 n4984 ; n4985
g2550 nor pi0215 n4985 ; n4986
g2551 nor n4848 n4986 ; n4987
g2552 and n3331 n4987 ; n4988
g2553 and n3556 n4849_not ; n4989
g2554 and n4866 n4989_not ; n4990
g2555 and n3331_not n4990 ; n4991
g2556 and pi0062 n4991_not ; n4992
g2557 and n4988_not n4992 ; n4993
g2558 nor n2537 n4990 ; n4994
g2559 and n2537 n4987_not ; n4995
g2560 and pi0056 n4994_not ; n4996
g2561 and n4995_not n4996 ; n4997
g2562 and n2572 n4987 ; n4998
g2563 and n2572_not n4990 ; n4999
g2564 and pi0055 n4999_not ; n5000
g2565 and n4998_not n5000 ; n5001
g2566 nor n3472 n4900 ; n5002
g2567 and pi0299 n4990_not ; n5003
g2568 and n5002 n5003_not ; n5004
g2569 and n2532_not n5004 ; n5005
g2570 and n2625_not n5004 ; n5006
g2571 and pi0299 n4987_not ; n5007
g2572 and n5002 n5007_not ; n5008
g2573 and n2625 n5008 ; n5009
g2574 nor n5006 n5009 ; n5010
g2575 and n2533 n5010_not ; n5011
g2576 and n2533_not n5004 ; n5012
g2577 and pi0092 n5012_not ; n5013
g2578 and n5011_not n5013 ; n5014
g2579 and pi0075 n5004 ; n5015
g2580 and pi0087 n5010 ; n5016
g2581 and pi0038 n5004 ; n5017
g2582 and pi0039 n5008_not ; n5018
g2583 and pi0877_not n3508 ; n5019
g2584 nor pi0169 n5019 ; n5020
g2585 nor pi0877 n3499 ; n5021
g2586 and pi0877 n3416_not ; n5022
g2587 and pi0169 n5021_not ; n5023
g2588 and n5022_not n5023 ; n5024
g2589 nor n5020 n5024 ; n5025
g2590 nor pi0228 n5025 ; n5026
g2591 and n3793_not n4856 ; n5027
g2592 and n5026_not n5027 ; n5028
g2593 and n4850 n5028_not ; n5029
g2594 nor n4863 n5029 ; n5030
g2595 nor pi0215 n5030 ; n5031
g2596 and n4923 n5031_not ; n5032
g2597 and n4943 n5032_not ; n5033
g2598 nor pi0038 n5018 ; n5034
g2599 and n5033_not n5034 ; n5035
g2600 nor pi0100 n5017 ; n5036
g2601 and n5035_not n5036 ; n5037
g2602 and n2530_not n5004 ; n5038
g2603 and n4954_not n4982 ; n5039
g2604 and n4850 n5039_not ; n5040
g2605 nor n4863 n5040 ; n5041
g2606 nor pi0215 n5041 ; n5042
g2607 nor n4848 n5042 ; n5043
g2608 and pi0299 n5043_not ; n5044
g2609 and n2530 n5002 ; n5045
g2610 and n5044_not n5045 ; n5046
g2611 and pi0100 n5038_not ; n5047
g2612 and n5046_not n5047 ; n5048
g2613 nor n5037 n5048 ; n5049
g2614 nor pi0087 n5049 ; n5050
g2615 nor pi0075 n5016 ; n5051
g2616 and n5050_not n5051 ; n5052
g2617 nor pi0092 n5015 ; n5053
g2618 and n5052_not n5053 ; n5054
g2619 and n2532 n5014_not ; n5055
g2620 and n5054_not n5055 ; n5056
g2621 nor pi0055 n5005 ; n5057
g2622 and n5056_not n5057 ; n5058
g2623 nor pi0056 n5001 ; n5059
g2624 and n5058_not n5059 ; n5060
g2625 nor pi0062 n4997 ; n5061
g2626 and n5060_not n5061 ; n5062
g2627 and pi0246 n3328 ; n5063
g2628 and n4993_not n5063 ; n5064
g2629 and n5062_not n5064 ; n5065
g2630 and pi0246 n4989 ; n5066
g2631 nor n3328 n5066 ; n5067
g2632 and n4866 n5067 ; n5068
g2633 nor n5065 n5068 ; n5069
g2634 and n4981_not n5069 ; po0161
g2635 and pi0215 pi1137 ; n5071
g2636 and pi0216 pi0280 ; n5072
g2637 nor pi0221 n5072 ; n5073
g2638 and pi0105_not pi0168 ; n5074
g2639 and pi0878 n2442_not ; n5075
g2640 and pi0105 n5075_not ; n5076
g2641 and pi0228 n5074_not ; n5077
g2642 and n5076_not n5077 ; n5078
g2643 nor pi0216 n5078 ; n5079
g2644 nor pi0168 pi0228 ; n5080
g2645 and n5079 n5080_not ; n5081
g2646 and n5073 n5081_not ; n5082
g2647 nor pi1137 n2452 ; n5083
g2648 and pi0933_not n2452 ; n5084
g2649 and pi0221 n5083_not ; n5085
g2650 and n5084_not n5085 ; n5086
g2651 nor n5082 n5086 ; n5087
g2652 nor pi0215 n5087 ; n5088
g2653 nor n5071 n5088 ; n5089
g2654 and n3331_not n5089 ; n5090
g2655 and pi0878_not n2521 ; n5091
g2656 and pi0168 n2521_not ; n5092
g2657 nor pi0228 n5091 ; n5093
g2658 and n5092_not n5093 ; n5094
g2659 and n5079 n5094_not ; n5095
g2660 and n5073 n5095_not ; n5096
g2661 nor n5086 n5096 ; n5097
g2662 nor pi0215 n5097 ; n5098
g2663 nor n5071 n5098 ; n5099
g2664 and n3331 n5099 ; n5100
g2665 and pi0062 n5090_not ; n5101
g2666 and n5100_not n5101 ; n5102
g2667 nor n2537 n5089 ; n5103
g2668 and n2537 n5099_not ; n5104
g2669 and pi0056 n5103_not ; n5105
g2670 and n5104_not n5105 ; n5106
g2671 and n2572_not n5089 ; n5107
g2672 and n2572 n5099 ; n5108
g2673 and pi0055 n5107_not ; n5109
g2674 and n5108_not n5109 ; n5110
g2675 and pi0223 pi1137 ; n5111
g2676 and pi0224 pi0280 ; n5112
g2677 nor pi0222 n5112 ; n5113
g2678 nor pi0224 n5075 ; n5114
g2679 and n5113 n5114_not ; n5115
g2680 nor pi1137 n2591 ; n5116
g2681 and pi0933_not n2591 ; n5117
g2682 and pi0222 n5116_not ; n5118
g2683 and n5117_not n5118 ; n5119
g2684 nor n5115 n5119 ; n5120
g2685 nor pi0223 n5120 ; n5121
g2686 nor n5111 n5121 ; n5122
g2687 nor pi0299 n5122 ; n5123
g2688 and pi0299 n5089_not ; n5124
g2689 nor n5123 n5124 ; n5125
g2690 and n2532_not n5125 ; n5126
g2691 and n2625_not n5125 ; n5127
g2692 and pi0299 n5099_not ; n5128
g2693 nor n5123 n5128 ; n5129
g2694 and n2625 n5129 ; n5130
g2695 nor n5127 n5130 ; n5131
g2696 and n2533 n5131_not ; n5132
g2697 and n2533_not n5125 ; n5133
g2698 and pi0092 n5133_not ; n5134
g2699 and n5132_not n5134 ; n5135
g2700 and pi0075 n5125 ; n5136
g2701 and pi0087 n5131 ; n5137
g2702 and pi0038 n5125 ; n5138
g2703 and pi0039 n5129_not ; n5139
g2704 nor pi0299 n5111 ; n5140
g2705 and pi0878 n3488 ; n5141
g2706 nor pi0224 n5141 ; n5142
g2707 and n5113 n5142_not ; n5143
g2708 nor n5119 n5143 ; n5144
g2709 and n5140 n5144 ; n5145
g2710 and pi0299 n5071_not ; n5146
g2711 and pi0878 n3499 ; n5147
g2712 nor pi0168 n5147 ; n5148
g2713 and pi0168 n3508 ; n5149
g2714 nor n5148 n5149 ; n5150
g2715 and pi0878 n5150_not ; n5151
g2716 and n3416_not n5148 ; n5152
g2717 nor n5151 n5152 ; n5153
g2718 nor pi0228 n5153 ; n5154
g2719 and n3497_not n5078 ; n5155
g2720 nor pi0216 n5155 ; n5156
g2721 and n5154_not n5156 ; n5157
g2722 and n5073 n5157_not ; n5158
g2723 nor n5086 n5158 ; n5159
g2724 nor pi0215 n5159 ; n5160
g2725 and n5146 n5160_not ; n5161
g2726 and n3488_not n5113 ; n5162
g2727 and n5144 n5162_not ; n5163
g2728 nor pi0223 n5163 ; n5164
g2729 and n5140 n5164_not ; n5165
g2730 nor pi0039 n5165 ; n5166
g2731 and n5145_not n5166 ; n5167
g2732 and n5161_not n5167 ; n5168
g2733 nor pi0038 n5139 ; n5169
g2734 and n5168_not n5169 ; n5170
g2735 nor pi0100 n5138 ; n5171
g2736 and n5170_not n5171 ; n5172
g2737 and n2530_not n5125 ; n5173
g2738 and pi0878_not n3394 ; n5174
g2739 and pi0168 n3394_not ; n5175
g2740 nor pi0228 n5174 ; n5176
g2741 and n5175_not n5176 ; n5177
g2742 and n5079 n5177_not ; n5178
g2743 and n5073 n5178_not ; n5179
g2744 nor n5086 n5179 ; n5180
g2745 nor pi0215 n5180 ; n5181
g2746 nor n5071 n5181 ; n5182
g2747 and pi0299 n5182_not ; n5183
g2748 and n2530 n5123_not ; n5184
g2749 and n5183_not n5184 ; n5185
g2750 and pi0100 n5173_not ; n5186
g2751 and n5185_not n5186 ; n5187
g2752 nor n5172 n5187 ; n5188
g2753 nor pi0087 n5188 ; n5189
g2754 nor pi0075 n5137 ; n5190
g2755 and n5189_not n5190 ; n5191
g2756 nor pi0092 n5136 ; n5192
g2757 and n5191_not n5192 ; n5193
g2758 and n2532 n5135_not ; n5194
g2759 and n5193_not n5194 ; n5195
g2760 nor pi0055 n5126 ; n5196
g2761 and n5195_not n5196 ; n5197
g2762 nor pi0056 n5110 ; n5198
g2763 and n5197_not n5198 ; n5199
g2764 nor pi0062 n5106 ; n5200
g2765 and n5199_not n5200 ; n5201
g2766 and pi0240_not n3328 ; n5202
g2767 and n5102_not n5202 ; n5203
g2768 and n5201_not n5203 ; n5204
g2769 and n3447_not n5079 ; n5205
g2770 and n5094_not n5205 ; n5206
g2771 and n5073 n5206_not ; n5207
g2772 nor n5086 n5207 ; n5208
g2773 nor pi0215 n5208 ; n5209
g2774 nor n5071 n5209 ; n5210
g2775 and n3331 n5210 ; n5211
g2776 and n3556 n5072_not ; n5212
g2777 and n5089 n5212_not ; n5213
g2778 and n3331_not n5213 ; n5214
g2779 and pi0062 n5214_not ; n5215
g2780 and n5211_not n5215 ; n5216
g2781 nor n2537 n5213 ; n5217
g2782 and n2537 n5210_not ; n5218
g2783 and pi0056 n5217_not ; n5219
g2784 and n5218_not n5219 ; n5220
g2785 and n2572 n5210 ; n5221
g2786 and n2572_not n5213 ; n5222
g2787 and pi0055 n5222_not ; n5223
g2788 and n5221_not n5223 ; n5224
g2789 nor n3472 n5123 ; n5225
g2790 and pi0299 n5213_not ; n5226
g2791 and n5225 n5226_not ; n5227
g2792 and n2532_not n5227 ; n5228
g2793 and n2625_not n5227 ; n5229
g2794 and pi0299 n5210_not ; n5230
g2795 and n5225 n5230_not ; n5231
g2796 and n2625 n5231 ; n5232
g2797 nor n5229 n5232 ; n5233
g2798 and n2533 n5233_not ; n5234
g2799 and n2533_not n5227 ; n5235
g2800 and pi0092 n5235_not ; n5236
g2801 and n5234_not n5236 ; n5237
g2802 and pi0075 n5227 ; n5238
g2803 and pi0087 n5233 ; n5239
g2804 and pi0038 n5227 ; n5240
g2805 and pi0039 n5231_not ; n5241
g2806 and pi0878_not n3508 ; n5242
g2807 nor pi0168 n5242 ; n5243
g2808 nor pi0878 n3499 ; n5244
g2809 and pi0878 n3416_not ; n5245
g2810 and pi0168 n5244_not ; n5246
g2811 and n5245_not n5246 ; n5247
g2812 nor n5243 n5247 ; n5248
g2813 nor pi0228 n5248 ; n5249
g2814 and n3793_not n5079 ; n5250
g2815 and n5249_not n5250 ; n5251
g2816 and n5073 n5251_not ; n5252
g2817 nor n5086 n5252 ; n5253
g2818 nor pi0215 n5253 ; n5254
g2819 and n5146 n5254_not ; n5255
g2820 and n5166 n5255_not ; n5256
g2821 nor pi0038 n5241 ; n5257
g2822 and n5256_not n5257 ; n5258
g2823 nor pi0100 n5240 ; n5259
g2824 and n5258_not n5259 ; n5260
g2825 and n2530_not n5227 ; n5261
g2826 and n5177_not n5205 ; n5262
g2827 and n5073 n5262_not ; n5263
g2828 nor n5086 n5263 ; n5264
g2829 nor pi0215 n5264 ; n5265
g2830 nor n5071 n5265 ; n5266
g2831 and pi0299 n5266_not ; n5267
g2832 and n2530 n5225 ; n5268
g2833 and n5267_not n5268 ; n5269
g2834 and pi0100 n5261_not ; n5270
g2835 and n5269_not n5270 ; n5271
g2836 nor n5260 n5271 ; n5272
g2837 nor pi0087 n5272 ; n5273
g2838 nor pi0075 n5239 ; n5274
g2839 and n5273_not n5274 ; n5275
g2840 nor pi0092 n5238 ; n5276
g2841 and n5275_not n5276 ; n5277
g2842 and n2532 n5237_not ; n5278
g2843 and n5277_not n5278 ; n5279
g2844 nor pi0055 n5228 ; n5280
g2845 and n5279_not n5280 ; n5281
g2846 nor pi0056 n5224 ; n5282
g2847 and n5281_not n5282 ; n5283
g2848 nor pi0062 n5220 ; n5284
g2849 and n5283_not n5284 ; n5285
g2850 and pi0240 n3328 ; n5286
g2851 and n5216_not n5286 ; n5287
g2852 and n5285_not n5287 ; n5288
g2853 and pi0240 n5212 ; n5289
g2854 nor n3328 n5289 ; n5290
g2855 and n5089 n5290 ; n5291
g2856 nor n5288 n5291 ; n5292
g2857 and n5204_not n5292 ; po0162
g2858 and pi0215 pi1136 ; n5294
g2859 and pi0216 pi0266 ; n5295
g2860 and pi0875 n2442_not ; n5296
g2861 and pi0105 n5296_not ; n5297
g2862 nor pi0105 pi0166 ; n5298
g2863 nor n5297 n5298 ; n5299
g2864 and pi0228 n5299 ; n5300
g2865 and pi0166 pi0228_not ; n5301
g2866 nor n5300 n5301 ; n5302
g2867 nor pi0216 n5302 ; n5303
g2868 nor n5295 n5303 ; n5304
g2869 nor pi0221 n5304 ; n5305
g2870 nor pi1136 n2452 ; n5306
g2871 and pi0928_not n2452 ; n5307
g2872 and pi0221 n5306_not ; n5308
g2873 and n5307_not n5308 ; n5309
g2874 nor n5305 n5309 ; n5310
g2875 nor pi0215 n5310 ; n5311
g2876 nor n5294 n5311 ; n5312
g2877 and n3328_not n5312 ; n5313
g2878 and n3331_not n5312 ; n5314
g2879 nor pi0166 n2521 ; n5315
g2880 and pi0875_not n2521 ; n5316
g2881 nor pi0228 n5315 ; n5317
g2882 and n5316_not n5317 ; n5318
g2883 nor n5300 n5318 ; n5319
g2884 nor pi0216 n5319 ; n5320
g2885 nor n5295 n5320 ; n5321
g2886 nor pi0221 n5321 ; n5322
g2887 nor n5309 n5322 ; n5323
g2888 nor pi0215 n5323 ; n5324
g2889 nor n5294 n5324 ; n5325
g2890 and n3331 n5325 ; n5326
g2891 and pi0062 n5314_not ; n5327
g2892 and n5326_not n5327 ; n5328
g2893 nor n2537 n5312 ; n5329
g2894 and n2537 n5325_not ; n5330
g2895 and pi0056 n5329_not ; n5331
g2896 and n5330_not n5331 ; n5332
g2897 and n2572_not n5312 ; n5333
g2898 and n2572 n5325 ; n5334
g2899 and pi0055 n5333_not ; n5335
g2900 and n5334_not n5335 ; n5336
g2901 and pi0223 pi1136 ; n5337
g2902 and pi0224 pi0266_not ; n5338
g2903 nor pi0224 pi0875 ; n5339
g2904 and n2442_not n5339 ; n5340
g2905 nor pi0222 n5338 ; n5341
g2906 and n5340_not n5341 ; n5342
g2907 nor pi1136 n2591 ; n5343
g2908 and pi0928_not n2591 ; n5344
g2909 and pi0222 n5343_not ; n5345
g2910 and n5344_not n5345 ; n5346
g2911 nor n5342 n5346 ; n5347
g2912 nor pi0223 n5347 ; n5348
g2913 nor n5337 n5348 ; n5349
g2914 nor pi0299 n5349 ; n5350
g2915 and n2604 n5296_not ; n5351
g2916 and n5350 n5351_not ; n5352
g2917 and pi0299 n5312_not ; n5353
g2918 nor n5352 n5353 ; n5354
g2919 and n2532_not n5354 ; n5355
g2920 and n2625_not n5354 ; n5356
g2921 and pi0299 n5325_not ; n5357
g2922 nor n5352 n5357 ; n5358
g2923 and n2625 n5358 ; n5359
g2924 nor n5356 n5359 ; n5360
g2925 and n2533 n5360_not ; n5361
g2926 and n2533_not n5354 ; n5362
g2927 and pi0092 n5362_not ; n5363
g2928 and n5361_not n5363 ; n5364
g2929 and pi0075 n5354 ; n5365
g2930 and pi0087 n5360 ; n5366
g2931 and pi0038 n5354 ; n5367
g2932 and pi0039 n5358_not ; n5368
g2933 and n2603 n3488_not ; n5369
g2934 and n5342 n5369_not ; n5370
g2935 nor pi0299 n5337 ; n5371
g2936 and n5346_not n5371 ; n5372
g2937 and n5370_not n5372 ; n5373
g2938 and n3498 n5299_not ; n5374
g2939 nor pi0216 n5374 ; n5375
g2940 and pi0166 n3499 ; n5376
g2941 nor pi0166 n3508 ; n5377
g2942 and pi0875 n5376_not ; n5378
g2943 and n5377_not n5378 ; n5379
g2944 and pi0166 pi0875_not ; n5380
g2945 and n3416_not n5380 ; n5381
g2946 nor n5379 n5381 ; n5382
g2947 nor pi0228 n5382 ; n5383
g2948 nor n3498 n5383 ; n5384
g2949 and n5375 n5384_not ; n5385
g2950 nor n5295 n5385 ; n5386
g2951 nor pi0221 n5386 ; n5387
g2952 nor n5309 n5387 ; n5388
g2953 nor pi0215 n5388 ; n5389
g2954 and pi0299 n5294_not ; n5390
g2955 and n5389_not n5390 ; n5391
g2956 and n5347 n5369_not ; n5392
g2957 nor pi0223 n5392 ; n5393
g2958 and n5371 n5393_not ; n5394
g2959 nor pi0039 n5394 ; n5395
g2960 and n5373_not n5395 ; n5396
g2961 and n5391_not n5396 ; n5397
g2962 nor pi0038 n5368 ; n5398
g2963 and n5397_not n5398 ; n5399
g2964 nor pi0100 n5367 ; n5400
g2965 and n5399_not n5400 ; n5401
g2966 and n2530_not n5354 ; n5402
g2967 and pi0875_not n3387 ; n5403
g2968 and pi0166 n5403_not ; n5404
g2969 nor n2638 n3387 ; n5405
g2970 and n2638 n3385_not ; n5406
g2971 and pi0875 n5406_not ; n5407
g2972 and n5405_not n5407 ; n5408
g2973 nor n5404 n5408 ; n5409
g2974 nor pi0228 n5409 ; n5410
g2975 nor n5300 n5410 ; n5411
g2976 nor pi0216 n5411 ; n5412
g2977 nor n5295 n5412 ; n5413
g2978 nor pi0221 n5413 ; n5414
g2979 nor n5309 n5414 ; n5415
g2980 nor pi0215 n5415 ; n5416
g2981 nor n5294 n5416 ; n5417
g2982 and pi0299 n5417_not ; n5418
g2983 and n2530 n5352_not ; n5419
g2984 and n5418_not n5419 ; n5420
g2985 and pi0100 n5402_not ; n5421
g2986 and n5420_not n5421 ; n5422
g2987 nor n5401 n5422 ; n5423
g2988 nor pi0087 n5423 ; n5424
g2989 nor pi0075 n5366 ; n5425
g2990 and n5424_not n5425 ; n5426
g2991 nor pi0092 n5365 ; n5427
g2992 and n5426_not n5427 ; n5428
g2993 and n2532 n5364_not ; n5429
g2994 and n5428_not n5429 ; n5430
g2995 nor pi0055 n5355 ; n5431
g2996 and n5430_not n5431 ; n5432
g2997 nor pi0056 n5336 ; n5433
g2998 and n5432_not n5433 ; n5434
g2999 nor pi0062 n5332 ; n5435
g3000 and n5434_not n5435 ; n5436
g3001 and n3328 n5328_not ; n5437
g3002 and n5436_not n5437 ; n5438
g3003 nor pi0245 n5313 ; n5439
g3004 and n5438_not n5439 ; n5440
g3005 and n3450_not n5312 ; n5441
g3006 and n3328_not n5441 ; n5442
g3007 nor n3447 n5300 ; n5443
g3008 and n5318_not n5443 ; n5444
g3009 nor pi0216 n5444 ; n5445
g3010 nor n5295 n5445 ; n5446
g3011 nor pi0221 n5446 ; n5447
g3012 nor n5309 n5447 ; n5448
g3013 nor pi0215 n5448 ; n5449
g3014 nor n5294 n5449 ; n5450
g3015 and n3331 n5450 ; n5451
g3016 and n3331_not n5441 ; n5452
g3017 and pi0062 n5452_not ; n5453
g3018 and n5451_not n5453 ; n5454
g3019 nor n2537 n5441 ; n5455
g3020 and n2537 n5450_not ; n5456
g3021 and pi0056 n5455_not ; n5457
g3022 and n5456_not n5457 ; n5458
g3023 and n2572 n5450 ; n5459
g3024 and n2572_not n5441 ; n5460
g3025 and pi0055 n5460_not ; n5461
g3026 and n5459_not n5461 ; n5462
g3027 and pi0299 n5441_not ; n5463
g3028 nor n5350 n5463 ; n5464
g3029 and n2532_not n5464 ; n5465
g3030 and n2625_not n5464 ; n5466
g3031 and pi0299 n5450_not ; n5467
g3032 nor n5350 n5467 ; n5468
g3033 and n2625 n5468 ; n5469
g3034 nor n5466 n5469 ; n5470
g3035 and n2533 n5470_not ; n5471
g3036 and n2533_not n5464 ; n5472
g3037 and pi0092 n5472_not ; n5473
g3038 and n5471_not n5473 ; n5474
g3039 and pi0075 n5464 ; n5475
g3040 and pi0087 n5470 ; n5476
g3041 and pi0038 n5464 ; n5477
g3042 and pi0039 n5468_not ; n5478
g3043 nor pi0166 n3499 ; n5479
g3044 and pi0166 n3508 ; n5480
g3045 nor pi0875 n5479 ; n5481
g3046 and n5480_not n5481 ; n5482
g3047 nor pi0166 n3416 ; n5483
g3048 and pi0875 n5483_not ; n5484
g3049 nor pi0228 n5482 ; n5485
g3050 and n5484_not n5485 ; n5486
g3051 and n5375 n5486_not ; n5487
g3052 nor n5295 n5487 ; n5488
g3053 nor pi0221 n5488 ; n5489
g3054 nor n5309 n5489 ; n5490
g3055 nor pi0215 n5490 ; n5491
g3056 and n5390 n5491_not ; n5492
g3057 and n5395 n5492_not ; n5493
g3058 nor pi0038 n5478 ; n5494
g3059 and n5493_not n5494 ; n5495
g3060 nor pi0100 n5477 ; n5496
g3061 and n5495_not n5496 ; n5497
g3062 and n2530_not n5464 ; n5498
g3063 and n5410_not n5443 ; n5499
g3064 nor pi0216 n5499 ; n5500
g3065 nor n5295 n5500 ; n5501
g3066 nor pi0221 n5501 ; n5502
g3067 nor n5309 n5502 ; n5503
g3068 nor pi0215 n5503 ; n5504
g3069 nor n5294 n5504 ; n5505
g3070 and pi0299 n5505_not ; n5506
g3071 and n2530 n5350_not ; n5507
g3072 and n5506_not n5507 ; n5508
g3073 and pi0100 n5498_not ; n5509
g3074 and n5508_not n5509 ; n5510
g3075 nor n5497 n5510 ; n5511
g3076 nor pi0087 n5511 ; n5512
g3077 nor pi0075 n5476 ; n5513
g3078 and n5512_not n5513 ; n5514
g3079 nor pi0092 n5475 ; n5515
g3080 and n5514_not n5515 ; n5516
g3081 and n2532 n5474_not ; n5517
g3082 and n5516_not n5517 ; n5518
g3083 nor pi0055 n5465 ; n5519
g3084 and n5518_not n5519 ; n5520
g3085 nor pi0056 n5462 ; n5521
g3086 and n5520_not n5521 ; n5522
g3087 nor pi0062 n5458 ; n5523
g3088 and n5522_not n5523 ; n5524
g3089 and n3328 n5454_not ; n5525
g3090 and n5524_not n5525 ; n5526
g3091 and pi0245 n5442_not ; n5527
g3092 and n5526_not n5527 ; n5528
g3093 or n5440 n5528 ; po0163
g3094 and pi0215 pi1135 ; n5530
g3095 and pi0216 pi0279 ; n5531
g3096 and pi0879 n2442_not ; n5532
g3097 and pi0105 n5532_not ; n5533
g3098 nor pi0105 pi0161 ; n5534
g3099 nor n5533 n5534 ; n5535
g3100 and pi0228 n5535 ; n5536
g3101 and pi0161 pi0228_not ; n5537
g3102 nor n5536 n5537 ; n5538
g3103 nor pi0216 n5538 ; n5539
g3104 nor n5531 n5539 ; n5540
g3105 nor pi0221 n5540 ; n5541
g3106 nor pi1135 n2452 ; n5542
g3107 and pi0938_not n2452 ; n5543
g3108 and pi0221 n5542_not ; n5544
g3109 and n5543_not n5544 ; n5545
g3110 nor n5541 n5545 ; n5546
g3111 nor pi0215 n5546 ; n5547
g3112 nor n5530 n5547 ; n5548
g3113 and n3328_not n5548 ; n5549
g3114 and n3331_not n5548 ; n5550
g3115 and pi0879_not n2521 ; n5551
g3116 nor n3335 n5537 ; n5552
g3117 nor n5551 n5552 ; n5553
g3118 nor n5536 n5553 ; n5554
g3119 nor pi0216 n5554 ; n5555
g3120 nor n5531 n5555 ; n5556
g3121 nor pi0221 n5556 ; n5557
g3122 nor n5545 n5557 ; n5558
g3123 nor pi0215 n5558 ; n5559
g3124 nor n5530 n5559 ; n5560
g3125 and n3331 n5560 ; n5561
g3126 and pi0062 n5550_not ; n5562
g3127 and n5561_not n5562 ; n5563
g3128 nor n2537 n5548 ; n5564
g3129 and n2537 n5560_not ; n5565
g3130 and pi0056 n5564_not ; n5566
g3131 and n5565_not n5566 ; n5567
g3132 and n2572_not n5548 ; n5568
g3133 and n2572 n5560 ; n5569
g3134 and pi0055 n5568_not ; n5570
g3135 and n5569_not n5570 ; n5571
g3136 and pi0223 pi1135 ; n5572
g3137 nor pi1135 n2591 ; n5573
g3138 and pi0938_not n2591 ; n5574
g3139 and pi0222 n5573_not ; n5575
g3140 and n5574_not n5575 ; n5576
g3141 and pi0224 pi0279_not ; n5577
g3142 nor pi0224 pi0879 ; n5578
g3143 and n2442_not n5578 ; n5579
g3144 nor pi0222 n5577 ; n5580
g3145 and n5579_not n5580 ; n5581
g3146 nor n5576 n5581 ; n5582
g3147 nor pi0223 n5582 ; n5583
g3148 nor n5572 n5583 ; n5584
g3149 nor pi0299 n5584 ; n5585
g3150 and n2604 n5532_not ; n5586
g3151 and n5585 n5586_not ; n5587
g3152 and pi0299 n5548_not ; n5588
g3153 nor n5587 n5588 ; n5589
g3154 and n2532_not n5589 ; n5590
g3155 and n2625_not n5589 ; n5591
g3156 and pi0299 n5560_not ; n5592
g3157 nor n5587 n5592 ; n5593
g3158 and n2625 n5593 ; n5594
g3159 nor n5591 n5594 ; n5595
g3160 and n2533 n5595_not ; n5596
g3161 and n2533_not n5589 ; n5597
g3162 and pi0092 n5597_not ; n5598
g3163 and n5596_not n5598 ; n5599
g3164 and pi0075 n5589 ; n5600
g3165 and pi0087 n5595 ; n5601
g3166 and pi0038 n5589 ; n5602
g3167 and pi0039 n5593_not ; n5603
g3168 nor pi0299 n5572 ; n5604
g3169 and n5369 n5576_not ; n5605
g3170 and n5583 n5605_not ; n5606
g3171 and n5604 n5606_not ; n5607
g3172 and n3498 n5535_not ; n5608
g3173 nor pi0216 n5608 ; n5609
g3174 and pi0161 n3499 ; n5610
g3175 nor pi0161 n3508 ; n5611
g3176 and pi0879 n5610_not ; n5612
g3177 and n5611_not n5612 ; n5613
g3178 and pi0161 pi0879_not ; n5614
g3179 and n3416_not n5614 ; n5615
g3180 nor n5613 n5615 ; n5616
g3181 nor pi0228 n5616 ; n5617
g3182 nor n3498 n5617 ; n5618
g3183 and n5609 n5618_not ; n5619
g3184 nor n5531 n5619 ; n5620
g3185 nor pi0221 n5620 ; n5621
g3186 nor n5545 n5621 ; n5622
g3187 nor pi0215 n5622 ; n5623
g3188 and pi0299 n5530_not ; n5624
g3189 and n5623_not n5624 ; n5625
g3190 nor pi0039 n5607 ; n5626
g3191 and n5625_not n5626 ; n5627
g3192 nor pi0038 n5603 ; n5628
g3193 and n5627_not n5628 ; n5629
g3194 nor pi0100 n5602 ; n5630
g3195 and n5629_not n5630 ; n5631
g3196 and n2530_not n5589 ; n5632
g3197 and pi0879_not n3387 ; n5633
g3198 and pi0161 n5633_not ; n5634
g3199 nor pi0152 pi0166 ; n5635
g3200 and n3385_not n5635 ; n5636
g3201 nor n3387 n5635 ; n5637
g3202 and pi0879 n5636_not ; n5638
g3203 and n5637_not n5638 ; n5639
g3204 nor n5634 n5639 ; n5640
g3205 nor pi0228 n5640 ; n5641
g3206 nor n5536 n5641 ; n5642
g3207 nor pi0216 n5642 ; n5643
g3208 nor n5531 n5643 ; n5644
g3209 nor pi0221 n5644 ; n5645
g3210 nor n5545 n5645 ; n5646
g3211 nor pi0215 n5646 ; n5647
g3212 nor n5530 n5647 ; n5648
g3213 and pi0299 n5648_not ; n5649
g3214 and n2530 n5587_not ; n5650
g3215 and n5649_not n5650 ; n5651
g3216 and pi0100 n5632_not ; n5652
g3217 and n5651_not n5652 ; n5653
g3218 nor n5631 n5653 ; n5654
g3219 nor pi0087 n5654 ; n5655
g3220 nor pi0075 n5601 ; n5656
g3221 and n5655_not n5656 ; n5657
g3222 nor pi0092 n5600 ; n5658
g3223 and n5657_not n5658 ; n5659
g3224 and n2532 n5599_not ; n5660
g3225 and n5659_not n5660 ; n5661
g3226 nor pi0055 n5590 ; n5662
g3227 and n5661_not n5662 ; n5663
g3228 nor pi0056 n5571 ; n5664
g3229 and n5663_not n5664 ; n5665
g3230 nor pi0062 n5567 ; n5666
g3231 and n5665_not n5666 ; n5667
g3232 and n3328 n5563_not ; n5668
g3233 and n5667_not n5668 ; n5669
g3234 nor pi0244 n5549 ; n5670
g3235 and n5669_not n5670 ; n5671
g3236 and n3450_not n5548 ; n5672
g3237 and n3328_not n5672 ; n5673
g3238 nor n3447 n5536 ; n5674
g3239 and n5553_not n5674 ; n5675
g3240 nor pi0216 n5675 ; n5676
g3241 nor n5531 n5676 ; n5677
g3242 nor pi0221 n5677 ; n5678
g3243 nor n5545 n5678 ; n5679
g3244 nor pi0215 n5679 ; n5680
g3245 nor n5530 n5680 ; n5681
g3246 and n3331 n5681 ; n5682
g3247 and n3331_not n5672 ; n5683
g3248 and pi0062 n5683_not ; n5684
g3249 and n5682_not n5684 ; n5685
g3250 nor n2537 n5672 ; n5686
g3251 and n2537 n5681_not ; n5687
g3252 and pi0056 n5686_not ; n5688
g3253 and n5687_not n5688 ; n5689
g3254 and n2572 n5681 ; n5690
g3255 and n2572_not n5672 ; n5691
g3256 and pi0055 n5691_not ; n5692
g3257 and n5690_not n5692 ; n5693
g3258 and pi0299 n5672_not ; n5694
g3259 nor n5585 n5694 ; n5695
g3260 and n2532_not n5695 ; n5696
g3261 and n2625_not n5695 ; n5697
g3262 and pi0299 n5681_not ; n5698
g3263 nor n5585 n5698 ; n5699
g3264 and n2625 n5699 ; n5700
g3265 nor n5697 n5700 ; n5701
g3266 and n2533 n5701_not ; n5702
g3267 and n2533_not n5695 ; n5703
g3268 and pi0092 n5703_not ; n5704
g3269 and n5702_not n5704 ; n5705
g3270 and pi0075 n5695 ; n5706
g3271 and pi0087 n5701 ; n5707
g3272 and pi0038 n5695 ; n5708
g3273 and pi0039 n5699_not ; n5709
g3274 and n5369_not n5582 ; n5710
g3275 nor pi0223 n5710 ; n5711
g3276 and n5604 n5711_not ; n5712
g3277 nor pi0161 n3499 ; n5713
g3278 and pi0161 n3508 ; n5714
g3279 nor pi0879 n5713 ; n5715
g3280 and n5714_not n5715 ; n5716
g3281 nor pi0161 n3416 ; n5717
g3282 and pi0879 n5717_not ; n5718
g3283 nor pi0228 n5716 ; n5719
g3284 and n5718_not n5719 ; n5720
g3285 and n5609 n5720_not ; n5721
g3286 nor n5531 n5721 ; n5722
g3287 nor pi0221 n5722 ; n5723
g3288 nor n5545 n5723 ; n5724
g3289 nor pi0215 n5724 ; n5725
g3290 and n5624 n5725_not ; n5726
g3291 nor pi0039 n5712 ; n5727
g3292 and n5726_not n5727 ; n5728
g3293 nor pi0038 n5709 ; n5729
g3294 and n5728_not n5729 ; n5730
g3295 nor pi0100 n5708 ; n5731
g3296 and n5730_not n5731 ; n5732
g3297 and n2530_not n5695 ; n5733
g3298 and n5641_not n5674 ; n5734
g3299 nor pi0216 n5734 ; n5735
g3300 nor n5531 n5735 ; n5736
g3301 nor pi0221 n5736 ; n5737
g3302 nor n5545 n5737 ; n5738
g3303 nor pi0215 n5738 ; n5739
g3304 nor n5530 n5739 ; n5740
g3305 and pi0299 n5740_not ; n5741
g3306 and n2530 n5585_not ; n5742
g3307 and n5741_not n5742 ; n5743
g3308 and pi0100 n5733_not ; n5744
g3309 and n5743_not n5744 ; n5745
g3310 nor n5732 n5745 ; n5746
g3311 nor pi0087 n5746 ; n5747
g3312 nor pi0075 n5707 ; n5748
g3313 and n5747_not n5748 ; n5749
g3314 nor pi0092 n5706 ; n5750
g3315 and n5749_not n5750 ; n5751
g3316 and n2532 n5705_not ; n5752
g3317 and n5751_not n5752 ; n5753
g3318 nor pi0055 n5696 ; n5754
g3319 and n5753_not n5754 ; n5755
g3320 nor pi0056 n5693 ; n5756
g3321 and n5755_not n5756 ; n5757
g3322 nor pi0062 n5689 ; n5758
g3323 and n5757_not n5758 ; n5759
g3324 and n3328 n5685_not ; n5760
g3325 and n5759_not n5760 ; n5761
g3326 and pi0244 n5673_not ; n5762
g3327 and n5761_not n5762 ; n5763
g3328 or n5671 n5763 ; po0164
g3329 and pi0216 pi0278 ; n5765
g3330 nor pi0221 n5765 ; n5766
g3331 and pi0105_not pi0152 ; n5767
g3332 and pi0846 n2442_not ; n5768
g3333 and pi0105 n5768 ; n5769
g3334 nor n5767 n5769 ; n5770
g3335 and pi0228 n5770_not ; n5771
g3336 and pi0152 pi0228_not ; n5772
g3337 nor n5771 n5772 ; n5773
g3338 nor pi0216 n5773 ; n5774
g3339 and n5766 n5774_not ; n5775
g3340 and pi0833 pi0930_not ; n5776
g3341 and pi0216_not pi0221 ; n5777
g3342 and n5776 n5777 ; n5778
g3343 and pi0221 n2452_not ; n5779
g3344 nor pi0215 n5779 ; n5780
g3345 and n5778_not n5780 ; n5781
g3346 and n5775_not n5781 ; n5782
g3347 nor n3450 n5782 ; n5783
g3348 nor n3328 n5783 ; n5784
g3349 nor n3331 n5783 ; n5785
g3350 nor n3447 n5771 ; n5786
g3351 nor pi0152 n2521 ; n5787
g3352 and pi0846_not n2521 ; n5788
g3353 nor pi0228 n5787 ; n5789
g3354 and n5788_not n5789 ; n5790
g3355 and n5786 n5790_not ; n5791
g3356 nor pi0216 n5791 ; n5792
g3357 and n5766 n5792_not ; n5793
g3358 and n5781 n5793_not ; n5794
g3359 and n3331 n5794 ; n5795
g3360 and pi0062 n5785_not ; n5796
g3361 and n5795_not n5796 ; n5797
g3362 and n2537 n5794_not ; n5798
g3363 and n2537_not n5783 ; n5799
g3364 and pi0056 n5799_not ; n5800
g3365 and n5798_not n5800 ; n5801
g3366 nor n2572 n5783 ; n5802
g3367 and n2572 n5794 ; n5803
g3368 and pi0055 n5802_not ; n5804
g3369 and n5803_not n5804 ; n5805
g3370 and pi0224 pi0278 ; n5806
g3371 nor pi0222 n5806 ; n5807
g3372 and pi0224_not n5768 ; n5808
g3373 and n5807 n5808_not ; n5809
g3374 and pi0222 pi0224_not ; n5810
g3375 and n5776 n5810 ; n5811
g3376 and n2593 n5811_not ; n5812
g3377 and n5809_not n5812 ; n5813
g3378 nor pi0299 n5813 ; n5814
g3379 and n3755_not n5814 ; n5815
g3380 and pi0299 n5783 ; n5816
g3381 nor n5815 n5816 ; n5817
g3382 and n2532_not n5817 ; n5818
g3383 and n2625_not n5817 ; n5819
g3384 and pi0299 n5794_not ; n5820
g3385 nor n5815 n5820 ; n5821
g3386 and n2625 n5821 ; n5822
g3387 nor n5819 n5822 ; n5823
g3388 and n2533 n5823_not ; n5824
g3389 and n2533_not n5817 ; n5825
g3390 and pi0092 n5825_not ; n5826
g3391 and n5824_not n5826 ; n5827
g3392 and pi0075 n5817 ; n5828
g3393 and pi0087 n5823 ; n5829
g3394 and pi0038 n5817 ; n5830
g3395 and pi0039 n5821_not ; n5831
g3396 and pi0846_not n3488 ; n5832
g3397 nor pi0224 n5832 ; n5833
g3398 and n5807 n5833_not ; n5834
g3399 nor n5811 n5834 ; n5835
g3400 and n2592_not n3470 ; n5836
g3401 and n5835 n5836 ; n5837
g3402 and pi0228 n5767_not ; n5838
g3403 and pi0105 n5832_not ; n5839
g3404 and n5838 n5839_not ; n5840
g3405 nor pi0216 n5840 ; n5841
g3406 and pi0152_not n3499 ; n5842
g3407 and pi0152 n3508_not ; n5843
g3408 nor pi0846 n5842 ; n5844
g3409 and n5843_not n5844 ; n5845
g3410 and pi0152_not pi0846 ; n5846
g3411 and n3416_not n5846 ; n5847
g3412 nor n5845 n5847 ; n5848
g3413 nor pi0228 n5848 ; n5849
g3414 and n5841 n5849_not ; n5850
g3415 and n5766 n5850_not ; n5851
g3416 nor n5778 n5851 ; n5852
g3417 and pi0215_not pi0299 ; n5853
g3418 and n5779_not n5853 ; n5854
g3419 and n5852 n5854 ; n5855
g3420 nor pi0039 n5837 ; n5856
g3421 and n5855_not n5856 ; n5857
g3422 nor pi0038 n5831 ; n5858
g3423 and n5857_not n5858 ; n5859
g3424 nor pi0100 n5830 ; n5860
g3425 and n5859_not n5860 ; n5861
g3426 and n2530_not n5817 ; n5862
g3427 and pi0846 n3393_not ; n5863
g3428 nor n3388 n5863 ; n5864
g3429 nor pi0228 n5864 ; n5865
g3430 and n5786 n5865_not ; n5866
g3431 nor pi0216 n5866 ; n5867
g3432 and n5766 n5867_not ; n5868
g3433 and n5781 n5868_not ; n5869
g3434 and pi0299 n5869_not ; n5870
g3435 and n2530 n5815_not ; n5871
g3436 and n5870_not n5871 ; n5872
g3437 and pi0100 n5862_not ; n5873
g3438 and n5872_not n5873 ; n5874
g3439 nor n5861 n5874 ; n5875
g3440 nor pi0087 n5875 ; n5876
g3441 nor pi0075 n5829 ; n5877
g3442 and n5876_not n5877 ; n5878
g3443 nor pi0092 n5828 ; n5879
g3444 and n5878_not n5879 ; n5880
g3445 and n2532 n5827_not ; n5881
g3446 and n5880_not n5881 ; n5882
g3447 nor pi0055 n5818 ; n5883
g3448 and n5882_not n5883 ; n5884
g3449 nor pi0056 n5805 ; n5885
g3450 and n5884_not n5885 ; n5886
g3451 nor pi0062 n5801 ; n5887
g3452 and n5886_not n5887 ; n5888
g3453 and n3328 n5797_not ; n5889
g3454 and n5888_not n5889 ; n5890
g3455 and pi0242 n5784_not ; n5891
g3456 and n5890_not n5891 ; n5892
g3457 and n3328_not n5782 ; n5893
g3458 and n3331_not n5782 ; n5894
g3459 nor n5771 n5790 ; n5895
g3460 nor pi0216 n5895 ; n5896
g3461 and n5766 n5896_not ; n5897
g3462 and n5781 n5897_not ; n5898
g3463 and n3331 n5898 ; n5899
g3464 and pi0062 n5894_not ; n5900
g3465 and n5899_not n5900 ; n5901
g3466 nor n2537 n5782 ; n5902
g3467 and n2537 n5898_not ; n5903
g3468 and pi0056 n5902_not ; n5904
g3469 and n5903_not n5904 ; n5905
g3470 and n2572_not n5782 ; n5906
g3471 and n2572 n5898 ; n5907
g3472 and pi0055 n5906_not ; n5908
g3473 and n5907_not n5908 ; n5909
g3474 and pi0299 n5782_not ; n5910
g3475 nor n5814 n5910 ; n5911
g3476 and n2532_not n5911 ; n5912
g3477 and n2625_not n5911 ; n5913
g3478 and pi0299 n5898_not ; n5914
g3479 nor n5814 n5914 ; n5915
g3480 and n2625 n5915 ; n5916
g3481 nor n5913 n5916 ; n5917
g3482 and n2533 n5917_not ; n5918
g3483 and n2533_not n5911 ; n5919
g3484 and pi0092 n5919_not ; n5920
g3485 and n5918_not n5920 ; n5921
g3486 and pi0075 n5911 ; n5922
g3487 and pi0087 n5917 ; n5923
g3488 and pi0038 n5911 ; n5924
g3489 and pi0039 n5915_not ; n5925
g3490 and n3487_not n5808 ; n5926
g3491 and n5807 n5926_not ; n5927
g3492 and n5811_not n5836 ; n5928
g3493 and n5927_not n5928 ; n5929
g3494 and n3488_not n5838 ; n5930
g3495 and pi0152 pi0846_not ; n5931
g3496 and n3416_not n5931 ; n5932
g3497 and pi0152 n3499 ; n5933
g3498 nor pi0152 n3508 ; n5934
g3499 and pi0846 n5933_not ; n5935
g3500 and n5934_not n5935 ; n5936
g3501 nor pi0228 n5932 ; n5937
g3502 and n5936_not n5937 ; n5938
g3503 and n5841 n5930_not ; n5939
g3504 and n5938_not n5939 ; n5940
g3505 and n5766 n5940_not ; n5941
g3506 nor n5778 n5941 ; n5942
g3507 and n5854 n5942 ; n5943
g3508 nor pi0039 n5929 ; n5944
g3509 and n5943_not n5944 ; n5945
g3510 nor pi0038 n5925 ; n5946
g3511 and n5945_not n5946 ; n5947
g3512 nor pi0100 n5924 ; n5948
g3513 and n5947_not n5948 ; n5949
g3514 and n2530_not n5911 ; n5950
g3515 nor n5771 n5865 ; n5951
g3516 nor pi0216 n5951 ; n5952
g3517 and n5766 n5952_not ; n5953
g3518 and n5781 n5953_not ; n5954
g3519 and pi0299 n5954_not ; n5955
g3520 and n2530 n5814_not ; n5956
g3521 and n5955_not n5956 ; n5957
g3522 and pi0100 n5950_not ; n5958
g3523 and n5957_not n5958 ; n5959
g3524 nor n5949 n5959 ; n5960
g3525 nor pi0087 n5960 ; n5961
g3526 nor pi0075 n5923 ; n5962
g3527 and n5961_not n5962 ; n5963
g3528 nor pi0092 n5922 ; n5964
g3529 and n5963_not n5964 ; n5965
g3530 and n2532 n5921_not ; n5966
g3531 and n5965_not n5966 ; n5967
g3532 nor pi0055 n5912 ; n5968
g3533 and n5967_not n5968 ; n5969
g3534 nor pi0056 n5909 ; n5970
g3535 and n5969_not n5970 ; n5971
g3536 nor pi0062 n5905 ; n5972
g3537 and n5971_not n5972 ; n5973
g3538 and n3328 n5901_not ; n5974
g3539 and n5973_not n5974 ; n5975
g3540 nor pi0242 n5893 ; n5976
g3541 and n5975_not n5976 ; n5977
g3542 nor n5892 n5977 ; n5978
g3543 nor pi1134 n5978 ; n5979
g3544 nor n5775 n5778 ; n5980
g3545 nor pi0215 n5980 ; n5981
g3546 and n3328_not n5981 ; n5982
g3547 and n3331_not n5981 ; n5983
g3548 nor n5778 n5897 ; n5984
g3549 nor pi0215 n5984 ; n5985
g3550 and n3331 n5985 ; n5986
g3551 and pi0062 n5983_not ; n5987
g3552 and n5986_not n5987 ; n5988
g3553 nor n2537 n5981 ; n5989
g3554 and n2537 n5985_not ; n5990
g3555 and pi0056 n5989_not ; n5991
g3556 and n5990_not n5991 ; n5992
g3557 and n2572_not n5981 ; n5993
g3558 and n2572 n5985 ; n5994
g3559 and pi0055 n5993_not ; n5995
g3560 and n5994_not n5995 ; n5996
g3561 and n2593 n5815 ; n5997
g3562 nor pi0299 n5997 ; n5998
g3563 and pi0223_not n5809 ; n5999
g3564 and n5998 n5999_not ; n6000
g3565 and pi0299 n5981_not ; n6001
g3566 nor n6000 n6001 ; n6002
g3567 and n2532_not n6002 ; n6003
g3568 and n2625_not n6002 ; n6004
g3569 and pi0299 n5985_not ; n6005
g3570 nor n6000 n6005 ; n6006
g3571 and n2625 n6006 ; n6007
g3572 nor n6004 n6007 ; n6008
g3573 and n2533 n6008_not ; n6009
g3574 and n2533_not n6002 ; n6010
g3575 and pi0092 n6010_not ; n6011
g3576 and n6009_not n6011 ; n6012
g3577 and pi0075 n6002 ; n6013
g3578 and pi0087 n6008 ; n6014
g3579 and pi0038 n6002 ; n6015
g3580 and pi0039 n6006_not ; n6016
g3581 and n3470 n5927 ; n6017
g3582 and n5853 n5942_not ; n6018
g3583 and n3470 n5835_not ; n6019
g3584 nor pi0039 n6019 ; n6020
g3585 and n6017_not n6020 ; n6021
g3586 and n6018_not n6021 ; n6022
g3587 nor pi0038 n6016 ; n6023
g3588 and n6022_not n6023 ; n6024
g3589 nor pi0100 n6015 ; n6025
g3590 and n6024_not n6025 ; n6026
g3591 and n2530_not n6002 ; n6027
g3592 nor n5778 n5953 ; n6028
g3593 nor pi0215 n6028 ; n6029
g3594 and pi0299 n6029_not ; n6030
g3595 and n2530 n6000_not ; n6031
g3596 and n6030_not n6031 ; n6032
g3597 and pi0100 n6027_not ; n6033
g3598 and n6032_not n6033 ; n6034
g3599 nor n6026 n6034 ; n6035
g3600 nor pi0087 n6035 ; n6036
g3601 nor pi0075 n6014 ; n6037
g3602 and n6036_not n6037 ; n6038
g3603 nor pi0092 n6013 ; n6039
g3604 and n6038_not n6039 ; n6040
g3605 and n2532 n6012_not ; n6041
g3606 and n6040_not n6041 ; n6042
g3607 nor pi0055 n6003 ; n6043
g3608 and n6042_not n6043 ; n6044
g3609 nor pi0056 n5996 ; n6045
g3610 and n6044_not n6045 ; n6046
g3611 nor pi0062 n5992 ; n6047
g3612 and n6046_not n6047 ; n6048
g3613 and n3328 n5988_not ; n6049
g3614 and n6048_not n6049 ; n6050
g3615 nor pi0242 n5982 ; n6051
g3616 and n6050_not n6051 ; n6052
g3617 and n3450_not n5981 ; n6053
g3618 and n3328_not n6053 ; n6054
g3619 nor n5778 n5793 ; n6055
g3620 nor pi0215 n6055 ; n6056
g3621 and n3331 n6056 ; n6057
g3622 and n3331_not n6053 ; n6058
g3623 and pi0062 n6058_not ; n6059
g3624 and n6057_not n6059 ; n6060
g3625 nor n2537 n6053 ; n6061
g3626 and n2537 n6056_not ; n6062
g3627 and pi0056 n6061_not ; n6063
g3628 and n6062_not n6063 ; n6064
g3629 and n2572 n6056 ; n6065
g3630 and n2572_not n6053 ; n6066
g3631 and pi0055 n6066_not ; n6067
g3632 and n6065_not n6067 ; n6068
g3633 and pi0299 n6053_not ; n6069
g3634 nor n5998 n6069 ; n6070
g3635 and n2532_not n6070 ; n6071
g3636 and n2625_not n6070 ; n6072
g3637 and pi0299 n6056_not ; n6073
g3638 nor n5998 n6073 ; n6074
g3639 and n2625 n6074 ; n6075
g3640 nor n6072 n6075 ; n6076
g3641 and n2533 n6076_not ; n6077
g3642 and n2533_not n6070 ; n6078
g3643 and pi0092 n6078_not ; n6079
g3644 and n6077_not n6079 ; n6080
g3645 and pi0075 n6070 ; n6081
g3646 and pi0087 n6076 ; n6082
g3647 and pi0038 n6070 ; n6083
g3648 and pi0039 n6074_not ; n6084
g3649 and n5852_not n5853 ; n6085
g3650 and n6020 n6085_not ; n6086
g3651 nor pi0038 n6084 ; n6087
g3652 and n6086_not n6087 ; n6088
g3653 nor pi0100 n6083 ; n6089
g3654 and n6088_not n6089 ; n6090
g3655 and n2530_not n6070 ; n6091
g3656 nor n5778 n5868 ; n6092
g3657 nor pi0215 n6092 ; n6093
g3658 and pi0299 n6093_not ; n6094
g3659 and n2530 n5998_not ; n6095
g3660 and n6094_not n6095 ; n6096
g3661 and pi0100 n6091_not ; n6097
g3662 and n6096_not n6097 ; n6098
g3663 nor n6090 n6098 ; n6099
g3664 nor pi0087 n6099 ; n6100
g3665 nor pi0075 n6082 ; n6101
g3666 and n6100_not n6101 ; n6102
g3667 nor pi0092 n6081 ; n6103
g3668 and n6102_not n6103 ; n6104
g3669 and n2532 n6080_not ; n6105
g3670 and n6104_not n6105 ; n6106
g3671 nor pi0055 n6071 ; n6107
g3672 and n6106_not n6107 ; n6108
g3673 nor pi0056 n6068 ; n6109
g3674 and n6108_not n6109 ; n6110
g3675 nor pi0062 n6064 ; n6111
g3676 and n6110_not n6111 ; n6112
g3677 and n3328 n6060_not ; n6113
g3678 and n6112_not n6113 ; n6114
g3679 and pi0242 n6054_not ; n6115
g3680 and n6114_not n6115 ; n6116
g3681 and pi1134 n6052_not ; n6117
g3682 and n6116_not n6117 ; n6118
g3683 nor n5979 n6118 ; po0165
g3684 and pi0057 pi0059 ; n6120
g3685 and n2521 n2538 ; n6121
g3686 nor n3328 n6121 ; n6122
g3687 nor n6120 n6122 ; n6123
g3688 and pi0057 n6123_not ; n6124
g3689 and n2512 n2625 ; n6125
g3690 and n2536 n6125 ; n6126
g3691 and pi0056 n6126_not ; n6127
g3692 and pi0054_not n2534 ; n6128
g3693 and n6125 n6128 ; n6129
g3694 and pi0074 n6129_not ; n6130
g3695 nor pi0055 n6130 ; n6131
g3696 and pi0087 n6125_not ; n6132
g3697 nor pi0075 n6132 ; n6133
g3698 nor pi0054 pi0092 ; n6134
g3699 and pi0039_not n2512 ; n6135
g3700 and pi0038 n6135_not ; n6136
g3701 nor pi0100 n6136 ; n6137
g3702 and pi0058 n2502 ; n6138
g3703 nor pi0090 n6138 ; n6139
g3704 and n2720 n2769 ; n6140
g3705 and n2874 n6140 ; n6141
g3706 and n2781 n6141_not ; n6142
g3707 nor n2776 n6142 ; n6143
g3708 nor pi0108 n6143 ; n6144
g3709 and n2775 n6144_not ; n6145
g3710 and pi0110_not n2889 ; n6146
g3711 and n6145_not n6146 ; n6147
g3712 nor n2759 n2766 ; n6148
g3713 and n6147_not n6148 ; n6149
g3714 nor pi0047 n6149 ; n6150
g3715 and n2700 n2762_not ; n6151
g3716 and n6150_not n6151 ; n6152
g3717 and n6139 n6152_not ; n6153
g3718 nor n2896 n6153 ; n6154
g3719 nor pi0093 n6154 ; n6155
g3720 and pi0841_not n2503 ; n6156
g3721 and pi0093 n6156_not ; n6157
g3722 nor n6155 n6157 ; n6158
g3723 nor pi0035 n6158 ; n6159
g3724 nor pi0070 n2729 ; n6160
g3725 and n6159_not n6160 ; n6161
g3726 nor pi0051 n6161 ; n6162
g3727 and n2748 n6162_not ; n6163
g3728 and n3168 n6163_not ; n6164
g3729 and n2746 n6164_not ; n6165
g3730 and n2744 n6165_not ; n6166
g3731 nor pi0198 pi0299 ; n6167
g3732 and pi0210_not pi0299 ; n6168
g3733 nor n6167 n6168 ; n6169
g3734 and pi0035_not n2508 ; n6170
g3735 and pi0040_not n6170 ; n6171
g3736 and n2915 n6171 ; n6172
g3737 and pi0032 n6172_not ; n6173
g3738 nor n6169 n6173 ; n6174
g3739 and n3412_not n6169 ; n6175
g3740 nor n6174 n6175 ; n6176
g3741 nor n6166 n6176 ; n6177
g3742 nor pi0095 n6177 ; n6178
g3743 nor n2741 n6178 ; n6179
g3744 nor pi0039 n6179 ; n6180
g3745 and pi0835 pi0984 ; n6181
g3746 nor pi0252 pi1001 ; n6182
g3747 nor pi0979 n6182 ; n6183
g3748 and n6181_not n6183 ; n6184
g3749 and pi0287_not n6184 ; n6185
g3750 and pi0835 pi0950 ; n6186
g3751 and n6185 n6186 ; n6187
g3752 and n2928 n6187 ; n6188
g3753 and pi0222 pi0224 ; n6189
g3754 and pi0603 pi0642_not ; n6190
g3755 nor pi0614 pi0616 ; n6191
g3756 and n6190 n6191 ; n6192
g3757 and pi0662_not pi0680 ; n6193
g3758 and pi0661_not n6193 ; n6194
g3759 and pi0681_not n6194 ; n6195
g3760 or n6192 n6195 ; po1101
g3761 nor pi0332 pi0468 ; n6197
g3762 and po1101 n6197_not ; n6198
g3763 nor pi0587 pi0602 ; n6199
g3764 nor pi0961 pi0967 ; n6200
g3765 nor pi0969 pi0971 ; n6201
g3766 nor pi0974 pi0977 ; n6202
g3767 and n6201 n6202 ; n6203
g3768 and n6199 n6200 ; n6204
g3769 and n6203 n6204 ; n6205
g3770 and n6197 n6205_not ; n6206
g3771 nor n6198 n6206 ; n6207
g3772 and n6188 n6189 ; n6208
g3773 and n6207_not n6208 ; n6209
g3774 and n2521 n6209_not ; n6210
g3775 nor pi0223 n6210 ; n6211
g3776 and pi1092 n6187 ; n6212
g3777 nor pi0824 pi0829 ; n6213
g3778 and pi0824 pi1091_not ; n6214
g3779 and pi1093 n2924_not ; n6215
g3780 and n6214_not n6215 ; n6216
g3781 nor n6213 n6216 ; n6217
g3782 and n6212 n6217 ; n6218
g3783 nor n6197 n6218 ; n6219
g3784 and po1101 n6219_not ; n6220
g3785 and n2521 n6220_not ; n6221
g3786 and n2512 n6197 ; n6222
g3787 and po1101 n6222 ; n6223
g3788 nor n6221 n6223 ; n6224
g3789 and n6205 n6224_not ; n6225
g3790 nor n6192 n6197 ; n6226
g3791 and n6195_not n6226 ; n6227
g3792 and n6218 n6227_not ; n6228
g3793 and n2521 n6228_not ; n6229
g3794 and n6205_not n6229 ; n6230
g3795 and pi0223 n6230_not ; n6231
g3796 and n6225_not n6231 ; n6232
g3797 nor pi0299 n6211 ; n6233
g3798 and n6232_not n6233 ; n6234
g3799 and pi0216 pi0221 ; n6235
g3800 nor pi0907 pi0947 ; n6236
g3801 nor pi0960 pi0963 ; n6237
g3802 nor pi0970 pi0972 ; n6238
g3803 nor pi0975 pi0978 ; n6239
g3804 and n6238 n6239 ; n6240
g3805 and n6237 n6240 ; n6241
g3806 and n6236 n6241 ; n6242
g3807 and n6197 n6242_not ; n6243
g3808 nor n6198 n6243 ; n6244
g3809 and n6188 n6235 ; n6245
g3810 and n6244_not n6245 ; n6246
g3811 and n2521 n6246_not ; n6247
g3812 nor pi0215 n6247 ; n6248
g3813 and n6229 n6242_not ; n6249
g3814 and n6224_not n6242 ; n6250
g3815 and pi0215 n6249_not ; n6251
g3816 and n6250_not n6251 ; n6252
g3817 and pi0299 n6248_not ; n6253
g3818 and n6252_not n6253 ; n6254
g3819 and pi0039 n6234_not ; n6255
g3820 and n6254_not n6255 ; n6256
g3821 nor n6180 n6256 ; n6257
g3822 nor pi0038 n6257 ; n6258
g3823 and n6137 n6258_not ; n6259
g3824 nor pi0142 n2669 ; n6260
g3825 and pi0299_not n6260 ; n6261
g3826 and pi0299 n2640 ; n6262
g3827 nor n6261 n6262 ; n6263
g3828 and n3385_not n6263 ; n6264
g3829 nor pi0041 pi0099 ; n6265
g3830 and pi0101_not n6265 ; n6266
g3831 nor pi0042 pi0043 ; n6267
g3832 and pi0052_not n6267 ; n6268
g3833 nor pi0113 pi0116 ; n6269
g3834 nor pi0114 pi0115 ; n6270
g3835 and n6269 n6270 ; n6271
g3836 and n6268 n6271 ; n6272
g3837 and n6266 n6272 ; n6273
g3838 nand pi0044_not n6273 ; po1057
g3839 and pi0683_not po1057 ; n6275
g3840 and pi0129 pi0250 ; n6276
g3841 and n2932 n6213_not ; n6277
g3842 and pi1093_not n6277 ; po0740
g3843 nor pi0250 po0740 ; n6279
g3844 nor n6276 n6279 ; n6280
g3845 nor n6275 n6280 ; n6281
g3846 and n6263_not po1057 ; n6282
g3847 and n6281 n6282 ; n6283
g3848 and pi0039_not n2521 ; n6284
g3849 and pi0038_not pi0100 ; n6285
g3850 and n6284 n6285 ; n6286
g3851 nor n6264 n6283 ; n6287
g3852 and n6286 n6287 ; n6288
g3853 nor pi0087 n6288 ; n6289
g3854 and n6259_not n6289 ; n6290
g3855 and n6133 n6134 ; n6291
g3856 and n6290_not n6291 ; n6292
g3857 nor pi0074 n6292 ; n6293
g3858 and n6131 n6293_not ; n6294
g3859 nor pi0056 n6294 ; n6295
g3860 nor n6127 n6295 ; n6296
g3861 nor pi0062 n6296 ; n6297
g3862 and n3330 n6125 ; n6298
g3863 and pi0062 n6298_not ; n6299
g3864 nor pi0059 n6299 ; n6300
g3865 and n6297_not n6300 ; n6301
g3866 nor pi0057 n6301 ; n6302
g3867 nor n6124 n6302 ; po0167
g3868 and pi0055_not n2529 ; n6304
g3869 and pi0059_not n6304 ; n6305
g3870 nor pi0228 n6305 ; n6306
g3871 and pi0057 n6306_not ; n6307
g3872 nor n6195 n6197 ; n6308
g3873 and pi0907_not n6197 ; n6309
g3874 nor n6308 n6309 ; n6310
g3875 nor pi0228 n2572 ; n6311
g3876 and pi0030 pi0228 ; n6312
g3877 nor n3335 n6312 ; n6313
g3878 nor n6311 n6313 ; n6314
g3879 and n6310 n6314 ; n6315
g3880 and n6307 n6315 ; n6316
g3881 nor pi0228 n6304 ; n6317
g3882 and n6315 n6317_not ; n6318
g3883 and pi0059 n6318_not ; n6319
g3884 and n6310 n6312 ; n6320
g3885 and n2529_not n6320 ; n6321
g3886 and pi0055 n6315_not ; n6322
g3887 and pi0054_not n2569 ; n6323
g3888 and pi0299 n6310 ; n6324
g3889 and pi0602_not n6197 ; n6325
g3890 nor n6308 n6325 ; n6326
g3891 and pi0299_not n6326 ; n6327
g3892 nor n6324 n6327 ; n6328
g3893 and n6312 n6328_not ; n6329
g3894 nor n6323 n6329 ; n6330
g3895 and n2610_not n6329 ; n6331
g3896 nor pi0039 n6313 ; n6332
g3897 and n6328_not n6332 ; n6333
g3898 and n2620 n6333 ; n6334
g3899 nor n6331 n6334 ; n6335
g3900 and n2569 n6335 ; n6336
g3901 and pi0054_not n6336 ; n6337
g3902 and pi0074 n6330_not ; n6338
g3903 and n6337_not n6338 ; n6339
g3904 nor n2569 n6329 ; n6340
g3905 nor n6336 n6340 ; n6341
g3906 and pi0054 n6341_not ; n6342
g3907 and pi0075_not n6335 ; n6343
g3908 and pi0075 n6329_not ; n6344
g3909 and pi0092 n6344_not ; n6345
g3910 and n6343_not n6345 ; n6346
g3911 and pi0075 n6335 ; n6347
g3912 and pi0087 n6329 ; n6348
g3913 and n2530_not n6329 ; n6349
g3914 and n6312 n6326 ; n6350
g3915 and n2521 n6280_not ; n6351
g3916 and pi0683 po1057 ; n6352
g3917 and n6351 n6352 ; n6353
g3918 and n6308_not n6353 ; n6354
g3919 and n6260 n6354 ; n6355
g3920 and pi0252 n6260_not ; n6356
g3921 and pi0252 n6222 ; n6357
g3922 and n6195_not n6357 ; n6358
g3923 and pi0252 n2521 ; n6359
g3924 and n6195 n6359 ; n6360
g3925 nor n6358 n6360 ; n6361
g3926 and n6356 n6361_not ; n6362
g3927 nor n6355 n6362 ; n6363
g3928 nor pi0228 n6325 ; n6364
g3929 and n6363_not n6364 ; n6365
g3930 nor pi0299 n6350 ; n6366
g3931 and n6365_not n6366 ; n6367
g3932 and pi0299 n6320_not ; n6368
g3933 and n2640 n6354_not ; n6369
g3934 and n2640_not n6361 ; n6370
g3935 nor pi0228 n6309 ; n6371
g3936 and n6369_not n6371 ; n6372
g3937 and n6370_not n6372 ; n6373
g3938 and n6368 n6373_not ; n6374
g3939 and n2530 n6374_not ; n6375
g3940 and n6367_not n6375 ; n6376
g3941 and pi0100 n6349_not ; n6377
g3942 and n6376_not n6377 ; n6378
g3943 and pi0215_not pi0221 ; n6379
g3944 and pi0287_not n2521 ; n6380
g3945 and pi0835 n6184 ; n6381
g3946 and n6380 n6381 ; n6382
g3947 and pi0824 pi1093 ; n6383
g3948 and n2932 n6383 ; n6384
g3949 and n6382 n6384 ; n6385
g3950 and pi1091_not n6385 ; n6386
g3951 and pi1091 n2923 ; n6387
g3952 and n6384 n6387_not ; n6388
g3953 nor n2928 n6388 ; n6389
g3954 and pi1091 n6389_not ; n6390
g3955 and n6382 n6390 ; n6391
g3956 nor n6386 n6391 ; n6392
g3957 and pi0216 n6392_not ; n6393
g3958 nor pi0829 n2923 ; n6394
g3959 and pi1091 n6394_not ; n6395
g3960 and n6385 n6395_not ; n6396
g3961 and pi0216_not n6396 ; n6397
g3962 nor n6393 n6397 ; n6398
g3963 nor pi0228 n6398 ; n6399
g3964 nor n6312 n6399 ; n6400
g3965 and n6379 n6400_not ; n6401
g3966 nor n6312 n6401 ; n6402
g3967 and n6310 n6402_not ; n6403
g3968 and pi0299 n6403_not ; n6404
g3969 and pi0222 pi0223_not ; n6405
g3970 nor pi0224 n6396 ; n6406
g3971 and pi0224 n6392 ; n6407
g3972 and n6405 n6406_not ; n6408
g3973 and n6407_not n6408 ; n6409
g3974 and pi0228_not n6409 ; n6410
g3975 nor n6312 n6410 ; n6411
g3976 and n6326 n6411_not ; n6412
g3977 nor pi0299 n6412 ; n6413
g3978 and pi0039 n6413_not ; n6414
g3979 and n6404_not n6414 ; n6415
g3980 and pi0158 pi0159 ; n6416
g3981 and pi0160 pi0197 ; n6417
g3982 and n6416 n6417 ; n6418
g3983 and pi0091 n2755_not ; n6419
g3984 nor pi0058 n6419 ; n6420
g3985 nor pi0091 pi0314 ; n6421
g3986 and n2765 n2766_not ; n6422
g3987 and pi0067 n2483 ; n6423
g3988 and pi0085 n2827 ; n6424
g3989 and n2469 n6424_not ; n6425
g3990 and n2831 n6425_not ; n6426
g3991 and n2478 n6426_not ; n6427
g3992 nor n2810 n2811 ; n6428
g3993 and n6427_not n6428 ; n6429
g3994 and n2479 n6429 ; n6430
g3995 nor n2807 n6430 ; n6431
g3996 and n2804 n6431_not ; n6432
g3997 and n2797 n6423_not ; n6433
g3998 and n6432_not n6433 ; n6434
g3999 and n2796 n6434_not ; n6435
g4000 nor pi0071 n6435 ; n6436
g4001 nand pi0064_not n2487 ; po1049
g4002 and n2791 po1049_not ; n6438
g4003 and n6436_not n6438 ; n6439
g4004 nor pi0081 n6439 ; n6440
g4005 and n2845 n6438 ; n6441
g4006 and n6440 n6441_not ; n6442
g4007 nor pi0102 n2786 ; n6443
g4008 and n2463 n6443 ; n6444
g4009 and n6442_not n6444 ; n6445
g4010 and n2785 n6445_not ; n6446
g4011 and n2877 n6446_not ; n6447
g4012 and n2719 n6447_not ; n6448
g4013 nor n2722 n6448 ; n6449
g4014 nor pi0086 n6449 ; n6450
g4015 and pi0046_not n2496 ; n6451
g4016 and n2783 n6451 ; n6452
g4017 and n6450_not n6452 ; n6453
g4018 and n2889 n6453_not ; n6454
g4019 and n6422 n6454_not ; n6455
g4020 and n6421 n6455_not ; n6456
g4021 and pi0091_not pi0314 ; n6457
g4022 and n6440_not n6444 ; n6458
g4023 and n2785 n6458_not ; n6459
g4024 and n2877 n6459_not ; n6460
g4025 and n2719 n6460_not ; n6461
g4026 nor n2722 n6461 ; n6462
g4027 nor pi0086 n6462 ; n6463
g4028 and n6452 n6463_not ; n6464
g4029 and n2889 n6464_not ; n6465
g4030 and n6422 n6465_not ; n6466
g4031 and n6457 n6466_not ; n6467
g4032 and n6420 n6467_not ; n6468
g4033 and n6456_not n6468 ; n6469
g4034 nor pi0090 n6469 ; n6470
g4035 nor n2896 n6470 ; n6471
g4036 nor pi0093 n6471 ; n6472
g4037 and pi0093 n2914_not ; n6473
g4038 nor pi0035 n6473 ; n6474
g4039 and n6472_not n6474 ; n6475
g4040 nor pi0070 n6475 ; n6476
g4041 and n3100 n6476_not ; n6477
g4042 nor pi0072 n6477 ; n6478
g4043 and pi0095_not n2510 ; n6479
g4044 and n2745_not n6479 ; n6480
g4045 and n6478_not n6480 ; n6481
g4046 nor n3181 n6481 ; n6482
g4047 and pi0841_not n2728 ; n6483
g4048 and n2962 n6483 ; n6484
g4049 and n2736 n6484 ; n6485
g4050 and pi0032 n6485 ; n6486
g4051 and pi0095_not n6486 ; n6487
g4052 and pi0210_not n6487 ; n6488
g4053 and n6482 n6488_not ; n6489
g4054 nor n6197 n6489 ; n6490
g4055 and pi0047_not n2493 ; n6491
g4056 nor n2888 n6453 ; n6492
g4057 and n6491 n6492_not ; n6493
g4058 and n6421 n6493_not ; n6494
g4059 nor n2888 n6464 ; n6495
g4060 and n6491 n6495_not ; n6496
g4061 and n6457 n6496_not ; n6497
g4062 and n6420 n6497_not ; n6498
g4063 and n6494_not n6498 ; n6499
g4064 nor pi0090 n6499 ; n6500
g4065 nor n2896 n6500 ; n6501
g4066 nor pi0093 n6501 ; n6502
g4067 and n6474 n6502_not ; n6503
g4068 nor pi0070 n6503 ; n6504
g4069 and n3100 n6504_not ; n6505
g4070 nor pi0072 n6505 ; n6506
g4071 and n6480 n6506_not ; n6507
g4072 nor n3181 n6507 ; n6508
g4073 and n6488_not n6508 ; n6509
g4074 and n6197 n6509_not ; n6510
g4075 nor n6490 n6510 ; n6511
g4076 and n6310 n6511_not ; n6512
g4077 and n6418 n6512_not ; n6513
g4078 and n6310 n6489_not ; n6514
g4079 nor n6418 n6514 ; n6515
g4080 nor pi0228 n6515 ; n6516
g4081 and n6513_not n6516 ; n6517
g4082 and n6368 n6517_not ; n6518
g4083 and pi0198_not n6487 ; n6519
g4084 and n6482 n6519_not ; n6520
g4085 nor pi0228 n6520 ; n6521
g4086 nor n6312 n6521 ; n6522
g4087 and n6326 n6522_not ; n6523
g4088 nor pi0299 n6523 ; n6524
g4089 and pi0145 pi0180 ; n6525
g4090 and pi0181 pi0182 ; n6526
g4091 and n6525 n6526 ; n6527
g4092 and pi0299_not n6527 ; n6528
g4093 nor n6524 n6528 ; n6529
g4094 nor n6197 n6520 ; n6530
g4095 and n6508 n6519_not ; n6531
g4096 and n6197 n6531_not ; n6532
g4097 nor n6530 n6532 ; n6533
g4098 and pi0228_not n6326 ; n6534
g4099 and n6533_not n6534 ; n6535
g4100 nor n6350 n6535 ; n6536
g4101 and n6527 n6536_not ; n6537
g4102 nor n6529 n6537 ; n6538
g4103 and pi0232 n6518_not ; n6539
g4104 and n6538_not n6539 ; n6540
g4105 and pi0228_not n6514 ; n6541
g4106 and n6368 n6541_not ; n6542
g4107 nor pi0232 n6542 ; n6543
g4108 and n6524_not n6543 ; n6544
g4109 nor n6540 n6544 ; n6545
g4110 nor pi0039 n6545 ; n6546
g4111 nor pi0038 n6415 ; n6547
g4112 and n6546_not n6547 ; n6548
g4113 and pi0038 n6329_not ; n6549
g4114 and n6333_not n6549 ; n6550
g4115 nor n6548 n6550 ; n6551
g4116 nor pi0100 n6551 ; n6552
g4117 nor pi0087 n6378 ; n6553
g4118 and n6552_not n6553 ; n6554
g4119 nor pi0075 n6348 ; n6555
g4120 and n6554_not n6555 ; n6556
g4121 nor pi0092 n6347 ; n6557
g4122 and n6556_not n6557 ; n6558
g4123 nor pi0054 n6346 ; n6559
g4124 and n6558_not n6559 ; n6560
g4125 nor pi0074 n6342 ; n6561
g4126 and n6560_not n6561 ; n6562
g4127 nor pi0055 n6339 ; n6563
g4128 and n6562_not n6563 ; n6564
g4129 and n2529 n6322_not ; n6565
g4130 and n6564_not n6565 ; n6566
g4131 nor pi0059 n6321 ; n6567
g4132 and n6566_not n6567 ; n6568
g4133 nor pi0057 n6319 ; n6569
g4134 and n6568_not n6569 ; n6570
g4135 nor n6316 n6570 ; po0171
g4136 and pi0947_not n6197 ; n6572
g4137 nor n6226 n6572 ; n6573
g4138 and n6314 n6573 ; n6574
g4139 and n6307 n6574 ; n6575
g4140 and n6317_not n6574 ; n6576
g4141 and pi0059 n6576_not ; n6577
g4142 and n6312 n6573 ; n6578
g4143 and n2529_not n6578 ; n6579
g4144 and pi0055 n6574_not ; n6580
g4145 and pi0299 n6573_not ; n6581
g4146 and pi0587_not n6197 ; n6582
g4147 nor n6226 n6582 ; n6583
g4148 nor pi0299 n6583 ; n6584
g4149 nor n6581 n6584 ; n6585
g4150 and n6312 n6585 ; n6586
g4151 nor n6323 n6586 ; n6587
g4152 and n2610_not n6586 ; n6588
g4153 and n6332 n6585 ; n6589
g4154 and n2620 n6589 ; n6590
g4155 nor n6588 n6590 ; n6591
g4156 and n2569 n6591 ; n6592
g4157 and pi0054_not n6592 ; n6593
g4158 and pi0074 n6587_not ; n6594
g4159 and n6593_not n6594 ; n6595
g4160 nor n2569 n6586 ; n6596
g4161 nor n6592 n6596 ; n6597
g4162 and pi0054 n6597_not ; n6598
g4163 and pi0075_not n6591 ; n6599
g4164 and pi0075 n6586_not ; n6600
g4165 and pi0092 n6600_not ; n6601
g4166 and n6599_not n6601 ; n6602
g4167 and pi0075 n6591 ; n6603
g4168 and pi0087 n6586 ; n6604
g4169 and n2530_not n6586 ; n6605
g4170 and pi0299 n6578_not ; n6606
g4171 and n6226_not n6353 ; n6607
g4172 and n2640 n6572_not ; n6608
g4173 and n6607 n6608 ; n6609
g4174 nor n6192 n6357 ; n6610
g4175 and n6192 n6359_not ; n6611
g4176 nor n6610 n6611 ; n6612
g4177 and n6192 n6197_not ; n6613
g4178 nor pi0947 n6613 ; n6614
g4179 nor n2640 n6614 ; n6615
g4180 and n6612 n6615 ; n6616
g4181 nor n6609 n6616 ; n6617
g4182 nor pi0228 n6617 ; n6618
g4183 and n6606 n6618_not ; n6619
g4184 and pi0228_not n2669 ; n6620
g4185 and n6582_not n6612 ; n6621
g4186 and n6620 n6621_not ; n6622
g4187 nor pi0587 n6613 ; n6623
g4188 and pi0142 n6612_not ; n6624
g4189 nor pi0142 n6607 ; n6625
g4190 nor pi0228 n6623 ; n6626
g4191 and n6625_not n6626 ; n6627
g4192 and n6624_not n6627 ; n6628
g4193 and n6312 n6583 ; n6629
g4194 nor n6620 n6629 ; n6630
g4195 and n6628_not n6630 ; n6631
g4196 nor n6622 n6631 ; n6632
g4197 nor pi0299 n6632 ; n6633
g4198 and n2530 n6619_not ; n6634
g4199 and n6633_not n6634 ; n6635
g4200 and pi0100 n6605_not ; n6636
g4201 and n6635_not n6636 ; n6637
g4202 and n6411_not n6583 ; n6638
g4203 nor pi0299 n6638 ; n6639
g4204 and pi0299 n6379 ; n6640
g4205 nor n6606 n6640 ; n6641
g4206 and n6401 n6573 ; n6642
g4207 nor n6641 n6642 ; n6643
g4208 and pi0039 n6639_not ; n6644
g4209 and n6643_not n6644 ; n6645
g4210 and n6511_not n6573 ; n6646
g4211 and n6418 n6646_not ; n6647
g4212 and n6489_not n6573 ; n6648
g4213 nor n6418 n6648 ; n6649
g4214 nor pi0228 n6649 ; n6650
g4215 and n6647_not n6650 ; n6651
g4216 and n6606 n6651_not ; n6652
g4217 and n6522_not n6583 ; n6653
g4218 and n6527_not n6653 ; n6654
g4219 and pi0228_not n6583 ; n6655
g4220 and n6533_not n6655 ; n6656
g4221 nor n6629 n6656 ; n6657
g4222 and n6527 n6657_not ; n6658
g4223 nor pi0299 n6654 ; n6659
g4224 and n6658_not n6659 ; n6660
g4225 and pi0232 n6652_not ; n6661
g4226 and n6660_not n6661 ; n6662
g4227 and pi0228_not n6648 ; n6663
g4228 and n6606 n6663_not ; n6664
g4229 nor pi0299 n6653 ; n6665
g4230 nor pi0232 n6664 ; n6666
g4231 and n6665_not n6666 ; n6667
g4232 nor n6662 n6667 ; n6668
g4233 nor pi0039 n6668 ; n6669
g4234 nor pi0038 n6645 ; n6670
g4235 and n6669_not n6670 ; n6671
g4236 and pi0038 n6586_not ; n6672
g4237 and n6589_not n6672 ; n6673
g4238 nor n6671 n6673 ; n6674
g4239 nor pi0100 n6674 ; n6675
g4240 nor pi0087 n6637 ; n6676
g4241 and n6675_not n6676 ; n6677
g4242 nor pi0075 n6604 ; n6678
g4243 and n6677_not n6678 ; n6679
g4244 nor pi0092 n6603 ; n6680
g4245 and n6679_not n6680 ; n6681
g4246 nor pi0054 n6602 ; n6682
g4247 and n6681_not n6682 ; n6683
g4248 nor pi0074 n6598 ; n6684
g4249 and n6683_not n6684 ; n6685
g4250 nor pi0055 n6595 ; n6686
g4251 and n6685_not n6686 ; n6687
g4252 and n2529 n6580_not ; n6688
g4253 and n6687_not n6688 ; n6689
g4254 nor pi0059 n6579 ; n6690
g4255 and n6689_not n6690 ; n6691
g4256 nor pi0057 n6577 ; n6692
g4257 and n6691_not n6692 ; n6693
g4258 nor n6575 n6693 ; po0172
g4259 and pi0030 n6197 ; n6695
g4260 and pi0228 n6695 ; n6696
g4261 and pi0970 n6696 ; n6697
g4262 and pi0228_not pi0970 ; n6698
g4263 and n6222 n6698 ; n6699
g4264 and n2572 n6699 ; n6700
g4265 and n6305 n6700 ; n6701
g4266 nor n6697 n6701 ; n6702
g4267 and pi0057 n6702_not ; n6703
g4268 and n6304 n6700 ; n6704
g4269 and pi0059 n6697_not ; n6705
g4270 and n6704_not n6705 ; n6706
g4271 and n2529_not n6697 ; n6707
g4272 and pi0055 n6697_not ; n6708
g4273 and n6700_not n6708 ; n6709
g4274 and pi0299 pi0970 ; n6710
g4275 and pi0299_not pi0967 ; n6711
g4276 nor n6710 n6711 ; n6712
g4277 and n6696 n6712_not ; n6713
g4278 nor n6323 n6713 ; n6714
g4279 and n2610_not n6713 ; n6715
g4280 and pi0299 n6697_not ; n6716
g4281 and n6699_not n6716 ; n6717
g4282 and pi0228 n6695_not ; n6718
g4283 nor pi0228 n6222 ; n6719
g4284 nor n6718 n6719 ; n6720
g4285 and pi0967 n6720 ; n6721
g4286 nor pi0299 n6721 ; n6722
g4287 nor pi0039 n6717 ; n6723
g4288 and n6722_not n6723 ; n6724
g4289 and n2620 n6724 ; n6725
g4290 nor n6715 n6725 ; n6726
g4291 and n2569 n6726 ; n6727
g4292 and pi0054_not n6727 ; n6728
g4293 and pi0074 n6714_not ; n6729
g4294 and n6728_not n6729 ; n6730
g4295 nor n2569 n6713 ; n6731
g4296 nor n6727 n6731 ; n6732
g4297 and pi0054 n6732_not ; n6733
g4298 and pi0075_not n6726 ; n6734
g4299 and pi0075 n6713_not ; n6735
g4300 and pi0092 n6735_not ; n6736
g4301 and n6734_not n6736 ; n6737
g4302 and pi0075 n6726 ; n6738
g4303 and pi0087 n6713 ; n6739
g4304 and n2530_not n6713 ; n6740
g4305 nor n2640 n6357 ; n6741
g4306 and n6197 n6353 ; n6742
g4307 and n2640 n6742_not ; n6743
g4308 nor pi0228 n6741 ; n6744
g4309 and n6743_not n6744 ; n6745
g4310 and pi0970 n6745 ; n6746
g4311 and n6716 n6746_not ; n6747
g4312 and n6260_not n6357 ; n6748
g4313 and n6260 n6742 ; n6749
g4314 nor pi0228 n6748 ; n6750
g4315 and n6749_not n6750 ; n6751
g4316 nor n6718 n6751 ; n6752
g4317 and pi0967 n6752 ; n6753
g4318 nor pi0299 n6753 ; n6754
g4319 and n2530 n6747_not ; n6755
g4320 and n6754_not n6755 ; n6756
g4321 and pi0100 n6740_not ; n6757
g4322 and n6756_not n6757 ; n6758
g4323 and n6379 n6398_not ; n6759
g4324 and n6197 n6759 ; n6760
g4325 nor pi0228 n6760 ; n6761
g4326 and n6710 n6761_not ; n6762
g4327 and n6197 n6409 ; n6763
g4328 nor pi0228 n6763 ; n6764
g4329 and n6711 n6764_not ; n6765
g4330 nor n6762 n6765 ; n6766
g4331 and pi0039 n6718_not ; n6767
g4332 and n6766_not n6767 ; n6768
g4333 and n6197 n6522_not ; n6769
g4334 nor n6527 n6769 ; n6770
g4335 nor n6520 n6527 ; n6771
g4336 and pi0228_not n6532 ; n6772
g4337 nor n6696 n6771 ; n6773
g4338 and n6772_not n6773 ; n6774
g4339 nor n6770 n6774 ; n6775
g4340 and pi0967 n6775 ; n6776
g4341 nor pi0299 n6776 ; n6777
g4342 and n6197 n6489_not ; n6778
g4343 and n6698 n6778 ; n6779
g4344 and n6716 n6779_not ; n6780
g4345 and pi0299 n6416 ; n6781
g4346 nor n6780 n6781 ; n6782
g4347 and n6417 n6510_not ; n6783
g4348 and n6417_not n6489 ; n6784
g4349 nor n6783 n6784 ; n6785
g4350 and n6197 n6785 ; n6786
g4351 and n6698 n6786 ; n6787
g4352 nor n6697 n6787 ; n6788
g4353 and n6416 n6788_not ; n6789
g4354 nor n6782 n6789 ; n6790
g4355 and pi0232 n6777_not ; n6791
g4356 and n6790_not n6791 ; n6792
g4357 and pi0967 n6769 ; n6793
g4358 nor pi0299 n6793 ; n6794
g4359 nor pi0232 n6780 ; n6795
g4360 and n6794_not n6795 ; n6796
g4361 nor n6792 n6796 ; n6797
g4362 nor pi0039 n6797 ; n6798
g4363 nor pi0038 n6768 ; n6799
g4364 and n6798_not n6799 ; n6800
g4365 and pi0039 n6713 ; n6801
g4366 and pi0038 n6801_not ; n6802
g4367 and n6724_not n6802 ; n6803
g4368 nor n6800 n6803 ; n6804
g4369 nor pi0100 n6804 ; n6805
g4370 nor pi0087 n6758 ; n6806
g4371 and n6805_not n6806 ; n6807
g4372 nor pi0075 n6739 ; n6808
g4373 and n6807_not n6808 ; n6809
g4374 nor pi0092 n6738 ; n6810
g4375 and n6809_not n6810 ; n6811
g4376 nor pi0054 n6737 ; n6812
g4377 and n6811_not n6812 ; n6813
g4378 nor pi0074 n6733 ; n6814
g4379 and n6813_not n6814 ; n6815
g4380 nor pi0055 n6730 ; n6816
g4381 and n6815_not n6816 ; n6817
g4382 and n2529 n6709_not ; n6818
g4383 and n6817_not n6818 ; n6819
g4384 nor pi0059 n6707 ; n6820
g4385 and n6819_not n6820 ; n6821
g4386 nor pi0057 n6706 ; n6822
g4387 and n6821_not n6822 ; n6823
g4388 nor n6703 n6823 ; po0173
g4389 and pi0972 n6696 ; n6825
g4390 and pi0228_not pi0972 ; n6826
g4391 and n6222 n6826 ; n6827
g4392 and n2572 n6827 ; n6828
g4393 and n6305 n6828 ; n6829
g4394 nor n6825 n6829 ; n6830
g4395 and pi0057 n6830_not ; n6831
g4396 and n6304 n6828 ; n6832
g4397 and pi0059 n6825_not ; n6833
g4398 and n6832_not n6833 ; n6834
g4399 and n2529_not n6825 ; n6835
g4400 and pi0055 n6825_not ; n6836
g4401 and n6828_not n6836 ; n6837
g4402 and pi0299_not pi0961 ; n6838
g4403 and pi0299 pi0972 ; n6839
g4404 nor n6838 n6839 ; n6840
g4405 and n6696 n6840_not ; n6841
g4406 nor n6323 n6841 ; n6842
g4407 and n2610_not n6841 ; n6843
g4408 and pi0299 n6825_not ; n6844
g4409 and n6827_not n6844 ; n6845
g4410 and pi0961 n6720 ; n6846
g4411 nor pi0299 n6846 ; n6847
g4412 nor pi0039 n6845 ; n6848
g4413 and n6847_not n6848 ; n6849
g4414 and n2620 n6849 ; n6850
g4415 nor n6843 n6850 ; n6851
g4416 and n2569 n6851 ; n6852
g4417 and pi0054_not n6852 ; n6853
g4418 and pi0074 n6842_not ; n6854
g4419 and n6853_not n6854 ; n6855
g4420 nor n2569 n6841 ; n6856
g4421 nor n6852 n6856 ; n6857
g4422 and pi0054 n6857_not ; n6858
g4423 and pi0075_not n6851 ; n6859
g4424 and pi0075 n6841_not ; n6860
g4425 and pi0092 n6860_not ; n6861
g4426 and n6859_not n6861 ; n6862
g4427 and pi0075 n6851 ; n6863
g4428 and pi0087 n6841 ; n6864
g4429 and n2530_not n6841 ; n6865
g4430 and pi0972 n6745 ; n6866
g4431 and n6844 n6866_not ; n6867
g4432 and pi0961 n6752 ; n6868
g4433 nor pi0299 n6868 ; n6869
g4434 and n2530 n6867_not ; n6870
g4435 and n6869_not n6870 ; n6871
g4436 and pi0100 n6865_not ; n6872
g4437 and n6871_not n6872 ; n6873
g4438 and n6764_not n6838 ; n6874
g4439 and n6761_not n6839 ; n6875
g4440 nor n6874 n6875 ; n6876
g4441 and n6767 n6876_not ; n6877
g4442 and pi0961 n6775 ; n6878
g4443 nor pi0299 n6878 ; n6879
g4444 and n6778 n6826 ; n6880
g4445 and n6844 n6880_not ; n6881
g4446 nor n6781 n6881 ; n6882
g4447 and n6786 n6826 ; n6883
g4448 nor n6825 n6883 ; n6884
g4449 and n6416 n6884_not ; n6885
g4450 nor n6882 n6885 ; n6886
g4451 and pi0232 n6879_not ; n6887
g4452 and n6886_not n6887 ; n6888
g4453 and pi0961 n6769 ; n6889
g4454 nor pi0299 n6889 ; n6890
g4455 nor pi0232 n6881 ; n6891
g4456 and n6890_not n6891 ; n6892
g4457 nor n6888 n6892 ; n6893
g4458 nor pi0039 n6893 ; n6894
g4459 nor pi0038 n6877 ; n6895
g4460 and n6894_not n6895 ; n6896
g4461 and pi0039 n6841 ; n6897
g4462 and pi0038 n6897_not ; n6898
g4463 and n6849_not n6898 ; n6899
g4464 nor n6896 n6899 ; n6900
g4465 nor pi0100 n6900 ; n6901
g4466 nor pi0087 n6873 ; n6902
g4467 and n6901_not n6902 ; n6903
g4468 nor pi0075 n6864 ; n6904
g4469 and n6903_not n6904 ; n6905
g4470 nor pi0092 n6863 ; n6906
g4471 and n6905_not n6906 ; n6907
g4472 nor pi0054 n6862 ; n6908
g4473 and n6907_not n6908 ; n6909
g4474 nor pi0074 n6858 ; n6910
g4475 and n6909_not n6910 ; n6911
g4476 nor pi0055 n6855 ; n6912
g4477 and n6911_not n6912 ; n6913
g4478 and n2529 n6837_not ; n6914
g4479 and n6913_not n6914 ; n6915
g4480 nor pi0059 n6835 ; n6916
g4481 and n6915_not n6916 ; n6917
g4482 nor pi0057 n6834 ; n6918
g4483 and n6917_not n6918 ; n6919
g4484 nor n6831 n6919 ; po0174
g4485 and pi0960 n6696 ; n6921
g4486 and pi0228_not pi0960 ; n6922
g4487 and n6222 n6922 ; n6923
g4488 and n2572 n6923 ; n6924
g4489 and n6305 n6924 ; n6925
g4490 nor n6921 n6925 ; n6926
g4491 and pi0057 n6926_not ; n6927
g4492 and n6304 n6924 ; n6928
g4493 and pi0059 n6921_not ; n6929
g4494 and n6928_not n6929 ; n6930
g4495 and n2529_not n6921 ; n6931
g4496 and pi0055 n6921_not ; n6932
g4497 and n6924_not n6932 ; n6933
g4498 and pi0299_not pi0977 ; n6934
g4499 and pi0299 pi0960 ; n6935
g4500 nor n6934 n6935 ; n6936
g4501 and n6696 n6936_not ; n6937
g4502 nor n6323 n6937 ; n6938
g4503 and n2610_not n6937 ; n6939
g4504 and pi0299 n6921_not ; n6940
g4505 and n6923_not n6940 ; n6941
g4506 and pi0977 n6720 ; n6942
g4507 nor pi0299 n6942 ; n6943
g4508 nor pi0039 n6941 ; n6944
g4509 and n6943_not n6944 ; n6945
g4510 and n2620 n6945 ; n6946
g4511 nor n6939 n6946 ; n6947
g4512 and n2569 n6947 ; n6948
g4513 and pi0054_not n6948 ; n6949
g4514 and pi0074 n6938_not ; n6950
g4515 and n6949_not n6950 ; n6951
g4516 nor n2569 n6937 ; n6952
g4517 nor n6948 n6952 ; n6953
g4518 and pi0054 n6953_not ; n6954
g4519 and pi0075_not n6947 ; n6955
g4520 and pi0075 n6937_not ; n6956
g4521 and pi0092 n6956_not ; n6957
g4522 and n6955_not n6957 ; n6958
g4523 and pi0075 n6947 ; n6959
g4524 and pi0087 n6937 ; n6960
g4525 and n2530_not n6937 ; n6961
g4526 and pi0960 n6745 ; n6962
g4527 and n6940 n6962_not ; n6963
g4528 and pi0977 n6752 ; n6964
g4529 nor pi0299 n6964 ; n6965
g4530 and n2530 n6963_not ; n6966
g4531 and n6965_not n6966 ; n6967
g4532 and pi0100 n6961_not ; n6968
g4533 and n6967_not n6968 ; n6969
g4534 and n6764_not n6934 ; n6970
g4535 and n6761_not n6935 ; n6971
g4536 nor n6970 n6971 ; n6972
g4537 and n6767 n6972_not ; n6973
g4538 and pi0977 n6775 ; n6974
g4539 nor pi0299 n6974 ; n6975
g4540 and n6778 n6922 ; n6976
g4541 and n6940 n6976_not ; n6977
g4542 nor n6781 n6977 ; n6978
g4543 and n6786 n6922 ; n6979
g4544 nor n6921 n6979 ; n6980
g4545 and n6416 n6980_not ; n6981
g4546 nor n6978 n6981 ; n6982
g4547 and pi0232 n6975_not ; n6983
g4548 and n6982_not n6983 ; n6984
g4549 and pi0977 n6769 ; n6985
g4550 nor pi0299 n6985 ; n6986
g4551 nor pi0232 n6977 ; n6987
g4552 and n6986_not n6987 ; n6988
g4553 nor n6984 n6988 ; n6989
g4554 nor pi0039 n6989 ; n6990
g4555 nor pi0038 n6973 ; n6991
g4556 and n6990_not n6991 ; n6992
g4557 and pi0039 n6937 ; n6993
g4558 and pi0038 n6993_not ; n6994
g4559 and n6945_not n6994 ; n6995
g4560 nor n6992 n6995 ; n6996
g4561 nor pi0100 n6996 ; n6997
g4562 nor pi0087 n6969 ; n6998
g4563 and n6997_not n6998 ; n6999
g4564 nor pi0075 n6960 ; n7000
g4565 and n6999_not n7000 ; n7001
g4566 nor pi0092 n6959 ; n7002
g4567 and n7001_not n7002 ; n7003
g4568 nor pi0054 n6958 ; n7004
g4569 and n7003_not n7004 ; n7005
g4570 nor pi0074 n6954 ; n7006
g4571 and n7005_not n7006 ; n7007
g4572 nor pi0055 n6951 ; n7008
g4573 and n7007_not n7008 ; n7009
g4574 and n2529 n6933_not ; n7010
g4575 and n7009_not n7010 ; n7011
g4576 nor pi0059 n6931 ; n7012
g4577 and n7011_not n7012 ; n7013
g4578 nor pi0057 n6930 ; n7014
g4579 and n7013_not n7014 ; n7015
g4580 nor n6927 n7015 ; po0175
g4581 and pi0963 n6696 ; n7017
g4582 and pi0228_not pi0963 ; n7018
g4583 and n6222 n7018 ; n7019
g4584 and n2572 n7019 ; n7020
g4585 and n6305 n7020 ; n7021
g4586 nor n7017 n7021 ; n7022
g4587 and pi0057 n7022_not ; n7023
g4588 and n6304 n7020 ; n7024
g4589 and pi0059 n7017_not ; n7025
g4590 and n7024_not n7025 ; n7026
g4591 and n2529_not n7017 ; n7027
g4592 and pi0055 n7017_not ; n7028
g4593 and n7020_not n7028 ; n7029
g4594 and pi0299_not pi0969 ; n7030
g4595 and pi0299 pi0963 ; n7031
g4596 nor n7030 n7031 ; n7032
g4597 and n6696 n7032_not ; n7033
g4598 nor n6323 n7033 ; n7034
g4599 and n2610_not n7033 ; n7035
g4600 and pi0299 n7017_not ; n7036
g4601 and n7019_not n7036 ; n7037
g4602 and pi0969 n6720 ; n7038
g4603 nor pi0299 n7038 ; n7039
g4604 nor pi0039 n7037 ; n7040
g4605 and n7039_not n7040 ; n7041
g4606 and n2620 n7041 ; n7042
g4607 nor n7035 n7042 ; n7043
g4608 and n2569 n7043 ; n7044
g4609 and pi0054_not n7044 ; n7045
g4610 and pi0074 n7034_not ; n7046
g4611 and n7045_not n7046 ; n7047
g4612 nor n2569 n7033 ; n7048
g4613 nor n7044 n7048 ; n7049
g4614 and pi0054 n7049_not ; n7050
g4615 and pi0075_not n7043 ; n7051
g4616 and pi0075 n7033_not ; n7052
g4617 and pi0092 n7052_not ; n7053
g4618 and n7051_not n7053 ; n7054
g4619 and pi0075 n7043 ; n7055
g4620 and pi0087 n7033 ; n7056
g4621 and n2530_not n7033 ; n7057
g4622 and pi0963 n6745 ; n7058
g4623 and n7036 n7058_not ; n7059
g4624 and pi0969 n6752 ; n7060
g4625 nor pi0299 n7060 ; n7061
g4626 and n2530 n7059_not ; n7062
g4627 and n7061_not n7062 ; n7063
g4628 and pi0100 n7057_not ; n7064
g4629 and n7063_not n7064 ; n7065
g4630 and n6764_not n7030 ; n7066
g4631 and n6761_not n7031 ; n7067
g4632 nor n7066 n7067 ; n7068
g4633 and n6767 n7068_not ; n7069
g4634 and pi0969 n6775 ; n7070
g4635 nor pi0299 n7070 ; n7071
g4636 and n6778 n7018 ; n7072
g4637 and n7036 n7072_not ; n7073
g4638 nor n6781 n7073 ; n7074
g4639 and n6786 n7018 ; n7075
g4640 nor n7017 n7075 ; n7076
g4641 and n6416 n7076_not ; n7077
g4642 nor n7074 n7077 ; n7078
g4643 and pi0232 n7071_not ; n7079
g4644 and n7078_not n7079 ; n7080
g4645 and pi0969 n6769 ; n7081
g4646 nor pi0299 n7081 ; n7082
g4647 nor pi0232 n7073 ; n7083
g4648 and n7082_not n7083 ; n7084
g4649 nor n7080 n7084 ; n7085
g4650 nor pi0039 n7085 ; n7086
g4651 nor pi0038 n7069 ; n7087
g4652 and n7086_not n7087 ; n7088
g4653 and pi0039 n7033 ; n7089
g4654 and pi0038 n7089_not ; n7090
g4655 and n7041_not n7090 ; n7091
g4656 nor n7088 n7091 ; n7092
g4657 nor pi0100 n7092 ; n7093
g4658 nor pi0087 n7065 ; n7094
g4659 and n7093_not n7094 ; n7095
g4660 nor pi0075 n7056 ; n7096
g4661 and n7095_not n7096 ; n7097
g4662 nor pi0092 n7055 ; n7098
g4663 and n7097_not n7098 ; n7099
g4664 nor pi0054 n7054 ; n7100
g4665 and n7099_not n7100 ; n7101
g4666 nor pi0074 n7050 ; n7102
g4667 and n7101_not n7102 ; n7103
g4668 nor pi0055 n7047 ; n7104
g4669 and n7103_not n7104 ; n7105
g4670 and n2529 n7029_not ; n7106
g4671 and n7105_not n7106 ; n7107
g4672 nor pi0059 n7027 ; n7108
g4673 and n7107_not n7108 ; n7109
g4674 nor pi0057 n7026 ; n7110
g4675 and n7109_not n7110 ; n7111
g4676 nor n7023 n7111 ; po0176
g4677 and pi0975 n6696 ; n7113
g4678 and pi0228_not pi0975 ; n7114
g4679 and n6222 n7114 ; n7115
g4680 and n2572 n7115 ; n7116
g4681 and n6305 n7116 ; n7117
g4682 nor n7113 n7117 ; n7118
g4683 and pi0057 n7118_not ; n7119
g4684 and n6304 n7116 ; n7120
g4685 and pi0059 n7113_not ; n7121
g4686 and n7120_not n7121 ; n7122
g4687 and n2529_not n7113 ; n7123
g4688 and pi0055 n7113_not ; n7124
g4689 and n7116_not n7124 ; n7125
g4690 and pi0299_not pi0971 ; n7126
g4691 and pi0299 pi0975 ; n7127
g4692 nor n7126 n7127 ; n7128
g4693 and n6696 n7128_not ; n7129
g4694 nor n6323 n7129 ; n7130
g4695 and n2610_not n7129 ; n7131
g4696 and pi0299 n7113_not ; n7132
g4697 and n7115_not n7132 ; n7133
g4698 and pi0971 n6720 ; n7134
g4699 nor pi0299 n7134 ; n7135
g4700 nor pi0039 n7133 ; n7136
g4701 and n7135_not n7136 ; n7137
g4702 and n2620 n7137 ; n7138
g4703 nor n7131 n7138 ; n7139
g4704 and n2569 n7139 ; n7140
g4705 and pi0054_not n7140 ; n7141
g4706 and pi0074 n7130_not ; n7142
g4707 and n7141_not n7142 ; n7143
g4708 nor n2569 n7129 ; n7144
g4709 nor n7140 n7144 ; n7145
g4710 and pi0054 n7145_not ; n7146
g4711 and pi0075_not n7139 ; n7147
g4712 and pi0075 n7129_not ; n7148
g4713 and pi0092 n7148_not ; n7149
g4714 and n7147_not n7149 ; n7150
g4715 and pi0075 n7139 ; n7151
g4716 and pi0087 n7129 ; n7152
g4717 and n2530_not n7129 ; n7153
g4718 and pi0975 n6745 ; n7154
g4719 and n7132 n7154_not ; n7155
g4720 and pi0971 n6752 ; n7156
g4721 nor pi0299 n7156 ; n7157
g4722 and n2530 n7155_not ; n7158
g4723 and n7157_not n7158 ; n7159
g4724 and pi0100 n7153_not ; n7160
g4725 and n7159_not n7160 ; n7161
g4726 and n6764_not n7126 ; n7162
g4727 and n6761_not n7127 ; n7163
g4728 nor n7162 n7163 ; n7164
g4729 and n6767 n7164_not ; n7165
g4730 and pi0971 n6775 ; n7166
g4731 nor pi0299 n7166 ; n7167
g4732 and n6778 n7114 ; n7168
g4733 and n7132 n7168_not ; n7169
g4734 nor n6781 n7169 ; n7170
g4735 and n6786 n7114 ; n7171
g4736 nor n7113 n7171 ; n7172
g4737 and n6416 n7172_not ; n7173
g4738 nor n7170 n7173 ; n7174
g4739 and pi0232 n7167_not ; n7175
g4740 and n7174_not n7175 ; n7176
g4741 and pi0971 n6769 ; n7177
g4742 nor pi0299 n7177 ; n7178
g4743 nor pi0232 n7169 ; n7179
g4744 and n7178_not n7179 ; n7180
g4745 nor n7176 n7180 ; n7181
g4746 nor pi0039 n7181 ; n7182
g4747 nor pi0038 n7165 ; n7183
g4748 and n7182_not n7183 ; n7184
g4749 and pi0039 n7129 ; n7185
g4750 and pi0038 n7185_not ; n7186
g4751 and n7137_not n7186 ; n7187
g4752 nor n7184 n7187 ; n7188
g4753 nor pi0100 n7188 ; n7189
g4754 nor pi0087 n7161 ; n7190
g4755 and n7189_not n7190 ; n7191
g4756 nor pi0075 n7152 ; n7192
g4757 and n7191_not n7192 ; n7193
g4758 nor pi0092 n7151 ; n7194
g4759 and n7193_not n7194 ; n7195
g4760 nor pi0054 n7150 ; n7196
g4761 and n7195_not n7196 ; n7197
g4762 nor pi0074 n7146 ; n7198
g4763 and n7197_not n7198 ; n7199
g4764 nor pi0055 n7143 ; n7200
g4765 and n7199_not n7200 ; n7201
g4766 and n2529 n7125_not ; n7202
g4767 and n7201_not n7202 ; n7203
g4768 nor pi0059 n7123 ; n7204
g4769 and n7203_not n7204 ; n7205
g4770 nor pi0057 n7122 ; n7206
g4771 and n7205_not n7206 ; n7207
g4772 nor n7119 n7207 ; po0177
g4773 and pi0978 n6696 ; n7209
g4774 and pi0228_not pi0978 ; n7210
g4775 and n2572 n7210 ; n7211
g4776 and n6222 n7211 ; n7212
g4777 and n6305 n7212 ; n7213
g4778 nor n7209 n7213 ; n7214
g4779 and pi0057 n7214_not ; n7215
g4780 and n6304 n7212 ; n7216
g4781 and pi0059 n7209_not ; n7217
g4782 and n7216_not n7217 ; n7218
g4783 and n2529_not n7209 ; n7219
g4784 and pi0055 n7209_not ; n7220
g4785 and n7212_not n7220 ; n7221
g4786 and pi0299_not pi0974 ; n7222
g4787 and pi0299 pi0978 ; n7223
g4788 nor n7222 n7223 ; n7224
g4789 and n6696 n7224_not ; n7225
g4790 nor n6323 n7225 ; n7226
g4791 and n6720 n7224_not ; n7227
g4792 nor pi0228 n2610 ; n7228
g4793 and n7227 n7228_not ; n7229
g4794 and n2569 n7229_not ; n7230
g4795 and pi0054_not n7230 ; n7231
g4796 and pi0074 n7226_not ; n7232
g4797 and n7231_not n7232 ; n7233
g4798 nor n2569 n7225 ; n7234
g4799 nor n7230 n7234 ; n7235
g4800 and pi0054 n7235_not ; n7236
g4801 nor pi0075 n7229 ; n7237
g4802 and pi0075 n7225_not ; n7238
g4803 and pi0092 n7238_not ; n7239
g4804 and n7237_not n7239 ; n7240
g4805 and pi0075 n7229_not ; n7241
g4806 and pi0087 n7225 ; n7242
g4807 and n2530_not n7225 ; n7243
g4808 and pi0299 n7209_not ; n7244
g4809 and pi0978 n6745 ; n7245
g4810 and n7244 n7245_not ; n7246
g4811 and pi0974 n6752 ; n7247
g4812 nor pi0299 n7247 ; n7248
g4813 and n2530 n7246_not ; n7249
g4814 and n7248_not n7249 ; n7250
g4815 and pi0100 n7243_not ; n7251
g4816 and n7250_not n7251 ; n7252
g4817 and pi0039 n7225 ; n7253
g4818 and pi0039_not n7227 ; n7254
g4819 and pi0038 n7253_not ; n7255
g4820 and n7254_not n7255 ; n7256
g4821 and n6764_not n7222 ; n7257
g4822 and n6761_not n7223 ; n7258
g4823 nor n7257 n7258 ; n7259
g4824 and n6767 n7259_not ; n7260
g4825 and pi0974 n6775 ; n7261
g4826 nor pi0299 n7261 ; n7262
g4827 and n6778 n7210 ; n7263
g4828 and n7244 n7263_not ; n7264
g4829 nor n6781 n7264 ; n7265
g4830 and n6786 n7210 ; n7266
g4831 nor n7209 n7266 ; n7267
g4832 and n6416 n7267_not ; n7268
g4833 nor n7265 n7268 ; n7269
g4834 and pi0232 n7262_not ; n7270
g4835 and n7269_not n7270 ; n7271
g4836 and pi0974 n6769 ; n7272
g4837 nor pi0299 n7272 ; n7273
g4838 nor pi0232 n7264 ; n7274
g4839 and n7273_not n7274 ; n7275
g4840 nor n7271 n7275 ; n7276
g4841 nor pi0039 n7276 ; n7277
g4842 nor pi0038 n7260 ; n7278
g4843 and n7277_not n7278 ; n7279
g4844 nor n7256 n7279 ; n7280
g4845 nor pi0100 n7280 ; n7281
g4846 nor pi0087 n7252 ; n7282
g4847 and n7281_not n7282 ; n7283
g4848 nor pi0075 n7242 ; n7284
g4849 and n7283_not n7284 ; n7285
g4850 nor pi0092 n7241 ; n7286
g4851 and n7285_not n7286 ; n7287
g4852 nor pi0054 n7240 ; n7288
g4853 and n7287_not n7288 ; n7289
g4854 nor pi0074 n7236 ; n7290
g4855 and n7289_not n7290 ; n7291
g4856 nor pi0055 n7233 ; n7292
g4857 and n7291_not n7292 ; n7293
g4858 and n2529 n7221_not ; n7294
g4859 and n7293_not n7294 ; n7295
g4860 nor pi0059 n7219 ; n7296
g4861 and n7295_not n7296 ; n7297
g4862 nor pi0057 n7218 ; n7298
g4863 and n7297_not n7298 ; n7299
g4864 nor n7215 n7299 ; po0178
g4865 and n2620 n6284 ; n7301
g4866 and pi0075 n7301_not ; n7302
g4867 and n2533 n2608 ; n7303
g4868 and n6284 n7303 ; n7304
g4869 and pi0092 n7304_not ; n7305
g4870 nor n7302 n7305 ; n7306
g4871 and pi0299 n6244_not ; n7307
g4872 and n6759 n7307 ; n7308
g4873 nor pi0299 n6207 ; n7309
g4874 and n6409 n7309 ; n7310
g4875 and pi0039 n7310_not ; n7311
g4876 and n7308_not n7311 ; n7312
g4877 and pi0299 n6489 ; n7313
g4878 and pi0299_not n6520 ; n7314
g4879 nor pi0232 n7313 ; n7315
g4880 and n7314_not n7315 ; n7316
g4881 and n6527 n6532 ; n7317
g4882 nor pi0299 n6530 ; n7318
g4883 and n6771_not n7318 ; n7319
g4884 and n7317_not n7319 ; n7320
g4885 and n6416_not n7313 ; n7321
g4886 and n6490_not n6781 ; n7322
g4887 and n6785_not n7322 ; n7323
g4888 and pi0232 n7321_not ; n7324
g4889 and n7320_not n7324 ; n7325
g4890 and n7323_not n7325 ; n7326
g4891 nor pi0039 n7316 ; n7327
g4892 and n7326_not n7327 ; n7328
g4893 nor n7312 n7328 ; n7329
g4894 nor pi0038 n7329 ; n7330
g4895 nor n6136 n7330 ; n7331
g4896 nor pi0100 n7331 ; n7332
g4897 and pi0038_not n6284 ; n7333
g4898 and pi0100 n7333_not ; n7334
g4899 and n6289 n7334_not ; n7335
g4900 and n7332_not n7335 ; n7336
g4901 and n2569 n7336_not ; n7337
g4902 and n7306 n7337_not ; n7338
g4903 nor pi0054 n7338 ; n7339
g4904 and pi0092_not n7304 ; n7340
g4905 and pi0054 n7340_not ; n7341
g4906 nor n7339 n7341 ; n7342
g4907 nor pi0074 n7342 ; n7343
g4908 nor n6130 n7343 ; n7344
g4909 nor pi0055 n7344 ; n7345
g4910 and n2535 n6125 ; n7346
g4911 and pi0055 n7346_not ; n7347
g4912 nor pi0056 n7347 ; n7348
g4913 and pi0062_not n7348 ; n7349
g4914 and n7345_not n7349 ; n7350
g4915 and n3328 n7350_not ; n7351
g4916 and n6123 n7351_not ; po0195
g4917 nor pi0954 po0195 ; n7353
g4918 and pi0024 pi0954 ; n7354
g4919 nor n7353 n7354 ; po0182
g4920 and n2531 n3335 ; n7356
g4921 and n3330 n7356 ; n7357
g4922 nor n2441 n7357 ; n7358
g4923 and pi0062 n7358_not ; n7359
g4924 and n2537 n3335 ; n7360
g4925 and pi0056 n2441_not ; n7361
g4926 and n7360_not n7361 ; n7362
g4927 and n2531 n6128 ; n7363
g4928 and n3335 n7363 ; n7364
g4929 and pi0074_not n7364 ; n7365
g4930 nor n2441 n7365 ; n7366
g4931 and pi0055 n7366_not ; n7367
g4932 nor n2441 n2532 ; n7368
g4933 and n3335 n3373 ; n7369
g4934 nor n2441 n7369 ; n7370
g4935 and pi0092 n7370_not ; n7371
g4936 and pi0075 n2441_not ; n7372
g4937 nor n2441 n7356 ; n7373
g4938 and pi0087 n7373_not ; n7374
g4939 and pi0100_not n4730 ; n7375
g4940 and n2521 n6356_not ; n7376
g4941 nor pi0299 n7376 ; n7377
g4942 and pi0299 n3394_not ; n7378
g4943 nor n7377 n7378 ; n7379
g4944 and pi0100 n3335 ; n7380
g4945 and n7379 n7380 ; n7381
g4946 nor pi0039 n7381 ; n7382
g4947 and n7375_not n7382 ; n7383
g4948 and pi0100_not n3335 ; n7384
g4949 and pi0039 n7384_not ; n7385
g4950 nor pi0038 n7385 ; n7386
g4951 and n7383_not n7386 ; n7387
g4952 nor n2441 n7387 ; n7388
g4953 nor pi0087 n7388 ; n7389
g4954 nor pi0075 n7374 ; n7390
g4955 and n7389_not n7390 ; n7391
g4956 nor pi0092 n7372 ; n7392
g4957 and n7391_not n7392 ; n7393
g4958 and n2532 n7371_not ; n7394
g4959 and n7393_not n7394 ; n7395
g4960 nor pi0055 n7368 ; n7396
g4961 and n7395_not n7396 ; n7397
g4962 nor pi0056 n7367 ; n7398
g4963 and n7397_not n7398 ; n7399
g4964 nor pi0062 n7362 ; n7400
g4965 and n7399_not n7400 ; n7401
g4966 nor n7359 n7401 ; n7402
g4967 and n3328 n7402_not ; n7403
g4968 and n2441 n3328_not ; n7404
g4969 or n7403 n7404 ; po0183
g4970 and pi0119 pi1056 ; n7406
g4971 and pi0228_not pi0252 ; n7407
g4972 nor pi0119 n7407 ; n7408
g4973 nor pi0468 n7408 ; n7409
g4974 nand n7406_not n7409 ; po0184
g4975 and pi0119 pi1077 ; n7411
g4976 nand n7409 n7411_not ; po0185
g4977 and pi0119 pi1073 ; n7413
g4978 nand n7409 n7413_not ; po0186
g4979 and pi0119 pi1041 ; n7415
g4980 nand n7409 n7415_not ; po0187
g4981 and pi0824 n2932 ; n7417
g4982 and pi0122_not pi1093 ; n7418
g4983 and n7417 n7418 ; n7419
g4984 and pi1091_not n7419 ; n7420
g4985 and pi0098_not n7420 ; n7421
g4986 and pi0567 n7421 ; n7422
g4987 nor pi0285 pi0286 ; n7423
g4988 and pi0289_not n7423 ; n7424
g4989 and pi0288_not n7424 ; n7425
g4990 nand pi0057_not n6305 ; po1038
g4991 and n7425_not po1038 ; n7427
g4992 and n7422 n7427 ; n7428
g4993 and pi0074_not n6134 ; n7429
g4994 and pi0122_not pi0829 ; n7430
g4995 and n2961 n6157_not ; n7431
g4996 and pi0841_not n2703 ; n7432
g4997 and pi0090 n7432 ; n7433
g4998 nor pi0093 n7433 ; n7434
g4999 and n7431 n7434_not ; n7435
g5000 nor pi0051 n7435 ; n7436
g5001 and pi0088_not pi0098 ; n7437
g5002 nor pi0050 pi0077 ; n7438
g5003 and pi0094_not n7438 ; n7439
g5004 and n2767 n7439 ; n7440
g5005 and n2495 n7437 ; n7441
g5006 and n7440 n7441 ; n7442
g5007 nor pi0097 n7442 ; n7443
g5008 and n2717 n7443_not ; n7444
g5009 and pi0035_not n2704 ; n7445
g5010 and pi0070_not n7445 ; n7446
g5011 and n7444 n7446 ; n7447
g5012 and n7436 n7447_not ; n7448
g5013 nor n2747 n7448 ; n7449
g5014 and pi0096_not n2519 ; n7450
g5015 and n7449 n7450 ; n7451
g5016 and n6277 n7451 ; n7452
g5017 and n7430_not n7452 ; n7453
g5018 nor pi0096 n7449 ; n7454
g5019 and pi0096 n6484_not ; n7455
g5020 and n2519 n7455_not ; n7456
g5021 and n2932 n7430 ; n7457
g5022 and n7456 n7457 ; n7458
g5023 and n7454_not n7458 ; n7459
g5024 nor n7453 n7459 ; n7460
g5025 nor pi1093 n7460 ; n7461
g5026 nor pi0087 n7461 ; n7462
g5027 and n2521 po0740 ; n7463
g5028 and pi0087 n7463_not ; n7464
g5029 and pi0075_not n2531 ; n7465
g5030 and n7464_not n7465 ; n7466
g5031 and n7462_not n7466 ; n7467
g5032 nor pi0567 n7467 ; n7468
g5033 and n7429 n7468_not ; n7469
g5034 nor pi0299 n2669 ; n7470
g5035 and pi0299 n2639_not ; n7471
g5036 nor n7470 n7471 ; n7472
g5037 and pi0232 n6197 ; n7473
g5038 and n7472 n7473 ; n7474
g5039 and n2610 n7474_not ; n7475
g5040 and n7421 n7475_not ; n7476
g5041 and pi0024_not n6359 ; n7477
g5042 and n2923_not po1057 ; n7478
g5043 and pi1093 n7457 ; n7479
g5044 and n7478 n7479 ; n7480
g5045 and n7477 n7480 ; n7481
g5046 and pi1091 n7481_not ; n7482
g5047 and n7475 n7482_not ; n7483
g5048 and pi0098_not n7417 ; n7484
g5049 and n7418 n7484 ; n7485
g5050 nor pi1091 n7485 ; n7486
g5051 and n7483 n7486_not ; n7487
g5052 and pi0075 n7476_not ; n7488
g5053 and n7487_not n7488 ; n7489
g5054 and pi1093 n2923 ; n7490
g5055 and n6277 n7490_not ; n7491
g5056 and n2521 n7491 ; n7492
g5057 and pi1091 n7492_not ; n7493
g5058 nor pi1091 n7463 ; n7494
g5059 and n2521 n7417 ; n7495
g5060 and pi0122 n7495 ; n7496
g5061 and pi0122_not n7484 ; n7497
g5062 nor n7496 n7497 ; n7498
g5063 and pi1093 n7498_not ; n7499
g5064 and n7494 n7499_not ; n7500
g5065 and n2625 n7493_not ; n7501
g5066 and n7500_not n7501 ; n7502
g5067 nor n7421 n7502 ; n7503
g5068 and pi0087 n7503_not ; n7504
g5069 and n2530_not n7421 ; n7505
g5070 and pi0228 n7474_not ; n7506
g5071 nor n7421 n7506 ; n7507
g5072 and n2521 n7480 ; n7508
g5073 and pi1091 n7508_not ; n7509
g5074 nor n7486 n7509 ; n7510
g5075 and n7506 n7510_not ; n7511
g5076 and n2530 n7507_not ; n7512
g5077 and n7511_not n7512 ; n7513
g5078 and pi0100 n7505_not ; n7514
g5079 and n7513_not n7514 ; n7515
g5080 and pi0038 n7421 ; n7516
g5081 and pi1093 n2923_not ; n7517
g5082 and n2747_not n7450 ; n7518
g5083 and n7436_not n7518 ; n7519
g5084 and n7417 n7519 ; n7520
g5085 and pi0829_not n7520 ; n7521
g5086 and pi0024_not n2756 ; n7522
g5087 and pi0046_not pi0097 ; n7523
g5088 and pi0108_not n7523 ; n7524
g5089 and n6491 n7524 ; n7525
g5090 and n2772 n7525 ; n7526
g5091 and pi0091_not n7526 ; n7527
g5092 nor n7522 n7527 ; n7528
g5093 and n2461 n7431 ; n7529
g5094 and n7528_not n7529 ; n7530
g5095 and n7436 n7530_not ; n7531
g5096 nor n2747 n7531 ; n7532
g5097 nor pi0096 n7532 ; n7533
g5098 and n2933 n7456 ; n7534
g5099 and n7533_not n7534 ; n7535
g5100 nor n7521 n7535 ; n7536
g5101 nor pi0122 n7536 ; n7537
g5102 and pi0122 n6277 ; n7538
g5103 and n7519 n7538 ; n7539
g5104 nor n7537 n7539 ; n7540
g5105 and n7517 n7540_not ; n7541
g5106 and pi1091 n7541_not ; n7542
g5107 and n7461_not n7542 ; n7543
g5108 nor pi0039 n7543 ; n7544
g5109 nor pi1091 n7461 ; n7545
g5110 and pi0122 n7520 ; n7546
g5111 nor n7497 n7546 ; n7547
g5112 and pi1093 n7547_not ; n7548
g5113 and n7545 n7548_not ; n7549
g5114 and n7544 n7549_not ; n7550
g5115 and pi0223_not n5810 ; n7551
g5116 and n7421 n7551_not ; n7552
g5117 and n2923_not n2925 ; n7553
g5118 and n6382 n7553 ; n7554
g5119 and n2926 n7554 ; n7555
g5120 and pi1091 n7555_not ; n7556
g5121 nor n7486 n7556 ; n7557
g5122 and n6198 n7557 ; n7558
g5123 and n6198_not n7421 ; n7559
g5124 nor n7558 n7559 ; n7560
g5125 and n6205 n7560 ; n7561
g5126 and n6227_not n7557 ; n7562
g5127 and n6227 n7421 ; n7563
g5128 nor n7562 n7563 ; n7564
g5129 and n6205_not n7564 ; n7565
g5130 and n7551 n7561_not ; n7566
g5131 and n7565_not n7566 ; n7567
g5132 nor pi0299 n7552 ; n7568
g5133 and n7567_not n7568 ; n7569
g5134 and pi0216_not n6379 ; n7570
g5135 and n7421 n7570_not ; n7571
g5136 and n6242 n7560 ; n7572
g5137 and n6242_not n7564 ; n7573
g5138 and n7570 n7572_not ; n7574
g5139 and n7573_not n7574 ; n7575
g5140 and pi0299 n7571_not ; n7576
g5141 and n7575_not n7576 ; n7577
g5142 and pi0039 n7569_not ; n7578
g5143 and n7577_not n7578 ; n7579
g5144 nor n7550 n7579 ; n7580
g5145 nor pi0038 n7580 ; n7581
g5146 nor pi0100 n7516 ; n7582
g5147 and n7581_not n7582 ; n7583
g5148 nor pi0087 n7515 ; n7584
g5149 and n7583_not n7584 ; n7585
g5150 nor pi0075 n7504 ; n7586
g5151 and n7585_not n7586 ; n7587
g5152 nor n7489 n7587 ; n7588
g5153 and pi0567 n7588_not ; n7589
g5154 and n7469 n7589_not ; n7590
g5155 and n7422 n7429_not ; n7591
g5156 nor n7590 n7591 ; n7592
g5157 and n7425_not n7592 ; n7593
g5158 and pi1091 n7478 ; n7594
g5159 and n7457 n7594 ; n7595
g5160 and n7477 n7595 ; n7596
g5161 and pi1093 n7596 ; n7597
g5162 and n7475 n7597 ; n7598
g5163 and pi0075 n7598_not ; n7599
g5164 nor n7543 n7545 ; n7600
g5165 nor pi0039 n7600 ; n7601
g5166 and pi1091 n7555 ; n7602
g5167 and n6244_not n7602 ; n7603
g5168 and pi0216_not n6640 ; n7604
g5169 and n7603 n7604 ; n7605
g5170 and n6207_not n7602 ; n7606
g5171 and pi0299_not n6405 ; n7607
g5172 and pi0224_not n7607 ; n7608
g5173 and n7606 n7608 ; n7609
g5174 and pi0039 n7605_not ; n7610
g5175 and n7609_not n7610 ; n7611
g5176 nor pi0038 n7611 ; n7612
g5177 and n7601_not n7612 ; n7613
g5178 nor pi0100 n7613 ; n7614
g5179 and n6384 n7519 ; n7615
g5180 and n7612 n7615 ; n7616
g5181 and n7542_not n7616 ; n7617
g5182 and n7614 n7617_not ; n7618
g5183 and pi1091 n7508 ; n7619
g5184 and pi0228 n7619 ; n7620
g5185 and n2530 n7474_not ; n7621
g5186 and n7620 n7621 ; n7622
g5187 and pi0100 n7622_not ; n7623
g5188 nor n7618 n7623 ; n7624
g5189 nor pi0087 n7624 ; n7625
g5190 and pi1091_not pi1093 ; n7626
g5191 and n7495_not n7626 ; n7627
g5192 nor n7492 n7626 ; n7628
g5193 and n2625 n7628_not ; n7629
g5194 and n7627_not n7629 ; n7630
g5195 and pi0087 n7630_not ; n7631
g5196 nor n7625 n7631 ; n7632
g5197 nor pi0075 n7632 ; n7633
g5198 nor n7599 n7633 ; n7634
g5199 and pi0567 n7634_not ; n7635
g5200 and n7469 n7635_not ; n7636
g5201 and n7425 n7636_not ; n7637
g5202 nor po1038 n7593 ; n7638
g5203 and n7637_not n7638 ; n7639
g5204 and pi0217 n7428_not ; n7640
g5205 and n7639_not n7640 ; n7641
g5206 nor pi1161 pi1162 ; n7642
g5207 and pi1163_not n7642 ; n7643
g5208 and pi0592_not n7422 ; n7644
g5209 and pi0592 n7422 ; n7645
g5210 nor pi0363 pi0372 ; n7646
g5211 and pi0363 pi0372 ; n7647
g5212 nor n7646 n7647 ; n7648
g5213 and pi0386 n7648_not ; n7649
g5214 and pi0386_not n7648 ; n7650
g5215 nor n7649 n7650 ; n7651
g5216 and pi0338 pi0388_not ; n7652
g5217 and pi0338_not pi0388 ; n7653
g5218 nor n7652 n7653 ; n7654
g5219 and pi0337 pi0339_not ; n7655
g5220 and pi0337_not pi0339 ; n7656
g5221 nor n7655 n7656 ; n7657
g5222 and pi0387 n7657 ; n7658
g5223 nor pi0387 n7657 ; n7659
g5224 nor n7658 n7659 ; n7660
g5225 and pi0380 n7660_not ; n7661
g5226 and pi0380_not n7660 ; n7662
g5227 nor n7661 n7662 ; n7663
g5228 and n7654 n7663_not ; n7664
g5229 and n7654_not n7663 ; n7665
g5230 nor n7664 n7665 ; n7666
g5231 and n7651 n7666 ; n7667
g5232 nor n7651 n7666 ; n7668
g5233 nor n7667 n7668 ; n7669
g5234 and pi1196 n7669_not ; n7670
g5235 nor pi0368 pi0389 ; n7671
g5236 and pi0368 pi0389 ; n7672
g5237 nor n7671 n7672 ; n7673
g5238 and pi0365 pi0447_not ; n7674
g5239 and pi0365_not pi0447 ; n7675
g5240 nor n7674 n7675 ; n7676
g5241 and pi0336 pi0383_not ; n7677
g5242 and pi0336_not pi0383 ; n7678
g5243 nor n7677 n7678 ; n7679
g5244 and pi0364 pi0366_not ; n7680
g5245 and pi0364_not pi0366 ; n7681
g5246 nor n7680 n7681 ; n7682
g5247 and n7679 n7682 ; n7683
g5248 nor n7679 n7682 ; n7684
g5249 nor n7683 n7684 ; n7685
g5250 and n7676 n7685 ; n7686
g5251 nor n7676 n7685 ; n7687
g5252 nor n7686 n7687 ; n7688
g5253 and pi0367 n7688_not ; n7689
g5254 and pi0367_not n7688 ; n7690
g5255 nor n7689 n7690 ; n7691
g5256 and n7673 n7691 ; n7692
g5257 nor n7673 n7691 ; n7693
g5258 and pi1197 n7692_not ; n7694
g5259 and n7693_not n7694 ; n7695
g5260 nor n7670 n7695 ; n7696
g5261 and pi0592 n7696_not ; n7697
g5262 and pi0379 pi0382_not ; n7698
g5263 and pi0379_not pi0382 ; n7699
g5264 nor n7698 n7699 ; n7700
g5265 and pi0376 pi0439_not ; n7701
g5266 and pi0376_not pi0439 ; n7702
g5267 nor n7701 n7702 ; n7703
g5268 and pi0381 n7703 ; n7704
g5269 nor pi0381 n7703 ; n7705
g5270 nor n7704 n7705 ; n7706
g5271 and pi0317 pi0385_not ; n7707
g5272 and pi0317_not pi0385 ; n7708
g5273 nor n7707 n7708 ; n7709
g5274 and pi0378 n7709 ; n7710
g5275 nor pi0378 n7709 ; n7711
g5276 nor n7710 n7711 ; n7712
g5277 and n7706 n7712_not ; n7713
g5278 and n7706_not n7712 ; n7714
g5279 nor n7713 n7714 ; n7715
g5280 and n7700 n7715 ; n7716
g5281 nor n7700 n7715 ; n7717
g5282 nor n7716 n7717 ; n7718
g5283 nor pi0377 n7718 ; n7719
g5284 and pi0377 n7718 ; n7720
g5285 nor n7719 n7720 ; n7721
g5286 and n7696 n7721_not ; n7722
g5287 and pi0592 n7722_not ; n7723
g5288 and n7422 n7723_not ; n7724
g5289 and pi1199 n7724_not ; n7725
g5290 nor n7697 n7725 ; n7726
g5291 and n7645 n7726 ; n7727
g5292 and pi1198_not n7727 ; n7728
g5293 and pi0384 pi0442_not ; n7729
g5294 and pi0384_not pi0442 ; n7730
g5295 nor n7729 n7730 ; n7731
g5296 and pi0440 n7731_not ; n7732
g5297 and pi0440_not n7731 ; n7733
g5298 nor n7732 n7733 ; n7734
g5299 nor pi0369 pi0374 ; n7735
g5300 and pi0369 pi0374 ; n7736
g5301 nor n7735 n7736 ; n7737
g5302 nor pi0370 n7737 ; n7738
g5303 and pi0370 n7737 ; n7739
g5304 nor n7738 n7739 ; n7740
g5305 nor pi0371 n7740 ; n7741
g5306 and pi0371 n7740 ; n7742
g5307 nor n7741 n7742 ; n7743
g5308 nor pi0373 n7743 ; n7744
g5309 and pi0373 n7743 ; n7745
g5310 nor n7744 n7745 ; n7746
g5311 and pi0375 n7746_not ; n7747
g5312 and pi0375_not n7746 ; n7748
g5313 nor n7747 n7748 ; n7749
g5314 nor n7734 n7749 ; n7750
g5315 and n7734 n7749 ; n7751
g5316 nor n7750 n7751 ; n7752
g5317 and n7727 n7752 ; n7753
g5318 nor n7644 n7728 ; n7754
g5319 and n7753_not n7754 ; n7755
g5320 nor pi0590 n7755 ; n7756
g5321 and pi0351 pi1199 ; n7757
g5322 and pi0345 pi0346_not ; n7758
g5323 and pi0345_not pi0346 ; n7759
g5324 nor n7758 n7759 ; n7760
g5325 and pi0323 n7760_not ; n7761
g5326 and pi0323_not n7760 ; n7762
g5327 nor n7761 n7762 ; n7763
g5328 and pi0358 pi0450_not ; n7764
g5329 and pi0358_not pi0450 ; n7765
g5330 nor n7764 n7765 ; n7766
g5331 and n7763 n7766_not ; n7767
g5332 and n7763_not n7766 ; n7768
g5333 nor n7767 n7768 ; n7769
g5334 nor pi0327 pi0362 ; n7770
g5335 and pi0327 pi0362 ; n7771
g5336 nor n7770 n7771 ; n7772
g5337 and pi0343 pi0344_not ; n7773
g5338 and pi0343_not pi0344 ; n7774
g5339 nor n7773 n7774 ; n7775
g5340 and n7772 n7775_not ; n7776
g5341 and n7772_not n7775 ; n7777
g5342 nor n7776 n7777 ; n7778
g5343 and n7769 n7778 ; n7779
g5344 nor n7769 n7778 ; n7780
g5345 and pi1197 n7779_not ; n7781
g5346 and n7780_not n7781 ; n7782
g5347 and pi0320 pi0460_not ; n7783
g5348 and pi0320_not pi0460 ; n7784
g5349 nor n7783 n7784 ; n7785
g5350 and pi0342 n7785_not ; n7786
g5351 and pi0342_not n7785 ; n7787
g5352 nor n7786 n7787 ; n7788
g5353 and pi0452 pi0455_not ; n7789
g5354 and pi0452_not pi0455 ; n7790
g5355 nor n7789 n7790 ; n7791
g5356 and pi0355 n7791 ; n7792
g5357 nor pi0355 n7791 ; n7793
g5358 nor n7792 n7793 ; n7794
g5359 and pi0361 pi0458_not ; n7795
g5360 and pi0361_not pi0458 ; n7796
g5361 nor n7795 n7796 ; n7797
g5362 and n7794 n7797 ; n7798
g5363 nor n7794 n7797 ; n7799
g5364 nor n7798 n7799 ; n7800
g5365 and pi0441_not n7800 ; n7801
g5366 and pi0441 n7800_not ; n7802
g5367 nor pi0592 n7801 ; n7803
g5368 and n7802_not n7803 ; n7804
g5369 and n7422 n7788 ; n7805
g5370 and n7804_not n7805 ; n7806
g5371 and pi0361 pi0441_not ; n7807
g5372 and pi0361_not pi0441 ; n7808
g5373 nor n7807 n7808 ; n7809
g5374 and n7788 n7809 ; n7810
g5375 nor n7788 n7809 ; n7811
g5376 nor n7810 n7811 ; n7812
g5377 and pi0458 n7812 ; n7813
g5378 nor pi0458 n7812 ; n7814
g5379 nor n7813 n7814 ; n7815
g5380 and n7794 n7815 ; n7816
g5381 nor n7794 n7815 ; n7817
g5382 nor n7816 n7817 ; n7818
g5383 and pi0592_not n7818 ; n7819
g5384 and n7422 n7788_not ; n7820
g5385 and n7819_not n7820 ; n7821
g5386 and pi1196 n7806_not ; n7822
g5387 and n7821_not n7822 ; n7823
g5388 nor pi1198 n7823 ; n7824
g5389 and pi1196 n7818 ; n7825
g5390 and pi0321 pi0347_not ; n7826
g5391 and pi0321_not pi0347 ; n7827
g5392 nor n7826 n7827 ; n7828
g5393 and pi0316 pi0349_not ; n7829
g5394 and pi0316_not pi0349 ; n7830
g5395 nor n7829 n7830 ; n7831
g5396 and pi0348 n7831 ; n7832
g5397 nor pi0348 n7831 ; n7833
g5398 nor n7832 n7833 ; n7834
g5399 and pi0315 pi0359_not ; n7835
g5400 and pi0315_not pi0359 ; n7836
g5401 nor n7835 n7836 ; n7837
g5402 and pi0322 n7837 ; n7838
g5403 nor pi0322 n7837 ; n7839
g5404 nor n7838 n7839 ; n7840
g5405 and n7834 n7840_not ; n7841
g5406 and n7834_not n7840 ; n7842
g5407 nor n7841 n7842 ; n7843
g5408 and n7828 n7843 ; n7844
g5409 nor n7828 n7843 ; n7845
g5410 nor n7844 n7845 ; n7846
g5411 and pi0350 n7846_not ; n7847
g5412 and pi0350_not n7846 ; n7848
g5413 nor n7847 n7848 ; n7849
g5414 and n7825_not n7849 ; n7850
g5415 and pi1198 n7644 ; n7851
g5416 and n7850 n7851 ; n7852
g5417 nor n7824 n7852 ; n7853
g5418 nor n7782 n7853 ; n7854
g5419 nor pi0592 n7854 ; n7855
g5420 and n7422 n7855_not ; n7856
g5421 nor n7757 n7856 ; n7857
g5422 and pi1199 n7645_not ; n7858
g5423 and pi0351 n7858 ; n7859
g5424 nor n7857 n7859 ; n7860
g5425 nor pi0461 n7860 ; n7861
g5426 and pi0351_not pi1199 ; n7862
g5427 nor n7856 n7862 ; n7863
g5428 and pi0351_not n7858 ; n7864
g5429 nor n7863 n7864 ; n7865
g5430 and pi0461 n7865_not ; n7866
g5431 nor n7861 n7866 ; n7867
g5432 nor pi0357 n7867 ; n7868
g5433 nor pi0461 n7865 ; n7869
g5434 and pi0461 n7860_not ; n7870
g5435 nor n7869 n7870 ; n7871
g5436 and pi0357 n7871_not ; n7872
g5437 nor n7868 n7872 ; n7873
g5438 nor pi0356 n7873 ; n7874
g5439 nor pi0357 n7871 ; n7875
g5440 and pi0357 n7867_not ; n7876
g5441 nor n7875 n7876 ; n7877
g5442 and pi0356 n7877_not ; n7878
g5443 and pi0360 pi0462_not ; n7879
g5444 and pi0360_not pi0462 ; n7880
g5445 nor n7879 n7880 ; n7881
g5446 and pi0352 pi0353_not ; n7882
g5447 and pi0352_not pi0353 ; n7883
g5448 nor n7882 n7883 ; n7884
g5449 and n7881 n7884 ; n7885
g5450 nor n7881 n7884 ; n7886
g5451 nor n7885 n7886 ; n7887
g5452 and pi0354 n7887_not ; n7888
g5453 and pi0354_not n7887 ; n7889
g5454 nor n7888 n7889 ; n7890
g5455 and n7874_not n7890 ; n7891
g5456 and n7878_not n7891 ; n7892
g5457 nor pi0356 n7877 ; n7893
g5458 and pi0356 n7873_not ; n7894
g5459 nor n7890 n7893 ; n7895
g5460 and n7894_not n7895 ; n7896
g5461 nor n7892 n7896 ; n7897
g5462 and pi0590 n7897_not ; n7898
g5463 nor pi0591 n7756 ; n7899
g5464 and n7898_not n7899 ; n7900
g5465 and pi0590 n7422 ; n7901
g5466 and pi1197 n7645_not ; n7902
g5467 and pi0318 pi0409_not ; n7903
g5468 and pi0318_not pi0409 ; n7904
g5469 nor n7903 n7904 ; n7905
g5470 and pi0401 pi0402_not ; n7906
g5471 and pi0401_not pi0402 ; n7907
g5472 nor n7906 n7907 ; n7908
g5473 and pi0406 n7908 ; n7909
g5474 nor pi0406 n7908 ; n7910
g5475 nor n7909 n7910 ; n7911
g5476 nor pi0403 pi0405 ; n7912
g5477 and pi0403 pi0405 ; n7913
g5478 nor n7912 n7913 ; n7914
g5479 and pi0325 pi0326_not ; n7915
g5480 and pi0325_not pi0326 ; n7916
g5481 nor n7915 n7916 ; n7917
g5482 and n7914 n7917 ; n7918
g5483 nor n7914 n7917 ; n7919
g5484 nor n7918 n7919 ; n7920
g5485 and n7911 n7920_not ; n7921
g5486 and n7911_not n7920 ; n7922
g5487 nor n7921 n7922 ; n7923
g5488 and n7905 n7923 ; n7924
g5489 nor n7905 n7923 ; n7925
g5490 nor n7924 n7925 ; n7926
g5491 and n7485 n7926_not ; n7927
g5492 and pi1091_not n7927 ; n7928
g5493 and pi0567 n7928 ; n7929
g5494 and pi0390 pi0410_not ; n7930
g5495 and pi0390_not pi0410 ; n7931
g5496 nor n7930 n7931 ; n7932
g5497 and pi0397 pi0412_not ; n7933
g5498 and pi0397_not pi0412 ; n7934
g5499 nor n7933 n7934 ; n7935
g5500 and pi0404 n7935 ; n7936
g5501 nor pi0404 n7935 ; n7937
g5502 nor n7936 n7937 ; n7938
g5503 and pi0319 pi0324_not ; n7939
g5504 and pi0319_not pi0324 ; n7940
g5505 nor n7939 n7940 ; n7941
g5506 and pi0456 n7941_not ; n7942
g5507 and pi0456_not n7941 ; n7943
g5508 nor n7942 n7943 ; n7944
g5509 and n7938 n7944_not ; n7945
g5510 and n7938_not n7944 ; n7946
g5511 nor n7945 n7946 ; n7947
g5512 and n7932 n7947 ; n7948
g5513 nor n7932 n7947 ; n7949
g5514 nor n7948 n7949 ; n7950
g5515 and pi0411 n7950 ; n7951
g5516 nor pi0411 n7950 ; n7952
g5517 nor n7951 n7952 ; n7953
g5518 and pi1196 n7953_not ; n7954
g5519 and pi0592_not n7929 ; n7955
g5520 and n7954_not n7955 ; n7956
g5521 and n7858 n7956_not ; n7957
g5522 and pi0592_not pi1196 ; n7958
g5523 and n7422 n7958_not ; n7959
g5524 and n7485 n7953 ; n7960
g5525 and pi1091_not n7960 ; n7961
g5526 and pi0567 n7961 ; n7962
g5527 and n7958 n7962 ; n7963
g5528 nor pi1199 n7959 ; n7964
g5529 and n7963_not n7964 ; n7965
g5530 nor n7957 n7965 ; n7966
g5531 nor pi1197 n7966 ; n7967
g5532 nor n7902 n7967 ; n7968
g5533 and pi0333 n7968_not ; n7969
g5534 and pi1198 n7645_not ; n7970
g5535 and n7966 n7970_not ; n7971
g5536 and pi0328 pi0408_not ; n7972
g5537 and pi0328_not pi0408 ; n7973
g5538 nor n7972 n7973 ; n7974
g5539 nor pi0394 pi0396 ; n7975
g5540 and pi0394 pi0396 ; n7976
g5541 nor n7975 n7976 ; n7977
g5542 and n7974 n7977_not ; n7978
g5543 and n7974_not n7977 ; n7979
g5544 nor n7978 n7979 ; n7980
g5545 and pi0398 pi0399_not ; n7981
g5546 and pi0398_not pi0399 ; n7982
g5547 nor n7981 n7982 ; n7983
g5548 and pi0395 n7983 ; n7984
g5549 nor pi0395 n7983 ; n7985
g5550 nor n7984 n7985 ; n7986
g5551 and pi0329 n7986_not ; n7987
g5552 and pi0329_not n7986 ; n7988
g5553 nor n7987 n7988 ; n7989
g5554 and pi0400 n7989_not ; n7990
g5555 and pi0400_not n7989 ; n7991
g5556 nor n7990 n7991 ; n7992
g5557 and n7980 n7992 ; n7993
g5558 nor n7980 n7992 ; n7994
g5559 nor n7993 n7994 ; n7995
g5560 nor n7971 n7995 ; n7996
g5561 nor pi0333 n7966 ; n7997
g5562 nor n7996 n7997 ; n7998
g5563 and n7969_not n7998 ; n7999
g5564 nor pi0391 n7999 ; n8000
g5565 nor pi0333 n7968 ; n8001
g5566 and n7966 n7996_not ; n8002
g5567 and n8001_not n8002 ; n8003
g5568 and pi0391 n8003_not ; n8004
g5569 nor n8000 n8004 ; n8005
g5570 nor pi0392 n8005 ; n8006
g5571 nor pi0391 n8003 ; n8007
g5572 and pi0391 n7999_not ; n8008
g5573 nor n8007 n8008 ; n8009
g5574 and pi0392 n8009_not ; n8010
g5575 nor n8006 n8010 ; n8011
g5576 nor pi0393 n8011 ; n8012
g5577 nor pi0392 n8009 ; n8013
g5578 and pi0392 n8005_not ; n8014
g5579 nor n8013 n8014 ; n8015
g5580 and pi0393 n8015_not ; n8016
g5581 and pi0407 pi0463_not ; n8017
g5582 and pi0407_not pi0463 ; n8018
g5583 nor n8017 n8018 ; n8019
g5584 and pi0335 pi0413_not ; n8020
g5585 and pi0335_not pi0413 ; n8021
g5586 nor n8020 n8021 ; n8022
g5587 and n8019 n8022 ; n8023
g5588 nor n8019 n8022 ; n8024
g5589 nor n8023 n8024 ; n8025
g5590 and pi0334 n8025_not ; n8026
g5591 and pi0334_not n8025 ; n8027
g5592 nor n8026 n8027 ; n8028
g5593 and n8012_not n8028 ; n8029
g5594 and n8016_not n8029 ; n8030
g5595 nor pi0393 n8015 ; n8031
g5596 and pi0393 n8011_not ; n8032
g5597 nor n8028 n8031 ; n8033
g5598 and n8032_not n8033 ; n8034
g5599 nor n8030 n8034 ; n8035
g5600 nor pi0590 n8035 ; n8036
g5601 and pi0591 n7901_not ; n8037
g5602 and n8036_not n8037 ; n8038
g5603 nor n7900 n8038 ; n8039
g5604 nor pi0588 n8039 ; n8040
g5605 nor pi0590 pi0591 ; n8041
g5606 and n7422 n8041_not ; n8042
g5607 nor pi0417 pi0418 ; n8043
g5608 and pi0417 pi0418 ; n8044
g5609 nor n8043 n8044 ; n8045
g5610 and pi0437 n8045 ; n8046
g5611 nor pi0437 n8045 ; n8047
g5612 nor n8046 n8047 ; n8048
g5613 and pi0453 pi0464_not ; n8049
g5614 and pi0453_not pi0464 ; n8050
g5615 nor n8049 n8050 ; n8051
g5616 and n8048 n8051 ; n8052
g5617 nor n8048 n8051 ; n8053
g5618 nor n8052 n8053 ; n8054
g5619 and pi0415 pi0431_not ; n8055
g5620 and pi0415_not pi0431 ; n8056
g5621 nor n8055 n8056 ; n8057
g5622 and pi0416 pi0438_not ; n8058
g5623 and pi0416_not pi0438 ; n8059
g5624 nor n8058 n8059 ; n8060
g5625 and n8057 n8060 ; n8061
g5626 nor n8057 n8060 ; n8062
g5627 nor n8061 n8062 ; n8063
g5628 and n8054 n8063_not ; n8064
g5629 and n8054_not n8063 ; n8065
g5630 and pi1197 n8064_not ; n8066
g5631 and n8065_not n8066 ; n8067
g5632 and pi0421 pi0454_not ; n8068
g5633 and pi0421_not pi0454 ; n8069
g5634 nor n8068 n8069 ; n8070
g5635 and pi0432 pi0459_not ; n8071
g5636 and pi0432_not pi0459 ; n8072
g5637 nor n8071 n8072 ; n8073
g5638 and n8070 n8073_not ; n8074
g5639 and n8070_not n8073 ; n8075
g5640 nor n8074 n8075 ; n8076
g5641 nor pi0419 pi0420 ; n8077
g5642 and pi0419 pi0420 ; n8078
g5643 nor n8077 n8078 ; n8079
g5644 and pi0423 pi0424_not ; n8080
g5645 and pi0423_not pi0424 ; n8081
g5646 nor n8080 n8081 ; n8082
g5647 and n8079 n8082_not ; n8083
g5648 and n8079_not n8082 ; n8084
g5649 nor n8083 n8084 ; n8085
g5650 and n8076 n8085 ; n8086
g5651 nor n8076 n8085 ; n8087
g5652 nor n8086 n8087 ; n8088
g5653 and pi0425 n8088_not ; n8089
g5654 and pi0425_not n8088 ; n8090
g5655 and pi1198 n8089_not ; n8091
g5656 and n8090_not n8091 ; n8092
g5657 nor n8067 n8092 ; n8093
g5658 nor pi0429 pi0435 ; n8094
g5659 and pi0429 pi0435 ; n8095
g5660 nor n8094 n8095 ; n8096
g5661 and pi0434 pi0446_not ; n8097
g5662 and pi0434_not pi0446 ; n8098
g5663 nor n8097 n8098 ; n8099
g5664 and pi0414 pi0422_not ; n8100
g5665 and pi0414_not pi0422 ; n8101
g5666 nor n8100 n8101 ; n8102
g5667 and n8099 n8102 ; n8103
g5668 nor n8099 n8102 ; n8104
g5669 nor n8103 n8104 ; n8105
g5670 and n8096 n8105 ; n8106
g5671 nor n8096 n8105 ; n8107
g5672 nor n8106 n8107 ; n8108
g5673 and pi0436 pi0443_not ; n8109
g5674 and pi0436_not pi0443 ; n8110
g5675 nor n8109 n8110 ; n8111
g5676 and pi0444_not n8111 ; n8112
g5677 and pi0444 n8111_not ; n8113
g5678 nor n8112 n8113 ; n8114
g5679 nor n8108 n8114 ; n8115
g5680 and n8108 n8114 ; n8116
g5681 and n7958 n8115_not ; n8117
g5682 and n8116_not n8117 ; n8118
g5683 and n8093 n8118_not ; n8119
g5684 and n7644 n8119 ; n8120
g5685 nor pi1199 n7645 ; n8121
g5686 and n8120_not n8121 ; n8122
g5687 and pi0433 pi0451_not ; n8123
g5688 and pi0433_not pi0451 ; n8124
g5689 nor n8123 n8124 ; n8125
g5690 and pi0449 n8125 ; n8126
g5691 nor pi0449 n8125 ; n8127
g5692 nor n8126 n8127 ; n8128
g5693 and pi0427_not pi0428 ; n8129
g5694 and pi0427 pi0428_not ; n8130
g5695 nor n8129 n8130 ; n8131
g5696 and pi0430 n8131_not ; n8132
g5697 and pi0430_not n8131 ; n8133
g5698 nor n8132 n8133 ; n8134
g5699 nor pi0426 n8134 ; n8135
g5700 and pi0426 n8134 ; n8136
g5701 nor n8135 n8136 ; n8137
g5702 nor pi0445 n8137 ; n8138
g5703 and pi0445 n8137 ; n8139
g5704 nor n8138 n8139 ; n8140
g5705 nor pi0448 n8140 ; n8141
g5706 and pi0448 n8140 ; n8142
g5707 nor n8141 n8142 ; n8143
g5708 and n8120 n8143_not ; n8144
g5709 nor n7645 n8144 ; n8145
g5710 and n8128 n8145_not ; n8146
g5711 and n8120 n8143 ; n8147
g5712 nor n7645 n8147 ; n8148
g5713 nor n8128 n8148 ; n8149
g5714 and pi1199 n8146_not ; n8150
g5715 and n8149_not n8150 ; n8151
g5716 and n8041 n8122_not ; n8152
g5717 and n8151_not n8152 ; n8153
g5718 and pi0588 n8042_not ; n8154
g5719 and n8153_not n8154 ; n8155
g5720 and n7427 n8155_not ; n8156
g5721 and n8040_not n8156 ; n8157
g5722 and n7636 n8041_not ; n8158
g5723 nor pi0087 n7623 ; n8159
g5724 and n7614_not n8159 ; n8160
g5725 and pi0087 pi0100_not ; n8161
g5726 and n2530 n8161 ; n8162
g5727 and n7493_not n8162 ; n8163
g5728 and n7494_not n8163 ; n8164
g5729 nor pi0075 n8164 ; n8165
g5730 and n8160_not n8165 ; n8166
g5731 nor n7599 n8166 ; n8167
g5732 and pi0567 n8167_not ; n8168
g5733 and n7469 n8168_not ; n8169
g5734 nor pi0592 n8169 ; n8170
g5735 and pi0592 n7636_not ; n8171
g5736 nor n8170 n8171 ; n8172
g5737 and n8093_not n8172 ; n8173
g5738 nor pi1196 n7636 ; n8174
g5739 nor pi0443 pi0592 ; n8175
g5740 nor n7636 n8175 ; n8176
g5741 and n8169_not n8175 ; n8177
g5742 nor n8176 n8177 ; n8178
g5743 nor pi0444 n8178 ; n8179
g5744 and pi0443 pi0592_not ; n8180
g5745 nor n7636 n8180 ; n8181
g5746 and n8169_not n8180 ; n8182
g5747 nor n8181 n8182 ; n8183
g5748 and pi0444 n8183_not ; n8184
g5749 nor n8179 n8184 ; n8185
g5750 nor pi0436 n8185 ; n8186
g5751 nor pi0444 n8183 ; n8187
g5752 and pi0444 n8178_not ; n8188
g5753 nor n8187 n8188 ; n8189
g5754 and pi0436 n8189_not ; n8190
g5755 and n8108 n8186_not ; n8191
g5756 and n8190_not n8191 ; n8192
g5757 nor pi0436 n8189 ; n8193
g5758 and pi0436 n8185_not ; n8194
g5759 nor n8108 n8193 ; n8195
g5760 and n8194_not n8195 ; n8196
g5761 and pi1196 n8192_not ; n8197
g5762 and n8196_not n8197 ; n8198
g5763 and n8093 n8174_not ; n8199
g5764 and n8198_not n8199 ; n8200
g5765 nor n8173 n8200 ; n8201
g5766 and pi1199_not n8201 ; n8202
g5767 and pi0428 n8201_not ; n8203
g5768 and pi0428_not n8172 ; n8204
g5769 nor n8203 n8204 ; n8205
g5770 nor pi0427 n8205 ; n8206
g5771 nor pi0428 n8201 ; n8207
g5772 and pi0428 n8172 ; n8208
g5773 nor n8207 n8208 ; n8209
g5774 and pi0427 n8209_not ; n8210
g5775 nor n8206 n8210 ; n8211
g5776 and pi0430 n8211_not ; n8212
g5777 nor pi0427 n8209 ; n8213
g5778 and pi0427 n8205_not ; n8214
g5779 nor n8213 n8214 ; n8215
g5780 nor pi0430 n8215 ; n8216
g5781 nor n8212 n8216 ; n8217
g5782 and pi0426 n8217_not ; n8218
g5783 and pi0430 n8215_not ; n8219
g5784 nor pi0430 n8211 ; n8220
g5785 nor n8219 n8220 ; n8221
g5786 nor pi0426 n8221 ; n8222
g5787 nor n8218 n8222 ; n8223
g5788 and pi0445 n8223_not ; n8224
g5789 and pi0426 n8221_not ; n8225
g5790 nor pi0426 n8217 ; n8226
g5791 nor n8225 n8226 ; n8227
g5792 nor pi0445 n8227 ; n8228
g5793 nor n8224 n8228 ; n8229
g5794 and pi0448 n8128_not ; n8230
g5795 and pi0448_not n8128 ; n8231
g5796 nor n8230 n8231 ; n8232
g5797 nor n8229 n8232 ; n8233
g5798 and pi0445 n8227_not ; n8234
g5799 nor pi0445 n8223 ; n8235
g5800 nor n8234 n8235 ; n8236
g5801 and n8232 n8236_not ; n8237
g5802 and pi1199 n8233_not ; n8238
g5803 and n8237_not n8238 ; n8239
g5804 and n8041 n8202_not ; n8240
g5805 and n8239_not n8240 ; n8241
g5806 and n7425 n8158_not ; n8242
g5807 and n8241_not n8242 ; n8243
g5808 nor n7592 n8041 ; n8244
g5809 and pi1196_not n7592 ; n8245
g5810 and n7592 n8175_not ; n8246
g5811 and pi0436_not pi0444 ; n8247
g5812 and pi0436 pi0444_not ; n8248
g5813 nor n8247 n8248 ; n8249
g5814 and n8108 n8249_not ; n8250
g5815 and n8108_not n8249 ; n8251
g5816 nor n8250 n8251 ; n8252
g5817 and n8177_not n8252 ; n8253
g5818 and n8246_not n8253 ; n8254
g5819 and n7592 n8180_not ; n8255
g5820 nor n8182 n8252 ; n8256
g5821 and n8255_not n8256 ; n8257
g5822 and pi1196 n8254_not ; n8258
g5823 and n8257_not n8258 ; n8259
g5824 nor n8245 n8259 ; n8260
g5825 and n8093 n8260_not ; n8261
g5826 and pi0592 n7592 ; n8262
g5827 nor n8170 n8262 ; n8263
g5828 nor n8093 n8263 ; n8264
g5829 nor n8261 n8264 ; n8265
g5830 nor pi1199 n8265 ; n8266
g5831 and pi0428_not n8263 ; n8267
g5832 and pi0428 n8265 ; n8268
g5833 and pi0427 n8267_not ; n8269
g5834 and n8268_not n8269 ; n8270
g5835 and pi0428_not n8265 ; n8271
g5836 and pi0428 n8263 ; n8272
g5837 nor pi0427 n8272 ; n8273
g5838 and n8271_not n8273 ; n8274
g5839 nor n8270 n8274 ; n8275
g5840 nor pi0430 n8275 ; n8276
g5841 and n8131 n8263 ; n8277
g5842 and n8131_not n8265 ; n8278
g5843 nor n8277 n8278 ; n8279
g5844 and pi0430 n8279 ; n8280
g5845 nor n8276 n8280 ; n8281
g5846 nor pi0426 n8281 ; n8282
g5847 and pi0430 n8275_not ; n8283
g5848 and pi0430_not n8279 ; n8284
g5849 nor n8283 n8284 ; n8285
g5850 and pi0426 n8285_not ; n8286
g5851 nor n8282 n8286 ; n8287
g5852 nor pi0445 n8287 ; n8288
g5853 nor pi0426 n8285 ; n8289
g5854 and pi0426 n8281_not ; n8290
g5855 nor n8289 n8290 ; n8291
g5856 and pi0445 n8291_not ; n8292
g5857 nor n8288 n8292 ; n8293
g5858 and pi0448 n8293 ; n8294
g5859 nor pi0445 n8291 ; n8295
g5860 and pi0445 n8287_not ; n8296
g5861 nor n8295 n8296 ; n8297
g5862 and pi0448_not n8297 ; n8298
g5863 nor n8128 n8294 ; n8299
g5864 and n8298_not n8299 ; n8300
g5865 and pi0448_not n8293 ; n8301
g5866 and pi0448 n8297 ; n8302
g5867 and n8128 n8301_not ; n8303
g5868 and n8302_not n8303 ; n8304
g5869 nor n8300 n8304 ; n8305
g5870 and pi1199 n8305_not ; n8306
g5871 and n8041 n8266_not ; n8307
g5872 and n8306_not n8307 ; n8308
g5873 nor n7425 n8244 ; n8309
g5874 and n8308_not n8309 ; n8310
g5875 nor n8243 n8310 ; n8311
g5876 and pi0588 n8311_not ; n8312
g5877 and pi0591 n7636 ; n8313
g5878 and n7825 n8172_not ; n8314
g5879 nor pi0350 pi0592 ; n8315
g5880 nor n7636 n8315 ; n8316
g5881 and n8169_not n8315 ; n8317
g5882 and n7846 n8317_not ; n8318
g5883 and n8316_not n8318 ; n8319
g5884 and pi0350 pi0592_not ; n8320
g5885 nor n7636 n8320 ; n8321
g5886 and n8169_not n8320 ; n8322
g5887 nor n7846 n8322 ; n8323
g5888 and n8321_not n8323 ; n8324
g5889 nor n7825 n8319 ; n8325
g5890 and n8324_not n8325 ; n8326
g5891 and pi1198 n8314_not ; n8327
g5892 and n8326_not n8327 ; n8328
g5893 nor pi0455 n8172 ; n8329
g5894 and pi0455 n7636_not ; n8330
g5895 nor n8329 n8330 ; n8331
g5896 nor pi0452 n8331 ; n8332
g5897 and pi0455 n8172_not ; n8333
g5898 nor pi0455 n7636 ; n8334
g5899 nor n8333 n8334 ; n8335
g5900 and pi0452 n8335_not ; n8336
g5901 nor n8332 n8336 ; n8337
g5902 nor pi0355 n8337 ; n8338
g5903 nor pi0452 n8335 ; n8339
g5904 and pi0452 n8331_not ; n8340
g5905 nor n8339 n8340 ; n8341
g5906 and pi0355 n8341_not ; n8342
g5907 nor n8338 n8342 ; n8343
g5908 and pi0458 n8343_not ; n8344
g5909 nor pi0355 n8341 ; n8345
g5910 and pi0355 n8337_not ; n8346
g5911 nor n8345 n8346 ; n8347
g5912 nor pi0458 n8347 ; n8348
g5913 and n7812 n8344_not ; n8349
g5914 and n8348_not n8349 ; n8350
g5915 and pi0458 n8347_not ; n8351
g5916 nor pi0458 n8343 ; n8352
g5917 nor n7812 n8351 ; n8353
g5918 and n8352_not n8353 ; n8354
g5919 and pi1196 n8350_not ; n8355
g5920 and n8354_not n8355 ; n8356
g5921 nor pi1198 n8174 ; n8357
g5922 and n8356_not n8357 ; n8358
g5923 nor n8328 n8358 ; n8359
g5924 nor n7782 n8359 ; n8360
g5925 and n7782 n8172 ; n8361
g5926 nor n8360 n8361 ; n8362
g5927 and n7862_not n8362 ; n8363
g5928 and pi1199 n8172_not ; n8364
g5929 and pi0351_not n8364 ; n8365
g5930 nor n8363 n8365 ; n8366
g5931 nor pi0461 n8366 ; n8367
g5932 and n7757_not n8362 ; n8368
g5933 and pi0351 n8364 ; n8369
g5934 nor n8368 n8369 ; n8370
g5935 and pi0461 n8370_not ; n8371
g5936 nor n8367 n8371 ; n8372
g5937 nor pi0357 n8372 ; n8373
g5938 nor pi0461 n8370 ; n8374
g5939 and pi0461 n8366_not ; n8375
g5940 nor n8374 n8375 ; n8376
g5941 and pi0357 n8376_not ; n8377
g5942 nor n8373 n8377 ; n8378
g5943 nor pi0356 n8378 ; n8379
g5944 nor pi0357 n8376 ; n8380
g5945 and pi0357 n8372_not ; n8381
g5946 nor n8380 n8381 ; n8382
g5947 and pi0356 n8382_not ; n8383
g5948 nor n8379 n8383 ; n8384
g5949 nor n7890 n8384 ; n8385
g5950 nor pi0356 n8382 ; n8386
g5951 and pi0356 n8378_not ; n8387
g5952 nor n8386 n8387 ; n8388
g5953 and n7890 n8388_not ; n8389
g5954 nor pi0591 n8385 ; n8390
g5955 and n8389_not n8390 ; n8391
g5956 and pi0590 n8313_not ; n8392
g5957 and n8391_not n8392 ; n8393
g5958 and pi1197 n8172_not ; n8394
g5959 and pi1198 n7995_not ; n8395
g5960 and n8172 n8395 ; n8396
g5961 and pi0075_not n7954 ; n8397
g5962 nor n7926 n8397 ; n8398
g5963 and n7617 n8398 ; n8399
g5964 and n7614 n8399_not ; n8400
g5965 and n8159 n8400_not ; n8401
g5966 and n7628_not n8162 ; n8402
g5967 and n7495 n7926_not ; n8403
g5968 and n7626 n8403_not ; n8404
g5969 and n8402 n8404_not ; n8405
g5970 and pi1196_not n8405 ; n8406
g5971 and n7495 n7953 ; n8407
g5972 and n7626 n8407_not ; n8408
g5973 and n8405 n8408_not ; n8409
g5974 nor pi0075 pi0592 ; n8410
g5975 and pi1199 n8410 ; n8411
g5976 and n8406_not n8411 ; n8412
g5977 and n8409_not n8412 ; n8413
g5978 and n8401_not n8413 ; n8414
g5979 nor n7634 n8410 ; n8415
g5980 and n8402 n8408_not ; n8416
g5981 and n7617 n7953 ; n8417
g5982 and n7614 n8417_not ; n8418
g5983 and n8159 n8418_not ; n8419
g5984 and pi1196 n8410 ; n8420
g5985 and n8416_not n8420 ; n8421
g5986 and n8419_not n8421 ; n8422
g5987 and pi1196_not n7633 ; n8423
g5988 nor n8422 n8423 ; n8424
g5989 nor pi1199 n8424 ; n8425
g5990 nor n8414 n8415 ; n8426
g5991 and n8425_not n8426 ; n8427
g5992 and pi0567 n8427_not ; n8428
g5993 and n7469 n8395_not ; n8429
g5994 and n8428_not n8429 ; n8430
g5995 nor n8396 n8430 ; n8431
g5996 and pi1197_not n8431 ; n8432
g5997 nor n8394 n8432 ; n8433
g5998 and pi0333 n8433_not ; n8434
g5999 and pi0333_not n8431 ; n8435
g6000 nor n8434 n8435 ; n8436
g6001 and pi0391 n8436_not ; n8437
g6002 and pi0333 n8431_not ; n8438
g6003 and pi0333_not n8433 ; n8439
g6004 nor n8438 n8439 ; n8440
g6005 and pi0391_not n8440 ; n8441
g6006 nor n8437 n8441 ; n8442
g6007 nor pi0392 n8442 ; n8443
g6008 nor pi0391 n8436 ; n8444
g6009 and pi0391 n8440 ; n8445
g6010 nor n8444 n8445 ; n8446
g6011 and pi0392 n8446_not ; n8447
g6012 nor n8443 n8447 ; n8448
g6013 nor pi0393 n8448 ; n8449
g6014 nor pi0392 n8446 ; n8450
g6015 and pi0392 n8442_not ; n8451
g6016 nor n8450 n8451 ; n8452
g6017 and pi0393 n8452_not ; n8453
g6018 nor n8449 n8453 ; n8454
g6019 and pi0334_not n8454 ; n8455
g6020 nor pi0393 n8452 ; n8456
g6021 and pi0393 n8448_not ; n8457
g6022 nor n8456 n8457 ; n8458
g6023 and pi0334 n8458 ; n8459
g6024 and n8025 n8455_not ; n8460
g6025 and n8459_not n8460 ; n8461
g6026 and pi0334_not n8458 ; n8462
g6027 and pi0334 n8454 ; n8463
g6028 nor n8025 n8462 ; n8464
g6029 and n8463_not n8464 ; n8465
g6030 and pi0591 n8461_not ; n8466
g6031 and n8465_not n8466 ; n8467
g6032 and pi0377 pi0592 ; n8468
g6033 nor n7636 n8468 ; n8469
g6034 and n8169_not n8468 ; n8470
g6035 nor n7718 n8470 ; n8471
g6036 and n8469_not n8471 ; n8472
g6037 and pi0377_not pi0592 ; n8473
g6038 nor n7636 n8473 ; n8474
g6039 and n8169_not n8473 ; n8475
g6040 and n7718 n8475_not ; n8476
g6041 and n8474_not n8476 ; n8477
g6042 nor n8472 n8477 ; n8478
g6043 and n7696 n8478_not ; n8479
g6044 and pi0592 n8169_not ; n8480
g6045 nor pi0592 n7636 ; n8481
g6046 nor n8480 n8481 ; n8482
g6047 and n7696_not n8482 ; n8483
g6048 nor n8479 n8483 ; n8484
g6049 and pi1199 n8484 ; n8485
g6050 and n7636 n7695_not ; n8486
g6051 and n7695 n8482 ; n8487
g6052 nor n8486 n8487 ; n8488
g6053 and n7669 n8488_not ; n8489
g6054 nor pi1196 n7695 ; n8490
g6055 and n8482 n8490_not ; n8491
g6056 and pi1196_not n8486 ; n8492
g6057 nor n8491 n8492 ; n8493
g6058 nor n7669 n8493 ; n8494
g6059 nor pi1199 n8489 ; n8495
g6060 and n8494_not n8495 ; n8496
g6061 nor n8485 n8496 ; n8497
g6062 nor pi0374 n8497 ; n8498
g6063 and pi1198_not pi1199 ; n8499
g6064 and n8484 n8499 ; n8500
g6065 and pi1198_not n8496 ; n8501
g6066 and pi1198 n8482_not ; n8502
g6067 nor n8500 n8502 ; n8503
g6068 and n8501_not n8503 ; n8504
g6069 and pi0374 n8504_not ; n8505
g6070 nor n8498 n8505 ; n8506
g6071 and pi0369 n8506_not ; n8507
g6072 nor pi0374 n8504 ; n8508
g6073 and pi0374 n8497_not ; n8509
g6074 nor n8508 n8509 ; n8510
g6075 nor pi0369 n8510 ; n8511
g6076 nor n8507 n8511 ; n8512
g6077 nor pi0370 n8512 ; n8513
g6078 nor pi0369 n8506 ; n8514
g6079 and pi0369 n8510_not ; n8515
g6080 nor n8514 n8515 ; n8516
g6081 and pi0370 n8516_not ; n8517
g6082 nor n8513 n8517 ; n8518
g6083 nor pi0371 n8518 ; n8519
g6084 nor pi0370 n8516 ; n8520
g6085 and pi0370 n8512_not ; n8521
g6086 nor n8520 n8521 ; n8522
g6087 and pi0371 n8522_not ; n8523
g6088 nor n8519 n8523 ; n8524
g6089 nor pi0373 n8524 ; n8525
g6090 nor pi0371 n8522 ; n8526
g6091 and pi0371 n8518_not ; n8527
g6092 nor n8526 n8527 ; n8528
g6093 and pi0373 n8528_not ; n8529
g6094 nor n8525 n8529 ; n8530
g6095 and pi0375_not n8530 ; n8531
g6096 nor pi0373 n8528 ; n8532
g6097 and pi0373 n8524_not ; n8533
g6098 nor n8532 n8533 ; n8534
g6099 and pi0375 n8534 ; n8535
g6100 and n7734 n8531_not ; n8536
g6101 and n8535_not n8536 ; n8537
g6102 and pi0375 n8530 ; n8538
g6103 and pi0375_not n8534 ; n8539
g6104 nor n7734 n8538 ; n8540
g6105 and n8539_not n8540 ; n8541
g6106 nor pi0591 n8537 ; n8542
g6107 and n8541_not n8542 ; n8543
g6108 nor pi0590 n8467 ; n8544
g6109 and n8543_not n8544 ; n8545
g6110 and n7425 n8545_not ; n8546
g6111 and n8393_not n8546 ; n8547
g6112 and pi0591 n7592_not ; n8548
g6113 and n7782 n8263_not ; n8549
g6114 and n7825 n8263_not ; n8550
g6115 and n7592 n8320_not ; n8551
g6116 and n8323 n8551_not ; n8552
g6117 and n7592 n8315_not ; n8553
g6118 and n8318 n8553_not ; n8554
g6119 nor n7825 n8552 ; n8555
g6120 and n8554_not n8555 ; n8556
g6121 and pi1198 n8550_not ; n8557
g6122 and n8556_not n8557 ; n8558
g6123 and pi0455 n8263_not ; n8559
g6124 and pi0455_not n7592 ; n8560
g6125 nor n8559 n8560 ; n8561
g6126 nor pi0452 n8561 ; n8562
g6127 nor pi0455 n8263 ; n8563
g6128 and pi0455 n7592 ; n8564
g6129 nor n8563 n8564 ; n8565
g6130 and pi0452 n8565_not ; n8566
g6131 and pi0355 n7815_not ; n8567
g6132 and pi0355_not n7815 ; n8568
g6133 nor n8567 n8568 ; n8569
g6134 nor n8562 n8569 ; n8570
g6135 and n8566_not n8570 ; n8571
g6136 nor pi0452 n8565 ; n8572
g6137 and pi0452 n8561_not ; n8573
g6138 and n8569 n8572_not ; n8574
g6139 and n8573_not n8574 ; n8575
g6140 and pi1196 n8571_not ; n8576
g6141 and n8575_not n8576 ; n8577
g6142 nor pi1198 n8245 ; n8578
g6143 and n8577_not n8578 ; n8579
g6144 nor n7782 n8558 ; n8580
g6145 and n8579_not n8580 ; n8581
g6146 nor n8549 n8581 ; n8582
g6147 nor n7862 n8582 ; n8583
g6148 and pi1199 n8263_not ; n8584
g6149 and pi0351_not n8584 ; n8585
g6150 nor n8583 n8585 ; n8586
g6151 nor pi0461 n8586 ; n8587
g6152 nor n7757 n8582 ; n8588
g6153 and pi0351 n8584 ; n8589
g6154 nor n8588 n8589 ; n8590
g6155 and pi0461 n8590_not ; n8591
g6156 nor n8587 n8591 ; n8592
g6157 nor pi0357 n8592 ; n8593
g6158 nor pi0461 n8590 ; n8594
g6159 and pi0461 n8586_not ; n8595
g6160 nor n8594 n8595 ; n8596
g6161 and pi0357 n8596_not ; n8597
g6162 nor n8593 n8597 ; n8598
g6163 nor pi0356 n8598 ; n8599
g6164 nor pi0357 n8596 ; n8600
g6165 and pi0357 n8592_not ; n8601
g6166 nor n8600 n8601 ; n8602
g6167 and pi0356 n8602_not ; n8603
g6168 nor n8599 n8603 ; n8604
g6169 nor n7890 n8604 ; n8605
g6170 nor pi0356 n8602 ; n8606
g6171 and pi0356 n8598_not ; n8607
g6172 nor n8606 n8607 ; n8608
g6173 and n7890 n8608_not ; n8609
g6174 nor pi0591 n8605 ; n8610
g6175 and n8609_not n8610 ; n8611
g6176 and pi0590 n8548_not ; n8612
g6177 and n8611_not n8612 ; n8613
g6178 and n7429_not n7962 ; n8614
g6179 and pi0038 n7961 ; n8615
g6180 nor pi0100 n8615 ; n8616
g6181 and n7545 n7953_not ; n8617
g6182 and n7550 n8617_not ; n8618
g6183 and n7570_not n7961 ; n8619
g6184 and pi0299 n8619_not ; n8620
g6185 and n6227_not n7602 ; n8621
g6186 nor n7961 n8621 ; n8622
g6187 and n6242_not n8622 ; n8623
g6188 and n6198 n7602 ; n8624
g6189 nor n7961 n8624 ; n8625
g6190 and n6242 n8625 ; n8626
g6191 and n7570 n8623_not ; n8627
g6192 and n8626_not n8627 ; n8628
g6193 and n8620 n8628_not ; n8629
g6194 and n7551_not n7961 ; n8630
g6195 nor pi0299 n8630 ; n8631
g6196 and n6205_not n8622 ; n8632
g6197 and n6205 n8625 ; n8633
g6198 and n7551 n8632_not ; n8634
g6199 and n8633_not n8634 ; n8635
g6200 and n8631 n8635_not ; n8636
g6201 and pi0039 n8629_not ; n8637
g6202 and n8636_not n8637 ; n8638
g6203 nor n8618 n8638 ; n8639
g6204 nor pi0038 n8639 ; n8640
g6205 and n8616 n8640_not ; n8641
g6206 and n7623 n7961_not ; n8642
g6207 nor n8641 n8642 ; n8643
g6208 nor pi0087 n8643 ; n8644
g6209 and n2625_not n7961 ; n8645
g6210 and pi0087 n8645_not ; n8646
g6211 and n7494 n7953_not ; n8647
g6212 and n7502 n8647_not ; n8648
g6213 and n8646 n8648_not ; n8649
g6214 nor n8644 n8649 ; n8650
g6215 nor pi0075 n8650 ; n8651
g6216 and n7475_not n7961 ; n8652
g6217 and pi0075 n8652_not ; n8653
g6218 nor pi1091 n7960 ; n8654
g6219 and n7483 n8654_not ; n8655
g6220 and n8653 n8655_not ; n8656
g6221 nor n8651 n8656 ; n8657
g6222 and pi0567 n8657_not ; n8658
g6223 and n7469 n8658_not ; n8659
g6224 and n7958 n8614_not ; n8660
g6225 and n8659_not n8660 ; n8661
g6226 nor pi1199 n8245 ; n8662
g6227 and n8661_not n8662 ; n8663
g6228 and n7484 n7926_not ; n8664
g6229 and n8614 n8664 ; n8665
g6230 and n7958 n8665_not ; n8666
g6231 and n7429_not n7929 ; n8667
g6232 nor pi0592 pi1196 ; n8668
g6233 and n8667_not n8668 ; n8669
g6234 nor n8666 n8669 ; n8670
g6235 nor n7469 n8670 ; n8671
g6236 and n7570_not n7928 ; n8672
g6237 and pi0299 n8672_not ; n8673
g6238 nor n8620 n8673 ; n8674
g6239 and n7926_not n7961 ; n8675
g6240 nor n8624 n8675 ; n8676
g6241 and n6242 n8676 ; n8677
g6242 nor n8621 n8675 ; n8678
g6243 and n6242_not n8678 ; n8679
g6244 and n7570 n8677_not ; n8680
g6245 and n8679_not n8680 ; n8681
g6246 nor n8674 n8681 ; n8682
g6247 and n7551_not n7928 ; n8683
g6248 nor pi0299 n8683 ; n8684
g6249 nor n8631 n8684 ; n8685
g6250 and n6205 n8676 ; n8686
g6251 and n6205_not n8678 ; n8687
g6252 and n7551 n8686_not ; n8688
g6253 and n8687_not n8688 ; n8689
g6254 nor n8685 n8689 ; n8690
g6255 and pi0039 n8682_not ; n8691
g6256 and n8690_not n8691 ; n8692
g6257 and n7520 n7926_not ; n8693
g6258 and pi0122 n8693_not ; n8694
g6259 nor pi0122 n8664 ; n8695
g6260 and pi1093 n8695_not ; n8696
g6261 and n8694_not n8696 ; n8697
g6262 and n7545 n8697_not ; n8698
g6263 and n8618 n8698_not ; n8699
g6264 nor n8692 n8699 ; n8700
g6265 nor pi0038 n8700 ; n8701
g6266 and pi0038 n7928 ; n8702
g6267 nor pi0100 n8702 ; n8703
g6268 nor n8616 n8703 ; n8704
g6269 nor n8701 n8704 ; n8705
g6270 and n2530_not n8675 ; n8706
g6271 nor pi0232 n8675 ; n8707
g6272 and n7620_not n8707 ; n8708
g6273 and n6197 n7471_not ; n8709
g6274 nor n7470 n8709 ; n8710
g6275 and pi0228 n8710 ; n8711
g6276 and n8675 n8711_not ; n8712
g6277 and n7470 n7619 ; n8713
g6278 nor pi1091 n8675 ; n8714
g6279 and n8710 n8714_not ; n8715
g6280 and n7509_not n8715 ; n8716
g6281 nor n8713 n8716 ; n8717
g6282 and pi0228 n8717_not ; n8718
g6283 and pi0232 n8712_not ; n8719
g6284 and n8718_not n8719 ; n8720
g6285 and n2530 n8708_not ; n8721
g6286 and n8720_not n8721 ; n8722
g6287 and pi0100 n8706_not ; n8723
g6288 and n8722_not n8723 ; n8724
g6289 nor n8705 n8724 ; n8725
g6290 nor pi0087 n8725 ; n8726
g6291 and n2625_not n7928 ; n8727
g6292 and pi0087 n8727_not ; n8728
g6293 nor n8646 n8728 ; n8729
g6294 and n7494 n7926 ; n8730
g6295 and n7502 n8730_not ; n8731
g6296 and n8647_not n8731 ; n8732
g6297 nor n8729 n8732 ; n8733
g6298 nor n8726 n8733 ; n8734
g6299 nor pi0075 n8734 ; n8735
g6300 and n7475_not n7928 ; n8736
g6301 and pi0075 n8736_not ; n8737
g6302 nor n8653 n8737 ; n8738
g6303 and n7483 n8714_not ; n8739
g6304 nor n8738 n8739 ; n8740
g6305 nor n8735 n8740 ; n8741
g6306 and n8666 n8741_not ; n8742
g6307 and n8728 n8731_not ; n8743
g6308 and n7623 n7928_not ; n8744
g6309 and n7544 n8698_not ; n8745
g6310 nor n7928 n8621 ; n8746
g6311 and n6242_not n8746 ; n8747
g6312 nor n7928 n8624 ; n8748
g6313 and n6242 n8748 ; n8749
g6314 and n7570 n8747_not ; n8750
g6315 and n8749_not n8750 ; n8751
g6316 and n8673 n8751_not ; n8752
g6317 and n6205_not n8746 ; n8753
g6318 and n6205 n8748 ; n8754
g6319 and n7551 n8753_not ; n8755
g6320 and n8754_not n8755 ; n8756
g6321 and n8684 n8756_not ; n8757
g6322 and pi0039 n8752_not ; n8758
g6323 and n8757_not n8758 ; n8759
g6324 nor n8745 n8759 ; n8760
g6325 nor pi0038 n8760 ; n8761
g6326 and n8703 n8761_not ; n8762
g6327 nor n8744 n8762 ; n8763
g6328 nor pi0087 n8763 ; n8764
g6329 nor n8743 n8764 ; n8765
g6330 nor pi0075 n8765 ; n8766
g6331 nor pi1091 n7927 ; n8767
g6332 and n7483 n8767_not ; n8768
g6333 and n8737 n8768_not ; n8769
g6334 nor n8766 n8769 ; n8770
g6335 and n8669 n8770_not ; n8771
g6336 nor n8742 n8771 ; n8772
g6337 and pi0567 n8772_not ; n8773
g6338 and pi1199 n8671_not ; n8774
g6339 and n8773_not n8774 ; n8775
g6340 nor n8395 n8663 ; n8776
g6341 and n8775_not n8776 ; n8777
g6342 and n8170 n8395 ; n8778
g6343 nor n8262 n8778 ; n8779
g6344 and n8777_not n8779 ; n8780
g6345 nor pi1197 n8780 ; n8781
g6346 and pi1197 n8263_not ; n8782
g6347 nor n8781 n8782 ; n8783
g6348 nor pi0333 n8783 ; n8784
g6349 and pi0333 n8780_not ; n8785
g6350 nor n8784 n8785 ; n8786
g6351 nor pi0391 n8786 ; n8787
g6352 nor pi0333 n8780 ; n8788
g6353 and pi0333 n8783_not ; n8789
g6354 nor n8788 n8789 ; n8790
g6355 and pi0391 n8790_not ; n8791
g6356 nor n8787 n8791 ; n8792
g6357 nor pi0392 n8792 ; n8793
g6358 nor pi0391 n8790 ; n8794
g6359 and pi0391 n8786_not ; n8795
g6360 nor n8794 n8795 ; n8796
g6361 and pi0392 n8796_not ; n8797
g6362 nor n8793 n8797 ; n8798
g6363 and pi0393 n8028 ; n8799
g6364 nor pi0393 n8028 ; n8800
g6365 nor n8799 n8800 ; n8801
g6366 nor n8798 n8801 ; n8802
g6367 nor pi0392 n8796 ; n8803
g6368 and pi0392 n8792_not ; n8804
g6369 nor n8803 n8804 ; n8805
g6370 and n8801 n8805_not ; n8806
g6371 and pi0591 n8802_not ; n8807
g6372 and n8806_not n8807 ; n8808
g6373 and pi0592_not n7592 ; n8809
g6374 nor n8480 n8809 ; n8810
g6375 and n7696_not n8810 ; n8811
g6376 and n7592_not n7696 ; n8812
g6377 nor pi1199 n8812 ; n8813
g6378 and n8811_not n8813 ; n8814
g6379 and n7592 n8473_not ; n8815
g6380 and n8476 n8815_not ; n8816
g6381 and n7592 n8468_not ; n8817
g6382 and n8471 n8817_not ; n8818
g6383 nor n8816 n8818 ; n8819
g6384 and n7696 n8819_not ; n8820
g6385 and pi1199 n8811_not ; n8821
g6386 and n8820_not n8821 ; n8822
g6387 nor n8814 n8822 ; n8823
g6388 nor pi0374 n8823 ; n8824
g6389 nor pi1198 n8823 ; n8825
g6390 and pi1198 n8810_not ; n8826
g6391 nor n8825 n8826 ; n8827
g6392 and pi0374 n8827_not ; n8828
g6393 nor n8824 n8828 ; n8829
g6394 and pi0369 n8829_not ; n8830
g6395 nor pi0374 n8827 ; n8831
g6396 and pi0374 n8823_not ; n8832
g6397 nor n8831 n8832 ; n8833
g6398 nor pi0369 n8833 ; n8834
g6399 nor n8830 n8834 ; n8835
g6400 nor pi0370 n8835 ; n8836
g6401 nor pi0369 n8829 ; n8837
g6402 and pi0369 n8833_not ; n8838
g6403 nor n8837 n8838 ; n8839
g6404 and pi0370 n8839_not ; n8840
g6405 nor n8836 n8840 ; n8841
g6406 nor pi0371 n8841 ; n8842
g6407 nor pi0370 n8839 ; n8843
g6408 and pi0370 n8835_not ; n8844
g6409 nor n8843 n8844 ; n8845
g6410 and pi0371 n8845_not ; n8846
g6411 nor n8842 n8846 ; n8847
g6412 and pi0375 n7734 ; n8848
g6413 nor pi0375 n7734 ; n8849
g6414 nor n8848 n8849 ; n8850
g6415 and pi0373 n8850_not ; n8851
g6416 and pi0373_not n8850 ; n8852
g6417 nor n8851 n8852 ; n8853
g6418 nor n8847 n8853 ; n8854
g6419 nor pi0371 n8845 ; n8855
g6420 and pi0371 n8841_not ; n8856
g6421 nor n8855 n8856 ; n8857
g6422 and n8853 n8857_not ; n8858
g6423 nor pi0591 n8854 ; n8859
g6424 and n8858_not n8859 ; n8860
g6425 nor pi0590 n8808 ; n8861
g6426 and n8860_not n8861 ; n8862
g6427 nor n7425 n8862 ; n8863
g6428 and n8613_not n8863 ; n8864
g6429 nor pi0588 n8864 ; n8865
g6430 and n8547_not n8865 ; n8866
g6431 nor po1038 n8312 ; n8867
g6432 and n8866_not n8867 ; n8868
g6433 nor pi0217 n8157 ; n8869
g6434 and n8868_not n8869 ; n8870
g6435 and n7641_not n7643 ; n8871
g6436 and n8870_not n8871 ; n8872
g6437 and pi1161 pi1163_not ; n8873
g6438 and n2926 n8873 ; n8874
g6439 and pi0031_not pi1162 ; n8875
g6440 and n8874 n8875 ; n8876
g6441 or n8872 n8876 ; po0189
g6442 and n2529 n3328 ; n8878
g6443 nor pi0055 pi0074 ; n8879
g6444 and n8878 n8879 ; n8880
g6445 and n6134 n8880 ; n8881
g6446 and pi0100 n2530 ; n8882
g6447 nor n6263 po1057 ; n8883
g6448 and n6351 n8883 ; n8884
g6449 and pi0137_not n8884 ; n8885
g6450 and pi0137_not pi0252 ; n8886
g6451 and pi0129 n2521 ; n8887
g6452 and po1057 n7474_not ; n8888
g6453 and n6263 n8888_not ; n8889
g6454 and n8886 n8889 ; n8890
g6455 and n8887 n8890 ; n8891
g6456 nor n8885 n8891 ; n8892
g6457 and n8882 n8892_not ; n8893
g6458 nor pi0024 pi0090 ; n8894
g6459 and n6171 n8894 ; n8895
g6460 and n2497 n2714 ; n8896
g6461 and n2701 n8896 ; n8897
g6462 and pi0050 n2777 ; n8898
g6463 and n2495 n8898 ; n8899
g6464 and pi0093_not n8897 ; n8900
g6465 and n8899 n8900 ; n8901
g6466 and n8895 n8901 ; n8902
g6467 and pi0829 pi1093_not ; n8903
g6468 and n2932 n8903 ; n8904
g6469 or n2928 n8904 ; po0840
g6470 nor n7425 po0840 ; n8906
g6471 nor pi0137 n8906 ; n8907
g6472 and n8902 n8907_not ; n8908
g6473 nor pi0068 pi0073 ; n8909
g6474 and n2462 n2804 ; n8910
g6475 and pi0103_not n2471 ; n8911
g6476 and n8910 n8911 ; n8912
g6477 nor pi0089 pi0102 ; n8913
g6478 and n7438 n8913 ; n8914
g6479 nor pi0045 pi0048 ; n8915
g6480 and n2466 n2797 ; n8916
g6481 nor pi0061 pi0104 ; n8917
g6482 and n8915 n8917 ; n8918
g6483 and n8916 n8918 ; n8919
g6484 nor pi0049 pi0066 ; n8920
g6485 nor pi0064 pi0081 ; n8921
g6486 and n2487 n8921 ; n8922
g6487 and pi0076 pi0084_not ; n8923
g6488 and n2479 n8923 ; n8924
g6489 and n8909 n8920 ; n8925
g6490 and n8924 n8925 ; n8926
g6491 and n8914 n8922 ; n8927
g6492 and n8926 n8927 ; n8928
g6493 and n8912 n8919 ; n8929
g6494 and n8928 n8929 ; n8930
g6495 and n2495 n8930 ; n8931
g6496 and n8897 n8931 ; n8932
g6497 and pi0024 n8932_not ; n8933
g6498 nor n8898 n8930 ; n8934
g6499 and n2499 n2702 ; n8935
g6500 and n8934_not n8935 ; n8936
g6501 nor pi0024 n8936 ; n8937
g6502 and n2507 n2736 ; n8938
g6503 and pi0137_not n7445 ; n8939
g6504 and n8938 n8939 ; n8940
g6505 and n8906_not n8940 ; n8941
g6506 and n8933_not n8941 ; n8942
g6507 and n8937_not n8942 ; n8943
g6508 nor n8908 n8943 ; n8944
g6509 nor pi0032 n8944 ; n8945
g6510 nor pi0024 pi0841 ; n8946
g6511 and pi0032 n8946_not ; n8947
g6512 and n2710 n8947 ; n8948
g6513 nor n8945 n8948 ; n8949
g6514 nor n6169 n8949 ; n8950
g6515 nor pi0032 n8902 ; n8951
g6516 and n6169 n6173_not ; n8952
g6517 and n8951_not n8952 ; n8953
g6518 nor n8950 n8953 ; n8954
g6519 and pi0095_not n2531 ; n8955
g6520 and n8954_not n8955 ; n8956
g6521 nor n8893 n8956 ; n8957
g6522 and n2533 n8957_not ; n8958
g6523 and pi0024_not n2505 ; n8959
g6524 and n2519 n2705 ; n8960
g6525 and pi0051_not n8960 ; n8961
g6526 and n8959 n8961 ; n8962
g6527 and po0840_not n8962 ; n8963
g6528 and pi0252 n8888_not ; n8964
g6529 and pi0087_not n2530 ; n8965
g6530 and pi0075 pi0100_not ; n8966
g6531 and n8965 n8966 ; n8967
g6532 and pi0137_not n8967 ; n8968
g6533 and n6282_not n8968 ; n8969
g6534 and n8964_not n8969 ; n8970
g6535 and n8963 n8970 ; n8971
g6536 nor n8958 n8971 ; n8972
g6537 and n8881 n8972_not ; po0190
g6538 nor pi0195 pi0196 ; n8974
g6539 and pi0138_not n8974 ; n8975
g6540 and pi0139_not n8975 ; n8976
g6541 and pi0118_not n8976 ; n8977
g6542 and pi0079_not n8977 ; n8978
g6543 and pi0034_not n8978 ; n8979
g6544 nor pi0033 n8979 ; n8980
g6545 and pi0149 pi0157 ; n8981
g6546 nor pi0149 pi0157 ; n8982
g6547 and n6197 n8982_not ; n8983
g6548 and n8981_not n8983 ; n8984
g6549 and pi0232 n8984 ; n8985
g6550 and pi0075 n8985_not ; n8986
g6551 and pi0100 n8985_not ; n8987
g6552 nor n8986 n8987 ; n8988
g6553 nor pi0075 pi0100 ; n8989
g6554 and n7473 n8989 ; n8990
g6555 and pi0164 n8990 ; n8991
g6556 and n8988 n8991_not ; n8992
g6557 nor pi0074 n8992 ; n8993
g6558 and pi0169 n8990 ; n8994
g6559 and n8988 n8994_not ; n8995
g6560 and pi0074 n8995_not ; n8996
g6561 nor n3328 n8993 ; n8997
g6562 and n8996_not n8997 ; n8998
g6563 and pi0054 n8992_not ; n8999
g6564 and pi0164 n7473 ; n9000
g6565 and pi0038 n9000 ; n9001
g6566 and n8989 n9001 ; n9002
g6567 and n8988 n9002_not ; n9003
g6568 and n8999_not n9003 ; n9004
g6569 nor pi0074 n9004 ; n9005
g6570 nor n8996 n9005 ; n9006
g6571 nor n2529 n9006 ; n9007
g6572 and n3328 n9007_not ; n9008
g6573 and pi0299 n8984_not ; n9009
g6574 and pi0178 pi0183 ; n9010
g6575 nor pi0178 pi0183 ; n9011
g6576 and n6197 n9011_not ; n9012
g6577 and n9010_not n9012 ; n9013
g6578 nor pi0299 n9013 ; n9014
g6579 and pi0232 n9009_not ; n9015
g6580 and n9014_not n9015 ; n9016
g6581 and pi0100 n9016_not ; n9017
g6582 and pi0075 n9016_not ; n9018
g6583 nor n9017 n9018 ; n9019
g6584 and pi0191 pi0299_not ; n9020
g6585 and pi0169 pi0299 ; n9021
g6586 nor n9020 n9021 ; n9022
g6587 and n8990 n9022_not ; n9023
g6588 and n9019 n9023_not ; n9024
g6589 and pi0074 n9024_not ; n9025
g6590 nor pi0055 n9025 ; n9026
g6591 nor pi0186 pi0299 ; n9027
g6592 and pi0164_not pi0299 ; n9028
g6593 nor n9027 n9028 ; n9029
g6594 and n7473 n9029 ; n9030
g6595 and n8989 n9030 ; n9031
g6596 and n9019 n9031_not ; n9032
g6597 and pi0054 n9032_not ; n9033
g6598 and pi0038 n9030 ; n9034
g6599 and pi0087 n9034_not ; n9035
g6600 and pi0216 n6379 ; n9036
g6601 and n6243 n6392_not ; n9037
g6602 and pi0154 n9037_not ; n9038
g6603 and n6243 n6396 ; n9039
g6604 nor pi0154 n9039 ; n9040
g6605 nor pi0152 n9040 ; n9041
g6606 and n9038_not n9041 ; n9042
g6607 and n6197 n7602 ; n9043
g6608 and n6242_not n9043 ; n9044
g6609 and pi0152 pi0154 ; n9045
g6610 and n9044 n9045 ; n9046
g6611 nor n9042 n9046 ; n9047
g6612 and n9036 n9047_not ; n9048
g6613 and pi0299 n9048_not ; n9049
g6614 and pi0176_not pi0232 ; n9050
g6615 and pi0224 n6405 ; n9051
g6616 and n6206 n6396 ; n9052
g6617 and n9051 n9052 ; n9053
g6618 and pi0174_not n9053 ; n9054
g6619 nor pi0299 n9054 ; n9055
g6620 and n9050 n9055_not ; n9056
g6621 and pi0176 pi0232 ; n9057
g6622 and n6206 n9051 ; n9058
g6623 and n7602 n9058 ; n9059
g6624 and pi0174 n9059 ; n9060
g6625 and n6392_not n9051 ; n9061
g6626 and n6206 n9061 ; n9062
g6627 and pi0174_not n9062 ; n9063
g6628 nor pi0299 n9060 ; n9064
g6629 and n9063_not n9064 ; n9065
g6630 and n9057 n9065_not ; n9066
g6631 nor n9056 n9066 ; n9067
g6632 and pi0039 n9049_not ; n9068
g6633 and n9067_not n9068 ; n9069
g6634 and n3181 n6197 ; n9070
g6635 and pi0180 n9070 ; n9071
g6636 and pi0090 n7432_not ; n9072
g6637 nor pi0072 pi0093 ; n9073
g6638 and n2707 n9073 ; n9074
g6639 and n9072_not n9074 ; n9075
g6640 nor pi0066 pi0084 ; n9076
g6641 and pi0068_not n2468 ; n9077
g6642 and pi0111_not n2467 ; n9078
g6643 and pi0036_not n9077 ; n9079
g6644 and n9078 n9079 ; n9080
g6645 and pi0102_not n8921 ; n9081
g6646 and n2466 n9081 ; n9082
g6647 and n2464 n9082 ; n9083
g6648 and pi0073 pi0082_not ; n9084
g6649 and n9076 n9084 ; n9085
g6650 and n9080 n9085 ; n9086
g6651 and n9083 n9086 ; n9087
g6652 and n2477 n9087 ; n9088
g6653 and n8935 n9088 ; n9089
g6654 and n2487 n9089 ; n9090
g6655 and n6139 n9090_not ; n9091
g6656 and n9075 n9091_not ; n9092
g6657 and n2518 n6197 ; n9093
g6658 and pi0040_not n9093 ; n9094
g6659 and n9092 n9094 ; n9095
g6660 and pi0183_not n9095 ; n9096
g6661 and pi0183 n6197 ; n9097
g6662 and n2504 n6139_not ; n9098
g6663 and n9072_not n9098 ; n9099
g6664 and n2485 n9083 ; n9100
g6665 and pi0060_not n9100 ; n9101
g6666 and pi0053 n9101_not ; n9102
g6667 and pi0060_not n8898 ; n9103
g6668 and n2719 n9103_not ; n9104
g6669 nor n9102 n9104 ; n9105
g6670 and n2494 n9088 ; n9106
g6671 and n2487 n9106_not ; n9107
g6672 and n9105_not n9107 ; n9108
g6673 and n2720 n9108_not ; n9109
g6674 and pi0090_not n2717 ; n9110
g6675 and n2504 n9110 ; n9111
g6676 and n2723 n9111 ; n9112
g6677 and n2487 n9112 ; n9113
g6678 and n9109 n9113 ; n9114
g6679 nor pi0070 n9114 ; n9115
g6680 and n9099_not n9115 ; n9116
g6681 and n2519 n3100 ; n9117
g6682 and n9116_not n9117 ; n9118
g6683 and n9115_not n9117 ; n9119
g6684 nor n6487 n9119 ; n9120
g6685 nor pi0198 n9120 ; n9121
g6686 nor n9118 n9121 ; n9122
g6687 and n9097 n9122_not ; n9123
g6688 nor pi0174 n9096 ; n9124
g6689 and n9123_not n9124 ; n9125
g6690 and n9104_not n9112 ; n9126
g6691 nor pi0070 n9126 ; n9127
g6692 and n9099_not n9127 ; n9128
g6693 and n9117 n9128_not ; n9129
g6694 nor n6519 n9129 ; n9130
g6695 and n6197 n9130_not ; n9131
g6696 and pi0183 n9131 ; n9132
g6697 and n6139_not n9075 ; n9133
g6698 and n9094 n9133 ; n9134
g6699 and pi0183_not n9134 ; n9135
g6700 and pi0174 n9135_not ; n9136
g6701 and n9132_not n9136 ; n9137
g6702 nor n9125 n9137 ; n9138
g6703 and pi0193 n9138_not ; n9139
g6704 and pi0040_not n6197 ; n9140
g6705 and pi0090_not n9074 ; n9141
g6706 and n9090 n9141 ; n9142
g6707 and n2518 n9142 ; n9143
g6708 and n9140 n9143 ; n9144
g6709 nor pi0174 pi0183 ; n9145
g6710 and n9144 n9145 ; n9146
g6711 nor n6519 n9119 ; n9147
g6712 and pi0174_not n9147 ; n9148
g6713 and n9117 n9127_not ; n9149
g6714 nor n6519 n9149 ; n9150
g6715 and pi0174 n9150 ; n9151
g6716 and n9097 n9151_not ; n9152
g6717 and n9148_not n9152 ; n9153
g6718 nor pi0193 n9146 ; n9154
g6719 and n9153_not n9154 ; n9155
g6720 nor n9139 n9155 ; n9156
g6721 nor pi0299 n9071 ; n9157
g6722 and n9156_not n9157 ; n9158
g6723 and pi0039_not pi0232 ; n9159
g6724 and pi0158 n9070 ; n9160
g6725 and pi0172 n9118 ; n9161
g6726 nor n6488 n9119 ; n9162
g6727 and pi0152_not n9162 ; n9163
g6728 and n9161_not n9163 ; n9164
g6729 and pi0172 n9129 ; n9165
g6730 nor n6488 n9149 ; n9166
g6731 and pi0152 n9165_not ; n9167
g6732 and n9166 n9167 ; n9168
g6733 and pi0149 n6197 ; n9169
g6734 and n9168_not n9169 ; n9170
g6735 and n9164_not n9170 ; n9171
g6736 and pi0152_not n9095 ; n9172
g6737 nor n9134 n9172 ; n9173
g6738 and pi0172 n9173_not ; n9174
g6739 nor pi0152 pi0172 ; n9175
g6740 and n9144 n9175 ; n9176
g6741 nor n9174 n9176 ; n9177
g6742 nor pi0149 n9177 ; n9178
g6743 and pi0299 n9160_not ; n9179
g6744 and n9178_not n9179 ; n9180
g6745 and n9171_not n9180 ; n9181
g6746 and n9159 n9181_not ; n9182
g6747 and n9158_not n9182 ; n9183
g6748 nor n9069 n9183 ; n9184
g6749 nor pi0038 n9184 ; n9185
g6750 and pi0299 n7473 ; n9186
g6751 and n6135_not n9186 ; n9187
g6752 nor pi0186 n9187 ; n9188
g6753 and n6284_not n7473 ; n9189
g6754 and pi0186 n9189_not ; n9190
g6755 and pi0164 n9190_not ; n9191
g6756 and n9188_not n9191 ; n9192
g6757 and pi0299_not n7473 ; n9193
g6758 and n6135_not n9193 ; n9194
g6759 and pi0164_not pi0186 ; n9195
g6760 and n9194 n9195 ; n9196
g6761 nor n9192 n9196 ; n9197
g6762 and pi0038 n9197_not ; n9198
g6763 nor pi0087 n9198 ; n9199
g6764 and n9185_not n9199 ; n9200
g6765 nor pi0100 n9035 ; n9201
g6766 and n9200_not n9201 ; n9202
g6767 nor n9017 n9202 ; n9203
g6768 and n2569 n9203_not ; n9204
g6769 and pi0075_not pi0092 ; n9205
g6770 and pi0100_not n9034 ; n9206
g6771 nor n9017 n9206 ; n9207
g6772 nor pi0038 pi0087 ; n9208
g6773 and pi0232 n3383_not ; n9209
g6774 nor pi0176 pi0299 ; n9210
g6775 and n6197 n9210_not ; n9211
g6776 and n9209 n9211 ; n9212
g6777 and pi0100_not n9208 ; n9213
g6778 and n9212 n9213 ; n9214
g6779 and n6135 n9214 ; n9215
g6780 and n9207 n9215_not ; n9216
g6781 and n9205 n9216_not ; n9217
g6782 nor n9018 n9217 ; n9218
g6783 and n9204_not n9218 ; n9219
g6784 nor pi0054 n9219 ; n9220
g6785 nor n9033 n9220 ; n9221
g6786 nor pi0074 n9221 ; n9222
g6787 and n9026 n9222_not ; n9223
g6788 and pi0055 n8996_not ; n9224
g6789 nor pi0092 n8986 ; n9225
g6790 and pi0038 n9000_not ; n9226
g6791 and n2568 n9226_not ; n9227
g6792 and pi0149 n7473 ; n9228
g6793 and n6135 n9228 ; n9229
g6794 nor pi0038 n9229 ; n9230
g6795 and n9227 n9230_not ; n9231
g6796 and n8161 n9001 ; n9232
g6797 nor n8987 n9232 ; n9233
g6798 and n9231_not n9233 ; n9234
g6799 nor pi0075 n9234 ; n9235
g6800 and n9225 n9235_not ; n9236
g6801 and pi0092 n9003 ; n9237
g6802 nor pi0054 n9237 ; n9238
g6803 and n9236_not n9238 ; n9239
g6804 nor n8999 n9239 ; n9240
g6805 nor pi0074 n9240 ; n9241
g6806 and n9224 n9241_not ; n9242
g6807 and n2529 n9242_not ; n9243
g6808 and n9223_not n9243 ; n9244
g6809 and n9008 n9244_not ; n9245
g6810 nor n8998 n9245 ; n9246
g6811 and n8980 n9246_not ; n9247
g6812 and pi0040_not n2487 ; n9248
g6813 and pi0038_not n9248 ; n9249
g6814 and n8989 n9249 ; n9250
g6815 and n2532 n9250 ; n9251
g6816 and n2529_not n9251 ; n9252
g6817 and n2716 n2720 ; n9253
g6818 and pi0053_not n9253 ; n9254
g6819 and n9101 n9254 ; n9255
g6820 and pi0058_not n9255 ; n9256
g6821 and n7445 n9256 ; n9257
g6822 and pi0032_not n2508 ; n9258
g6823 and n9257 n9258 ; n9259
g6824 and pi0095_not n9259 ; n9260
g6825 nor pi0039 n9228 ; n9261
g6826 and n9260 n9261 ; n9262
g6827 and n9248 n9262_not ; n9263
g6828 nor pi0038 n9263 ; n9264
g6829 and n9227 n9264_not ; n9265
g6830 nor pi0038 n9248 ; n9266
g6831 nor pi0100 n9266 ; n9267
g6832 and n9226_not n9267 ; n9268
g6833 and pi0087 n9268 ; n9269
g6834 nor n8987 n9269 ; n9270
g6835 and n9265_not n9270 ; n9271
g6836 nor pi0075 n9271 ; n9272
g6837 and n9225 n9272_not ; n9273
g6838 and pi0075_not n9268 ; n9274
g6839 and pi0092 n8988 ; n9275
g6840 and n9274_not n9275 ; n9276
g6841 nor pi0054 n9276 ; n9277
g6842 and n9273_not n9277 ; n9278
g6843 nor n8999 n9278 ; n9279
g6844 nor pi0074 n9279 ; n9280
g6845 and n9224 n9280_not ; n9281
g6846 and n2609 n9260 ; n9282
g6847 and n9212_not n9282 ; n9283
g6848 and n2608 n9248 ; n9284
g6849 and n9283_not n9284 ; n9285
g6850 and n9207 n9285_not ; n9286
g6851 and n9205 n9286_not ; n9287
g6852 and pi0087 n9284_not ; n9288
g6853 and n9207 n9288 ; n9289
g6854 and n9036_not n9248 ; n9290
g6855 and pi0299 n9290_not ; n9291
g6856 and n6383 n6395_not ; n9292
g6857 and n6212 n9292 ; n9293
g6858 nor n6188 n9293 ; n9294
g6859 and n9260 n9294_not ; n9295
g6860 and n6198 n9295 ; n9296
g6861 and n9248 n9296_not ; n9297
g6862 and n6197 n9295 ; n9298
g6863 and n9248 n9298_not ; n9299
g6864 nor n6242 n9299 ; n9300
g6865 and n9297 n9300_not ; n9301
g6866 and n9291 n9301_not ; n9302
g6867 and n9051_not n9248 ; n9303
g6868 nor n9297 n9303 ; n9304
g6869 nor n6205 n9299 ; n9305
g6870 and n9303_not n9305 ; n9306
g6871 nor n9304 n9306 ; n9307
g6872 nor pi0299 n9307 ; n9308
g6873 nor n9302 n9308 ; n9309
g6874 nor pi0232 n9309 ; n9310
g6875 and n9260 n9293 ; n9311
g6876 and n6197 n9311 ; n9312
g6877 and n9248 n9312_not ; n9313
g6878 nor n6205 n9313 ; n9314
g6879 and n9303_not n9314 ; n9315
g6880 and pi0174 n9315 ; n9316
g6881 nor n9304 n9316 ; n9317
g6882 nor pi0299 n9317 ; n9318
g6883 and n9248 n9311_not ; n9319
g6884 and n6243 n9319_not ; n9320
g6885 and pi0152 n9320 ; n9321
g6886 and n9297 n9321_not ; n9322
g6887 and pi0154 n9322_not ; n9323
g6888 and n6188 n9260 ; n9324
g6889 and n6227_not n9324 ; n9325
g6890 and n9248 n9325_not ; n9326
g6891 and n6197 n9326 ; n9327
g6892 and pi0152_not n9327 ; n9328
g6893 nor pi0154 n9301 ; n9329
g6894 and n9328_not n9329 ; n9330
g6895 and n9036 n9323_not ; n9331
g6896 and n9330_not n9331 ; n9332
g6897 and n9291 n9332_not ; n9333
g6898 nor n9318 n9333 ; n9334
g6899 and n6206 n9324 ; n9335
g6900 and n9051 n9248 ; n9336
g6901 and n9335_not n9336 ; n9337
g6902 nor n9303 n9337 ; n9338
g6903 and pi0299_not n9338 ; n9339
g6904 and n9334 n9339_not ; n9340
g6905 and n9050 n9340_not ; n9341
g6906 and n9057 n9334_not ; n9342
g6907 and pi0039 n9310_not ; n9343
g6908 and n9342_not n9343 ; n9344
g6909 and n9341_not n9344 ; n9345
g6910 and pi0095 n9248_not ; n9346
g6911 nor n2442 n9346 ; n9347
g6912 nor pi0040 pi0479 ; n9348
g6913 and n2487 n9259_not ; n9349
g6914 and n9348 n9349 ; n9350
g6915 nor n9347 n9350 ; n9351
g6916 and pi0032 n9248_not ; n9352
g6917 and n2487 n2506_not ; n9353
g6918 and n2487 n9257_not ; n9354
g6919 and pi0070 n9354_not ; n9355
g6920 and n2487 n9255_not ; n9356
g6921 and pi0058 n9356_not ; n9357
g6922 and n2487 n2716_not ; n9358
g6923 nor n2487 n2720 ; n9359
g6924 and n2716 n9359_not ; n9360
g6925 and n9109_not n9360 ; n9361
g6926 nor pi0058 n9358 ; n9362
g6927 and n9361_not n9362 ; n9363
g6928 nor n9357 n9363 ; n9364
g6929 nor pi0090 n9364 ; n9365
g6930 and pi0841_not n9256 ; n9366
g6931 and n2487 n9366_not ; n9367
g6932 and pi0090 n9367_not ; n9368
g6933 and n2504 n9368_not ; n9369
g6934 and n9365_not n9369 ; n9370
g6935 and n2487 n2504_not ; n9371
g6936 nor pi0070 n9371 ; n9372
g6937 and n9370_not n9372 ; n9373
g6938 nor n9355 n9373 ; n9374
g6939 nor pi0051 n9374 ; n9375
g6940 and pi0051 n2487_not ; n9376
g6941 and n2506 n9376_not ; n9377
g6942 and n9375_not n9377 ; n9378
g6943 nor n9353 n9378 ; n9379
g6944 nor pi0040 n9379 ; n9380
g6945 nor pi0032 n9380 ; n9381
g6946 nor n9352 n9381 ; n9382
g6947 nor pi0095 n9382 ; n9383
g6948 nor n9351 n9383 ; n9384
g6949 and n9141 n9366 ; n9385
g6950 and n9248 n9385_not ; n9386
g6951 and pi0032 n9386_not ; n9387
g6952 nor n9381 n9387 ; n9388
g6953 nor pi0095 n9388 ; n9389
g6954 and pi0198_not n9389 ; n9390
g6955 and n9384 n9390_not ; n9391
g6956 and n6197_not n9391 ; n9392
g6957 and n9105 n9253 ; n9393
g6958 and n2487 n9393_not ; n9394
g6959 nor pi0058 n9394 ; n9395
g6960 nor n9357 n9395 ; n9396
g6961 nor pi0090 n9396 ; n9397
g6962 and n9369 n9397_not ; n9398
g6963 and n9372 n9398_not ; n9399
g6964 nor n9355 n9399 ; n9400
g6965 nor pi0051 n9400 ; n9401
g6966 and n9377 n9401_not ; n9402
g6967 nor n9353 n9402 ; n9403
g6968 nor pi0040 n9403 ; n9404
g6969 nor pi0032 n9404 ; n9405
g6970 nor n9387 n9405 ; n9406
g6971 nor pi0095 n9406 ; n9407
g6972 and pi0198_not n9407 ; n9408
g6973 and n6197 n9346_not ; n9409
g6974 nor n9352 n9405 ; n9410
g6975 nor pi0095 n9410 ; n9411
g6976 and n9409 n9411_not ; n9412
g6977 and n9408_not n9412 ; n9413
g6978 nor n9392 n9413 ; n9414
g6979 nor pi0183 n9414 ; n9415
g6980 nor pi0040 n9352 ; n9416
g6981 and n2487 n6170_not ; n9417
g6982 nor pi0032 n9417 ; n9418
g6983 and pi0093 n2487_not ; n9419
g6984 and n6170 n9419_not ; n9420
g6985 and n2487 n9357_not ; n9421
g6986 nor pi0090 n9421 ; n9422
g6987 nor n9368 n9422 ; n9423
g6988 nor pi0093 n9423 ; n9424
g6989 and n9420 n9424_not ; n9425
g6990 and n9418 n9425_not ; n9426
g6991 and n9416 n9426_not ; n9427
g6992 nor pi0095 n9427 ; n9428
g6993 and n9409 n9428_not ; n9429
g6994 nor n9392 n9429 ; n9430
g6995 and pi0183 n9430_not ; n9431
g6996 nor n9415 n9431 ; n9432
g6997 and pi0095_not n9432 ; n9433
g6998 nor pi0174 n9351 ; n9434
g6999 and n9433_not n9434 ; n9435
g7000 nor n9097 n9391 ; n9436
g7001 and pi0090_not n9089 ; n9437
g7002 and n9423 n9437_not ; n9438
g7003 nor pi0093 n9438 ; n9439
g7004 and n9420 n9439_not ; n9440
g7005 and n9418 n9440_not ; n9441
g7006 and n9416 n9441_not ; n9442
g7007 nor pi0095 n9442 ; n9443
g7008 nor n9351 n9443 ; n9444
g7009 and n6197 n9444_not ; n9445
g7010 and pi0183 n9445 ; n9446
g7011 and pi0174 n9446_not ; n9447
g7012 and n9436_not n9447 ; n9448
g7013 nor pi0180 n9448 ; n9449
g7014 and n9435_not n9449 ; n9450
g7015 nor pi0174 n9432 ; n9451
g7016 and n9409 n9443_not ; n9452
g7017 nor n9392 n9452 ; n9453
g7018 and pi0183 n9453_not ; n9454
g7019 nor n9346 n9383 ; n9455
g7020 and n9390_not n9455 ; n9456
g7021 and n9140 n9456 ; n9457
g7022 nor n9392 n9457 ; n9458
g7023 nor pi0183 n9458 ; n9459
g7024 nor n9454 n9459 ; n9460
g7025 and pi0174 n9460_not ; n9461
g7026 and pi0180 n9451_not ; n9462
g7027 and n9461_not n9462 ; n9463
g7028 nor n9450 n9463 ; n9464
g7029 nor pi0193 n9464 ; n9465
g7030 nor pi0040 n2487 ; n9466
g7031 and pi0032 n9466_not ; n9467
g7032 and n2461 n2504 ; n9468
g7033 nor n2487 n9468 ; n9469
g7034 and n7445 n9363 ; n9470
g7035 nor n9469 n9470 ; n9471
g7036 nor pi0070 n9471 ; n9472
g7037 nor n9355 n9472 ; n9473
g7038 nor pi0051 n9473 ; n9474
g7039 and n9377 n9474_not ; n9475
g7040 nor pi0040 n9353 ; n9476
g7041 and n9475_not n9476 ; n9477
g7042 nor pi0032 n9477 ; n9478
g7043 nor n9467 n9478 ; n9479
g7044 nor n2736 n9248 ; n9480
g7045 nor n9479 n9480 ; n9481
g7046 nor pi0095 n9481 ; n9482
g7047 nor n9351 n9482 ; n9483
g7048 nor n9346 n9482 ; n9484
g7049 and pi0095 n9466_not ; n9485
g7050 nor pi0040 n9386 ; n9486
g7051 and pi0032 n9486_not ; n9487
g7052 nor n9478 n9487 ; n9488
g7053 nor pi0095 n9488 ; n9489
g7054 nor n9485 n9489 ; n9490
g7055 and n9484 n9490_not ; n9491
g7056 nor pi0198 n9491 ; n9492
g7057 and n6197 n9492_not ; n9493
g7058 and n6197 n9248_not ; n9494
g7059 nor n9493 n9494 ; n9495
g7060 and n9483 n9495_not ; n9496
g7061 nor n9392 n9496 ; n9497
g7062 nor pi0183 n9497 ; n9498
g7063 and n2704 n6170 ; n9499
g7064 and n8935 n9499 ; n9500
g7065 and pi0032_not n9500 ; n9501
g7066 and n9088 n9501 ; n9502
g7067 and n9248 n9502_not ; n9503
g7068 nor pi0095 n9503 ; n9504
g7069 and n6197 n9504_not ; n9505
g7070 and n9351_not n9505 ; n9506
g7071 nor n9392 n9506 ; n9507
g7072 and pi0183 n9507_not ; n9508
g7073 and pi0174 n9508_not ; n9509
g7074 and n9498_not n9509 ; n9510
g7075 nor n6197 n9391 ; n9511
g7076 and n7445 n9395 ; n9512
g7077 nor n9469 n9512 ; n9513
g7078 nor pi0070 n9513 ; n9514
g7079 nor n9355 n9514 ; n9515
g7080 nor pi0051 n9515 ; n9516
g7081 and n9377 n9516_not ; n9517
g7082 nor n9353 n9517 ; n9518
g7083 nor pi0040 n9518 ; n9519
g7084 nor pi0032 n9519 ; n9520
g7085 nor n9352 n9520 ; n9521
g7086 nor pi0095 n9521 ; n9522
g7087 nor n9351 n9522 ; n9523
g7088 nor n9387 n9520 ; n9524
g7089 nor pi0095 n9524 ; n9525
g7090 and pi0198_not n9525 ; n9526
g7091 and n9523 n9526_not ; n9527
g7092 and n6197 n9527_not ; n9528
g7093 nor n9511 n9528 ; n9529
g7094 and pi0183_not n9529 ; n9530
g7095 nor pi0095 n9248 ; n9531
g7096 nor n9351 n9531 ; n9532
g7097 and n6197 n9532 ; n9533
g7098 nor n9392 n9533 ; n9534
g7099 and pi0183 n9534_not ; n9535
g7100 nor pi0174 n9530 ; n9536
g7101 and n9535_not n9536 ; n9537
g7102 nor pi0180 n9537 ; n9538
g7103 and n9510_not n9538 ; n9539
g7104 and n9409 n9504_not ; n9540
g7105 nor n9392 n9540 ; n9541
g7106 and pi0183 n9541_not ; n9542
g7107 and n9484 n9493 ; n9543
g7108 nor n9392 n9543 ; n9544
g7109 nor pi0183 n9544 ; n9545
g7110 and pi0174 n9542_not ; n9546
g7111 and n9545_not n9546 ; n9547
g7112 nor n9494 n9511 ; n9548
g7113 and pi0183 n9548 ; n9549
g7114 and pi0040_not n9518 ; n9550
g7115 nor pi0032 n9550 ; n9551
g7116 nor n9467 n9551 ; n9552
g7117 nor pi0095 n9552 ; n9553
g7118 nor n9485 n9553 ; n9554
g7119 and pi0198 n9554_not ; n9555
g7120 nor n9487 n9551 ; n9556
g7121 nor pi0095 n9556 ; n9557
g7122 nor n9485 n9557 ; n9558
g7123 nor pi0198 n9558 ; n9559
g7124 nor n9555 n9559 ; n9560
g7125 and n9140 n9560_not ; n9561
g7126 nor n9392 n9561 ; n9562
g7127 nor pi0183 n9562 ; n9563
g7128 nor pi0174 n9549 ; n9564
g7129 and n9563_not n9564 ; n9565
g7130 and pi0180 n9547_not ; n9566
g7131 and n9565_not n9566 ; n9567
g7132 and pi0193 n9539_not ; n9568
g7133 and n9567_not n9568 ; n9569
g7134 nor n9465 n9569 ; n9570
g7135 nor pi0299 n9570 ; n9571
g7136 and pi0158 pi0299 ; n9572
g7137 and pi0210_not n9389 ; n9573
g7138 and n9384 n9573_not ; n9574
g7139 and n6197_not n9574 ; n9575
g7140 and pi0210_not n9407 ; n9576
g7141 and n9412 n9576_not ; n9577
g7142 nor n9575 n9577 ; n9578
g7143 nor pi0152 n9578 ; n9579
g7144 nor n6197 n9574 ; n9580
g7145 and n9455 n9573_not ; n9581
g7146 and n6197 n9581_not ; n9582
g7147 nor n9580 n9582 ; n9583
g7148 and pi0152 n9583 ; n9584
g7149 nor pi0172 n9579 ; n9585
g7150 and n9584_not n9585 ; n9586
g7151 nor n9346 n9525 ; n9587
g7152 nor pi0210 n9587 ; n9588
g7153 and n6197 n9588_not ; n9589
g7154 nor n9346 n9522 ; n9590
g7155 and n9589 n9590 ; n9591
g7156 nor n9575 n9591 ; n9592
g7157 nor pi0152 n9592 ; n9593
g7158 nor pi0210 n9491 ; n9594
g7159 and n6197 n9594_not ; n9595
g7160 and n9484 n9595 ; n9596
g7161 nor n9575 n9596 ; n9597
g7162 and pi0152 n9597_not ; n9598
g7163 and pi0172 n9593_not ; n9599
g7164 and n9598_not n9599 ; n9600
g7165 nor n9586 n9600 ; n9601
g7166 and n9572 n9601_not ; n9602
g7167 and pi0158_not pi0299 ; n9603
g7168 nor n9351 n9411 ; n9604
g7169 and n9576_not n9604 ; n9605
g7170 and n6197 n9605 ; n9606
g7171 nor pi0152 n9606 ; n9607
g7172 and pi0152 n9574_not ; n9608
g7173 nor pi0172 n9607 ; n9609
g7174 and n9608_not n9609 ; n9610
g7175 nor n9494 n9595 ; n9611
g7176 and n9483 n9611_not ; n9612
g7177 and pi0152 n9612_not ; n9613
g7178 nor n9494 n9589 ; n9614
g7179 and n9523 n9614_not ; n9615
g7180 nor pi0152 n9615 ; n9616
g7181 and pi0172 n9616_not ; n9617
g7182 and n9613_not n9617 ; n9618
g7183 and n9575_not n9603 ; n9619
g7184 and n9610_not n9619 ; n9620
g7185 and n9618_not n9620 ; n9621
g7186 nor pi0149 n9621 ; n9622
g7187 and n9602_not n9622 ; n9623
g7188 nor n9452 n9575 ; n9624
g7189 and pi0152 n9624_not ; n9625
g7190 nor n9429 n9575 ; n9626
g7191 nor pi0152 n9626 ; n9627
g7192 nor pi0172 n9625 ; n9628
g7193 and n9627_not n9628 ; n9629
g7194 nor n9540 n9575 ; n9630
g7195 and pi0152 n9630_not ; n9631
g7196 nor n9494 n9580 ; n9632
g7197 and pi0152_not n9632 ; n9633
g7198 and pi0172 n9631_not ; n9634
g7199 and n9633_not n9634 ; n9635
g7200 nor n9629 n9635 ; n9636
g7201 and n9572 n9636_not ; n9637
g7202 nor n9506 n9575 ; n9638
g7203 and pi0152 n9638_not ; n9639
g7204 nor n9533 n9575 ; n9640
g7205 nor pi0152 n9640 ; n9641
g7206 and pi0172 n9639_not ; n9642
g7207 and n9641_not n9642 ; n9643
g7208 nor n9351 n9428 ; n9644
g7209 and n6197 n9644_not ; n9645
g7210 nor n9580 n9645 ; n9646
g7211 and pi0152_not n9646 ; n9647
g7212 nor n9445 n9580 ; n9648
g7213 and pi0152 n9648 ; n9649
g7214 nor pi0172 n9647 ; n9650
g7215 and n9649_not n9650 ; n9651
g7216 nor n9643 n9651 ; n9652
g7217 and n9603 n9652_not ; n9653
g7218 and pi0149 n9637_not ; n9654
g7219 and n9653_not n9654 ; n9655
g7220 nor n9623 n9655 ; n9656
g7221 nor n9571 n9656 ; n9657
g7222 and pi0232 n9657_not ; n9658
g7223 and n6169_not n9389 ; n9659
g7224 and n9384 n9659_not ; n9660
g7225 nor pi0232 n9660 ; n9661
g7226 nor pi0039 n9661 ; n9662
g7227 and n9658_not n9662 ; n9663
g7228 nor n9345 n9663 ; n9664
g7229 nor pi0038 n9664 ; n9665
g7230 nor n9198 n9665 ; n9666
g7231 nor pi0100 n9666 ; n9667
g7232 nor pi0087 n9017 ; n9668
g7233 and n9667_not n9668 ; n9669
g7234 and n2569 n9289_not ; n9670
g7235 and n9669_not n9670 ; n9671
g7236 nor n9018 n9287 ; n9672
g7237 and n9671_not n9672 ; n9673
g7238 nor pi0054 n9673 ; n9674
g7239 nor n9033 n9674 ; n9675
g7240 nor pi0074 n9675 ; n9676
g7241 and n9026 n9676_not ; n9677
g7242 and n2529 n9281_not ; n9678
g7243 and n9677_not n9678 ; n9679
g7244 and n9008 n9252_not ; n9680
g7245 and n9679_not n9680 ; n9681
g7246 nor n8998 n9681 ; n9682
g7247 nor n8980 n9682 ; n9683
g7248 nor pi0954 n9247 ; n9684
g7249 and n9683_not n9684 ; n9685
g7250 and pi0033 n9246_not ; n9686
g7251 nor pi0033 n9682 ; n9687
g7252 and pi0954 n9686_not ; n9688
g7253 and n9687_not n9688 ; n9689
g7254 nor n9685 n9689 ; po0191
g7255 and pi0197 n8982 ; n9691
g7256 nor pi0197 n8982 ; n9692
g7257 nor n9691 n9692 ; n9693
g7258 and pi0162 n6197 ; n9694
g7259 and n9693 n9694_not ; n9695
g7260 and n9691 n9694 ; n9696
g7261 nor pi0162 pi0197 ; n9697
g7262 and n8983 n9697_not ; n9698
g7263 and n6197 n9698_not ; n9699
g7264 and n9696_not n9699 ; n9700
g7265 nor n9693 n9700 ; n9701
g7266 nor n9695 n9701 ; n9702
g7267 and pi0232 n9702 ; n9703
g7268 and n8989_not n9703 ; n9704
g7269 and pi0167 n7473 ; n9705
g7270 and n8989 n9705 ; n9706
g7271 nor n9704 n9706 ; n9707
g7272 and pi0074_not n9707 ; n9708
g7273 and pi0148 n8990 ; n9709
g7274 and pi0074 n9709_not ; n9710
g7275 and n9704_not n9710 ; n9711
g7276 nor n9708 n9711 ; n9712
g7277 and n3328_not n9712 ; n9713
g7278 nor pi0054 n9704 ; n9714
g7279 and pi0038 n9706 ; n9715
g7280 and n9714 n9715_not ; n9716
g7281 and pi0074_not n9716 ; n9717
g7282 and n9712 n9717_not ; n9718
g7283 nor n2529 n9718 ; n9719
g7284 and n3328 n9719_not ; n9720
g7285 and pi0140 pi0145 ; n9721
g7286 and n9011 n9721_not ; n9722
g7287 nor pi0140 pi0145 ; n9723
g7288 and n6197 n9723_not ; n9724
g7289 and n9722 n9724 ; n9725
g7290 nor n9721 n9723 ; n9726
g7291 and n9012 n9726_not ; n9727
g7292 nor pi0299 n9725 ; n9728
g7293 and n9727_not n9728 ; n9729
g7294 and pi0299 n9702_not ; n9730
g7295 and pi0232 n9729_not ; n9731
g7296 and n9730_not n9731 ; n9732
g7297 and pi0100 n9732_not ; n9733
g7298 and pi0075 n9732_not ; n9734
g7299 nor n9733 n9734 ; n9735
g7300 and pi0141 pi0299_not ; n9736
g7301 and pi0148 pi0299 ; n9737
g7302 nor n9736 n9737 ; n9738
g7303 and n7473 n9738_not ; n9739
g7304 and n8989 n9739_not ; n9740
g7305 and n9735 n9740_not ; n9741
g7306 and pi0074 n9741_not ; n9742
g7307 nor pi0055 n9742 ; n9743
g7308 and pi0188 pi0299_not ; n9744
g7309 and pi0167 pi0299 ; n9745
g7310 nor n9744 n9745 ; n9746
g7311 and n7473 n9746_not ; n9747
g7312 nor pi0100 n9747 ; n9748
g7313 and pi0075_not n9748 ; n9749
g7314 and n9735 n9749_not ; n9750
g7315 and pi0054 n9750_not ; n9751
g7316 nor pi0188 n9187 ; n9752
g7317 and pi0188 n9194 ; n9753
g7318 nor pi0167 n9753 ; n9754
g7319 and pi0167 pi0188 ; n9755
g7320 and n9189_not n9755 ; n9756
g7321 nor n9752 n9756 ; n9757
g7322 and n9754_not n9757 ; n9758
g7323 and pi0038 n9758_not ; n9759
g7324 and pi0038_not pi0155 ; n9760
g7325 and pi0161 n9044_not ; n9761
g7326 nor pi0161 n9037 ; n9762
g7327 and n9036 n9762_not ; n9763
g7328 and n9761_not n9763 ; n9764
g7329 and n9760 n9764_not ; n9765
g7330 nor pi0038 pi0155 ; n9766
g7331 and pi0161_not n9036 ; n9767
g7332 and n9039 n9767 ; n9768
g7333 and n9766 n9768_not ; n9769
g7334 nor n9765 n9769 ; n9770
g7335 and pi0299 n9770_not ; n9771
g7336 nor pi0177 pi0299 ; n9772
g7337 and pi0144_not n9053 ; n9773
g7338 and n9772 n9773_not ; n9774
g7339 and pi0144_not n9062 ; n9775
g7340 and pi0177 pi0299_not ; n9776
g7341 and pi0144 n9059 ; n9777
g7342 and n9776 n9777_not ; n9778
g7343 and n9775_not n9778 ; n9779
g7344 and pi0232 n9774_not ; n9780
g7345 and n9779_not n9780 ; n9781
g7346 nor pi0038 n9781 ; n9782
g7347 nor n9771 n9782 ; n9783
g7348 and pi0039 n9783_not ; n9784
g7349 nor pi0146 n9095 ; n9785
g7350 and pi0146 n9144_not ; n9786
g7351 nor pi0161 n9786 ; n9787
g7352 and n9785_not n9787 ; n9788
g7353 and pi0146_not pi0161 ; n9789
g7354 and n9134 n9789 ; n9790
g7355 nor n9788 n9790 ; n9791
g7356 nor pi0162 n9791 ; n9792
g7357 and pi0159_not pi0299 ; n9793
g7358 and pi0159 pi0299 ; n9794
g7359 and pi0162_not n9070 ; n9795
g7360 and n9794 n9795_not ; n9796
g7361 nor n9793 n9796 ; n9797
g7362 nor n9694 n9797 ; n9798
g7363 and pi0159 n3181 ; n9799
g7364 and pi0146_not n9129 ; n9800
g7365 and n9166 n9800_not ; n9801
g7366 and pi0161 n9801_not ; n9802
g7367 and pi0146_not n9118 ; n9803
g7368 and n9162 n9803_not ; n9804
g7369 nor pi0161 n9804 ; n9805
g7370 and pi0299 n9799_not ; n9806
g7371 and n9802_not n9806 ; n9807
g7372 and n9805_not n9807 ; n9808
g7373 nor n9798 n9808 ; n9809
g7374 nor n9792 n9809 ; n9810
g7375 and pi0181 n9070 ; n9811
g7376 and pi0140 n6197_not ; n9812
g7377 and pi0142_not n9134 ; n9813
g7378 nor pi0140 n9813 ; n9814
g7379 and pi0142_not n9129 ; n9815
g7380 and pi0140 n9815_not ; n9816
g7381 and n9150 n9816 ; n9817
g7382 nor n9814 n9817 ; n9818
g7383 and pi0144 n9818_not ; n9819
g7384 and pi0142_not n9095 ; n9820
g7385 and pi0142 n9144 ; n9821
g7386 nor pi0140 n9821 ; n9822
g7387 and n9820_not n9822 ; n9823
g7388 and pi0142_not n9118 ; n9824
g7389 and pi0140 n9147 ; n9825
g7390 and n9824_not n9825 ; n9826
g7391 nor n9823 n9826 ; n9827
g7392 nor pi0144 n9827 ; n9828
g7393 nor n9812 n9819 ; n9829
g7394 and n9828_not n9829 ; n9830
g7395 nor pi0299 n9811 ; n9831
g7396 and n9830_not n9831 ; n9832
g7397 and pi0232 n9810_not ; n9833
g7398 and n9832_not n9833 ; n9834
g7399 and n2530 n9834_not ; n9835
g7400 nor n9759 n9784 ; n9836
g7401 and n9835_not n9836 ; n9837
g7402 nor pi0100 n9837 ; n9838
g7403 nor n9733 n9838 ; n9839
g7404 nor pi0087 n9839 ; n9840
g7405 nor n2608 n9748 ; n9841
g7406 and n9733_not n9841 ; n9842
g7407 and pi0087 n9842_not ; n9843
g7408 nor n9840 n9843 ; n9844
g7409 and n2569 n9844_not ; n9845
g7410 and pi0038 n9746_not ; n9846
g7411 and pi0155 pi0299 ; n9847
g7412 nor n9776 n9847 ; n9848
g7413 and n2530 n9848_not ; n9849
g7414 and n2512 n9849 ; n9850
g7415 nor n9846 n9850 ; n9851
g7416 and n7473 n9851_not ; n9852
g7417 nor pi0100 n9852 ; n9853
g7418 nor n9733 n9853 ; n9854
g7419 nor pi0087 n9854 ; n9855
g7420 nor n9843 n9855 ; n9856
g7421 and n9205 n9856_not ; n9857
g7422 nor n9734 n9857 ; n9858
g7423 and n9845_not n9858 ; n9859
g7424 nor pi0054 n9859 ; n9860
g7425 nor n9751 n9860 ; n9861
g7426 nor pi0074 n9861 ; n9862
g7427 and n9743 n9862_not ; n9863
g7428 and pi0055 n9711_not ; n9864
g7429 and pi0054 n9707 ; n9865
g7430 and pi0038 n9705 ; n9866
g7431 and pi0092_not pi0162 ; n9867
g7432 and n9159 n9867 ; n9868
g7433 and n9208 n9868 ; n9869
g7434 and n6222 n9869 ; n9870
g7435 nor n9866 n9870 ; n9871
g7436 and n8989 n9871_not ; n9872
g7437 and n9714 n9872_not ; n9873
g7438 nor n9865 n9873 ; n9874
g7439 nor pi0074 n9874 ; n9875
g7440 and n9864 n9875_not ; n9876
g7441 and n2529 n9876_not ; n9877
g7442 and n9863_not n9877 ; n9878
g7443 and n9720 n9878_not ; n9879
g7444 nor n9713 n9879 ; n9880
g7445 and pi0034 n9880 ; n9881
g7446 nor n2529 n9251 ; n9882
g7447 and n3328 n9882_not ; n9883
g7448 nor n9720 n9883 ; n9884
g7449 and n9250_not n9716 ; n9885
g7450 nor n6134 n9885 ; n9886
g7451 and pi0075 n9703_not ; n9887
g7452 and pi0100 n9703_not ; n9888
g7453 and n9282 n9694_not ; n9889
g7454 and n9249 n9889_not ; n9890
g7455 nor pi0100 n9890 ; n9891
g7456 and pi0232_not n9282 ; n9892
g7457 nor n9891 n9892 ; n9893
g7458 nor n9866 n9893 ; n9894
g7459 nor n9888 n9894 ; n9895
g7460 nor pi0075 n9895 ; n9896
g7461 nor pi0092 n9887 ; n9897
g7462 and n9896_not n9897 ; n9898
g7463 nor n9886 n9898 ; n9899
g7464 nor n9865 n9899 ; n9900
g7465 nor pi0074 n9900 ; n9901
g7466 and n9864 n9901_not ; n9902
g7467 and pi0146 n9646 ; n9903
g7468 nor pi0146 n9640 ; n9904
g7469 nor pi0161 n9903 ; n9905
g7470 and n9904_not n9905 ; n9906
g7471 and pi0146 n9648 ; n9907
g7472 nor pi0146 n9638 ; n9908
g7473 and pi0161 n9907_not ; n9909
g7474 and n9908_not n9909 ; n9910
g7475 nor n9906 n9910 ; n9911
g7476 and pi0162 n9911_not ; n9912
g7477 nor pi0161 n9606 ; n9913
g7478 and pi0161 n9574_not ; n9914
g7479 and pi0146 n9913_not ; n9915
g7480 and n9914_not n9915 ; n9916
g7481 nor pi0161 n9615 ; n9917
g7482 and pi0161 n9612_not ; n9918
g7483 nor pi0146 n9917 ; n9919
g7484 and n9918_not n9919 ; n9920
g7485 nor pi0162 n9575 ; n9921
g7486 and n9916_not n9921 ; n9922
g7487 and n9920_not n9922 ; n9923
g7488 nor n9912 n9923 ; n9924
g7489 and n9793 n9924_not ; n9925
g7490 and pi0142 n9391 ; n9926
g7491 nor pi0142 n9497 ; n9927
g7492 nor pi0140 n9926 ; n9928
g7493 and n9927_not n9928 ; n9929
g7494 and pi0142 n9445_not ; n9930
g7495 and n9511_not n9930 ; n9931
g7496 nor pi0142 n9507 ; n9932
g7497 and pi0140 n9931_not ; n9933
g7498 and n9932_not n9933 ; n9934
g7499 nor n9929 n9934 ; n9935
g7500 nor pi0181 n9935 ; n9936
g7501 nor pi0142 n9544 ; n9937
g7502 and pi0142 n9458_not ; n9938
g7503 nor pi0140 n9938 ; n9939
g7504 and n9937_not n9939 ; n9940
g7505 and pi0142 n9453_not ; n9941
g7506 nor pi0142 n9541 ; n9942
g7507 and pi0140 n9941_not ; n9943
g7508 and n9942_not n9943 ; n9944
g7509 nor n9940 n9944 ; n9945
g7510 and pi0181 n9945_not ; n9946
g7511 and pi0144 n9946_not ; n9947
g7512 and n9936_not n9947 ; n9948
g7513 and n9408_not n9604 ; n9949
g7514 and n6197 n9949_not ; n9950
g7515 and pi0142 n9950_not ; n9951
g7516 and n9511_not n9951 ; n9952
g7517 and pi0142_not n9529 ; n9953
g7518 nor pi0140 n9952 ; n9954
g7519 and n9953_not n9954 ; n9955
g7520 and pi0142 n9645_not ; n9956
g7521 and n9511_not n9956 ; n9957
g7522 nor pi0142 n9534 ; n9958
g7523 and pi0140 n9957_not ; n9959
g7524 and n9958_not n9959 ; n9960
g7525 nor n9955 n9960 ; n9961
g7526 nor pi0181 n9961 ; n9962
g7527 and pi0142 n9414_not ; n9963
g7528 nor pi0142 n9562 ; n9964
g7529 nor pi0140 n9963 ; n9965
g7530 and n9964_not n9965 ; n9966
g7531 and pi0142_not n9548 ; n9967
g7532 and pi0142 n9430_not ; n9968
g7533 and pi0140 n9967_not ; n9969
g7534 and n9968_not n9969 ; n9970
g7535 nor n9966 n9970 ; n9971
g7536 and pi0181 n9971_not ; n9972
g7537 nor pi0144 n9962 ; n9973
g7538 and n9972_not n9973 ; n9974
g7539 nor pi0299 n9974 ; n9975
g7540 and n9948_not n9975 ; n9976
g7541 and pi0146 n9583 ; n9977
g7542 nor pi0146 n9597 ; n9978
g7543 and pi0161 n9977_not ; n9979
g7544 and n9978_not n9979 ; n9980
g7545 and pi0146 n9578_not ; n9981
g7546 nor pi0146 n9592 ; n9982
g7547 nor pi0161 n9981 ; n9983
g7548 and n9982_not n9983 ; n9984
g7549 nor pi0162 n9980 ; n9985
g7550 and n9984_not n9985 ; n9986
g7551 and pi0146_not n9632 ; n9987
g7552 and pi0146 n9626_not ; n9988
g7553 nor pi0161 n9987 ; n9989
g7554 and n9988_not n9989 ; n9990
g7555 and pi0146 n9624_not ; n9991
g7556 nor pi0146 n9630 ; n9992
g7557 and pi0161 n9991_not ; n9993
g7558 and n9992_not n9993 ; n9994
g7559 and pi0162 n9990_not ; n9995
g7560 and n9994_not n9995 ; n9996
g7561 and n9794 n9986_not ; n9997
g7562 and n9996_not n9997 ; n9998
g7563 nor n9925 n9998 ; n9999
g7564 and n9976_not n9999 ; n10000
g7565 and pi0232 n10000_not ; n10001
g7566 nor n9661 n10001 ; n10002
g7567 and n2530 n10002_not ; n10003
g7568 and pi0144 n9307 ; n10004
g7569 nor pi0144 n9304 ; n10005
g7570 and n9338_not n10005 ; n10006
g7571 and n9772 n10006_not ; n10007
g7572 and n10004_not n10007 ; n10008
g7573 nor n9304 n9315 ; n10009
g7574 and n9776 n10005_not ; n10010
g7575 and n10009_not n10010 ; n10011
g7576 nor n10008 n10011 ; n10012
g7577 and pi0232 n10012_not ; n10013
g7578 nor n9310 n10013 ; n10014
g7579 nor pi0038 n10014 ; n10015
g7580 and pi0161_not n9327 ; n10016
g7581 nor n9301 n10016 ; n10017
g7582 and n9036 n10017_not ; n10018
g7583 and n9291 n9766 ; n10019
g7584 and n10018_not n10019 ; n10020
g7585 and pi0161 n9320 ; n10021
g7586 and n9036 n9297 ; n10022
g7587 and n10021_not n10022 ; n10023
g7588 and n9291 n9760 ; n10024
g7589 and n10023_not n10024 ; n10025
g7590 nor n10020 n10025 ; n10026
g7591 and pi0232 n10026_not ; n10027
g7592 nor n10015 n10027 ; n10028
g7593 and pi0039 n10028_not ; n10029
g7594 nor pi0087 n9759 ; n10030
g7595 and n10029_not n10030 ; n10031
g7596 and n10003_not n10031 ; n10032
g7597 and pi0038 n9747_not ; n10033
g7598 nor n9266 n10033 ; n10034
g7599 and pi0087 n10034 ; n10035
g7600 nor pi0100 n10035 ; n10036
g7601 and n10032_not n10036 ; n10037
g7602 nor n9733 n10037 ; n10038
g7603 and n2569 n10038_not ; n10039
g7604 and pi0038_not n9848 ; n10040
g7605 and n7473 n10040_not ; n10041
g7606 and n9282 n10041_not ; n10042
g7607 and n10034 n10042_not ; n10043
g7608 nor pi0100 n10043 ; n10044
g7609 nor n9733 n10044 ; n10045
g7610 and n9205 n10045_not ; n10046
g7611 nor n9734 n10046 ; n10047
g7612 and n10039_not n10047 ; n10048
g7613 nor pi0054 n10048 ; n10049
g7614 nor n9751 n10049 ; n10050
g7615 nor pi0074 n10050 ; n10051
g7616 and n9743 n10051_not ; n10052
g7617 and n2529 n9902_not ; n10053
g7618 and n10052_not n10053 ; n10054
g7619 nor n9884 n10054 ; n10055
g7620 nor n9713 n10055 ; n10056
g7621 and pi0034_not n10056 ; n10057
g7622 nor pi0033 pi0954 ; n10058
g7623 nor n9881 n10058 ; n10059
g7624 and n10057_not n10059 ; n10060
g7625 nor pi0034 n8978 ; n10061
g7626 and n9880 n10061 ; n10062
g7627 and n10056 n10061_not ; n10063
g7628 and n10058 n10062_not ; n10064
g7629 and n10063_not n10064 ; n10065
g7630 nor n10060 n10065 ; po0192
g7631 and n2529 n2572 ; n10067
g7632 and n8962 n10067 ; n10068
g7633 and pi0055_not n10068 ; n10069
g7634 and pi0059 n10069_not ; n10070
g7635 and pi0024_not n7340 ; n10071
g7636 and pi0054 n10071_not ; n10072
g7637 and pi0137 n8884 ; n10073
g7638 and n2923 n2930 ; n10074
g7639 and n7417 n10074_not ; n10075
g7640 and pi0683 n10075 ; n10076
g7641 and pi0252 po1057 ; n10077
g7642 and n10076_not n10077 ; n10078
g7643 and pi0146 n7471 ; n10079
g7644 and pi0142 n7470 ; n10080
g7645 nor n10079 n10080 ; n10081
g7646 and n7472_not n10081 ; n10082
g7647 nor n10078 n10082 ; n10083
g7648 nor n7474 n10083 ; n10084
g7649 nor n8886 n10084 ; n10085
g7650 and n6263 n8889_not ; n10086
g7651 and n10078_not n10086 ; n10087
g7652 nor n10085 n10087 ; n10088
g7653 and n8887 n10088_not ; n10089
g7654 nor n10073 n10089 ; n10090
g7655 and n8882 n10090_not ; n10091
g7656 and pi0090_not n6138 ; n10092
g7657 nor pi0093 n10092 ; n10093
g7658 nor n6157 n10093 ; n10094
g7659 nor pi0035 n10094 ; n10095
g7660 and pi0035 n2915_not ; n10096
g7661 and n8938 n10096_not ; n10097
g7662 and n10095_not n10097 ; n10098
g7663 and pi0032_not n10098 ; n10099
g7664 and pi0032 pi0093_not ; n10100
g7665 and n8895 n10100 ; n10101
g7666 and n7432 n10101 ; n10102
g7667 nor n10099 n10102 ; n10103
g7668 nor pi0095 n6169 ; n10104
g7669 and n10103_not n10104 ; n10105
g7670 and n6169 n10095_not ; n10106
g7671 nor pi0137 n6169 ; n10107
g7672 and n2924 n7479 ; n10108
g7673 nor n7425 n10107 ; n10109
g7674 and n10108 n10109 ; n10110
g7675 nor pi0122 po0740 ; n10111
g7676 and n7425 n10107_not ; n10112
g7677 and n10111 n10112 ; n10113
g7678 nor n10110 n10113 ; n10114
g7679 and n10106_not n10114 ; n10115
g7680 and n2704 n8932 ; n10116
g7681 and n10095 n10116_not ; n10117
g7682 and n2518 n10097 ; n10118
g7683 and n10117_not n10118 ; n10119
g7684 and n10115_not n10119 ; n10120
g7685 nor n2743 n10098 ; n10121
g7686 and pi1082 n2518 ; n10122
g7687 and n10121_not n10122 ; n10123
g7688 nor pi0038 n10120 ; n10124
g7689 and n10123_not n10124 ; n10125
g7690 and n10105_not n10125 ; n10126
g7691 and pi0038 n8962_not ; n10127
g7692 nor pi0039 pi0100 ; n10128
g7693 and n10127_not n10128 ; n10129
g7694 and n10126_not n10129 ; n10130
g7695 nor n10091 n10130 ; n10131
g7696 and n2533 n10131_not ; n10132
g7697 and pi0137 po0840_not ; n10133
g7698 and n6282_not n10133 ; n10134
g7699 nor n8964 n10134 ; n10135
g7700 and n8967 n10135_not ; n10136
g7701 and n8962 n10136 ; n10137
g7702 nor n10132 n10137 ; n10138
g7703 nor pi0092 n10138 ; n10139
g7704 nor pi0054 n10139 ; n10140
g7705 and n2529 n8879 ; n10141
g7706 and n10072_not n10141 ; n10142
g7707 and n10140_not n10142 ; n10143
g7708 nor pi0059 n10143 ; n10144
g7709 nor pi0057 n10070 ; n10145
g7710 and n10144_not n10145 ; po0193
g7711 and n2717 n2771 ; n10147
g7712 and pi0065_not n2462 ; n10148
g7713 and n2487 n10148 ; n10149
g7714 and n9081 n10149 ; n10150
g7715 and pi0069_not n10150 ; n10151
g7716 nor pi0067 pi0071 ; n10152
g7717 and pi0083_not n2802 ; n10153
g7718 and pi0036 pi0103_not ; n10154
g7719 and n10152 n10154 ; n10155
g7720 and n10151 n10155 ; n10156
g7721 and n10153 n10156 ; n10157
g7722 and n10147 n10157 ; n10158
g7723 and pi0058_not n7522 ; n10159
g7724 nor n10158 n10159 ; n10160
g7725 and n2704 n6479 ; n10161
g7726 and n6170 n10161 ; n10162
g7727 and n2532 po1038_not ; n10163
g7728 and n3373 n10163 ; n10164
g7729 and pi0092_not n10164 ; n10165
g7730 and n10162 n10165 ; n10166
g7731 and po0740 n10166 ; n10167
g7732 and n10160_not n10167 ; po0194
g7733 nor pi0081 n2789 ; n10169
g7734 nor pi0045 pi0073 ; n10170
g7735 and n8920 n10170 ; n10171
g7736 and pi0071_not n2487 ; n10172
g7737 and pi0104_not n2472 ; n10173
g7738 and n10172 n10173 ; n10174
g7739 nor pi0048 pi0065 ; n10175
g7740 nor pi0082 pi0084 ; n10176
g7741 and pi0089 n10176 ; n10177
g7742 and n10175 n10177 ; n10178
g7743 and n10171 n10178 ; n10179
g7744 and n9080 n10179 ; n10180
g7745 and n10174 n10180 ; n10181
g7746 and pi0332 n10181 ; n10182
g7747 nor pi0064 n10182 ; n10183
g7748 and n6479 n9468 ; n10184
g7749 and n2501 n10184 ; n10185
g7750 and n2508 n10185 ; n10186
g7751 nor pi0039 pi0841 ; n10187
g7752 and n2465 n10187 ; n10188
g7753 and n10183_not n10188 ; n10189
g7754 and n10186 n10189 ; n10190
g7755 and n10169 n10190 ; n10191
g7756 nor pi0038 n10191 ; n10192
g7757 and pi0039_not n2519 ; n10193
g7758 and pi0024 n10193 ; n10194
g7759 and n2709 n10194 ; n10195
g7760 and pi0038 n10195_not ; n10196
g7761 and n2571 po1038_not ; n10197
g7762 and n10192_not n10197 ; n10198
g7763 and n10196_not n10198 ; po0196
g7764 and pi0038_not n10197 ; n10200
g7765 and pi0786 pi1082_not ; n10201
g7766 nor pi0984 n2932 ; n10202
g7767 and pi0835 n10202_not ; n10203
g7768 and n6183 n10203_not ; n10204
g7769 and n6217 n10204_not ; n10205
g7770 and pi1093 n10205 ; n10206
g7771 and n6184 n6380 ; n10207
g7772 and n10206_not n10207 ; n10208
g7773 and pi0223_not n10208 ; n10209
g7774 and n6198 n10205 ; n10210
g7775 and n10207 n10210_not ; n10211
g7776 and n6205 n10211 ; n10212
g7777 and n6227_not n10205 ; n10213
g7778 and n10207 n10213_not ; n10214
g7779 and n6205_not n10214 ; n10215
g7780 nor pi0299 n10212 ; n10216
g7781 and n10215_not n10216 ; n10217
g7782 and n10209_not n10217 ; n10218
g7783 and pi0215_not n10208 ; n10219
g7784 and n6242 n10211 ; n10220
g7785 and n6242_not n10214 ; n10221
g7786 and pi0299 n10220_not ; n10222
g7787 and n10221_not n10222 ; n10223
g7788 and n10219_not n10223 ; n10224
g7789 nor n10201 n10218 ; n10225
g7790 and n10224_not n10225 ; n10226
g7791 and n5853 n6244_not ; n10227
g7792 and n3470 n6207_not ; n10228
g7793 nor n10227 n10228 ; n10229
g7794 and po0740 n10201 ; n10230
g7795 and n10229_not n10230 ; n10231
g7796 and n6382 n10231 ; n10232
g7797 nor n10226 n10232 ; n10233
g7798 and pi0039 n10233_not ; n10234
g7799 nor pi0039 pi0095 ; n10235
g7800 and n6169 n6486 ; n10236
g7801 nor pi0986 po0740 ; n10237
g7802 and pi0252 n10237_not ; n10238
g7803 and pi0314 n10238_not ; n10239
g7804 and pi0108 n2714 ; n10240
g7805 and n2773 n10240 ; n10241
g7806 and pi0841_not n2494 ; n10242
g7807 and n2720 n10242 ; n10243
g7808 and n2714 n2774_not ; n10244
g7809 and n8921 n9076 ; n10245
g7810 nor pi0065 pi0069 ; n10246
g7811 and n10245 n10246 ; n10247
g7812 and pi0048 pi0049_not ; n10248
g7813 nor pi0068 pi0082 ; n10249
g7814 and n10248 n10249 ; n10250
g7815 and n10170 n10250 ; n10251
g7816 and n8910 n8914 ; n10252
g7817 and n9078 n10252 ; n10253
g7818 and n10247 n10251 ; n10254
g7819 and n10253 n10254 ; n10255
g7820 and n10174 n10255 ; n10256
g7821 and pi0097_not n10243 ; n10257
g7822 and n10256 n10257 ; n10258
g7823 and n10244 n10258 ; n10259
g7824 nor pi0047 n10241 ; n10260
g7825 and n10259_not n10260 ; n10261
g7826 and n6151 n10239 ; n10262
g7827 and n10261_not n10262 ; n10263
g7828 nor pi0047 pi0841 ; n10264
g7829 and n10256 n10264 ; n10265
g7830 nor n2760 n10265 ; n10266
g7831 and n2500 n2700 ; n10267
g7832 and n10239_not n10267 ; n10268
g7833 and n10266_not n10268 ; n10269
g7834 nor n10263 n10269 ; n10270
g7835 and n2704 n10270_not ; n10271
g7836 nor pi0035 n10271 ; n10272
g7837 and pi0035 n6483_not ; n10273
g7838 and n2508 n10273_not ; n10274
g7839 and n2510 n10274 ; n10275
g7840 and n10272_not n10275 ; n10276
g7841 nor n10236 n10276 ; n10277
g7842 and n10235 n10277_not ; n10278
g7843 nor n10234 n10278 ; n10279
g7844 and n10200 n10279_not ; po0197
g7845 and pi0093_not pi0102 ; n10281
g7846 and n2461 n10281 ; n10282
g7847 and n2464 n10282 ; n10283
g7848 and n6170 n10283 ; n10284
g7849 and n2501 n10284 ; n10285
g7850 and n2490 n10285 ; n10286
g7851 and n6479 n10286 ; n10287
g7852 and pi1082 n10287_not ; n10288
g7853 and n2518 n3411_not ; n10289
g7854 nor pi0040 n10286 ; n10290
g7855 and n10289 n10290_not ; n10291
g7856 nor pi1082 n10291 ; n10292
g7857 and n10165 n10288_not ; n10293
g7858 and n10292_not n10293 ; po0198
g7859 and pi0189_not n6197 ; n10295
g7860 and pi0144 n10295 ; n10296
g7861 and pi0174_not n10296 ; n10297
g7862 nor pi0299 n10297 ; n10298
g7863 and pi0166_not n6197 ; n10299
g7864 and pi0161 n10299 ; n10300
g7865 and pi0152_not n10300 ; n10301
g7866 nor n7470 n10301 ; n10302
g7867 and pi0232 n10298_not ; n10303
g7868 and n10302_not n10303 ; n10304
g7869 nor pi0072 n10304 ; n10305
g7870 and pi0039 n10305_not ; n10306
g7871 nor pi0041 pi0072 ; n10307
g7872 nor pi0039 n10307 ; n10308
g7873 nor n10306 n10308 ; n10309
g7874 and n2620_not n10309 ; n10310
g7875 nor n7506 n10307 ; n10311
g7876 and n2924_not n10307 ; n10312
g7877 and n7506 n10312_not ; n10313
g7878 and pi0041_not pi0072 ; n10314
g7879 and n2924 n10314_not ; n10315
g7880 and pi0044_not n2521 ; n10316
g7881 and pi0101_not n10316 ; n10317
g7882 and n7479 n10317 ; n10318
g7883 and n7477 n10318 ; n10319
g7884 and pi0041 n10319_not ; n10320
g7885 and pi0099_not n6272 ; n10321
g7886 and pi0072_not pi0101 ; n10322
g7887 nor pi0041 n10322 ; n10323
g7888 and pi0252 n6479 ; n10324
g7889 and pi0024_not n2709 ; n10325
g7890 and n7479 n10324 ; n10326
g7891 and n10325 n10326 ; n10327
g7892 and pi0044_not n10327 ; n10328
g7893 and n10323 n10328 ; n10329
g7894 and n10321_not n10329 ; n10330
g7895 and n10315 n10330_not ; n10331
g7896 and n10320_not n10331 ; n10332
g7897 and n10313 n10332_not ; n10333
g7898 nor n10311 n10333 ; n10334
g7899 nor pi0039 n10334 ; n10335
g7900 and n2620 n10306_not ; n10336
g7901 and n10335_not n10336 ; n10337
g7902 and pi0075 n10310_not ; n10338
g7903 and n10337_not n10338 ; n10339
g7904 and n2608_not n10308 ; n10340
g7905 and pi0228_not n10307 ; n10341
g7906 and n2709 n6479 ; n10342
g7907 and pi0044_not n10342 ; n10343
g7908 and n10323 n10343 ; n10344
g7909 nor n10314 n10344 ; n10345
g7910 and pi0041 n10317_not ; n10346
g7911 and pi0228 n10345 ; n10347
g7912 and n10346_not n10347 ; n10348
g7913 and n2625 n10341_not ; n10349
g7914 and n10348_not n10349 ; n10350
g7915 and pi0087 n10340_not ; n10351
g7916 and n10306_not n10351 ; n10352
g7917 and n10350_not n10352 ; n10353
g7918 and pi0038 n10309_not ; n10354
g7919 and pi0041 n10318_not ; n10355
g7920 and n2924 n10321_not ; n10356
g7921 nor n10315 n10356 ; n10357
g7922 nor pi0072 n7479 ; n10358
g7923 nor n10345 n10358 ; n10359
g7924 and n10321_not n10359 ; n10360
g7925 nor n10355 n10357 ; n10361
g7926 and n10360_not n10361 ; n10362
g7927 and n10313 n10362_not ; n10363
g7928 nor n10311 n10363 ; n10364
g7929 nor pi0039 n10364 ; n10365
g7930 nor n10306 n10365 ; n10366
g7931 and n6285 n10366_not ; n10367
g7932 and pi0287 n2521 ; n10368
g7933 and n10304 n10368 ; n10369
g7934 nor n10305 n10369 ; n10370
g7935 and pi0039 n10370_not ; n10371
g7936 and pi0901 pi0959_not ; n10372
g7937 and pi0480_not pi0949 ; n10373
g7938 and n2717 n2780 ; n10374
g7939 and n2708 n10374 ; n10375
g7940 and n10373_not n10375 ; n10376
g7941 and n2708 n10373 ; n10377
g7942 and n2700 n2759_not ; n10378
g7943 and pi0109_not n6451 ; n10379
g7944 and n2780 n10379 ; n10380
g7945 nor pi0110 n10380 ; n10381
g7946 and pi0047_not n10377 ; n10382
g7947 and n10378 n10382 ; n10383
g7948 and n10381_not n10383 ; n10384
g7949 and n10372 n10376_not ; n10385
g7950 and n10384_not n10385 ; n10386
g7951 and n2701 n2758 ; n10387
g7952 and pi0110 n10387 ; n10388
g7953 and n10377 n10388 ; n10389
g7954 nor n10372 n10389 ; n10390
g7955 and pi0250_not pi0252 ; n10391
g7956 and n6479 n10391 ; n10392
g7957 and n10390_not n10392 ; n10393
g7958 and n10386_not n10393 ; n10394
g7959 and pi0072_not n10394 ; n10395
g7960 and n10162 n10388 ; n10396
g7961 and n10373 n10391_not ; n10397
g7962 and n10396 n10397 ; n10398
g7963 nor n10395 n10398 ; n10399
g7964 nor pi0044 n10399 ; n10400
g7965 and pi0101_not n10400 ; n10401
g7966 and pi0041 n10401_not ; n10402
g7967 and pi0044 pi0072 ; n10403
g7968 and n6479 n10391_not ; n10404
g7969 and n10389 n10404 ; n10405
g7970 nor pi0072 n10405 ; n10406
g7971 and n10394_not n10406 ; n10407
g7972 nor pi0044 n10407 ; n10408
g7973 nor n10403 n10408 ; n10409
g7974 and pi0101_not n10409 ; n10410
g7975 and n10323 n10410_not ; n10411
g7976 nor n10402 n10411 ; n10412
g7977 nor pi0228 n10412 ; n10413
g7978 nor pi0072 n7451 ; n10414
g7979 and n7457_not n10414 ; n10415
g7980 and n6479 n7455_not ; n10416
g7981 and n7454_not n10416 ; n10417
g7982 and pi0072_not n7457 ; n10418
g7983 and n10417_not n10418 ; n10419
g7984 nor pi1093 n10415 ; n10420
g7985 and n10419_not n10420 ; n10421
g7986 and n10414 n10421_not ; n10422
g7987 nor pi0044 n10422 ; n10423
g7988 nor n10403 n10423 ; n10424
g7989 and pi0101_not n10424 ; n10425
g7990 and n10323 n10425_not ; n10426
g7991 and n7451 n7457_not ; n10427
g7992 nor pi1093 n7459 ; n10428
g7993 and n10427_not n10428 ; n10429
g7994 nor pi0044 n10429 ; n10430
g7995 and pi1093 n7451_not ; n10431
g7996 and n10430 n10431_not ; n10432
g7997 and pi0101_not n10432 ; n10433
g7998 and pi0041 n10433_not ; n10434
g7999 nor n2924 n10434 ; n10435
g8000 and n10426_not n10435 ; n10436
g8001 and n2935 n7443_not ; n10437
g8002 and n2937 n10437 ; n10438
g8003 nor n7522 n10438 ; n10439
g8004 and n2461 n10439_not ; n10440
g8005 and n7434 n10440_not ; n10441
g8006 and n7431 n10441_not ; n10442
g8007 nor pi0051 n10442 ; n10443
g8008 nor n2747 n10443 ; n10444
g8009 nor pi0096 n10444 ; n10445
g8010 and n10416 n10418 ; n10446
g8011 and n10445_not n10446 ; n10447
g8012 nor n10427 n10447 ; n10448
g8013 and pi1093 n10448 ; n10449
g8014 and n10430 n10449_not ; n10450
g8015 and pi0101_not n10450 ; n10451
g8016 and pi0041 n10451_not ; n10452
g8017 and pi0072_not n10448 ; n10453
g8018 and pi1093 n10453_not ; n10454
g8019 nor n10421 n10454 ; n10455
g8020 nor pi0044 n10455 ; n10456
g8021 nor n10403 n10456 ; n10457
g8022 and pi0101_not n10457 ; n10458
g8023 and n10323 n10458_not ; n10459
g8024 and n2924 n10459_not ; n10460
g8025 and n10452_not n10460 ; n10461
g8026 and pi0228 n10436_not ; n10462
g8027 and n10461_not n10462 ; n10463
g8028 nor pi0039 n10413 ; n10464
g8029 and n10463_not n10464 ; n10465
g8030 and n2608 n10371_not ; n10466
g8031 and n10465_not n10466 ; n10467
g8032 nor pi0087 n10354 ; n10468
g8033 and n10367_not n10468 ; n10469
g8034 and n10467_not n10469 ; n10470
g8035 nor pi0075 n10353 ; n10471
g8036 and n10470_not n10471 ; n10472
g8037 nor n10339 n10472 ; n10473
g8038 and n7429 n10473_not ; n10474
g8039 nor n7429 n10309 ; n10475
g8040 nor po1038 n10475 ; n10476
g8041 and n10474_not n10476 ; n10477
g8042 and pi0039 pi0232 ; n10478
g8043 and n10301 n10478 ; n10479
g8044 nor pi0072 n10308 ; n10480
g8045 and po1038 n10480 ; n10481
g8046 and n10479_not n10481 ; n10482
g8047 nor n10477 n10482 ; po0199
g8048 and pi0211 pi0214 ; n10484
g8049 and pi0212 n10484 ; n10485
g8050 nor pi0219 n10485 ; n10486
g8051 and pi0207 pi0208 ; n10487
g8052 and pi0042 pi0072_not ; n10488
g8053 and n2620_not n10488 ; n10489
g8054 nor n7506 n10488 ; n10490
g8055 and pi0115_not n2924 ; n10491
g8056 and n10488 n10491_not ; n10492
g8057 and n7506 n10492_not ; n10493
g8058 and pi0114 n10488_not ; n10494
g8059 and n10491 n10494_not ; n10495
g8060 and n6266 n10328 ; n10496
g8061 and pi0113_not n10496 ; n10497
g8062 and pi0116_not n10497 ; n10498
g8063 and n10488 n10498_not ; n10499
g8064 and n6265 n10317 ; n10500
g8065 and n6269 n10500 ; n10501
g8066 and n7479 n10501 ; n10502
g8067 nor pi0114 n6268 ; n10503
g8068 and n10502 n10503 ; n10504
g8069 and n7477 n10504 ; n10505
g8070 and pi0042_not n10505 ; n10506
g8071 nor pi0114 n10499 ; n10507
g8072 and n10506_not n10507 ; n10508
g8073 and n10495 n10508_not ; n10509
g8074 and n10493 n10509_not ; n10510
g8075 and n2620 n10490_not ; n10511
g8076 and n10510_not n10511 ; n10512
g8077 nor pi0039 n10489 ; n10513
g8078 and n10512_not n10513 ; n10514
g8079 and pi0072_not pi0199 ; n10515
g8080 nor pi0232 n10515 ; n10516
g8081 nor pi0299 n10516 ; n10517
g8082 nor pi0072 n10295 ; n10518
g8083 and pi0199 n10518 ; n10519
g8084 and pi0232 n10519_not ; n10520
g8085 and n10517 n10520_not ; n10521
g8086 and pi0166_not n7473 ; n10522
g8087 nor pi0072 n10522 ; n10523
g8088 and pi0299 n10523 ; n10524
g8089 and pi0039 n10524_not ; n10525
g8090 and n10521_not n10525 ; n10526
g8091 nor n10514 n10526 ; n10527
g8092 and pi0075 n10527_not ; n10528
g8093 nor pi0039 n10488 ; n10529
g8094 and n2608_not n10529 ; n10530
g8095 and n6266 n10343 ; n10531
g8096 and pi0228 n10531 ; n10532
g8097 and n6271 n10532 ; n10533
g8098 and n10488 n10533_not ; n10534
g8099 and pi0228 n10501 ; n10535
g8100 and pi0115_not n10535 ; n10536
g8101 and pi0114_not n10536 ; n10537
g8102 and pi0042_not n10537 ; n10538
g8103 and n2625 n10534_not ; n10539
g8104 and n10538_not n10539 ; n10540
g8105 and pi0087 n10530_not ; n10541
g8106 and n10540_not n10541 ; n10542
g8107 and n10526_not n10542 ; n10543
g8108 and pi0115 n10488_not ; n10544
g8109 and pi0042 pi0114_not ; n10545
g8110 and pi0072 pi0116 ; n10546
g8111 and pi0072 pi0113 ; n10547
g8112 and pi0072 n6265_not ; n10548
g8113 and pi0099_not n10411 ; n10549
g8114 nor n10548 n10549 ; n10550
g8115 nor pi0113 n10550 ; n10551
g8116 nor n10547 n10551 ; n10552
g8117 nor pi0116 n10552 ; n10553
g8118 nor n10546 n10553 ; n10554
g8119 and n10545 n10554_not ; n10555
g8120 and n6265 n10401 ; n10556
g8121 and pi0113_not n10556 ; n10557
g8122 and pi0116_not n10557 ; n10558
g8123 nor pi0042 n10558 ; n10559
g8124 nor n10494 n10559 ; n10560
g8125 and n10555_not n10560 ; n10561
g8126 nor pi0115 n10561 ; n10562
g8127 nor pi0228 n10544 ; n10563
g8128 and n10562_not n10563 ; n10564
g8129 and pi0099_not n10459 ; n10565
g8130 nor n10548 n10565 ; n10566
g8131 nor pi0113 n10566 ; n10567
g8132 nor n10547 n10567 ; n10568
g8133 nor pi0116 n10568 ; n10569
g8134 nor n10546 n10569 ; n10570
g8135 and n10545 n10570_not ; n10571
g8136 and n6265 n10451 ; n10572
g8137 and n6269 n10572 ; n10573
g8138 nor pi0042 n10573 ; n10574
g8139 nor n10494 n10574 ; n10575
g8140 and n10571_not n10575 ; n10576
g8141 and n10491 n10576_not ; n10577
g8142 nor pi0115 n2924 ; n10578
g8143 and n6265 n10433 ; n10579
g8144 and n6269 n10579 ; n10580
g8145 and pi0042_not n10580 ; n10581
g8146 and pi0099_not n10426 ; n10582
g8147 nor n10548 n10582 ; n10583
g8148 nor pi0113 n10583 ; n10584
g8149 nor n10547 n10584 ; n10585
g8150 nor pi0116 n10585 ; n10586
g8151 nor n10546 n10586 ; n10587
g8152 and pi0042 n10587 ; n10588
g8153 nor pi0114 n10581 ; n10589
g8154 and n10588_not n10589 ; n10590
g8155 nor n10494 n10590 ; n10591
g8156 and n10578 n10591_not ; n10592
g8157 and pi0228 n10544_not ; n10593
g8158 and n10592_not n10593 ; n10594
g8159 and n10577_not n10594 ; n10595
g8160 nor pi0039 n10564 ; n10596
g8161 and n10595_not n10596 ; n10597
g8162 and pi0232 pi0299 ; n10598
g8163 and n10299 n10368 ; n10599
g8164 and n10523_not n10598 ; n10600
g8165 and n10599_not n10600 ; n10601
g8166 and pi0232 pi0299_not ; n10602
g8167 and n6197 n10368 ; n10603
g8168 and pi0189_not n10603 ; n10604
g8169 nor n10518 n10604 ; n10605
g8170 and pi0199 n10605_not ; n10606
g8171 and n10602 n10606_not ; n10607
g8172 and pi0072 pi0232_not ; n10608
g8173 and pi0299 n10608_not ; n10609
g8174 and n10516 n10609_not ; n10610
g8175 nor n10601 n10610 ; n10611
g8176 and n10607_not n10611 ; n10612
g8177 and pi0039 n10612_not ; n10613
g8178 nor n10597 n10613 ; n10614
g8179 and n2608 n10614_not ; n10615
g8180 and n6269 n10531 ; n10616
g8181 nor pi0072 n10616 ; n10617
g8182 nor n10358 n10617 ; n10618
g8183 and pi0042 n10618_not ; n10619
g8184 and pi0042_not n10504 ; n10620
g8185 nor pi0114 n10619 ; n10621
g8186 and n10620_not n10621 ; n10622
g8187 and n10495 n10622_not ; n10623
g8188 and n10493 n10623_not ; n10624
g8189 nor n10490 n10624 ; n10625
g8190 nor pi0039 n10625 ; n10626
g8191 nor n10526 n10626 ; n10627
g8192 and n6285 n10627_not ; n10628
g8193 nor n10526 n10529 ; n10629
g8194 and pi0038 n10629_not ; n10630
g8195 nor pi0087 n10630 ; n10631
g8196 and n10628_not n10631 ; n10632
g8197 and n10615_not n10632 ; n10633
g8198 nor pi0075 n10543 ; n10634
g8199 and n10633_not n10634 ; n10635
g8200 and n7429 n10528_not ; n10636
g8201 and n10635_not n10636 ; n10637
g8202 nor n10487 n10637 ; n10638
g8203 and pi0072_not pi0200 ; n10639
g8204 nor pi0232 n10639 ; n10640
g8205 nor pi0299 n10640 ; n10641
g8206 and pi0200 n10518 ; n10642
g8207 and pi0232 n10642_not ; n10643
g8208 and n10641 n10643_not ; n10644
g8209 and pi0039 n10644_not ; n10645
g8210 and n10521_not n10645 ; n10646
g8211 nor n10529 n10646 ; n10647
g8212 and n7429_not n10647 ; n10648
g8213 and n10487 n10648_not ; n10649
g8214 and n10526 n10645 ; n10650
g8215 nor n10514 n10650 ; n10651
g8216 and pi0075 n10651_not ; n10652
g8217 nor n10626 n10650 ; n10653
g8218 and n6285 n10653_not ; n10654
g8219 and pi0038 n10647_not ; n10655
g8220 nor pi0087 n10655 ; n10656
g8221 nor n10631 n10656 ; n10657
g8222 and pi0232 n10606_not ; n10658
g8223 and pi0200 n10605_not ; n10659
g8224 and n10658 n10659_not ; n10660
g8225 and pi0299_not n10660 ; n10661
g8226 and n10610 n10639_not ; n10662
g8227 nor n10601 n10662 ; n10663
g8228 and n10661_not n10663 ; n10664
g8229 and pi0039 n10664_not ; n10665
g8230 nor n10597 n10665 ; n10666
g8231 and n2608 n10666_not ; n10667
g8232 nor n10654 n10657 ; n10668
g8233 and n10667_not n10668 ; n10669
g8234 and n10541 n10650_not ; n10670
g8235 and n10540_not n10670 ; n10671
g8236 nor pi0075 n10671 ; n10672
g8237 and n10669_not n10672 ; n10673
g8238 and n7429 n10652_not ; n10674
g8239 and n10673_not n10674 ; n10675
g8240 and n10649 n10675_not ; n10676
g8241 nor n10638 n10676 ; n10677
g8242 and n7429_not n10629 ; n10678
g8243 nor n10486 n10678 ; n10679
g8244 and n10677_not n10679 ; n10680
g8245 and pi0039 n10521_not ; n10681
g8246 nor n10514 n10681 ; n10682
g8247 and pi0075 n10682_not ; n10683
g8248 and n10542 n10681_not ; n10684
g8249 nor n10626 n10681 ; n10685
g8250 and n6285 n10685_not ; n10686
g8251 nor n10529 n10681 ; n10687
g8252 and pi0038 n10687_not ; n10688
g8253 and n10517 n10658_not ; n10689
g8254 and pi0039 n10689_not ; n10690
g8255 nor n10597 n10690 ; n10691
g8256 and n2608 n10691_not ; n10692
g8257 nor pi0087 n10688 ; n10693
g8258 and n10686_not n10693 ; n10694
g8259 and n10692_not n10694 ; n10695
g8260 nor pi0075 n10684 ; n10696
g8261 and n10695_not n10696 ; n10697
g8262 and n7429 n10683_not ; n10698
g8263 and n10697_not n10698 ; n10699
g8264 and n7429_not n10687 ; n10700
g8265 nor n10487 n10700 ; n10701
g8266 and n10699_not n10701 ; n10702
g8267 nor n10514 n10646 ; n10703
g8268 and pi0075 n10703_not ; n10704
g8269 and n10542 n10646_not ; n10705
g8270 nor n10517 n10641 ; n10706
g8271 nor n10660 n10706 ; n10707
g8272 and pi0039 n10707_not ; n10708
g8273 nor n10597 n10708 ; n10709
g8274 and n2608 n10709_not ; n10710
g8275 nor n10626 n10646 ; n10711
g8276 and n6285 n10711_not ; n10712
g8277 and n10656 n10712_not ; n10713
g8278 and n10710_not n10713 ; n10714
g8279 nor pi0075 n10705 ; n10715
g8280 and n10714_not n10715 ; n10716
g8281 and n7429 n10704_not ; n10717
g8282 and n10716_not n10717 ; n10718
g8283 and n10649 n10718_not ; n10719
g8284 nor n10702 n10719 ; n10720
g8285 and n10486 n10720_not ; n10721
g8286 nor po1038 n10680 ; n10722
g8287 and n10721_not n10722 ; n10723
g8288 and n10486_not n10523 ; n10724
g8289 and pi0039 n10724_not ; n10725
g8290 and po1038 n10529_not ; n10726
g8291 and n10725_not n10726 ; n10727
g8292 or n10723 n10727 ; po0200
g8293 and pi0043 pi0072_not ; n10729
g8294 nor n7506 n10729 ; n10730
g8295 and pi0042_not n6270 ; n10731
g8296 and n2924 n10731 ; n10732
g8297 and n10729 n10732_not ; n10733
g8298 and n7506 n10733_not ; n10734
g8299 nor pi0072 n10498 ; n10735
g8300 and pi0043 n10735 ; n10736
g8301 and pi0043_not pi0052 ; n10737
g8302 and n7477 n10502 ; n10738
g8303 and n10737 n10738 ; n10739
g8304 nor n10736 n10739 ; n10740
g8305 and n10732 n10740_not ; n10741
g8306 and n10734 n10741_not ; n10742
g8307 nor n10730 n10742 ; n10743
g8308 nor pi0039 n10743 ; n10744
g8309 and n2620 n10744_not ; n10745
g8310 nor pi0039 n10729 ; n10746
g8311 nor n2620 n10746 ; n10747
g8312 nor n10745 n10747 ; n10748
g8313 nor n10645 n10748 ; n10749
g8314 and pi0075 n10749_not ; n10750
g8315 and n2608_not n10746 ; n10751
g8316 nor pi0043 n10501 ; n10752
g8317 and pi0043 n10617_not ; n10753
g8318 and pi0228 n10731 ; n10754
g8319 and n10753_not n10754 ; n10755
g8320 and n10752_not n10755 ; n10756
g8321 and n10729 n10754_not ; n10757
g8322 and n2625 n10757_not ; n10758
g8323 and n10756_not n10758 ; n10759
g8324 and pi0087 n10751_not ; n10760
g8325 and n10759_not n10760 ; n10761
g8326 and n10645_not n10761 ; n10762
g8327 and n10502 n10737 ; n10763
g8328 and pi0043 n10618_not ; n10764
g8329 nor n10763 n10764 ; n10765
g8330 and n10732 n10765_not ; n10766
g8331 and n10734 n10766_not ; n10767
g8332 nor n10730 n10767 ; n10768
g8333 nor pi0039 n10768 ; n10769
g8334 nor n10645 n10769 ; n10770
g8335 and n6285 n10770_not ; n10771
g8336 nor n10645 n10746 ; n10772
g8337 and pi0038 n10772_not ; n10773
g8338 and pi0232 n10659_not ; n10774
g8339 and n10641 n10774_not ; n10775
g8340 and pi0039 n10775_not ; n10776
g8341 nor pi0228 n10558 ; n10777
g8342 nor n2924 n10579 ; n10778
g8343 and n2924 n10572_not ; n10779
g8344 nor n10778 n10779 ; n10780
g8345 and n6269 n10780 ; n10781
g8346 and pi0228 n10781_not ; n10782
g8347 nor n10777 n10782 ; n10783
g8348 nor pi0043 n10783 ; n10784
g8349 nor n10729 n10731 ; n10785
g8350 nor n2924 n10587 ; n10786
g8351 and n2924 n10570_not ; n10787
g8352 nor n10786 n10787 ; n10788
g8353 and pi0228 n10788_not ; n10789
g8354 nor pi0228 n10554 ; n10790
g8355 nor n10789 n10790 ; n10791
g8356 and pi0043 n10731 ; n10792
g8357 and n10791_not n10792 ; n10793
g8358 nor n10784 n10785 ; n10794
g8359 and n10793_not n10794 ; n10795
g8360 nor pi0039 n10795 ; n10796
g8361 nor n10776 n10796 ; n10797
g8362 and n2608 n10797_not ; n10798
g8363 nor pi0087 n10773 ; n10799
g8364 and n10771_not n10799 ; n10800
g8365 and n10798_not n10800 ; n10801
g8366 nor pi0075 n10762 ; n10802
g8367 and n10801_not n10802 ; n10803
g8368 and n7429 n10750_not ; n10804
g8369 and n10803_not n10804 ; n10805
g8370 and n7429_not n10772 ; n10806
g8371 nor n10487 n10806 ; n10807
g8372 and n10805_not n10807 ; n10808
g8373 nor pi0199 pi0200 ; n10809
g8374 nor pi0299 n10809 ; n10810
g8375 nor pi0072 n10810 ; n10811
g8376 nor pi0232 n10811 ; n10812
g8377 nor pi0299 n10812 ; n10813
g8378 and n10518 n10809 ; n10814
g8379 and pi0232 n10814_not ; n10815
g8380 and n10813 n10815_not ; n10816
g8381 and pi0039 n10816_not ; n10817
g8382 nor n10746 n10817 ; n10818
g8383 and n7429_not n10818 ; n10819
g8384 nor n10748 n10817 ; n10820
g8385 and pi0075 n10820_not ; n10821
g8386 nor n10769 n10817 ; n10822
g8387 and n6285 n10822_not ; n10823
g8388 and pi0038 n10818_not ; n10824
g8389 and n10605_not n10809 ; n10825
g8390 and pi0232 n10825_not ; n10826
g8391 and n10813 n10826_not ; n10827
g8392 and pi0039 n10827_not ; n10828
g8393 nor n10796 n10828 ; n10829
g8394 and n2608 n10829_not ; n10830
g8395 nor pi0087 n10824 ; n10831
g8396 and n10823_not n10831 ; n10832
g8397 and n10830_not n10832 ; n10833
g8398 nor n2531 n10818 ; n10834
g8399 and n10761 n10834_not ; n10835
g8400 nor pi0075 n10835 ; n10836
g8401 and n10833_not n10836 ; n10837
g8402 and n7429 n10821_not ; n10838
g8403 and n10837_not n10838 ; n10839
g8404 and n10487 n10819_not ; n10840
g8405 and n10839_not n10840 ; n10841
g8406 nor n10808 n10841 ; n10842
g8407 and pi0212 pi0214 ; n10843
g8408 nor pi0211 pi0219 ; n10844
g8409 and n10843 n10844_not ; n10845
g8410 nor pi0211 n10843 ; n10846
g8411 nor n10845 n10846 ; n10847
g8412 nor n10842 n10847 ; n10848
g8413 and n10525 n10644_not ; n10849
g8414 nor n10748 n10849 ; n10850
g8415 and pi0075 n10850_not ; n10851
g8416 and n10761 n10849_not ; n10852
g8417 nor n10769 n10849 ; n10853
g8418 and n6285 n10853_not ; n10854
g8419 nor n10746 n10849 ; n10855
g8420 and pi0038 n10855_not ; n10856
g8421 and n10602 n10659_not ; n10857
g8422 and n10609_not n10640 ; n10858
g8423 nor n10601 n10858 ; n10859
g8424 and n10857_not n10859 ; n10860
g8425 and pi0039 n10860_not ; n10861
g8426 nor n10796 n10861 ; n10862
g8427 and n2608 n10862_not ; n10863
g8428 nor pi0087 n10856 ; n10864
g8429 and n10854_not n10864 ; n10865
g8430 and n10863_not n10865 ; n10866
g8431 nor pi0075 n10852 ; n10867
g8432 and n10866_not n10867 ; n10868
g8433 and n7429 n10851_not ; n10869
g8434 and n10868_not n10869 ; n10870
g8435 and n7429_not n10855 ; n10871
g8436 nor n10487 n10871 ; n10872
g8437 and n10870_not n10872 ; n10873
g8438 and n10524_not n10817 ; n10874
g8439 nor n10746 n10874 ; n10875
g8440 and n7429_not n10875 ; n10876
g8441 nor n10748 n10874 ; n10877
g8442 and pi0075 n10877_not ; n10878
g8443 and n10761 n10874_not ; n10879
g8444 nor n10769 n10874 ; n10880
g8445 and n6285 n10880_not ; n10881
g8446 and pi0038 n10875_not ; n10882
g8447 and n10602 n10825_not ; n10883
g8448 nor n10601 n10812 ; n10884
g8449 and n10883_not n10884 ; n10885
g8450 and pi0039 n10885_not ; n10886
g8451 nor n10796 n10886 ; n10887
g8452 and n2608 n10887_not ; n10888
g8453 nor pi0087 n10882 ; n10889
g8454 and n10881_not n10889 ; n10890
g8455 and n10888_not n10890 ; n10891
g8456 nor pi0075 n10879 ; n10892
g8457 and n10891_not n10892 ; n10893
g8458 and n7429 n10878_not ; n10894
g8459 and n10893_not n10894 ; n10895
g8460 and n10487 n10876_not ; n10896
g8461 and n10895_not n10896 ; n10897
g8462 nor n10873 n10897 ; n10898
g8463 and n10847 n10898_not ; n10899
g8464 nor po1038 n10848 ; n10900
g8465 and n10899_not n10900 ; n10901
g8466 and n10523 n10847 ; n10902
g8467 and pi0039 n10902_not ; n10903
g8468 and po1038 n10746_not ; n10904
g8469 and n10903_not n10904 ; n10905
g8470 or n10901 n10905 ; po0201
g8471 and pi0072_not n7474 ; n10907
g8472 and pi0039 n10907_not ; n10908
g8473 and pi0044 pi0072_not ; n10909
g8474 nor pi0039 n10909 ; n10910
g8475 nor n10908 n10910 ; n10911
g8476 and n2620_not n10911 ; n10912
g8477 nor n7506 n10909 ; n10913
g8478 nor pi0039 n10913 ; n10914
g8479 and n2924_not n10909 ; n10915
g8480 and n7506 n10915_not ; n10916
g8481 and n7594 n10403_not ; n10917
g8482 and n7479 n10316 ; n10918
g8483 and n7477 n10918 ; n10919
g8484 and pi0044 n10327_not ; n10920
g8485 nor n10919 n10920 ; n10921
g8486 and n10917 n10921_not ; n10922
g8487 and n10916 n10922_not ; n10923
g8488 and n10914 n10923_not ; n10924
g8489 and pi0039 n7474 ; n10925
g8490 and pi0072_not n10925 ; n10926
g8491 nor n10924 n10926 ; n10927
g8492 and n2620 n10927_not ; n10928
g8493 and pi0075 n10912_not ; n10929
g8494 and n10928_not n10929 ; n10930
g8495 and pi0228 n2608 ; n10931
g8496 and n10316 n10931 ; n10932
g8497 and n10342 n10931 ; n10933
g8498 and n10909 n10933_not ; n10934
g8499 nor pi0039 n10934 ; n10935
g8500 and n10932_not n10935 ; n10936
g8501 and pi0087 n10908_not ; n10937
g8502 and n10936_not n10937 ; n10938
g8503 and pi0038 n10911_not ; n10939
g8504 and n7479 n10342 ; n10940
g8505 and pi0044 n10940_not ; n10941
g8506 nor n10918 n10941 ; n10942
g8507 and n10917 n10942_not ; n10943
g8508 and n10916 n10943_not ; n10944
g8509 and n10914 n10944_not ; n10945
g8510 and n6285 n10926_not ; n10946
g8511 and n10945_not n10946 ; n10947
g8512 and pi0287 n10342 ; n10948
g8513 nor pi0072 n10948 ; n10949
g8514 and n10925 n10949 ; n10950
g8515 and pi0044 n10407 ; n10951
g8516 nor pi0228 n10951 ; n10952
g8517 and n10400_not n10952 ; n10953
g8518 and pi0044 n10455 ; n10954
g8519 and n2924 n10450_not ; n10955
g8520 and n10954_not n10955 ; n10956
g8521 and pi0044 n10422 ; n10957
g8522 nor n2924 n10432 ; n10958
g8523 and n10957_not n10958 ; n10959
g8524 nor n10956 n10959 ; n10960
g8525 and pi0228 n10960_not ; n10961
g8526 nor pi0039 n10953 ; n10962
g8527 and n10961_not n10962 ; n10963
g8528 and n2608 n10950_not ; n10964
g8529 and n10963_not n10964 ; n10965
g8530 nor pi0087 n10939 ; n10966
g8531 and n10947_not n10966 ; n10967
g8532 and n10965_not n10967 ; n10968
g8533 nor pi0075 n10938 ; n10969
g8534 and n10968_not n10969 ; n10970
g8535 nor n10930 n10970 ; n10971
g8536 and n7429 n10971_not ; n10972
g8537 nor n7429 n10911 ; n10973
g8538 nor po1038 n10973 ; n10974
g8539 and n10972_not n10974 ; n10975
g8540 and n2639 n7473 ; n10976
g8541 and pi0072_not n10976 ; n10977
g8542 and pi0039 n10977_not ; n10978
g8543 and po1038 n10910_not ; n10979
g8544 and n10978_not n10979 ; n10980
g8545 or n10975 n10980 ; po0202
g8546 and pi0038_not pi0039 ; n10982
g8547 and n10197 n10982 ; n10983
g8548 and pi0979 n10983 ; n10984
g8549 and n6380 n10984 ; po0203
g8550 nor pi0102 pi0104 ; n10986
g8551 and pi0111_not n10986 ; n10987
g8552 nor pi0049 pi0076 ; n10988
g8553 and n8909 n10988 ; n10989
g8554 and pi0061 pi0082_not ; n10990
g8555 nor pi0083 pi0089 ; n10991
g8556 and n10990 n10991 ; n10992
g8557 and n7438 n8915 ; n10993
g8558 and n10992 n10993 ; n10994
g8559 and n10172 n10987 ; n10995
g8560 and n10989 n10995 ; n10996
g8561 and n8912 n10994 ; n10997
g8562 and n10247 n10997 ; n10998
g8563 and n10996 n10998 ; n10999
g8564 and n8935 n10999 ; n11000
g8565 and pi0841_not n11000 ; n11001
g8566 and n2702 n2888 ; n11002
g8567 and pi0024 n11002 ; n11003
g8568 nor n11001 n11003 ; n11004
g8569 and n10166 n11004_not ; po0204
g8570 and pi0082_not n2474 ; n11006
g8571 and pi0084_not pi0104 ; n11007
g8572 and n2805 n11007 ; n11008
g8573 and n10171 n11008 ; n11009
g8574 and n11006 n11009 ; n11010
g8575 nor pi0036 n11010 ; n11011
g8576 and n8916 n9081 ; n11012
g8577 nor pi0067 pi0103 ; n11013
g8578 and n2487 n11013 ; n11014
g8579 and pi0098_not n11014 ; n11015
g8580 and n11012 n11015 ; n11016
g8581 and n11011_not n11016 ; n11017
g8582 and n2803_not n11017 ; n11018
g8583 nor pi0088 n11018 ; n11019
g8584 and n2871_not n7438 ; n11020
g8585 and n2754 n11019_not ; n11021
g8586 and n11020 n11021 ; n11022
g8587 and n2700 n11022 ; n11023
g8588 nor n10159 n11023 ; n11024
g8589 and n10162 n11024_not ; n11025
g8590 and n7490 n11025_not ; n11026
g8591 and pi0036_not n11017 ; n11027
g8592 nor pi0088 n11027 ; n11028
g8593 and n11020 n11028_not ; n11029
g8594 and n10186 n11029 ; n11030
g8595 and pi0824_not n2932 ; n11031
g8596 and n11030 n11031 ; n11032
g8597 and n2932_not n11025 ; n11033
g8598 and pi0829 n11032_not ; n11034
g8599 and n11033_not n11034 ; n11035
g8600 and n2923_not n11035 ; n11036
g8601 nor n11026 n11036 ; n11037
g8602 and pi1091 n11037_not ; n11038
g8603 and n7417_not n11025 ; n11039
g8604 nor pi0829 n11039 ; n11040
g8605 nor n11035 n11040 ; n11041
g8606 nor pi1093 n11041 ; n11042
g8607 and n7417 n10162 ; n11043
g8608 and n10160_not n11043 ; n11044
g8609 nor n6394 n7626 ; n11045
g8610 nor n11044 n11045 ; n11046
g8611 and n11039_not n11046 ; n11047
g8612 and n10165 n11047_not ; n11048
g8613 and n11042_not n11048 ; n11049
g8614 and n11038_not n11049 ; po0205
g8615 and pi0072_not pi0841 ; n11051
g8616 and n2705 n11051 ; n11052
g8617 and pi0051_not n11052 ; n11053
g8618 and n10256 n11053 ; n11054
g8619 and n10165 n11054 ; n11055
g8620 and n10185 n11055 ; po0206
g8621 and n2464 n2487 ; n11057
g8622 and pi0103_not n2804 ; n11058
g8623 and n10245 n11058 ; n11059
g8624 and n8909 n8916 ; n11060
g8625 and n11059 n11060 ; n11061
g8626 and pi0045_not pi0049 ; n11062
g8627 and n10987 n11062 ; n11063
g8628 and n11057 n11063 ; n11064
g8629 and n11061 n11064 ; n11065
g8630 and n11006 n11065 ; n11066
g8631 and n2706 n8935 ; n11067
g8632 and n11066 n11067 ; n11068
g8633 and n10161 n11052 ; n11069
g8634 and n11068 n11069 ; n11070
g8635 nor pi0074 n11070 ; n11071
g8636 and pi0074 n8962_not ; n11072
g8637 and n7363 po1038_not ; n11073
g8638 and n11071_not n11073 ; n11074
g8639 and n11072_not n11074 ; po0207
g8640 and pi0024 n8897 ; n11076
g8641 nor n10374 n11076 ; n11077
g8642 nor pi0252 n8888 ; n11078
g8643 and pi0252 po0840_not ; n11079
g8644 nor n11078 n11079 ; n11080
g8645 and pi0024 pi0094_not ; n11081
g8646 and n8899_not n11081 ; n11082
g8647 and n10162 n11080 ; n11083
g8648 and n11082_not n11083 ; n11084
g8649 and n11077_not n11084 ; n11085
g8650 and n2962 n7450 ; n11086
g8651 and pi0024 pi0090_not ; n11087
g8652 and n11086 n11087 ; n11088
g8653 and n11080_not n11088 ; n11089
g8654 and n8901 n11089 ; n11090
g8655 nor n11085 n11090 ; n11091
g8656 nor pi0100 n11091 ; n11092
g8657 and pi0100 n6263_not ; n11093
g8658 and n6353 n11093 ; n11094
g8659 nor n11092 n11094 ; n11095
g8660 and n2530 n2533 ; n11096
g8661 and n11095_not n11096 ; n11097
g8662 and n6282 n8967 ; n11098
g8663 and n8963 n11098 ; n11099
g8664 nor n11097 n11099 ; n11100
g8665 and n8881 n11100_not ; po0208
g8666 and n9082 n11057 ; n11102
g8667 and n2467 n11102 ; n11103
g8668 and pi0069_not n11103 ; n11104
g8669 and n2804 n11104 ; n11105
g8670 and n2700 n10166 ; n11106
g8671 and n2754 n11106 ; n11107
g8672 and n2807 n11105 ; n11108
g8673 and n11107 n11108 ; po0209
g8674 and pi0219_not n10846 ; n11110
g8675 and pi0052 pi0072_not ; n11111
g8676 nor pi0039 n11111 ; n11112
g8677 nor n10525 n11112 ; n11113
g8678 nor n7429 n11113 ; n11114
g8679 and n10601_not n10609 ; n11115
g8680 and pi0039 n11115_not ; n11116
g8681 and n6267 n6270 ; n11117
g8682 nor n11111 n11117 ; n11118
g8683 and pi0052_not n10558 ; n11119
g8684 and pi0052 n10554 ; n11120
g8685 and n11117 n11119_not ; n11121
g8686 and n11120_not n11121 ; n11122
g8687 nor pi0228 n11118 ; n11123
g8688 and n11122_not n11123 ; n11124
g8689 and pi0114_not n6267 ; n11125
g8690 and pi0052_not n10573 ; n11126
g8691 and pi0052 n10570 ; n11127
g8692 and n10491 n11126_not ; n11128
g8693 and n11127_not n11128 ; n11129
g8694 and pi0052_not n10580 ; n11130
g8695 and pi0052 n10587 ; n11131
g8696 and n10578 n11130_not ; n11132
g8697 and n11131_not n11132 ; n11133
g8698 nor n11129 n11133 ; n11134
g8699 and n11125 n11134_not ; n11135
g8700 and pi0228 n11118_not ; n11136
g8701 and n11135_not n11136 ; n11137
g8702 nor pi0039 n11124 ; n11138
g8703 and n11137_not n11138 ; n11139
g8704 nor n11116 n11139 ; n11140
g8705 and n2608 n11140_not ; n11141
g8706 and pi0038 n11113_not ; n11142
g8707 and n7506 n10491 ; n11143
g8708 and n11125 n11143 ; n11144
g8709 and n7479 n11144 ; n11145
g8710 and n10616 n11145 ; n11146
g8711 and n11111 n11146_not ; n11147
g8712 nor pi0039 n11147 ; n11148
g8713 nor n10525 n11148 ; n11149
g8714 and n6285 n11149_not ; n11150
g8715 nor n11142 n11150 ; n11151
g8716 and n11141_not n11151 ; n11152
g8717 nor pi0087 n11152 ; n11153
g8718 and n2608_not n11113 ; n11154
g8719 and pi0087 n11154_not ; n11155
g8720 and pi0228 n11117 ; n11156
g8721 and pi0052_not n10501 ; n11157
g8722 and pi0052 n10617 ; n11158
g8723 nor n11157 n11158 ; n11159
g8724 and n11156 n11159_not ; n11160
g8725 and n11111 n11156_not ; n11161
g8726 nor n11160 n11161 ; n11162
g8727 and pi0039_not n11162 ; n11163
g8728 and n2608 n10525_not ; n11164
g8729 and n11163_not n11164 ; n11165
g8730 and n11155 n11165_not ; n11166
g8731 and n10487 n11166_not ; n11167
g8732 and n11153_not n11167 ; n11168
g8733 nor n10817 n11112 ; n11169
g8734 and n2608_not n11169 ; n11170
g8735 and n2608 n10874_not ; n11171
g8736 and n11163_not n11171 ; n11172
g8737 and n11155 n11170_not ; n11173
g8738 and n11172_not n11173 ; n11174
g8739 nor n10886 n11139 ; n11175
g8740 and n2608 n11175_not ; n11176
g8741 nor n10874 n11148 ; n11177
g8742 and n6285 n11177_not ; n11178
g8743 and pi0038 n11169_not ; n11179
g8744 and n11113_not n11179 ; n11180
g8745 nor n11178 n11180 ; n11181
g8746 and n11176_not n11181 ; n11182
g8747 nor pi0087 n11182 ; n11183
g8748 nor n10487 n11174 ; n11184
g8749 and n11183_not n11184 ; n11185
g8750 nor n11168 n11185 ; n11186
g8751 nor pi0075 n11186 ; n11187
g8752 and n10498 n11144 ; n11188
g8753 and n2620 n11188 ; n11189
g8754 and pi0039_not n11111 ; n11190
g8755 and n11189_not n11190 ; n11191
g8756 nor pi0039 n11191 ; n11192
g8757 and n10487_not n10874 ; n11193
g8758 and n10487 n10525 ; n11194
g8759 and pi0075 n11194_not ; n11195
g8760 and n11193_not n11195 ; n11196
g8761 and n11192_not n11196 ; n11197
g8762 and n7429 n11197_not ; n11198
g8763 and n11187_not n11198 ; n11199
g8764 and n11110 n11114_not ; n11200
g8765 and n11199_not n11200 ; n11201
g8766 nor n7429 n10487 ; n11202
g8767 and n11169 n11202 ; n11203
g8768 nor n7429 n11190 ; n11204
g8769 and pi0075 n11191 ; n11205
g8770 and pi0100 n11190_not ; n11206
g8771 and pi0038 n11190_not ; n11207
g8772 and pi0038_not n11162 ; n11208
g8773 nor n11207 n11208 ; n11209
g8774 nor pi0100 n11209 ; n11210
g8775 and pi0100_not n10982 ; n11211
g8776 and pi0087 n11211_not ; n11212
g8777 and n11206_not n11212 ; n11213
g8778 and n11210_not n11213 ; n11214
g8779 and pi0100 n11147_not ; n11215
g8780 and pi0100_not n11139 ; n11216
g8781 nor pi0039 n11215 ; n11217
g8782 and n11216_not n11217 ; n11218
g8783 nor pi0038 n11218 ; n11219
g8784 nor pi0087 n11207 ; n11220
g8785 and n11219_not n11220 ; n11221
g8786 nor n11214 n11221 ; n11222
g8787 nor pi0075 n11222 ; n11223
g8788 and n7429 n11205_not ; n11224
g8789 and n11223_not n11224 ; n11225
g8790 and n10487 n11204_not ; n11226
g8791 and n11225_not n11226 ; n11227
g8792 and n2608 n10817_not ; n11228
g8793 and n11163_not n11228 ; n11229
g8794 nor n11170 n11229 ; n11230
g8795 and pi0087 n11230_not ; n11231
g8796 nor n10828 n11139 ; n11232
g8797 and n2608 n11232_not ; n11233
g8798 nor n10817 n11148 ; n11234
g8799 and n6285 n11234_not ; n11235
g8800 nor pi0087 n11179 ; n11236
g8801 and n11235_not n11236 ; n11237
g8802 and n11233_not n11237 ; n11238
g8803 nor pi0075 n11231 ; n11239
g8804 and n11238_not n11239 ; n11240
g8805 and n2620_not n11169 ; n11241
g8806 and n11111 n11188_not ; n11242
g8807 nor pi0039 n11242 ; n11243
g8808 and n2620 n10817_not ; n11244
g8809 and n11243_not n11244 ; n11245
g8810 and pi0075 n11241_not ; n11246
g8811 and n11245_not n11246 ; n11247
g8812 and n7429 n10487_not ; n11248
g8813 and n11247_not n11248 ; n11249
g8814 and n11240_not n11249 ; n11250
g8815 nor n11227 n11250 ; n11251
g8816 nor n11110 n11251 ; n11252
g8817 nor po1038 n11203 ; n11253
g8818 and n11201_not n11253 ; n11254
g8819 and n11252_not n11254 ; n11255
g8820 and pi0039 n11110 ; n11256
g8821 and n10523 n11256 ; n11257
g8822 and po1038 n11190_not ; n11258
g8823 and n11257_not n11258 ; n11259
g8824 nor n11255 n11259 ; po0210
g8825 nor pi0287 pi0979 ; n11261
g8826 and n6181 n11261 ; n11262
g8827 and pi0039 n11262_not ; n11263
g8828 and pi0024 n10162 ; n11264
g8829 and pi0053 n2720 ; n11265
g8830 and n2717 n11265 ; n11266
g8831 and n2721 n11266 ; n11267
g8832 and n11264 n11267 ; n11268
g8833 nor pi0039 n11268 ; n11269
g8834 and n10200 n11263_not ; n11270
g8835 and n11269_not n11270 ; n11271
g8836 and n3402_not n11271 ; po0211
g8837 and n8897 n9254 ; n11273
g8838 nor pi0060 pi0085 ; n11274
g8839 and pi0106 n11274 ; n11275
g8840 and n2479 n8913 ; n11276
g8841 and n11275 n11276 ; n11277
g8842 and n10989 n11277 ; n11278
g8843 and n8919 n11059 ; n11279
g8844 and n11278 n11279 ; n11280
g8845 and n11057 n11280 ; n11281
g8846 and n11273 n11281 ; n11282
g8847 and pi0841_not n2704 ; n11283
g8848 and n8960 n11283 ; n11284
g8849 and n2611 n2706 ; n11285
g8850 and n11284 n11285 ; n11286
g8851 and n11282 n11286 ; n11287
g8852 nor pi0054 n11287 ; n11288
g8853 and n2621 n10195 ; n11289
g8854 and pi0054 n11289_not ; n11290
g8855 and n8880 n11288_not ; n11291
g8856 and n11290_not n11291 ; po0212
g8857 and pi0054_not n11289 ; n11293
g8858 and pi0074_not n11293 ; n11294
g8859 and pi0055 n11294_not ; n11295
g8860 and pi0045 n2479 ; n11296
g8861 and n2487 n11296 ; n11297
g8862 and n11061 n11297 ; n11298
g8863 and n2476 n11298 ; n11299
g8864 and n6479 n9500 ; n11300
g8865 and n2465 n2572 ; n11301
g8866 and n11300 n11301 ; n11302
g8867 and n11299 n11302 ; n11303
g8868 nor pi0055 n11303 ; n11304
g8869 and n8878 n11304_not ; n11305
g8870 and n11295_not n11305 ; po0213
g8871 and n2518 n2537 ; n11307
g8872 and n6172 n11307 ; n11308
g8873 and pi0056 n11308_not ; n11309
g8874 and pi0056 pi0062_not ; n11310
g8875 and pi0055 n10068 ; n11311
g8876 nor n11310 n11311 ; n11312
g8877 and n3328 n11309_not ; n11313
g8878 and n11312_not n11313 ; po0214
g8879 and n6304 n11294 ; n11315
g8880 and pi0057 n11315_not ; n11316
g8881 and n6485 n11307 ; n11317
g8882 and pi0056_not pi0062 ; n11318
g8883 and pi0924_not n11318 ; n11319
g8884 nor n11310 n11319 ; n11320
g8885 and n11317 n11320_not ; n11321
g8886 nor pi0057 n11321 ; n11322
g8887 nor pi0059 n11316 ; n11323
g8888 and n11322_not n11323 ; po0215
g8889 and pi0093_not n11086 ; n11325
g8890 and n10165 n11325 ; n11326
g8891 and n7433 n11326 ; po0216
g8892 and pi0059 n11315_not ; n11328
g8893 and pi0924 n11318 ; n11329
g8894 and n11317 n11329 ; n11330
g8895 nor pi0059 n11330 ; n11331
g8896 nor pi0057 n11328 ; n11332
g8897 and n11331_not n11332 ; po0217
g8898 and pi0039 pi0979_not ; n11334
g8899 and n6181_not n11334 ; n11335
g8900 and n6182 n11335 ; n11336
g8901 and n6380 n11336 ; n11337
g8902 and pi0039_not n11264 ; n11338
g8903 and n11273 n11338 ; n11339
g8904 and n2718 n11339 ; n11340
g8905 nor n11337 n11340 ; n11341
g8906 and n10200 n11341_not ; po0218
g8907 and pi0841 n11000 ; n11343
g8908 and pi0024_not n11273 ; n11344
g8909 and n2718 n11344 ; n11345
g8910 nor n11343 n11345 ; n11346
g8911 and n10166 n11346_not ; po0219
g8912 and pi0057 n10069_not ; n11348
g8913 and n11308 n11318 ; n11349
g8914 nor pi0057 n11349 ; n11350
g8915 nor pi0059 n11348 ; n11351
g8916 and n11350_not n11351 ; po0220
g8917 and n2861 n8935 ; n11353
g8918 and n9100 n11353 ; n11354
g8919 and pi0999 n11354 ; n11355
g8920 and pi0024_not n11002 ; n11356
g8921 nor n11355 n11356 ; n11357
g8922 and n10166 n11357_not ; po0221
g8923 and pi0063_not pi0107 ; n11359
g8924 and n9100 n11359 ; n11360
g8925 nor pi0841 n11360 ; n11361
g8926 and n2486 n11359 ; n11362
g8927 nor pi0064 n11362 ; n11363
g8928 and n2465 n11363_not ; n11364
g8929 and n10169 n11364 ; n11365
g8930 and pi0841 n11365_not ; n11366
g8931 and n11107 n11361_not ; n11367
g8932 and n11366_not n11367 ; po0222
g8933 and pi0039 n10201 ; n11369
g8934 and n10200 n11369 ; n11370
g8935 and n10217_not n11370 ; n11371
g8936 and n10223_not n11371 ; po0223
g8937 and pi0199 pi0299_not ; n11373
g8938 and n2570 n2608 ; n11374
g8939 and pi0314 n2464 ; n11375
g8940 and n11300 n11375 ; n11376
g8941 and pi0081 pi0102_not ; n11377
g8942 and n11376 n11377 ; n11378
g8943 and n2489 n11378 ; n11379
g8944 and n2609 n11373 ; n11380
g8945 and n11374 n11380 ; n11381
g8946 and n11379 n11381 ; n11382
g8947 nor pi0219 n11382 ; n11383
g8948 nor pi0199 pi0299 ; n11384
g8949 and n2572 n11379 ; n11385
g8950 and n11384_not n11385 ; n11386
g8951 and pi0219 n11386_not ; n11387
g8952 nor po1038 n11383 ; n11388
g8953 and n11387_not n11388 ; po0224
g8954 and pi0083 pi0103_not ; n11390
g8955 and n11102 n11390 ; n11391
g8956 and n10165 n11391 ; n11392
g8957 and n11376 n11392 ; n11393
g8958 and n2484 n11393 ; po0225
g8959 and n6244_not n6396 ; n11395
g8960 and n3310 n5853 ; n11396
g8961 and n11395 n11396 ; n11397
g8962 and n6207_not n6396 ; n11398
g8963 and n3351 n3470 ; n11399
g8964 and n11398 n11399 ; n11400
g8965 nor n11397 n11400 ; n11401
g8966 and n10983 n11401_not ; po0226
g8967 and pi0069 n11058 ; n11403
g8968 and n10153 n11403 ; n11404
g8969 nor pi0071 n11404 ; n11405
g8970 nor pi0081 pi0314 ; n11406
g8971 and n2465 n11406 ; n11407
g8972 and n6438 n11407 ; n11408
g8973 and n11405_not n11408 ; n11409
g8974 and pi0071 pi0314 ; n11410
g8975 and n7438 n11410 ; n11411
g8976 and n10150 n11411 ; n11412
g8977 and n2485 n11412 ; n11413
g8978 nor n11409 n11413 ; n11414
g8979 and n11107 n11414_not ; po0227
g8980 and n2505 n2749 ; n11416
g8981 and pi0096_not n11416 ; n11417
g8982 and n10194 n11417 ; n11418
g8983 and pi0198 pi0589 ; n11419
g8984 and n3471 n6207_not ; n11420
g8985 and n11419 n11420 ; n11421
g8986 and pi0210 pi0589 ; n11422
g8987 and pi0221_not n5853 ; n11423
g8988 and pi0216_not n11423 ; n11424
g8989 and n6244_not n11424 ; n11425
g8990 and n11422 n11425 ; n11426
g8991 nor n11421 n11426 ; n11427
g8992 and pi0593_not n6381 ; n11428
g8993 and n6389_not n11428 ; n11429
g8994 and n11427_not n11429 ; n11430
g8995 nor pi0287 n11430 ; n11431
g8996 and pi0039 n11431_not ; n11432
g8997 and n2521 n11432 ; n11433
g8998 nor n11418 n11433 ; n11434
g8999 and n10200 n11434_not ; po0228
g9000 and n2469 n2481 ; n11436
g9001 and n6424 n11436 ; n11437
g9002 and n11014 n11437 ; n11438
g9003 and pi0064_not n8916 ; n11439
g9004 and n11438 n11439 ; n11440
g9005 nor pi0081 n11440 ; n11441
g9006 and pi0050_not n8935 ; n11442
g9007 and n6444 n11442 ; n11443
g9008 and pi0199_not pi0200 ; n11444
g9009 and pi0299_not n11444 ; n11445
g9010 and pi0211 pi0219_not ; n11446
g9011 and pi0299 n11446 ; n11447
g9012 nor n11445 n11447 ; n11448
g9013 and pi0314 n11448_not ; n11449
g9014 and n10162 n11449 ; n11450
g9015 and n11441_not n11450 ; n11451
g9016 and n11443 n11451 ; n11452
g9017 and n11012 n11448 ; n11453
g9018 and n11376 n11453 ; n11454
g9019 and n11438 n11454 ; n11455
g9020 nor n11452 n11455 ; n11456
g9021 and n10165 n11456_not ; po0229
g9022 and pi0024 n2709 ; n11458
g9023 and pi0072 n11458 ; n11459
g9024 and pi0088 n10147 ; n11460
g9025 and n6388 n9141 ; n11461
g9026 and n11460 n11461 ; n11462
g9027 and n2870 n11462 ; n11463
g9028 nor n11459 n11463 ; n11464
g9029 and n6479 n11464_not ; n11465
g9030 nor pi0039 n11465 ; n11466
g9031 and n7604 n11395 ; n11467
g9032 and n7608 n11398 ; n11468
g9033 and pi0039 n11467_not ; n11469
g9034 and n11468_not n11469 ; n11470
g9035 and n10200 n11470_not ; n11471
g9036 and n11466_not n11471 ; po0230
g9037 and pi0314_not pi1050 ; n11473
g9038 and n9090 n10162 ; n11474
g9039 and n11473 n11474 ; n11475
g9040 nor pi0039 n11475 ; n11476
g9041 and n9051 n11398 ; n11477
g9042 nor pi0299 n11477 ; n11478
g9043 and n9036 n11395 ; n11479
g9044 and pi0299 n11479_not ; n11480
g9045 nor n11478 n11480 ; n11481
g9046 and pi0039 n11481_not ; n11482
g9047 and n10200 n11476_not ; n11483
g9048 and n11482_not n11483 ; po0231
g9049 and pi0074 n11293 ; n11485
g9050 and n2964 n7526 ; n11486
g9051 nor pi0096 n11486 ; n11487
g9052 nor pi0096 pi1093 ; n11488
g9053 and n7417 n11488 ; n11489
g9054 nor pi0096 n6169 ; n11490
g9055 and pi0479 n11490_not ; n11491
g9056 and n3373 n7429 ; n11492
g9057 and n11489_not n11492 ; n11493
g9058 nor po0840 n11491 ; n11494
g9059 and n11493 n11494 ; n11495
g9060 and n11487_not n11495 ; n11496
g9061 and n7456 n11496 ; n11497
g9062 nor n11485 n11497 ; n11498
g9063 nor po1038 n11498 ; po0232
g9064 and n2620 n10195 ; n11500
g9065 and pi0075 n11500_not ; n11501
g9066 and pi0096 pi1093_not ; n11502
g9067 and n2931 n11487_not ; n11503
g9068 nor n11502 n11503 ; n11504
g9069 and n2610 n11504_not ; n11505
g9070 and n7534 n11505 ; n11506
g9071 nor pi0075 n11506 ; n11507
g9072 and n8881 n11501_not ; n11508
g9073 and n11507_not n11508 ; po0233
g9074 and n8930 n10186 ; n11510
g9075 and n10111_not n11510 ; n11511
g9076 and po1057 n11511_not ; n11512
g9077 and n2519 n10375 ; n11513
g9078 and pi0252 n2933 ; n11514
g9079 and n11513 n11514_not ; n11515
g9080 and pi0137_not n11515 ; n11516
g9081 and pi0137_not n2924 ; n11517
g9082 nor pi0094 n8931 ; n11518
g9083 nor n8897 n10374 ; n11519
g9084 and n10162 n11518_not ; n11520
g9085 and n11519_not n11520 ; n11521
g9086 nor n2933 n11521 ; n11522
g9087 and pi0252_not n11521 ; n11523
g9088 and pi0252 n11510 ; n11524
g9089 and n2933 n11524_not ; n11525
g9090 and n11523_not n11525 ; n11526
g9091 nor n11522 n11526 ; n11527
g9092 and pi0122 n11527_not ; n11528
g9093 and n7417 n11522 ; n11529
g9094 nor n6277 n11513 ; n11530
g9095 nor n11526 n11530 ; n11531
g9096 and n11529_not n11531 ; n11532
g9097 nor pi0122 n11532 ; n11533
g9098 nor n11528 n11533 ; n11534
g9099 nor pi1093 n11534 ; n11535
g9100 nor pi0122 n11515 ; n11536
g9101 nor n11528 n11536 ; n11537
g9102 and pi1093 n11537_not ; n11538
g9103 nor n11535 n11538 ; n11539
g9104 and n2924 n11539_not ; n11540
g9105 nor n11517 n11540 ; n11541
g9106 nor n11516 n11541 ; n11542
g9107 and pi0122_not n11513 ; n11543
g9108 and pi1093 n11521_not ; n11544
g9109 nor n7418 n11544 ; n11545
g9110 nor n11543 n11545 ; n11546
g9111 nor n11535 n11546 ; n11547
g9112 nor n2924 n11547 ; n11548
g9113 nor pi0137 n2924 ; n11549
g9114 nor n11548 n11549 ; n11550
g9115 and pi0252 pi1092 ; n11551
g9116 and pi1093_not n11551 ; n11552
g9117 and n2925 n11552 ; n11553
g9118 nor pi0137 n11553 ; n11554
g9119 and n11513 n11554 ; n11555
g9120 nor n11550 n11555 ; n11556
g9121 nor n11542 n11556 ; n11557
g9122 nor po1057 n11557 ; n11558
g9123 and pi0137_not po1057 ; n11559
g9124 nor n11512 n11559 ; n11560
g9125 and n11558_not n11560 ; n11561
g9126 nor pi0210 n11561 ; n11562
g9127 nor n11540 n11548 ; n11563
g9128 nor po1057 n11563 ; n11564
g9129 nor n11512 n11564 ; n11565
g9130 and pi0210 n11565_not ; n11566
g9131 nor n11562 n11566 ; n11567
g9132 and n2638 n10299 ; n11568
g9133 nor n11567 n11568 ; n11569
g9134 nor pi0210 n11557 ; n11570
g9135 and pi0210 n11563_not ; n11571
g9136 nor n11570 n11571 ; n11572
g9137 and n11568 n11572_not ; n11573
g9138 and pi0299 n11573_not ; n11574
g9139 and n11569_not n11574 ; n11575
g9140 nor pi0198 n11561 ; n11576
g9141 and pi0198 n11565_not ; n11577
g9142 nor n11576 n11577 ; n11578
g9143 and n2669 n6197 ; n11579
g9144 nor n11578 n11579 ; n11580
g9145 and pi0198 n11563_not ; n11581
g9146 nor pi0198 n11557 ; n11582
g9147 nor n11581 n11582 ; n11583
g9148 and n11579 n11583_not ; n11584
g9149 nor pi0299 n11584 ; n11585
g9150 and n11580_not n11585 ; n11586
g9151 nor n11575 n11586 ; n11587
g9152 and pi0232 n11587_not ; n11588
g9153 and pi0299 n11567_not ; n11589
g9154 nor pi0299 n11578 ; n11590
g9155 nor pi0232 n11589 ; n11591
g9156 and n11590_not n11591 ; n11592
g9157 nor n11588 n11592 ; n11593
g9158 and n7425 n11593_not ; n11594
g9159 and n2924_not n11544 ; n11595
g9160 and n2933 n11513_not ; n11596
g9161 nor n11514 n11522 ; n11597
g9162 and n11596_not n11597 ; n11598
g9163 and n7418 n11598_not ; n11599
g9164 nor n11528 n11599 ; n11600
g9165 and n2924 n11600_not ; n11601
g9166 nor pi1093 n11527 ; n11602
g9167 nor n11595 n11602 ; n11603
g9168 and n11601_not n11603 ; n11604
g9169 and po1057_not n11604 ; n11605
g9170 and po1057 n11510 ; n11606
g9171 and n10108_not n11606 ; n11607
g9172 nor n11605 n11607 ; n11608
g9173 and pi0210 n11608_not ; n11609
g9174 and n8904 n11559 ; n11610
g9175 and pi0137 n11602 ; n11611
g9176 nor pi0137 n11598 ; n11612
g9177 and pi1093_not n11612 ; n11613
g9178 nor n11544 n11611 ; n11614
g9179 and n11613_not n11614 ; n11615
g9180 and po1057_not n11615 ; n11616
g9181 nor n11606 n11616 ; n11617
g9182 nor n2924 n11610 ; n11618
g9183 and n11617_not n11618 ; n11619
g9184 and pi0137 n7418_not ; n11620
g9185 and n2933 n11620_not ; n11621
g9186 and n11510 n11621_not ; n11622
g9187 and po1057 n11622_not ; n11623
g9188 and pi0137 n11600_not ; n11624
g9189 nor n11611 n11612 ; n11625
g9190 and n11624_not n11625 ; n11626
g9191 nor po1057 n11626 ; n11627
g9192 and n2924 n11623_not ; n11628
g9193 and n11627_not n11628 ; n11629
g9194 nor n11619 n11629 ; n11630
g9195 nor pi0210 n11630 ; n11631
g9196 nor n11609 n11631 ; n11632
g9197 nor n11568 n11632 ; n11633
g9198 and n2924_not n11615 ; n11634
g9199 and n2924 n11626 ; n11635
g9200 nor n11634 n11635 ; n11636
g9201 and pi0210_not n11636 ; n11637
g9202 and pi0210 n11604_not ; n11638
g9203 and n11568 n11638_not ; n11639
g9204 and n11637_not n11639 ; n11640
g9205 and pi0299 n11640_not ; n11641
g9206 and n11633_not n11641 ; n11642
g9207 and pi0198 n11608_not ; n11643
g9208 nor pi0198 n11630 ; n11644
g9209 nor n11643 n11644 ; n11645
g9210 nor n11579 n11645 ; n11646
g9211 nor pi0198 n11636 ; n11647
g9212 and pi0198 n11604 ; n11648
g9213 nor n11647 n11648 ; n11649
g9214 and n11579 n11649_not ; n11650
g9215 nor pi0299 n11650 ; n11651
g9216 and n11646_not n11651 ; n11652
g9217 nor n11642 n11652 ; n11653
g9218 and pi0232 n11653_not ; n11654
g9219 nor pi0299 n11645 ; n11655
g9220 and pi0299 n11632_not ; n11656
g9221 nor pi0232 n11655 ; n11657
g9222 and n11656_not n11657 ; n11658
g9223 nor n7425 n11658 ; n11659
g9224 and n11654_not n11659 ; n11660
g9225 nor n11594 n11660 ; n11661
g9226 and n10165 n11661_not ; po0234
g9227 and pi0086 n8897 ; n11663
g9228 and n2778 n11663 ; n11664
g9229 and pi0314 n11664_not ; n11665
g9230 and n2769 n2784 ; n11666
g9231 nor pi0086 n11666 ; n11667
g9232 and n6452 n11667_not ; n11668
g9233 and n2702 n11668 ; n11669
g9234 nor pi0314 n11669 ; n11670
g9235 and n10166 n11665_not ; n11671
g9236 and n11670_not n11671 ; po0235
g9237 and pi0119 pi0232 ; n11673
g9238 and pi0468_not n11673 ; po0236
g9239 and pi0163 n9700_not ; n11675
g9240 nor pi0163 n9696 ; n11676
g9241 and n9698_not n11676 ; n11677
g9242 nor n11675 n11677 ; n11678
g9243 and pi0232 n11678 ; n11679
g9244 and n8989_not n11679 ; n11680
g9245 and pi0074 n11680_not ; n11681
g9246 and pi0075 n11679_not ; n11682
g9247 and pi0100 n11679_not ; n11683
g9248 nor n11682 n11683 ; n11684
g9249 and pi0147 n7473 ; n11685
g9250 and n8989 n11685 ; n11686
g9251 and n11684 n11686_not ; n11687
g9252 nor n3328 n11681 ; n11688
g9253 and n11687 n11688 ; n11689
g9254 and pi0054 n11687_not ; n11690
g9255 nor pi0038 pi0040 ; n11691
g9256 and pi0038 n11685_not ; n11692
g9257 nor pi0100 n11692 ; n11693
g9258 and n11691_not n11693 ; n11694
g9259 nor n11683 n11694 ; n11695
g9260 nor pi0075 n11695 ; n11696
g9261 nor n11682 n11696 ; n11697
g9262 nor pi0054 n11697 ; n11698
g9263 nor n11690 n11698 ; n11699
g9264 nor pi0074 n11699 ; n11700
g9265 nor n11681 n11700 ; n11701
g9266 nor n2529 n11701 ; n11702
g9267 and n3328 n11702_not ; n11703
g9268 and n9722_not n9724 ; n11704
g9269 and pi0184_not n11704 ; n11705
g9270 and pi0184 n6197 ; n11706
g9271 and n11704_not n11706 ; n11707
g9272 nor pi0299 n11705 ; n11708
g9273 and n11707_not n11708 ; n11709
g9274 and pi0299 n11678_not ; n11710
g9275 and pi0232 n11709_not ; n11711
g9276 and n11710_not n11711 ; n11712
g9277 and n8989_not n11712 ; n11713
g9278 and pi0074 n11713_not ; n11714
g9279 nor pi0055 n11714 ; n11715
g9280 nor pi0187 pi0299 ; n11716
g9281 and pi0147_not pi0299 ; n11717
g9282 nor n11716 n11717 ; n11718
g9283 and n7473 n11718 ; n11719
g9284 and n8989 n11719_not ; n11720
g9285 and pi0054 n11720_not ; n11721
g9286 and n11713_not n11721 ; n11722
g9287 and pi0075 n11712_not ; n11723
g9288 and pi0100 n11712_not ; n11724
g9289 and pi0038 n11719_not ; n11725
g9290 nor pi0100 n11725 ; n11726
g9291 nor pi0179 pi0299 ; n11727
g9292 and pi0156_not pi0299 ; n11728
g9293 nor n11727 n11728 ; n11729
g9294 and n7473 n11729 ; n11730
g9295 and n2518 n2609 ; n11731
g9296 and n11730 n11731 ; n11732
g9297 and n2509 n11732 ; n11733
g9298 and n11691 n11733_not ; n11734
g9299 and n11726 n11734_not ; n11735
g9300 nor n11724 n11735 ; n11736
g9301 and n9205 n11736_not ; n11737
g9302 nor pi0187 n9187 ; n11738
g9303 and pi0187 n9189_not ; n11739
g9304 and pi0147 n11739_not ; n11740
g9305 and n11738_not n11740 ; n11741
g9306 and pi0147_not pi0187 ; n11742
g9307 and n9194 n11742 ; n11743
g9308 nor n11741 n11743 ; n11744
g9309 and pi0038 n11744_not ; n11745
g9310 and n2509 n9093 ; n11746
g9311 and n6242_not n9036 ; n11747
g9312 and pi0156 n6188 ; n11748
g9313 and pi0166_not n9293 ; n11749
g9314 nor n11748 n11749 ; n11750
g9315 and n11747 n11750_not ; n11751
g9316 and n11746 n11751 ; n11752
g9317 and pi0040_not pi0299 ; n11753
g9318 and n11752_not n11753 ; n11754
g9319 and pi0189_not n9293 ; n11755
g9320 and pi0179 n6188 ; n11756
g9321 nor n11755 n11756 ; n11757
g9322 and n6205_not n9051 ; n11758
g9323 and n11757_not n11758 ; n11759
g9324 and n11746 n11759 ; n11760
g9325 nor pi0040 pi0299 ; n11761
g9326 and n11760_not n11761 ; n11762
g9327 and pi0039 n11754_not ; n11763
g9328 and n11762_not n11763 ; n11764
g9329 nor pi0175 pi0299 ; n11765
g9330 and pi0184 n9147 ; n11766
g9331 nor pi0184 n9143 ; n11767
g9332 nor pi0189 n11767 ; n11768
g9333 and n11766_not n11768 ; n11769
g9334 and pi0032_not pi0095 ; n11770
g9335 and pi0479_not n11770 ; n11771
g9336 and n2509 n11771 ; n11772
g9337 and pi0182 n11772 ; n11773
g9338 and pi0184 pi0189 ; n11774
g9339 and n9150_not n11774 ; n11775
g9340 nor n11773 n11775 ; n11776
g9341 and n11769_not n11776 ; n11777
g9342 and n6197 n11777_not ; n11778
g9343 nor pi0040 n11778 ; n11779
g9344 and n11765 n11779_not ; n11780
g9345 and n6197 n11772 ; n11781
g9346 and pi0153 n9093 ; n11782
g9347 and n9133 n11782 ; n11783
g9348 and n9143 n10299 ; n11784
g9349 nor pi0040 pi0163 ; n11785
g9350 and n11784_not n11785 ; n11786
g9351 and n11783_not n11786 ; n11787
g9352 and n11781_not n11787 ; n11788
g9353 and pi0040 n6197_not ; n11789
g9354 and pi0166 n6197 ; n11790
g9355 nor pi0040 n11772 ; n11791
g9356 and n9166 n11791 ; n11792
g9357 and n11790 n11792_not ; n11793
g9358 and n9162 n11791 ; n11794
g9359 and n10299 n11794_not ; n11795
g9360 nor pi0153 n11793 ; n11796
g9361 and n11795_not n11796 ; n11797
g9362 nor pi0210 n9120 ; n11798
g9363 and n9118_not n11791 ; n11799
g9364 and n11798_not n11799 ; n11800
g9365 and n10299 n11800_not ; n11801
g9366 and n9129_not n11792 ; n11802
g9367 and n11790 n11802_not ; n11803
g9368 and pi0153 n11803_not ; n11804
g9369 and n11801_not n11804 ; n11805
g9370 nor n11797 n11805 ; n11806
g9371 and pi0163 n11789_not ; n11807
g9372 and n11806_not n11807 ; n11808
g9373 and pi0160 n11808_not ; n11809
g9374 and pi0153 n9118 ; n11810
g9375 and n9162 n11810_not ; n11811
g9376 and n10299 n11811_not ; n11812
g9377 and pi0153 n9129 ; n11813
g9378 and n9166 n11813_not ; n11814
g9379 and n11790 n11814_not ; n11815
g9380 and pi0040_not pi0163 ; n11816
g9381 and n11815_not n11816 ; n11817
g9382 and n11812_not n11817 ; n11818
g9383 nor pi0160 n11787 ; n11819
g9384 and n11818_not n11819 ; n11820
g9385 nor n11809 n11820 ; n11821
g9386 and pi0299 n11788_not ; n11822
g9387 and n11821_not n11822 ; n11823
g9388 and n9121_not n11799 ; n11824
g9389 and n10295 n11824_not ; n11825
g9390 and pi0189 n6197 ; n11826
g9391 and n9130 n11791 ; n11827
g9392 and n11826 n11827_not ; n11828
g9393 and pi0182 pi0184 ; n11829
g9394 and n11789_not n11829 ; n11830
g9395 and n11828_not n11830 ; n11831
g9396 and n11825_not n11831 ; n11832
g9397 and pi0175 pi0299_not ; n11833
g9398 and pi0189 n9133_not ; n11834
g9399 nor pi0189 n9092 ; n11835
g9400 and n2518 n11834_not ; n11836
g9401 and n11835_not n11836 ; n11837
g9402 nor n11773 n11837 ; n11838
g9403 and n6197 n11838_not ; n11839
g9404 nor pi0184 n11839 ; n11840
g9405 and pi0189 n9131 ; n11841
g9406 and n9122_not n10295 ; n11842
g9407 and pi0182_not pi0184 ; n11843
g9408 and n11841_not n11843 ; n11844
g9409 and n11842_not n11844 ; n11845
g9410 nor n11840 n11845 ; n11846
g9411 nor pi0040 n11846 ; n11847
g9412 and n11832_not n11833 ; n11848
g9413 and n11847_not n11848 ; n11849
g9414 nor n11780 n11849 ; n11850
g9415 and n11823_not n11850 ; n11851
g9416 nor pi0039 n11851 ; n11852
g9417 and pi0232 n11764_not ; n11853
g9418 and n11852_not n11853 ; n11854
g9419 nor pi0040 pi0232 ; n11855
g9420 nor pi0038 n11855 ; n11856
g9421 and n11854_not n11856 ; n11857
g9422 nor n11745 n11857 ; n11858
g9423 and n2568 n11858_not ; n11859
g9424 and pi0087 n11691_not ; n11860
g9425 and n11726 n11860 ; n11861
g9426 nor n11724 n11861 ; n11862
g9427 and n11859_not n11862 ; n11863
g9428 and n2569 n11863_not ; n11864
g9429 nor n11723 n11737 ; n11865
g9430 and n11864_not n11865 ; n11866
g9431 nor pi0054 n11866 ; n11867
g9432 nor n11722 n11867 ; n11868
g9433 nor pi0074 n11868 ; n11869
g9434 and n11715 n11869_not ; n11870
g9435 and pi0055 n11681_not ; n11871
g9436 and pi0163 pi0232 ; n11872
g9437 and pi0092_not n2609 ; n11873
g9438 and n11872 n11873 ; n11874
g9439 and n11746 n11874 ; n11875
g9440 and n11691 n11875_not ; n11876
g9441 and pi0075_not n11693 ; n11877
g9442 and n11876_not n11877 ; n11878
g9443 and n11684 n11878_not ; n11879
g9444 nor pi0054 n11879 ; n11880
g9445 nor n11690 n11880 ; n11881
g9446 nor pi0074 n11881 ; n11882
g9447 and n11871 n11882_not ; n11883
g9448 and n2529 n11883_not ; n11884
g9449 and n11870_not n11884 ; n11885
g9450 and n11703 n11885_not ; n11886
g9451 nor n11689 n11886 ; n11887
g9452 and pi0079 n11887 ; n11888
g9453 and n2487 n9260_not ; n11889
g9454 nor pi0040 n11889 ; n11890
g9455 and n6197_not n9260 ; n11891
g9456 and n9248 n11891_not ; n11892
g9457 and n11872 n11892 ; n11893
g9458 and n11890 n11893_not ; n11894
g9459 nor pi0039 n11894 ; n11895
g9460 and pi0039 n9466_not ; n11896
g9461 and n9208 n11896_not ; n11897
g9462 and n11895_not n11897 ; n11898
g9463 and pi0087 n2487_not ; n11899
g9464 and n11691 n11899 ; n11900
g9465 and n11693 n11900_not ; n11901
g9466 and n11898_not n11901 ; n11902
g9467 nor n11683 n11902 ; n11903
g9468 and n2569 n11903_not ; n11904
g9469 and n9284_not n11695 ; n11905
g9470 and n9205 n11905_not ; n11906
g9471 nor n11682 n11906 ; n11907
g9472 and n11904_not n11907 ; n11908
g9473 nor pi0054 n11908 ; n11909
g9474 nor n11690 n11909 ; n11910
g9475 nor pi0074 n11910 ; n11911
g9476 and n11871 n11911_not ; n11912
g9477 and n11726 n11900_not ; n11913
g9478 and n2487 n11730 ; n11914
g9479 and n11890 n11914_not ; n11915
g9480 nor pi0039 n11915 ; n11916
g9481 and n11897 n11916_not ; n11917
g9482 and n11913 n11917_not ; n11918
g9483 nor n11724 n11918 ; n11919
g9484 and n9205 n11919_not ; n11920
g9485 and pi0087 n11913 ; n11921
g9486 nor pi0040 n9297 ; n11922
g9487 and n6242 n11922_not ; n11923
g9488 and n6227 n9466 ; n11924
g9489 and n2487 n9295_not ; n11925
g9490 nor pi0040 n11925 ; n11926
g9491 and n6227_not n11926 ; n11927
g9492 nor n11924 n11927 ; n11928
g9493 and n6242_not n11928 ; n11929
g9494 nor n11923 n11929 ; n11930
g9495 and n9291 n11930 ; n11931
g9496 and n6205 n11922_not ; n11932
g9497 and n6205_not n11928 ; n11933
g9498 nor n11932 n11933 ; n11934
g9499 and n9051 n11934_not ; n11935
g9500 nor n9051 n9466 ; n11936
g9501 nor pi0299 n11936 ; n11937
g9502 and n11935_not n11937 ; n11938
g9503 nor pi0232 n11931 ; n11939
g9504 and n11938_not n11939 ; n11940
g9505 nor pi0189 n11922 ; n11941
g9506 and n2487 n9311_not ; n11942
g9507 and n9140 n11942_not ; n11943
g9508 and n6198 n11926 ; n11944
g9509 nor n11924 n11944 ; n11945
g9510 and n11943_not n11945 ; n11946
g9511 and pi0189 n6205_not ; n11947
g9512 and n11946 n11947 ; n11948
g9513 nor n11941 n11948 ; n11949
g9514 and pi0179 n11949_not ; n11950
g9515 and pi0189 n11928_not ; n11951
g9516 and n9140 n9324 ; n11952
g9517 and n2487_not n9140 ; n11953
g9518 nor n11952 n11953 ; n11954
g9519 and n11945 n11954 ; n11955
g9520 nor pi0189 n11955 ; n11956
g9521 nor pi0179 n6205 ; n11957
g9522 and n11951_not n11957 ; n11958
g9523 and n11956_not n11958 ; n11959
g9524 nor n11932 n11959 ; n11960
g9525 and n11950_not n11960 ; n11961
g9526 and n9051 n11961_not ; n11962
g9527 nor n11936 n11962 ; n11963
g9528 nor pi0299 n11963 ; n11964
g9529 and n9036_not n9466 ; n11965
g9530 and pi0299 n11965_not ; n11966
g9531 nor pi0166 n6242 ; n11967
g9532 nor n11930 n11967 ; n11968
g9533 and n11955 n11967 ; n11969
g9534 and n9036 n11969_not ; n11970
g9535 and n11968_not n11970 ; n11971
g9536 and n11966 n11971_not ; n11972
g9537 nor n11964 n11972 ; n11973
g9538 and pi0156_not pi0232 ; n11974
g9539 and n11973_not n11974 ; n11975
g9540 and pi0166 n6242_not ; n11976
g9541 and n11946 n11976 ; n11977
g9542 nor n11922 n11976 ; n11978
g9543 and n9036 n11978_not ; n11979
g9544 and n11977_not n11979 ; n11980
g9545 and n11966 n11980_not ; n11981
g9546 nor n11964 n11981 ; n11982
g9547 and pi0156 pi0232 ; n11983
g9548 and n11982_not n11983 ; n11984
g9549 and pi0039 n11940_not ; n11985
g9550 and n11975_not n11985 ; n11986
g9551 and n11984_not n11986 ; n11987
g9552 nor n2442 n9485 ; n11988
g9553 and n9348 n9349_not ; n11989
g9554 nor n11988 n11989 ; n11990
g9555 nor pi0040 n9456 ; n11991
g9556 nor pi0095 n11991 ; n11992
g9557 nor n11990 n11992 ; n11993
g9558 and pi0299_not n11993 ; n11994
g9559 nor pi0040 n9581 ; n11995
g9560 nor pi0095 n11995 ; n11996
g9561 nor n11990 n11996 ; n11997
g9562 and pi0299 n11997 ; n11998
g9563 nor pi0232 n11994 ; n11999
g9564 and n11998_not n11999 ; n12000
g9565 and n6197_not n11993 ; n12001
g9566 nor pi0040 n9427 ; n12002
g9567 nor pi0095 n12002 ; n12003
g9568 nor pi0040 n9442 ; n12004
g9569 and pi0189 n12004 ; n12005
g9570 and n12003 n12005_not ; n12006
g9571 and pi0182_not n11990 ; n12007
g9572 and pi0182 n9485 ; n12008
g9573 and n6197 n12008_not ; n12009
g9574 and n12007_not n12009 ; n12010
g9575 and n12006_not n12010 ; n12011
g9576 and pi0184 n12011_not ; n12012
g9577 and pi0040_not n9403 ; n12013
g9578 nor pi0032 n12013 ; n12014
g9579 nor n9487 n12014 ; n12015
g9580 nor pi0095 n12015 ; n12016
g9581 nor n9485 n12016 ; n12017
g9582 nor pi0198 n12017 ; n12018
g9583 nor n9467 n12014 ; n12019
g9584 nor pi0095 n12019 ; n12020
g9585 nor n9485 n12020 ; n12021
g9586 and pi0198 n12021_not ; n12022
g9587 and n10295 n12018_not ; n12023
g9588 and n12022_not n12023 ; n12024
g9589 and n11826 n11991 ; n12025
g9590 and pi0182 pi0184_not ; n12026
g9591 and n12024_not n12026 ; n12027
g9592 and n12025_not n12027 ; n12028
g9593 nor n12012 n12028 ; n12029
g9594 and n11765 n12029_not ; n12030
g9595 and pi0095 pi0182_not ; n12031
g9596 nor pi0040 n9503 ; n12032
g9597 and pi0095_not pi0189 ; n12033
g9598 and n2487 n12033_not ; n12034
g9599 and n12032 n12034_not ; n12035
g9600 nor n12031 n12035 ; n12036
g9601 and n11706 n12036_not ; n12037
g9602 and n12007_not n12037 ; n12038
g9603 and n9560 n10295 ; n12039
g9604 nor pi0198 n9490 ; n12040
g9605 nor pi0095 n9479 ; n12041
g9606 nor n9485 n12041 ; n12042
g9607 and pi0198 n12042_not ; n12043
g9608 and n11826 n12040_not ; n12044
g9609 and n12043_not n12044 ; n12045
g9610 and pi0182 n12039_not ; n12046
g9611 and n12045_not n12046 ; n12047
g9612 nor n9489 n11990 ; n12048
g9613 nor pi0198 n12048 ; n12049
g9614 nor n11990 n12041 ; n12050
g9615 and pi0198 n12050_not ; n12051
g9616 and n11826 n12049_not ; n12052
g9617 and n12051_not n12052 ; n12053
g9618 nor pi0182 n12053 ; n12054
g9619 nor n12047 n12054 ; n12055
g9620 nor n9560 n12031 ; n12056
g9621 and n10295 n11990_not ; n12057
g9622 and n12056_not n12057 ; n12058
g9623 nor n12055 n12058 ; n12059
g9624 nor pi0184 n12059 ; n12060
g9625 and n11833 n12038_not ; n12061
g9626 and n12060_not n12061 ; n12062
g9627 nor n12030 n12062 ; n12063
g9628 nor n12001 n12063 ; n12064
g9629 and n6197_not n11997 ; n12065
g9630 nor pi0095 n12032 ; n12066
g9631 and pi0166 n12066_not ; n12067
g9632 nor n11474 n12066 ; n12068
g9633 and pi0153 n12067_not ; n12069
g9634 and n12068_not n12069 ; n12070
g9635 and pi0166 n12004 ; n12071
g9636 and n12003 n12071_not ; n12072
g9637 and pi0153_not n12072 ; n12073
g9638 and pi0160_not n6197 ; n12074
g9639 and n12070_not n12074 ; n12075
g9640 and n11990_not n12075 ; n12076
g9641 and n12073_not n12076 ; n12077
g9642 and n6197 n9485_not ; n12078
g9643 and n12067 n12078 ; n12079
g9644 and n9466 n10299 ; n12080
g9645 and pi0153 n12080_not ; n12081
g9646 and n12079_not n12081 ; n12082
g9647 and n12072_not n12078 ; n12083
g9648 nor pi0153 n12083 ; n12084
g9649 and pi0160 n12082_not ; n12085
g9650 and n12084_not n12085 ; n12086
g9651 and pi0163 n12077_not ; n12087
g9652 and n12086_not n12087 ; n12088
g9653 and pi0210 n12050_not ; n12089
g9654 nor pi0210 n12048 ; n12090
g9655 and n11790 n12089_not ; n12091
g9656 and n12090_not n12091 ; n12092
g9657 nor n9557 n11990 ; n12093
g9658 nor pi0210 n12093 ; n12094
g9659 nor n9553 n11990 ; n12095
g9660 and pi0210 n12095_not ; n12096
g9661 and n10299 n12094_not ; n12097
g9662 and n12096_not n12097 ; n12098
g9663 and pi0153 n12092_not ; n12099
g9664 and n12098_not n12099 ; n12100
g9665 and pi0166 n11997 ; n12101
g9666 nor n11990 n12020 ; n12102
g9667 and pi0210 n12102_not ; n12103
g9668 nor n11990 n12016 ; n12104
g9669 nor pi0210 n12104 ; n12105
g9670 and n10299 n12103_not ; n12106
g9671 and n12105_not n12106 ; n12107
g9672 nor pi0153 n12107 ; n12108
g9673 and n12101_not n12108 ; n12109
g9674 nor pi0160 n12100 ; n12110
g9675 and n12109_not n12110 ; n12111
g9676 and pi0210 n9554_not ; n12112
g9677 nor pi0210 n9558 ; n12113
g9678 and n10299 n12112_not ; n12114
g9679 and n12113_not n12114 ; n12115
g9680 nor pi0210 n9490 ; n12116
g9681 and pi0210 n12042_not ; n12117
g9682 and n11790 n12116_not ; n12118
g9683 and n12117_not n12118 ; n12119
g9684 and pi0153 n12115_not ; n12120
g9685 and n12119_not n12120 ; n12121
g9686 and n11790 n11995 ; n12122
g9687 nor pi0210 n12017 ; n12123
g9688 and pi0210 n12021_not ; n12124
g9689 and n10299 n12123_not ; n12125
g9690 and n12124_not n12125 ; n12126
g9691 nor pi0153 n12126 ; n12127
g9692 and n12122_not n12127 ; n12128
g9693 and pi0160 n12121_not ; n12129
g9694 and n12128_not n12129 ; n12130
g9695 nor pi0163 n12130 ; n12131
g9696 and n12111_not n12131 ; n12132
g9697 nor n12088 n12132 ; n12133
g9698 and pi0299 n12065_not ; n12134
g9699 and n12133_not n12134 ; n12135
g9700 and n10295_not n11993 ; n12136
g9701 and pi0198 n12102_not ; n12137
g9702 nor pi0198 n12104 ; n12138
g9703 and n10295 n12137_not ; n12139
g9704 and n12138_not n12139 ; n12140
g9705 nor pi0182 pi0184 ; n12141
g9706 and n11765 n12141 ; n12142
g9707 and n12140_not n12142 ; n12143
g9708 and n12136_not n12143 ; n12144
g9709 nor n12064 n12144 ; n12145
g9710 and n12135_not n12145 ; n12146
g9711 and pi0232 n12146_not ; n12147
g9712 nor pi0039 n12000 ; n12148
g9713 and n12147_not n12148 ; n12149
g9714 nor pi0038 n11987 ; n12150
g9715 and n12149_not n12150 ; n12151
g9716 nor n11745 n12151 ; n12152
g9717 and n2568 n12152_not ; n12153
g9718 nor n11724 n11921 ; n12154
g9719 and n12153_not n12154 ; n12155
g9720 and n2569 n12155_not ; n12156
g9721 nor n11723 n11920 ; n12157
g9722 and n12156_not n12157 ; n12158
g9723 nor pi0054 n12158 ; n12159
g9724 nor n11722 n12159 ; n12160
g9725 nor pi0074 n12160 ; n12161
g9726 and n11715 n12161_not ; n12162
g9727 and n2529 n11912_not ; n12163
g9728 and n12162_not n12163 ; n12164
g9729 and n9252_not n11703 ; n12165
g9730 and n12164_not n12165 ; n12166
g9731 nor n11689 n12166 ; n12167
g9732 and pi0079_not n12167 ; n12168
g9733 and pi0034_not n10058 ; n12169
g9734 nor n11888 n12169 ; n12170
g9735 and n12168_not n12170 ; n12171
g9736 nor pi0079 n8977 ; n12172
g9737 and n11887 n12172 ; n12173
g9738 and n12167 n12172_not ; n12174
g9739 and n12169 n12173_not ; n12175
g9740 and n12174_not n12175 ; n12176
g9741 or n12171 n12176 ; po0237
g9742 and pi0098 pi1092 ; n12178
g9743 and pi1093 n12178 ; n12179
g9744 and pi0567_not n2926 ; n12180
g9745 nor n12179 n12180 ; n12181
g9746 nor pi0080 n12181 ; n12182
g9747 and pi0217 n12182_not ; n12183
g9748 and n7425 n12181 ; n12184
g9749 and n8041_not n12181 ; n12185
g9750 and pi0588 n12185_not ; n12186
g9751 and pi0592 n8093_not ; n12187
g9752 and n7422 n8119_not ; n12188
g9753 and n12187_not n12188 ; n12189
g9754 and n12181 n12189_not ; n12190
g9755 nor pi1199 n12190 ; n12191
g9756 and pi0428 n12190_not ; n12192
g9757 and n7644_not n12181 ; n12193
g9758 nor pi0428 n12193 ; n12194
g9759 nor n12192 n12194 ; n12195
g9760 nor pi0427 n12195 ; n12196
g9761 nor pi0428 n12190 ; n12197
g9762 and pi0428 n12193_not ; n12198
g9763 nor n12197 n12198 ; n12199
g9764 and pi0427 n12199_not ; n12200
g9765 nor n12196 n12200 ; n12201
g9766 nor pi0430 n12201 ; n12202
g9767 nor pi0427 n12199 ; n12203
g9768 and pi0427 n12195_not ; n12204
g9769 nor n12203 n12204 ; n12205
g9770 and pi0430 n12205_not ; n12206
g9771 nor n12202 n12206 ; n12207
g9772 nor pi0426 n12207 ; n12208
g9773 nor pi0430 n12205 ; n12209
g9774 and pi0430 n12201_not ; n12210
g9775 nor n12209 n12210 ; n12211
g9776 and pi0426 n12211_not ; n12212
g9777 nor n12208 n12212 ; n12213
g9778 nor pi0445 n12213 ; n12214
g9779 nor pi0426 n12211 ; n12215
g9780 and pi0426 n12207_not ; n12216
g9781 nor n12215 n12216 ; n12217
g9782 and pi0445 n12217_not ; n12218
g9783 nor n12214 n12218 ; n12219
g9784 and pi0448 n12219_not ; n12220
g9785 nor pi0445 n12217 ; n12221
g9786 and pi0445 n12213_not ; n12222
g9787 nor n12221 n12222 ; n12223
g9788 nor pi0448 n12223 ; n12224
g9789 and n8128 n12220_not ; n12225
g9790 and n12224_not n12225 ; n12226
g9791 nor pi0448 n12219 ; n12227
g9792 and pi0448 n12223_not ; n12228
g9793 nor n8128 n12227 ; n12229
g9794 and n12228_not n12229 ; n12230
g9795 and pi1199 n12226_not ; n12231
g9796 and n12230_not n12231 ; n12232
g9797 and n8041 n12191_not ; n12233
g9798 and n12232_not n12233 ; n12234
g9799 and n12186 n12234_not ; n12235
g9800 and pi0591 n12181_not ; n12236
g9801 and pi0590 n12236_not ; n12237
g9802 and n7645_not n12181 ; n12238
g9803 and n7854 n12238 ; n12239
g9804 and n7757_not n12239 ; n12240
g9805 nor n12193 n12240 ; n12241
g9806 and pi0461 n12241_not ; n12242
g9807 and n7862_not n12239 ; n12243
g9808 nor n12193 n12243 ; n12244
g9809 nor pi0461 n12244 ; n12245
g9810 nor n12242 n12245 ; n12246
g9811 and pi0357 n12246_not ; n12247
g9812 and pi0461 n12244_not ; n12248
g9813 nor pi0461 n12241 ; n12249
g9814 nor n12248 n12249 ; n12250
g9815 nor pi0357 n12250 ; n12251
g9816 nor n12247 n12251 ; n12252
g9817 and pi0356 n12252_not ; n12253
g9818 and pi0357 n12250_not ; n12254
g9819 nor pi0357 n12246 ; n12255
g9820 nor n12254 n12255 ; n12256
g9821 nor pi0356 n12256 ; n12257
g9822 nor n12253 n12257 ; n12258
g9823 and pi0354 n12258 ; n12259
g9824 and pi0356 n12256_not ; n12260
g9825 nor pi0356 n12252 ; n12261
g9826 nor n12260 n12261 ; n12262
g9827 and pi0354_not n12262 ; n12263
g9828 nor n7887 n12259 ; n12264
g9829 and n12263_not n12264 ; n12265
g9830 and pi0354 n12262 ; n12266
g9831 and pi0354_not n12258 ; n12267
g9832 and n7887 n12266_not ; n12268
g9833 and n12267_not n12268 ; n12269
g9834 nor pi0591 n12265 ; n12270
g9835 and n12269_not n12270 ; n12271
g9836 and n12237 n12271_not ; n12272
g9837 nor pi1197 n8395 ; n12273
g9838 nor n12193 n12273 ; n12274
g9839 and pi0592 n12181_not ; n12275
g9840 nor pi1196 n12181 ; n12276
g9841 nor n12275 n12276 ; n12277
g9842 and pi0397 pi0404_not ; n12278
g9843 and pi0397_not pi0404 ; n12279
g9844 nor n12278 n12279 ; n12280
g9845 and pi0411 n12280_not ; n12281
g9846 and pi0411_not n12280 ; n12282
g9847 nor n12281 n12282 ; n12283
g9848 and n7932_not n12283 ; n12284
g9849 and n7932 n12283_not ; n12285
g9850 nor n12284 n12285 ; n12286
g9851 and n7417 n12286_not ; n12287
g9852 nor n12178 n12287 ; n12288
g9853 nor pi0412 n12288 ; n12289
g9854 and n7417 n12286 ; n12290
g9855 nor n12178 n12290 ; n12291
g9856 and pi0412 n12291_not ; n12292
g9857 and n7944 n12289_not ; n12293
g9858 and n12292_not n12293 ; n12294
g9859 and pi0412 n12288_not ; n12295
g9860 nor pi0412 n12291 ; n12296
g9861 nor n7944 n12295 ; n12297
g9862 and n12296_not n12297 ; n12298
g9863 nor pi0122 n12294 ; n12299
g9864 and n12298_not n12299 ; n12300
g9865 nor n12178 n12300 ; n12301
g9866 and n7626 n12301_not ; n12302
g9867 and pi1091 n12179 ; n12303
g9868 nor n12302 n12303 ; n12304
g9869 and pi0567 n12304_not ; n12305
g9870 nor n12180 n12305 ; n12306
g9871 and n7958 n12306_not ; n12307
g9872 and n12277 n12307_not ; n12308
g9873 nor pi1199 n12308 ; n12309
g9874 and pi0122_not n7417 ; n12310
g9875 nor n12178 n12310 ; n12311
g9876 nor n7626 n12303 ; n12312
g9877 and n7417 n7926 ; n12313
g9878 nor pi0122 n12178 ; n12314
g9879 and n12313_not n12314 ; n12315
g9880 nor n12312 n12315 ; n12316
g9881 and n12311_not n12316 ; n12317
g9882 and pi0567 n12317 ; n12318
g9883 nor n12180 n12318 ; n12319
g9884 and n12305_not n12319 ; n12320
g9885 and n7958 n12320_not ; n12321
g9886 and n8668 n12319_not ; n12322
g9887 nor n12275 n12322 ; n12323
g9888 and n12321_not n12323 ; n12324
g9889 and pi1199 n12324_not ; n12325
g9890 nor n12309 n12325 ; n12326
g9891 and n12273 n12326_not ; n12327
g9892 nor n12274 n12327 ; n12328
g9893 and pi0333 n12328_not ; n12329
g9894 and n8395 n12193_not ; n12330
g9895 nor n8395 n12326 ; n12331
g9896 nor n12330 n12331 ; n12332
g9897 nor pi0333 n12332 ; n12333
g9898 nor n12329 n12333 ; n12334
g9899 and pi0391 n12334_not ; n12335
g9900 nor pi0333 n12328 ; n12336
g9901 and pi0333 n12332_not ; n12337
g9902 nor n12336 n12337 ; n12338
g9903 nor pi0391 n12338 ; n12339
g9904 and pi0392 n8801 ; n12340
g9905 nor pi0392 n8801 ; n12341
g9906 nor n12340 n12341 ; n12342
g9907 nor n12335 n12342 ; n12343
g9908 and n12339_not n12343 ; n12344
g9909 and pi0391 n12338_not ; n12345
g9910 nor pi0391 n12334 ; n12346
g9911 and n12342 n12345_not ; n12347
g9912 and n12346_not n12347 ; n12348
g9913 and pi0591 n12344_not ; n12349
g9914 and n12348_not n12349 ; n12350
g9915 nor n7644 n7755 ; n12351
g9916 and n7422 n7726_not ; n12352
g9917 nor pi1198 n12352 ; n12353
g9918 nor n7970 n12353 ; n12354
g9919 and n12351_not n12354 ; n12355
g9920 and n12181 n12355_not ; n12356
g9921 nor pi0591 n12356 ; n12357
g9922 nor pi0590 n12357 ; n12358
g9923 and n12350_not n12358 ; n12359
g9924 nor pi0588 n12272 ; n12360
g9925 and n12359_not n12360 ; n12361
g9926 nor n7425 n12235 ; n12362
g9927 and n12361_not n12362 ; n12363
g9928 and pi0080_not po1038 ; n12364
g9929 and n12184_not n12364 ; n12365
g9930 and n12363_not n12365 ; n12366
g9931 and pi0567 n7429 ; n12367
g9932 nor n7420 n12179 ; n12368
g9933 and pi0122_not n12368 ; n12369
g9934 and n7626 n12369_not ; n12370
g9935 and n2625 n12303_not ; n12371
g9936 and n12370_not n12371 ; n12372
g9937 and pi0824 pi0950 ; n12373
g9938 and pi0110_not n2701 ; n12374
g9939 and pi0088_not n2495 ; n12375
g9940 and n10379 n12375 ; n12376
g9941 and n12374 n12376 ; n12377
g9942 and n7440 n12377 ; n12378
g9943 and n7446 n12378 ; n12379
g9944 and pi0051 n12379 ; n12380
g9945 and pi0090 pi0093 ; n12381
g9946 nor pi0841 n2704 ; n12382
g9947 and n12381_not n12382 ; n12383
g9948 and n2962 n12383 ; n12384
g9949 and n12378 n12384 ; n12385
g9950 nor n12380 n12385 ; n12386
g9951 and n7450 n12373 ; n12387
g9952 and n12386_not n12387 ; n12388
g9953 nor pi0098 n12388 ; n12389
g9954 and pi1092 n12389_not ; n12390
g9955 and pi0087_not n12371 ; n12391
g9956 and n12390_not n12391 ; n12392
g9957 and n2520 n12373 ; n12393
g9958 and n12379 n12393 ; n12394
g9959 nor pi0098 n12394 ; n12395
g9960 and pi1092 n12395_not ; n12396
g9961 and pi0087 n12371 ; n12397
g9962 and n12396_not n12397 ; n12398
g9963 nor n12392 n12398 ; n12399
g9964 and pi0122 n12399_not ; n12400
g9965 nor n12372 n12400 ; n12401
g9966 nor pi0075 n12401 ; n12402
g9967 and n7465_not n12368 ; n12403
g9968 and n12367 n12403_not ; n12404
g9969 and n12402_not n12404 ; n12405
g9970 nor n7429 n12368 ; n12406
g9971 nor n12180 n12406 ; n12407
g9972 and n12405_not n12407 ; n12408
g9973 nor pi0592 n12408 ; n12409
g9974 nor n12275 n12409 ; n12410
g9975 and n8093_not n12410 ; n12411
g9976 and n8093 n12276_not ; n12412
g9977 nor pi0443 n12181 ; n12413
g9978 and pi0443 n12410_not ; n12414
g9979 nor n12413 n12414 ; n12415
g9980 and n8249 n12415 ; n12416
g9981 and pi0443 n12181_not ; n12417
g9982 nor pi0443 n12410 ; n12418
g9983 nor n12417 n12418 ; n12419
g9984 and n8249_not n12419 ; n12420
g9985 nor n12416 n12420 ; n12421
g9986 and pi0435 n12421_not ; n12422
g9987 and pi0444_not n12419 ; n12423
g9988 and pi0444 n12415 ; n12424
g9989 nor pi0436 n12423 ; n12425
g9990 and n12424_not n12425 ; n12426
g9991 and pi0444_not n12415 ; n12427
g9992 and pi0444 n12419 ; n12428
g9993 and pi0436 n12427_not ; n12429
g9994 and n12428_not n12429 ; n12430
g9995 nor n12426 n12430 ; n12431
g9996 and pi0435_not n12431 ; n12432
g9997 nor n12422 n12432 ; n12433
g9998 and pi0429_not n12433 ; n12434
g9999 nor pi0435 n12421 ; n12435
g10000 and pi0435 n12431 ; n12436
g10001 nor n12435 n12436 ; n12437
g10002 and pi0429 n12437 ; n12438
g10003 and n8105 n12434_not ; n12439
g10004 and n12438_not n12439 ; n12440
g10005 and pi0429_not n12437 ; n12441
g10006 and pi0429 n12433 ; n12442
g10007 nor n8105 n12441 ; n12443
g10008 and n12442_not n12443 ; n12444
g10009 and pi1196 n12440_not ; n12445
g10010 and n12444_not n12445 ; n12446
g10011 and n12412 n12446_not ; n12447
g10012 nor n12411 n12447 ; n12448
g10013 and pi1199_not n12448 ; n12449
g10014 and pi0428 n12448_not ; n12450
g10015 and pi0428_not n12410 ; n12451
g10016 nor n12450 n12451 ; n12452
g10017 nor pi0427 n12452 ; n12453
g10018 nor pi0428 n12448 ; n12454
g10019 and pi0428 n12410 ; n12455
g10020 nor n12454 n12455 ; n12456
g10021 and pi0427 n12456_not ; n12457
g10022 nor n12453 n12457 ; n12458
g10023 and pi0430 n12458_not ; n12459
g10024 nor pi0427 n12456 ; n12460
g10025 and pi0427 n12452_not ; n12461
g10026 nor n12460 n12461 ; n12462
g10027 nor pi0430 n12462 ; n12463
g10028 nor n12459 n12463 ; n12464
g10029 and pi0426 n12464_not ; n12465
g10030 and pi0430 n12462_not ; n12466
g10031 nor pi0430 n12458 ; n12467
g10032 nor n12466 n12467 ; n12468
g10033 nor pi0426 n12468 ; n12469
g10034 nor n12465 n12469 ; n12470
g10035 and pi0445 n12470_not ; n12471
g10036 and pi0426 n12468_not ; n12472
g10037 nor pi0426 n12464 ; n12473
g10038 nor n12472 n12473 ; n12474
g10039 nor pi0445 n12474 ; n12475
g10040 nor n12471 n12475 ; n12476
g10041 and pi0448 n12476 ; n12477
g10042 and pi0445 n12474_not ; n12478
g10043 nor pi0445 n12470 ; n12479
g10044 nor n12478 n12479 ; n12480
g10045 and pi0448_not n12480 ; n12481
g10046 nor n8128 n12477 ; n12482
g10047 and n12481_not n12482 ; n12483
g10048 and pi0448_not n12476 ; n12484
g10049 and pi0448 n12480 ; n12485
g10050 and n8128 n12484_not ; n12486
g10051 and n12485_not n12486 ; n12487
g10052 and pi1199 n12483_not ; n12488
g10053 and n12487_not n12488 ; n12489
g10054 and n8041 n12449_not ; n12490
g10055 and n12489_not n12490 ; n12491
g10056 and n12186 n12491_not ; n12492
g10057 and n7850 n12181 ; n12493
g10058 and n7850_not n12410 ; n12494
g10059 nor n12493 n12494 ; n12495
g10060 and pi1198 n12495_not ; n12496
g10061 nor pi1198 n12276 ; n12497
g10062 and n7791 n12181 ; n12498
g10063 and n7791_not n12410 ; n12499
g10064 nor n12498 n12499 ; n12500
g10065 nor pi0355 n12500 ; n12501
g10066 and pi0455 n12181_not ; n12502
g10067 nor pi0455 n12410 ; n12503
g10068 nor n12502 n12503 ; n12504
g10069 nor pi0452 n12504 ; n12505
g10070 nor pi0455 n12181 ; n12506
g10071 and pi0455 n12410_not ; n12507
g10072 nor n12506 n12507 ; n12508
g10073 and pi0452 n12508_not ; n12509
g10074 nor n12505 n12509 ; n12510
g10075 and pi0355 n12510 ; n12511
g10076 nor n12501 n12511 ; n12512
g10077 and pi0458_not n12512 ; n12513
g10078 and pi0355 n12500_not ; n12514
g10079 and pi0355_not n12510 ; n12515
g10080 nor n12514 n12515 ; n12516
g10081 and pi0458 n12516 ; n12517
g10082 and n7812 n12513_not ; n12518
g10083 and n12517_not n12518 ; n12519
g10084 and pi0458_not n12516 ; n12520
g10085 and pi0458 n12512 ; n12521
g10086 nor n7812 n12520 ; n12522
g10087 and n12521_not n12522 ; n12523
g10088 and pi1196 n12519_not ; n12524
g10089 and n12523_not n12524 ; n12525
g10090 and n12497 n12525_not ; n12526
g10091 nor n12496 n12526 ; n12527
g10092 nor n7782 n12527 ; n12528
g10093 and n7782 n12410 ; n12529
g10094 nor n12528 n12529 ; n12530
g10095 and n7757_not n12530 ; n12531
g10096 and pi1199 n12410_not ; n12532
g10097 and pi0351 n12532 ; n12533
g10098 nor n12531 n12533 ; n12534
g10099 nor pi0461 n12534 ; n12535
g10100 and n7862_not n12530 ; n12536
g10101 and pi0351_not n12532 ; n12537
g10102 nor n12536 n12537 ; n12538
g10103 and pi0461 n12538_not ; n12539
g10104 nor n12535 n12539 ; n12540
g10105 nor pi0357 n12540 ; n12541
g10106 nor pi0461 n12538 ; n12542
g10107 and pi0461 n12534_not ; n12543
g10108 nor n12542 n12543 ; n12544
g10109 and pi0357 n12544_not ; n12545
g10110 nor n12541 n12545 ; n12546
g10111 nor pi0356 n12546 ; n12547
g10112 nor pi0357 n12544 ; n12548
g10113 and pi0357 n12540_not ; n12549
g10114 nor n12548 n12549 ; n12550
g10115 and pi0356 n12550_not ; n12551
g10116 nor n12547 n12551 ; n12552
g10117 nor pi0354 n12552 ; n12553
g10118 nor pi0356 n12550 ; n12554
g10119 and pi0356 n12546_not ; n12555
g10120 nor n12554 n12555 ; n12556
g10121 and pi0354 n12556_not ; n12557
g10122 nor n7887 n12553 ; n12558
g10123 and n12557_not n12558 ; n12559
g10124 nor pi0354 n12556 ; n12560
g10125 and pi0354 n12552_not ; n12561
g10126 and n7887 n12560_not ; n12562
g10127 and n12561_not n12562 ; n12563
g10128 nor pi0591 n12559 ; n12564
g10129 and n12563_not n12564 ; n12565
g10130 and n12237 n12565_not ; n12566
g10131 and n12273_not n12410 ; n12567
g10132 and n7429 n12180_not ; n12568
g10133 nor n12306 n12568 ; n12569
g10134 and pi0075 n12304 ; n12570
g10135 and pi0411_not n12178 ; n12571
g10136 and n7950 n12571_not ; n12572
g10137 and pi0411 n12396 ; n12573
g10138 and n12572 n12573_not ; n12574
g10139 and pi0411_not n12396 ; n12575
g10140 nor n7950 n12178 ; n12576
g10141 nor n7952 n12576 ; n12577
g10142 nor n12575 n12577 ; n12578
g10143 nor n12574 n12578 ; n12579
g10144 and pi0122 n12579 ; n12580
g10145 nor n12300 n12580 ; n12581
g10146 and n7626 n12581_not ; n12582
g10147 and n12397 n12582_not ; n12583
g10148 and pi0411 n12390 ; n12584
g10149 and n12572 n12584_not ; n12585
g10150 and pi0411_not n12390 ; n12586
g10151 nor n12577 n12586 ; n12587
g10152 nor n12585 n12587 ; n12588
g10153 and pi0122 n12588 ; n12589
g10154 nor n12300 n12589 ; n12590
g10155 and n7626 n12590_not ; n12591
g10156 and n12391 n12591_not ; n12592
g10157 and n2625_not n12304 ; n12593
g10158 nor n12583 n12593 ; n12594
g10159 and n12592_not n12594 ; n12595
g10160 nor pi0075 n12595 ; n12596
g10161 and n12367 n12570_not ; n12597
g10162 and n12596_not n12597 ; n12598
g10163 nor n12569 n12598 ; n12599
g10164 and n7958 n12599_not ; n12600
g10165 nor n12276 n12600 ; n12601
g10166 nor pi1199 n12601 ; n12602
g10167 nor n12320 n12568 ; n12603
g10168 nor n7465 n12317 ; n12604
g10169 and n12302_not n12604 ; n12605
g10170 and n2625 n12316_not ; n12606
g10171 and n12302_not n12606 ; n12607
g10172 and pi0122_not n12313 ; n12608
g10173 and n7926 n12390 ; n12609
g10174 and n7926_not n12178 ; n12610
g10175 nor n12609 n12610 ; n12611
g10176 and n12391 n12611 ; n12612
g10177 nor n7950 n12586 ; n12613
g10178 nor n12585 n12613 ; n12614
g10179 and n12612 n12614_not ; n12615
g10180 and n7926 n12396 ; n12616
g10181 and n12397 n12616_not ; n12617
g10182 and n12579_not n12617 ; n12618
g10183 nor n12615 n12618 ; n12619
g10184 nor n12300 n12608 ; n12620
g10185 and n12619_not n12620 ; n12621
g10186 nor n12607 n12621 ; n12622
g10187 nor pi0075 n12622 ; n12623
g10188 and n12367 n12605_not ; n12624
g10189 and n12623_not n12624 ; n12625
g10190 nor n12603 n12625 ; n12626
g10191 and n7958 n12626_not ; n12627
g10192 nor n12319 n12568 ; n12628
g10193 nor n12610 n12616 ; n12629
g10194 and n12397 n12629 ; n12630
g10195 nor n12612 n12630 ; n12631
g10196 and pi0122 n12631_not ; n12632
g10197 nor n12606 n12632 ; n12633
g10198 nor pi0075 n12633 ; n12634
g10199 and n12367 n12604_not ; n12635
g10200 and n12634_not n12635 ; n12636
g10201 nor n12628 n12636 ; n12637
g10202 and n8668 n12637_not ; n12638
g10203 nor n12627 n12638 ; n12639
g10204 and pi1199 n12639_not ; n12640
g10205 nor n12275 n12640 ; n12641
g10206 and n12602_not n12641 ; n12642
g10207 and n12273 n12642 ; n12643
g10208 nor n12567 n12643 ; n12644
g10209 and pi0333 n12644_not ; n12645
g10210 and n8395 n12410_not ; n12646
g10211 nor n8395 n12642 ; n12647
g10212 nor n12646 n12647 ; n12648
g10213 and pi0333_not n12648 ; n12649
g10214 nor n12645 n12649 ; n12650
g10215 and pi0391 n12650_not ; n12651
g10216 and pi0333 n12648_not ; n12652
g10217 and pi0333_not n12644 ; n12653
g10218 nor n12652 n12653 ; n12654
g10219 and pi0391_not n12654 ; n12655
g10220 nor n12651 n12655 ; n12656
g10221 and pi0392 n12656_not ; n12657
g10222 and pi0391_not n12650 ; n12658
g10223 and pi0391 n12654_not ; n12659
g10224 nor n12658 n12659 ; n12660
g10225 and pi0392_not n12660 ; n12661
g10226 nor n12657 n12661 ; n12662
g10227 and pi0393 n12662_not ; n12663
g10228 nor pi0392 n12656 ; n12664
g10229 and pi0392 n12660 ; n12665
g10230 nor n12664 n12665 ; n12666
g10231 nor pi0393 n12666 ; n12667
g10232 nor n12663 n12667 ; n12668
g10233 nor n8028 n12668 ; n12669
g10234 and pi0393 n12666_not ; n12670
g10235 nor pi0393 n12662 ; n12671
g10236 nor n12670 n12671 ; n12672
g10237 and n8028 n12672_not ; n12673
g10238 and pi0591 n12669_not ; n12674
g10239 and n12673_not n12674 ; n12675
g10240 nor pi0592 n12181 ; n12676
g10241 and pi0592 n12408_not ; n12677
g10242 nor n12676 n12677 ; n12678
g10243 and n7722_not n12678 ; n12679
g10244 and n7722 n12181 ; n12680
g10245 nor n12679 n12680 ; n12681
g10246 and pi1199 n12681 ; n12682
g10247 and n7670 n12678 ; n12683
g10248 nor pi1197 n12181 ; n12684
g10249 nor n7670 n12684 ; n12685
g10250 and pi0367 n12181_not ; n12686
g10251 nor pi0367 n12678 ; n12687
g10252 nor n12686 n12687 ; n12688
g10253 and n7673 n12688_not ; n12689
g10254 nor pi0367 n12181 ; n12690
g10255 and pi0367 n12678_not ; n12691
g10256 nor n12690 n12691 ; n12692
g10257 nor n7673 n12692 ; n12693
g10258 nor n12689 n12693 ; n12694
g10259 and n7676 n12694_not ; n12695
g10260 and n7673_not n12688 ; n12696
g10261 and n7673 n12692 ; n12697
g10262 nor n12696 n12697 ; n12698
g10263 and n7676_not n12698 ; n12699
g10264 nor n7685 n12695 ; n12700
g10265 and n12699_not n12700 ; n12701
g10266 nor n7676 n12694 ; n12702
g10267 and n7676 n12698 ; n12703
g10268 and n7685 n12702_not ; n12704
g10269 and n12703_not n12704 ; n12705
g10270 and pi1197 n12701_not ; n12706
g10271 and n12705_not n12706 ; n12707
g10272 and n12685 n12707_not ; n12708
g10273 nor pi1199 n12683 ; n12709
g10274 and n12708_not n12709 ; n12710
g10275 nor n12682 n12710 ; n12711
g10276 nor pi0374 n12711 ; n12712
g10277 and n8499 n12681 ; n12713
g10278 and pi1198_not n12710 ; n12714
g10279 and pi1198 n12678_not ; n12715
g10280 nor n12713 n12715 ; n12716
g10281 and n12714_not n12716 ; n12717
g10282 and pi0374 n12717_not ; n12718
g10283 nor n12712 n12718 ; n12719
g10284 and pi0369 n12719_not ; n12720
g10285 nor pi0374 n12717 ; n12721
g10286 and pi0374 n12711_not ; n12722
g10287 nor n12721 n12722 ; n12723
g10288 nor pi0369 n12723 ; n12724
g10289 and pi0371 n8853 ; n12725
g10290 nor pi0371 n8853 ; n12726
g10291 nor n12725 n12726 ; n12727
g10292 and pi0370 n12727_not ; n12728
g10293 and pi0370_not n12727 ; n12729
g10294 nor n12728 n12729 ; n12730
g10295 and n12720_not n12730 ; n12731
g10296 and n12724_not n12731 ; n12732
g10297 nor pi0369 n12719 ; n12733
g10298 and pi0369 n12723_not ; n12734
g10299 nor n12730 n12733 ; n12735
g10300 and n12734_not n12735 ; n12736
g10301 nor pi0591 n12732 ; n12737
g10302 and n12736_not n12737 ; n12738
g10303 nor pi0590 n12675 ; n12739
g10304 and n12738_not n12739 ; n12740
g10305 nor pi0588 n12740 ; n12741
g10306 and n12566_not n12741 ; n12742
g10307 nor n7425 n12742 ; n12743
g10308 and n12492_not n12743 ; n12744
g10309 and n7429_not n12181 ; n12745
g10310 and pi0075 n12179 ; n12746
g10311 nor n12303 n12396 ; n12747
g10312 and n8162 n12312_not ; n12748
g10313 and n12747_not n12748 ; n12749
g10314 nor n12303 n12390 ; n12750
g10315 and n2610 n12312_not ; n12751
g10316 and n12750_not n12751 ; n12752
g10317 and n2625_not n12179 ; n12753
g10318 nor n12749 n12753 ; n12754
g10319 and n12752_not n12754 ; n12755
g10320 nor pi0075 n12755 ; n12756
g10321 nor n12746 n12756 ; n12757
g10322 and pi0567 n12757_not ; n12758
g10323 and n12568 n12758_not ; n12759
g10324 nor n12745 n12759 ; n12760
g10325 and pi0592_not n12760 ; n12761
g10326 nor n12275 n12761 ; n12762
g10327 and n8093_not n12762 ; n12763
g10328 and pi0443 n12762_not ; n12764
g10329 nor n12413 n12764 ; n12765
g10330 and n8249 n12765 ; n12766
g10331 nor pi0443 n12762 ; n12767
g10332 nor n12417 n12767 ; n12768
g10333 and n8249_not n12768 ; n12769
g10334 nor n12766 n12769 ; n12770
g10335 and pi0435 n12770_not ; n12771
g10336 and pi0444_not n12768 ; n12772
g10337 and pi0444 n12765 ; n12773
g10338 nor pi0436 n12772 ; n12774
g10339 and n12773_not n12774 ; n12775
g10340 and pi0444_not n12765 ; n12776
g10341 and pi0444 n12768 ; n12777
g10342 and pi0436 n12776_not ; n12778
g10343 and n12777_not n12778 ; n12779
g10344 nor n12775 n12779 ; n12780
g10345 and pi0435_not n12780 ; n12781
g10346 nor n12771 n12781 ; n12782
g10347 and pi0429_not n12782 ; n12783
g10348 nor pi0435 n12770 ; n12784
g10349 and pi0435 n12780 ; n12785
g10350 nor n12784 n12785 ; n12786
g10351 and pi0429 n12786 ; n12787
g10352 and n8105 n12783_not ; n12788
g10353 and n12787_not n12788 ; n12789
g10354 and pi0429_not n12786 ; n12790
g10355 and pi0429 n12782 ; n12791
g10356 nor n8105 n12790 ; n12792
g10357 and n12791_not n12792 ; n12793
g10358 and pi1196 n12789_not ; n12794
g10359 and n12793_not n12794 ; n12795
g10360 and n12412 n12795_not ; n12796
g10361 nor n12763 n12796 ; n12797
g10362 and pi1199_not n12797 ; n12798
g10363 nor pi0428 n12797 ; n12799
g10364 and pi0428 n12762 ; n12800
g10365 nor n12799 n12800 ; n12801
g10366 nor pi0427 n12801 ; n12802
g10367 and pi0428 n12797_not ; n12803
g10368 and pi0428_not n12762 ; n12804
g10369 nor n12803 n12804 ; n12805
g10370 and pi0427 n12805_not ; n12806
g10371 nor n12802 n12806 ; n12807
g10372 and pi0430 n12807_not ; n12808
g10373 nor pi0427 n12805 ; n12809
g10374 and pi0427 n12801_not ; n12810
g10375 nor n12809 n12810 ; n12811
g10376 nor pi0430 n12811 ; n12812
g10377 nor n12808 n12812 ; n12813
g10378 and pi0426 n12813_not ; n12814
g10379 and pi0430 n12811_not ; n12815
g10380 nor pi0430 n12807 ; n12816
g10381 nor n12815 n12816 ; n12817
g10382 nor pi0426 n12817 ; n12818
g10383 nor n12814 n12818 ; n12819
g10384 and pi0445 n12819_not ; n12820
g10385 and pi0426 n12817_not ; n12821
g10386 nor pi0426 n12813 ; n12822
g10387 nor n12821 n12822 ; n12823
g10388 nor pi0445 n12823 ; n12824
g10389 nor n12820 n12824 ; n12825
g10390 and pi0448 n12825 ; n12826
g10391 and pi0445 n12823_not ; n12827
g10392 nor pi0445 n12819 ; n12828
g10393 nor n12827 n12828 ; n12829
g10394 and pi0448_not n12829 ; n12830
g10395 and n8128 n12826_not ; n12831
g10396 and n12830_not n12831 ; n12832
g10397 and pi0448 n12829 ; n12833
g10398 and pi0448_not n12825 ; n12834
g10399 nor n8128 n12833 ; n12835
g10400 and n12834_not n12835 ; n12836
g10401 and pi1199 n12832_not ; n12837
g10402 and n12836_not n12837 ; n12838
g10403 and n8041 n12798_not ; n12839
g10404 and n12838_not n12839 ; n12840
g10405 and n12186 n12840_not ; n12841
g10406 nor n12273 n12762 ; n12842
g10407 and n8410 n12568 ; n12843
g10408 nor n12181 n12843 ; n12844
g10409 and n7958 n12745_not ; n12845
g10410 nor n12303 n12579 ; n12846
g10411 and n12748 n12846_not ; n12847
g10412 nor n12303 n12588 ; n12848
g10413 and n12751 n12848_not ; n12849
g10414 nor n12753 n12847 ; n12850
g10415 and n12849_not n12850 ; n12851
g10416 and n7926 n12749 ; n12852
g10417 and n12611_not n12752 ; n12853
g10418 nor n12852 n12853 ; n12854
g10419 and n12851 n12854 ; n12855
g10420 and n12845 n12855_not ; n12856
g10421 and n12629_not n12749 ; n12857
g10422 nor n12753 n12857 ; n12858
g10423 and n12853_not n12858 ; n12859
g10424 and n8668 n12745_not ; n12860
g10425 and n12859_not n12860 ; n12861
g10426 nor n12856 n12861 ; n12862
g10427 and pi0075_not pi0567 ; n12863
g10428 and n12862_not n12863 ; n12864
g10429 and pi1199 n12844_not ; n12865
g10430 and n12864_not n12865 ; n12866
g10431 nor pi0075 n12851 ; n12867
g10432 nor n12746 n12867 ; n12868
g10433 and pi0567 n12868_not ; n12869
g10434 and n12568 n12869_not ; n12870
g10435 and n12845 n12870_not ; n12871
g10436 and pi1199_not n12277 ; n12872
g10437 and n12871_not n12872 ; n12873
g10438 nor n8395 n12866 ; n12874
g10439 and n12873_not n12874 ; n12875
g10440 and pi1197_not n12875 ; n12876
g10441 nor n12842 n12876 ; n12877
g10442 nor pi0333 n12877 ; n12878
g10443 and n8395 n12762_not ; n12879
g10444 nor n12875 n12879 ; n12880
g10445 and pi0333 n12880_not ; n12881
g10446 nor n12878 n12881 ; n12882
g10447 nor pi0391 n12882 ; n12883
g10448 and pi0333 n12877_not ; n12884
g10449 nor pi0333 n12880 ; n12885
g10450 nor n12884 n12885 ; n12886
g10451 and pi0391 n12886_not ; n12887
g10452 nor n12883 n12887 ; n12888
g10453 nor pi0392 n12888 ; n12889
g10454 nor pi0391 n12886 ; n12890
g10455 and pi0391 n12882_not ; n12891
g10456 nor n12890 n12891 ; n12892
g10457 and pi0392 n12892_not ; n12893
g10458 nor n12889 n12893 ; n12894
g10459 nor pi0393 n12894 ; n12895
g10460 nor pi0392 n12892 ; n12896
g10461 and pi0392 n12888_not ; n12897
g10462 nor n12896 n12897 ; n12898
g10463 and pi0393 n12898_not ; n12899
g10464 nor n8028 n12895 ; n12900
g10465 and n12899_not n12900 ; n12901
g10466 nor pi0393 n12898 ; n12902
g10467 and pi0393 n12894_not ; n12903
g10468 and n8028 n12902_not ; n12904
g10469 and n12903_not n12904 ; n12905
g10470 and pi0591 n12901_not ; n12906
g10471 and n12905_not n12906 ; n12907
g10472 and pi0592 n12760 ; n12908
g10473 nor n12676 n12908 ; n12909
g10474 and n7722_not n12909 ; n12910
g10475 and pi1199 n12680_not ; n12911
g10476 and n12910_not n12911 ; n12912
g10477 and n7673 n7688 ; n12913
g10478 nor n7673 n7688 ; n12914
g10479 nor n12913 n12914 ; n12915
g10480 and pi0367 n12915_not ; n12916
g10481 and pi0367_not n12915 ; n12917
g10482 nor n12916 n12917 ; n12918
g10483 and n12181 n12918_not ; n12919
g10484 and n12909 n12918 ; n12920
g10485 and pi1197 n12919_not ; n12921
g10486 and n12920_not n12921 ; n12922
g10487 and n12685 n12922_not ; n12923
g10488 and n7670 n12909 ; n12924
g10489 nor pi1199 n12924 ; n12925
g10490 and n12923_not n12925 ; n12926
g10491 nor n12912 n12926 ; n12927
g10492 nor pi0374 n12927 ; n12928
g10493 nor pi1198 n12927 ; n12929
g10494 and pi1198 n12909_not ; n12930
g10495 nor n12929 n12930 ; n12931
g10496 and pi0374 n12931_not ; n12932
g10497 nor n12928 n12932 ; n12933
g10498 nor pi0369 n12933 ; n12934
g10499 nor pi0374 n12931 ; n12935
g10500 and pi0374 n12927_not ; n12936
g10501 nor n12935 n12936 ; n12937
g10502 and pi0369 n12937_not ; n12938
g10503 nor n12730 n12934 ; n12939
g10504 and n12938_not n12939 ; n12940
g10505 and pi0369 n12933_not ; n12941
g10506 nor pi0369 n12937 ; n12942
g10507 and n12730 n12941_not ; n12943
g10508 and n12942_not n12943 ; n12944
g10509 nor pi0591 n12940 ; n12945
g10510 and n12944_not n12945 ; n12946
g10511 nor pi0590 n12946 ; n12947
g10512 and n12907_not n12947 ; n12948
g10513 and n7850_not n12762 ; n12949
g10514 nor n12493 n12949 ; n12950
g10515 and pi1198 n12950_not ; n12951
g10516 and n7791_not n12762 ; n12952
g10517 nor n12498 n12952 ; n12953
g10518 and pi0355 n12953_not ; n12954
g10519 nor pi0455 n12762 ; n12955
g10520 nor n12502 n12955 ; n12956
g10521 nor pi0452 n12956 ; n12957
g10522 and pi0455 n12762_not ; n12958
g10523 nor n12506 n12958 ; n12959
g10524 and pi0452 n12959_not ; n12960
g10525 nor n12957 n12960 ; n12961
g10526 and pi0355_not n12961 ; n12962
g10527 nor n12954 n12962 ; n12963
g10528 and pi0458_not n12963 ; n12964
g10529 nor pi0355 n12953 ; n12965
g10530 and pi0355 n12961 ; n12966
g10531 nor n12965 n12966 ; n12967
g10532 and pi0458 n12967 ; n12968
g10533 nor n7812 n12964 ; n12969
g10534 and n12968_not n12969 ; n12970
g10535 and pi0458_not n12967 ; n12971
g10536 and pi0458 n12963 ; n12972
g10537 and n7812 n12971_not ; n12973
g10538 and n12972_not n12973 ; n12974
g10539 and pi1196 n12970_not ; n12975
g10540 and n12974_not n12975 ; n12976
g10541 and n12497 n12976_not ; n12977
g10542 nor n12951 n12977 ; n12978
g10543 nor n7782 n12978 ; n12979
g10544 and n7782 n12762 ; n12980
g10545 nor n12979 n12980 ; n12981
g10546 and n7757_not n12981 ; n12982
g10547 and pi1199 n12762_not ; n12983
g10548 and pi0351 n12983 ; n12984
g10549 nor n12982 n12984 ; n12985
g10550 nor pi0461 n12985 ; n12986
g10551 and n7862_not n12981 ; n12987
g10552 and pi0351_not n12983 ; n12988
g10553 nor n12987 n12988 ; n12989
g10554 and pi0461 n12989_not ; n12990
g10555 nor n12986 n12990 ; n12991
g10556 nor pi0357 n12991 ; n12992
g10557 nor pi0461 n12989 ; n12993
g10558 and pi0461 n12985_not ; n12994
g10559 nor n12993 n12994 ; n12995
g10560 and pi0357 n12995_not ; n12996
g10561 nor n12992 n12996 ; n12997
g10562 nor pi0356 n12997 ; n12998
g10563 nor pi0357 n12995 ; n12999
g10564 and pi0357 n12991_not ; n13000
g10565 nor n12999 n13000 ; n13001
g10566 and pi0356 n13001_not ; n13002
g10567 nor n12998 n13002 ; n13003
g10568 nor pi0354 n13003 ; n13004
g10569 nor pi0356 n13001 ; n13005
g10570 and pi0356 n12997_not ; n13006
g10571 nor n13005 n13006 ; n13007
g10572 and pi0354 n13007_not ; n13008
g10573 nor n7887 n13004 ; n13009
g10574 and n13008_not n13009 ; n13010
g10575 nor pi0354 n13007 ; n13011
g10576 and pi0354 n13003_not ; n13012
g10577 and n7887 n13011_not ; n13013
g10578 and n13012_not n13013 ; n13014
g10579 nor pi0591 n13010 ; n13015
g10580 and n13014_not n13015 ; n13016
g10581 and n12237 n13016_not ; n13017
g10582 nor pi0588 n12948 ; n13018
g10583 and n13017_not n13018 ; n13019
g10584 and n7425 n13019_not ; n13020
g10585 and n12841_not n13020 ; n13021
g10586 nor pi0080 po1038 ; n13022
g10587 and n12744_not n13022 ; n13023
g10588 and n13021_not n13023 ; n13024
g10589 nor pi0217 n12366 ; n13025
g10590 and n13024_not n13025 ; n13026
g10591 and n7643 n12183_not ; n13027
g10592 and n13026_not n13027 ; po0238
g10593 and po1038_not n11302 ; n13029
g10594 and pi0081 pi0314_not ; n13030
g10595 and n2489 n13030 ; n13031
g10596 and pi0068 pi0081_not ; n13032
g10597 and n2480 n13032 ; n13033
g10598 and n11014 n13033 ; n13034
g10599 and n11439 n13034 ; n13035
g10600 and n2800 n13035 ; n13036
g10601 nor n13031 n13036 ; n13037
g10602 and n13029 n13037_not ; po0239
g10603 and pi0069 pi0314 ; n13039
g10604 and n2792 n13039 ; n13040
g10605 and pi0066 pi0073_not ; n13041
g10606 and n2468 n13041 ; n13042
g10607 and n2482 n13042 ; n13043
g10608 nor n13040 n13043 ; n13044
g10609 and n11103 n11107 ; n13045
g10610 and n13044_not n13045 ; po0240
g10611 and n2480 n2799 ; n13047
g10612 and pi0084 n9077 ; n13048
g10613 and n13047 n13048 ; n13049
g10614 and n2467 n13049 ; n13050
g10615 and n2499 n11102 ; n13051
g10616 and n2702 n13051 ; n13052
g10617 and n13050 n13052 ; n13053
g10618 and pi0314 n13053_not ; n13054
g10619 nor pi0083 n13049 ; n13055
g10620 and n13052 n13055_not ; n13056
g10621 and n2795 n13056 ; n13057
g10622 nor pi0314 n13057 ; n13058
g10623 and n10166 n13054_not ; n13059
g10624 and n13058_not n13059 ; po0241
g10625 and pi0211 pi0299 ; n13061
g10626 and pi0219 pi0299 ; n13062
g10627 nor n13061 n13062 ; n13063
g10628 and n10810_not n13063 ; n13064
g10629 and po1038_not n13064 ; n13065
g10630 and n11385 n13065 ; po0242
g10631 and n6423 n11104 ; n13067
g10632 and pi0314_not n11105 ; n13068
g10633 and n11437 n13068 ; n13069
g10634 nor n13067 n13069 ; n13070
g10635 and n11107 n13070_not ; po0243
g10636 and n7603 n11396 ; n13072
g10637 and n7606 n11399 ; n13073
g10638 nor n13072 n13073 ; n13074
g10639 and n10983 n13074_not ; po0244
g10640 and n2845 n13051 ; n13076
g10641 and pi0314 n10166 ; n13077
g10642 and n2702 n13077 ; n13078
g10643 and n13076 n13078 ; po0245
g10644 and n2708 n7417 ; n13080
g10645 and pi1093_not n2519 ; n13081
g10646 and n2572 n13081 ; n13082
g10647 and n13080 n13082 ; n13083
g10648 and n11460 n13083 ; n13084
g10649 and n2870 n13084 ; n13085
g10650 nor n7425 n13085 ; n13086
g10651 and n7417 n11030 ; n13087
g10652 nor pi1093 n13087 ; n13088
g10653 and n7439 n12376 ; n13089
g10654 and n11027 n13089 ; n13090
g10655 and n11043 n12374 ; n13091
g10656 and n13090 n13091 ; n13092
g10657 and pi1093 n13092_not ; n13093
g10658 and n2572 n10074_not ; n13094
g10659 and n13093_not n13094 ; n13095
g10660 and n13088_not n13095 ; n13096
g10661 and n7425 n13096_not ; n13097
g10662 nor po1038 n13086 ; n13098
g10663 and n13097_not n13098 ; po0246
g10664 and n2465 n8921 ; n13100
g10665 and n8935 n13100 ; n13101
g10666 and n10181 n13101 ; n13102
g10667 and pi0841 n7445 ; n13103
g10668 and n13102 n13103 ; n13104
g10669 nor pi0070 n13104 ; n13105
g10670 and pi0070 n8959_not ; n13106
g10671 and n2520 n10165 ; n13107
g10672 and n13105_not n13107 ; n13108
g10673 and n13106_not n13108 ; po0247
g10674 and pi1050_not n9090 ; n13110
g10675 nor pi0090 n13110 ; n13111
g10676 and n11326 n13111_not ; n13112
g10677 and n2896_not n13112 ; n13113
g10678 and n7433_not n13113 ; po0248
g10679 and pi0058_not n2756 ; n13115
g10680 nor n10158 n13115 ; n13116
g10681 and n2928 n10162 ; n13117
g10682 and n13116_not n13117 ; n13118
g10683 and pi0024 n2938 ; n13119
g10684 and n2928_not n13119 ; n13120
g10685 and n11086 n13120 ; n13121
g10686 and n2756 n13121 ; n13122
g10687 nor pi0039 n13122 ; n13123
g10688 and n13118_not n13123 ; n13124
g10689 and n10197 n13124_not ; n13125
g10690 and n7612 n13125 ; po0249
g10691 and pi0092 n2521 ; n13127
g10692 and n3373 n11473 ; n13128
g10693 and n13127 n13128 ; n13129
g10694 and n5853 n6235 ; n13130
g10695 and n7603 n13130 ; n13131
g10696 and n3470 n6189 ; n13132
g10697 and n7606 n13132 ; n13133
g10698 nor n13131 n13133 ; n13134
g10699 and n2534 n11211 ; n13135
g10700 and n13134_not n13135 ; n13136
g10701 nor n13129 n13136 ; n13137
g10702 and n10163 n13137_not ; po0250
g10703 and pi0093 n11086 ; n13139
g10704 and n2914 n13139 ; n13140
g10705 nor pi0092 n13140 ; n13141
g10706 and pi1050_not n2521 ; n13142
g10707 and pi0092 n13142_not ; n13143
g10708 and n10164 n13141_not ; n13144
g10709 and n13143_not n13144 ; po0251
g10710 and n11068 n11284 ; n13146
g10711 nor n8888 n13146 ; n13147
g10712 and n2924 n13146 ; n13148
g10713 and pi1093 n13148_not ; n13149
g10714 and n2933 n13149_not ; n13150
g10715 and n10243 n11066 ; n13151
g10716 nor n2780 n13151 ; n13152
g10717 and n2717 n10162 ; n13153
g10718 and pi0252 n13153 ; n13154
g10719 and n13152_not n13154 ; n13155
g10720 nor n13150 n13155 ; n13156
g10721 nor po0840 n13156 ; n13157
g10722 nor n13146 n13157 ; n13158
g10723 and pi0252 n13156 ; n13159
g10724 nor n13158 n13159 ; n13160
g10725 and n8888 n13160_not ; n13161
g10726 and n10165 n13147_not ; n13162
g10727 and n13161_not n13162 ; po0252
g10728 and n2517 n11770 ; n13164
g10729 and n11458 n13164 ; n13165
g10730 and pi0332_not n10162 ; n13166
g10731 and n11283 n13166 ; n13167
g10732 and n13102 n13167 ; n13168
g10733 nor pi0039 n13168 ; n13169
g10734 and n13165_not n13169 ; n13170
g10735 and n11422_not n11425 ; n13171
g10736 and n6392_not n13171 ; n13172
g10737 nor n6207 n6392 ; n13173
g10738 and n3471 n11419_not ; n13174
g10739 and n13173 n13174 ; n13175
g10740 and pi0039 n13172_not ; n13176
g10741 and n13175_not n13176 ; n13177
g10742 and n10200 n13170_not ; n13178
g10743 and n13177_not n13178 ; po0253
g10744 and n10325 n13164 ; n13180
g10745 and pi0479 po0840_not ; n13181
g10746 and n3183 n13181 ; n13182
g10747 and pi0096 n2510 ; n13183
g10748 and n2961 n13183 ; n13184
g10749 and n13181_not n13184 ; n13185
g10750 and n2916 n13185 ; n13186
g10751 nor n13182 n13186 ; n13187
g10752 nor pi0095 n13187 ; n13188
g10753 nor n13180 n13188 ; n13189
g10754 and n10165 n13189_not ; po0254
g10755 and pi0039 pi0593 ; n13191
g10756 and n11427_not n13191 ; n13192
g10757 and n6392_not n13192 ; n13193
g10758 and n6169 n13181 ; n13194
g10759 nor po0740 n13194 ; n13195
g10760 and pi0096_not n10193 ; n13196
g10761 and n13195_not n13196 ; n13197
g10762 and n11486 n13197 ; n13198
g10763 nor n13193 n13198 ; n13199
g10764 and n10200 n13199_not ; po0255
g10765 and pi0092_not n11474 ; n13201
g10766 nor n13127 n13201 ; n13202
g10767 and pi0314 pi1050 ; n13203
g10768 and n10164 n13203 ; n13204
g10769 and n13202_not n13204 ; po0256
g10770 and pi0072_not pi0152 ; n13206
g10771 and n10300 n13206 ; n13207
g10772 and pi0299 n13207 ; n13208
g10773 and pi0072_not pi0174 ; n13209
g10774 and pi0299_not n13209 ; n13210
g10775 and n10296 n13210 ; n13211
g10776 nor n13208 n13211 ; n13212
g10777 and pi0232 n13212_not ; n13213
g10778 and pi0039 n13213_not ; n13214
g10779 and pi0072_not pi0099 ; n13215
g10780 nor pi0039 n13215 ; n13216
g10781 nor n13214 n13216 ; n13217
g10782 and n2620_not n13217 ; n13218
g10783 nor n7506 n13215 ; n13219
g10784 and n2924_not n13215 ; n13220
g10785 and n7506 n13220_not ; n13221
g10786 and n10329_not n13215 ; n13222
g10787 and n6266 n10919 ; n13223
g10788 nor n13222 n13223 ; n13224
g10789 and n10356 n13224_not ; n13225
g10790 and n13221 n13225_not ; n13226
g10791 nor n13219 n13226 ; n13227
g10792 nor pi0039 n13227 ; n13228
g10793 and n2620 n13214_not ; n13229
g10794 and n13228_not n13229 ; n13230
g10795 and pi0075 n13218_not ; n13231
g10796 and n13230_not n13231 ; n13232
g10797 and pi0228 n10500 ; n13233
g10798 and pi0228 n10344 ; n13234
g10799 and n13215 n13234_not ; n13235
g10800 and n2531 n13235_not ; n13236
g10801 and n13233_not n13236 ; n13237
g10802 nor n2531 n13217 ; n13238
g10803 and pi0087 n13238_not ; n13239
g10804 and n13237_not n13239 ; n13240
g10805 and pi0038 n13217_not ; n13241
g10806 and n10478 n13212_not ; n13242
g10807 and n10948_not n13242 ; n13243
g10808 and pi0041 pi0072 ; n13244
g10809 and pi0099 n13244_not ; n13245
g10810 and n10411_not n13245 ; n13246
g10811 nor pi0228 n10556 ; n13247
g10812 and n13246_not n13247 ; n13248
g10813 and n10459_not n13245 ; n13249
g10814 and n10779 n13249_not ; n13250
g10815 and n10426_not n13245 ; n13251
g10816 and n10778 n13251_not ; n13252
g10817 nor n13250 n13252 ; n13253
g10818 and pi0228 n13253_not ; n13254
g10819 nor pi0039 n13248 ; n13255
g10820 and n13254_not n13255 ; n13256
g10821 and n2608 n13243_not ; n13257
g10822 and n13256_not n13257 ; n13258
g10823 and n10359_not n13215 ; n13259
g10824 and n6265 n10318 ; n13260
g10825 nor n13259 n13260 ; n13261
g10826 and n10356 n13261_not ; n13262
g10827 and n13221 n13262_not ; n13263
g10828 nor n13219 n13263 ; n13264
g10829 nor pi0039 n13264 ; n13265
g10830 nor n13214 n13265 ; n13266
g10831 and n6285 n13266_not ; n13267
g10832 nor pi0087 n13241 ; n13268
g10833 and n13267_not n13268 ; n13269
g10834 and n13258_not n13269 ; n13270
g10835 nor pi0075 n13240 ; n13271
g10836 and n13270_not n13271 ; n13272
g10837 nor n13232 n13272 ; n13273
g10838 and n7429 n13273_not ; n13274
g10839 nor n7429 n13217 ; n13275
g10840 nor po1038 n13275 ; n13276
g10841 and n13274_not n13276 ; n13277
g10842 and pi0232 n13207 ; n13278
g10843 and pi0039 n13278_not ; n13279
g10844 and po1038 n13216_not ; n13280
g10845 and n13279_not n13280 ; n13281
g10846 or n13277 n13281 ; po0257
g10847 nor n6263 n6281 ; n13283
g10848 and n7473_not n10078 ; n13284
g10849 and pi0129 n13284_not ; n13285
g10850 and n7472 n13285_not ; n13286
g10851 and pi0129 n10078_not ; n13287
g10852 nor n10081 n13287 ; n13288
g10853 nor n13283 n13288 ; n13289
g10854 and n13286_not n13289 ; n13290
g10855 and pi0075_not n2609 ; n13291
g10856 and n6285 n13291 ; n13292
g10857 and n13290_not n13292 ; n13293
g10858 and pi0024_not n8967 ; n13294
g10859 and po0840 n13294 ; n13295
g10860 and n8964_not n13295 ; n13296
g10861 nor n13293 n13296 ; n13297
g10862 and n8881 n13297_not ; n13298
g10863 and n2521 n13298 ; po0258
g10864 nor pi0039 n10322 ; n13300
g10865 and pi0152 n3389 ; n13301
g10866 and n6197 n13301 ; n13302
g10867 and pi0072_not n13302 ; n13303
g10868 and pi0299 n13303_not ; n13304
g10869 and pi0144_not pi0174 ; n13305
g10870 and n10295 n13305 ; n13306
g10871 and pi0072_not n13306 ; n13307
g10872 nor pi0299 n13307 ; n13308
g10873 and pi0232 n13304_not ; n13309
g10874 and n13308_not n13309 ; n13310
g10875 and pi0039 n13310_not ; n13311
g10876 nor n13300 n13311 ; n13312
g10877 and n2620_not n13312 ; n13313
g10878 nor n7506 n10322 ; n13314
g10879 and n2924_not n10322 ; n13315
g10880 and n7506 n13315_not ; n13316
g10881 and n2924 n6273_not ; n13317
g10882 and n10322 n10328_not ; n13318
g10883 nor n10319 n13318 ; n13319
g10884 and n13317 n13319_not ; n13320
g10885 and n13316 n13320_not ; n13321
g10886 nor n13314 n13321 ; n13322
g10887 nor pi0039 n13322 ; n13323
g10888 and n2620 n13311_not ; n13324
g10889 and n13323_not n13324 ; n13325
g10890 and pi0075 n13313_not ; n13326
g10891 and n13325_not n13326 ; n13327
g10892 and n10343 n10931 ; n13328
g10893 and n10322 n13328_not ; n13329
g10894 and pi0101_not n10932 ; n13330
g10895 nor pi0039 n13329 ; n13331
g10896 and n13330_not n13331 ; n13332
g10897 and pi0087 n13311_not ; n13333
g10898 and n13332_not n13333 ; n13334
g10899 and pi0038 n13312_not ; n13335
g10900 and n10949 n13302 ; n13336
g10901 and pi0299 n13336_not ; n13337
g10902 and n10949 n13306 ; n13338
g10903 nor pi0299 n13338 ; n13339
g10904 and n10478 n13337_not ; n13340
g10905 and n13339_not n13340 ; n13341
g10906 and pi0101 n10409 ; n13342
g10907 nor pi0228 n10401 ; n13343
g10908 and n13342_not n13343 ; n13344
g10909 and pi0101 n10457 ; n13345
g10910 and n2924 n10451_not ; n13346
g10911 and n13345_not n13346 ; n13347
g10912 and pi0101 n10424 ; n13348
g10913 nor n2924 n10433 ; n13349
g10914 and n13348_not n13349 ; n13350
g10915 nor n13347 n13350 ; n13351
g10916 and pi0228 n13351_not ; n13352
g10917 nor pi0039 n13344 ; n13353
g10918 and n13352_not n13353 ; n13354
g10919 and n2608 n13341_not ; n13355
g10920 and n13354_not n13355 ; n13356
g10921 and pi0044_not n10940 ; n13357
g10922 and n10322 n13357_not ; n13358
g10923 nor n10318 n13358 ; n13359
g10924 and n13317 n13359_not ; n13360
g10925 and n13316 n13360_not ; n13361
g10926 nor n13314 n13361 ; n13362
g10927 nor pi0039 n13362 ; n13363
g10928 nor n13311 n13363 ; n13364
g10929 and n6285 n13364_not ; n13365
g10930 nor pi0087 n13335 ; n13366
g10931 and n13365_not n13366 ; n13367
g10932 and n13356_not n13367 ; n13368
g10933 nor pi0075 n13334 ; n13369
g10934 and n13368_not n13369 ; n13370
g10935 nor n13327 n13370 ; n13371
g10936 and n7429 n13371_not ; n13372
g10937 nor n7429 n13312 ; n13373
g10938 nor po1038 n13373 ; n13374
g10939 and n13372_not n13374 ; n13375
g10940 and pi0232 n13303 ; n13376
g10941 and pi0039 n13376_not ; n13377
g10942 and po1038 n13300_not ; n13378
g10943 and n13377_not n13378 ; n13379
g10944 or n13375 n13379 ; po0259
g10945 and n2851 n8922 ; n13381
g10946 and n13029 n13381 ; po0260
g10947 and pi0109 n2765 ; n13383
g10948 and n2699 n13383 ; n13384
g10949 and pi0314 n13384_not ; n13385
g10950 nor pi0109 n13076 ; n13386
g10951 and n6422 n13386_not ; n13387
g10952 nor pi0314 n13387 ; n13388
g10953 and n11106 n13385_not ; n13389
g10954 and n13388_not n13389 ; po0261
g10955 and n7425 n8888_not ; n13391
g10956 and n10075 n13391_not ; n13392
g10957 and n10396 n13392_not ; n13393
g10958 and po1057 n13092_not ; n13394
g10959 nor pi0110 n13090 ; n13395
g10960 and pi0047_not n11043 ; n13396
g10961 and n13395_not n13396 ; n13397
g10962 and n10378 n13397 ; n13398
g10963 nor po1057 n13398 ; n13399
g10964 nor n7474 n10074 ; n13400
g10965 and n13394_not n13400 ; n13401
g10966 and n13399_not n13401 ; n13402
g10967 and n7474 n10074_not ; n13403
g10968 and n13398 n13403 ; n13404
g10969 nor n13402 n13404 ; n13405
g10970 nor n7425 n13405 ; n13406
g10971 nor n13393 n13406 ; n13407
g10972 and n10165 n13407_not ; po0262
g10973 and pi0024 n11282 ; n13409
g10974 nor pi0053 n11281 ; n13410
g10975 and n2723 n13410_not ; n13411
g10976 and pi0024_not n2717 ; n13412
g10977 and n13411 n13412 ; n13413
g10978 nor n13409 n13413 ; n13414
g10979 and pi0841 n13414_not ; n13415
g10980 and n8946 n11267 ; n13416
g10981 nor n13415 n13416 ; n13417
g10982 and n10166 n13417_not ; po0264
g10983 and pi0999_not n10166 ; n13419
g10984 and n11354 n13419 ; po0265
g10985 and pi0097_not n7442 ; n13421
g10986 nor pi0108 n13421 ; n13422
g10987 and n2701 n13422_not ; n13423
g10988 and n10244 n13423 ; n13424
g10989 nor pi0314 n13424 ; n13425
g10990 and pi0314 n7444_not ; n13426
g10991 and n7446 n10238_not ; n13427
g10992 and n13426_not n13427 ; n13428
g10993 and n13425_not n13428 ; n13429
g10994 and n7446 n10238 ; n13430
g10995 and n13424 n13430 ; n13431
g10996 nor pi0051 n13431 ; n13432
g10997 and n13429_not n13432 ; n13433
g10998 and n2625 n7518 ; n13434
g10999 and n13433_not n13434 ; n13435
g11000 nor pi0087 n13435 ; n13436
g11001 and n6133 n8881 ; n13437
g11002 and n13436_not n13437 ; po0266
g11003 and n2784 n11442 ; n13439
g11004 and n13077 n13439 ; po0267
g11005 nor pi0082 pi0109 ; n13441
g11006 and pi0111 n13441 ; n13442
g11007 and n12374 n13442 ; n13443
g11008 and n2499 n13443 ; n13444
g11009 and n11105 n13444 ; n13445
g11010 and n2801 n13445 ; n13446
g11011 and pi0314 n13446 ; n13447
g11012 and n8888 n10075 ; n13448
g11013 and n10388 n13448 ; n13449
g11014 nor n13447 n13449 ; n13450
g11015 and n10166 n13450_not ; po0268
g11016 and pi0072 n10325 ; n13452
g11017 and pi0314_not n13446 ; n13453
g11018 and n9141 n13453 ; n13454
g11019 nor n13452 n13454 ; n13455
g11020 and n6479 n10165 ; n13456
g11021 and n13455_not n13456 ; po0269
g11022 nand pi0124 pi0468_not ; po0270
g11023 and pi0072_not pi0113 ; n13459
g11024 and pi0039_not n13459 ; n13460
g11025 and pi0038 n13460_not ; n13461
g11026 and n2924 n7506 ; n13462
g11027 and n7479 n10531 ; n13463
g11028 nor n6272 n13463 ; n13464
g11029 and n13462 n13464_not ; n13465
g11030 and n13459 n13465_not ; n13466
g11031 and n6272_not n13462 ; n13467
g11032 and pi0113_not n13467 ; n13468
g11033 and n13260 n13468 ; n13469
g11034 nor n13466 n13469 ; n13470
g11035 nor pi0039 n13470 ; n13471
g11036 and n6285 n13471_not ; n13472
g11037 and pi0113 n10550 ; n13473
g11038 nor pi0228 n10557 ; n13474
g11039 and n13473_not n13474 ; n13475
g11040 and pi0113_not n10780 ; n13476
g11041 nor n2924 n10426 ; n13477
g11042 nor pi0099 n13477 ; n13478
g11043 and n10460_not n13478 ; n13479
g11044 and pi0113 n10548_not ; n13480
g11045 and n13479_not n13480 ; n13481
g11046 and pi0228 n13476_not ; n13482
g11047 and n13481_not n13482 ; n13483
g11048 nor pi0039 n13475 ; n13484
g11049 and n13483_not n13484 ; n13485
g11050 and n2608 n13485_not ; n13486
g11051 nor n13461 n13472 ; n13487
g11052 and n13486_not n13487 ; n13488
g11053 nor pi0087 n13488 ; n13489
g11054 and n2608_not n13460 ; n13490
g11055 and n10532_not n13459 ; n13491
g11056 and pi0113_not n13233 ; n13492
g11057 nor n13491 n13492 ; n13493
g11058 and n2531 n13493_not ; n13494
g11059 and pi0087 n13490_not ; n13495
g11060 and n13494_not n13495 ; n13496
g11061 nor n13489 n13496 ; n13497
g11062 nor pi0075 n13497 ; n13498
g11063 and n7477 n13469 ; n13499
g11064 nor n6272 n10496 ; n13500
g11065 and n13462 n13500_not ; n13501
g11066 and n13459 n13501_not ; n13502
g11067 nor n13499 n13502 ; n13503
g11068 and n2610 n13503_not ; n13504
g11069 and n2620_not n13460 ; n13505
g11070 and pi0075 n13505_not ; n13506
g11071 and n13504_not n13506 ; n13507
g11072 nor n13498 n13507 ; n13508
g11073 and n8881 n13508_not ; n13509
g11074 nor n8881 n13460 ; n13510
g11075 nor n13509 n13510 ; po0271
g11076 and pi0072_not pi0114 ; n13512
g11077 and pi0039_not n13512 ; n13513
g11078 and n2620_not n13513 ; n13514
g11079 nor n11143 n13512 ; n13515
g11080 and pi0114 n10735 ; n13516
g11081 and n11143 n13516_not ; n13517
g11082 and n10505_not n13517 ; n13518
g11083 and n2610 n13515_not ; n13519
g11084 and n13518_not n13519 ; n13520
g11085 and pi0075 n13514_not ; n13521
g11086 and n13520_not n13521 ; n13522
g11087 nor n2608 n13513 ; n13523
g11088 and pi0228 n10616 ; n13524
g11089 and pi0115_not n13524 ; n13525
g11090 and n13512 n13525_not ; n13526
g11091 and n2608 n13526_not ; n13527
g11092 and n10537_not n13527 ; n13528
g11093 and n11212 n13523_not ; n13529
g11094 and n13528_not n13529 ; n13530
g11095 and pi0038 n13513_not ; n13531
g11096 and pi0114 n10618_not ; n13532
g11097 and n11143 n13532_not ; n13533
g11098 and n10504_not n13533 ; n13534
g11099 nor pi0039 n13515 ; n13535
g11100 and n13534_not n13535 ; n13536
g11101 and n6285 n13536_not ; n13537
g11102 nor pi0114 n10783 ; n13538
g11103 and pi0114 n10791_not ; n13539
g11104 nor n13538 n13539 ; n13540
g11105 nor pi0115 n13540 ; n13541
g11106 and pi0115 n13512_not ; n13542
g11107 nor pi0039 n13542 ; n13543
g11108 and n13541_not n13543 ; n13544
g11109 and n2608 n13544_not ; n13545
g11110 nor pi0087 n13531 ; n13546
g11111 and n13537_not n13546 ; n13547
g11112 and n13545_not n13547 ; n13548
g11113 nor pi0075 n13530 ; n13549
g11114 and n13548_not n13549 ; n13550
g11115 nor n13522 n13550 ; n13551
g11116 and n8881 n13551_not ; n13552
g11117 nor n8881 n13513 ; n13553
g11118 nor n13552 n13553 ; po0272
g11119 and pi0072_not pi0115 ; n13555
g11120 and pi0039_not n13555 ; n13556
g11121 and n2620_not n13556 ; n13557
g11122 nor n13462 n13555 ; n13558
g11123 and pi0115 n10735 ; n13559
g11124 and pi0052_not n11125 ; n13560
g11125 nor pi0115 n13560 ; n13561
g11126 and n10502 n13561 ; n13562
g11127 and n7477 n13562 ; n13563
g11128 and n13462 n13559_not ; n13564
g11129 and n13563_not n13564 ; n13565
g11130 and n2610 n13558_not ; n13566
g11131 and n13565_not n13566 ; n13567
g11132 and pi0075 n13557_not ; n13568
g11133 and n13567_not n13568 ; n13569
g11134 nor n2608 n13556 ; n13570
g11135 and n13524_not n13555 ; n13571
g11136 and n2608 n13571_not ; n13572
g11137 and n10536_not n13572 ; n13573
g11138 and n11212 n13570_not ; n13574
g11139 and n13573_not n13574 ; n13575
g11140 and pi0038 n13556_not ; n13576
g11141 and pi0115 n10618_not ; n13577
g11142 and n13462 n13577_not ; n13578
g11143 and n13562_not n13578 ; n13579
g11144 nor pi0039 n13558 ; n13580
g11145 and n13579_not n13580 ; n13581
g11146 and n6285 n13581_not ; n13582
g11147 nor pi0115 n10783 ; n13583
g11148 and pi0115 n10791_not ; n13584
g11149 nor pi0039 n13583 ; n13585
g11150 and n13584_not n13585 ; n13586
g11151 and n2608 n13586_not ; n13587
g11152 nor pi0087 n13576 ; n13588
g11153 and n13582_not n13588 ; n13589
g11154 and n13587_not n13589 ; n13590
g11155 nor pi0075 n13575 ; n13591
g11156 and n13590_not n13591 ; n13592
g11157 nor n13569 n13592 ; n13593
g11158 and n8881 n13593_not ; n13594
g11159 nor n8881 n13556 ; n13595
g11160 nor n13594 n13595 ; po0273
g11161 and pi0072_not pi0116 ; n13597
g11162 and pi0039_not n13597 ; n13598
g11163 and pi0038 n13598_not ; n13599
g11164 and pi0113_not n10532 ; n13600
g11165 and n13597 n13600_not ; n13601
g11166 nor pi0038 n13601 ; n13602
g11167 and n10535_not n13602 ; n13603
g11168 nor n13599 n13603 ; n13604
g11169 nor pi0100 n13604 ; n13605
g11170 and pi0100 n13598_not ; n13606
g11171 and n11212 n13606_not ; n13607
g11172 and n13605_not n13607 ; n13608
g11173 and n2924_not n10580 ; n13609
g11174 and pi0116 n10585 ; n13610
g11175 nor n2924 n13610 ; n13611
g11176 and n2924 n10568_not ; n13612
g11177 and pi0116 n13612_not ; n13613
g11178 nor n10573 n13613 ; n13614
g11179 nor n13611 n13614 ; n13615
g11180 and pi0228 n13609_not ; n13616
g11181 and n13615_not n13616 ; n13617
g11182 and pi0116 n10552 ; n13618
g11183 and n10777 n13618_not ; n13619
g11184 nor pi0039 n13619 ; n13620
g11185 and n13617_not n13620 ; n13621
g11186 and n2608 n13621_not ; n13622
g11187 and n13462_not n13597 ; n13623
g11188 and pi0113_not n13463 ; n13624
g11189 and n13597 n13624_not ; n13625
g11190 nor n10502 n13625 ; n13626
g11191 and n13467 n13626_not ; n13627
g11192 nor n13623 n13627 ; n13628
g11193 nor pi0039 n13628 ; n13629
g11194 and n6285 n13629_not ; n13630
g11195 nor pi0087 n13599 ; n13631
g11196 and n13630_not n13631 ; n13632
g11197 and n13622_not n13632 ; n13633
g11198 nor pi0075 n13608 ; n13634
g11199 and n13633_not n13634 ; n13635
g11200 and n10497_not n13597 ; n13636
g11201 nor n10738 n13636 ; n13637
g11202 and n13467 n13637_not ; n13638
g11203 nor n13623 n13638 ; n13639
g11204 and n2610 n13639_not ; n13640
g11205 and n2620_not n13598 ; n13641
g11206 and pi0075 n13641_not ; n13642
g11207 and n13640_not n13642 ; n13643
g11208 nor n13635 n13643 ; n13644
g11209 and n8881 n13644_not ; n13645
g11210 nor n8881 n13598 ; n13646
g11211 nor n13645 n13646 ; po0274
g11212 and n3686 n7379 ; n13648
g11213 nor n3685 n13648 ; n13649
g11214 nor pi0038 n13649 ; n13650
g11215 nor pi0087 n13650 ; n13651
g11216 and n6133 n13651_not ; n13652
g11217 nor pi0092 n13652 ; n13653
g11218 nor pi0054 n7305 ; n13654
g11219 and pi0074_not n13654 ; n13655
g11220 and n13653_not n13655 ; n13656
g11221 nor pi0055 n13656 ; n13657
g11222 nor n7347 n13657 ; n13658
g11223 nor pi0056 n13658 ; n13659
g11224 nor n6127 n13659 ; n13660
g11225 nor pi0062 n13660 ; n13661
g11226 and pi0057_not n6300 ; n13662
g11227 and n13661_not n13662 ; po0275
g11228 and pi0079_not n12169 ; n13664
g11229 and pi0163 n6197 ; n13665
g11230 nor n11678 n13665 ; n13666
g11231 nor pi0150 n13666 ; n13667
g11232 and pi0150 n9699 ; n13668
g11233 and n11676 n13668 ; n13669
g11234 nor n13667 n13669 ; n13670
g11235 and pi0232 n13670_not ; n13671
g11236 and n8989_not n13671 ; n13672
g11237 and pi0074 n13672_not ; n13673
g11238 and pi0165 n7473 ; n13674
g11239 nor pi0038 pi0054 ; n13675
g11240 nor n13674 n13675 ; n13676
g11241 and n8989 n13676 ; n13677
g11242 nor pi0074 n13672 ; n13678
g11243 and n13677_not n13678 ; n13679
g11244 nor n13673 n13679 ; n13680
g11245 nor n2529 n13680 ; n13681
g11246 and n3328 n13681_not ; n13682
g11247 nor n9883 n13682 ; n13683
g11248 and pi0055 n13673_not ; n13684
g11249 and pi0150 n7473 ; n13685
g11250 and pi0092_not n9282 ; n13686
g11251 and n13685 n13686 ; n13687
g11252 and n9248 n13675 ; n13688
g11253 and n13687_not n13688 ; n13689
g11254 nor n13676 n13689 ; n13690
g11255 and n8989 n13690_not ; n13691
g11256 and n13678 n13691_not ; n13692
g11257 and n13684 n13692_not ; n13693
g11258 nor pi0184 n11704 ; n13694
g11259 and pi0185 n13694_not ; n13695
g11260 and pi0185_not n13694 ; n13696
g11261 and n6197 n13695_not ; n13697
g11262 and n13696_not n13697 ; n13698
g11263 nor pi0299 n13698 ; n13699
g11264 and pi0299 n13670 ; n13700
g11265 and pi0232 n13699_not ; n13701
g11266 and n13700_not n13701 ; n13702
g11267 and n8989_not n13702 ; n13703
g11268 and pi0074 n13703_not ; n13704
g11269 nor pi0055 n13704 ; n13705
g11270 nor pi0143 pi0299 ; n13706
g11271 and pi0165_not pi0299 ; n13707
g11272 nor n13706 n13707 ; n13708
g11273 and n7473 n13708 ; n13709
g11274 and n8989 n13709_not ; n13710
g11275 and pi0054 n13710_not ; n13711
g11276 and n13703_not n13711 ; n13712
g11277 and pi0075 n13702_not ; n13713
g11278 and pi0100 n13702_not ; n13714
g11279 and pi0038 n13709_not ; n13715
g11280 nor pi0100 n13715 ; n13716
g11281 and pi0157_not pi0299 ; n13717
g11282 nor pi0178 pi0299 ; n13718
g11283 nor n13717 n13718 ; n13719
g11284 and n7473 n13719 ; n13720
g11285 and n9282 n13720 ; n13721
g11286 and n9249 n13721_not ; n13722
g11287 and n13716 n13722_not ; n13723
g11288 nor n13714 n13723 ; n13724
g11289 and n9205 n13724_not ; n13725
g11290 nor pi0143 n9187 ; n13726
g11291 and pi0143 n9189_not ; n13727
g11292 and pi0165 n13727_not ; n13728
g11293 and n13726_not n13728 ; n13729
g11294 and pi0143 pi0165_not ; n13730
g11295 and n9194 n13730 ; n13731
g11296 and pi0038 n13731_not ; n13732
g11297 and n13729_not n13732 ; n13733
g11298 and n2568 n13733_not ; n13734
g11299 and pi0232_not n9532 ; n13735
g11300 nor n6197 n9532 ; n13736
g11301 and n6197 n9574_not ; n13737
g11302 nor n13736 n13737 ; n13738
g11303 and pi0151 pi0168 ; n13739
g11304 and n13738_not n13739 ; n13740
g11305 and n6197_not n9532 ; n13741
g11306 and pi0151 pi0168_not ; n13742
g11307 and n9606_not n13742 ; n13743
g11308 and pi0168_not n9615 ; n13744
g11309 and pi0168 n9612 ; n13745
g11310 nor pi0151 n13744 ; n13746
g11311 and n13745_not n13746 ; n13747
g11312 nor n13743 n13747 ; n13748
g11313 nor n13741 n13748 ; n13749
g11314 and pi0150 n13740_not ; n13750
g11315 and n13749_not n13750 ; n13751
g11316 and pi0168 n6197 ; n13752
g11317 and n9532 n13752_not ; n13753
g11318 and pi0168 n9506 ; n13754
g11319 nor pi0151 n13753 ; n13755
g11320 and n13754_not n13755 ; n13756
g11321 nor n9645 n13736 ; n13757
g11322 and pi0168_not n13757 ; n13758
g11323 nor n9445 n13736 ; n13759
g11324 and pi0168 n13759 ; n13760
g11325 and pi0151 n13758_not ; n13761
g11326 and n13760_not n13761 ; n13762
g11327 nor pi0150 n13756 ; n13763
g11328 and n13762_not n13763 ; n13764
g11329 and pi0299 n13764_not ; n13765
g11330 and n13751_not n13765 ; n13766
g11331 nor n9506 n13741 ; n13767
g11332 nor pi0173 n13767 ; n13768
g11333 and pi0173 n13759 ; n13769
g11334 nor pi0185 n13768 ; n13770
g11335 and n13769_not n13770 ; n13771
g11336 and n6197 n9391_not ; n13772
g11337 and pi0173 n13736_not ; n13773
g11338 and n13772_not n13773 ; n13774
g11339 nor n9496 n13741 ; n13775
g11340 nor pi0173 n13775 ; n13776
g11341 and pi0185 n13774_not ; n13777
g11342 and n13776_not n13777 ; n13778
g11343 and pi0190 n13771_not ; n13779
g11344 and n13778_not n13779 ; n13780
g11345 nor pi0173 n9527 ; n13781
g11346 and pi0173 n9949_not ; n13782
g11347 and n6197 n13781_not ; n13783
g11348 and n13782_not n13783 ; n13784
g11349 and pi0185 n13741_not ; n13785
g11350 and n13784_not n13785 ; n13786
g11351 and pi0173 n13757 ; n13787
g11352 and pi0173_not n9532 ; n13788
g11353 nor pi0185 n13788 ; n13789
g11354 and n13787_not n13789 ; n13790
g11355 nor pi0190 n13790 ; n13791
g11356 and n13786_not n13791 ; n13792
g11357 nor pi0299 n13792 ; n13793
g11358 and n13780_not n13793 ; n13794
g11359 and pi0232 n13794_not ; n13795
g11360 and n13766_not n13795 ; n13796
g11361 nor pi0039 n13735 ; n13797
g11362 and n13796_not n13797 ; n13798
g11363 and pi0168 n9311 ; n13799
g11364 and pi0157 n9324 ; n13800
g11365 nor n13799 n13800 ; n13801
g11366 and n6197 n11747 ; n13802
g11367 and n13801_not n13802 ; n13803
g11368 and pi0299 n13803_not ; n13804
g11369 nor n13718 n13804 ; n13805
g11370 and n9248 n13805_not ; n13806
g11371 and pi0178 n9338_not ; n13807
g11372 nor pi0190 n13807 ; n13808
g11373 nor pi0299 n13808 ; n13809
g11374 nor n13806 n13809 ; n13810
g11375 and n6205 n9248_not ; n13811
g11376 and n9051 n13811_not ; n13812
g11377 and pi0178_not n13812 ; n13813
g11378 and n9314_not n13813 ; n13814
g11379 nor pi0299 n9303 ; n13815
g11380 and pi0178 n13812 ; n13816
g11381 and n9305_not n13816 ; n13817
g11382 and pi0190 n13815 ; n13818
g11383 and n13814_not n13818 ; n13819
g11384 and n13817_not n13819 ; n13820
g11385 and pi0232 n13820_not ; n13821
g11386 and n13810_not n13821 ; n13822
g11387 and pi0232_not n9248 ; n13823
g11388 and pi0039 n13823_not ; n13824
g11389 and n13822_not n13824 ; n13825
g11390 nor pi0038 n13825 ; n13826
g11391 and n13798_not n13826 ; n13827
g11392 and n13734 n13827_not ; n13828
g11393 and n8161 n13715_not ; n13829
g11394 and n9249_not n13829 ; n13830
g11395 nor n13714 n13830 ; n13831
g11396 and n13828_not n13831 ; n13832
g11397 and n2569 n13832_not ; n13833
g11398 nor n13713 n13725 ; n13834
g11399 and n13833_not n13834 ; n13835
g11400 nor pi0054 n13835 ; n13836
g11401 nor n13712 n13836 ; n13837
g11402 nor pi0074 n13837 ; n13838
g11403 and n13705 n13838_not ; n13839
g11404 and n2529 n13693_not ; n13840
g11405 and n13839_not n13840 ; n13841
g11406 nor n13683 n13841 ; n13842
g11407 and n8989 n13674 ; n13843
g11408 nor n8989 n13671 ; n13844
g11409 nor n3328 n13843 ; n13845
g11410 and n13844_not n13845 ; n13846
g11411 and n13673_not n13846 ; n13847
g11412 nor n13842 n13847 ; n13848
g11413 and pi0118 n13848 ; n13849
g11414 and n8965 n13720_not ; n13850
g11415 and n2521 n13850 ; n13851
g11416 and n13716 n13851_not ; n13852
g11417 nor n13714 n13852 ; n13853
g11418 and n9205 n13853_not ; n13854
g11419 and n7309 n9061 ; n13855
g11420 and n6244_not n13130 ; n13856
g11421 and n6392_not n13856 ; n13857
g11422 nor pi0232 n13857 ; n13858
g11423 and n13855_not n13858 ; n13859
g11424 and n6198 n6392_not ; n13860
g11425 and pi0157 n9039_not ; n13861
g11426 and pi0157_not n9044 ; n13862
g11427 and pi0168 n13862_not ; n13863
g11428 nor pi0157 pi0168 ; n13864
g11429 and n9037_not n13864 ; n13865
g11430 nor n13861 n13865 ; n13866
g11431 and n13863_not n13866 ; n13867
g11432 nor n13860 n13867 ; n13868
g11433 and n13130 n13868_not ; n13869
g11434 nor pi0178 n6205 ; n13870
g11435 and n9043 n13870 ; n13871
g11436 nor n13860 n13871 ; n13872
g11437 and pi0190 n13872_not ; n13873
g11438 and pi0178 n9052_not ; n13874
g11439 and n13860_not n13874 ; n13875
g11440 nor pi0178 n13173 ; n13876
g11441 nor pi0190 n13875 ; n13877
g11442 and n13876_not n13877 ; n13878
g11443 nor n13873 n13878 ; n13879
g11444 and n13132 n13879_not ; n13880
g11445 and pi0232 n13880_not ; n13881
g11446 and n13869_not n13881 ; n13882
g11447 and pi0039 n13859_not ; n13883
g11448 and n13882_not n13883 ; n13884
g11449 nor n6169 n9120 ; n13885
g11450 nor pi0232 n9118 ; n13886
g11451 and n13885_not n13886 ; n13887
g11452 nor n9118 n11798 ; n13888
g11453 nor n6197 n13888 ; n13889
g11454 and n9142 n13742 ; n13890
g11455 and pi0168 n9133_not ; n13891
g11456 nor pi0168 n9092 ; n13892
g11457 nor pi0151 n13891 ; n13893
g11458 and n13892_not n13893 ; n13894
g11459 nor n13890 n13894 ; n13895
g11460 and n9094 n13895_not ; n13896
g11461 and pi0150 n13896_not ; n13897
g11462 and pi0151_not n9129 ; n13898
g11463 and n9166 n13898_not ; n13899
g11464 and n13752 n13899_not ; n13900
g11465 and pi0151_not n9118 ; n13901
g11466 and n9162 n13901_not ; n13902
g11467 nor pi0168 n13902 ; n13903
g11468 nor pi0150 n13900 ; n13904
g11469 and n13903_not n13904 ; n13905
g11470 nor n13897 n13905 ; n13906
g11471 and pi0299 n13889_not ; n13907
g11472 and n13906_not n13907 ; n13908
g11473 nor n6197 n9122 ; n13909
g11474 and n6479 n9142 ; n13910
g11475 and pi0173 n13910 ; n13911
g11476 and pi0173_not n6479 ; n13912
g11477 and n9092 n13912 ; n13913
g11478 nor n13911 n13913 ; n13914
g11479 and pi0190_not n6197 ; n13915
g11480 and n13914_not n13915 ; n13916
g11481 and pi0173_not pi0190 ; n13917
g11482 and n9134 n13917 ; n13918
g11483 and pi0185 n13918_not ; n13919
g11484 and n13916_not n13919 ; n13920
g11485 and pi0173 n9150 ; n13921
g11486 and pi0190 n9131 ; n13922
g11487 and n13921_not n13922 ; n13923
g11488 and pi0173_not n9118 ; n13924
g11489 and n9147 n13924_not ; n13925
g11490 nor pi0190 n13925 ; n13926
g11491 nor pi0185 n13923 ; n13927
g11492 and n13926_not n13927 ; n13928
g11493 nor n13920 n13928 ; n13929
g11494 nor pi0299 n13909 ; n13930
g11495 and n13929_not n13930 ; n13931
g11496 nor n13908 n13931 ; n13932
g11497 and pi0232 n13932_not ; n13933
g11498 nor pi0039 n13887 ; n13934
g11499 and n13933_not n13934 ; n13935
g11500 nor n13884 n13935 ; n13936
g11501 nor pi0038 n13936 ; n13937
g11502 and n13734 n13937_not ; n13938
g11503 nor n13714 n13829 ; n13939
g11504 and n13938_not n13939 ; n13940
g11505 and n2569 n13940_not ; n13941
g11506 nor n13713 n13854 ; n13942
g11507 and n13941_not n13942 ; n13943
g11508 nor pi0054 n13943 ; n13944
g11509 nor n13712 n13944 ; n13945
g11510 nor pi0074 n13945 ; n13946
g11511 and n13705 n13946_not ; n13947
g11512 and pi0054 n13674 ; n13948
g11513 and pi0092_not n8989 ; n13949
g11514 and n8965 n13949 ; n13950
g11515 and n13685_not n13950 ; n13951
g11516 and n13948_not n13951 ; n13952
g11517 and n2521 n13952 ; n13953
g11518 and n13679 n13953_not ; n13954
g11519 and n13684 n13954_not ; n13955
g11520 and n2529 n13955_not ; n13956
g11521 and n13947_not n13956 ; n13957
g11522 and n13682 n13957_not ; n13958
g11523 nor n13847 n13958 ; n13959
g11524 and pi0118_not n13959 ; n13960
g11525 nor n13664 n13960 ; n13961
g11526 and n13849_not n13961 ; n13962
g11527 nor pi0118 n8976 ; n13963
g11528 and n13959 n13963_not ; n13964
g11529 and n13848 n13963 ; n13965
g11530 and n13664 n13964_not ; n13966
g11531 and n13965_not n13966 ; n13967
g11532 or n13962 n13967 ; po0276
g11533 and pi0128 pi0228 ; n13969
g11534 and n10163_not n13969 ; n13970
g11535 and n7384 n8965 ; n13971
g11536 nor n13969 n13971 ; n13972
g11537 and pi0075 n13972_not ; n13973
g11538 and pi0087 n13969_not ; n13974
g11539 and n2530 n3335 ; n13975
g11540 nor n13969 n13975 ; n13976
g11541 and pi0100 n13976_not ; n13977
g11542 and n2603_not n3470 ; n13978
g11543 and n7606 n13978 ; n13979
g11544 and n3448_not n5853 ; n13980
g11545 and n7603 n13980 ; n13981
g11546 nor n13979 n13981 ; n13982
g11547 and pi0039 n13982_not ; n13983
g11548 and pi0299 n6418 ; n13984
g11549 nor n6528 n13984 ; n13985
g11550 and n7473 n13985_not ; n13986
g11551 and pi0109 n13986_not ; n13987
g11552 and n2928_not n11668 ; n13988
g11553 and n2770 n10157 ; n13989
g11554 and n11667 n13989_not ; n13990
g11555 and n2783 n13990_not ; n13991
g11556 nor pi0097 n13991 ; n13992
g11557 and pi0046_not n2928 ; n13993
g11558 and n2936 n13993 ; n13994
g11559 and n13992_not n13994 ; n13995
g11560 nor n13987 n13988 ; n13996
g11561 and n13995_not n13996 ; n13997
g11562 nor n6422 n13986 ; n13998
g11563 and n6491_not n13986 ; n13999
g11564 nor n13998 n13999 ; n14000
g11565 and n13997_not n14000 ; n14001
g11566 nor pi0091 n14001 ; n14002
g11567 and n2938 n6419_not ; n14003
g11568 and n14002_not n14003 ; n14004
g11569 nor n2752 n14004 ; n14005
g11570 and pi0039_not n11086 ; n14006
g11571 and n14005_not n14006 ; n14007
g11572 nor n13983 n14007 ; n14008
g11573 nor pi0038 n14008 ; n14009
g11574 and pi0228_not n14009 ; n14010
g11575 nor n13969 n14010 ; n14011
g11576 nor pi0100 n14011 ; n14012
g11577 nor pi0087 n13977 ; n14013
g11578 and n14012_not n14013 ; n14014
g11579 nor pi0075 n13974 ; n14015
g11580 and n14014_not n14015 ; n14016
g11581 nor pi0092 n13973 ; n14017
g11582 and n14016_not n14017 ; n14018
g11583 and pi0092 n13969_not ; n14019
g11584 and n7369_not n14019 ; n14020
g11585 and n10163 n14020_not ; n14021
g11586 and n14018_not n14021 ; n14022
g11587 or n13970 n14022 ; po0277
g11588 nor pi0031 pi0080 ; n14024
g11589 and pi0818 n14024 ; n14025
g11590 and n7420 n7429_not ; n14026
g11591 nor n7425 n14026 ; n14027
g11592 nor pi0120 n7429 ; n14028
g11593 and pi1093_not n14028 ; n14029
g11594 and n14027 n14029_not ; n14030
g11595 and pi0120 n7420_not ; n14031
g11596 and pi0120_not pi1093 ; n14032
g11597 and pi1091_not n12310 ; n14033
g11598 and n14032 n14033_not ; n14034
g11599 nor n14031 n14034 ; n14035
g11600 and n2521 n7595 ; n14036
g11601 and n7619_not n14031 ; n14037
g11602 and n14036 n14037_not ; n14038
g11603 and n7619 n14032_not ; n14039
g11604 nor n14038 n14039 ; n14040
g11605 and n2530 n7506 ; n14041
g11606 and n14040_not n14041 ; n14042
g11607 and pi0100 n14035_not ; n14043
g11608 and n14042_not n14043 ; n14044
g11609 and pi0038 n7420 ; n14045
g11610 and pi1093_not n7460 ; n14046
g11611 and pi0120 n14046 ; n14047
g11612 nor pi0039 n14047 ; n14048
g11613 and pi0122 n7452_not ; n14049
g11614 and n7534 n10445_not ; n14050
g11615 and n7417 n7451 ; n14051
g11616 and pi0829_not n14051 ; n14052
g11617 nor pi0122 n14052 ; n14053
g11618 and n14050_not n14053 ; n14054
g11619 nor n2923 n14049 ; n14055
g11620 and n14054_not n14055 ; n14056
g11621 and n2930 n14056_not ; n14057
g11622 and n7626 n14051_not ; n14058
g11623 and n12310_not n14058 ; n14059
g11624 nor n14057 n14059 ; n14060
g11625 and n14048 n14060 ; n14061
g11626 and n7570_not n14035 ; n14062
g11627 and n6198_not n14035 ; n14063
g11628 and n7602_not n14031 ; n14064
g11629 and pi1091 pi1092 ; n14065
g11630 and n7554 n14065 ; n14066
g11631 and n14034 n14066_not ; n14067
g11632 nor n14064 n14067 ; n14068
g11633 and n6198 n14068 ; n14069
g11634 nor n14063 n14069 ; n14070
g11635 and n6242 n14070 ; n14071
g11636 and n6227 n14035_not ; n14072
g11637 nor n6227 n14068 ; n14073
g11638 nor n14072 n14073 ; n14074
g11639 nor n6242 n14074 ; n14075
g11640 and n7570 n14071_not ; n14076
g11641 and n14075_not n14076 ; n14077
g11642 and pi0299 n14062_not ; n14078
g11643 and n14077_not n14078 ; n14079
g11644 and n6205 n14070 ; n14080
g11645 nor n6205 n14074 ; n14081
g11646 and n7551 n14080_not ; n14082
g11647 and n14081_not n14082 ; n14083
g11648 and n7551_not n14035 ; n14084
g11649 nor pi0299 n14084 ; n14085
g11650 and n14083_not n14085 ; n14086
g11651 and pi0039 n14079_not ; n14087
g11652 and n14086_not n14087 ; n14088
g11653 nor n14061 n14088 ; n14089
g11654 nor pi0038 n14089 ; n14090
g11655 nor pi0120 pi1093 ; n14091
g11656 and pi0038 n14091 ; n14092
g11657 nor pi0100 n14092 ; n14093
g11658 and n14045_not n14093 ; n14094
g11659 and n14090_not n14094 ; n14095
g11660 nor n14044 n14095 ; n14096
g11661 nor pi0087 n14096 ; n14097
g11662 and n7631 n14091_not ; n14098
g11663 and n2625_not n7420 ; n14099
g11664 and n7626 n12310_not ; n14100
g11665 and n7496_not n14100 ; n14101
g11666 and n7629 n14101_not ; n14102
g11667 and pi0087 n14099_not ; n14103
g11668 and n14102_not n14103 ; n14104
g11669 and n14098 n14104 ; n14105
g11670 nor n14097 n14105 ; n14106
g11671 nor pi0075 n14106 ; n14107
g11672 and n7474 n14035 ; n14108
g11673 and n7596_not n14034 ; n14109
g11674 nor pi1091 n7419 ; n14110
g11675 nor n7482 n14110 ; n14111
g11676 and pi0120 n14111_not ; n14112
g11677 nor n7474 n14112 ; n14113
g11678 and n14109_not n14113 ; n14114
g11679 nor n14108 n14114 ; n14115
g11680 and n2610 n14115_not ; n14116
g11681 and n2610_not n14035 ; n14117
g11682 and pi0075 n14117_not ; n14118
g11683 and n14116_not n14118 ; n14119
g11684 and n7429 n14119_not ; n14120
g11685 and n14107_not n14120 ; n14121
g11686 and n14030 n14121_not ; n14122
g11687 and n7599 n14091_not ; n14123
g11688 nor n14057 n14058 ; n14124
g11689 and n14048 n14124 ; n14125
g11690 and pi1093 n6198_not ; n14126
g11691 and n6242 n14126 ; n14127
g11692 and n6227 n6242_not ; n14128
g11693 and n7570 n14128_not ; n14129
g11694 and n14127_not n14129 ; n14130
g11695 and n7602 n14130 ; n14131
g11696 and pi0299 n14091_not ; n14132
g11697 and n14131_not n14132 ; n14133
g11698 and n6205 n14126 ; n14134
g11699 and n6205_not n6227 ; n14135
g11700 and n7551 n14135_not ; n14136
g11701 and n14134_not n14136 ; n14137
g11702 and n7602 n14137 ; n14138
g11703 nor pi0299 n14091 ; n14139
g11704 and n14138_not n14139 ; n14140
g11705 and pi0039 n14133_not ; n14141
g11706 and n14140_not n14141 ; n14142
g11707 nor n14125 n14142 ; n14143
g11708 nor pi0038 n14143 ; n14144
g11709 and n14093 n14144_not ; n14145
g11710 and pi0120 n7619 ; n14146
g11711 and pi0120_not n14036 ; n14147
g11712 nor n14146 n14147 ; n14148
g11713 and n14041 n14148_not ; n14149
g11714 and pi0100 n14091_not ; n14150
g11715 and n14149_not n14150 ; n14151
g11716 nor n14145 n14151 ; n14152
g11717 nor pi0087 n14152 ; n14153
g11718 nor n14098 n14153 ; n14154
g11719 nor pi0075 n14154 ; n14155
g11720 and n7429 n14123_not ; n14156
g11721 and n14155_not n14156 ; n14157
g11722 and n7425 n14029_not ; n14158
g11723 and n14157_not n14158 ; n14159
g11724 nor n14122 n14159 ; n14160
g11725 and n14025 n14160_not ; n14161
g11726 nor po1038 n14161 ; n14162
g11727 and n7425_not n14035 ; n14163
g11728 and pi0120 n14163_not ; n14164
g11729 and n14025 n14091_not ; n14165
g11730 and n14163_not n14165 ; n14166
g11731 and po1038 n14166_not ; n14167
g11732 and n14164_not n14167 ; n14168
g11733 nor n7643 n14168 ; n14169
g11734 and pi0951 pi0982 ; n14170
g11735 and pi1092 n14170 ; n14171
g11736 and pi1093 n14171 ; n14172
g11737 nor pi0120 n14172 ; n14173
g11738 nor n14163 n14173 ; n14174
g11739 and n14167 n14174_not ; n14175
g11740 and n7643 n14175_not ; n14176
g11741 nor n14169 n14176 ; n14177
g11742 nor n14162 n14177 ; n14178
g11743 and n14028 n14172_not ; n14179
g11744 nor n2610 n14173 ; n14180
g11745 and pi0120 n7597 ; n14181
g11746 and pi1091_not n14172 ; n14182
g11747 nor pi0120 n14182 ; n14183
g11748 and n2930 n14171 ; n14184
g11749 nor pi0093 pi0122 ; n14185
g11750 and n2506 n14185 ; n14186
g11751 and n2925 n8894 ; n14187
g11752 and n14186 n14187 ; n14188
g11753 and n2962 n14188 ; n14189
g11754 and n10324 n14189 ; n14190
g11755 and n7478 n14190 ; n14191
g11756 and n2703 n14191 ; n14192
g11757 and n14184 n14192_not ; n14193
g11758 and n14183 n14193_not ; n14194
g11759 nor n14181 n14194 ; n14195
g11760 nor n7474 n14195 ; n14196
g11761 and n7474 n14173 ; n14197
g11762 and n2610 n14197_not ; n14198
g11763 and n14196_not n14198 ; n14199
g11764 and pi0075 n14180_not ; n14200
g11765 and n14199_not n14200 ; n14201
g11766 and n2625_not n14173 ; n14202
g11767 and pi0087 n14202_not ; n14203
g11768 and pi0950 n2521 ; n14204
g11769 nor n2923 n6213 ; n14205
g11770 and n14204 n14205 ; n14206
g11771 and n14184 n14206_not ; n14207
g11772 and pi0824 n14204 ; n14208
g11773 and n14182 n14208_not ; n14209
g11774 nor n14207 n14209 ; n14210
g11775 nor pi0120 n14210 ; n14211
g11776 nor n7627 n7628 ; n14212
g11777 and pi0120 n14212_not ; n14213
g11778 and n2625 n14213_not ; n14214
g11779 and n14211_not n14214 ; n14215
g11780 and n14203 n14215_not ; n14216
g11781 and n7430 n7478 ; n14217
g11782 and n14204 n14217 ; n14218
g11783 and n14184 n14218_not ; n14219
g11784 and n14183 n14219_not ; n14220
g11785 nor n14146 n14220 ; n14221
g11786 and pi0039_not n7506 ; n14222
g11787 and n14221_not n14222 ; n14223
g11788 and pi0100 n14223_not ; n14224
g11789 nor pi0038 n14224 ; n14225
g11790 and n14041_not n14173 ; n14226
g11791 nor n14225 n14226 ; n14227
g11792 and n7551_not n14173 ; n14228
g11793 nor pi0299 n14228 ; n14229
g11794 nor n8621 n14173 ; n14230
g11795 and n6205_not n14230 ; n14231
g11796 nor n8624 n14173 ; n14232
g11797 and n6205 n14232 ; n14233
g11798 and n7551 n14231_not ; n14234
g11799 and n14233_not n14234 ; n14235
g11800 and n14229 n14235_not ; n14236
g11801 and n7570_not n14173 ; n14237
g11802 and pi0299 n14237_not ; n14238
g11803 and n6242_not n14230 ; n14239
g11804 and n6242 n14232 ; n14240
g11805 and n7570 n14239_not ; n14241
g11806 and n14240_not n14241 ; n14242
g11807 and n14238 n14242_not ; n14243
g11808 nor n14236 n14243 ; n14244
g11809 and pi0039 n14244_not ; n14245
g11810 and n2771 n7437 ; n14246
g11811 and n2767 n14246 ; n14247
g11812 and n9110 n14247 ; n14248
g11813 and n7431 n14248 ; n14249
g11814 and n7436 n14249_not ; n14250
g11815 and pi0950 n7518 ; n14251
g11816 and n14250_not n14251 ; n14252
g11817 and pi0824 n14252 ; n14253
g11818 and n14171 n14253_not ; n14254
g11819 and pi0829_not n14254 ; n14255
g11820 nor pi0097 n14247 ; n14256
g11821 and n2935 n14256_not ; n14257
g11822 and n2937 n14257 ; n14258
g11823 nor n7522 n14258 ; n14259
g11824 and n2461 n14259_not ; n14260
g11825 and n7434 n14260_not ; n14261
g11826 and n7431 n14261_not ; n14262
g11827 nor pi0051 n14262 ; n14263
g11828 nor n2747 n14263 ; n14264
g11829 nor pi0096 n14264 ; n14265
g11830 and pi0072_not pi0950 ; n14266
g11831 and n10416 n14266 ; n14267
g11832 and n14265_not n14267 ; n14268
g11833 and n7430 n14171 ; n14269
g11834 and n14268_not n14269 ; n14270
g11835 and pi0829 pi1092 ; n14271
g11836 and pi0122 n14170 ; n14272
g11837 and n14271 n14272 ; n14273
g11838 and n14252_not n14273 ; n14274
g11839 nor n14255 n14274 ; n14275
g11840 and n14270_not n14275 ; n14276
g11841 and n7517 n14276_not ; n14277
g11842 and n2923 n14172 ; n14278
g11843 nor n14277 n14278 ; n14279
g11844 and pi1091 n14279_not ; n14280
g11845 and n14182 n14253_not ; n14281
g11846 nor pi0120 n14281 ; n14282
g11847 and n14280_not n14282 ; n14283
g11848 and n14046_not n14124 ; n14284
g11849 and pi0120 n14284 ; n14285
g11850 nor pi0039 n14283 ; n14286
g11851 and n14285_not n14286 ; n14287
g11852 nor n14245 n14287 ; n14288
g11853 and n2608 n14288_not ; n14289
g11854 nor n14227 n14289 ; n14290
g11855 nor pi0087 n14290 ; n14291
g11856 nor pi0075 n14216 ; n14292
g11857 and n14291_not n14292 ; n14293
g11858 nor n14201 n14293 ; n14294
g11859 and n7429 n14294_not ; n14295
g11860 and n7425 n14295_not ; n14296
g11861 nor n14035 n14173 ; n14297
g11862 nor n2530 n14297 ; n14298
g11863 and n7506_not n14297 ; n14299
g11864 and n12310_not n14182 ; n14300
g11865 nor n14219 n14300 ; n14301
g11866 nor pi0120 n14301 ; n14302
g11867 nor n14037 n14302 ; n14303
g11868 and n7506 n14303_not ; n14304
g11869 and n2530 n14299_not ; n14305
g11870 and n14304_not n14305 ; n14306
g11871 and pi0100 n14298_not ; n14307
g11872 and n14306_not n14307 ; n14308
g11873 and pi0038 n14297_not ; n14309
g11874 and n14046_not n14060 ; n14310
g11875 and pi0120 n14310 ; n14311
g11876 and n14100 n14254 ; n14312
g11877 nor pi0120 n14312 ; n14313
g11878 and n14280_not n14313 ; n14314
g11879 nor n14311 n14314 ; n14315
g11880 nor pi0039 n14315 ; n14316
g11881 and n7554_not n14184 ; n14317
g11882 nor n14300 n14317 ; n14318
g11883 nor pi0120 n14318 ; n14319
g11884 nor n14064 n14319 ; n14320
g11885 and n6198 n14320_not ; n14321
g11886 and n6198_not n14297 ; n14322
g11887 nor n14321 n14322 ; n14323
g11888 and n6205 n14323_not ; n14324
g11889 nor n6227 n14320 ; n14325
g11890 and n6227 n14297 ; n14326
g11891 nor n14325 n14326 ; n14327
g11892 nor n6205 n14327 ; n14328
g11893 and n7551 n14324_not ; n14329
g11894 and n14328_not n14329 ; n14330
g11895 and n14084_not n14229 ; n14331
g11896 and n14330_not n14331 ; n14332
g11897 and n6242 n14323_not ; n14333
g11898 nor n6242 n14327 ; n14334
g11899 and n7570 n14333_not ; n14335
g11900 and n14334_not n14335 ; n14336
g11901 and n7420 n7570_not ; n14337
g11902 and n14238 n14337_not ; n14338
g11903 and n14336_not n14338 ; n14339
g11904 and pi0039 n14332_not ; n14340
g11905 and n14339_not n14340 ; n14341
g11906 nor n14316 n14341 ; n14342
g11907 nor pi0038 n14342 ; n14343
g11908 nor pi0100 n14309 ; n14344
g11909 and n14343_not n14344 ; n14345
g11910 nor n14308 n14345 ; n14346
g11911 nor pi0087 n14346 ; n14347
g11912 nor n14102 n14214 ; n14348
g11913 nor n14207 n14300 ; n14349
g11914 and n14211 n14349_not ; n14350
g11915 nor n14348 n14350 ; n14351
g11916 and n14099_not n14203 ; n14352
g11917 and n14351_not n14352 ; n14353
g11918 nor n14347 n14353 ; n14354
g11919 nor pi0075 n14354 ; n14355
g11920 and n7474 n14297_not ; n14356
g11921 nor n14193 n14300 ; n14357
g11922 nor pi0120 n14357 ; n14358
g11923 and n14113 n14358_not ; n14359
g11924 nor n14356 n14359 ; n14360
g11925 and n2610 n14360_not ; n14361
g11926 nor n2610 n14297 ; n14362
g11927 and pi0075 n14362_not ; n14363
g11928 and n14361_not n14363 ; n14364
g11929 and n7429 n14364_not ; n14365
g11930 and n14355_not n14365 ; n14366
g11931 and n14030 n14366_not ; n14367
g11932 nor n14296 n14367 ; n14368
g11933 and n14176 n14179_not ; n14369
g11934 and n14368_not n14369 ; n14370
g11935 and n7420_not n7623 ; n14371
g11936 nor pi0039 n14310 ; n14372
g11937 and n7420 n7551_not ; n14373
g11938 nor n7556 n14110 ; n14374
g11939 and n6198 n14374_not ; n14375
g11940 nor n6198 n7420 ; n14376
g11941 nor n14375 n14376 ; n14377
g11942 and n6205 n14377_not ; n14378
g11943 nor n6227 n14374 ; n14379
g11944 and n6227 n7420_not ; n14380
g11945 nor n14379 n14380 ; n14381
g11946 nor n6205 n14381 ; n14382
g11947 and n7551 n14378_not ; n14383
g11948 and n14382_not n14383 ; n14384
g11949 nor pi0299 n14373 ; n14385
g11950 and n14384_not n14385 ; n14386
g11951 and n6242 n14377_not ; n14387
g11952 nor n6242 n14381 ; n14388
g11953 and n7570 n14387_not ; n14389
g11954 and n14388_not n14389 ; n14390
g11955 and pi0299 n14337_not ; n14391
g11956 and n14390_not n14391 ; n14392
g11957 nor n14386 n14392 ; n14393
g11958 and pi0039 n14393_not ; n14394
g11959 nor pi0038 n14394 ; n14395
g11960 and n14372_not n14395 ; n14396
g11961 nor pi0100 n14045 ; n14397
g11962 and n14396_not n14397 ; n14398
g11963 nor n14371 n14398 ; n14399
g11964 nor pi0087 n14399 ; n14400
g11965 nor n14104 n14400 ; n14401
g11966 nor pi0075 n14401 ; n14402
g11967 and n7420 n7475_not ; n14403
g11968 and n7475 n14111 ; n14404
g11969 and pi0075 n14403_not ; n14405
g11970 and n14404_not n14405 ; n14406
g11971 nor n14402 n14406 ; n14407
g11972 and n14027 n14407_not ; n14408
g11973 nor n7429 n14163 ; n14409
g11974 nor pi0039 n14284 ; n14410
g11975 and n7612 n14410_not ; n14411
g11976 nor pi0100 n14411 ; n14412
g11977 nor n7623 n14412 ; n14413
g11978 nor pi0087 n14413 ; n14414
g11979 nor n7631 n14414 ; n14415
g11980 nor pi0075 n14415 ; n14416
g11981 nor n7599 n14416 ; n14417
g11982 and n7425 n14028_not ; n14418
g11983 and n14417_not n14418 ; n14419
g11984 nor n14408 n14409 ; n14420
g11985 and n14419_not n14420 ; n14421
g11986 and pi0120 n14169 ; n14422
g11987 and n14421_not n14422 ; n14423
g11988 nor n14370 n14423 ; n14424
g11989 nor n14025 n14424 ; n14425
g11990 or n14178 n14425 ; po0278
g11991 nor pi0134 pi0135 ; n14427
g11992 and pi0136_not n14427 ; n14428
g11993 and pi0130_not n14428 ; n14429
g11994 and pi0132_not n14429 ; n14430
g11995 and pi0126_not n14430 ; n14431
g11996 and pi0121_not n14431 ; n14432
g11997 nor pi0125 pi0133 ; n14433
g11998 and pi0121 n14433_not ; n14434
g11999 and pi0121_not n14433 ; n14435
g12000 nor n14434 n14435 ; n14436
g12001 nor n14432 n14436 ; n14437
g12002 and n2478 n10152 ; n14438
g12003 and pi0051_not n14438 ; n14439
g12004 and pi0087_not n14439 ; n14440
g12005 and n14437_not n14440 ; n14441
g12006 and pi0051 pi0146 ; n14442
g12007 and pi0051 n6197 ; n14443
g12008 and pi0146_not n14443 ; n14444
g12009 and pi0161 n14444_not ; n14445
g12010 and n6197 n14439_not ; n14446
g12011 nor n14442 n14445 ; n14447
g12012 and n14446 n14447 ; n14448
g12013 nor pi0087 n14448 ; n14449
g12014 and pi0087 n13665_not ; n14450
g12015 and pi0232 n14450_not ; n14451
g12016 and n14449_not n14451 ; n14452
g12017 and po1038 n14441_not ; n14453
g12018 and n14452_not n14453 ; n14454
g12019 nor pi0087 n2570 ; n14455
g12020 and n14439_not n14455 ; n14456
g12021 and pi0142_not n14443 ; n14457
g12022 and pi0144 n14457_not ; n14458
g12023 and pi0051 pi0142 ; n14459
g12024 and n14446 n14459_not ; n14460
g12025 and n14458_not n14460 ; n14461
g12026 nor pi0299 n14461 ; n14462
g12027 and pi0299 n14448_not ; n14463
g12028 and pi0232 n14462_not ; n14464
g12029 and n14463_not n14464 ; n14465
g12030 and n14456 n14465_not ; n14466
g12031 and pi0100 n14439 ; n14467
g12032 and n2535 n14467_not ; n14468
g12033 and pi0100 n14465 ; n14469
g12034 and pi0038 n14465_not ; n14470
g12035 nor pi0100 n14470 ; n14471
g12036 and pi0038 n14439_not ; n14472
g12037 nor pi0100 n14472 ; n14473
g12038 nor n14471 n14473 ; n14474
g12039 nor pi0161 n14444 ; n14475
g12040 and n2705 n7445 ; n14476
g12041 and pi0024_not pi0314 ; n14477
g12042 and n14476 n14477 ; n14478
g12043 and n2467 n10151 ; n14479
g12044 and n13047 n14479 ; n14480
g12045 and pi0050_not pi0077 ; n14481
g12046 and n2495 n14481 ; n14482
g12047 and n14480 n14482 ; n14483
g12048 and n8897 n14478 ; n14484
g12049 and n14483 n14484 ; n14485
g12050 and n2519 n14485 ; n14486
g12051 and n2770 n14480 ; n14487
g12052 and pi0058_not n14476 ; n14488
g12053 and n9253 n14488 ; n14489
g12054 and n14487 n14489 ; n14490
g12055 and pi0072 n6479 ; n14491
g12056 and n14490 n14491 ; n14492
g12057 and n14438 n14476_not ; n14493
g12058 nor pi0051 n14493 ; n14494
g12059 and pi0024_not n11663 ; n14495
g12060 and n14487 n14495 ; n14496
g12061 and pi0086 n14487 ; n14497
g12062 nor n14483 n14497 ; n14498
g12063 and n11076 n14498_not ; n14499
g12064 and n14438 n14496_not ; n14500
g12065 and n14499_not n14500 ; n14501
g12066 and n14494 n14501_not ; n14502
g12067 and n2519 n14502 ; n14503
g12068 and n14439 n14503_not ; n14504
g12069 and n14492_not n14504 ; n14505
g12070 and n14486_not n14505 ; n14506
g12071 nor n6197 n14506 ; n14507
g12072 and pi0072 n10342 ; n14508
g12073 nor n14443 n14508 ; n14509
g12074 and n6197 n14509_not ; n14510
g12075 nor n14507 n14510 ; n14511
g12076 and n14475 n14511_not ; n14512
g12077 and n14439 n14486_not ; n14513
g12078 and n14503_not n14513 ; n14514
g12079 nor n6197 n14514 ; n14515
g12080 nor n14446 n14515 ; n14516
g12081 and n14492_not n14516 ; n14517
g12082 and pi0146 n14517 ; n14518
g12083 and pi0051_not n6197 ; n14519
g12084 and n14438 n14492_not ; n14520
g12085 and n14519 n14520_not ; n14521
g12086 nor pi0146 n14521 ; n14522
g12087 and n14507_not n14522 ; n14523
g12088 and pi0161 n14518_not ; n14524
g12089 and n14523_not n14524 ; n14525
g12090 nor n14512 n14525 ; n14526
g12091 and n9572 n14526_not ; n14527
g12092 and n6197_not n14506 ; n14528
g12093 and pi0051_not n14478 ; n14529
g12094 and n13439 n14529 ; n14530
g12095 nor pi0072 n14530 ; n14531
g12096 and n6480 n14531_not ; n14532
g12097 and n6197 n14532_not ; n14533
g12098 nor n14528 n14533 ; n14534
g12099 nor pi0146 n14534 ; n14535
g12100 and n2519 n6197 ; n14536
g12101 and n14530 n14536 ; n14537
g12102 and n14511 n14537_not ; n14538
g12103 and pi0146 n14538 ; n14539
g12104 nor pi0161 n14535 ; n14540
g12105 and n14539_not n14540 ; n14541
g12106 and n14519 n14520 ; n14542
g12107 and n14486_not n14542 ; n14543
g12108 nor n14443 n14543 ; n14544
g12109 and pi0146 n14439_not ; n14545
g12110 nor n14544 n14545 ; n14546
g12111 and pi0161 n14546_not ; n14547
g12112 and n14528_not n14547 ; n14548
g12113 nor n14541 n14548 ; n14549
g12114 and n9603 n14549_not ; n14550
g12115 nor n14527 n14550 ; n14551
g12116 and pi0156 n14551_not ; n14552
g12117 and pi0144 n14517_not ; n14553
g12118 nor pi0144 n14511 ; n14554
g12119 nor n14553 n14554 ; n14555
g12120 nor n14457 n14555 ; n14556
g12121 and pi0180 n14556_not ; n14557
g12122 nor pi0142 n14534 ; n14558
g12123 and pi0142 n14538 ; n14559
g12124 nor pi0144 n14558 ; n14560
g12125 and n14559_not n14560 ; n14561
g12126 and n14486_not n14517 ; n14562
g12127 and n14458 n14562_not ; n14563
g12128 nor pi0180 n14563 ; n14564
g12129 and n14561_not n14564 ; n14565
g12130 and pi0179 n14557_not ; n14566
g12131 and n14565_not n14566 ; n14567
g12132 and n14458 n14506_not ; n14568
g12133 nor pi0024 n11664 ; n14569
g12134 and pi0024 n11669_not ; n14570
g12135 nor n14569 n14570 ; n14571
g12136 nor pi0314 n14571 ; n14572
g12137 and pi0314 n11669_not ; n14573
g12138 nor n14572 n14573 ; n14574
g12139 and n7445 n8960 ; n14575
g12140 and n14574 n14575 ; n14576
g12141 nor pi0051 n14576 ; n14577
g12142 and n14508_not n14577 ; n14578
g12143 and n6197 n14578_not ; n14579
g12144 nor n14507 n14579 ; n14580
g12145 and pi0142 n14580 ; n14581
g12146 and n2708 n14574 ; n14582
g12147 nor pi0072 n14582 ; n14583
g12148 and n6480 n14583_not ; n14584
g12149 and n6197 n14584_not ; n14585
g12150 nor n14528 n14585 ; n14586
g12151 nor pi0142 n14586 ; n14587
g12152 nor pi0144 n14581 ; n14588
g12153 and n14587_not n14588 ; n14589
g12154 nor pi0180 n14568 ; n14590
g12155 and n14589_not n14590 ; n14591
g12156 and n14505_not n14519 ; n14592
g12157 nor n14507 n14592 ; n14593
g12158 and n6197 n14504_not ; n14594
g12159 nor pi0142 n14594 ; n14595
g12160 nor pi0051 n14438 ; n14596
g12161 and n6197 n14596 ; n14597
g12162 nor n14536 n14597 ; n14598
g12163 and n2519 n14502_not ; n14599
g12164 nor n14598 n14599 ; n14600
g12165 and pi0142 n14600_not ; n14601
g12166 nor n14595 n14601 ; n14602
g12167 nor n14516 n14602 ; n14603
g12168 and n14593 n14603_not ; n14604
g12169 and pi0144 n14604_not ; n14605
g12170 and n2708 n14571 ; n14606
g12171 nor pi0072 n14606 ; n14607
g12172 and n6480 n14607_not ; n14608
g12173 and n6197 n14608_not ; n14609
g12174 nor n14528 n14609 ; n14610
g12175 nor pi0142 n14610 ; n14611
g12176 and n14536 n14606 ; n14612
g12177 nor n14510 n14612 ; n14613
g12178 and n14507_not n14613 ; n14614
g12179 and pi0142 n14614 ; n14615
g12180 nor pi0144 n14615 ; n14616
g12181 and n14611_not n14616 ; n14617
g12182 and pi0180 n14605_not ; n14618
g12183 and n14617_not n14618 ; n14619
g12184 nor pi0179 n14619 ; n14620
g12185 and n14591_not n14620 ; n14621
g12186 nor n14567 n14621 ; n14622
g12187 nor pi0299 n14622 ; n14623
g12188 and pi0146 n14614 ; n14624
g12189 nor pi0146 n14610 ; n14625
g12190 and n9572 n14624_not ; n14626
g12191 and n14625_not n14626 ; n14627
g12192 nor pi0146 n14586 ; n14628
g12193 and pi0146 n14580 ; n14629
g12194 and n9603 n14628_not ; n14630
g12195 and n14629_not n14630 ; n14631
g12196 nor pi0161 n14627 ; n14632
g12197 and n14631_not n14632 ; n14633
g12198 nor pi0146 n14594 ; n14634
g12199 and pi0146 n14600_not ; n14635
g12200 nor n14634 n14635 ; n14636
g12201 nor n14516 n14636 ; n14637
g12202 and n14593 n14637_not ; n14638
g12203 and n9572 n14638_not ; n14639
g12204 and n9603 n14444_not ; n14640
g12205 and n14506_not n14640 ; n14641
g12206 and pi0161 n14641_not ; n14642
g12207 and n14639_not n14642 ; n14643
g12208 nor pi0156 n14643 ; n14644
g12209 and n14633_not n14644 ; n14645
g12210 nor n14552 n14645 ; n14646
g12211 and n14623_not n14646 ; n14647
g12212 and n9159 n14647_not ; n14648
g12213 and n2519 n14490 ; n14649
g12214 nor n6640 n7607 ; n14650
g12215 and n14649 n14650_not ; n14651
g12216 and pi0232_not n14439 ; n14652
g12217 and n14651_not n14652 ; n14653
g12218 and n14439 n14649_not ; n14654
g12219 nor pi0051 n14654 ; n14655
g12220 nor pi0287 n14655 ; n14656
g12221 and pi0287_not n6197 ; n14657
g12222 nor n14597 n14657 ; n14658
g12223 nor n14656 n14658 ; n14659
g12224 nor n14460 n14659 ; n14660
g12225 and n9051 n14660_not ; n14661
g12226 and n14438 n14661 ; n14662
g12227 nor n14439 n14457 ; n14663
g12228 nor n6405 n14663 ; n14664
g12229 and pi0144 n14664_not ; n14665
g12230 and pi0051 n6197_not ; n14666
g12231 nor n14655 n14666 ; n14667
g12232 and n6405 n14459_not ; n14668
g12233 and n14667 n14668 ; n14669
g12234 and n14665 n14669_not ; n14670
g12235 and n14662_not n14670 ; n14671
g12236 nor n6197 n14654 ; n14672
g12237 nor n6222 n14672 ; n14673
g12238 nor pi0142 n14673 ; n14674
g12239 and n2515 n7450 ; n14675
g12240 nor pi0051 n14675 ; n14676
g12241 and n6197 n14676_not ; n14677
g12242 nor n14672 n14677 ; n14678
g12243 and pi0142 n14678_not ; n14679
g12244 and n6405 n14674_not ; n14680
g12245 and n14679_not n14680 ; n14681
g12246 nor n9051 n14681 ; n14682
g12247 and pi0051_not n14657 ; n14683
g12248 nor n14678 n14683 ; n14684
g12249 and pi0224 n14457_not ; n14685
g12250 and n14684 n14685 ; n14686
g12251 nor n14682 n14686 ; n14687
g12252 and n6405_not n14597 ; n14688
g12253 nor n14664 n14688 ; n14689
g12254 and n14665_not n14689 ; n14690
g12255 and n14687_not n14690 ; n14691
g12256 and pi0181 n14671_not ; n14692
g12257 and n14691_not n14692 ; n14693
g12258 and n14681_not n14690 ; n14694
g12259 nor pi0181 n14670 ; n14695
g12260 and n14694_not n14695 ; n14696
g12261 nor pi0299 n14696 ; n14697
g12262 and n14693_not n14697 ; n14698
g12263 nor n14444 n14654 ; n14699
g12264 and pi0161 n14699_not ; n14700
g12265 nor pi0146 n14673 ; n14701
g12266 and pi0146 n14678_not ; n14702
g12267 nor pi0161 n14701 ; n14703
g12268 and n14702_not n14703 ; n14704
g12269 nor n14700 n14704 ; n14705
g12270 and n6379 n14705_not ; n14706
g12271 nor n14439 n14448 ; n14707
g12272 nor n6379 n14707 ; n14708
g12273 and n9793 n14708_not ; n14709
g12274 and n14706_not n14709 ; n14710
g12275 nor n9036 n14706 ; n14711
g12276 and n14475 n14684 ; n14712
g12277 and n14649 n14657_not ; n14713
g12278 and n14439 n14713_not ; n14714
g12279 and n14445 n14714_not ; n14715
g12280 nor n14712 n14715 ; n14716
g12281 and pi0216 n14716_not ; n14717
g12282 nor n14711 n14717 ; n14718
g12283 and n9794 n14708_not ; n14719
g12284 and n14718_not n14719 ; n14720
g12285 and pi0232 n14710_not ; n14721
g12286 and n14698_not n14721 ; n14722
g12287 and n14720_not n14722 ; n14723
g12288 and pi0039 n14653_not ; n14724
g12289 and n14723_not n14724 ; n14725
g12290 nor pi0039 pi0232 ; n14726
g12291 and n14506_not n14726 ; n14727
g12292 nor n14725 n14727 ; n14728
g12293 and n14648_not n14728 ; n14729
g12294 nor pi0038 n14729 ; n14730
g12295 nor n14474 n14730 ; n14731
g12296 and n14468 n14469_not ; n14732
g12297 and n14731_not n14732 ; n14733
g12298 nor pi0184 pi0299 ; n14734
g12299 and pi0163_not pi0299 ; n14735
g12300 nor n14734 n14735 ; n14736
g12301 and n7473 n14736 ; n14737
g12302 and pi0087 n14737_not ; n14738
g12303 nor n14437 n14738 ; n14739
g12304 and n14466_not n14739 ; n14740
g12305 and n14733_not n14740 ; n14741
g12306 and n14455 n14465_not ; n14742
g12307 and pi0158_not n14463 ; n14743
g12308 and n14445 n14537_not ; n14744
g12309 and n6197 n14513_not ; n14745
g12310 and pi0146_not n14745 ; n14746
g12311 and n14438 n14485_not ; n14747
g12312 nor pi0051 n14747 ; n14748
g12313 and n2519 n14748_not ; n14749
g12314 nor n14598 n14749 ; n14750
g12315 and pi0146 n14750 ; n14751
g12316 nor pi0161 n14746 ; n14752
g12317 and n14751_not n14752 ; n14753
g12318 nor n14744 n14753 ; n14754
g12319 and n9572 n14754_not ; n14755
g12320 and pi0232 n14743_not ; n14756
g12321 and n14755_not n14756 ; n14757
g12322 and pi0156_not n2530 ; n14758
g12323 and n14757_not n14758 ; n14759
g12324 and pi0159_not n14463 ; n14760
g12325 and pi0181_not n14461 ; n14761
g12326 nor pi0144 n14460 ; n14762
g12327 and n14661_not n14762 ; n14763
g12328 and n9051 n14657 ; n14764
g12329 and pi0142 n2521_not ; n14765
g12330 nor pi0142 n14675 ; n14766
g12331 and n14764 n14765_not ; n14767
g12332 and n14766_not n14767 ; n14768
g12333 and n14458 n14768_not ; n14769
g12334 and pi0181 n14763_not ; n14770
g12335 and n14769_not n14770 ; n14771
g12336 nor pi0299 n14761 ; n14772
g12337 and n14771_not n14772 ; n14773
g12338 and n9036_not n14448 ; n14774
g12339 and n14475 n14659_not ; n14775
g12340 and n6197 n6380 ; n14776
g12341 and n14445 n14776_not ; n14777
g12342 and n9036 n14775_not ; n14778
g12343 and n14777_not n14778 ; n14779
g12344 and n9794 n14774_not ; n14780
g12345 and n14779_not n14780 ; n14781
g12346 and n10478 n14760_not ; n14782
g12347 and n14781_not n14782 ; n14783
g12348 and n14773_not n14783 ; n14784
g12349 and n6197 n14577_not ; n14785
g12350 and n14442_not n14785 ; n14786
g12351 and pi0161 n14786_not ; n14787
g12352 and n6197 n14514_not ; n14788
g12353 and pi0146_not n14788 ; n14789
g12354 and n14476 n14747 ; n14790
g12355 and n14501 n14790 ; n14791
g12356 and n14494 n14791_not ; n14792
g12357 and n2519 n14792_not ; n14793
g12358 nor n14598 n14793 ; n14794
g12359 and pi0146 n14794 ; n14795
g12360 nor pi0161 n14789 ; n14796
g12361 and n14795_not n14796 ; n14797
g12362 nor n14787 n14797 ; n14798
g12363 and n9572 n14798_not ; n14799
g12364 and n14445 n14612_not ; n14800
g12365 nor pi0161 n14636 ; n14801
g12366 nor n14800 n14801 ; n14802
g12367 and n9603 n14802_not ; n14803
g12368 and pi0232 n14803_not ; n14804
g12369 and n14799_not n14804 ; n14805
g12370 and pi0156 n14805_not ; n14806
g12371 and pi0142_not n14788 ; n14807
g12372 and pi0142 n14794 ; n14808
g12373 nor pi0144 n14807 ; n14809
g12374 and n14808_not n14809 ; n14810
g12375 and n14459_not n14785 ; n14811
g12376 and pi0144 n14811_not ; n14812
g12377 and pi0180 n14810_not ; n14813
g12378 and n14812_not n14813 ; n14814
g12379 and n14458 n14612_not ; n14815
g12380 nor pi0144 n14602 ; n14816
g12381 nor pi0180 n14816 ; n14817
g12382 and n14815_not n14817 ; n14818
g12383 and pi0179 n14818_not ; n14819
g12384 and n14814_not n14819 ; n14820
g12385 and pi0180_not n14461 ; n14821
g12386 and pi0142_not n14745 ; n14822
g12387 and pi0142 n14750 ; n14823
g12388 nor pi0144 n14822 ; n14824
g12389 and n14823_not n14824 ; n14825
g12390 and n14458 n14537_not ; n14826
g12391 and pi0180 n14825_not ; n14827
g12392 and n14826_not n14827 ; n14828
g12393 nor pi0179 n14821 ; n14829
g12394 and n14828_not n14829 ; n14830
g12395 nor n14820 n14830 ; n14831
g12396 nor pi0299 n14831 ; n14832
g12397 nor pi0039 n14806 ; n14833
g12398 and n14832_not n14833 ; n14834
g12399 nor pi0038 n14784 ; n14835
g12400 and n14834_not n14835 ; n14836
g12401 and n14471 n14759_not ; n14837
g12402 and n14836_not n14837 ; n14838
g12403 and n2535 n14469_not ; n14839
g12404 and n14838_not n14839 ; n14840
g12405 and n14437 n14738_not ; n14841
g12406 and n14742_not n14841 ; n14842
g12407 and n14840_not n14842 ; n14843
g12408 nor po1038 n14843 ; n14844
g12409 and n14741_not n14844 ; n14845
g12410 or n14454 n14845 ; po0279
g12411 and n7420 n7427 ; n14847
g12412 and n7429 n14407 ; n14848
g12413 and n14027 n14848_not ; n14849
g12414 and n7429 n14417 ; n14850
g12415 and n7425 n14850_not ; n14851
g12416 nor po1038 n14849 ; n14852
g12417 and n14851_not n14852 ; n14853
g12418 or n14847 n14853 ; po0280
g12419 and pi0110 n10075 ; n14855
g12420 and n10976_not n14855 ; n14856
g12421 and po1057 n14856 ; n14857
g12422 nor pi0039 n14857 ; n14858
g12423 and pi0110_not n9293 ; n14859
g12424 and n6244_not n6379 ; n14860
g12425 and n14859 n14860 ; n14861
g12426 and pi0039 n14861_not ; n14862
g12427 and po1038 n14858_not ; n14863
g12428 and n14862_not n14863 ; n14864
g12429 and pi0110 n13448 ; n14865
g12430 nor pi0039 n14865 ; n14866
g12431 and n6207_not n7607 ; n14867
g12432 and n14859 n14867 ; n14868
g12433 and pi0299 n14861 ; n14869
g12434 and pi0039 n14868_not ; n14870
g12435 and n14869_not n14870 ; n14871
g12436 nor n14866 n14871 ; n14872
g12437 and pi0038_not n2571 ; n14873
g12438 nor n14872 n14873 ; n14874
g12439 and pi0090 n10387_not ; n14875
g12440 nor pi0111 n6429 ; n14876
g12441 and pi0036_not n2809 ; n14877
g12442 and n14876_not n14877 ; n14878
g12443 and n2468 n14878_not ; n14879
g12444 nor n2793 n2798 ; n14880
g12445 and n14879_not n14880 ; n14881
g12446 nor pi0083 n14881 ; n14882
g12447 and n2795 n14882_not ; n14883
g12448 nor pi0071 n14883 ; n14884
g12449 and n6438 n14884_not ; n14885
g12450 nor pi0081 n14885 ; n14886
g12451 and n11443 n14886_not ; n14887
g12452 nor pi0090 n14887 ; n14888
g12453 and n2707 n14888_not ; n14889
g12454 and n9073 n14875_not ; n14890
g12455 and n14889 n14890 ; n14891
g12456 and pi0072 n2708 ; n14892
g12457 and n10387 n14892 ; n14893
g12458 nor n14891 n14893 ; n14894
g12459 and n6479 n14894_not ; n14895
g12460 nor pi0110 n14895 ; n14896
g12461 and n13448 n14896_not ; n14897
g12462 and n2897 n14889 ; n14898
g12463 nor pi0072 n14898 ; n14899
g12464 and n6480 n13448_not ; n14900
g12465 and n14899_not n14900 ; n14901
g12466 nor pi0039 n14901 ; n14902
g12467 and n14897_not n14902 ; n14903
g12468 nor n14871 n14903 ; n14904
g12469 and n14873 n14904_not ; n14905
g12470 nor po1038 n14874 ; n14906
g12471 and n14905_not n14906 ; n14907
g12472 nor n14864 n14907 ; po0281
g12473 and pi0125_not n14432 ; n14909
g12474 and pi0125 pi0133 ; n14910
g12475 nor n14433 n14910 ; n14911
g12476 nor n14909 n14911 ; n14912
g12477 and n14439 n14912_not ; n14913
g12478 and pi0172 n14443 ; n14914
g12479 and pi0152_not n14597 ; n14915
g12480 nor n14914 n14915 ; n14916
g12481 and pi0232 n14916_not ; n14917
g12482 nor n14913 n14917 ; n14918
g12483 nor pi0087 n14918 ; n14919
g12484 and pi0087 n7473 ; n14920
g12485 and pi0162 n14920 ; n14921
g12486 and po1038 n14921_not ; n14922
g12487 and n14919_not n14922 ; n14923
g12488 and pi0193 n14443 ; n14924
g12489 and pi0174_not n14597 ; n14925
g12490 nor pi0299 n14924 ; n14926
g12491 and n14925_not n14926 ; n14927
g12492 and pi0299 n14916 ; n14928
g12493 and pi0232 n14927_not ; n14929
g12494 and n14928_not n14929 ; n14930
g12495 and n14455 n14930_not ; n14931
g12496 and pi0140 pi0299_not ; n14932
g12497 and pi0162 pi0299 ; n14933
g12498 nor n14932 n14933 ; n14934
g12499 and n7473 n14934_not ; n14935
g12500 and pi0087 n14935_not ; n14936
g12501 and pi0100 n14930 ; n14937
g12502 nor pi0232 n14508 ; n14938
g12503 nor pi0039 n14938 ; n14939
g12504 nor pi0299 n7551 ; n14940
g12505 and pi0299 n7570_not ; n14941
g12506 nor n14940 n14941 ; n14942
g12507 and n2521 n14942 ; n14943
g12508 nor pi0232 n14943 ; n14944
g12509 and pi0039 n14944_not ; n14945
g12510 and n7570_not n14916 ; n14946
g12511 and n2521 n6197_not ; n14947
g12512 and n6197 n14654_not ; n14948
g12513 nor n14947 n14948 ; n14949
g12514 nor pi0152 n14949 ; n14950
g12515 nor n14677 n14947 ; n14951
g12516 and pi0152 n14951_not ; n14952
g12517 nor n14950 n14952 ; n14953
g12518 and pi0051 pi0172_not ; n14954
g12519 nor n14953 n14954 ; n14955
g12520 nor pi0216 n14955 ; n14956
g12521 and n6379 n14956 ; n14957
g12522 nor n14946 n14957 ; n14958
g12523 and n9603 n14958_not ; n14959
g12524 nor n6379 n14916 ; n14960
g12525 and n14649 n14657 ; n14961
g12526 nor n14446 n14961 ; n14962
g12527 and pi0152_not n14962 ; n14963
g12528 and n14657 n14675 ; n14964
g12529 nor n14443 n14964 ; n14965
g12530 and pi0152 n14965 ; n14966
g12531 and pi0172 n14963_not ; n14967
g12532 and n14966_not n14967 ; n14968
g12533 nor pi0152 n14659 ; n14969
g12534 and pi0152 n14776_not ; n14970
g12535 nor pi0172 n14969 ; n14971
g12536 and n14970_not n14971 ; n14972
g12537 and pi0216 n14968_not ; n14973
g12538 and n14972_not n14973 ; n14974
g12539 and n6379 n14974_not ; n14975
g12540 and n14956_not n14975 ; n14976
g12541 and n9572 n14960_not ; n14977
g12542 and n14976_not n14977 ; n14978
g12543 nor n7551 n14446 ; n14979
g12544 and n6197 n14655 ; n14980
g12545 nor n14947 n14980 ; n14981
g12546 nor n14979 n14981 ; n14982
g12547 and pi0174_not n14982 ; n14983
g12548 and n2521 n7551 ; n14984
g12549 and pi0174 n14984 ; n14985
g12550 nor n14924 n14985 ; n14986
g12551 and n14983_not n14986 ; n14987
g12552 nor pi0180 n14987 ; n14988
g12553 and n7551 n14949 ; n14989
g12554 and pi0224 n14961_not ; n14990
g12555 and n6405 n14990_not ; n14991
g12556 nor n14446 n14991 ; n14992
g12557 nor n14989 n14992 ; n14993
g12558 and pi0174_not n14993 ; n14994
g12559 and pi0224 n14965 ; n14995
g12560 and n6405 n14995_not ; n14996
g12561 and n7551 n14951 ; n14997
g12562 and n14996 n14997_not ; n14998
g12563 nor n14443 n14998 ; n14999
g12564 and pi0174 n14999_not ; n15000
g12565 and pi0193 n14994_not ; n15001
g12566 and n15000_not n15001 ; n15002
g12567 nor n7551 n14764 ; n15003
g12568 and n2521 n15003_not ; n15004
g12569 and pi0174 n15004 ; n15005
g12570 and pi0224 n14659_not ; n15006
g12571 and pi0224_not n14981 ; n15007
g12572 and n6405 n15006_not ; n15008
g12573 and n15007_not n15008 ; n15009
g12574 nor n14688 n15009 ; n15010
g12575 nor pi0174 n15010 ; n15011
g12576 nor pi0193 n15005 ; n15012
g12577 and n15011_not n15012 ; n15013
g12578 and pi0180 n15013_not ; n15014
g12579 and n15002_not n15014 ; n15015
g12580 nor pi0299 n14988 ; n15016
g12581 and n15015_not n15016 ; n15017
g12582 nor n14959 n14978 ; n15018
g12583 and n15017_not n15018 ; n15019
g12584 and pi0232 n15019_not ; n15020
g12585 and n14945 n15020_not ; n15021
g12586 nor pi0038 n14939 ; n15022
g12587 and n15021_not n15022 ; n15023
g12588 and pi0038 n14930_not ; n15024
g12589 nor pi0100 n15024 ; n15025
g12590 and pi0152_not n14521 ; n15026
g12591 and pi0152_not n6197 ; n15027
g12592 and n14508 n15027_not ; n15028
g12593 nor pi0197 n15026 ; n15029
g12594 and n15028_not n15029 ; n15030
g12595 and n6197_not n14508 ; n15031
g12596 nor n14519 n15031 ; n15032
g12597 nor n14543 n15032 ; n15033
g12598 and pi0152_not pi0197 ; n15034
g12599 and n15033_not n15034 ; n15035
g12600 nor n15030 n15035 ; n15036
g12601 nor n14914 n15036 ; n15037
g12602 nor n6197 n14508 ; n15038
g12603 nor n14533 n15038 ; n15039
g12604 and pi0172_not n15039 ; n15040
g12605 nor n14443 n14537 ; n15041
g12606 and n14508_not n15041 ; n15042
g12607 and pi0172 n15042_not ; n15043
g12608 and pi0152 pi0197 ; n15044
g12609 and n15043_not n15044 ; n15045
g12610 and n15040_not n15045 ; n15046
g12611 nor n15037 n15046 ; n15047
g12612 and n9766 n15047_not ; n15048
g12613 and n14505 n14542 ; n15049
g12614 nor n15038 n15049 ; n15050
g12615 and pi0152_not n15050 ; n15051
g12616 and n14509 n14612_not ; n15052
g12617 and pi0152 n15052_not ; n15053
g12618 and pi0172 n15051_not ; n15054
g12619 and n15053_not n15054 ; n15055
g12620 nor n14609 n15038 ; n15056
g12621 and pi0152 n15056 ; n15057
g12622 nor n14592 n15031 ; n15058
g12623 nor pi0152 n15058 ; n15059
g12624 nor pi0172 n15059 ; n15060
g12625 and n15057_not n15060 ; n15061
g12626 nor pi0197 n15055 ; n15062
g12627 and n15061_not n15062 ; n15063
g12628 nor n14585 n15038 ; n15064
g12629 and pi0172_not n15064 ; n15065
g12630 nor n14578 n15038 ; n15066
g12631 and pi0172 n15066 ; n15067
g12632 and pi0152 n15067_not ; n15068
g12633 and n15065_not n15068 ; n15069
g12634 and n6197 n14506 ; n15070
g12635 nor n15032 n15070 ; n15071
g12636 nor pi0152 n14914 ; n15072
g12637 and n15071_not n15072 ; n15073
g12638 and pi0197 n15073_not ; n15074
g12639 and n15069_not n15074 ; n15075
g12640 and n9760 n15063_not ; n15076
g12641 and n15075_not n15076 ; n15077
g12642 nor n15048 n15077 ; n15078
g12643 and pi0299 n15078_not ; n15079
g12644 and pi0145_not n14508 ; n15080
g12645 and pi0145 n15039 ; n15081
g12646 and pi0174 n15080_not ; n15082
g12647 and n15081_not n15082 ; n15083
g12648 nor n14521 n15031 ; n15084
g12649 nor pi0145 n15084 ; n15085
g12650 and pi0145 n15033 ; n15086
g12651 nor pi0174 n15085 ; n15087
g12652 and n15086_not n15087 ; n15088
g12653 nor n15083 n15088 ; n15089
g12654 nor pi0193 n15089 ; n15090
g12655 and pi0145_not n14537 ; n15091
g12656 nor n15041 n15091 ; n15092
g12657 nor n14508 n15092 ; n15093
g12658 and pi0174 n15093_not ; n15094
g12659 nor n14443 n14486 ; n15095
g12660 and pi0145 n15095_not ; n15096
g12661 and n14542 n15096_not ; n15097
g12662 nor pi0174 n15097 ; n15098
g12663 and n15038_not n15098 ; n15099
g12664 and pi0193 n15099_not ; n15100
g12665 and n15094_not n15100 ; n15101
g12666 nor n15090 n15101 ; n15102
g12667 and n9772 n15102_not ; n15103
g12668 and pi0193 n15050 ; n15104
g12669 nor pi0193 n15058 ; n15105
g12670 nor pi0145 n15104 ; n15106
g12671 and n15105_not n15106 ; n15107
g12672 and pi0145 n14924_not ; n15108
g12673 and n15071_not n15108 ; n15109
g12674 nor pi0174 n15109 ; n15110
g12675 and n15107_not n15110 ; n15111
g12676 and pi0145 n15066 ; n15112
g12677 nor pi0145 n15052 ; n15113
g12678 and pi0193 n15113_not ; n15114
g12679 and n15112_not n15114 ; n15115
g12680 and pi0145_not n15056 ; n15116
g12681 and pi0145 n15064 ; n15117
g12682 nor pi0193 n15116 ; n15118
g12683 and n15117_not n15118 ; n15119
g12684 and pi0174 n15115_not ; n15120
g12685 and n15119_not n15120 ; n15121
g12686 and n9776 n15111_not ; n15122
g12687 and n15121_not n15122 ; n15123
g12688 nor n15103 n15123 ; n15124
g12689 nor pi0038 n15124 ; n15125
g12690 nor n15079 n15125 ; n15126
g12691 and n9159 n15126_not ; n15127
g12692 and n15023_not n15025 ; n15128
g12693 and n15127_not n15128 ; n15129
g12694 and n2535 n14937_not ; n15130
g12695 and n15129_not n15130 ; n15131
g12696 and n14912 n14936_not ; n15132
g12697 and n14931_not n15132 ; n15133
g12698 and n15131_not n15133 ; n15134
g12699 and n14456 n14930_not ; n15135
g12700 nor n14473 n15025 ; n15136
g12701 nor n14515 n14612 ; n15137
g12702 and pi0145 n15137 ; n15138
g12703 and n14536 n14582 ; n15139
g12704 nor n14515 n15139 ; n15140
g12705 and pi0145_not n15140 ; n15141
g12706 nor pi0174 n15138 ; n15142
g12707 and n15141_not n15142 ; n15143
g12708 nor n14515 n14794 ; n15144
g12709 nor pi0145 n14513 ; n15145
g12710 nor n6197 n14513 ; n15146
g12711 nor n14446 n15146 ; n15147
g12712 and n14503_not n15147 ; n15148
g12713 and n15145_not n15148 ; n15149
g12714 and n2519 n15149 ; n15150
g12715 and pi0174 n15144_not ; n15151
g12716 and n15150_not n15151 ; n15152
g12717 and pi0193 n15152_not ; n15153
g12718 and n15143_not n15153 ; n15154
g12719 and pi0174 n15149_not ; n15155
g12720 and pi0051_not n15138 ; n15156
g12721 nor pi0145 n14515 ; n15157
g12722 and n14785_not n15157 ; n15158
g12723 nor pi0174 n15156 ; n15159
g12724 and n15158_not n15159 ; n15160
g12725 nor pi0193 n15155 ; n15161
g12726 and n15160_not n15161 ; n15162
g12727 and n9772 n15154_not ; n15163
g12728 and n15162_not n15163 ; n15164
g12729 and pi0145 n14597_not ; n15165
g12730 nor pi0174 n15091 ; n15166
g12731 and pi0145_not pi0174 ; n15167
g12732 and n14750_not n15167 ; n15168
g12733 nor n15165 n15168 ; n15169
g12734 and n15166_not n15169 ; n15170
g12735 and pi0193 n14515_not ; n15171
g12736 and n15170_not n15171 ; n15172
g12737 nor n14443 n14515 ; n15173
g12738 and pi0145 n14438 ; n15174
g12739 nor n15166 n15174 ; n15175
g12740 and n15173 n15175_not ; n15176
g12741 nor n14515 n14745 ; n15177
g12742 and pi0174 n15177 ; n15178
g12743 nor n15176 n15178 ; n15179
g12744 nor pi0193 n15179 ; n15180
g12745 and n9776 n15172_not ; n15181
g12746 and n15180_not n15181 ; n15182
g12747 nor n15164 n15182 ; n15183
g12748 nor pi0038 n15183 ; n15184
g12749 and pi0172_not n14443 ; n15185
g12750 and pi0172_not n15148 ; n15186
g12751 nor n14515 n14600 ; n15187
g12752 and pi0172 n15187 ; n15188
g12753 and pi0152 n15186_not ; n15189
g12754 and n15188_not n15189 ; n15190
g12755 nor pi0152 n15137 ; n15191
g12756 and pi0197 n15185_not ; n15192
g12757 and n15190_not n15192 ; n15193
g12758 and n15191_not n15193 ; n15194
g12759 nor pi0152 n15140 ; n15195
g12760 and pi0152 n15144_not ; n15196
g12761 and pi0172 n15196_not ; n15197
g12762 and n15195_not n15197 ; n15198
g12763 and pi0152_not n14785 ; n15199
g12764 nor n14514 n15027 ; n15200
g12765 nor pi0172 n15200 ; n15201
g12766 and n15199_not n15201 ; n15202
g12767 nor n15198 n15202 ; n15203
g12768 nor pi0197 n15203 ; n15204
g12769 and pi0299 n9766 ; n15205
g12770 and n15194_not n15205 ; n15206
g12771 and n15204_not n15206 ; n15207
g12772 and pi0152 n14597 ; n15208
g12773 nor n14515 n15208 ; n15209
g12774 and pi0172 n15209_not ; n15210
g12775 nor pi0172 n14915 ; n15211
g12776 and n14516_not n15211 ; n15212
g12777 and pi0197 n15210_not ; n15213
g12778 and n15212_not n15213 ; n15214
g12779 and pi0152 n15177 ; n15215
g12780 nor n14515 n14537 ; n15216
g12781 and pi0152_not n15216 ; n15217
g12782 and n14443_not n15217 ; n15218
g12783 nor pi0172 n15215 ; n15219
g12784 and n15218_not n15219 ; n15220
g12785 nor n14515 n14750 ; n15221
g12786 and pi0152 n15221 ; n15222
g12787 and pi0172 n15222_not ; n15223
g12788 and n15217_not n15223 ; n15224
g12789 nor pi0197 n15224 ; n15225
g12790 and n15220_not n15225 ; n15226
g12791 and pi0299 n9760 ; n15227
g12792 and n15214_not n15227 ; n15228
g12793 and n15226_not n15228 ; n15229
g12794 nor n15207 n15229 ; n15230
g12795 and n15184_not n15230 ; n15231
g12796 and n9159 n15231_not ; n15232
g12797 and n14439_not n14916 ; n15233
g12798 nor n9036 n15233 ; n15234
g12799 nor n14654 n15027 ; n15235
g12800 and pi0152_not n14677 ; n15236
g12801 nor n15235 n15236 ; n15237
g12802 nor pi0172 n15237 ; n15238
g12803 and pi0152_not n14673 ; n15239
g12804 and pi0152 n14667 ; n15240
g12805 and pi0172 n15240_not ; n15241
g12806 and n15239_not n15241 ; n15242
g12807 and n9036 n15238_not ; n15243
g12808 and n15242_not n15243 ; n15244
g12809 and n9603 n15244_not ; n15245
g12810 and pi0152 n14914_not ; n15246
g12811 and n14714_not n15246 ; n15247
g12812 and n14684 n15072 ; n15248
g12813 and n9036 n15247_not ; n15249
g12814 and n15248_not n15249 ; n15250
g12815 and n9572 n15250_not ; n15251
g12816 nor n15245 n15251 ; n15252
g12817 nor n15234 n15252 ; n15253
g12818 and pi0180 n14714 ; n15254
g12819 and n9051 n14649 ; n15255
g12820 and n14439 n15255_not ; n15256
g12821 and pi0174 n15256_not ; n15257
g12822 and n15254_not n15257 ; n15258
g12823 and n9051 n14678 ; n15259
g12824 nor n6197 n14438 ; n15260
g12825 nor n9051 n15260 ; n15261
g12826 and pi0051_not n15261 ; n15262
g12827 nor n15259 n15262 ; n15263
g12828 and pi0180 n14683 ; n15264
g12829 nor pi0174 n15264 ; n15265
g12830 and n15263 n15265 ; n15266
g12831 nor pi0193 n15258 ; n15267
g12832 and n15266_not n15267 ; n15268
g12833 and n14666_not n15261 ; n15269
g12834 and n9051 n14673 ; n15270
g12835 nor n15269 n15270 ; n15271
g12836 nor pi0174 n15271 ; n15272
g12837 nor n14443 n15256 ; n15273
g12838 and pi0174 n15273_not ; n15274
g12839 nor pi0180 n15274 ; n15275
g12840 and n15272_not n15275 ; n15276
g12841 and n9051 n14672_not ; n15277
g12842 and n10603_not n15277 ; n15278
g12843 nor n15269 n15278 ; n15279
g12844 nor pi0174 n15279 ; n15280
g12845 nor pi0051 n14714 ; n15281
g12846 and n6197 n15281_not ; n15282
g12847 nor n15256 n15282 ; n15283
g12848 and pi0174 n15283_not ; n15284
g12849 and pi0180 n15284_not ; n15285
g12850 and n15280_not n15285 ; n15286
g12851 and pi0193 n15286_not ; n15287
g12852 and n15276_not n15287 ; n15288
g12853 nor pi0299 n15268 ; n15289
g12854 and n15288_not n15289 ; n15290
g12855 nor n15253 n15290 ; n15291
g12856 and pi0232 n15291_not ; n15292
g12857 nor pi0299 n15256 ; n15293
g12858 and n9036 n14649 ; n15294
g12859 and n14439 n15294_not ; n15295
g12860 and pi0299 n15295_not ; n15296
g12861 nor n15293 n15296 ; n15297
g12862 nor pi0232 n15297 ; n15298
g12863 and pi0039 n15298_not ; n15299
g12864 and n15292_not n15299 ; n15300
g12865 nor pi0232 n14514 ; n15301
g12866 nor pi0039 n15301 ; n15302
g12867 nor pi0038 n15302 ; n15303
g12868 and n15300_not n15303 ; n15304
g12869 nor n15136 n15304 ; n15305
g12870 and n15232_not n15305 ; n15306
g12871 and n14468 n14937_not ; n15307
g12872 and n15306_not n15307 ; n15308
g12873 nor n14912 n14936 ; n15309
g12874 and n15135_not n15309 ; n15310
g12875 and n15308_not n15310 ; n15311
g12876 nor po1038 n15311 ; n15312
g12877 and n15134_not n15312 ; n15313
g12878 or n14923 n15313 ; po0282
g12879 and pi0175 n14443 ; n15315
g12880 and pi0189_not n14597 ; n15316
g12881 nor pi0299 n15315 ; n15317
g12882 and n15316_not n15317 ; n15318
g12883 nor pi0051 n14597 ; n15319
g12884 nor n10299 n14438 ; n15320
g12885 nor pi0051 n15320 ; n15321
g12886 and pi0153 n14443 ; n15322
g12887 nor n15321 n15322 ; n15323
g12888 nor n15319 n15323 ; n15324
g12889 and pi0299 n15324_not ; n15325
g12890 and pi0232 n15318_not ; n15326
g12891 and n15325_not n15326 ; n15327
g12892 and n2608_not n15327 ; n15328
g12893 and pi0126_not n14435 ; n15329
g12894 and pi0126 n14435_not ; n15330
g12895 nor n15329 n15330 ; n15331
g12896 nor n14431 n15331 ; n15332
g12897 and n2608_not n14439 ; n15333
g12898 and n15332_not n15333 ; n15334
g12899 and pi0182 n14714 ; n15335
g12900 and pi0189 n15256_not ; n15336
g12901 and n15335_not n15336 ; n15337
g12902 and pi0182 n14683 ; n15338
g12903 nor pi0189 n15338 ; n15339
g12904 and n15263 n15339 ; n15340
g12905 nor n15337 n15340 ; n15341
g12906 and n11765 n15341_not ; n15342
g12907 nor pi0189 n15271 ; n15343
g12908 and pi0189 n15273_not ; n15344
g12909 nor pi0182 n15344 ; n15345
g12910 and n15343_not n15345 ; n15346
g12911 nor pi0189 n15279 ; n15347
g12912 and pi0189 n15283_not ; n15348
g12913 and pi0182 n15348_not ; n15349
g12914 and n15347_not n15349 ; n15350
g12915 nor n15346 n15350 ; n15351
g12916 and n11833 n15351_not ; n15352
g12917 nor n9036 n15323 ; n15353
g12918 and pi0166_not n14684 ; n15354
g12919 and pi0166 n14714_not ; n15355
g12920 nor n15354 n15355 ; n15356
g12921 and pi0160 n15322_not ; n15357
g12922 and n15356_not n15357 ; n15358
g12923 nor n10299 n14654 ; n15359
g12924 and pi0166_not n14677 ; n15360
g12925 nor n15359 n15360 ; n15361
g12926 nor pi0153 n15361 ; n15362
g12927 and pi0166_not n14673 ; n15363
g12928 and pi0166 n14667 ; n15364
g12929 and pi0153 n15364_not ; n15365
g12930 and n15363_not n15365 ; n15366
g12931 nor n15362 n15366 ; n15367
g12932 nor pi0160 n15367 ; n15368
g12933 and n9036 n15358_not ; n15369
g12934 and n15368_not n15369 ; n15370
g12935 and pi0299 n15353_not ; n15371
g12936 and n15370_not n15371 ; n15372
g12937 nor n15342 n15352 ; n15373
g12938 and n15372_not n15373 ; n15374
g12939 and pi0232 n15374_not ; n15375
g12940 and n15299 n15375_not ; n15376
g12941 and pi0189_not n15173 ; n15377
g12942 and pi0178 n15377_not ; n15378
g12943 and pi0189 n14516 ; n15379
g12944 and n15378 n15379_not ; n15380
g12945 and pi0189 n15148 ; n15381
g12946 and n14612_not n15377 ; n15382
g12947 nor pi0178 n15381 ; n15383
g12948 and n15382_not n15383 ; n15384
g12949 and pi0181 n15380_not ; n15385
g12950 and n15384_not n15385 ; n15386
g12951 and pi0189 n15177 ; n15387
g12952 and pi0189_not n15216 ; n15388
g12953 and pi0178 n15388_not ; n15389
g12954 nor n15378 n15389 ; n15390
g12955 nor n15387 n15390 ; n15391
g12956 nor n10295 n14514 ; n15392
g12957 and pi0189_not n14785 ; n15393
g12958 nor n15392 n15393 ; n15394
g12959 nor pi0178 n15394 ; n15395
g12960 nor pi0181 n15391 ; n15396
g12961 and n15395_not n15396 ; n15397
g12962 and n11765 n15386_not ; n15398
g12963 and n15397_not n15398 ; n15399
g12964 nor pi0189 n14612 ; n15400
g12965 and pi0189 n14600_not ; n15401
g12966 nor pi0178 n15401 ; n15402
g12967 and n15400_not n15402 ; n15403
g12968 and pi0178 n11826 ; n15404
g12969 and n14596 n15404 ; n15405
g12970 and pi0181 n15405_not ; n15406
g12971 and n14515_not n15406 ; n15407
g12972 and n15403_not n15407 ; n15408
g12973 and pi0189 n15221 ; n15409
g12974 and n15389 n15409_not ; n15410
g12975 and pi0189_not n15140 ; n15411
g12976 and pi0189 n15144 ; n15412
g12977 nor pi0178 n15412 ; n15413
g12978 and n15411_not n15413 ; n15414
g12979 nor pi0181 n15410 ; n15415
g12980 and n15414_not n15415 ; n15416
g12981 and n11833 n15408_not ; n15417
g12982 and n15416_not n15417 ; n15418
g12983 and pi0166 n14597 ; n15419
g12984 nor n14515 n15419 ; n15420
g12985 and pi0153 n15420_not ; n15421
g12986 nor pi0153 n15324 ; n15422
g12987 and n14516_not n15422 ; n15423
g12988 and pi0157 n15421_not ; n15424
g12989 and n15423_not n15424 ; n15425
g12990 and pi0153 pi0166 ; n15426
g12991 and n15187_not n15426 ; n15427
g12992 nor pi0166 n15137 ; n15428
g12993 and pi0166 n15148_not ; n15429
g12994 and pi0051 n10299 ; n15430
g12995 nor n15429 n15430 ; n15431
g12996 nor pi0153 n15431 ; n15432
g12997 nor pi0157 n15427 ; n15433
g12998 and n15432_not n15433 ; n15434
g12999 and n15428_not n15434 ; n15435
g13000 and n9794 n15425_not ; n15436
g13001 and n15435_not n15436 ; n15437
g13002 nor pi0166 n15216 ; n15438
g13003 and pi0166 n15177_not ; n15439
g13004 nor n15430 n15439 ; n15440
g13005 nor pi0153 n15440 ; n15441
g13006 and n15221_not n15426 ; n15442
g13007 and pi0157 n15442_not ; n15443
g13008 and n15438_not n15443 ; n15444
g13009 and n15441_not n15444 ; n15445
g13010 nor pi0166 n15140 ; n15446
g13011 and pi0166 n15144_not ; n15447
g13012 and pi0153 n15447_not ; n15448
g13013 and n15446_not n15448 ; n15449
g13014 and pi0166_not n14785 ; n15450
g13015 nor n10299 n14514 ; n15451
g13016 nor pi0153 n15451 ; n15452
g13017 and n15450_not n15452 ; n15453
g13018 nor n15449 n15453 ; n15454
g13019 nor pi0157 n15454 ; n15455
g13020 and n9793 n15445_not ; n15456
g13021 and n15455_not n15456 ; n15457
g13022 nor n15418 n15437 ; n15458
g13023 and n15399_not n15458 ; n15459
g13024 and n15457_not n15459 ; n15460
g13025 and pi0232 n15460_not ; n15461
g13026 and n15302 n15461_not ; n15462
g13027 nor n15332 n15376 ; n15463
g13028 and n15462_not n15463 ; n15464
g13029 and pi0189_not n14982 ; n15465
g13030 and pi0189 n14984 ; n15466
g13031 nor pi0182 n15466 ; n15467
g13032 and n15465_not n15467 ; n15468
g13033 and n14443_not n15468 ; n15469
g13034 and pi0189_not n14993 ; n15470
g13035 and pi0189 n14999_not ; n15471
g13036 and pi0182 n15470_not ; n15472
g13037 and n15471_not n15472 ; n15473
g13038 nor n15469 n15473 ; n15474
g13039 and n11833 n15474_not ; n15475
g13040 nor pi0189 n15010 ; n15476
g13041 and pi0189 n15004 ; n15477
g13042 and pi0182 n15477_not ; n15478
g13043 and n15476_not n15478 ; n15479
g13044 nor n15468 n15479 ; n15480
g13045 and n11765 n15480_not ; n15481
g13046 and pi0160_not pi0216 ; n15482
g13047 and n6379 n15482_not ; n15483
g13048 and n15324 n15483_not ; n15484
g13049 and pi0166_not n14659 ; n15485
g13050 and pi0166 n14776 ; n15486
g13051 nor pi0153 n15485 ; n15487
g13052 and n15486_not n15487 ; n15488
g13053 and pi0166 n14965_not ; n15489
g13054 nor pi0166 n14962 ; n15490
g13055 and pi0153 n15490_not ; n15491
g13056 and n15489_not n15491 ; n15492
g13057 and pi0160 n15488_not ; n15493
g13058 and n15492_not n15493 ; n15494
g13059 and pi0216 n15494_not ; n15495
g13060 nor pi0166 n14949 ; n15496
g13061 and pi0166 n14951_not ; n15497
g13062 nor n15496 n15497 ; n15498
g13063 and pi0051 pi0153_not ; n15499
g13064 nor n15498 n15499 ; n15500
g13065 nor pi0216 n15500 ; n15501
g13066 and n6379 n15495_not ; n15502
g13067 and n15501_not n15502 ; n15503
g13068 and pi0299 n15484_not ; n15504
g13069 and n15503_not n15504 ; n15505
g13070 nor n15475 n15481 ; n15506
g13071 and n15505_not n15506 ; n15507
g13072 and pi0232 n15507_not ; n15508
g13073 and n14945 n15508_not ; n15509
g13074 and pi0153_not n15064 ; n15510
g13075 and pi0153 n15066 ; n15511
g13076 and pi0157 n15511_not ; n15512
g13077 and n15510_not n15512 ; n15513
g13078 and pi0153_not n15039 ; n15514
g13079 and pi0153 n15042_not ; n15515
g13080 nor pi0157 n15515 ; n15516
g13081 and n15514_not n15516 ; n15517
g13082 nor n15513 n15517 ; n15518
g13083 and pi0166 n15518_not ; n15519
g13084 and pi0157 n15071 ; n15520
g13085 and pi0157_not n15033 ; n15521
g13086 nor pi0166 n15322 ; n15522
g13087 and n15520_not n15522 ; n15523
g13088 and n15521_not n15523 ; n15524
g13089 nor n15519 n15524 ; n15525
g13090 and n9794 n15525_not ; n15526
g13091 and pi0166_not n15050 ; n15527
g13092 and pi0166 n15052_not ; n15528
g13093 and pi0153 n15527_not ; n15529
g13094 and n15528_not n15529 ; n15530
g13095 and pi0166 n15056 ; n15531
g13096 nor pi0166 n15058 ; n15532
g13097 nor pi0153 n15532 ; n15533
g13098 and n15531_not n15533 ; n15534
g13099 nor n15530 n15534 ; n15535
g13100 and pi0157 n15535_not ; n15536
g13101 and pi0166 n14508 ; n15537
g13102 nor pi0166 n15084 ; n15538
g13103 nor pi0157 n15322 ; n15539
g13104 and n15537_not n15539 ; n15540
g13105 and n15538_not n15540 ; n15541
g13106 nor n15536 n15541 ; n15542
g13107 and n9793 n15542_not ; n15543
g13108 nor pi0189 n15084 ; n15544
g13109 and pi0189 n14508 ; n15545
g13110 nor pi0178 n15545 ; n15546
g13111 and n14443_not n15546 ; n15547
g13112 and n15544_not n15547 ; n15548
g13113 nor pi0181 n15548 ; n15549
g13114 and pi0189 n15052_not ; n15550
g13115 and pi0189_not n15050 ; n15551
g13116 and pi0178 n15551_not ; n15552
g13117 and n15550_not n15552 ; n15553
g13118 and n15549 n15553_not ; n15554
g13119 and pi0189 n15042 ; n15555
g13120 nor pi0189 n15033 ; n15556
g13121 and n14443_not n15556 ; n15557
g13122 nor n15555 n15557 ; n15558
g13123 nor pi0178 n15558 ; n15559
g13124 and pi0189_not n15071 ; n15560
g13125 and n15066 n15377_not ; n15561
g13126 and pi0178 n15560_not ; n15562
g13127 and n15561_not n15562 ; n15563
g13128 and pi0181 n15559_not ; n15564
g13129 and n15563_not n15564 ; n15565
g13130 and n11833 n15554_not ; n15566
g13131 and n15565_not n15566 ; n15567
g13132 and n15084 n15546 ; n15568
g13133 nor pi0189 n15058 ; n15569
g13134 and pi0189 n15056 ; n15570
g13135 and pi0178 n15569_not ; n15571
g13136 and n15570_not n15571 ; n15572
g13137 and n15549 n15568_not ; n15573
g13138 and n15572_not n15573 ; n15574
g13139 and pi0189 n15064 ; n15575
g13140 nor n15560 n15575 ; n15576
g13141 and pi0178 n15576_not ; n15577
g13142 and pi0189 n15039_not ; n15578
g13143 nor pi0178 n15556 ; n15579
g13144 and n15578_not n15579 ; n15580
g13145 nor n15577 n15580 ; n15581
g13146 and pi0181 n15581_not ; n15582
g13147 and n11765 n15574_not ; n15583
g13148 and n15582_not n15583 ; n15584
g13149 nor n15543 n15567 ; n15585
g13150 and n15526_not n15585 ; n15586
g13151 and n15584_not n15586 ; n15587
g13152 and pi0232 n15587_not ; n15588
g13153 and n14939 n15588_not ; n15589
g13154 and n15332 n15509_not ; n15590
g13155 and n15589_not n15590 ; n15591
g13156 and n2608 n15464_not ; n15592
g13157 and n15591_not n15592 ; n15593
g13158 and n2535 n15334_not ; n15594
g13159 and n15328_not n15594 ; n15595
g13160 and n15593_not n15595 ; n15596
g13161 and n14455 n15327_not ; n15597
g13162 and pi0150_not pi0299 ; n15598
g13163 nor pi0185 pi0299 ; n15599
g13164 nor n15598 n15599 ; n15600
g13165 and n7473 n15600 ; n15601
g13166 and pi0087 n15601_not ; n15602
g13167 nor n15597 n15602 ; n15603
g13168 and n14440 n15332_not ; n15604
g13169 nor n15603 n15604 ; n15605
g13170 nor po1038 n15605 ; n15606
g13171 and n15596_not n15606 ; n15607
g13172 and pi0232 n15319_not ; n15608
g13173 and n15332 n15608_not ; n15609
g13174 nor pi0232 n14439 ; n15610
g13175 nor n15323 n15610 ; n15611
g13176 and n15609_not n15611 ; n15612
g13177 nor pi0087 n15612 ; n15613
g13178 and pi0087 n13685_not ; n15614
g13179 and po1038 n15614_not ; n15615
g13180 and n15613_not n15615 ; n15616
g13181 nor n15607 n15616 ; po0283
g13182 and n2537 n8887 ; n15618
g13183 and n2529 n15618 ; n15619
g13184 nor n3328 n15619 ; n15620
g13185 nor n2529 n15618 ; n15621
g13186 and pi0129 n7301 ; n15622
g13187 and n6323 n15622 ; n15623
g13188 and pi0074 n15623_not ; n15624
g13189 and pi0054 n2611 ; n15625
g13190 and n8887 n15625 ; n15626
g13191 and pi0092 pi0129_not ; n15627
g13192 and pi0075 n15622 ; n15628
g13193 nor n2625 n8965 ; n15629
g13194 and n8887 n15629_not ; n15630
g13195 nor n2568 n15630 ; n15631
g13196 and pi0129 n6135 ; n15632
g13197 and pi0038 n15632_not ; n15633
g13198 and pi0039 n8887 ; n15634
g13199 nor n2729 n3106 ; n15635
g13200 and n2788 n2859_not ; n15636
g13201 and n2462 n15636_not ; n15637
g13202 and n2873 n15637_not ; n15638
g13203 and n2785 n15638_not ; n15639
g13204 and n2877 n15639_not ; n15640
g13205 and n2719 n15640_not ; n15641
g13206 nor n2722 n15641 ; n15642
g13207 nor pi0086 n15642 ; n15643
g13208 and n2783 n15643_not ; n15644
g13209 nor pi0097 n15644 ; n15645
g13210 nor n2776 n15645 ; n15646
g13211 nor pi0108 n15646 ; n15647
g13212 and n2775 n15647_not ; n15648
g13213 and n2889 n15648_not ; n15649
g13214 nor n2766 n15649 ; n15650
g13215 and n2765 n15650_not ; n15651
g13216 and n2764 n15651_not ; n15652
g13217 and po0740 n15652 ; n15653
g13218 and pi0250 n7474_not ; n15654
g13219 and n10077 n15654 ; n15655
g13220 and n2781 n15644_not ; n15656
g13221 nor n2776 n15656 ; n15657
g13222 nor pi0108 n15657 ; n15658
g13223 and n2775 n15658_not ; n15659
g13224 and n2889 n15659_not ; n15660
g13225 nor n2766 n15660 ; n15661
g13226 and n2765 n15661_not ; n15662
g13227 and n2764 n15662_not ; n15663
g13228 and po0740_not n15663 ; n15664
g13229 and n15653_not n15655 ; n15665
g13230 and n15664_not n15665 ; n15666
g13231 and pi0127_not n15652 ; n15667
g13232 and pi0127 n15663 ; n15668
g13233 nor n15655 n15667 ; n15669
g13234 and n15668_not n15669 ; n15670
g13235 nor n15666 n15670 ; n15671
g13236 and n2757 n15671_not ; n15672
g13237 and n3108 n15672_not ; n15673
g13238 and n2504 n15673_not ; n15674
g13239 and n15635 n15674_not ; n15675
g13240 nor pi0070 n15675 ; n15676
g13241 nor n3099 n15676 ; n15677
g13242 nor pi0051 n15677 ; n15678
g13243 and n2748 n15678_not ; n15679
g13244 and n3168 n15679_not ; n15680
g13245 nor n2745 n15680 ; n15681
g13246 and n2510 n15681_not ; n15682
g13247 and n3413 n15682_not ; n15683
g13248 nor pi0095 n15683 ; n15684
g13249 and pi0039_not pi0129 ; n15685
g13250 and n2741_not n15685 ; n15686
g13251 and n15684_not n15686 ; n15687
g13252 nor pi0038 n15634 ; n15688
g13253 and n15687_not n15688 ; n15689
g13254 nor n15633 n15689 ; n15690
g13255 and n2568 n15690_not ; n15691
g13256 nor pi0075 n15631 ; n15692
g13257 and n15691_not n15692 ; n15693
g13258 nor pi0092 n15628 ; n15694
g13259 and n15693_not n15694 ; n15695
g13260 and n13654 n15627_not ; n15696
g13261 and n15695_not n15696 ; n15697
g13262 nor pi0074 n15626 ; n15698
g13263 and n15697_not n15698 ; n15699
g13264 nor pi0055 n15624 ; n15700
g13265 and n15699_not n15700 ; n15701
g13266 and pi0055 n2570 ; n15702
g13267 and n15622 n15702 ; n15703
g13268 nor n15701 n15703 ; n15704
g13269 nor pi0056 n15704 ; n15705
g13270 nor n11310 n11318 ; n15706
g13271 and n15705_not n15706 ; n15707
g13272 nor n15621 n15707 ; n15708
g13273 and n3328 n15708_not ; n15709
g13274 nor n6120 n15620 ; n15710
g13275 and n15709_not n15710 ; po0284
g13276 nor n6130 n7347 ; n15712
g13277 and n8888 n10391 ; n15713
g13278 and po0740 n15713 ; n15714
g13279 nor pi0129 n15713 ; n15715
g13280 and n8967 n15714_not ; n15716
g13281 and n15715_not n15716 ; n15717
g13282 and n2521 n15717 ; n15718
g13283 nor pi0038 n3418 ; n15719
g13284 and n6137 n15719_not ; n15720
g13285 and n6280_not n6286 ; n15721
g13286 nor pi0087 n15721 ; n15722
g13287 and n15720_not n15722 ; n15723
g13288 and n6133 n15723_not ; n15724
g13289 and n6134 n15718_not ; n15725
g13290 and n15724_not n15725 ; n15726
g13291 nor n7305 n7341 ; n15727
g13292 and n15726_not n15727 ; n15728
g13293 and n8879 n15728_not ; n15729
g13294 and n15712 n15729_not ; n15730
g13295 nor pi0056 n15730 ; n15731
g13296 nor n6127 n15731 ; n15732
g13297 nor pi0062 n15732 ; n15733
g13298 nor n6299 n15733 ; n15734
g13299 and n3328 n15734_not ; n15735
g13300 and n6123 n15735_not ; po0286
g13301 and pi0087 n9747_not ; n15737
g13302 and n7473 n9022_not ; n15738
g13303 and n14596 n15738_not ; n15739
g13304 nor n15319 n15739 ; n15740
g13305 and n14455 n15740_not ; n15741
g13306 nor n15737 n15741 ; n15742
g13307 nor n14440 n15742 ; n15743
g13308 and pi0132_not n15329 ; n15744
g13309 and pi0130 n15744_not ; n15745
g13310 and pi0130_not n15744 ; n15746
g13311 nor n15745 n15746 ; n15747
g13312 nor n14429 n15747 ; n15748
g13313 and pi0100 n15740 ; n15749
g13314 and n2535 n15749_not ; n15750
g13315 and n10982_not n15739 ; n15751
g13316 nor pi0051 n15297 ; n15752
g13317 nor pi0232 n15752 ; n15753
g13318 and n10982 n15753_not ; n15754
g13319 nor pi0191 pi0299 ; n15755
g13320 nor pi0051 n15256 ; n15756
g13321 and pi0140 n15282 ; n15757
g13322 and n15756 n15757_not ; n15758
g13323 and n15755 n15758_not ; n15759
g13324 and pi0051_not n15263 ; n15760
g13325 and pi0140 n14657 ; n15761
g13326 and n15760 n15761_not ; n15762
g13327 and n9020 n15762_not ; n15763
g13328 and pi0169 n6197 ; n15764
g13329 and n9036_not n14596 ; n15765
g13330 and n15764_not n15765 ; n15766
g13331 and pi0162 n9036 ; n15767
g13332 nor pi0051 n14678 ; n15768
g13333 and n14657_not n15768 ; n15769
g13334 and pi0169 n15769_not ; n15770
g13335 nor pi0169 n15281 ; n15771
g13336 and n15767 n15771_not ; n15772
g13337 and n15770_not n15772 ; n15773
g13338 and n2521_not n15764 ; n15774
g13339 nor n14655 n15764 ; n15775
g13340 and pi0162_not n9036 ; n15776
g13341 and n15775_not n15776 ; n15777
g13342 and n15774_not n15777 ; n15778
g13343 and pi0299 n15766_not ; n15779
g13344 and n15778_not n15779 ; n15780
g13345 and n15773_not n15780 ; n15781
g13346 nor n15759 n15763 ; n15782
g13347 and n15781_not n15782 ; n15783
g13348 and pi0232 n15783_not ; n15784
g13349 and n15754 n15784_not ; n15785
g13350 nor pi0100 n15751 ; n15786
g13351 and n15785_not n15786 ; n15787
g13352 and n14467_not n15750 ; n15788
g13353 and n15787_not n15788 ; n15789
g13354 nor n15743 n15748 ; n15790
g13355 and n15789_not n15790 ; n15791
g13356 nor n14676 n15764 ; n15792
g13357 and pi0169 n14948 ; n15793
g13358 nor n15792 n15793 ; n15794
g13359 nor pi0216 n15794 ; n15795
g13360 and n14666_not n14962 ; n15796
g13361 and pi0169 n15796 ; n15797
g13362 nor pi0051 n14964 ; n15798
g13363 and pi0169_not n15798 ; n15799
g13364 and pi0162 pi0216 ; n15800
g13365 and n15797_not n15800 ; n15801
g13366 and n15799_not n15801 ; n15802
g13367 nor n15795 n15802 ; n15803
g13368 and n6379 n15803_not ; n15804
g13369 and pi0169 n14597 ; n15805
g13370 nor pi0051 n15805 ; n15806
g13371 nor n7570 n15767 ; n15807
g13372 and n15806_not n15807 ; n15808
g13373 nor n15804 n15808 ; n15809
g13374 and pi0299 n15809_not ; n15810
g13375 and n7551 n14675 ; n15811
g13376 nor pi0051 n15811 ; n15812
g13377 and pi0140_not n15812 ; n15813
g13378 and n14675 n14996 ; n15814
g13379 nor pi0051 n15814 ; n15815
g13380 and pi0140 n15815 ; n15816
g13381 and n15755 n15813_not ; n15817
g13382 and n15816_not n15817 ; n15818
g13383 nor n6197 n14676 ; n15819
g13384 nor n14948 n15819 ; n15820
g13385 and n7551 n15820_not ; n15821
g13386 nor n7551 n15319 ; n15822
g13387 nor n15821 n15822 ; n15823
g13388 and pi0140_not n15823 ; n15824
g13389 and pi0224 n15796_not ; n15825
g13390 nor pi0224 n15820 ; n15826
g13391 nor n15825 n15826 ; n15827
g13392 and n6405 n15827_not ; n15828
g13393 nor n6405 n15319 ; n15829
g13394 nor n15828 n15829 ; n15830
g13395 and pi0140 n15830 ; n15831
g13396 and n9020 n15824_not ; n15832
g13397 and n15831_not n15832 ; n15833
g13398 nor n15810 n15818 ; n15834
g13399 and n15833_not n15834 ; n15835
g13400 and pi0232 n15835_not ; n15836
g13401 and n14675 n14942 ; n15837
g13402 nor pi0051 n15837 ; n15838
g13403 nor pi0232 n15838 ; n15839
g13404 and pi0039 n15839_not ; n15840
g13405 and n15836_not n15840 ; n15841
g13406 nor pi0232 n14578 ; n15842
g13407 nor pi0039 n15842 ; n15843
g13408 and n6197_not n14578 ; n15844
g13409 nor n15070 n15844 ; n15845
g13410 nor n9022 n15845 ; n15846
g13411 and n9022 n14578 ; n15847
g13412 and pi0232 n15847_not ; n15848
g13413 and n15846_not n15848 ; n15849
g13414 and n15843 n15849_not ; n15850
g13415 nor n15841 n15850 ; n15851
g13416 nor pi0038 n15851 ; n15852
g13417 and pi0038 n15740_not ; n15853
g13418 nor pi0100 n15853 ; n15854
g13419 and n15852_not n15854 ; n15855
g13420 and n15750 n15855_not ; n15856
g13421 and n15742 n15748 ; n15857
g13422 and n15856_not n15857 ; n15858
g13423 nor n15791 n15858 ; n15859
g13424 nor po1038 n15859 ; n15860
g13425 and pi0087 n9705_not ; n15861
g13426 and pi0169 n7473 ; n15862
g13427 and pi0087_not n14596 ; n15863
g13428 and n15862_not n15863 ; n15864
g13429 nor pi0051 pi0087 ; n15865
g13430 and n15805_not n15865 ; n15866
g13431 and n15748 n15866 ; n15867
g13432 and po1038 n15861_not ; n15868
g13433 and n15864_not n15868 ; n15869
g13434 and n15867_not n15869 ; n15870
g13435 nor n15860 n15870 ; po0287
g13436 nor pi0100 n14009 ; n15872
g13437 nor pi0087 n7334 ; n15873
g13438 and n15872_not n15873 ; n15874
g13439 nor pi0075 n15874 ; n15875
g13440 nor n7302 n15875 ; n15876
g13441 nor pi0092 n15876 ; n15877
g13442 and n8880 n13654 ; n15878
g13443 and n15877_not n15878 ; po0288
g13444 and pi0164 n14920 ; n15880
g13445 and pi0051 pi0151_not ; n15881
g13446 nor n13752 n14443 ; n15882
g13447 nor n15881 n15882 ; n15883
g13448 and n14446 n15883 ; n15884
g13449 and pi0232 n15884 ; n15885
g13450 and pi0132 n15329_not ; n15886
g13451 nor n15744 n15886 ; n15887
g13452 nor n14430 n15887 ; n15888
g13453 and n14439 n15888_not ; n15889
g13454 nor n15885 n15889 ; n15890
g13455 nor pi0087 n15890 ; n15891
g13456 and po1038 n15880_not ; n15892
g13457 and n15891_not n15892 ; n15893
g13458 and pi0173 n14443 ; n15894
g13459 and pi0190 n14597 ; n15895
g13460 nor pi0299 n15894 ; n15896
g13461 and n15895_not n15896 ; n15897
g13462 and pi0299 n15884_not ; n15898
g13463 and pi0232 n15897_not ; n15899
g13464 and n15898_not n15899 ; n15900
g13465 and n14455 n15900_not ; n15901
g13466 and pi0087 n9030_not ; n15902
g13467 and n2608_not n15900 ; n15903
g13468 and n13752_not n14608 ; n15904
g13469 and pi0168 n14592 ; n15905
g13470 nor pi0151 n15905 ; n15906
g13471 and n15904_not n15906 ; n15907
g13472 nor n6197 n14608 ; n15908
g13473 and pi0168 n15049_not ; n15909
g13474 and n15908_not n15909 ; n15910
g13475 and n6197_not n14608 ; n15911
g13476 and n14613 n15911_not ; n15912
g13477 nor pi0168 n15912 ; n15913
g13478 and pi0151 n15910_not ; n15914
g13479 and n15913_not n15914 ; n15915
g13480 nor pi0160 n15907 ; n15916
g13481 and n15915_not n15916 ; n15917
g13482 and pi0151 n14578 ; n15918
g13483 nor pi0151 n14584 ; n15919
g13484 nor pi0168 n15918 ; n15920
g13485 and n15919_not n15920 ; n15921
g13486 and pi0168 n15881_not ; n15922
g13487 and n14506_not n15922 ; n15923
g13488 and n6197 n15923_not ; n15924
g13489 and n15921_not n15924 ; n15925
g13490 and pi0160 n15908_not ; n15926
g13491 and n15925_not n15926 ; n15927
g13492 and pi0299 n15917_not ; n15928
g13493 and n15927_not n15928 ; n15929
g13494 and pi0190 pi0299_not ; n15930
g13495 and pi0051 pi0173_not ; n15931
g13496 and pi0182 n14486 ; n15932
g13497 and n14505 n15932_not ; n15933
g13498 and n6197 n15931_not ; n15934
g13499 and n15933_not n15934 ; n15935
g13500 and n15930 n15935_not ; n15936
g13501 and n15911_not n15936 ; n15937
g13502 nor pi0190 pi0299 ; n15938
g13503 and pi0182_not n14608 ; n15939
g13504 and pi0182 n15908_not ; n15940
g13505 and n14585_not n15940 ; n15941
g13506 nor pi0173 n15939 ; n15942
g13507 and n15941_not n15942 ; n15943
g13508 nor pi0182 n15912 ; n15944
g13509 nor n14579 n15911 ; n15945
g13510 and pi0182 n15945_not ; n15946
g13511 and pi0173 n15944_not ; n15947
g13512 and n15946_not n15947 ; n15948
g13513 nor n15943 n15948 ; n15949
g13514 and n15938 n15949_not ; n15950
g13515 and pi0232 n15937_not ; n15951
g13516 and n15929_not n15951 ; n15952
g13517 and n15950_not n15952 ; n15953
g13518 and pi0232_not n14608 ; n15954
g13519 nor n15953 n15954 ; n15955
g13520 nor pi0039 n15955 ; n15956
g13521 and pi0183_not n14979 ; n15957
g13522 and pi0183 n15010_not ; n15958
g13523 nor pi0183 n14981 ; n15959
g13524 nor pi0173 n15959 ; n15960
g13525 and n15958_not n15960 ; n15961
g13526 nor pi0183 n14989 ; n15962
g13527 and pi0173 n14993_not ; n15963
g13528 and n15962_not n15963 ; n15964
g13529 nor n15957 n15964 ; n15965
g13530 and n15961_not n15965 ; n15966
g13531 and n15930 n15966_not ; n15967
g13532 nor pi0183 n7551 ; n15968
g13533 nor pi0173 n15968 ; n15969
g13534 and n15004 n15969 ; n15970
g13535 and pi0183 n14999 ; n15971
g13536 nor pi0183 n14443 ; n15972
g13537 and n14984_not n15972 ; n15973
g13538 and pi0173 n15973_not ; n15974
g13539 and n15971_not n15974 ; n15975
g13540 and n15938 n15970_not ; n15976
g13541 and n15975_not n15976 ; n15977
g13542 and pi0149_not pi0216 ; n15978
g13543 and n6379 n15978_not ; n15979
g13544 and n15884 n15979_not ; n15980
g13545 and pi0168_not n14776 ; n15981
g13546 and pi0168 n14659 ; n15982
g13547 nor pi0151 n15982 ; n15983
g13548 and n15981_not n15983 ; n15984
g13549 nor pi0168 n14965 ; n15985
g13550 and pi0168 n14962_not ; n15986
g13551 and pi0151 n15986_not ; n15987
g13552 and n15985_not n15987 ; n15988
g13553 and pi0149 n15984_not ; n15989
g13554 and n15988_not n15989 ; n15990
g13555 and pi0216 n15990_not ; n15991
g13556 and pi0168 n14949_not ; n15992
g13557 nor pi0168 n14951 ; n15993
g13558 nor n15992 n15993 ; n15994
g13559 nor n15881 n15994 ; n15995
g13560 nor pi0216 n15995 ; n15996
g13561 and n6379 n15991_not ; n15997
g13562 and n15996_not n15997 ; n15998
g13563 and pi0299 n15980_not ; n15999
g13564 and n15998_not n15999 ; n16000
g13565 nor n15967 n15977 ; n16001
g13566 and n16000_not n16001 ; n16002
g13567 and pi0232 n16002_not ; n16003
g13568 and n14945 n16003_not ; n16004
g13569 nor n15956 n16004 ; n16005
g13570 and n2608 n16005_not ; n16006
g13571 and n2535 n15903_not ; n16007
g13572 and n16006_not n16007 ; n16008
g13573 and n15888 n15902_not ; n16009
g13574 and n15901_not n16009 ; n16010
g13575 and n16008_not n16010 ; n16011
g13576 and n14456 n15900_not ; n16012
g13577 and n14439_not n15898 ; n16013
g13578 nor n13130 n16013 ; n16014
g13579 nor pi0168 n14667 ; n16015
g13580 and pi0168 n14673_not ; n16016
g13581 and pi0151 n16015_not ; n16017
g13582 and n16016_not n16017 ; n16018
g13583 and pi0168 n14677 ; n16019
g13584 nor n13752 n14654 ; n16020
g13585 nor pi0151 n16020 ; n16021
g13586 and n16019_not n16021 ; n16022
g13587 nor pi0149 n16022 ; n16023
g13588 and n16018_not n16023 ; n16024
g13589 nor n14714 n15883 ; n16025
g13590 nor pi0168 n16025 ; n16026
g13591 nor n14965 n15881 ; n16027
g13592 nor n14678 n16027 ; n16028
g13593 and pi0168 n16028_not ; n16029
g13594 and pi0149 n16026_not ; n16030
g13595 and n16029_not n16030 ; n16031
g13596 and n9036 n16024_not ; n16032
g13597 and n16031_not n16032 ; n16033
g13598 nor n16014 n16033 ; n16034
g13599 nor pi0183 n15271 ; n16035
g13600 and pi0183 n15279_not ; n16036
g13601 and pi0173 n16036_not ; n16037
g13602 and n16035_not n16037 ; n16038
g13603 and pi0183 n14683 ; n16039
g13604 nor pi0173 n16039 ; n16040
g13605 and n15263 n16040 ; n16041
g13606 nor n16038 n16041 ; n16042
g13607 and n15930 n16042_not ; n16043
g13608 and pi0183 n14714 ; n16044
g13609 and n15894_not n15938 ; n16045
g13610 and n15256_not n16045 ; n16046
g13611 and n16044_not n16046 ; n16047
g13612 nor n16034 n16047 ; n16048
g13613 and n16043_not n16048 ; n16049
g13614 and pi0232 n16049_not ; n16050
g13615 nor n15298 n16050 ; n16051
g13616 and pi0039 n16051_not ; n16052
g13617 and pi0232_not n14513 ; n16053
g13618 and pi0182 n15147 ; n16054
g13619 and n14513_not n16045 ; n16055
g13620 and n16054_not n16055 ; n16056
g13621 and pi0182_not n14537 ; n16057
g13622 nor n15146 n15931 ; n16058
g13623 and n16057_not n16058 ; n16059
g13624 and n15930 n16059_not ; n16060
g13625 and pi0168_not n14597 ; n16061
g13626 nor n15146 n16061 ; n16062
g13627 and pi0151 n16062_not ; n16063
g13628 nor pi0151 n15884 ; n16064
g13629 and n15147_not n16064 ; n16065
g13630 and pi0160 n16063_not ; n16066
g13631 and n16065_not n16066 ; n16067
g13632 nor pi0151 n14513 ; n16068
g13633 and pi0151 n14750 ; n16069
g13634 nor pi0168 n16068 ; n16070
g13635 and n16069_not n16070 ; n16071
g13636 and pi0151_not n14443 ; n16072
g13637 and pi0168 n16072_not ; n16073
g13638 and n14537_not n16073 ; n16074
g13639 nor n16071 n16074 ; n16075
g13640 nor pi0160 n15146 ; n16076
g13641 and n16075_not n16076 ; n16077
g13642 and pi0299 n16067_not ; n16078
g13643 and n16077_not n16078 ; n16079
g13644 and pi0232 n16056_not ; n16080
g13645 and n16060_not n16080 ; n16081
g13646 and n16079_not n16081 ; n16082
g13647 nor pi0039 n16053 ; n16083
g13648 and n16082_not n16083 ; n16084
g13649 and n2608 n16084_not ; n16085
g13650 and n16052_not n16085 ; n16086
g13651 and n2535 n15333_not ; n16087
g13652 and n15903_not n16087 ; n16088
g13653 and n16086_not n16088 ; n16089
g13654 nor n15888 n15902 ; n16090
g13655 and n16012_not n16090 ; n16091
g13656 and n16089_not n16091 ; n16092
g13657 nor po1038 n16092 ; n16093
g13658 and n16011_not n16093 ; n16094
g13659 or n15893 n16094 ; po0289
g13660 nor pi0133 n14909 ; n16096
g13661 and pi0145 n14714 ; n16097
g13662 and n15293 n16097_not ; n16098
g13663 and pi0197 n14657 ; n16099
g13664 and n15294 n16099_not ; n16100
g13665 and n14439 n16100_not ; n16101
g13666 and pi0299 n16101_not ; n16102
g13667 nor n16098 n16102 ; n16103
g13668 and pi0232 n16103_not ; n16104
g13669 and n15299 n16104_not ; n16105
g13670 and n9212_not n14503 ; n16106
g13671 and pi0039_not n14439 ; n16107
g13672 and n16106_not n16107 ; n16108
g13673 nor pi0038 n16108 ; n16109
g13674 and n16105_not n16109 ; n16110
g13675 and n14473 n16110_not ; n16111
g13676 and n14468 n16111_not ; n16112
g13677 nor n14456 n16112 ; n16113
g13678 nor n16096 n16113 ; n16114
g13679 nor pi0183 pi0299 ; n16115
g13680 and pi0149_not pi0299 ; n16116
g13681 nor n16115 n16116 ; n16117
g13682 and n7473 n16117 ; n16118
g13683 and pi0087 n16118_not ; n16119
g13684 and n9209_not n14532 ; n16120
g13685 nor n6197 n14532 ; n16121
g13686 nor n14585 n16121 ; n16122
g13687 and n9209 n16122 ; n16123
g13688 and pi0039_not pi0176 ; n16124
g13689 and n16120_not n16124 ; n16125
g13690 and n16123_not n16125 ; n16126
g13691 nor n5777 n16099 ; n16127
g13692 and n6640 n16127_not ; n16128
g13693 nor pi0145 n7551 ; n16129
g13694 nor pi0299 n16129 ; n16130
g13695 and n15003_not n16130 ; n16131
g13696 nor n16128 n16131 ; n16132
g13697 and n2521 n16132_not ; n16133
g13698 and pi0232 n16133_not ; n16134
g13699 nor n14944 n16134 ; n16135
g13700 and pi0039 n16135_not ; n16136
g13701 and pi0154 pi0232 ; n16137
g13702 and pi0299 n16137 ; n16138
g13703 and n14532 n16138_not ; n16139
g13704 and n16122 n16138 ; n16140
g13705 nor pi0039 pi0176 ; n16141
g13706 and n16139_not n16141 ; n16142
g13707 and n16140_not n16142 ; n16143
g13708 and n11374 n16136_not ; n16144
g13709 and n16126_not n16144 ; n16145
g13710 and n16143_not n16145 ; n16146
g13711 and pi0087_not n16096 ; n16147
g13712 and n16146_not n16147 ; n16148
g13713 nor n16114 n16119 ; n16149
g13714 and n16148_not n16149 ; n16150
g13715 nor po1038 n16150 ; n16151
g13716 and pi0149 n14920 ; n16152
g13717 and n14440 n16096_not ; n16153
g13718 and po1038 n16152_not ; n16154
g13719 and n16153_not n16154 ; n16155
g13720 or n16151 n16155 ; po0290
g13721 and po1038 n15865 ; n16157
g13722 and pi0136_not n15746 ; n16158
g13723 and pi0135_not n16158 ; n16159
g13724 and pi0134 n16159_not ; n16160
g13725 and n14438 n16160_not ; n16161
g13726 and pi0171 n6197 ; n16162
g13727 and n14438_not n16162 ; n16163
g13728 and pi0232 n16163 ; n16164
g13729 and n16157 n16164_not ; n16165
g13730 and n16161_not n16165 ; n16166
g13731 and pi0192 pi0299_not ; n16167
g13732 and pi0171 pi0299 ; n16168
g13733 nor n16167 n16168 ; n16169
g13734 and n7473 n16169_not ; n16170
g13735 and n14596 n16170_not ; n16171
g13736 nor n15319 n16171 ; n16172
g13737 and n14455 n16172_not ; n16173
g13738 and n2608_not n16172 ; n16174
g13739 and n2535 n16174_not ; n16175
g13740 nor pi0051 n16163 ; n16176
g13741 and pi0164_not pi0216 ; n16177
g13742 and n6379 n16177_not ; n16178
g13743 nor n16176 n16178 ; n16179
g13744 nor n14676 n16162 ; n16180
g13745 and pi0171 n14948 ; n16181
g13746 nor n16180 n16181 ; n16182
g13747 nor pi0216 n16182 ; n16183
g13748 and pi0171 n15796 ; n16184
g13749 and pi0171_not n15798 ; n16185
g13750 and pi0164 pi0216 ; n16186
g13751 and n16184_not n16186 ; n16187
g13752 and n16185_not n16187 ; n16188
g13753 nor n16183 n16188 ; n16189
g13754 and n6379 n16189_not ; n16190
g13755 nor n16179 n16190 ; n16191
g13756 and pi0299 n16191_not ; n16192
g13757 nor pi0192 pi0299 ; n16193
g13758 and n15812_not n16193 ; n16194
g13759 and pi0039 pi0186 ; n16195
g13760 and n15823_not n16167 ; n16196
g13761 nor n16194 n16195 ; n16197
g13762 and n16196_not n16197 ; n16198
g13763 and n15815_not n16193 ; n16199
g13764 and n15830_not n16167 ; n16200
g13765 and pi0186 n16199_not ; n16201
g13766 and n16200_not n16201 ; n16202
g13767 nor n16198 n16202 ; n16203
g13768 nor n16192 n16203 ; n16204
g13769 and pi0232 n16204_not ; n16205
g13770 and n15840 n16205_not ; n16206
g13771 and pi0232 n16169_not ; n16207
g13772 nor n14578 n16207 ; n16208
g13773 and n15845 n16207 ; n16209
g13774 nor pi0039 n16208 ; n16210
g13775 and n16209_not n16210 ; n16211
g13776 and n2608 n16206_not ; n16212
g13777 and n16211_not n16212 ; n16213
g13778 and n16175 n16213_not ; n16214
g13779 and n16160 n16173_not ; n16215
g13780 and n16214_not n16215 ; n16216
g13781 and n14455 n16171 ; n16217
g13782 and pi0039 pi0186_not ; n16218
g13783 and n15760_not n16167 ; n16219
g13784 and n15756_not n16193 ; n16220
g13785 nor n16219 n16220 ; n16221
g13786 and n15765 n16162_not ; n16222
g13787 and pi0299 n16222_not ; n16223
g13788 nor n14655 n16162 ; n16224
g13789 and n4192 n6197 ; n16225
g13790 and n9036 n16224_not ; n16226
g13791 and n16225_not n16226 ; n16227
g13792 and n16223 n16227_not ; n16228
g13793 and n16221 n16228_not ; n16229
g13794 and pi0232 n16229_not ; n16230
g13795 nor n15753 n16230 ; n16231
g13796 and n16218 n16231_not ; n16232
g13797 nor pi0039 n16171 ; n16233
g13798 and n14657_not n15760 ; n16234
g13799 and n16167 n16234_not ; n16235
g13800 and n15282_not n15756 ; n16236
g13801 and n16193 n16236_not ; n16237
g13802 nor n16235 n16237 ; n16238
g13803 and n16228_not n16238 ; n16239
g13804 and pi0232 n16239_not ; n16240
g13805 nor n15753 n16240 ; n16241
g13806 and n16195 n16241_not ; n16242
g13807 nor pi0164 n16233 ; n16243
g13808 and n16232_not n16243 ; n16244
g13809 and n16242_not n16244 ; n16245
g13810 nor pi0171 n15281 ; n16246
g13811 and pi0171 n15769_not ; n16247
g13812 and n9036 n16246_not ; n16248
g13813 and n16247_not n16248 ; n16249
g13814 and n16223 n16249_not ; n16250
g13815 and n16221 n16250_not ; n16251
g13816 and pi0232 n16251_not ; n16252
g13817 nor n15753 n16252 ; n16253
g13818 and n16218 n16253_not ; n16254
g13819 and n16238 n16250_not ; n16255
g13820 and pi0232 n16255_not ; n16256
g13821 nor n15753 n16256 ; n16257
g13822 and n16195 n16257_not ; n16258
g13823 and pi0164 n16233_not ; n16259
g13824 and n16254_not n16259 ; n16260
g13825 and n16258_not n16260 ; n16261
g13826 and n2608 n16245_not ; n16262
g13827 and n16261_not n16262 ; n16263
g13828 and n15333_not n16175 ; n16264
g13829 and n16263_not n16264 ; n16265
g13830 nor n16160 n16217 ; n16266
g13831 and n16265_not n16266 ; n16267
g13832 nor po1038 n16216 ; n16268
g13833 and n16267_not n16268 ; n16269
g13834 or n16166 n16269 ; po0291
g13835 and pi0135 n16158_not ; n16271
g13836 and pi0134 n16159 ; n16272
g13837 nor n16271 n16272 ; n16273
g13838 and pi0170 n6197 ; n16274
g13839 and n10598 n16274 ; n16275
g13840 and n14596 n16275_not ; n16276
g13841 and pi0194 n9193 ; n16277
g13842 and n16276 n16277_not ; n16278
g13843 and n14455 n16278 ; n16279
g13844 and pi0185 n15282 ; n16280
g13845 and n15756 n16280_not ; n16281
g13846 and n10982_not n16276 ; n16282
g13847 nor pi0194 n16282 ; n16283
g13848 and n16281_not n16283 ; n16284
g13849 and pi0185_not n15760 ; n16285
g13850 and pi0170 n7473 ; n16286
g13851 nor n9193 n16286 ; n16287
g13852 and n14596 n16287 ; n16288
g13853 and n10982_not n16288 ; n16289
g13854 and pi0194 n16289_not ; n16290
g13855 and n16234_not n16290 ; n16291
g13856 and n16285_not n16291 ; n16292
g13857 nor n16284 n16292 ; n16293
g13858 nor pi0299 n16293 ; n16294
g13859 and n15765 n16274_not ; n16295
g13860 and pi0150 pi0299 ; n16296
g13861 nor pi0170 n15281 ; n16297
g13862 and pi0170 n15769_not ; n16298
g13863 and n9036 n16297_not ; n16299
g13864 and n16298_not n16299 ; n16300
g13865 and n16296 n16300_not ; n16301
g13866 nor n14655 n16274 ; n16302
g13867 and n4415 n6197 ; n16303
g13868 and n9036 n16302_not ; n16304
g13869 and n16303_not n16304 ; n16305
g13870 and n15598 n16305_not ; n16306
g13871 nor n16301 n16306 ; n16307
g13872 nor n16283 n16290 ; n16308
g13873 nor n16295 n16308 ; n16309
g13874 and n16307_not n16309 ; n16310
g13875 nor n16294 n16310 ; n16311
g13876 and pi0232 n16311_not ; n16312
g13877 nor n15754 n16308 ; n16313
g13878 nor n16312 n16313 ; n16314
g13879 nor pi0100 n16314 ; n16315
g13880 nor n15319 n16278 ; n16316
g13881 and pi0100 n16316 ; n16317
g13882 and n2535 n16317_not ; n16318
g13883 and n14467_not n16318 ; n16319
g13884 and n16315_not n16319 ; n16320
g13885 and n16273 n16279_not ; n16321
g13886 and n16320_not n16321 ; n16322
g13887 nor n15319 n16276 ; n16323
g13888 and pi0038 n16323_not ; n16324
g13889 and n14438_not n16274 ; n16325
g13890 nor pi0051 n16325 ; n16326
g13891 and n6379_not n16326 ; n16327
g13892 and pi0170 n14948 ; n16328
g13893 nor n14676 n16274 ; n16329
g13894 and n7570 n16328_not ; n16330
g13895 and n16329_not n16330 ; n16331
g13896 nor n9036 n16331 ; n16332
g13897 and pi0170_not n15798 ; n16333
g13898 and pi0170 n15796 ; n16334
g13899 and pi0216 n16334_not ; n16335
g13900 and n16333_not n16335 ; n16336
g13901 nor n16332 n16336 ; n16337
g13902 and n16296 n16327_not ; n16338
g13903 and n16337_not n16338 ; n16339
g13904 and n7570_not n16326 ; n16340
g13905 and n15598 n16340_not ; n16341
g13906 and n16331_not n16341 ; n16342
g13907 nor n16339 n16342 ; n16343
g13908 and pi0185_not n15812 ; n16344
g13909 and pi0185 n15815 ; n16345
g13910 nor pi0299 n16344 ; n16346
g13911 and n16345_not n16346 ; n16347
g13912 and n16343 n16347_not ; n16348
g13913 and pi0232 n16348_not ; n16349
g13914 and n15840 n16349_not ; n16350
g13915 nor pi0299 n14578 ; n16351
g13916 and pi0170 n15845_not ; n16352
g13917 and pi0170_not n14578 ; n16353
g13918 and n10598 n16353_not ; n16354
g13919 and n16352_not n16354 ; n16355
g13920 and n15843 n16355_not ; n16356
g13921 and n16351_not n16356 ; n16357
g13922 nor n16350 n16357 ; n16358
g13923 nor pi0038 n16358 ; n16359
g13924 nor pi0194 n16324 ; n16360
g13925 and n16359_not n16360 ; n16361
g13926 nor n15319 n16288 ; n16362
g13927 and pi0038 n16362_not ; n16363
g13928 and pi0185_not n15823 ; n16364
g13929 and pi0185 n15830 ; n16365
g13930 nor pi0299 n16364 ; n16366
g13931 and n16365_not n16366 ; n16367
g13932 and n16343 n16367_not ; n16368
g13933 and pi0232 n16368_not ; n16369
g13934 and n15840 n16369_not ; n16370
g13935 and n10602 n15845 ; n16371
g13936 and n16356 n16371_not ; n16372
g13937 nor n16370 n16372 ; n16373
g13938 nor pi0038 n16373 ; n16374
g13939 and pi0194 n16363_not ; n16375
g13940 and n16374_not n16375 ; n16376
g13941 nor n16361 n16376 ; n16377
g13942 nor pi0100 n16377 ; n16378
g13943 and n16318 n16378_not ; n16379
g13944 and n14455 n16316_not ; n16380
g13945 nor n16273 n16380 ; n16381
g13946 and n16379_not n16381 ; n16382
g13947 nor po1038 n16322 ; n16383
g13948 and n16382_not n16383 ; n16384
g13949 and n14438 n16273 ; n16385
g13950 and n14438_not n16286 ; n16386
g13951 and n16157 n16386_not ; n16387
g13952 and n16385_not n16387 ; n16388
g13953 or n16384 n16388 ; po0292
g13954 and pi0136 n15746_not ; n16390
g13955 nor n16158 n16390 ; n16391
g13956 nor n14428 n16391 ; n16392
g13957 and n14596_not n16392 ; n16393
g13958 and pi0148 n7473 ; n16394
g13959 nor n14438 n16394 ; n16395
g13960 nor n16393 n16395 ; n16396
g13961 and n16157 n16396_not ; n16397
g13962 and n9739 n14438_not ; n16398
g13963 nor pi0051 n16398 ; n16399
g13964 and n14455 n16399 ; n16400
g13965 nor n2608 n16399 ; n16401
g13966 nor n9738 n15845 ; n16402
g13967 and n9738 n14578 ; n16403
g13968 and pi0232 n16403_not ; n16404
g13969 and n16402_not n16404 ; n16405
g13970 and n15843 n16405_not ; n16406
g13971 and pi0184_not n15823 ; n16407
g13972 and pi0184 n15830 ; n16408
g13973 and n9736 n16407_not ; n16409
g13974 and n16408_not n16409 ; n16410
g13975 nor pi0141 pi0299 ; n16411
g13976 and pi0184_not n15812 ; n16412
g13977 and pi0184 n15815 ; n16413
g13978 and n16411 n16412_not ; n16414
g13979 and n16413_not n16414 ; n16415
g13980 and pi0287_not n13665 ; n16416
g13981 and pi0216 n16416_not ; n16417
g13982 and n6379 n16417_not ; n16418
g13983 and n14675 n16418 ; n16419
g13984 nor pi0051 pi0148 ; n16420
g13985 and n16419_not n16420 ; n16421
g13986 and n6379_not n15319 ; n16422
g13987 nor n7570 n15319 ; n16423
g13988 nor pi0163 n16423 ; n16424
g13989 and pi0163 n6379 ; n16425
g13990 and n15796 n16425 ; n16426
g13991 nor n16422 n16424 ; n16427
g13992 and n16426_not n16427 ; n16428
g13993 and n7570 n15820_not ; n16429
g13994 and pi0148 n16428_not ; n16430
g13995 and n16429_not n16430 ; n16431
g13996 and pi0299 n16421_not ; n16432
g13997 and n16431_not n16432 ; n16433
g13998 nor n16415 n16433 ; n16434
g13999 and n16410_not n16434 ; n16435
g14000 and pi0232 n16435_not ; n16436
g14001 and n15840 n16436_not ; n16437
g14002 and n2608 n16437_not ; n16438
g14003 and n16406_not n16438 ; n16439
g14004 and n2535 n16401_not ; n16440
g14005 and n16439_not n16440 ; n16441
g14006 and n16392 n16400_not ; n16442
g14007 and n16441_not n16442 ; n16443
g14008 and n14438_not n16400 ; n16444
g14009 nor n11211 n14438 ; n16445
g14010 and n16399 n16445 ; n16446
g14011 and pi0184 n15282 ; n16447
g14012 and n15756 n16447_not ; n16448
g14013 and n16411 n16448_not ; n16449
g14014 and pi0184 n14657 ; n16450
g14015 and n15760 n16450_not ; n16451
g14016 and n9736 n16451_not ; n16452
g14017 and n6197_not n15765 ; n16453
g14018 and n9036 n15768 ; n16454
g14019 and pi0148 n16453_not ; n16455
g14020 and n16454_not n16455 ; n16456
g14021 and pi0051_not n15294 ; n16457
g14022 nor pi0148 n16457 ; n16458
g14023 nor n16416 n16458 ; n16459
g14024 and pi0148_not n14596 ; n16460
g14025 nor n16459 n16460 ; n16461
g14026 nor n16456 n16461 ; n16462
g14027 and pi0299 n16462_not ; n16463
g14028 nor n16449 n16452 ; n16464
g14029 and n16463_not n16464 ; n16465
g14030 and pi0232 n16465_not ; n16466
g14031 and pi0100_not n15754 ; n16467
g14032 and n16466_not n16467 ; n16468
g14033 nor n16446 n16468 ; n16469
g14034 and n2535 n16469_not ; n16470
g14035 nor n16392 n16444 ; n16471
g14036 and n16470_not n16471 ; n16472
g14037 nor po1038 n16472 ; n16473
g14038 and n16443_not n16473 ; n16474
g14039 or n16397 n16474 ; po0293
g14040 and pi0039_not pi0137 ; n16476
g14041 and n10368 n14873 ; n16477
g14042 and n6168 n11568 ; n16478
g14043 nor pi0299 po1038 ; n16479
g14044 and pi0198_not n11579 ; n16480
g14045 and n16479 n16480 ; n16481
g14046 nor n16478 n16481 ; n16482
g14047 nor n16477 n16482 ; n16483
g14048 and pi0210_not n11568 ; n16484
g14049 and po1038 n16484 ; n16485
g14050 nor n16483 n16485 ; n16486
g14051 and n10478 n16486_not ; n16487
g14052 or n16476 n16487 ; po0294
g14053 and n9739_not n13910 ; n16489
g14054 nor pi0039 n16489 ; n16490
g14055 nor pi0232 n11481 ; n16491
g14056 and n6198 n6396 ; n16492
g14057 and n9051 n16492 ; n16493
g14058 and n9736 n16493_not ; n16494
g14059 and n6198_not n9737 ; n16495
g14060 nor n9736 n11481 ; n16496
g14061 nor n16494 n16495 ; n16497
g14062 and n16496_not n16497 ; n16498
g14063 and pi0232 n16498_not ; n16499
g14064 nor n16491 n16499 ; n16500
g14065 and pi0039 n16500_not ; n16501
g14066 and n10200 n16490_not ; n16502
g14067 and n16501_not n16502 ; n16503
g14068 and pi0138_not n16503 ; n16504
g14069 and n9250 n9282_not ; n16505
g14070 and pi0092 n16505_not ; n16506
g14071 and n2532 n16506_not ; n16507
g14072 nor pi0075 n9288 ; n16508
g14073 nor n9326 n11892 ; n16509
g14074 and n9337 n16509_not ; n16510
g14075 and n13815 n16510_not ; n16511
g14076 nor n6242 n9326 ; n16512
g14077 and n9036 n16509_not ; n16513
g14078 and n16512_not n16513 ; n16514
g14079 and n9291 n16514_not ; n16515
g14080 nor n16511 n16515 ; n16516
g14081 nor pi0232 n16516 ; n16517
g14082 and pi0141_not n16511 ; n16518
g14083 and n9305_not n16510 ; n16519
g14084 and n13815 n16519_not ; n16520
g14085 and pi0141 n16520 ; n16521
g14086 nor n9300 n16509 ; n16522
g14087 nor n9290 n16522 ; n16523
g14088 and pi0148 n16523_not ; n16524
g14089 nor n9737 n16515 ; n16525
g14090 nor n16524 n16525 ; n16526
g14091 nor n16518 n16521 ; n16527
g14092 and n16526_not n16527 ; n16528
g14093 and pi0232 n16528_not ; n16529
g14094 nor n16517 n16529 ; n16530
g14095 and pi0039 n16530_not ; n16531
g14096 and pi0299 n9605_not ; n16532
g14097 nor pi0299 n9949 ; n16533
g14098 nor pi0232 n16532 ; n16534
g14099 and n16533_not n16534 ; n16535
g14100 nor pi0039 n16535 ; n16536
g14101 nor n6197 n9949 ; n16537
g14102 nor n13772 n16537 ; n16538
g14103 nor pi0299 n16538 ; n16539
g14104 and pi0141 n16539 ; n16540
g14105 and pi0148 n6197 ; n16541
g14106 nor n9605 n16541 ; n16542
g14107 and pi0148 n13737 ; n16543
g14108 nor n16542 n16543 ; n16544
g14109 and pi0299 n16544_not ; n16545
g14110 and pi0141_not n16533 ; n16546
g14111 and pi0232 n16546_not ; n16547
g14112 and n16540_not n16547 ; n16548
g14113 and n16545_not n16548 ; n16549
g14114 and n16536 n16549_not ; n16550
g14115 and n2608 n16531_not ; n16551
g14116 and n16550_not n16551 ; n16552
g14117 nor pi0087 n16552 ; n16553
g14118 and n16508 n16553_not ; n16554
g14119 nor pi0092 n16554 ; n16555
g14120 and n16507 n16555_not ; n16556
g14121 nor pi0055 n16556 ; n16557
g14122 and n9251 n13686_not ; n16558
g14123 and pi0055 n16558_not ; n16559
g14124 nor n16557 n16559 ; n16560
g14125 and n2529 n16560_not ; n16561
g14126 and n9883 n16561_not ; n16562
g14127 and pi0138 n16562 ; n16563
g14128 and pi0118_not n13664 ; n16564
g14129 and pi0139_not n16564 ; n16565
g14130 nor n16504 n16565 ; n16566
g14131 and n16563_not n16566 ; n16567
g14132 nor pi0138 n8974 ; n16568
g14133 and n16503 n16568_not ; n16569
g14134 and n16562 n16568 ; n16570
g14135 and n16565 n16569_not ; n16571
g14136 and n16570_not n16571 ; n16572
g14137 nor n16567 n16572 ; po0295
g14138 and n13910 n15738_not ; n16574
g14139 nor pi0039 n16574 ; n16575
g14140 and n11477_not n15755 ; n16576
g14141 and n6198_not n9021 ; n16577
g14142 and n9020 n16493_not ; n16578
g14143 nor n11480 n16577 ; n16579
g14144 nor n16576 n16578 ; n16580
g14145 and n16579 n16580 ; n16581
g14146 and pi0232 n16581_not ; n16582
g14147 nor n16491 n16582 ; n16583
g14148 and pi0039 n16583_not ; n16584
g14149 and n10200 n16575_not ; n16585
g14150 and n16584_not n16585 ; n16586
g14151 and pi0139_not n16586 ; n16587
g14152 and pi0169_not n9326 ; n16588
g14153 nor n16522 n16588 ; n16589
g14154 and n9036 n16589_not ; n16590
g14155 and n9291 n16590_not ; n16591
g14156 and pi0191_not n16511 ; n16592
g14157 and pi0191 n16520 ; n16593
g14158 nor n16591 n16592 ; n16594
g14159 and n16593_not n16594 ; n16595
g14160 and pi0232 n16595_not ; n16596
g14161 nor n16517 n16596 ; n16597
g14162 and pi0039 n16597_not ; n16598
g14163 and pi0191 n16539 ; n16599
g14164 nor n9605 n15764 ; n16600
g14165 and pi0169 n13737 ; n16601
g14166 nor n16600 n16601 ; n16602
g14167 and pi0299 n16602_not ; n16603
g14168 and pi0191_not n16533 ; n16604
g14169 and pi0232 n16604_not ; n16605
g14170 and n16599_not n16605 ; n16606
g14171 and n16603_not n16606 ; n16607
g14172 and n16536 n16607_not ; n16608
g14173 and n2608 n16598_not ; n16609
g14174 and n16608_not n16609 ; n16610
g14175 nor pi0087 n16610 ; n16611
g14176 and n16508 n16611_not ; n16612
g14177 nor pi0092 n16612 ; n16613
g14178 and n16507 n16613_not ; n16614
g14179 nor pi0055 n16614 ; n16615
g14180 nor n16559 n16615 ; n16616
g14181 and n2529 n16616_not ; n16617
g14182 and n9883 n16617_not ; n16618
g14183 and pi0139 n16618 ; n16619
g14184 nor n16564 n16587 ; n16620
g14185 and n16619_not n16620 ; n16621
g14186 nor pi0139 n8975 ; n16622
g14187 and n16586 n16622_not ; n16623
g14188 and n16618 n16622 ; n16624
g14189 and n16564 n16623_not ; n16625
g14190 and n16624_not n16625 ; n16626
g14191 nor n16621 n16626 ; po0296
g14192 and pi0641_not pi1158 ; n16628
g14193 and pi0641 pi1158_not ; n16629
g14194 nor n16628 n16629 ; n16630
g14195 and pi0788 n16630_not ; n16631
g14196 and pi0648_not pi1159 ; n16632
g14197 and pi0648 pi1159_not ; n16633
g14198 nor n16632 n16633 ; n16634
g14199 and pi0789 n16634_not ; n16635
g14200 and pi0627 pi1154 ; n16636
g14201 nor pi0627 pi1154 ; n16637
g14202 and pi0781 n16636_not ; n16638
g14203 and n16637_not n16638 ; n16639
g14204 and pi0140 n2571_not ; n16640
g14205 and n2926 n6284 ; n16641
g14206 nor pi0140 n16641 ; n16642
g14207 and pi0665 pi1091 ; n16643
g14208 and pi0680 n16643_not ; n16644
g14209 and n2926 n16644 ; n16645
g14210 and n6284 n16645 ; n16646
g14211 and pi0038 n16646_not ; n16647
g14212 and n16642_not n16647 ; n16648
g14213 and n6184_not n6380 ; n16649
g14214 nor pi0120 n16649 ; n16650
g14215 and pi0120 n2521_not ; n16651
g14216 nor n16650 n16651 ; n16652
g14217 and n2926 n16652 ; n16653
g14218 and n2603 n16653 ; n16654
g14219 and n16644 n16654 ; n16655
g14220 nor pi0661 pi0681 ; n16656
g14221 and pi0662_not n16656 ; n16657
g14222 and n16643_not n16653 ; n16658
g14223 and n6192_not n16658 ; n16659
g14224 nor pi0824 n16649 ; n16660
g14225 and n6380 n10204_not ; n16661
g14226 and pi1092 n16661 ; n16662
g14227 nor n11031 n16662 ; n16663
g14228 nor n16660 n16663 ; n16664
g14229 and pi1093 n16664 ; n16665
g14230 nor pi0120 n16665 ; n16666
g14231 and n2521 n2926 ; n16667
g14232 and pi0120 n16667_not ; n16668
g14233 nor pi1091 n16668 ; n16669
g14234 and n16666_not n16669 ; n16670
g14235 and n2926 n16649 ; n16671
g14236 and n2923 n16671 ; n16672
g14237 and pi0829 n16662_not ; n16673
g14238 nor pi0829 n16664 ; n16674
g14239 and n7517 n16673_not ; n16675
g14240 and n16674_not n16675 ; n16676
g14241 nor n16672 n16676 ; n16677
g14242 and pi1091 n16677_not ; n16678
g14243 nor pi0120 n16678 ; n16679
g14244 nor n16668 n16679 ; n16680
g14245 nor n16670 n16680 ; n16681
g14246 and n6197_not n16681 ; n16682
g14247 and n6197 n16653_not ; n16683
g14248 nor n16682 n16683 ; n16684
g14249 and pi0665 n16670_not ; n16685
g14250 nor n16681 n16685 ; n16686
g14251 nor n16658 n16686 ; n16687
g14252 and n16684 n16687_not ; n16688
g14253 and n6192 n16688 ; n16689
g14254 nor n16659 n16689 ; n16690
g14255 and n16657_not n16690 ; n16691
g14256 and n16657 n16688_not ; n16692
g14257 and pi0680 n16692_not ; n16693
g14258 and n16691_not n16693 ; n16694
g14259 and n6205 n16694_not ; n16695
g14260 and n6195 n16686 ; n16696
g14261 and n6197 n16681_not ; n16697
g14262 and n6197_not n16653 ; n16698
g14263 nor n16697 n16698 ; n16699
g14264 and n6192_not n16699 ; n16700
g14265 and n6192 n16681 ; n16701
g14266 nor n16700 n16701 ; n16702
g14267 and n16644 n16702 ; n16703
g14268 and n16657_not n16703 ; n16704
g14269 nor n16696 n16704 ; n16705
g14270 and n6205_not n16705 ; n16706
g14271 nor n2603 n16695 ; n16707
g14272 and n16706_not n16707 ; n16708
g14273 nor n16655 n16708 ; n16709
g14274 nor pi0223 n16709 ; n16710
g14275 and n6187 n14205 ; n16711
g14276 and n16667 n16711_not ; n16712
g14277 and pi0120 n16712_not ; n16713
g14278 nor pi0120 n16671 ; n16714
g14279 and pi1091 n16713_not ; n16715
g14280 and n16714_not n16715 ; n16716
g14281 and pi0120 pi0824 ; n16717
g14282 and n6187 n16717 ; n16718
g14283 and n16669 n16718_not ; n16719
g14284 and n16714_not n16719 ; n16720
g14285 nor n16716 n16720 ; n16721
g14286 and n6197 n16721_not ; n16722
g14287 nor n16698 n16722 ; n16723
g14288 and n6205_not n16723 ; n16724
g14289 and n6197_not n16721 ; n16725
g14290 and n16658 n16725_not ; n16726
g14291 nor n16659 n16726 ; n16727
g14292 and pi0680 n16727_not ; n16728
g14293 and n16724_not n16728 ; n16729
g14294 and n16657 n16726_not ; n16730
g14295 and pi0223 n16730_not ; n16731
g14296 and n16729 n16731 ; n16732
g14297 nor n16710 n16732 ; n16733
g14298 nor pi0299 n16733 ; n16734
g14299 and n6242_not n16705 ; n16735
g14300 and n6242 n16694_not ; n16736
g14301 nor n3448 n16735 ; n16737
g14302 and n16736_not n16737 ; n16738
g14303 and n16644 n16653 ; n16739
g14304 and n3448 n16739 ; n16740
g14305 nor n16738 n16740 ; n16741
g14306 nor pi0215 n16741 ; n16742
g14307 and n6242_not n16723 ; n16743
g14308 and n16728 n16743_not ; n16744
g14309 and pi0215 n16730_not ; n16745
g14310 and n16744 n16745 ; n16746
g14311 nor n16742 n16746 ; n16747
g14312 and pi0299 n16747_not ; n16748
g14313 nor n16734 n16748 ; n16749
g14314 and pi0140 n16749_not ; n16750
g14315 and pi0039 pi0140 ; n16751
g14316 and n16644_not n16654 ; n16752
g14317 nor pi0680 n16702 ; n16753
g14318 and n16643 n16680 ; n16754
g14319 and n6226_not n16754 ; n16755
g14320 and n16643 n16698 ; n16756
g14321 and n6192_not n16756 ; n16757
g14322 nor n16755 n16757 ; n16758
g14323 nor n16657 n16758 ; n16759
g14324 and n16657 n16754 ; n16760
g14325 and pi0680 n16760_not ; n16761
g14326 and n16759_not n16761 ; n16762
g14327 nor n16753 n16762 ; n16763
g14328 nor n6205 n16763 ; n16764
g14329 and pi0616 n16653_not ; n16765
g14330 and pi0614 n16653_not ; n16766
g14331 nor pi0603 n16653 ; n16767
g14332 and pi0603 n16684_not ; n16768
g14333 nor n16767 n16768 ; n16769
g14334 nor pi0642 n16769 ; n16770
g14335 nor n6190 n16653 ; n16771
g14336 nor n16770 n16771 ; n16772
g14337 nor pi0614 n16772 ; n16773
g14338 nor n16766 n16773 ; n16774
g14339 nor pi0616 n16774 ; n16775
g14340 nor n16765 n16775 ; n16776
g14341 nor pi0680 n16776 ; n16777
g14342 and n16643 n16653 ; n16778
g14343 and n6197 n16778_not ; n16779
g14344 nor n6197 n16754 ; n16780
g14345 nor n16779 n16780 ; n16781
g14346 and n6192 n16781 ; n16782
g14347 and n6192_not n16778 ; n16783
g14348 and pi0680 n16783_not ; n16784
g14349 and n16782_not n16784 ; n16785
g14350 nor n16777 n16785 ; n16786
g14351 and n16657_not n16786 ; n16787
g14352 and pi0680 n16781_not ; n16788
g14353 and n16657 n16788_not ; n16789
g14354 and n16777_not n16789 ; n16790
g14355 nor n16787 n16790 ; n16791
g14356 and n6205 n16791 ; n16792
g14357 nor n2603 n16764 ; n16793
g14358 and n16792_not n16793 ; n16794
g14359 nor pi0223 n16752 ; n16795
g14360 and n16794_not n16795 ; n16796
g14361 nor n16683 n16725 ; n16797
g14362 and n6190 n16797_not ; n16798
g14363 nor n16771 n16798 ; n16799
g14364 nor pi0614 n16799 ; n16800
g14365 nor n16766 n16800 ; n16801
g14366 nor pi0616 n16801 ; n16802
g14367 nor n16765 n16802 ; n16803
g14368 nor pi0680 n16803 ; n16804
g14369 and pi0665 n16716 ; n16805
g14370 nor n6197 n16805 ; n16806
g14371 nor n16779 n16806 ; n16807
g14372 and n6195 n16807_not ; n16808
g14373 and n16784 n16807_not ; n16809
g14374 nor n16808 n16809 ; n16810
g14375 and n16804_not n16810 ; n16811
g14376 and n6205 n16811 ; n16812
g14377 and pi0616_not n16800 ; n16813
g14378 nor n16723 n16813 ; n16814
g14379 nor pi0680 n16814 ; n16815
g14380 and pi0680 n16805_not ; n16816
g14381 and n16757_not n16816 ; n16817
g14382 nor n16815 n16817 ; n16818
g14383 and n16810 n16818 ; n16819
g14384 and n6205_not n16819 ; n16820
g14385 and pi0223 n16812_not ; n16821
g14386 and n16820_not n16821 ; n16822
g14387 nor n16796 n16822 ; n16823
g14388 nor pi0299 n16823 ; n16824
g14389 and n3448 n16652 ; n16825
g14390 and n2926 n16644_not ; n16826
g14391 and n16825 n16826 ; n16827
g14392 nor n6242 n16763 ; n16828
g14393 and n6242 n16791 ; n16829
g14394 nor n3448 n16828 ; n16830
g14395 and n16829_not n16830 ; n16831
g14396 nor pi0215 n16827 ; n16832
g14397 and n16831_not n16832 ; n16833
g14398 and n6242 n16811 ; n16834
g14399 and n6242_not n16819 ; n16835
g14400 and pi0215 n16834_not ; n16836
g14401 and n16835_not n16836 ; n16837
g14402 nor n16833 n16837 ; n16838
g14403 and pi0299 n16838_not ; n16839
g14404 nor n16824 n16839 ; n16840
g14405 and pi0039 n16840 ; n16841
g14406 nor n16751 n16841 ; n16842
g14407 nor n16750 n16842 ; n16843
g14408 nor pi0102 n11299 ; n16844
g14409 nor pi0098 n2787 ; n16845
g14410 and n16844_not n16845 ; n16846
g14411 and n7438 n12375 ; n16847
g14412 and n16846 n16847 ; n16848
g14413 and n8897 n9141 ; n16849
g14414 and n16848 n16849 ; n16850
g14415 nor pi0040 n16850 ; n16851
g14416 and n10289 n16851_not ; n16852
g14417 nor pi0252 n16852 ; n16853
g14418 and n2763 n2938 ; n16854
g14419 and n8896 n16848 ; n16855
g14420 nor pi0047 n16855 ; n16856
g14421 and pi0314 n10241 ; n16857
g14422 and n16856 n16857_not ; n16858
g14423 and n16854 n16858_not ; n16859
g14424 nor pi0035 n16859 ; n16860
g14425 and pi0040_not n10274 ; n16861
g14426 and n16860_not n16861 ; n16862
g14427 and pi0252 n2743_not ; n16863
g14428 and n16862_not n16863 ; n16864
g14429 nor n16853 n16864 ; n16865
g14430 and n2518 n16865 ; n16866
g14431 and pi1092 n12373_not ; n16867
g14432 and n16866 n16867 ; n16868
g14433 nor pi0088 n16846 ; n16869
g14434 and n11020 n16869_not ; n16870
g14435 and pi0252_not n9500 ; n16871
g14436 and n16870 n16871 ; n16872
g14437 and n2500 n16870 ; n16873
g14438 nor pi0047 n16857 ; n16874
g14439 and n16873_not n16874 ; n16875
g14440 and n16854 n16875_not ; n16876
g14441 nor pi0035 n16876 ; n16877
g14442 and pi0252 n10274 ; n16878
g14443 and n16877_not n16878 ; n16879
g14444 nor pi0040 n16872 ; n16880
g14445 and n16879_not n16880 ; n16881
g14446 and n7417 n10289 ; n16882
g14447 and n16881_not n16882 ; n16883
g14448 nor n16868 n16883 ; n16884
g14449 and pi1093 n16884_not ; n16885
g14450 nor n2923 n16885 ; n16886
g14451 and pi1092 n2930 ; n16887
g14452 and n2923 n16887 ; po1106
g14453 and n16866 po1106 ; n16889
g14454 nor n2924 n16889 ; n16890
g14455 nor n16886 n16890 ; n16891
g14456 and pi1091_not n16885 ; n16892
g14457 nor n16891 n16892 ; n16893
g14458 and pi0665 n16892_not ; n16894
g14459 nor n16893 n16894 ; n16895
g14460 nor pi0198 n16895 ; n16896
g14461 nor n3411 n16881 ; n16897
g14462 nor pi0032 n16897 ; n16898
g14463 and pi0032 n6485_not ; n16899
g14464 and pi0095_not n2932 ; n16900
g14465 and n16899_not n16900 ; n16901
g14466 and n16898_not n16901 ; n16902
g14467 and pi0824 n16902 ; n16903
g14468 nor n16868 n16903 ; n16904
g14469 and n7626 n16904_not ; n16905
g14470 nor pi0032 n16865 ; n16906
g14471 and n16901 n16906_not ; n16907
g14472 and pi0824_not pi0829 ; n16908
g14473 and n16907 n16908 ; n16909
g14474 and n16904 n16909_not ; n16910
g14475 and pi1093 n16910_not ; n16911
g14476 nor n2923 n16911 ; n16912
g14477 nor n16890 n16912 ; n16913
g14478 nor n16905 n16913 ; n16914
g14479 and pi0665 n16905_not ; n16915
g14480 nor n16914 n16915 ; n16916
g14481 and pi0198 n16916_not ; n16917
g14482 nor n16896 n16917 ; n16918
g14483 and pi0680 n16918 ; n16919
g14484 nor pi0299 n16919 ; n16920
g14485 and pi0210 n16916_not ; n16921
g14486 nor pi0210 n16895 ; n16922
g14487 nor n16921 n16922 ; n16923
g14488 and pi0680 n16923 ; n16924
g14489 and pi0299 n16924_not ; n16925
g14490 nor n16920 n16925 ; n16926
g14491 and pi0140 n16926 ; n16927
g14492 and pi0198_not n16893 ; n16928
g14493 and pi0198 n16914 ; n16929
g14494 nor n16928 n16929 ; n16930
g14495 and pi0665 n16913 ; n16931
g14496 and pi0198 n16931_not ; n16932
g14497 and pi0665 n16891 ; n16933
g14498 nor pi0198 n16933 ; n16934
g14499 nor n16932 n16934 ; n16935
g14500 and pi0680 n16935_not ; n16936
g14501 and n16930 n16936_not ; n16937
g14502 nor pi0299 n16937 ; n16938
g14503 and pi0210_not n16893 ; n16939
g14504 and pi0210 n16914 ; n16940
g14505 nor n16939 n16940 ; n16941
g14506 nor pi0210 n16933 ; n16942
g14507 and pi0210 n16931_not ; n16943
g14508 nor n16942 n16943 ; n16944
g14509 and pi0680 n16944_not ; n16945
g14510 and n16941 n16945_not ; n16946
g14511 and pi0299 n16946_not ; n16947
g14512 nor n16938 n16947 ; n16948
g14513 nor pi0140 n16948 ; n16949
g14514 nor pi0039 n16927 ; n16950
g14515 and n16949_not n16950 ; n16951
g14516 nor n16843 n16951 ; n16952
g14517 nor pi0038 n16952 ; n16953
g14518 nor pi0738 n16648 ; n16954
g14519 and n16953_not n16954 ; n16955
g14520 and pi0299 n16941_not ; n16956
g14521 nor pi0299 n16930 ; n16957
g14522 nor n16956 n16957 ; n16958
g14523 nor pi0039 n16958 ; n16959
g14524 and pi0681 n16814_not ; n16960
g14525 and pi0661 n16814 ; n16961
g14526 nor n6193 n16803 ; n16962
g14527 and n6193 n16721 ; n16963
g14528 nor n6197 n16963 ; n16964
g14529 and n16962_not n16964 ; n16965
g14530 nor n16722 n16965 ; n16966
g14531 nor pi0661 n16966 ; n16967
g14532 nor pi0681 n16961 ; n16968
g14533 and n16967_not n16968 ; n16969
g14534 nor n16960 n16969 ; n16970
g14535 nor n6205 n16970 ; n16971
g14536 and pi0681 n16803_not ; n16972
g14537 and pi0680 n16797_not ; n16973
g14538 nor pi0680 n16653 ; n16974
g14539 and pi0616 n16657 ; n16975
g14540 and n16974_not n16975 ; n16976
g14541 and n16973_not n16976 ; n16977
g14542 and pi0616 n16653 ; n16978
g14543 and n16657_not n16978 ; n16979
g14544 nor n16977 n16979 ; n16980
g14545 nor pi0616 n16657 ; n16981
g14546 and n16801 n16981 ; n16982
g14547 and pi0680_not n16802 ; n16983
g14548 and pi0616_not n16657 ; n16984
g14549 and n16973_not n16984 ; n16985
g14550 and n16983_not n16985 ; n16986
g14551 nor n16982 n16986 ; n16987
g14552 and pi0681_not n16980 ; n16988
g14553 and n16987 n16988 ; n16989
g14554 nor n16972 n16989 ; n16990
g14555 and n6205 n16990_not ; n16991
g14556 nor n16971 n16991 ; n16992
g14557 and pi0223 n16992_not ; n16993
g14558 and pi0681 n16776_not ; n16994
g14559 and pi0680 n16684_not ; n16995
g14560 and pi0614 n16657 ; n16996
g14561 and n16974_not n16996 ; n16997
g14562 and n16995_not n16997 ; n16998
g14563 and pi0614 n16653 ; n16999
g14564 and n16657_not n16999 ; n17000
g14565 nor n16998 n17000 ; n17001
g14566 nor pi0614 n6195 ; n17002
g14567 nor pi0616 n16772 ; n17003
g14568 and n16765_not n17002 ; n17004
g14569 and n17003_not n17004 ; n17005
g14570 and pi0614_not n6195 ; n17006
g14571 and n16684 n17006 ; n17007
g14572 nor n17005 n17007 ; n17008
g14573 and pi0681_not n17001 ; n17009
g14574 and n17008 n17009 ; n17010
g14575 nor n16994 n17010 ; n17011
g14576 and n6205 n17011_not ; n17012
g14577 and pi0681 n16702_not ; n17013
g14578 and n6194 n16681_not ; n17014
g14579 and n6194_not n16702 ; n17015
g14580 nor pi0681 n17014 ; n17016
g14581 and n17015_not n17016 ; n17017
g14582 nor n17013 n17017 ; n17018
g14583 nor n6205 n17018 ; n17019
g14584 nor n17012 n17019 ; n17020
g14585 and n2603_not n17020 ; n17021
g14586 nor pi0223 n16654 ; n17022
g14587 and n17021_not n17022 ; n17023
g14588 nor n16993 n17023 ; n17024
g14589 nor pi0299 n17024 ; n17025
g14590 and n3448 n16653 ; n17026
g14591 and n6241 n17011_not ; n17027
g14592 nor n6241 n17018 ; n17028
g14593 and n6236 n17028_not ; n17029
g14594 and n17027_not n17029 ; n17030
g14595 and n3448_not n17030 ; n17031
g14596 and n6236_not n17018 ; n17032
g14597 and n3448_not n17032 ; n17033
g14598 nor pi0215 n17026 ; n17034
g14599 and n17033_not n17034 ; n17035
g14600 and n17031_not n17035 ; n17036
g14601 and n6236_not n16970 ; n17037
g14602 nor n6241 n16970 ; n17038
g14603 and n6241 n16990_not ; n17039
g14604 and n6236 n17039_not ; n17040
g14605 and n17038_not n17040 ; n17041
g14606 nor n17037 n17041 ; n17042
g14607 and pi0215 n17042 ; n17043
g14608 nor n17036 n17043 ; n17044
g14609 and pi0299 n17044_not ; n17045
g14610 nor n17025 n17045 ; n17046
g14611 and pi0039 n17046_not ; n17047
g14612 nor n16959 n17047 ; n17048
g14613 nor pi0038 n17048 ; n17049
g14614 and n2926 n6135 ; n17050
g14615 and pi0038 n17050_not ; n17051
g14616 nor n17049 n17051 ; n17052
g14617 and pi0140_not pi0738 ; n17053
g14618 and n17052_not n17053 ; n17054
g14619 and n2571 n17054_not ; n17055
g14620 and n16955_not n17055 ; n17056
g14621 nor n16640 n17056 ; n17057
g14622 nor pi0778 n17057 ; n17058
g14623 and n2571 n17052 ; n17059
g14624 nor pi0140 n17059 ; n17060
g14625 and pi0625_not n17060 ; n17061
g14626 and pi0625 n17057 ; n17062
g14627 and pi1153 n17061_not ; n17063
g14628 and n17062_not n17063 ; n17064
g14629 and pi0625_not n17057 ; n17065
g14630 and pi0625 n17060 ; n17066
g14631 nor pi1153 n17066 ; n17067
g14632 and n17065_not n17067 ; n17068
g14633 nor n17064 n17068 ; n17069
g14634 and pi0778 n17069_not ; n17070
g14635 nor n17058 n17070 ; n17071
g14636 and pi0660 pi1155 ; n17072
g14637 nor pi0660 pi1155 ; n17073
g14638 and pi0785 n17072_not ; n17074
g14639 and n17073_not n17074 ; n17075
g14640 nor n17071 n17075 ; n17076
g14641 and n17060_not n17075 ; n17077
g14642 nor n17076 n17077 ; n17078
g14643 and n16639_not n17078 ; n17079
g14644 and n16639 n17060 ; n17080
g14645 nor n17079 n17080 ; n17081
g14646 and n16635_not n17081 ; n17082
g14647 and n16635 n17060_not ; n17083
g14648 nor n17082 n17083 ; n17084
g14649 and n16631_not n17084 ; n17085
g14650 and n16631 n17060 ; n17086
g14651 nor n17085 n17086 ; n17087
g14652 and pi0792_not n17087 ; n17088
g14653 and pi0628_not n17060 ; n17089
g14654 and pi0628 n17087_not ; n17090
g14655 and pi1156 n17089_not ; n17091
g14656 and n17090_not n17091 ; n17092
g14657 and pi0628 n17060 ; n17093
g14658 nor pi0628 n17087 ; n17094
g14659 nor pi1156 n17093 ; n17095
g14660 and n17094_not n17095 ; n17096
g14661 nor n17092 n17096 ; n17097
g14662 and pi0792 n17097_not ; n17098
g14663 nor n17088 n17098 ; n17099
g14664 nor pi0787 n17099 ; n17100
g14665 and pi0647_not n17060 ; n17101
g14666 and pi0647 n17099 ; n17102
g14667 and pi1157 n17101_not ; n17103
g14668 and n17102_not n17103 ; n17104
g14669 and pi0647_not n17099 ; n17105
g14670 and pi0647 n17060 ; n17106
g14671 nor pi1157 n17106 ; n17107
g14672 and n17105_not n17107 ; n17108
g14673 nor n17104 n17108 ; n17109
g14674 and pi0787 n17109_not ; n17110
g14675 nor n17100 n17110 ; n17111
g14676 and pi0644_not n17111 ; n17112
g14677 and pi0619_not n17060 ; n17113
g14678 and pi0608_not pi1153 ; n17114
g14679 and pi0608 pi1153_not ; n17115
g14680 nor n17114 n17115 ; n17116
g14681 and pi0778 n17116_not ; n17117
g14682 and pi0621 n16891 ; n17118
g14683 nor pi0210 n17118 ; n17119
g14684 and pi0621 n16913 ; n17120
g14685 and pi0210 n17120_not ; n17121
g14686 nor n17119 n17121 ; n17122
g14687 and pi0603 n17122_not ; n17123
g14688 and n16941 n17123_not ; n17124
g14689 and pi0299 n17124_not ; n17125
g14690 nor pi0198 n17118 ; n17126
g14691 and pi0198 n17120_not ; n17127
g14692 nor n17126 n17127 ; n17128
g14693 and pi0621 n16892_not ; n17129
g14694 nor n16893 n17129 ; n17130
g14695 and pi0198_not n17130 ; n17131
g14696 and pi0621 n16905_not ; n17132
g14697 nor n16914 n17132 ; n17133
g14698 and pi0198 n17133 ; n17134
g14699 nor n17131 n17134 ; n17135
g14700 nor pi0603 n17135 ; n17136
g14701 nor n17128 n17136 ; n17137
g14702 and pi0299_not n17137 ; n17138
g14703 nor n17125 n17138 ; n17139
g14704 nor pi0039 n17139 ; n17140
g14705 nor n6195 n16702 ; n17141
g14706 and n6195 n16681 ; n17142
g14707 nor n17141 n17142 ; n17143
g14708 and pi0621 pi1091 ; n17144
g14709 and n16680 n17144 ; n17145
g14710 and pi0621 n16670_not ; n17146
g14711 nor n16681 n17146 ; n17147
g14712 and pi0603_not n17147 ; n17148
g14713 and pi0603_not n16699 ; n17149
g14714 and n6197 n17145 ; n17150
g14715 and n16698 n17144 ; n17151
g14716 and pi0603 n17151_not ; n17152
g14717 and n17150_not n17152 ; n17153
g14718 nor n17149 n17153 ; n17154
g14719 nor n17145 n17148 ; n17155
g14720 and n17154_not n17155 ; n17156
g14721 and n17143 n17156_not ; n17157
g14722 nor n6242 n17157 ; n17158
g14723 and n16653 n17144 ; n17159
g14724 and n6197 n17159_not ; n17160
g14725 nor n6197 n17145 ; n17161
g14726 nor n17160 n17161 ; n17162
g14727 and pi0603 n17162_not ; n17163
g14728 and n16684 n17163_not ; n17164
g14729 and n6195 n17164_not ; n17165
g14730 nor pi0614 pi0642 ; n17166
g14731 and pi0616_not n17166 ; n17167
g14732 and pi0603 n17144_not ; n17168
g14733 and n16653 n17168_not ; n17169
g14734 and n17167_not n17169 ; n17170
g14735 and n16767_not n17167 ; n17171
g14736 and n17163_not n17171 ; n17172
g14737 nor n17170 n17172 ; n17173
g14738 and n6195_not n17173 ; n17174
g14739 nor n17165 n17174 ; n17175
g14740 and n6242 n17175_not ; n17176
g14741 nor n3448 n17158 ; n17177
g14742 and n17176_not n17177 ; n17178
g14743 and n3448 n17169 ; n17179
g14744 nor n17178 n17179 ; n17180
g14745 nor pi0215 n17180 ; n17181
g14746 and n2926 n17168_not ; n17182
g14747 and n16723_not n17182 ; n17183
g14748 and n6192 n16716_not ; n17184
g14749 and n17183 n17184_not ; n17185
g14750 nor n6195 n17185 ; n17186
g14751 and n16721_not n17182 ; n17187
g14752 and n6195 n17187_not ; n17188
g14753 nor n17186 n17188 ; n17189
g14754 nor n6242 n17189 ; n17190
g14755 and pi0621 n16716 ; n17191
g14756 nor n6197 n17191 ; n17192
g14757 nor n17160 n17192 ; n17193
g14758 and pi0603 n17193_not ; n17194
g14759 and n17171 n17194_not ; n17195
g14760 nor n17170 n17195 ; n17196
g14761 nor n6195 n17196 ; n17197
g14762 and n6195 n16797 ; n17198
g14763 and n17194_not n17198 ; n17199
g14764 nor n17197 n17199 ; n17200
g14765 and n6242 n17200 ; n17201
g14766 and pi0215 n17190_not ; n17202
g14767 and n17201_not n17202 ; n17203
g14768 nor n17181 n17203 ; n17204
g14769 and pi0299 n17204_not ; n17205
g14770 nor n6205 n17157 ; n17206
g14771 and n6205 n17175_not ; n17207
g14772 nor n2603 n17206 ; n17208
g14773 and n17207_not n17208 ; n17209
g14774 and n2603 n17169 ; n17210
g14775 nor n17209 n17210 ; n17211
g14776 nor pi0223 n17211 ; n17212
g14777 nor n6205 n17189 ; n17213
g14778 and n6205 n17200 ; n17214
g14779 and pi0223 n17213_not ; n17215
g14780 and n17214_not n17215 ; n17216
g14781 nor n17212 n17216 ; n17217
g14782 nor pi0299 n17217 ; n17218
g14783 nor n17205 n17218 ; n17219
g14784 and pi0039 n17219 ; n17220
g14785 nor n17140 n17220 ; n17221
g14786 and pi0761_not n17221 ; n17222
g14787 and pi0761 n17048 ; n17223
g14788 nor pi0140 n17222 ; n17224
g14789 and n17223_not n17224 ; n17225
g14790 and pi0603 n17135_not ; n17226
g14791 nor pi0299 n17226 ; n17227
g14792 nor pi0210 n17130 ; n17228
g14793 and pi0210 n17133_not ; n17229
g14794 nor n17228 n17229 ; n17230
g14795 and pi0603 n17230 ; n17231
g14796 and pi0299 n17231_not ; n17232
g14797 nor n17227 n17232 ; n17233
g14798 nor pi0039 n17233 ; n17234
g14799 and n16653 n17168 ; n17235
g14800 and n16725_not n17235 ; n17236
g14801 and n16723_not n17235 ; n17237
g14802 and n16725 n17167 ; n17238
g14803 and n17237 n17238_not ; n17239
g14804 and n6195_not n17239 ; n17240
g14805 nor n17236 n17240 ; n17241
g14806 nor n16743 n17241 ; n17242
g14807 and pi0215 n17242_not ; n17243
g14808 and n2926 n17168 ; n17244
g14809 and n16825 n17244 ; n17245
g14810 and n16684 n17168 ; n17246
g14811 and n6195 n17246 ; n17247
g14812 and n17167_not n17235 ; n17248
g14813 and n17167 n17246 ; n17249
g14814 nor n17248 n17249 ; n17250
g14815 nor n6195 n17250 ; n17251
g14816 nor n17247 n17251 ; n17252
g14817 and n6242 n17252 ; n17253
g14818 and n17143 n17168 ; n17254
g14819 nor n6242 n17254 ; n17255
g14820 nor n3448 n17253 ; n17256
g14821 and n17255_not n17256 ; n17257
g14822 nor pi0215 n17245 ; n17258
g14823 and n17257_not n17258 ; n17259
g14824 and pi0299 n17243_not ; n17260
g14825 and n17259_not n17260 ; n17261
g14826 nor n16724 n17241 ; n17262
g14827 and pi0223 n17262_not ; n17263
g14828 and n6205 n17252 ; n17264
g14829 nor n6205 n17254 ; n17265
g14830 nor n2603 n17264 ; n17266
g14831 and n17265_not n17266 ; n17267
g14832 and n16654 n17168 ; n17268
g14833 nor pi0223 n17268 ; n17269
g14834 and n17267_not n17269 ; n17270
g14835 nor pi0299 n17263 ; n17271
g14836 and n17270_not n17271 ; n17272
g14837 nor n17261 n17272 ; n17273
g14838 and pi0039 n17273 ; n17274
g14839 nor n17234 n17274 ; n17275
g14840 and pi0140 pi0761_not ; n17276
g14841 and n17275 n17276 ; n17277
g14842 nor n17225 n17277 ; n17278
g14843 nor pi0038 n17278 ; n17279
g14844 and n6284 n17244 ; n17280
g14845 and pi0761_not n17280 ; n17281
g14846 nor n16642 n17281 ; n17282
g14847 and pi0038 n17282_not ; n17283
g14848 nor n17279 n17283 ; n17284
g14849 and n2571 n17284 ; n17285
g14850 nor n16640 n17285 ; n17286
g14851 nor n17117 n17286 ; n17287
g14852 and n17060_not n17117 ; n17288
g14853 nor n17287 n17288 ; n17289
g14854 nor pi0785 n17289 ; n17290
g14855 and pi0609 n17117_not ; n17291
g14856 nor n17060 n17291 ; n17292
g14857 and pi0609 n17287 ; n17293
g14858 nor n17292 n17293 ; n17294
g14859 and pi1155 n17294_not ; n17295
g14860 nor pi0609 n17117 ; n17296
g14861 nor n17060 n17296 ; n17297
g14862 and pi0609_not n17287 ; n17298
g14863 nor n17297 n17298 ; n17299
g14864 nor pi1155 n17299 ; n17300
g14865 nor n17295 n17300 ; n17301
g14866 and pi0785 n17301_not ; n17302
g14867 nor n17290 n17302 ; n17303
g14868 nor pi0781 n17303 ; n17304
g14869 and pi0618_not n17060 ; n17305
g14870 and pi0618 n17303 ; n17306
g14871 and pi1154 n17305_not ; n17307
g14872 and n17306_not n17307 ; n17308
g14873 and pi0618_not n17303 ; n17309
g14874 and pi0618 n17060 ; n17310
g14875 nor pi1154 n17310 ; n17311
g14876 and n17309_not n17311 ; n17312
g14877 nor n17308 n17312 ; n17313
g14878 and pi0781 n17313_not ; n17314
g14879 nor n17304 n17314 ; n17315
g14880 and pi0619 n17315 ; n17316
g14881 and pi1159 n17113_not ; n17317
g14882 and n17316_not n17317 ; n17318
g14883 and pi0738 n17284_not ; n17319
g14884 and n16721_not n17235 ; n17320
g14885 nor n16805 n17320 ; n17321
g14886 and n6195 n17321 ; n17322
g14887 and pi0680 n16657_not ; n17323
g14888 nor n16756 n16805 ; n17324
g14889 and n17237_not n17324 ; n17325
g14890 and n17167_not n17325 ; n17326
g14891 and pi0603_not n16756 ; n17327
g14892 and n17321 n17327_not ; n17328
g14893 and n17167 n17328 ; n17329
g14894 nor n17326 n17329 ; n17330
g14895 and n17323 n17330_not ; n17331
g14896 nor n17322 n17331 ; n17332
g14897 and n16815_not n17332 ; n17333
g14898 nor n6205 n17333 ; n17334
g14899 and n16808 n17236_not ; n17335
g14900 nor n16643 n17168 ; n17336
g14901 and n16653 n17336_not ; n17337
g14902 and pi0616 n17337_not ; n17338
g14903 and pi0614 n17337_not ; n17339
g14904 and pi0642 n17337_not ; n17340
g14905 nor pi0642 n16807 ; n17341
g14906 and n17236_not n17341 ; n17342
g14907 and n17328 n17342 ; n17343
g14908 nor n17340 n17343 ; n17344
g14909 nor pi0614 n17344 ; n17345
g14910 nor n17339 n17345 ; n17346
g14911 nor pi0616 n17346 ; n17347
g14912 nor n17338 n17347 ; n17348
g14913 and n17323 n17348_not ; n17349
g14914 nor n16804 n17335 ; n17350
g14915 and n17349_not n17350 ; n17351
g14916 and n6205 n17351_not ; n17352
g14917 and pi0223 n17334_not ; n17353
g14918 and n17352_not n17353 ; n17354
g14919 and pi0680 n17336 ; n17355
g14920 and n16653 n17355_not ; n17356
g14921 and n2603 n17356_not ; n17357
g14922 and n16769 n17336_not ; n17358
g14923 nor pi0642 n17358 ; n17359
g14924 nor n17340 n17359 ; n17360
g14925 nor pi0614 n17360 ; n17361
g14926 nor n17339 n17361 ; n17362
g14927 nor pi0616 n17362 ; n17363
g14928 nor n17338 n17363 ; n17364
g14929 and n17323 n17364_not ; n17365
g14930 nor pi0603 n16781 ; n17366
g14931 and pi0603 pi0665_not ; n17367
g14932 and n17144 n17367 ; n17368
g14933 nor n16768 n17368 ; n17369
g14934 and n17366_not n17369 ; n17370
g14935 and n6195 n17370_not ; n17371
g14936 nor n16777 n17371 ; n17372
g14937 and n17365_not n17372 ; n17373
g14938 and n6205 n17373 ; n17374
g14939 and pi0603 n17147 ; n17375
g14940 and pi0603 pi0621_not ; n17376
g14941 and n16754 n17376_not ; n17377
g14942 and n6195 n17377_not ; n17378
g14943 and n17375_not n17378 ; n17379
g14944 and n16702 n17336_not ; n17380
g14945 and n17323 n17380_not ; n17381
g14946 nor n16753 n17379 ; n17382
g14947 and n17381_not n17382 ; n17383
g14948 and n6205_not n17383 ; n17384
g14949 nor n2603 n17384 ; n17385
g14950 and n17374_not n17385 ; n17386
g14951 nor pi0223 n17357 ; n17387
g14952 and n17386_not n17387 ; n17388
g14953 nor n17354 n17388 ; n17389
g14954 nor pi0299 n17389 ; n17390
g14955 and n3448 n17356_not ; n17391
g14956 nor n6242 n17383 ; n17392
g14957 and n6242 n17373_not ; n17393
g14958 nor n17392 n17393 ; n17394
g14959 nor n3448 n17394 ; n17395
g14960 nor pi0215 n17391 ; n17396
g14961 and n17395_not n17396 ; n17397
g14962 and n6242 n17351_not ; n17398
g14963 nor n6242 n17333 ; n17399
g14964 and pi0215 n17399_not ; n17400
g14965 and n17398_not n17400 ; n17401
g14966 nor n17397 n17401 ; n17402
g14967 and pi0299 n17402_not ; n17403
g14968 nor n17390 n17403 ; n17404
g14969 and pi0140_not n17404 ; n17405
g14970 and n17026 n17355 ; n17406
g14971 and n16643_not n17169 ; n17407
g14972 and pi0616 n17407_not ; n17408
g14973 and n17323 n17408_not ; n17409
g14974 and n17166_not n17407 ; n17410
g14975 and pi0603 pi0665 ; n17411
g14976 nor pi0603 n16658 ; n17412
g14977 nor n17411 n17412 ; n17413
g14978 and n17163_not n17413 ; n17414
g14979 and n17166 n17414 ; n17415
g14980 nor pi0616 n17410 ; n17416
g14981 and n17415_not n17416 ; n17417
g14982 and n17409 n17417_not ; n17418
g14983 and n16684 n17371 ; n17419
g14984 nor n17418 n17419 ; n17420
g14985 and n6242 n17420 ; n17421
g14986 and n16687_not n17154 ; n17422
g14987 and pi0616 n17422_not ; n17423
g14988 and pi0665_not n17145 ; n17424
g14989 and pi0603 n17424_not ; n17425
g14990 nor n16687 n16699 ; n17426
g14991 nor pi0603 n17426 ; n17427
g14992 nor n17425 n17427 ; n17428
g14993 and n17166 n17428 ; n17429
g14994 and n17167 n17428_not ; n17430
g14995 and n17422 n17430_not ; n17431
g14996 nor pi0616 n17429 ; n17432
g14997 and n17431_not n17432 ; n17433
g14998 nor n17423 n17433 ; n17434
g14999 nor n16657 n17434 ; n17435
g15000 and n16696 n17425_not ; n17436
g15001 nor n17323 n17436 ; n17437
g15002 nor n17435 n17437 ; n17438
g15003 nor n6242 n17438 ; n17439
g15004 nor n3448 n17421 ; n17440
g15005 and n17439_not n17440 ; n17441
g15006 nor pi0215 n17406 ; n17442
g15007 and n17441_not n17442 ; n17443
g15008 nor n16643 n17196 ; n17444
g15009 nor pi0616 n17444 ; n17445
g15010 and n17409 n17445_not ; n17446
g15011 and n17199 n17413 ; n17447
g15012 nor n17446 n17447 ; n17448
g15013 and n6242 n17448_not ; n17449
g15014 and n17183 n17413 ; n17450
g15015 and pi0616 n17450_not ; n17451
g15016 and pi0614 pi0616_not ; n17452
g15017 and n17450_not n17452 ; n17453
g15018 and n17194_not n17413 ; n17454
g15019 nor pi0642 n17454 ; n17455
g15020 and n17450 n17455_not ; n17456
g15021 and n6191 n17456_not ; n17457
g15022 nor n17453 n17457 ; n17458
g15023 and n17451_not n17458 ; n17459
g15024 nor n16657 n17459 ; n17460
g15025 and n16721_not n17355 ; n17461
g15026 nor n17323 n17461 ; n17462
g15027 nor n17460 n17462 ; n17463
g15028 and n6242_not n17463 ; n17464
g15029 and pi0215 n17449_not ; n17465
g15030 and n17464_not n17465 ; n17466
g15031 nor n17443 n17466 ; n17467
g15032 and pi0299 n17467_not ; n17468
g15033 and n16645 n17168_not ; n17469
g15034 nor n17244 n17469 ; n17470
g15035 and n16653 n17470_not ; n17471
g15036 and n2603 n17471_not ; n17472
g15037 and n6205_not n17438 ; n17473
g15038 and n6205 n17420_not ; n17474
g15039 nor n2603 n17474 ; n17475
g15040 and n17473_not n17475 ; n17476
g15041 and n17269 n17472_not ; n17477
g15042 and n17476_not n17477 ; n17478
g15043 and n6205 n17448 ; n17479
g15044 nor n6205 n17463 ; n17480
g15045 and pi0223 n17479_not ; n17481
g15046 and n17480_not n17481 ; n17482
g15047 nor pi0299 n17482 ; n17483
g15048 and n17478_not n17483 ; n17484
g15049 nor n17468 n17484 ; n17485
g15050 and pi0140 n17485 ; n17486
g15051 and pi0761 n17486_not ; n17487
g15052 and n17405_not n17487 ; n17488
g15053 nor n16644 n17168 ; n17489
g15054 and n16667 n17489 ; n17490
g15055 and n16650_not n17490 ; n17491
g15056 and n2603 n17491 ; n17492
g15057 and n16643 n17376_not ; n17493
g15058 and n16758_not n17493 ; n17494
g15059 and n17323 n17494_not ; n17495
g15060 and n16702 n17168_not ; n17496
g15061 nor pi0680 n17496 ; n17497
g15062 nor n17378 n17495 ; n17498
g15063 and n17497_not n17498 ; n17499
g15064 and n6205_not n17499 ; n17500
g15065 and pi0680_not n17173 ; n17501
g15066 and n16781 n17493 ; n17502
g15067 and n6195 n17502_not ; n17503
g15068 and n16778 n17376_not ; n17504
g15069 and n17167_not n17504 ; n17505
g15070 and n16643 n17172 ; n17506
g15071 and n17323 n17505_not ; n17507
g15072 and n17506_not n17507 ; n17508
g15073 nor n17501 n17503 ; n17509
g15074 and n17508_not n17509 ; n17510
g15075 and n6205 n17510 ; n17511
g15076 nor n17500 n17511 ; n17512
g15077 nor n2603 n17512 ; n17513
g15078 nor pi0223 n17492 ; n17514
g15079 and n17513_not n17514 ; n17515
g15080 and n16644_not n17197 ; n17516
g15081 and n6195 n17376_not ; n17517
g15082 and n16807 n17517 ; n17518
g15083 nor n17516 n17518 ; n17519
g15084 and n6205 n17519_not ; n17520
g15085 nor pi0680 n17185 ; n17521
g15086 nor n16816 n17376 ; n17522
g15087 and n6195 n17522_not ; n17523
g15088 nor n17196 n17324 ; n17524
g15089 and n17323 n17524_not ; n17525
g15090 nor n17521 n17523 ; n17526
g15091 and n17525_not n17526 ; n17527
g15092 and n6205_not n17527 ; n17528
g15093 and pi0223 n17520_not ; n17529
g15094 and n17528_not n17529 ; n17530
g15095 nor n17515 n17530 ; n17531
g15096 nor pi0299 n17531 ; n17532
g15097 and n3448 n17491 ; n17533
g15098 and n6242_not n17499 ; n17534
g15099 and n6242 n17510 ; n17535
g15100 nor n17534 n17535 ; n17536
g15101 nor n3448 n17536 ; n17537
g15102 nor pi0215 n17533 ; n17538
g15103 and n17537_not n17538 ; n17539
g15104 and n6242 n17519_not ; n17540
g15105 and n6242_not n17527 ; n17541
g15106 and pi0215 n17540_not ; n17542
g15107 and n17541_not n17542 ; n17543
g15108 nor n17539 n17543 ; n17544
g15109 and pi0299 n17544_not ; n17545
g15110 nor n17532 n17545 ; n17546
g15111 nor pi0140 n17546 ; n17547
g15112 and n16653 n17493_not ; n17548
g15113 and n17167_not n17548 ; n17549
g15114 and n17323 n17549_not ; n17550
g15115 and n16727 n17236_not ; n17551
g15116 and n17167 n17551_not ; n17552
g15117 and n17550 n17552_not ; n17553
g15118 and pi0680 n16730_not ; n17554
g15119 and n17241 n17554_not ; n17555
g15120 nor n17553 n17555 ; n17556
g15121 and n6205 n17556_not ; n17557
g15122 nor n17240 n17320 ; n17558
g15123 and n16658 n16723_not ; n17559
g15124 and n16727_not n17554 ; n17560
g15125 and n17559 n17560 ; n17561
g15126 and n17558 n17561_not ; n17562
g15127 and n6205_not n17562 ; n17563
g15128 and pi0223 n17563_not ; n17564
g15129 and n17557_not n17564 ; n17565
g15130 and pi0680_not n17250 ; n17566
g15131 nor n17246 n17414 ; n17567
g15132 and n17167 n17567_not ; n17568
g15133 and n17550 n17568_not ; n17569
g15134 and n6195 n16688_not ; n17570
g15135 and n17246_not n17570 ; n17571
g15136 nor n17566 n17571 ; n17572
g15137 and n17569_not n17572 ; n17573
g15138 and n6205 n17573 ; n17574
g15139 nor n17375 n17428 ; n17575
g15140 and n17167 n17575_not ; n17576
g15141 and n16699_not n17168 ; n17577
g15142 nor n17426 n17577 ; n17578
g15143 nor n17167 n17578 ; n17579
g15144 and n17323 n17579_not ; n17580
g15145 and n17576_not n17580 ; n17581
g15146 nor n16696 n17323 ; n17582
g15147 and n17254_not n17582 ; n17583
g15148 nor n17581 n17583 ; n17584
g15149 and n6205_not n17584 ; n17585
g15150 nor n2603 n17574 ; n17586
g15151 and n17585_not n17586 ; n17587
g15152 nor pi0223 n17472 ; n17588
g15153 and n17587_not n17588 ; n17589
g15154 nor pi0299 n17565 ; n17590
g15155 and n17589_not n17590 ; n17591
g15156 and n3448 n17471 ; n17592
g15157 and n6242_not n17584 ; n17593
g15158 and n6242 n17573 ; n17594
g15159 nor n17593 n17594 ; n17595
g15160 nor n3448 n17595 ; n17596
g15161 nor pi0215 n17592 ; n17597
g15162 and n17596_not n17597 ; n17598
g15163 nor n6242 n17562 ; n17599
g15164 and n6242 n17556 ; n17600
g15165 and pi0215 n17599_not ; n17601
g15166 and n17600_not n17601 ; n17602
g15167 nor n17598 n17602 ; n17603
g15168 and pi0299 n17603_not ; n17604
g15169 nor n17591 n17604 ; n17605
g15170 and pi0140 n17605 ; n17606
g15171 nor pi0761 n17547 ; n17607
g15172 and n17606_not n17607 ; n17608
g15173 nor n17488 n17608 ; n17609
g15174 and pi0039 n17609_not ; n17610
g15175 and pi0680 n17233 ; n17611
g15176 nor n16948 n17611 ; n17612
g15177 nor pi0140 n17612 ; n17613
g15178 and pi0603 n17128_not ; n17614
g15179 nor pi0603 n16918 ; n17615
g15180 nor n17411 n17614 ; n17616
g15181 and n17615_not n17616 ; n17617
g15182 and pi0680 n17617 ; n17618
g15183 nor pi0299 n17618 ; n17619
g15184 nor pi0603 n16923 ; n17620
g15185 nor n17123 n17411 ; n17621
g15186 and n17620_not n17621 ; n17622
g15187 and pi0680 n17622 ; n17623
g15188 and pi0299 n17623_not ; n17624
g15189 nor n17619 n17624 ; n17625
g15190 and pi0140 n17625_not ; n17626
g15191 and pi0761 n17613_not ; n17627
g15192 and n17626_not n17627 ; n17628
g15193 and n16948 n17139 ; n17629
g15194 and pi0140_not n17629 ; n17630
g15195 nor n16926 n17233 ; n17631
g15196 and pi0140 n17631 ; n17632
g15197 nor pi0761 n17632 ; n17633
g15198 and n17630_not n17633 ; n17634
g15199 nor pi0039 n17634 ; n17635
g15200 and n17628_not n17635 ; n17636
g15201 nor pi0038 n17636 ; n17637
g15202 and n17610_not n17637 ; n17638
g15203 and pi0140 n17470_not ; n17639
g15204 and n2521 n17639 ; n17640
g15205 nor pi0140 n17490 ; n17641
g15206 nor pi0761 n17640 ; n17642
g15207 and n17641_not n17642 ; n17643
g15208 nor pi0140 n16667 ; n17644
g15209 and n16667 n17355 ; n17645
g15210 and pi0761 n17644_not ; n17646
g15211 and n17645_not n17646 ; n17647
g15212 nor n17643 n17647 ; n17648
g15213 nor pi0039 n17648 ; n17649
g15214 and pi0038 n16751_not ; n17650
g15215 and n17649_not n17650 ; n17651
g15216 nor n17638 n17651 ; n17652
g15217 nor pi0738 n17652 ; n17653
g15218 and n2571 n17319_not ; n17654
g15219 and n17653_not n17654 ; n17655
g15220 nor n16640 n17655 ; n17656
g15221 and pi0625_not n17656 ; n17657
g15222 and pi0625 n17286 ; n17658
g15223 nor pi1153 n17658 ; n17659
g15224 and n17657_not n17659 ; n17660
g15225 nor pi0608 n17064 ; n17661
g15226 and n17660_not n17661 ; n17662
g15227 and pi0625_not n17286 ; n17663
g15228 and pi0625 n17656 ; n17664
g15229 and pi1153 n17663_not ; n17665
g15230 and n17664_not n17665 ; n17666
g15231 and pi0608 n17068_not ; n17667
g15232 and n17666_not n17667 ; n17668
g15233 nor n17662 n17668 ; n17669
g15234 and pi0778 n17669_not ; n17670
g15235 and pi0778_not n17656 ; n17671
g15236 nor n17670 n17671 ; n17672
g15237 nor pi0609 n17672 ; n17673
g15238 and pi0609 n17071 ; n17674
g15239 nor pi1155 n17674 ; n17675
g15240 and n17673_not n17675 ; n17676
g15241 nor pi0660 n17295 ; n17677
g15242 and n17676_not n17677 ; n17678
g15243 and pi0609_not n17071 ; n17679
g15244 and pi0609 n17672_not ; n17680
g15245 and pi1155 n17679_not ; n17681
g15246 and n17680_not n17681 ; n17682
g15247 and pi0660 n17300_not ; n17683
g15248 and n17682_not n17683 ; n17684
g15249 nor n17678 n17684 ; n17685
g15250 and pi0785 n17685_not ; n17686
g15251 nor pi0785 n17672 ; n17687
g15252 nor n17686 n17687 ; n17688
g15253 nor pi0618 n17688 ; n17689
g15254 and pi0618 n17078 ; n17690
g15255 nor pi1154 n17690 ; n17691
g15256 and n17689_not n17691 ; n17692
g15257 nor pi0627 n17308 ; n17693
g15258 and n17692_not n17693 ; n17694
g15259 and pi0618_not n17078 ; n17695
g15260 and pi0618 n17688_not ; n17696
g15261 and pi1154 n17695_not ; n17697
g15262 and n17696_not n17697 ; n17698
g15263 and pi0627 n17312_not ; n17699
g15264 and n17698_not n17699 ; n17700
g15265 nor n17694 n17700 ; n17701
g15266 and pi0781 n17701_not ; n17702
g15267 nor pi0781 n17688 ; n17703
g15268 nor n17702 n17703 ; n17704
g15269 nor pi0619 n17704 ; n17705
g15270 and pi0619 n17081_not ; n17706
g15271 nor pi1159 n17706 ; n17707
g15272 and n17705_not n17707 ; n17708
g15273 nor pi0648 n17318 ; n17709
g15274 and n17708_not n17709 ; n17710
g15275 and pi0619_not n17315 ; n17711
g15276 and pi0619 n17060 ; n17712
g15277 nor pi1159 n17712 ; n17713
g15278 and n17711_not n17713 ; n17714
g15279 and pi0619 n17704_not ; n17715
g15280 nor pi0619 n17081 ; n17716
g15281 and pi1159 n17716_not ; n17717
g15282 and n17715_not n17717 ; n17718
g15283 and pi0648 n17714_not ; n17719
g15284 and n17718_not n17719 ; n17720
g15285 nor n17710 n17720 ; n17721
g15286 and pi0789 n17721_not ; n17722
g15287 nor pi0789 n17704 ; n17723
g15288 nor n17722 n17723 ; n17724
g15289 and pi0788_not n17724 ; n17725
g15290 and pi0626_not n17724 ; n17726
g15291 and pi0626 n17084_not ; n17727
g15292 nor pi0641 n17727 ; n17728
g15293 and n17726_not n17728 ; n17729
g15294 nor pi0641 pi1158 ; n17730
g15295 nor pi0789 n17315 ; n17731
g15296 nor n17318 n17714 ; n17732
g15297 and pi0789 n17732_not ; n17733
g15298 nor n17731 n17733 ; n17734
g15299 and pi0626_not n17734 ; n17735
g15300 and pi0626 n17060 ; n17736
g15301 nor pi1158 n17736 ; n17737
g15302 and n17735_not n17737 ; n17738
g15303 nor n17730 n17738 ; n17739
g15304 nor n17729 n17739 ; n17740
g15305 and pi0626 n17724 ; n17741
g15306 nor pi0626 n17084 ; n17742
g15307 and pi0641 n17742_not ; n17743
g15308 and n17741_not n17743 ; n17744
g15309 and pi0641 pi1158 ; n17745
g15310 and pi0626_not n17060 ; n17746
g15311 and pi0626 n17734 ; n17747
g15312 and pi1158 n17746_not ; n17748
g15313 and n17747_not n17748 ; n17749
g15314 nor n17745 n17749 ; n17750
g15315 nor n17744 n17750 ; n17751
g15316 nor n17740 n17751 ; n17752
g15317 and pi0788 n17752_not ; n17753
g15318 nor n17725 n17753 ; n17754
g15319 and pi0628_not n17754 ; n17755
g15320 nor n17738 n17749 ; n17756
g15321 and pi0788 n17756_not ; n17757
g15322 nor pi0788 n17734 ; n17758
g15323 nor n17757 n17758 ; n17759
g15324 and pi0628 n17759 ; n17760
g15325 nor pi1156 n17760 ; n17761
g15326 and n17755_not n17761 ; n17762
g15327 nor pi0629 n17092 ; n17763
g15328 and n17762_not n17763 ; n17764
g15329 and pi0628 n17754 ; n17765
g15330 and pi0628_not n17759 ; n17766
g15331 and pi1156 n17766_not ; n17767
g15332 and n17765_not n17767 ; n17768
g15333 and pi0629 n17096_not ; n17769
g15334 and n17768_not n17769 ; n17770
g15335 nor n17764 n17770 ; n17771
g15336 and pi0792 n17771_not ; n17772
g15337 and pi0792_not n17754 ; n17773
g15338 nor n17772 n17773 ; n17774
g15339 nor pi0647 n17774 ; n17775
g15340 and pi0629_not pi1156 ; n17776
g15341 and pi0629 pi1156_not ; n17777
g15342 nor n17776 n17777 ; n17778
g15343 and pi0792 n17778_not ; n17779
g15344 and n17759 n17779_not ; n17780
g15345 and n17060 n17779 ; n17781
g15346 nor n17780 n17781 ; n17782
g15347 and pi0647 n17782_not ; n17783
g15348 nor pi1157 n17783 ; n17784
g15349 and n17775_not n17784 ; n17785
g15350 nor pi0630 n17104 ; n17786
g15351 and n17785_not n17786 ; n17787
g15352 and pi0647 n17774_not ; n17788
g15353 nor pi0647 n17782 ; n17789
g15354 and pi1157 n17789_not ; n17790
g15355 and n17788_not n17790 ; n17791
g15356 and pi0630 n17108_not ; n17792
g15357 and n17791_not n17792 ; n17793
g15358 nor n17787 n17793 ; n17794
g15359 and pi0787 n17794_not ; n17795
g15360 nor pi0787 n17774 ; n17796
g15361 nor n17795 n17796 ; n17797
g15362 and pi0644 n17797_not ; n17798
g15363 and pi0715 n17112_not ; n17799
g15364 and n17798_not n17799 ; n17800
g15365 and pi0630_not pi1157 ; n17801
g15366 and pi0630 pi1157_not ; n17802
g15367 nor n17801 n17802 ; n17803
g15368 and pi0787 n17803_not ; n17804
g15369 and n17782 n17804_not ; n17805
g15370 and n17060_not n17804 ; n17806
g15371 nor n17805 n17806 ; n17807
g15372 and pi0644 n17807 ; n17808
g15373 and pi0644_not n17060 ; n17809
g15374 nor pi0715 n17809 ; n17810
g15375 and n17808_not n17810 ; n17811
g15376 and pi1160 n17811_not ; n17812
g15377 and n17800_not n17812 ; n17813
g15378 nor pi0644 n17797 ; n17814
g15379 and pi0644 n17111 ; n17815
g15380 nor pi0715 n17815 ; n17816
g15381 and n17814_not n17816 ; n17817
g15382 and pi0644_not n17807 ; n17818
g15383 and pi0644 n17060 ; n17819
g15384 and pi0715 n17819_not ; n17820
g15385 and n17818_not n17820 ; n17821
g15386 nor pi1160 n17821 ; n17822
g15387 and n17817_not n17822 ; n17823
g15388 and pi0790 n17813_not ; n17824
g15389 and n17823_not n17824 ; n17825
g15390 and pi0790_not n17797 ; n17826
g15391 nor po1038 n17826 ; n17827
g15392 and n17825_not n17827 ; n17828
g15393 and pi0140_not po1038 ; n17829
g15394 nor pi0832 n17829 ; n17830
g15395 and n17828_not n17830 ; n17831
g15396 nor pi0140 n2926 ; n17832
g15397 and pi0647_not n17832 ; n17833
g15398 and pi0738_not n16645 ; n17834
g15399 nor n17832 n17834 ; n17835
g15400 and pi0778_not n17835 ; n17836
g15401 and pi0625_not n17834 ; n17837
g15402 nor n17835 n17837 ; n17838
g15403 and pi1153 n17838_not ; n17839
g15404 nor pi1153 n17832 ; n17840
g15405 and n17837_not n17840 ; n17841
g15406 nor n17839 n17841 ; n17842
g15407 and pi0778 n17842_not ; n17843
g15408 nor n17836 n17843 ; n17844
g15409 and n2926 n17075 ; n17845
g15410 and n17844 n17845_not ; n17846
g15411 and n2926 n16639 ; n17847
g15412 and n17846 n17847_not ; n17848
g15413 and n2926 n16635 ; n17849
g15414 and n17848 n17849_not ; n17850
g15415 and n2926 n16631 ; n17851
g15416 and n17850 n17851_not ; n17852
g15417 and pi0628_not pi1156 ; n17853
g15418 and pi0628 pi1156_not ; n17854
g15419 nor n17853 n17854 ; n17855
g15420 and pi0792 n17855_not ; n17856
g15421 and n2926 n17856 ; n17857
g15422 and n17852 n17857_not ; n17858
g15423 and pi0647 n17858 ; n17859
g15424 and pi1157 n17833_not ; n17860
g15425 and n17859_not n17860 ; n17861
g15426 and pi0628_not n2926 ; n17862
g15427 and n17852 n17862_not ; n17863
g15428 and pi1156 n17863_not ; n17864
g15429 and pi0626_not pi1158 ; n17865
g15430 and pi0626 pi1158_not ; n17866
g15431 nor n17865 n17866 ; n17867
g15432 and pi0626_not pi0641 ; n17868
g15433 and pi0626 pi0641_not ; n17869
g15434 nor n17868 n17869 ; n17870
g15435 nor n17867 n17870 ; n17871
g15436 and n17850 n17871 ; n17872
g15437 and pi0626_not n17832 ; n17873
g15438 and n2926 n17117 ; n17874
g15439 and pi0761_not n17244 ; n17875
g15440 nor n17832 n17875 ; n17876
g15441 nor n17874 n17876 ; n17877
g15442 nor pi0785 n17877 ; n17878
g15443 and n2926 n17291_not ; n17879
g15444 nor n17876 n17879 ; n17880
g15445 and pi1155 n17880_not ; n17881
g15446 and pi0609 n2926 ; n17882
g15447 and n17877 n17882_not ; n17883
g15448 nor pi1155 n17883 ; n17884
g15449 nor n17881 n17884 ; n17885
g15450 and pi0785 n17885_not ; n17886
g15451 nor n17878 n17886 ; n17887
g15452 nor pi0781 n17887 ; n17888
g15453 and pi0618_not n2926 ; n17889
g15454 and n17887 n17889_not ; n17890
g15455 and pi1154 n17890_not ; n17891
g15456 and pi0618 n2926 ; n17892
g15457 and n17887 n17892_not ; n17893
g15458 nor pi1154 n17893 ; n17894
g15459 nor n17891 n17894 ; n17895
g15460 and pi0781 n17895_not ; n17896
g15461 nor n17888 n17896 ; n17897
g15462 nor pi0789 n17897 ; n17898
g15463 and pi0619_not n17832 ; n17899
g15464 and pi0619 n17897 ; n17900
g15465 and pi1159 n17899_not ; n17901
g15466 and n17900_not n17901 ; n17902
g15467 and pi0619_not n17897 ; n17903
g15468 and pi0619 n17832 ; n17904
g15469 nor pi1159 n17904 ; n17905
g15470 and n17903_not n17905 ; n17906
g15471 nor n17902 n17906 ; n17907
g15472 and pi0789 n17907_not ; n17908
g15473 nor n17898 n17908 ; n17909
g15474 and pi0626 n17909 ; n17910
g15475 and pi1158 n17873_not ; n17911
g15476 and n17910_not n17911 ; n17912
g15477 and pi0626_not n17909 ; n17913
g15478 and pi0626 n17832 ; n17914
g15479 nor pi1158 n17914 ; n17915
g15480 and n17913_not n17915 ; n17916
g15481 nor n17912 n17916 ; n17917
g15482 and n16630_not n17917 ; n17918
g15483 nor n17872 n17918 ; n17919
g15484 and pi0788 n17919_not ; n17920
g15485 and pi0618 n17846 ; n17921
g15486 and pi0609 n17844 ; n17922
g15487 nor n17168 n17835 ; n17923
g15488 and pi0625 n17923 ; n17924
g15489 and n17876 n17923_not ; n17925
g15490 nor n17924 n17925 ; n17926
g15491 and n17840 n17926_not ; n17927
g15492 nor pi0608 n17839 ; n17928
g15493 and n17927_not n17928 ; n17929
g15494 and pi1153 n17876 ; n17930
g15495 and n17924_not n17930 ; n17931
g15496 and pi0608 n17841_not ; n17932
g15497 and n17931_not n17932 ; n17933
g15498 nor n17929 n17933 ; n17934
g15499 and pi0778 n17934_not ; n17935
g15500 nor pi0778 n17925 ; n17936
g15501 nor n17935 n17936 ; n17937
g15502 nor pi0609 n17937 ; n17938
g15503 nor pi1155 n17922 ; n17939
g15504 and n17938_not n17939 ; n17940
g15505 nor pi0660 n17881 ; n17941
g15506 and n17940_not n17941 ; n17942
g15507 and pi0609_not n17844 ; n17943
g15508 and pi0609 n17937_not ; n17944
g15509 and pi1155 n17943_not ; n17945
g15510 and n17944_not n17945 ; n17946
g15511 and pi0660 n17884_not ; n17947
g15512 and n17946_not n17947 ; n17948
g15513 nor n17942 n17948 ; n17949
g15514 and pi0785 n17949_not ; n17950
g15515 nor pi0785 n17937 ; n17951
g15516 nor n17950 n17951 ; n17952
g15517 nor pi0618 n17952 ; n17953
g15518 nor pi1154 n17921 ; n17954
g15519 and n17953_not n17954 ; n17955
g15520 nor pi0627 n17891 ; n17956
g15521 and n17955_not n17956 ; n17957
g15522 and pi0618_not n17846 ; n17958
g15523 and pi0618 n17952_not ; n17959
g15524 and pi1154 n17958_not ; n17960
g15525 and n17959_not n17960 ; n17961
g15526 and pi0627 n17894_not ; n17962
g15527 and n17961_not n17962 ; n17963
g15528 nor n17957 n17963 ; n17964
g15529 and pi0781 n17964_not ; n17965
g15530 nor pi0781 n17952 ; n17966
g15531 nor n17965 n17966 ; n17967
g15532 and pi0789_not n17967 ; n17968
g15533 and pi0788 n17867_not ; n17969
g15534 nor n16631 n17969 ; n17970
g15535 nor pi0619 n17967 ; n17971
g15536 and pi0619 n17848 ; n17972
g15537 nor pi1159 n17972 ; n17973
g15538 and n17971_not n17973 ; n17974
g15539 nor pi0648 n17902 ; n17975
g15540 and n17974_not n17975 ; n17976
g15541 and pi0619_not n17848 ; n17977
g15542 and pi0619 n17967_not ; n17978
g15543 and pi1159 n17977_not ; n17979
g15544 and n17978_not n17979 ; n17980
g15545 and pi0648 n17906_not ; n17981
g15546 and n17980_not n17981 ; n17982
g15547 and pi0789 n17976_not ; n17983
g15548 and n17982_not n17983 ; n17984
g15549 and n17968_not n17970 ; n17985
g15550 and n17984_not n17985 ; n17986
g15551 nor n17920 n17986 ; n17987
g15552 nor pi0628 n17987 ; n17988
g15553 nor pi0788 n17909 ; n17989
g15554 and pi0788 n17917_not ; n17990
g15555 nor n17989 n17990 ; n17991
g15556 and pi0628 n17991 ; n17992
g15557 nor pi1156 n17992 ; n17993
g15558 and n17988_not n17993 ; n17994
g15559 nor pi0629 n17864 ; n17995
g15560 and n17994_not n17995 ; n17996
g15561 and pi0628 n2926 ; n17997
g15562 and n17852 n17997_not ; n17998
g15563 nor pi1156 n17998 ; n17999
g15564 and pi0628_not n17991 ; n18000
g15565 and pi0628 n17987_not ; n18001
g15566 and pi1156 n18000_not ; n18002
g15567 and n18001_not n18002 ; n18003
g15568 and pi0629 n17999_not ; n18004
g15569 and n18003_not n18004 ; n18005
g15570 nor n17996 n18005 ; n18006
g15571 and pi0792 n18006_not ; n18007
g15572 nor pi0792 n17987 ; n18008
g15573 nor n18007 n18008 ; n18009
g15574 nor pi0647 n18009 ; n18010
g15575 and n17779_not n17991 ; n18011
g15576 and n17779 n17832 ; n18012
g15577 nor n18011 n18012 ; n18013
g15578 and pi0647 n18013_not ; n18014
g15579 nor pi1157 n18014 ; n18015
g15580 and n18010_not n18015 ; n18016
g15581 nor pi0630 n17861 ; n18017
g15582 and n18016_not n18017 ; n18018
g15583 and pi0647_not n17858 ; n18019
g15584 and pi0647 n17832 ; n18020
g15585 nor pi1157 n18020 ; n18021
g15586 and n18019_not n18021 ; n18022
g15587 and pi0647 n18009_not ; n18023
g15588 nor pi0647 n18013 ; n18024
g15589 and pi1157 n18024_not ; n18025
g15590 and n18023_not n18025 ; n18026
g15591 and pi0630 n18022_not ; n18027
g15592 and n18026_not n18027 ; n18028
g15593 nor n18018 n18028 ; n18029
g15594 and pi0787 n18029_not ; n18030
g15595 nor pi0787 n18009 ; n18031
g15596 nor n18030 n18031 ; n18032
g15597 nor pi0790 n18032 ; n18033
g15598 nor pi0787 n17858 ; n18034
g15599 nor n17861 n18022 ; n18035
g15600 and pi0787 n18035_not ; n18036
g15601 nor n18034 n18036 ; n18037
g15602 and pi0644_not n18037 ; n18038
g15603 and pi0644 n18032_not ; n18039
g15604 and pi0715 n18038_not ; n18040
g15605 and n18039_not n18040 ; n18041
g15606 and n17804 n17832_not ; n18042
g15607 and n17804_not n18013 ; n18043
g15608 nor n18042 n18043 ; n18044
g15609 and pi0644 n18044 ; n18045
g15610 and pi0644_not n17832 ; n18046
g15611 nor pi0715 n18046 ; n18047
g15612 and n18045_not n18047 ; n18048
g15613 and pi1160 n18048_not ; n18049
g15614 and n18041_not n18049 ; n18050
g15615 and pi0644_not n18044 ; n18051
g15616 and pi0644 n17832 ; n18052
g15617 and pi0715 n18052_not ; n18053
g15618 and n18051_not n18053 ; n18054
g15619 and pi0644 n18037 ; n18055
g15620 nor pi0644 n18032 ; n18056
g15621 nor pi0715 n18055 ; n18057
g15622 and n18056_not n18057 ; n18058
g15623 nor pi1160 n18054 ; n18059
g15624 and n18058_not n18059 ; n18060
g15625 nor n18050 n18060 ; n18061
g15626 and pi0790 n18061_not ; n18062
g15627 and pi0832 n18033_not ; n18063
g15628 and n18062_not n18063 ; n18064
g15629 nor n17831 n18064 ; po0297
g15630 nor pi0141 n17059 ; n18066
g15631 and n16635 n18066_not ; n18067
g15632 and pi0141 n2571_not ; n18068
g15633 nor pi0141 n16641 ; n18069
g15634 and n16647 n18069_not ; n18070
g15635 and pi0039_not n16948 ; n18071
g15636 nor n16841 n18071 ; n18072
g15637 and pi0141_not n18072 ; n18073
g15638 and pi0039 n16749_not ; n18074
g15639 and pi0039_not n16926 ; n18075
g15640 nor n18074 n18075 ; n18076
g15641 and pi0141 n18076_not ; n18077
g15642 nor pi0038 n18077 ; n18078
g15643 and n18073_not n18078 ; n18079
g15644 and pi0706 n18070_not ; n18080
g15645 and n18079_not n18080 ; n18081
g15646 nor pi0141 pi0706 ; n18082
g15647 and n17052_not n18082 ; n18083
g15648 and n2571 n18083_not ; n18084
g15649 and n18081_not n18084 ; n18085
g15650 nor n18068 n18085 ; n18086
g15651 nor pi0778 n18086 ; n18087
g15652 and pi0625_not n18066 ; n18088
g15653 and pi0625 n18086 ; n18089
g15654 and pi1153 n18088_not ; n18090
g15655 and n18089_not n18090 ; n18091
g15656 and pi0625_not n18086 ; n18092
g15657 and pi0625 n18066 ; n18093
g15658 nor pi1153 n18093 ; n18094
g15659 and n18092_not n18094 ; n18095
g15660 nor n18091 n18095 ; n18096
g15661 and pi0778 n18096_not ; n18097
g15662 nor n18087 n18097 ; n18098
g15663 nor n17075 n18098 ; n18099
g15664 and n17075 n18066_not ; n18100
g15665 nor n18099 n18100 ; n18101
g15666 and n16639_not n18101 ; n18102
g15667 and n16639 n18066 ; n18103
g15668 nor n18102 n18103 ; n18104
g15669 and n16635_not n18104 ; n18105
g15670 nor n18067 n18105 ; n18106
g15671 and n16631_not n18106 ; n18107
g15672 and n16631 n18066 ; n18108
g15673 nor n18107 n18108 ; n18109
g15674 and pi0792_not n18109 ; n18110
g15675 and pi0628_not n18066 ; n18111
g15676 and pi0628 n18109_not ; n18112
g15677 and pi1156 n18111_not ; n18113
g15678 and n18112_not n18113 ; n18114
g15679 and pi0628 n18066 ; n18115
g15680 nor pi0628 n18109 ; n18116
g15681 nor pi1156 n18115 ; n18117
g15682 and n18116_not n18117 ; n18118
g15683 nor n18114 n18118 ; n18119
g15684 and pi0792 n18119_not ; n18120
g15685 nor n18110 n18120 ; n18121
g15686 nor pi0787 n18121 ; n18122
g15687 and pi0647_not n18066 ; n18123
g15688 and pi0647 n18121 ; n18124
g15689 and pi1157 n18123_not ; n18125
g15690 and n18124_not n18125 ; n18126
g15691 and pi0647_not n18121 ; n18127
g15692 and pi0647 n18066 ; n18128
g15693 nor pi1157 n18128 ; n18129
g15694 and n18127_not n18129 ; n18130
g15695 nor n18126 n18130 ; n18131
g15696 and pi0787 n18131_not ; n18132
g15697 nor n18122 n18132 ; n18133
g15698 and pi0644_not n18133 ; n18134
g15699 and pi0618_not n18066 ; n18135
g15700 and pi0749 n17280 ; n18136
g15701 nor n18069 n18136 ; n18137
g15702 and pi0038 n18137_not ; n18138
g15703 and pi0749_not n17046 ; n18139
g15704 and pi0141 n17273 ; n18140
g15705 nor n18139 n18140 ; n18141
g15706 and pi0039 n18141_not ; n18142
g15707 and pi0141_not n17221 ; n18143
g15708 and pi0141 n17234 ; n18144
g15709 and pi0749 n18144_not ; n18145
g15710 and n18143_not n18145 ; n18146
g15711 and pi0039_not n16958 ; n18147
g15712 nor pi0141 pi0749 ; n18148
g15713 and n18147_not n18148 ; n18149
g15714 nor n18146 n18149 ; n18150
g15715 nor pi0038 n18150 ; n18151
g15716 and n18142_not n18151 ; n18152
g15717 nor n18138 n18152 ; n18153
g15718 and n2571 n18153 ; n18154
g15719 nor n18068 n18154 ; n18155
g15720 nor n17117 n18155 ; n18156
g15721 and n17117 n18066_not ; n18157
g15722 nor n18156 n18157 ; n18158
g15723 nor pi0785 n18158 ; n18159
g15724 nor n17291 n18066 ; n18160
g15725 and pi0609 n18156 ; n18161
g15726 nor n18160 n18161 ; n18162
g15727 and pi1155 n18162_not ; n18163
g15728 nor n17296 n18066 ; n18164
g15729 and pi0609_not n18156 ; n18165
g15730 nor n18164 n18165 ; n18166
g15731 nor pi1155 n18166 ; n18167
g15732 nor n18163 n18167 ; n18168
g15733 and pi0785 n18168_not ; n18169
g15734 nor n18159 n18169 ; n18170
g15735 and pi0618 n18170 ; n18171
g15736 and pi1154 n18135_not ; n18172
g15737 and n18171_not n18172 ; n18173
g15738 nor pi0706 n18153 ; n18174
g15739 and pi0039_not n17645 ; n18175
g15740 and pi0038 n18175_not ; n18176
g15741 and n18137 n18176 ; n18177
g15742 nor pi0141 n17629 ; n18178
g15743 and pi0141 n17631_not ; n18179
g15744 and pi0749 n18179_not ; n18180
g15745 and n18178_not n18180 ; n18181
g15746 and pi0141_not n17612 ; n18182
g15747 and pi0141 n17625 ; n18183
g15748 nor pi0749 n18182 ; n18184
g15749 and n18183_not n18184 ; n18185
g15750 nor pi0039 n18181 ; n18186
g15751 and n18185_not n18186 ; n18187
g15752 and pi0141 n17605 ; n18188
g15753 nor pi0141 n17546 ; n18189
g15754 and pi0749 n18189_not ; n18190
g15755 and n18188_not n18190 ; n18191
g15756 and pi0141_not n17404 ; n18192
g15757 and pi0141 n17485 ; n18193
g15758 nor pi0749 n18193 ; n18194
g15759 and n18192_not n18194 ; n18195
g15760 and pi0039 n18191_not ; n18196
g15761 and n18195_not n18196 ; n18197
g15762 nor pi0038 n18187 ; n18198
g15763 and n18197_not n18198 ; n18199
g15764 and pi0706 n18177_not ; n18200
g15765 and n18199_not n18200 ; n18201
g15766 and n2571 n18174_not ; n18202
g15767 and n18201_not n18202 ; n18203
g15768 nor n18068 n18203 ; n18204
g15769 and pi0625_not n18204 ; n18205
g15770 and pi0625 n18155 ; n18206
g15771 nor pi1153 n18206 ; n18207
g15772 and n18205_not n18207 ; n18208
g15773 nor pi0608 n18091 ; n18209
g15774 and n18208_not n18209 ; n18210
g15775 and pi0625_not n18155 ; n18211
g15776 and pi0625 n18204 ; n18212
g15777 and pi1153 n18211_not ; n18213
g15778 and n18212_not n18213 ; n18214
g15779 and pi0608 n18095_not ; n18215
g15780 and n18214_not n18215 ; n18216
g15781 nor n18210 n18216 ; n18217
g15782 and pi0778 n18217_not ; n18218
g15783 and pi0778_not n18204 ; n18219
g15784 nor n18218 n18219 ; n18220
g15785 nor pi0609 n18220 ; n18221
g15786 and pi0609 n18098 ; n18222
g15787 nor pi1155 n18222 ; n18223
g15788 and n18221_not n18223 ; n18224
g15789 nor pi0660 n18163 ; n18225
g15790 and n18224_not n18225 ; n18226
g15791 and pi0609_not n18098 ; n18227
g15792 and pi0609 n18220_not ; n18228
g15793 and pi1155 n18227_not ; n18229
g15794 and n18228_not n18229 ; n18230
g15795 and pi0660 n18167_not ; n18231
g15796 and n18230_not n18231 ; n18232
g15797 nor n18226 n18232 ; n18233
g15798 and pi0785 n18233_not ; n18234
g15799 nor pi0785 n18220 ; n18235
g15800 nor n18234 n18235 ; n18236
g15801 nor pi0618 n18236 ; n18237
g15802 and pi0618 n18101 ; n18238
g15803 nor pi1154 n18238 ; n18239
g15804 and n18237_not n18239 ; n18240
g15805 nor pi0627 n18173 ; n18241
g15806 and n18240_not n18241 ; n18242
g15807 and pi0618_not n18170 ; n18243
g15808 and pi0618 n18066 ; n18244
g15809 nor pi1154 n18244 ; n18245
g15810 and n18243_not n18245 ; n18246
g15811 and pi0618_not n18101 ; n18247
g15812 and pi0618 n18236_not ; n18248
g15813 and pi1154 n18247_not ; n18249
g15814 and n18248_not n18249 ; n18250
g15815 and pi0627 n18246_not ; n18251
g15816 and n18250_not n18251 ; n18252
g15817 nor n18242 n18252 ; n18253
g15818 and pi0781 n18253_not ; n18254
g15819 nor pi0781 n18236 ; n18255
g15820 nor n18254 n18255 ; n18256
g15821 nor pi0619 n18256 ; n18257
g15822 and pi0619 n18104_not ; n18258
g15823 nor pi1159 n18258 ; n18259
g15824 and n18257_not n18259 ; n18260
g15825 and pi0619_not n18066 ; n18261
g15826 nor pi0781 n18170 ; n18262
g15827 nor n18173 n18246 ; n18263
g15828 and pi0781 n18263_not ; n18264
g15829 nor n18262 n18264 ; n18265
g15830 and pi0619 n18265 ; n18266
g15831 and pi1159 n18261_not ; n18267
g15832 and n18266_not n18267 ; n18268
g15833 nor pi0648 n18268 ; n18269
g15834 and n18260_not n18269 ; n18270
g15835 and pi0619 n18256_not ; n18271
g15836 nor pi0619 n18104 ; n18272
g15837 and pi1159 n18272_not ; n18273
g15838 and n18271_not n18273 ; n18274
g15839 and pi0619_not n18265 ; n18275
g15840 and pi0619 n18066 ; n18276
g15841 nor pi1159 n18276 ; n18277
g15842 and n18275_not n18277 ; n18278
g15843 and pi0648 n18278_not ; n18279
g15844 and n18274_not n18279 ; n18280
g15845 nor n18270 n18280 ; n18281
g15846 and pi0789 n18281_not ; n18282
g15847 nor pi0789 n18256 ; n18283
g15848 nor n18282 n18283 ; n18284
g15849 and pi0788_not n18284 ; n18285
g15850 and pi0626_not n18284 ; n18286
g15851 and pi0626 n18106_not ; n18287
g15852 nor pi0641 n18287 ; n18288
g15853 and n18286_not n18288 ; n18289
g15854 nor pi0789 n18265 ; n18290
g15855 nor n18268 n18278 ; n18291
g15856 and pi0789 n18291_not ; n18292
g15857 nor n18290 n18292 ; n18293
g15858 and pi0626_not n18293 ; n18294
g15859 and pi0626 n18066 ; n18295
g15860 nor pi1158 n18295 ; n18296
g15861 and n18294_not n18296 ; n18297
g15862 nor n17730 n18297 ; n18298
g15863 nor n18289 n18298 ; n18299
g15864 and pi0626 n18284 ; n18300
g15865 nor pi0626 n18106 ; n18301
g15866 and pi0641 n18301_not ; n18302
g15867 and n18300_not n18302 ; n18303
g15868 and pi0626_not n18066 ; n18304
g15869 and pi0626 n18293 ; n18305
g15870 and pi1158 n18304_not ; n18306
g15871 and n18305_not n18306 ; n18307
g15872 nor n17745 n18307 ; n18308
g15873 nor n18303 n18308 ; n18309
g15874 nor n18299 n18309 ; n18310
g15875 and pi0788 n18310_not ; n18311
g15876 nor n18285 n18311 ; n18312
g15877 and pi0628_not n18312 ; n18313
g15878 nor n18297 n18307 ; n18314
g15879 and pi0788 n18314_not ; n18315
g15880 nor pi0788 n18293 ; n18316
g15881 nor n18315 n18316 ; n18317
g15882 and pi0628 n18317 ; n18318
g15883 nor pi1156 n18318 ; n18319
g15884 and n18313_not n18319 ; n18320
g15885 nor pi0629 n18114 ; n18321
g15886 and n18320_not n18321 ; n18322
g15887 and pi0628 n18312 ; n18323
g15888 and pi0628_not n18317 ; n18324
g15889 and pi1156 n18324_not ; n18325
g15890 and n18323_not n18325 ; n18326
g15891 and pi0629 n18118_not ; n18327
g15892 and n18326_not n18327 ; n18328
g15893 nor n18322 n18328 ; n18329
g15894 and pi0792 n18329_not ; n18330
g15895 and pi0792_not n18312 ; n18331
g15896 nor n18330 n18331 ; n18332
g15897 nor pi0647 n18332 ; n18333
g15898 and n17779_not n18317 ; n18334
g15899 and n17779 n18066 ; n18335
g15900 nor n18334 n18335 ; n18336
g15901 and pi0647 n18336_not ; n18337
g15902 nor pi1157 n18337 ; n18338
g15903 and n18333_not n18338 ; n18339
g15904 nor pi0630 n18126 ; n18340
g15905 and n18339_not n18340 ; n18341
g15906 and pi0647 n18332_not ; n18342
g15907 nor pi0647 n18336 ; n18343
g15908 and pi1157 n18343_not ; n18344
g15909 and n18342_not n18344 ; n18345
g15910 and pi0630 n18130_not ; n18346
g15911 and n18345_not n18346 ; n18347
g15912 nor n18341 n18347 ; n18348
g15913 and pi0787 n18348_not ; n18349
g15914 nor pi0787 n18332 ; n18350
g15915 nor n18349 n18350 ; n18351
g15916 and pi0644 n18351_not ; n18352
g15917 and pi0715 n18134_not ; n18353
g15918 and n18352_not n18353 ; n18354
g15919 and n17804 n18066_not ; n18355
g15920 and n17804_not n18336 ; n18356
g15921 nor n18355 n18356 ; n18357
g15922 and pi0644 n18357 ; n18358
g15923 and pi0644_not n18066 ; n18359
g15924 nor pi0715 n18359 ; n18360
g15925 and n18358_not n18360 ; n18361
g15926 and pi1160 n18361_not ; n18362
g15927 and n18354_not n18362 ; n18363
g15928 nor pi0644 n18351 ; n18364
g15929 and pi0644 n18133 ; n18365
g15930 nor pi0715 n18365 ; n18366
g15931 and n18364_not n18366 ; n18367
g15932 and pi0644_not n18357 ; n18368
g15933 and pi0644 n18066 ; n18369
g15934 and pi0715 n18369_not ; n18370
g15935 and n18368_not n18370 ; n18371
g15936 nor pi1160 n18371 ; n18372
g15937 and n18367_not n18372 ; n18373
g15938 and pi0790 n18363_not ; n18374
g15939 and n18373_not n18374 ; n18375
g15940 and pi0790_not n18351 ; n18376
g15941 nor po1038 n18376 ; n18377
g15942 and n18375_not n18377 ; n18378
g15943 and pi0141_not po1038 ; n18379
g15944 nor pi0832 n18379 ; n18380
g15945 and n18378_not n18380 ; n18381
g15946 nor pi0141 n2926 ; n18382
g15947 and pi0647_not n18382 ; n18383
g15948 and pi0706 n16645 ; n18384
g15949 nor n18382 n18384 ; n18385
g15950 and pi0778_not n18385 ; n18386
g15951 and pi0625_not n18384 ; n18387
g15952 nor n18385 n18387 ; n18388
g15953 and pi1153 n18388_not ; n18389
g15954 nor pi1153 n18382 ; n18390
g15955 and n18387_not n18390 ; n18391
g15956 nor n18389 n18391 ; n18392
g15957 and pi0778 n18392_not ; n18393
g15958 nor n18386 n18393 ; n18394
g15959 and n17845_not n18394 ; n18395
g15960 and n17847_not n18395 ; n18396
g15961 and n17849_not n18396 ; n18397
g15962 and n17851_not n18397 ; n18398
g15963 and n17857_not n18398 ; n18399
g15964 and pi0647 n18399 ; n18400
g15965 and pi1157 n18383_not ; n18401
g15966 and n18400_not n18401 ; n18402
g15967 and n17862_not n18398 ; n18403
g15968 and pi1156 n18403_not ; n18404
g15969 and n17871 n18397 ; n18405
g15970 and pi0626_not n18382 ; n18406
g15971 and pi0749 n17244 ; n18407
g15972 nor n18382 n18407 ; n18408
g15973 nor n17874 n18408 ; n18409
g15974 nor pi0785 n18409 ; n18410
g15975 nor n17879 n18408 ; n18411
g15976 and pi1155 n18411_not ; n18412
g15977 and n17882_not n18409 ; n18413
g15978 nor pi1155 n18413 ; n18414
g15979 nor n18412 n18414 ; n18415
g15980 and pi0785 n18415_not ; n18416
g15981 nor n18410 n18416 ; n18417
g15982 nor pi0781 n18417 ; n18418
g15983 and n17889_not n18417 ; n18419
g15984 and pi1154 n18419_not ; n18420
g15985 and n17892_not n18417 ; n18421
g15986 nor pi1154 n18421 ; n18422
g15987 nor n18420 n18422 ; n18423
g15988 and pi0781 n18423_not ; n18424
g15989 nor n18418 n18424 ; n18425
g15990 nor pi0789 n18425 ; n18426
g15991 and pi0619_not n18382 ; n18427
g15992 and pi0619 n18425 ; n18428
g15993 and pi1159 n18427_not ; n18429
g15994 and n18428_not n18429 ; n18430
g15995 and pi0619_not n18425 ; n18431
g15996 and pi0619 n18382 ; n18432
g15997 nor pi1159 n18432 ; n18433
g15998 and n18431_not n18433 ; n18434
g15999 nor n18430 n18434 ; n18435
g16000 and pi0789 n18435_not ; n18436
g16001 nor n18426 n18436 ; n18437
g16002 and pi0626 n18437 ; n18438
g16003 and pi1158 n18406_not ; n18439
g16004 and n18438_not n18439 ; n18440
g16005 and pi0626_not n18437 ; n18441
g16006 and pi0626 n18382 ; n18442
g16007 nor pi1158 n18442 ; n18443
g16008 and n18441_not n18443 ; n18444
g16009 nor n18440 n18444 ; n18445
g16010 and n16630_not n18445 ; n18446
g16011 nor n18405 n18446 ; n18447
g16012 and pi0788 n18447_not ; n18448
g16013 and pi0618 n18395 ; n18449
g16014 and pi0609 n18394 ; n18450
g16015 nor n17168 n18385 ; n18451
g16016 and pi0625 n18451 ; n18452
g16017 and n18408 n18451_not ; n18453
g16018 nor n18452 n18453 ; n18454
g16019 and n18390 n18454_not ; n18455
g16020 nor pi0608 n18389 ; n18456
g16021 and n18455_not n18456 ; n18457
g16022 and pi1153 n18408 ; n18458
g16023 and n18452_not n18458 ; n18459
g16024 and pi0608 n18391_not ; n18460
g16025 and n18459_not n18460 ; n18461
g16026 nor n18457 n18461 ; n18462
g16027 and pi0778 n18462_not ; n18463
g16028 nor pi0778 n18453 ; n18464
g16029 nor n18463 n18464 ; n18465
g16030 nor pi0609 n18465 ; n18466
g16031 nor pi1155 n18450 ; n18467
g16032 and n18466_not n18467 ; n18468
g16033 nor pi0660 n18412 ; n18469
g16034 and n18468_not n18469 ; n18470
g16035 and pi0609_not n18394 ; n18471
g16036 and pi0609 n18465_not ; n18472
g16037 and pi1155 n18471_not ; n18473
g16038 and n18472_not n18473 ; n18474
g16039 and pi0660 n18414_not ; n18475
g16040 and n18474_not n18475 ; n18476
g16041 nor n18470 n18476 ; n18477
g16042 and pi0785 n18477_not ; n18478
g16043 nor pi0785 n18465 ; n18479
g16044 nor n18478 n18479 ; n18480
g16045 nor pi0618 n18480 ; n18481
g16046 nor pi1154 n18449 ; n18482
g16047 and n18481_not n18482 ; n18483
g16048 nor pi0627 n18420 ; n18484
g16049 and n18483_not n18484 ; n18485
g16050 and pi0618_not n18395 ; n18486
g16051 and pi0618 n18480_not ; n18487
g16052 and pi1154 n18486_not ; n18488
g16053 and n18487_not n18488 ; n18489
g16054 and pi0627 n18422_not ; n18490
g16055 and n18489_not n18490 ; n18491
g16056 nor n18485 n18491 ; n18492
g16057 and pi0781 n18492_not ; n18493
g16058 nor pi0781 n18480 ; n18494
g16059 nor n18493 n18494 ; n18495
g16060 and pi0789_not n18495 ; n18496
g16061 nor pi0619 n18495 ; n18497
g16062 and pi0619 n18396 ; n18498
g16063 nor pi1159 n18498 ; n18499
g16064 and n18497_not n18499 ; n18500
g16065 nor pi0648 n18430 ; n18501
g16066 and n18500_not n18501 ; n18502
g16067 and pi0619_not n18396 ; n18503
g16068 and pi0619 n18495_not ; n18504
g16069 and pi1159 n18503_not ; n18505
g16070 and n18504_not n18505 ; n18506
g16071 and pi0648 n18434_not ; n18507
g16072 and n18506_not n18507 ; n18508
g16073 and pi0789 n18502_not ; n18509
g16074 and n18508_not n18509 ; n18510
g16075 and n17970 n18496_not ; n18511
g16076 and n18510_not n18511 ; n18512
g16077 nor n18448 n18512 ; n18513
g16078 nor pi0628 n18513 ; n18514
g16079 nor pi0788 n18437 ; n18515
g16080 and pi0788 n18445_not ; n18516
g16081 nor n18515 n18516 ; n18517
g16082 and pi0628 n18517 ; n18518
g16083 nor pi1156 n18518 ; n18519
g16084 and n18514_not n18519 ; n18520
g16085 nor pi0629 n18404 ; n18521
g16086 and n18520_not n18521 ; n18522
g16087 and n17997_not n18398 ; n18523
g16088 nor pi1156 n18523 ; n18524
g16089 and pi0628_not n18517 ; n18525
g16090 and pi0628 n18513_not ; n18526
g16091 and pi1156 n18525_not ; n18527
g16092 and n18526_not n18527 ; n18528
g16093 and pi0629 n18524_not ; n18529
g16094 and n18528_not n18529 ; n18530
g16095 nor n18522 n18530 ; n18531
g16096 and pi0792 n18531_not ; n18532
g16097 nor pi0792 n18513 ; n18533
g16098 nor n18532 n18533 ; n18534
g16099 nor pi0647 n18534 ; n18535
g16100 and n17779_not n18517 ; n18536
g16101 and n17779 n18382 ; n18537
g16102 nor n18536 n18537 ; n18538
g16103 and pi0647 n18538_not ; n18539
g16104 nor pi1157 n18539 ; n18540
g16105 and n18535_not n18540 ; n18541
g16106 nor pi0630 n18402 ; n18542
g16107 and n18541_not n18542 ; n18543
g16108 and pi0647_not n18399 ; n18544
g16109 and pi0647 n18382 ; n18545
g16110 nor pi1157 n18545 ; n18546
g16111 and n18544_not n18546 ; n18547
g16112 and pi0647 n18534_not ; n18548
g16113 nor pi0647 n18538 ; n18549
g16114 and pi1157 n18549_not ; n18550
g16115 and n18548_not n18550 ; n18551
g16116 and pi0630 n18547_not ; n18552
g16117 and n18551_not n18552 ; n18553
g16118 nor n18543 n18553 ; n18554
g16119 and pi0787 n18554_not ; n18555
g16120 nor pi0787 n18534 ; n18556
g16121 nor n18555 n18556 ; n18557
g16122 nor pi0790 n18557 ; n18558
g16123 nor pi0787 n18399 ; n18559
g16124 nor n18402 n18547 ; n18560
g16125 and pi0787 n18560_not ; n18561
g16126 nor n18559 n18561 ; n18562
g16127 and pi0644_not n18562 ; n18563
g16128 and pi0644 n18557_not ; n18564
g16129 and pi0715 n18563_not ; n18565
g16130 and n18564_not n18565 ; n18566
g16131 and n17804 n18382_not ; n18567
g16132 and n17804_not n18538 ; n18568
g16133 nor n18567 n18568 ; n18569
g16134 and pi0644 n18569 ; n18570
g16135 and pi0644_not n18382 ; n18571
g16136 nor pi0715 n18571 ; n18572
g16137 and n18570_not n18572 ; n18573
g16138 and pi1160 n18573_not ; n18574
g16139 and n18566_not n18574 ; n18575
g16140 and pi0644_not n18569 ; n18576
g16141 and pi0644 n18382 ; n18577
g16142 and pi0715 n18577_not ; n18578
g16143 and n18576_not n18578 ; n18579
g16144 and pi0644 n18562 ; n18580
g16145 nor pi0644 n18557 ; n18581
g16146 nor pi0715 n18580 ; n18582
g16147 and n18581_not n18582 ; n18583
g16148 nor pi1160 n18579 ; n18584
g16149 and n18583_not n18584 ; n18585
g16150 nor n18575 n18585 ; n18586
g16151 and pi0790 n18586_not ; n18587
g16152 and pi0832 n18558_not ; n18588
g16153 and n18587_not n18588 ; n18589
g16154 nor n18381 n18589 ; po0298
g16155 and n2571 n17051_not ; n18591
g16156 and pi0142 n18591_not ; n18592
g16157 and pi0039 n17025_not ; n18593
g16158 and pi0142 n18147_not ; n18594
g16159 and n18593_not n18594 ; n18595
g16160 and pi0142 n16970_not ; n18596
g16161 nor n6242 n18596 ; n18597
g16162 and pi0142 n16990_not ; n18598
g16163 and n6242 n18598_not ; n18599
g16164 and pi0215 n18599_not ; n18600
g16165 and n18597_not n18600 ; n18601
g16166 and pi0142 n16653_not ; n18602
g16167 and n3448 n18602_not ; n18603
g16168 and pi0142 n17018_not ; n18604
g16169 nor n6242 n18604 ; n18605
g16170 and pi0142 n17011_not ; n18606
g16171 and n6242 n18606_not ; n18607
g16172 nor n18605 n18607 ; n18608
g16173 nor n3448 n18608 ; n18609
g16174 nor pi0215 n18603 ; n18610
g16175 and n18609_not n18610 ; n18611
g16176 nor n18601 n18611 ; n18612
g16177 and pi0039 pi0299 ; n18613
g16178 and n18612_not n18613 ; n18614
g16179 nor n18595 n18614 ; n18615
g16180 and n14873 n18615_not ; n18616
g16181 nor n18592 n18616 ; n18617
g16182 and n16639 n18617_not ; n18618
g16183 and pi0142 n2571_not ; n18619
g16184 and pi0039 pi0142 ; n18620
g16185 and pi0038 n18620_not ; n18621
g16186 and pi0142 n16667_not ; n18622
g16187 and pi0735 n16645 ; n18623
g16188 and n2521 n18623 ; n18624
g16189 nor n18622 n18624 ; n18625
g16190 nor pi0039 n18625 ; n18626
g16191 and n18621 n18626_not ; n18627
g16192 nor pi0142 n16926 ; n18628
g16193 and pi0142 n16948 ; n18629
g16194 and pi0735 n18628_not ; n18630
g16195 and n18629_not n18630 ; n18631
g16196 and pi0142 pi0735_not ; n18632
g16197 and n16958_not n18632 ; n18633
g16198 nor n18631 n18633 ; n18634
g16199 nor pi0039 n18634 ; n18635
g16200 and n16652 n18623 ; n18636
g16201 nor n18602 n18636 ; n18637
g16202 and n3448 n18637 ; n18638
g16203 nor pi0142 n16694 ; n18639
g16204 and pi0142 n16791_not ; n18640
g16205 nor n18639 n18640 ; n18641
g16206 and pi0735 n18641_not ; n18642
g16207 nor pi0735 n18606 ; n18643
g16208 nor n18642 n18643 ; n18644
g16209 and n6242 n18644 ; n18645
g16210 and pi0142_not n16705 ; n18646
g16211 and pi0142 n16763 ; n18647
g16212 nor n18646 n18647 ; n18648
g16213 and pi0735 n18648_not ; n18649
g16214 nor pi0735 n18604 ; n18650
g16215 nor n18649 n18650 ; n18651
g16216 and n6242_not n18651 ; n18652
g16217 nor n3448 n18652 ; n18653
g16218 and n18645_not n18653 ; n18654
g16219 nor pi0215 n18638 ; n18655
g16220 and n18654_not n18655 ; n18656
g16221 nor pi0735 n18598 ; n18657
g16222 and pi0142_not n17560 ; n18658
g16223 and pi0142 n16811_not ; n18659
g16224 and pi0735 n18658_not ; n18660
g16225 and n18659_not n18660 ; n18661
g16226 nor n18657 n18661 ; n18662
g16227 and n6242 n18662_not ; n18663
g16228 nor pi0735 n18596 ; n18664
g16229 and pi0142 n16819_not ; n18665
g16230 and n17559 n18658 ; n18666
g16231 and pi0735 n18666_not ; n18667
g16232 and n18665_not n18667 ; n18668
g16233 nor n18664 n18668 ; n18669
g16234 nor n6242 n18669 ; n18670
g16235 and pi0215 n18663_not ; n18671
g16236 and n18670_not n18671 ; n18672
g16237 and pi0299 n18672_not ; n18673
g16238 and n18656_not n18673 ; n18674
g16239 and n6205 n18662_not ; n18675
g16240 nor n6205 n18669 ; n18676
g16241 and pi0223 n18675_not ; n18677
g16242 and n18676_not n18677 ; n18678
g16243 and n2603 n18637 ; n18679
g16244 and n6205 n18644 ; n18680
g16245 and n6205_not n18651 ; n18681
g16246 nor n2603 n18681 ; n18682
g16247 and n18680_not n18682 ; n18683
g16248 nor pi0223 n18679 ; n18684
g16249 and n18683_not n18684 ; n18685
g16250 nor pi0299 n18678 ; n18686
g16251 and n18685_not n18686 ; n18687
g16252 and pi0039 n18674_not ; n18688
g16253 and n18687_not n18688 ; n18689
g16254 nor pi0038 n18635 ; n18690
g16255 and n18689_not n18690 ; n18691
g16256 and n2571 n18627_not ; n18692
g16257 and n18691_not n18692 ; n18693
g16258 nor n18619 n18693 ; n18694
g16259 nor pi0778 n18694 ; n18695
g16260 and pi0625_not n18694 ; n18696
g16261 and pi0625 n18617 ; n18697
g16262 nor pi1153 n18697 ; n18698
g16263 and n18696_not n18698 ; n18699
g16264 and pi0625_not n18617 ; n18700
g16265 and pi0625 n18694 ; n18701
g16266 and pi1153 n18700_not ; n18702
g16267 and n18701_not n18702 ; n18703
g16268 nor n18699 n18703 ; n18704
g16269 and pi0778 n18704_not ; n18705
g16270 nor n18695 n18705 ; n18706
g16271 and n17075_not n18706 ; n18707
g16272 and n17075 n18617 ; n18708
g16273 nor n18707 n18708 ; n18709
g16274 and n16639_not n18709 ; n18710
g16275 nor n18618 n18710 ; n18711
g16276 and n16635_not n18711 ; n18712
g16277 and n16635 n18617 ; n18713
g16278 nor n18712 n18713 ; n18714
g16279 nor n16631 n18714 ; n18715
g16280 and n16631 n18617 ; n18716
g16281 nor n18715 n18716 ; n18717
g16282 and pi0792_not n18717 ; n18718
g16283 and pi0628_not n18617 ; n18719
g16284 and pi0628 n18717_not ; n18720
g16285 and pi1156 n18719_not ; n18721
g16286 and n18720_not n18721 ; n18722
g16287 and pi0628 n18617 ; n18723
g16288 nor pi0628 n18717 ; n18724
g16289 nor pi1156 n18723 ; n18725
g16290 and n18724_not n18725 ; n18726
g16291 nor n18722 n18726 ; n18727
g16292 and pi0792 n18727_not ; n18728
g16293 nor n18718 n18728 ; n18729
g16294 nor pi0787 n18729 ; n18730
g16295 and pi0647_not n18617 ; n18731
g16296 and pi0647 n18729 ; n18732
g16297 and pi1157 n18731_not ; n18733
g16298 and n18732_not n18733 ; n18734
g16299 and pi0647_not n18729 ; n18735
g16300 and pi0647 n18617 ; n18736
g16301 nor pi1157 n18736 ; n18737
g16302 and n18735_not n18737 ; n18738
g16303 nor n18734 n18738 ; n18739
g16304 and pi0787 n18739_not ; n18740
g16305 nor n18730 n18740 ; n18741
g16306 and pi0644_not n18741 ; n18742
g16307 and pi0618_not n18617 ; n18743
g16308 and pi0743 n17244 ; n18744
g16309 and n2521 n18744 ; n18745
g16310 nor n18622 n18745 ; n18746
g16311 nor pi0039 n18746 ; n18747
g16312 and n18621 n18747_not ; n18748
g16313 and pi0142 pi0743_not ; n18749
g16314 and n16930_not n18749 ; n18750
g16315 nor pi0142 n17226 ; n18751
g16316 and pi0142 n17137_not ; n18752
g16317 and pi0743 n18751_not ; n18753
g16318 and n18752_not n18753 ; n18754
g16319 nor pi0299 n18750 ; n18755
g16320 and n18754_not n18755 ; n18756
g16321 nor pi0142 n17231 ; n18757
g16322 and pi0142 n16941_not ; n18758
g16323 nor pi0743 n18758 ; n18759
g16324 and pi0142 n17124 ; n18760
g16325 nor n18757 n18759 ; n18761
g16326 and n18760_not n18761 ; n18762
g16327 and pi0299 n18762_not ; n18763
g16328 nor n18756 n18763 ; n18764
g16329 and pi0039_not n18764 ; n18765
g16330 nor pi0743 n18596 ; n18766
g16331 and pi0142 n17189_not ; n18767
g16332 and pi0743 n17558 ; n18768
g16333 and n18767_not n18768 ; n18769
g16334 nor n18766 n18769 ; n18770
g16335 nor n6205 n18770 ; n18771
g16336 nor pi0743 n18598 ; n18772
g16337 and pi0142 n17200 ; n18773
g16338 and pi0743 n17241 ; n18774
g16339 and n18773_not n18774 ; n18775
g16340 nor n18772 n18775 ; n18776
g16341 and n6205 n18776_not ; n18777
g16342 and pi0223 n18777_not ; n18778
g16343 and n18771_not n18778 ; n18779
g16344 nor pi0743 n18604 ; n18780
g16345 and pi0142 n17157_not ; n18781
g16346 and pi0743 n17254_not ; n18782
g16347 and n18781_not n18782 ; n18783
g16348 nor n18780 n18783 ; n18784
g16349 and n6205_not n18784 ; n18785
g16350 and pi0142_not n17252 ; n18786
g16351 and pi0142 n17175 ; n18787
g16352 nor n18786 n18787 ; n18788
g16353 and pi0743 n18788_not ; n18789
g16354 nor pi0743 n18606 ; n18790
g16355 nor n18789 n18790 ; n18791
g16356 and n6205 n18791 ; n18792
g16357 nor n2603 n18785 ; n18793
g16358 and n18792_not n18793 ; n18794
g16359 and pi0743 n17235 ; n18795
g16360 nor n18602 n18795 ; n18796
g16361 and n2603 n18796 ; n18797
g16362 nor pi0223 n18797 ; n18798
g16363 and n18794_not n18798 ; n18799
g16364 nor pi0299 n18779 ; n18800
g16365 and n18799_not n18800 ; n18801
g16366 and n3448 n18796_not ; n18802
g16367 and n6242_not n18784 ; n18803
g16368 and n6242 n18791 ; n18804
g16369 nor n18803 n18804 ; n18805
g16370 nor n3448 n18805 ; n18806
g16371 nor pi0215 n18802 ; n18807
g16372 and n18806_not n18807 ; n18808
g16373 and n6242_not n18770 ; n18809
g16374 and n6242 n18776 ; n18810
g16375 and pi0215 n18810_not ; n18811
g16376 and n18809_not n18811 ; n18812
g16377 nor n18808 n18812 ; n18813
g16378 and pi0299 n18813_not ; n18814
g16379 and pi0039 n18801_not ; n18815
g16380 and n18814_not n18815 ; n18816
g16381 nor pi0038 n18765 ; n18817
g16382 and n18816_not n18817 ; n18818
g16383 and n2571 n18748_not ; n18819
g16384 and n18818_not n18819 ; n18820
g16385 nor n18619 n18820 ; n18821
g16386 nor n17117 n18821 ; n18822
g16387 and n17117 n18617_not ; n18823
g16388 nor n18822 n18823 ; n18824
g16389 nor pi0785 n18824 ; n18825
g16390 nor n17291 n18617 ; n18826
g16391 and pi0609 n18822 ; n18827
g16392 nor n18826 n18827 ; n18828
g16393 and pi1155 n18828_not ; n18829
g16394 nor n17296 n18617 ; n18830
g16395 and pi0609_not n18822 ; n18831
g16396 nor n18830 n18831 ; n18832
g16397 nor pi1155 n18832 ; n18833
g16398 nor n18829 n18833 ; n18834
g16399 and pi0785 n18834_not ; n18835
g16400 nor n18825 n18835 ; n18836
g16401 and pi0618 n18836 ; n18837
g16402 and pi1154 n18743_not ; n18838
g16403 and n18837_not n18838 ; n18839
g16404 and pi0609 n18706 ; n18840
g16405 and pi0625_not n18821 ; n18841
g16406 and pi0735_not n18764 ; n18842
g16407 and n16937 n18752 ; n18843
g16408 and n16919_not n18751 ; n18844
g16409 nor n18843 n18844 ; n18845
g16410 and pi0743 n18845_not ; n18846
g16411 and pi0142 n16937_not ; n18847
g16412 and n17226_not n18847 ; n18848
g16413 and pi0142_not n17618 ; n18849
g16414 nor pi0743 n18848 ; n18850
g16415 and n18849_not n18850 ; n18851
g16416 nor pi0299 n18851 ; n18852
g16417 and n18846_not n18852 ; n18853
g16418 and n16924_not n18757 ; n18854
g16419 and n16945_not n18760 ; n18855
g16420 nor n18854 n18855 ; n18856
g16421 and pi0743 n18856_not ; n18857
g16422 and pi0142_not n17623 ; n18858
g16423 and pi0142 n16946_not ; n18859
g16424 and n17231_not n18859 ; n18860
g16425 nor pi0743 n18860 ; n18861
g16426 and n18858_not n18861 ; n18862
g16427 and pi0299 n18857_not ; n18863
g16428 and n18862_not n18863 ; n18864
g16429 nor n18853 n18864 ; n18865
g16430 and pi0735 n18865_not ; n18866
g16431 nor pi0039 n18842 ; n18867
g16432 and n18866_not n18867 ; n18868
g16433 nor pi0142 n17556 ; n18869
g16434 and pi0142 n17519_not ; n18870
g16435 and pi0743 n18869_not ; n18871
g16436 and n18870_not n18871 ; n18872
g16437 and pi0142_not n17448 ; n18873
g16438 and pi0142 n17351 ; n18874
g16439 nor pi0743 n18873 ; n18875
g16440 and n18874_not n18875 ; n18876
g16441 nor n18872 n18876 ; n18877
g16442 and pi0735 n18877_not ; n18878
g16443 and pi0735_not n18776 ; n18879
g16444 nor n18878 n18879 ; n18880
g16445 and n6205 n18880 ; n18881
g16446 and pi0142_not n17562 ; n18882
g16447 and pi0142 n17527 ; n18883
g16448 and pi0743 n18882_not ; n18884
g16449 and n18883_not n18884 ; n18885
g16450 nor pi0142 n17463 ; n18886
g16451 and pi0142 n17333 ; n18887
g16452 nor pi0743 n18887 ; n18888
g16453 and n18886_not n18888 ; n18889
g16454 nor n18885 n18889 ; n18890
g16455 and pi0735 n18890_not ; n18891
g16456 and pi0735_not n18770 ; n18892
g16457 nor n18891 n18892 ; n18893
g16458 and n6205_not n18893 ; n18894
g16459 and pi0223 n18881_not ; n18895
g16460 and n18894_not n18895 ; n18896
g16461 and pi0735_not n18796 ; n18897
g16462 and n17645_not n18746 ; n18898
g16463 nor n16650 n18898 ; n18899
g16464 and pi0735 n18899_not ; n18900
g16465 and n18602_not n18900 ; n18901
g16466 nor n18897 n18901 ; n18902
g16467 and n2603 n18902_not ; n18903
g16468 and pi0142 n17510 ; n18904
g16469 nor pi0142 n17573 ; n18905
g16470 and pi0743 n18904_not ; n18906
g16471 and n18905_not n18906 ; n18907
g16472 and pi0142_not n17420 ; n18908
g16473 and pi0142 n17373 ; n18909
g16474 nor pi0743 n18908 ; n18910
g16475 and n18909_not n18910 ; n18911
g16476 nor n18907 n18911 ; n18912
g16477 and pi0735 n18912_not ; n18913
g16478 and pi0735_not n18791 ; n18914
g16479 nor n18913 n18914 ; n18915
g16480 and n6205 n18915_not ; n18916
g16481 nor pi0142 n17584 ; n18917
g16482 and pi0142 n17499 ; n18918
g16483 and pi0743 n18918_not ; n18919
g16484 and n18917_not n18919 ; n18920
g16485 nor pi0142 n17438 ; n18921
g16486 and pi0142 n17383 ; n18922
g16487 nor pi0743 n18922 ; n18923
g16488 and n18921_not n18923 ; n18924
g16489 nor n18920 n18924 ; n18925
g16490 and pi0735 n18925_not ; n18926
g16491 and pi0735_not n18784 ; n18927
g16492 nor n18926 n18927 ; n18928
g16493 nor n6205 n18928 ; n18929
g16494 nor n2603 n18929 ; n18930
g16495 and n18916_not n18930 ; n18931
g16496 nor pi0223 n18903 ; n18932
g16497 and n18931_not n18932 ; n18933
g16498 nor n18896 n18933 ; n18934
g16499 nor pi0299 n18934 ; n18935
g16500 and n6242 n18880 ; n18936
g16501 and n6242_not n18893 ; n18937
g16502 and pi0215 n18936_not ; n18938
g16503 and n18937_not n18938 ; n18939
g16504 and n3448 n18902_not ; n18940
g16505 nor n6242 n18928 ; n18941
g16506 and n6242 n18915_not ; n18942
g16507 nor n3448 n18941 ; n18943
g16508 and n18942_not n18943 ; n18944
g16509 nor pi0215 n18940 ; n18945
g16510 and n18944_not n18945 ; n18946
g16511 nor n18939 n18946 ; n18947
g16512 and pi0299 n18947_not ; n18948
g16513 and pi0039 n18935_not ; n18949
g16514 and n18948_not n18949 ; n18950
g16515 nor n18868 n18950 ; n18951
g16516 nor pi0038 n18951 ; n18952
g16517 and pi0735 n17645 ; n18953
g16518 and n18746 n18953_not ; n18954
g16519 nor pi0039 n18954 ; n18955
g16520 and n18621 n18955_not ; n18956
g16521 and n2571 n18956_not ; n18957
g16522 and n18952_not n18957 ; n18958
g16523 nor n18619 n18958 ; n18959
g16524 and pi0625 n18959 ; n18960
g16525 and pi1153 n18841_not ; n18961
g16526 and n18960_not n18961 ; n18962
g16527 and pi0608 n18699_not ; n18963
g16528 and n18962_not n18963 ; n18964
g16529 and pi0625_not n18959 ; n18965
g16530 and pi0625 n18821 ; n18966
g16531 nor pi1153 n18966 ; n18967
g16532 and n18965_not n18967 ; n18968
g16533 nor pi0608 n18703 ; n18969
g16534 and n18968_not n18969 ; n18970
g16535 nor n18964 n18970 ; n18971
g16536 and pi0778 n18971_not ; n18972
g16537 and pi0778_not n18959 ; n18973
g16538 nor n18972 n18973 ; n18974
g16539 nor pi0609 n18974 ; n18975
g16540 nor pi1155 n18840 ; n18976
g16541 and n18975_not n18976 ; n18977
g16542 nor pi0660 n18829 ; n18978
g16543 and n18977_not n18978 ; n18979
g16544 and pi0609_not n18706 ; n18980
g16545 and pi0609 n18974_not ; n18981
g16546 and pi1155 n18980_not ; n18982
g16547 and n18981_not n18982 ; n18983
g16548 and pi0660 n18833_not ; n18984
g16549 and n18983_not n18984 ; n18985
g16550 nor n18979 n18985 ; n18986
g16551 and pi0785 n18986_not ; n18987
g16552 nor pi0785 n18974 ; n18988
g16553 nor n18987 n18988 ; n18989
g16554 nor pi0618 n18989 ; n18990
g16555 and pi0618 n18709_not ; n18991
g16556 nor pi1154 n18991 ; n18992
g16557 and n18990_not n18992 ; n18993
g16558 nor pi0627 n18839 ; n18994
g16559 and n18993_not n18994 ; n18995
g16560 and pi0618_not n18836 ; n18996
g16561 and pi0618 n18617 ; n18997
g16562 nor pi1154 n18997 ; n18998
g16563 and n18996_not n18998 ; n18999
g16564 and pi0618 n18989_not ; n19000
g16565 nor pi0618 n18709 ; n19001
g16566 and pi1154 n19001_not ; n19002
g16567 and n19000_not n19002 ; n19003
g16568 and pi0627 n18999_not ; n19004
g16569 and n19003_not n19004 ; n19005
g16570 nor n18995 n19005 ; n19006
g16571 and pi0781 n19006_not ; n19007
g16572 nor pi0781 n18989 ; n19008
g16573 nor n19007 n19008 ; n19009
g16574 nor pi0619 n19009 ; n19010
g16575 and pi0619 n18711 ; n19011
g16576 nor pi1159 n19011 ; n19012
g16577 and n19010_not n19012 ; n19013
g16578 and pi0619_not n18617 ; n19014
g16579 nor pi0781 n18836 ; n19015
g16580 nor n18839 n18999 ; n19016
g16581 and pi0781 n19016_not ; n19017
g16582 nor n19015 n19017 ; n19018
g16583 and pi0619 n19018 ; n19019
g16584 and pi1159 n19014_not ; n19020
g16585 and n19019_not n19020 ; n19021
g16586 nor pi0648 n19021 ; n19022
g16587 and n19013_not n19022 ; n19023
g16588 and pi0619 n19009_not ; n19024
g16589 and pi0619_not n18711 ; n19025
g16590 and pi1159 n19025_not ; n19026
g16591 and n19024_not n19026 ; n19027
g16592 and pi0619_not n19018 ; n19028
g16593 and pi0619 n18617 ; n19029
g16594 nor pi1159 n19029 ; n19030
g16595 and n19028_not n19030 ; n19031
g16596 and pi0648 n19031_not ; n19032
g16597 and n19027_not n19032 ; n19033
g16598 nor n19023 n19033 ; n19034
g16599 and pi0789 n19034_not ; n19035
g16600 nor pi0789 n19009 ; n19036
g16601 nor n19035 n19036 ; n19037
g16602 and pi0788_not n19037 ; n19038
g16603 and pi0626_not n19037 ; n19039
g16604 and pi0626 n18714 ; n19040
g16605 nor pi0641 n19040 ; n19041
g16606 and n19039_not n19041 ; n19042
g16607 nor pi0789 n19018 ; n19043
g16608 nor n19021 n19031 ; n19044
g16609 and pi0789 n19044_not ; n19045
g16610 nor n19043 n19045 ; n19046
g16611 and pi0626_not n19046 ; n19047
g16612 and pi0626 n18617 ; n19048
g16613 nor pi1158 n19048 ; n19049
g16614 and n19047_not n19049 ; n19050
g16615 nor n17730 n19050 ; n19051
g16616 nor n19042 n19051 ; n19052
g16617 and pi0626 n19037 ; n19053
g16618 and pi0626_not n18714 ; n19054
g16619 and pi0641 n19054_not ; n19055
g16620 and n19053_not n19055 ; n19056
g16621 and pi0626_not n18617 ; n19057
g16622 and pi0626 n19046 ; n19058
g16623 and pi1158 n19057_not ; n19059
g16624 and n19058_not n19059 ; n19060
g16625 nor n17745 n19060 ; n19061
g16626 nor n19056 n19061 ; n19062
g16627 nor n19052 n19062 ; n19063
g16628 and pi0788 n19063_not ; n19064
g16629 nor n19038 n19064 ; n19065
g16630 and pi0628_not n19065 ; n19066
g16631 nor n19050 n19060 ; n19067
g16632 and pi0788 n19067_not ; n19068
g16633 nor pi0788 n19046 ; n19069
g16634 nor n19068 n19069 ; n19070
g16635 and pi0628 n19070 ; n19071
g16636 nor pi1156 n19071 ; n19072
g16637 and n19066_not n19072 ; n19073
g16638 nor pi0629 n18722 ; n19074
g16639 and n19073_not n19074 ; n19075
g16640 and pi0628 n19065 ; n19076
g16641 and pi0628_not n19070 ; n19077
g16642 and pi1156 n19077_not ; n19078
g16643 and n19076_not n19078 ; n19079
g16644 and pi0629 n18726_not ; n19080
g16645 and n19079_not n19080 ; n19081
g16646 nor n19075 n19081 ; n19082
g16647 and pi0792 n19082_not ; n19083
g16648 and pi0792_not n19065 ; n19084
g16649 nor n19083 n19084 ; n19085
g16650 nor pi0647 n19085 ; n19086
g16651 and n17779_not n19070 ; n19087
g16652 and n17779 n18617 ; n19088
g16653 nor n19087 n19088 ; n19089
g16654 and pi0647 n19089_not ; n19090
g16655 nor pi1157 n19090 ; n19091
g16656 and n19086_not n19091 ; n19092
g16657 nor pi0630 n18734 ; n19093
g16658 and n19092_not n19093 ; n19094
g16659 and pi0647 n19085_not ; n19095
g16660 nor pi0647 n19089 ; n19096
g16661 and pi1157 n19096_not ; n19097
g16662 and n19095_not n19097 ; n19098
g16663 and pi0630 n18738_not ; n19099
g16664 and n19098_not n19099 ; n19100
g16665 nor n19094 n19100 ; n19101
g16666 and pi0787 n19101_not ; n19102
g16667 nor pi0787 n19085 ; n19103
g16668 nor n19102 n19103 ; n19104
g16669 and pi0644 n19104_not ; n19105
g16670 and pi0715 n18742_not ; n19106
g16671 and n19105_not n19106 ; n19107
g16672 and n17804 n18617_not ; n19108
g16673 and n17804_not n19089 ; n19109
g16674 nor n19108 n19109 ; n19110
g16675 and pi0644 n19110 ; n19111
g16676 and pi0644_not n18617 ; n19112
g16677 nor pi0715 n19112 ; n19113
g16678 and n19111_not n19113 ; n19114
g16679 and pi1160 n19114_not ; n19115
g16680 and n19107_not n19115 ; n19116
g16681 nor pi0644 n19104 ; n19117
g16682 and pi0644 n18741 ; n19118
g16683 nor pi0715 n19118 ; n19119
g16684 and n19117_not n19119 ; n19120
g16685 and pi0644_not n19110 ; n19121
g16686 and pi0644 n18617 ; n19122
g16687 and pi0715 n19122_not ; n19123
g16688 and n19121_not n19123 ; n19124
g16689 nor pi1160 n19124 ; n19125
g16690 and n19120_not n19125 ; n19126
g16691 and pi0790 n19116_not ; n19127
g16692 and n19126_not n19127 ; n19128
g16693 and pi0790_not n19104 ; n19129
g16694 and n6305 n19129_not ; n19130
g16695 and n19128_not n19130 ; n19131
g16696 nor pi0142 n6305 ; n19132
g16697 nor pi0057 n19132 ; n19133
g16698 and n19131_not n19133 ; n19134
g16699 and pi0057 pi0142 ; n19135
g16700 nor pi0832 n19135 ; n19136
g16701 and n19134_not n19136 ; n19137
g16702 and pi0142 n2926_not ; n19138
g16703 and pi0628 pi1156 ; n19139
g16704 nor pi0628 pi1156 ; n19140
g16705 and pi0792 n19139_not ; n19141
g16706 and n19140_not n19141 ; n19142
g16707 and pi0625_not pi1153 ; n19143
g16708 and pi0625 pi1153_not ; n19144
g16709 nor n19143 n19144 ; n19145
g16710 and pi0778 n19145_not ; n19146
g16711 and n18623 n19146_not ; n19147
g16712 nor n19138 n19147 ; n19148
g16713 nor n16631 n16635 ; n19149
g16714 nor n16639 n17075 ; n19150
g16715 and n19149 n19150 ; n19151
g16716 and n19148_not n19151 ; n19152
g16717 and n19142_not n19152 ; n19153
g16718 and pi0647 n19153 ; n19154
g16719 and pi1157 n19138_not ; n19155
g16720 and n19154_not n19155 ; n19156
g16721 and pi0628 n19152 ; n19157
g16722 nor n19138 n19157 ; n19158
g16723 and pi1156 n19158_not ; n19159
g16724 and pi0626_not n19138 ; n19160
g16725 and n17117_not n18744 ; n19161
g16726 and pi0609 n19161 ; n19162
g16727 and pi1155 n19138_not ; n19163
g16728 and n19162_not n19163 ; n19164
g16729 and pi0609_not n19161 ; n19165
g16730 nor pi1155 n19138 ; n19166
g16731 and n19165_not n19166 ; n19167
g16732 nor n19164 n19167 ; n19168
g16733 and pi0785 n19168_not ; n19169
g16734 nor pi0785 n19138 ; n19170
g16735 and n19161_not n19170 ; n19171
g16736 nor n19169 n19171 ; n19172
g16737 nor pi0781 n19172 ; n19173
g16738 and pi0618_not n19138 ; n19174
g16739 and pi0618 n19172 ; n19175
g16740 and pi1154 n19174_not ; n19176
g16741 and n19175_not n19176 ; n19177
g16742 and pi0618_not n19172 ; n19178
g16743 and pi0618 n19138 ; n19179
g16744 nor pi1154 n19179 ; n19180
g16745 and n19178_not n19180 ; n19181
g16746 nor n19177 n19181 ; n19182
g16747 and pi0781 n19182_not ; n19183
g16748 nor n19173 n19183 ; n19184
g16749 nor pi0789 n19184 ; n19185
g16750 and pi0619_not n19138 ; n19186
g16751 and pi0619 n19184 ; n19187
g16752 and pi1159 n19186_not ; n19188
g16753 and n19187_not n19188 ; n19189
g16754 and pi0619_not n19184 ; n19190
g16755 and pi0619 n19138 ; n19191
g16756 nor pi1159 n19191 ; n19192
g16757 and n19190_not n19192 ; n19193
g16758 nor n19189 n19193 ; n19194
g16759 and pi0789 n19194_not ; n19195
g16760 nor n19185 n19195 ; n19196
g16761 and pi0626 n19196 ; n19197
g16762 and pi1158 n19160_not ; n19198
g16763 and n19197_not n19198 ; n19199
g16764 and pi0626_not n19196 ; n19200
g16765 and pi0626 n19138 ; n19201
g16766 nor pi1158 n19201 ; n19202
g16767 and n19200_not n19202 ; n19203
g16768 nor n19199 n19203 ; n19204
g16769 and n16630_not n19204 ; n19205
g16770 and n16635 n19138_not ; n19206
g16771 nor n17075 n19148 ; n19207
g16772 and n16639_not n19207 ; n19208
g16773 nor n19138 n19208 ; n19209
g16774 and n17871 n19206_not ; n19210
g16775 and n19209_not n19210 ; n19211
g16776 nor n19205 n19211 ; n19212
g16777 and pi0788 n19212_not ; n19213
g16778 nor n19138 n19207 ; n19214
g16779 and pi0618 n19214_not ; n19215
g16780 and pi0625 n18623 ; n19216
g16781 and pi1153 n19138_not ; n19217
g16782 and n19216_not n19217 ; n19218
g16783 and pi0735 n17469 ; n19219
g16784 and pi0625 n19219 ; n19220
g16785 nor n18744 n19138 ; n19221
g16786 and n19219_not n19221 ; n19222
g16787 nor n19220 n19222 ; n19223
g16788 nor pi1153 n19223 ; n19224
g16789 nor pi0608 n19218 ; n19225
g16790 and n19224_not n19225 ; n19226
g16791 nor n18744 n19220 ; n19227
g16792 and pi1153 n19227_not ; n19228
g16793 nor pi0625 pi1153 ; n19229
g16794 and n18623 n19229 ; n19230
g16795 nor n19138 n19230 ; n19231
g16796 and n19228_not n19231 ; n19232
g16797 and pi0608 n19232_not ; n19233
g16798 nor n19226 n19233 ; n19234
g16799 and pi0778 n19234_not ; n19235
g16800 nor pi0778 n19222 ; n19236
g16801 nor n19235 n19236 ; n19237
g16802 nor pi0609 n19237 ; n19238
g16803 and pi0609 n19148_not ; n19239
g16804 nor pi1155 n19239 ; n19240
g16805 and n19238_not n19240 ; n19241
g16806 nor pi0660 n19164 ; n19242
g16807 and n19241_not n19242 ; n19243
g16808 and pi0609 n19237_not ; n19244
g16809 nor pi0609 n19148 ; n19245
g16810 and pi1155 n19245_not ; n19246
g16811 and n19244_not n19246 ; n19247
g16812 and pi0660 n19167_not ; n19248
g16813 and n19247_not n19248 ; n19249
g16814 nor n19243 n19249 ; n19250
g16815 and pi0785 n19250_not ; n19251
g16816 nor pi0785 n19237 ; n19252
g16817 nor n19251 n19252 ; n19253
g16818 nor pi0618 n19253 ; n19254
g16819 nor pi1154 n19215 ; n19255
g16820 and n19254_not n19255 ; n19256
g16821 nor pi0627 n19177 ; n19257
g16822 and n19256_not n19257 ; n19258
g16823 nor pi0618 n19214 ; n19259
g16824 and pi0618 n19253_not ; n19260
g16825 and pi1154 n19259_not ; n19261
g16826 and n19260_not n19261 ; n19262
g16827 and pi0627 n19181_not ; n19263
g16828 and n19262_not n19263 ; n19264
g16829 nor n19258 n19264 ; n19265
g16830 and pi0781 n19265_not ; n19266
g16831 nor pi0781 n19253 ; n19267
g16832 nor n19266 n19267 ; n19268
g16833 and pi0789_not n19268 ; n19269
g16834 nor pi0619 n19268 ; n19270
g16835 and pi0619 n19209_not ; n19271
g16836 nor pi1159 n19271 ; n19272
g16837 and n19270_not n19272 ; n19273
g16838 nor pi0648 n19189 ; n19274
g16839 and n19273_not n19274 ; n19275
g16840 and pi0619 n19268_not ; n19276
g16841 nor pi0619 n19209 ; n19277
g16842 and pi1159 n19277_not ; n19278
g16843 and n19276_not n19278 ; n19279
g16844 and pi0648 n19193_not ; n19280
g16845 and n19279_not n19280 ; n19281
g16846 and pi0789 n19275_not ; n19282
g16847 and n19281_not n19282 ; n19283
g16848 and n17970 n19269_not ; n19284
g16849 and n19283_not n19284 ; n19285
g16850 nor n19213 n19285 ; n19286
g16851 and pi0628_not n19286 ; n19287
g16852 nor pi0788 n19196 ; n19288
g16853 and pi0788 n19204_not ; n19289
g16854 nor n19288 n19289 ; n19290
g16855 and pi0628 n19290_not ; n19291
g16856 nor pi1156 n19291 ; n19292
g16857 and n19287_not n19292 ; n19293
g16858 nor pi0629 n19159 ; n19294
g16859 and n19293_not n19294 ; n19295
g16860 and pi0628_not n19152 ; n19296
g16861 nor n19138 n19296 ; n19297
g16862 nor pi1156 n19297 ; n19298
g16863 and pi0628 n19286 ; n19299
g16864 nor pi0628 n19290 ; n19300
g16865 and pi1156 n19300_not ; n19301
g16866 and n19299_not n19301 ; n19302
g16867 and pi0629 n19298_not ; n19303
g16868 and n19302_not n19303 ; n19304
g16869 nor n19295 n19304 ; n19305
g16870 and pi0792 n19305_not ; n19306
g16871 and pi0792_not n19286 ; n19307
g16872 nor n19306 n19307 ; n19308
g16873 and pi0647_not n19308 ; n19309
g16874 and n17779_not n19290 ; n19310
g16875 and n17779 n19138 ; n19311
g16876 nor n19310 n19311 ; n19312
g16877 and pi0647 n19312_not ; n19313
g16878 nor pi1157 n19313 ; n19314
g16879 and n19309_not n19314 ; n19315
g16880 nor pi0630 n19156 ; n19316
g16881 and n19315_not n19316 ; n19317
g16882 and pi0647_not n19153 ; n19318
g16883 nor pi1157 n19138 ; n19319
g16884 and n19318_not n19319 ; n19320
g16885 nor pi0647 n19312 ; n19321
g16886 and pi0647 n19308 ; n19322
g16887 and pi1157 n19321_not ; n19323
g16888 and n19322_not n19323 ; n19324
g16889 and pi0630 n19320_not ; n19325
g16890 and n19324_not n19325 ; n19326
g16891 nor n19317 n19326 ; n19327
g16892 and pi0787 n19327_not ; n19328
g16893 and pi0787_not n19308 ; n19329
g16894 nor n19328 n19329 ; n19330
g16895 nor pi0790 n19330 ; n19331
g16896 and n17804 n19138_not ; n19332
g16897 and n17804_not n19312 ; n19333
g16898 nor n19332 n19333 ; n19334
g16899 and pi0644 n19334 ; n19335
g16900 and pi0644_not n19138 ; n19336
g16901 nor pi0715 n19336 ; n19337
g16902 and n19335_not n19337 ; n19338
g16903 and pi0647_not pi1157 ; n19339
g16904 and pi0647 pi1157_not ; n19340
g16905 nor n19339 n19340 ; n19341
g16906 and pi0787 n19341_not ; n19342
g16907 and n19153 n19342_not ; n19343
g16908 nor n19138 n19343 ; n19344
g16909 nor pi0644 n19344 ; n19345
g16910 and pi0644 n19330_not ; n19346
g16911 and pi0715 n19345_not ; n19347
g16912 and n19346_not n19347 ; n19348
g16913 and pi1160 n19338_not ; n19349
g16914 and n19348_not n19349 ; n19350
g16915 and pi0644_not n19334 ; n19351
g16916 and pi0644 n19138 ; n19352
g16917 and pi0715 n19352_not ; n19353
g16918 and n19351_not n19353 ; n19354
g16919 and pi0644 n19344_not ; n19355
g16920 nor pi0644 n19330 ; n19356
g16921 nor pi0715 n19355 ; n19357
g16922 and n19356_not n19357 ; n19358
g16923 nor pi1160 n19354 ; n19359
g16924 and n19358_not n19359 ; n19360
g16925 nor n19350 n19360 ; n19361
g16926 and pi0790 n19361_not ; n19362
g16927 and pi0832 n19331_not ; n19363
g16928 and n19362_not n19363 ; n19364
g16929 nor n19137 n19364 ; po0299
g16930 nor pi0143 n17059 ; n19366
g16931 and n16635 n19366_not ; n19367
g16932 and pi0143 n2571_not ; n19368
g16933 nor pi0143 n17052 ; n19369
g16934 and pi0687_not n19369 ; n19370
g16935 nor pi0143 n16641 ; n19371
g16936 and n16647 n19371_not ; n19372
g16937 and pi0143_not n18072 ; n19373
g16938 and pi0143 n18076_not ; n19374
g16939 nor pi0038 n19374 ; n19375
g16940 and n19373_not n19375 ; n19376
g16941 and pi0687 n19372_not ; n19377
g16942 and n19376_not n19377 ; n19378
g16943 and n2571 n19370_not ; n19379
g16944 and n19378_not n19379 ; n19380
g16945 nor n19368 n19380 ; n19381
g16946 nor pi0778 n19381 ; n19382
g16947 and pi0625_not n19366 ; n19383
g16948 and pi0625 n19381 ; n19384
g16949 and pi1153 n19383_not ; n19385
g16950 and n19384_not n19385 ; n19386
g16951 and pi0625_not n19381 ; n19387
g16952 and pi0625 n19366 ; n19388
g16953 nor pi1153 n19388 ; n19389
g16954 and n19387_not n19389 ; n19390
g16955 nor n19386 n19390 ; n19391
g16956 and pi0778 n19391_not ; n19392
g16957 nor n19382 n19392 ; n19393
g16958 nor n17075 n19393 ; n19394
g16959 and n17075 n19366_not ; n19395
g16960 nor n19394 n19395 ; n19396
g16961 and n16639_not n19396 ; n19397
g16962 and n16639 n19366 ; n19398
g16963 nor n19397 n19398 ; n19399
g16964 and n16635_not n19399 ; n19400
g16965 nor n19367 n19400 ; n19401
g16966 and n16631_not n19401 ; n19402
g16967 and n16631 n19366 ; n19403
g16968 nor n19402 n19403 ; n19404
g16969 and pi0792_not n19404 ; n19405
g16970 and pi0628_not n19366 ; n19406
g16971 and pi0628 n19404_not ; n19407
g16972 and pi1156 n19406_not ; n19408
g16973 and n19407_not n19408 ; n19409
g16974 and pi0628 n19366 ; n19410
g16975 nor pi0628 n19404 ; n19411
g16976 nor pi1156 n19410 ; n19412
g16977 and n19411_not n19412 ; n19413
g16978 nor n19409 n19413 ; n19414
g16979 and pi0792 n19414_not ; n19415
g16980 nor n19405 n19415 ; n19416
g16981 nor pi0787 n19416 ; n19417
g16982 and pi0647_not n19366 ; n19418
g16983 and pi0647 n19416 ; n19419
g16984 and pi1157 n19418_not ; n19420
g16985 and n19419_not n19420 ; n19421
g16986 and pi0647_not n19416 ; n19422
g16987 and pi0647 n19366 ; n19423
g16988 nor pi1157 n19423 ; n19424
g16989 and n19422_not n19424 ; n19425
g16990 nor n19421 n19425 ; n19426
g16991 and pi0787 n19426_not ; n19427
g16992 nor n19417 n19427 ; n19428
g16993 and pi0644_not n19428 ; n19429
g16994 and pi0618_not n19366 ; n19430
g16995 and pi0774 n19369_not ; n19431
g16996 and n6135 n17244 ; n19432
g16997 and pi0038 n19432 ; n19433
g16998 and pi0038_not n17275 ; n19434
g16999 and pi0143 n19434_not ; n19435
g17000 nor pi0038 n17221 ; n19436
g17001 and n6284 n17182 ; n19437
g17002 and pi0038 n19437_not ; n19438
g17003 nor n19436 n19438 ; n19439
g17004 nor pi0143 pi0774 ; n19440
g17005 and n19439 n19440 ; n19441
g17006 nor n19435 n19441 ; n19442
g17007 nor n19433 n19442 ; n19443
g17008 nor n19431 n19443 ; n19444
g17009 and n2571 n19444_not ; n19445
g17010 nor n19368 n19445 ; n19446
g17011 nor n17117 n19446 ; n19447
g17012 and n17117 n19366_not ; n19448
g17013 nor n19447 n19448 ; n19449
g17014 nor pi0785 n19449 ; n19450
g17015 nor n17291 n19366 ; n19451
g17016 and pi0609 n19447 ; n19452
g17017 nor n19451 n19452 ; n19453
g17018 and pi1155 n19453_not ; n19454
g17019 nor n17296 n19366 ; n19455
g17020 and pi0609_not n19447 ; n19456
g17021 nor n19455 n19456 ; n19457
g17022 nor pi1155 n19457 ; n19458
g17023 nor n19454 n19458 ; n19459
g17024 and pi0785 n19459_not ; n19460
g17025 nor n19450 n19460 ; n19461
g17026 and pi0618 n19461 ; n19462
g17027 and pi1154 n19430_not ; n19463
g17028 and n19462_not n19463 ; n19464
g17029 nor pi0039 n17625 ; n19465
g17030 and pi0039 n17485_not ; n19466
g17031 nor n19465 n19466 ; n19467
g17032 and pi0038_not n19467 ; n19468
g17033 and pi0143 n19468 ; n19469
g17034 and pi0038 n18175 ; n19470
g17035 and n16641 n17355_not ; n19471
g17036 and pi0038 n19471 ; n19472
g17037 and pi0039 n17404_not ; n19473
g17038 nor pi0039 n17612 ; n19474
g17039 nor n19473 n19474 ; n19475
g17040 nor pi0038 n19475 ; n19476
g17041 nor n19472 n19476 ; n19477
g17042 and pi0143_not n19477 ; n19478
g17043 and pi0774 n19470_not ; n19479
g17044 and n19469_not n19479 ; n19480
g17045 and n19478_not n19480 ; n19481
g17046 nor pi0039 n17629 ; n19482
g17047 and pi0038_not n19482 ; n19483
g17048 and pi0039 n17546_not ; n19484
g17049 and pi0039_not n17490 ; n19485
g17050 and pi0038 n19485_not ; n19486
g17051 nor n19483 n19486 ; n19487
g17052 and n19484_not n19487 ; n19488
g17053 nor pi0143 n19488 ; n19489
g17054 and n6284 n17470_not ; n19490
g17055 and pi0038 n19490_not ; n19491
g17056 and pi0039 n17605_not ; n19492
g17057 and n16926_not n17234 ; n19493
g17058 nor n19492 n19493 ; n19494
g17059 nor pi0038 n19494 ; n19495
g17060 nor n19491 n19495 ; n19496
g17061 and pi0143 n19496 ; n19497
g17062 nor pi0774 n19489 ; n19498
g17063 and n19497_not n19498 ; n19499
g17064 and pi0687 n19499_not ; n19500
g17065 and n19481_not n19500 ; n19501
g17066 and pi0687_not n19444 ; n19502
g17067 and n2571 n19501_not ; n19503
g17068 and n19502_not n19503 ; n19504
g17069 nor n19368 n19504 ; n19505
g17070 and pi0625_not n19505 ; n19506
g17071 and pi0625 n19446 ; n19507
g17072 nor pi1153 n19507 ; n19508
g17073 and n19506_not n19508 ; n19509
g17074 nor pi0608 n19386 ; n19510
g17075 and n19509_not n19510 ; n19511
g17076 and pi0625_not n19446 ; n19512
g17077 and pi0625 n19505 ; n19513
g17078 and pi1153 n19512_not ; n19514
g17079 and n19513_not n19514 ; n19515
g17080 and pi0608 n19390_not ; n19516
g17081 and n19515_not n19516 ; n19517
g17082 nor n19511 n19517 ; n19518
g17083 and pi0778 n19518_not ; n19519
g17084 and pi0778_not n19505 ; n19520
g17085 nor n19519 n19520 ; n19521
g17086 nor pi0609 n19521 ; n19522
g17087 and pi0609 n19393 ; n19523
g17088 nor pi1155 n19523 ; n19524
g17089 and n19522_not n19524 ; n19525
g17090 nor pi0660 n19454 ; n19526
g17091 and n19525_not n19526 ; n19527
g17092 and pi0609_not n19393 ; n19528
g17093 and pi0609 n19521_not ; n19529
g17094 and pi1155 n19528_not ; n19530
g17095 and n19529_not n19530 ; n19531
g17096 and pi0660 n19458_not ; n19532
g17097 and n19531_not n19532 ; n19533
g17098 nor n19527 n19533 ; n19534
g17099 and pi0785 n19534_not ; n19535
g17100 nor pi0785 n19521 ; n19536
g17101 nor n19535 n19536 ; n19537
g17102 nor pi0618 n19537 ; n19538
g17103 and pi0618 n19396 ; n19539
g17104 nor pi1154 n19539 ; n19540
g17105 and n19538_not n19540 ; n19541
g17106 nor pi0627 n19464 ; n19542
g17107 and n19541_not n19542 ; n19543
g17108 and pi0618_not n19461 ; n19544
g17109 and pi0618 n19366 ; n19545
g17110 nor pi1154 n19545 ; n19546
g17111 and n19544_not n19546 ; n19547
g17112 and pi0618_not n19396 ; n19548
g17113 and pi0618 n19537_not ; n19549
g17114 and pi1154 n19548_not ; n19550
g17115 and n19549_not n19550 ; n19551
g17116 and pi0627 n19547_not ; n19552
g17117 and n19551_not n19552 ; n19553
g17118 nor n19543 n19553 ; n19554
g17119 and pi0781 n19554_not ; n19555
g17120 nor pi0781 n19537 ; n19556
g17121 nor n19555 n19556 ; n19557
g17122 nor pi0619 n19557 ; n19558
g17123 and pi0619 n19399_not ; n19559
g17124 nor pi1159 n19559 ; n19560
g17125 and n19558_not n19560 ; n19561
g17126 and pi0619_not n19366 ; n19562
g17127 nor pi0781 n19461 ; n19563
g17128 nor n19464 n19547 ; n19564
g17129 and pi0781 n19564_not ; n19565
g17130 nor n19563 n19565 ; n19566
g17131 and pi0619 n19566 ; n19567
g17132 and pi1159 n19562_not ; n19568
g17133 and n19567_not n19568 ; n19569
g17134 nor pi0648 n19569 ; n19570
g17135 and n19561_not n19570 ; n19571
g17136 and pi0619 n19557_not ; n19572
g17137 nor pi0619 n19399 ; n19573
g17138 and pi1159 n19573_not ; n19574
g17139 and n19572_not n19574 ; n19575
g17140 and pi0619_not n19566 ; n19576
g17141 and pi0619 n19366 ; n19577
g17142 nor pi1159 n19577 ; n19578
g17143 and n19576_not n19578 ; n19579
g17144 and pi0648 n19579_not ; n19580
g17145 and n19575_not n19580 ; n19581
g17146 nor n19571 n19581 ; n19582
g17147 and pi0789 n19582_not ; n19583
g17148 nor pi0789 n19557 ; n19584
g17149 nor n19583 n19584 ; n19585
g17150 and pi0788_not n19585 ; n19586
g17151 and pi0626_not n19585 ; n19587
g17152 and pi0626 n19401_not ; n19588
g17153 nor pi0641 n19588 ; n19589
g17154 and n19587_not n19589 ; n19590
g17155 nor pi0789 n19566 ; n19591
g17156 nor n19569 n19579 ; n19592
g17157 and pi0789 n19592_not ; n19593
g17158 nor n19591 n19593 ; n19594
g17159 and pi0626_not n19594 ; n19595
g17160 and pi0626 n19366 ; n19596
g17161 nor pi1158 n19596 ; n19597
g17162 and n19595_not n19597 ; n19598
g17163 nor n17730 n19598 ; n19599
g17164 nor n19590 n19599 ; n19600
g17165 and pi0626 n19585 ; n19601
g17166 nor pi0626 n19401 ; n19602
g17167 and pi0641 n19602_not ; n19603
g17168 and n19601_not n19603 ; n19604
g17169 and pi0626_not n19366 ; n19605
g17170 and pi0626 n19594 ; n19606
g17171 and pi1158 n19605_not ; n19607
g17172 and n19606_not n19607 ; n19608
g17173 nor n17745 n19608 ; n19609
g17174 nor n19604 n19609 ; n19610
g17175 nor n19600 n19610 ; n19611
g17176 and pi0788 n19611_not ; n19612
g17177 nor n19586 n19612 ; n19613
g17178 and pi0628_not n19613 ; n19614
g17179 nor n19598 n19608 ; n19615
g17180 and pi0788 n19615_not ; n19616
g17181 nor pi0788 n19594 ; n19617
g17182 nor n19616 n19617 ; n19618
g17183 and pi0628 n19618 ; n19619
g17184 nor pi1156 n19619 ; n19620
g17185 and n19614_not n19620 ; n19621
g17186 nor pi0629 n19409 ; n19622
g17187 and n19621_not n19622 ; n19623
g17188 and pi0628 n19613 ; n19624
g17189 and pi0628_not n19618 ; n19625
g17190 and pi1156 n19625_not ; n19626
g17191 and n19624_not n19626 ; n19627
g17192 and pi0629 n19413_not ; n19628
g17193 and n19627_not n19628 ; n19629
g17194 nor n19623 n19629 ; n19630
g17195 and pi0792 n19630_not ; n19631
g17196 and pi0792_not n19613 ; n19632
g17197 nor n19631 n19632 ; n19633
g17198 nor pi0647 n19633 ; n19634
g17199 and n17779_not n19618 ; n19635
g17200 and n17779 n19366 ; n19636
g17201 nor n19635 n19636 ; n19637
g17202 and pi0647 n19637_not ; n19638
g17203 nor pi1157 n19638 ; n19639
g17204 and n19634_not n19639 ; n19640
g17205 nor pi0630 n19421 ; n19641
g17206 and n19640_not n19641 ; n19642
g17207 and pi0647 n19633_not ; n19643
g17208 nor pi0647 n19637 ; n19644
g17209 and pi1157 n19644_not ; n19645
g17210 and n19643_not n19645 ; n19646
g17211 and pi0630 n19425_not ; n19647
g17212 and n19646_not n19647 ; n19648
g17213 nor n19642 n19648 ; n19649
g17214 and pi0787 n19649_not ; n19650
g17215 nor pi0787 n19633 ; n19651
g17216 nor n19650 n19651 ; n19652
g17217 and pi0644 n19652_not ; n19653
g17218 and pi0715 n19429_not ; n19654
g17219 and n19653_not n19654 ; n19655
g17220 and n17804 n19366_not ; n19656
g17221 and n17804_not n19637 ; n19657
g17222 nor n19656 n19657 ; n19658
g17223 and pi0644 n19658 ; n19659
g17224 and pi0644_not n19366 ; n19660
g17225 nor pi0715 n19660 ; n19661
g17226 and n19659_not n19661 ; n19662
g17227 and pi1160 n19662_not ; n19663
g17228 and n19655_not n19663 ; n19664
g17229 nor pi0644 n19652 ; n19665
g17230 and pi0644 n19428 ; n19666
g17231 nor pi0715 n19666 ; n19667
g17232 and n19665_not n19667 ; n19668
g17233 and pi0644_not n19658 ; n19669
g17234 and pi0644 n19366 ; n19670
g17235 and pi0715 n19670_not ; n19671
g17236 and n19669_not n19671 ; n19672
g17237 nor pi1160 n19672 ; n19673
g17238 and n19668_not n19673 ; n19674
g17239 and pi0790 n19664_not ; n19675
g17240 and n19674_not n19675 ; n19676
g17241 and pi0790_not n19652 ; n19677
g17242 nor po1038 n19677 ; n19678
g17243 and n19676_not n19678 ; n19679
g17244 and pi0143_not po1038 ; n19680
g17245 nor pi0832 n19680 ; n19681
g17246 and n19679_not n19681 ; n19682
g17247 nor pi0143 n2926 ; n19683
g17248 and pi0647_not n19683 ; n19684
g17249 and pi0687 n16645 ; n19685
g17250 nor n19683 n19685 ; n19686
g17251 and pi0778_not n19686 ; n19687
g17252 and pi0625_not n19685 ; n19688
g17253 nor n19686 n19688 ; n19689
g17254 and pi1153 n19689_not ; n19690
g17255 nor pi1153 n19683 ; n19691
g17256 and n19688_not n19691 ; n19692
g17257 nor n19690 n19692 ; n19693
g17258 and pi0778 n19693_not ; n19694
g17259 nor n19687 n19694 ; n19695
g17260 and n17845_not n19695 ; n19696
g17261 and n17847_not n19696 ; n19697
g17262 and n17849_not n19697 ; n19698
g17263 and n17851_not n19698 ; n19699
g17264 and n17857_not n19699 ; n19700
g17265 and pi0647 n19700 ; n19701
g17266 and pi1157 n19684_not ; n19702
g17267 and n19701_not n19702 ; n19703
g17268 and n17862_not n19699 ; n19704
g17269 and pi1156 n19704_not ; n19705
g17270 and n17871 n19698 ; n19706
g17271 and pi0626_not n19683 ; n19707
g17272 and pi0774_not n17244 ; n19708
g17273 nor n19683 n19708 ; n19709
g17274 nor n17874 n19709 ; n19710
g17275 nor pi0785 n19710 ; n19711
g17276 nor n17879 n19709 ; n19712
g17277 and pi1155 n19712_not ; n19713
g17278 and n17882_not n19710 ; n19714
g17279 nor pi1155 n19714 ; n19715
g17280 nor n19713 n19715 ; n19716
g17281 and pi0785 n19716_not ; n19717
g17282 nor n19711 n19717 ; n19718
g17283 nor pi0781 n19718 ; n19719
g17284 and n17889_not n19718 ; n19720
g17285 and pi1154 n19720_not ; n19721
g17286 and n17892_not n19718 ; n19722
g17287 nor pi1154 n19722 ; n19723
g17288 nor n19721 n19723 ; n19724
g17289 and pi0781 n19724_not ; n19725
g17290 nor n19719 n19725 ; n19726
g17291 nor pi0789 n19726 ; n19727
g17292 and pi0619_not n19683 ; n19728
g17293 and pi0619 n19726 ; n19729
g17294 and pi1159 n19728_not ; n19730
g17295 and n19729_not n19730 ; n19731
g17296 and pi0619_not n19726 ; n19732
g17297 and pi0619 n19683 ; n19733
g17298 nor pi1159 n19733 ; n19734
g17299 and n19732_not n19734 ; n19735
g17300 nor n19731 n19735 ; n19736
g17301 and pi0789 n19736_not ; n19737
g17302 nor n19727 n19737 ; n19738
g17303 and pi0626 n19738 ; n19739
g17304 and pi1158 n19707_not ; n19740
g17305 and n19739_not n19740 ; n19741
g17306 and pi0626_not n19738 ; n19742
g17307 and pi0626 n19683 ; n19743
g17308 nor pi1158 n19743 ; n19744
g17309 and n19742_not n19744 ; n19745
g17310 nor n19741 n19745 ; n19746
g17311 and n16630_not n19746 ; n19747
g17312 nor n19706 n19747 ; n19748
g17313 and pi0788 n19748_not ; n19749
g17314 and pi0618 n19696 ; n19750
g17315 and pi0609 n19695 ; n19751
g17316 nor n17168 n19686 ; n19752
g17317 and pi0625 n19752 ; n19753
g17318 and n19709 n19752_not ; n19754
g17319 nor n19753 n19754 ; n19755
g17320 and n19691 n19755_not ; n19756
g17321 nor pi0608 n19690 ; n19757
g17322 and n19756_not n19757 ; n19758
g17323 and pi1153 n19709 ; n19759
g17324 and n19753_not n19759 ; n19760
g17325 and pi0608 n19692_not ; n19761
g17326 and n19760_not n19761 ; n19762
g17327 nor n19758 n19762 ; n19763
g17328 and pi0778 n19763_not ; n19764
g17329 nor pi0778 n19754 ; n19765
g17330 nor n19764 n19765 ; n19766
g17331 nor pi0609 n19766 ; n19767
g17332 nor pi1155 n19751 ; n19768
g17333 and n19767_not n19768 ; n19769
g17334 nor pi0660 n19713 ; n19770
g17335 and n19769_not n19770 ; n19771
g17336 and pi0609_not n19695 ; n19772
g17337 and pi0609 n19766_not ; n19773
g17338 and pi1155 n19772_not ; n19774
g17339 and n19773_not n19774 ; n19775
g17340 and pi0660 n19715_not ; n19776
g17341 and n19775_not n19776 ; n19777
g17342 nor n19771 n19777 ; n19778
g17343 and pi0785 n19778_not ; n19779
g17344 nor pi0785 n19766 ; n19780
g17345 nor n19779 n19780 ; n19781
g17346 nor pi0618 n19781 ; n19782
g17347 nor pi1154 n19750 ; n19783
g17348 and n19782_not n19783 ; n19784
g17349 nor pi0627 n19721 ; n19785
g17350 and n19784_not n19785 ; n19786
g17351 and pi0618_not n19696 ; n19787
g17352 and pi0618 n19781_not ; n19788
g17353 and pi1154 n19787_not ; n19789
g17354 and n19788_not n19789 ; n19790
g17355 and pi0627 n19723_not ; n19791
g17356 and n19790_not n19791 ; n19792
g17357 nor n19786 n19792 ; n19793
g17358 and pi0781 n19793_not ; n19794
g17359 nor pi0781 n19781 ; n19795
g17360 nor n19794 n19795 ; n19796
g17361 and pi0789_not n19796 ; n19797
g17362 nor pi0619 n19796 ; n19798
g17363 and pi0619 n19697 ; n19799
g17364 nor pi1159 n19799 ; n19800
g17365 and n19798_not n19800 ; n19801
g17366 nor pi0648 n19731 ; n19802
g17367 and n19801_not n19802 ; n19803
g17368 and pi0619_not n19697 ; n19804
g17369 and pi0619 n19796_not ; n19805
g17370 and pi1159 n19804_not ; n19806
g17371 and n19805_not n19806 ; n19807
g17372 and pi0648 n19735_not ; n19808
g17373 and n19807_not n19808 ; n19809
g17374 and pi0789 n19803_not ; n19810
g17375 and n19809_not n19810 ; n19811
g17376 and n17970 n19797_not ; n19812
g17377 and n19811_not n19812 ; n19813
g17378 nor n19749 n19813 ; n19814
g17379 nor pi0628 n19814 ; n19815
g17380 nor pi0788 n19738 ; n19816
g17381 and pi0788 n19746_not ; n19817
g17382 nor n19816 n19817 ; n19818
g17383 and pi0628 n19818 ; n19819
g17384 nor pi1156 n19819 ; n19820
g17385 and n19815_not n19820 ; n19821
g17386 nor pi0629 n19705 ; n19822
g17387 and n19821_not n19822 ; n19823
g17388 and n17997_not n19699 ; n19824
g17389 nor pi1156 n19824 ; n19825
g17390 and pi0628_not n19818 ; n19826
g17391 and pi0628 n19814_not ; n19827
g17392 and pi1156 n19826_not ; n19828
g17393 and n19827_not n19828 ; n19829
g17394 and pi0629 n19825_not ; n19830
g17395 and n19829_not n19830 ; n19831
g17396 nor n19823 n19831 ; n19832
g17397 and pi0792 n19832_not ; n19833
g17398 nor pi0792 n19814 ; n19834
g17399 nor n19833 n19834 ; n19835
g17400 nor pi0647 n19835 ; n19836
g17401 and n17779_not n19818 ; n19837
g17402 and n17779 n19683 ; n19838
g17403 nor n19837 n19838 ; n19839
g17404 and pi0647 n19839_not ; n19840
g17405 nor pi1157 n19840 ; n19841
g17406 and n19836_not n19841 ; n19842
g17407 nor pi0630 n19703 ; n19843
g17408 and n19842_not n19843 ; n19844
g17409 and pi0647_not n19700 ; n19845
g17410 and pi0647 n19683 ; n19846
g17411 nor pi1157 n19846 ; n19847
g17412 and n19845_not n19847 ; n19848
g17413 and pi0647 n19835_not ; n19849
g17414 nor pi0647 n19839 ; n19850
g17415 and pi1157 n19850_not ; n19851
g17416 and n19849_not n19851 ; n19852
g17417 and pi0630 n19848_not ; n19853
g17418 and n19852_not n19853 ; n19854
g17419 nor n19844 n19854 ; n19855
g17420 and pi0787 n19855_not ; n19856
g17421 nor pi0787 n19835 ; n19857
g17422 nor n19856 n19857 ; n19858
g17423 nor pi0790 n19858 ; n19859
g17424 nor pi0787 n19700 ; n19860
g17425 nor n19703 n19848 ; n19861
g17426 and pi0787 n19861_not ; n19862
g17427 nor n19860 n19862 ; n19863
g17428 and pi0644_not n19863 ; n19864
g17429 and pi0644 n19858_not ; n19865
g17430 and pi0715 n19864_not ; n19866
g17431 and n19865_not n19866 ; n19867
g17432 and n17804 n19683_not ; n19868
g17433 and n17804_not n19839 ; n19869
g17434 nor n19868 n19869 ; n19870
g17435 and pi0644 n19870 ; n19871
g17436 and pi0644_not n19683 ; n19872
g17437 nor pi0715 n19872 ; n19873
g17438 and n19871_not n19873 ; n19874
g17439 and pi1160 n19874_not ; n19875
g17440 and n19867_not n19875 ; n19876
g17441 and pi0644_not n19870 ; n19877
g17442 and pi0644 n19683 ; n19878
g17443 and pi0715 n19878_not ; n19879
g17444 and n19877_not n19879 ; n19880
g17445 and pi0644 n19863 ; n19881
g17446 nor pi0644 n19858 ; n19882
g17447 nor pi0715 n19881 ; n19883
g17448 and n19882_not n19883 ; n19884
g17449 nor pi1160 n19880 ; n19885
g17450 and n19884_not n19885 ; n19886
g17451 nor n19876 n19886 ; n19887
g17452 and pi0790 n19887_not ; n19888
g17453 and pi0832 n19859_not ; n19889
g17454 and n19888_not n19889 ; n19890
g17455 nor n19682 n19890 ; po0300
g17456 and pi0144 n17059_not ; n19892
g17457 and n16635 n19892_not ; n19893
g17458 and n17075 n19892_not ; n19894
g17459 and pi0736 n2571 ; n19895
g17460 nor n19892 n19895 ; n19896
g17461 nor pi0144 n16641 ; n19897
g17462 and n16641 n16644_not ; n19898
g17463 and pi0038 n19898_not ; n19899
g17464 and n19897_not n19899 ; n19900
g17465 and pi0144_not n18076 ; n19901
g17466 and pi0144 n18072_not ; n19902
g17467 nor pi0038 n19901 ; n19903
g17468 and n19902_not n19903 ; n19904
g17469 and n19895 n19900_not ; n19905
g17470 and n19904_not n19905 ; n19906
g17471 nor n19896 n19906 ; n19907
g17472 and pi0778_not n19907 ; n19908
g17473 nor pi0625 n19892 ; n19909
g17474 and pi0625 n19907_not ; n19910
g17475 and pi1153 n19909_not ; n19911
g17476 and n19910_not n19911 ; n19912
g17477 nor pi0625 n19907 ; n19913
g17478 and pi0625 n19892_not ; n19914
g17479 nor pi1153 n19914 ; n19915
g17480 and n19913_not n19915 ; n19916
g17481 nor n19912 n19916 ; n19917
g17482 and pi0778 n19917_not ; n19918
g17483 nor n19908 n19918 ; n19919
g17484 and n17075_not n19919 ; n19920
g17485 nor n19894 n19920 ; n19921
g17486 and n16639_not n19921 ; n19922
g17487 and n16639 n19892 ; n19923
g17488 nor n19922 n19923 ; n19924
g17489 and n16635_not n19924 ; n19925
g17490 nor n19893 n19925 ; n19926
g17491 and n16631_not n19926 ; n19927
g17492 and n16631 n19892 ; n19928
g17493 nor n19927 n19928 ; n19929
g17494 nor pi0792 n19929 ; n19930
g17495 nor pi0628 n19892 ; n19931
g17496 and pi0628 n19929 ; n19932
g17497 and pi1156 n19931_not ; n19933
g17498 and n19932_not n19933 ; n19934
g17499 and pi0628 n19892_not ; n19935
g17500 and pi0628_not n19929 ; n19936
g17501 nor pi1156 n19935 ; n19937
g17502 and n19936_not n19937 ; n19938
g17503 nor n19934 n19938 ; n19939
g17504 and pi0792 n19939_not ; n19940
g17505 nor n19930 n19940 ; n19941
g17506 nor pi0787 n19941 ; n19942
g17507 nor pi0647 n19892 ; n19943
g17508 and pi0647 n19941 ; n19944
g17509 and pi1157 n19943_not ; n19945
g17510 and n19944_not n19945 ; n19946
g17511 and pi0647 n19892_not ; n19947
g17512 and pi0647_not n19941 ; n19948
g17513 nor pi1157 n19947 ; n19949
g17514 and n19948_not n19949 ; n19950
g17515 nor n19946 n19950 ; n19951
g17516 and pi0787 n19951_not ; n19952
g17517 nor n19942 n19952 ; n19953
g17518 and pi0644_not n19953 ; n19954
g17519 nor pi0619 n19892 ; n19955
g17520 and n17117 n19892_not ; n19956
g17521 and pi0144 n2571_not ; n19957
g17522 nor pi0758 n17046 ; n19958
g17523 and pi0758 n17219 ; n19959
g17524 nor n19958 n19959 ; n19960
g17525 and pi0039 n19960_not ; n19961
g17526 and pi0758_not n16958 ; n19962
g17527 and pi0758 n17139 ; n19963
g17528 nor pi0039 n19962 ; n19964
g17529 and n19963_not n19964 ; n19965
g17530 nor n19961 n19965 ; n19966
g17531 and pi0144 n19966_not ; n19967
g17532 and pi0144_not pi0758 ; n19968
g17533 and n17275 n19968 ; n19969
g17534 nor n19967 n19969 ; n19970
g17535 nor pi0038 n19970 ; n19971
g17536 and pi0758 n17168 ; n19972
g17537 and n16641 n19972_not ; n19973
g17538 and pi0038 n19897_not ; n19974
g17539 and n19973_not n19974 ; n19975
g17540 nor n19971 n19975 ; n19976
g17541 and n2571 n19976_not ; n19977
g17542 nor n19957 n19977 ; n19978
g17543 and n17117_not n19978 ; n19979
g17544 nor n19956 n19979 ; n19980
g17545 and pi0785_not n19980 ; n19981
g17546 nor pi0609 n19892 ; n19982
g17547 and pi0609 n19980_not ; n19983
g17548 and pi1155 n19982_not ; n19984
g17549 and n19983_not n19984 ; n19985
g17550 nor pi0609 n19980 ; n19986
g17551 and pi0609 n19892_not ; n19987
g17552 nor pi1155 n19987 ; n19988
g17553 and n19986_not n19988 ; n19989
g17554 nor n19985 n19989 ; n19990
g17555 and pi0785 n19990_not ; n19991
g17556 nor n19981 n19991 ; n19992
g17557 nor pi0781 n19992 ; n19993
g17558 nor pi0618 n19892 ; n19994
g17559 and pi0618 n19992 ; n19995
g17560 and pi1154 n19994_not ; n19996
g17561 and n19995_not n19996 ; n19997
g17562 and pi0618 n19892_not ; n19998
g17563 and pi0618_not n19992 ; n19999
g17564 nor pi1154 n19998 ; n20000
g17565 and n19999_not n20000 ; n20001
g17566 nor n19997 n20001 ; n20002
g17567 and pi0781 n20002_not ; n20003
g17568 nor n19993 n20003 ; n20004
g17569 and pi0619 n20004 ; n20005
g17570 and pi1159 n19955_not ; n20006
g17571 and n20005_not n20006 ; n20007
g17572 and pi0736_not n19976 ; n20008
g17573 nor pi0144 n17605 ; n20009
g17574 and pi0144 n17546 ; n20010
g17575 and pi0758 n20010_not ; n20011
g17576 and n20009_not n20011 ; n20012
g17577 and pi0144 n17404_not ; n20013
g17578 nor pi0144 n17485 ; n20014
g17579 nor pi0758 n20014 ; n20015
g17580 and n20013_not n20015 ; n20016
g17581 and pi0039 n20012_not ; n20017
g17582 and n20016_not n20017 ; n20018
g17583 and pi0144_not n17631 ; n20019
g17584 and pi0144 n17629 ; n20020
g17585 and pi0758 n20019_not ; n20021
g17586 and n20020_not n20021 ; n20022
g17587 nor pi0144 n17625 ; n20023
g17588 and pi0144 n17612_not ; n20024
g17589 nor pi0758 n20023 ; n20025
g17590 and n20024_not n20025 ; n20026
g17591 nor pi0039 n20022 ; n20027
g17592 and n20026_not n20027 ; n20028
g17593 nor pi0038 n20028 ; n20029
g17594 and n20018_not n20029 ; n20030
g17595 and pi0736 n19470_not ; n20031
g17596 and n19975_not n20031 ; n20032
g17597 and n20030_not n20032 ; n20033
g17598 and n2571 n20033_not ; n20034
g17599 and n20008_not n20034 ; n20035
g17600 nor n19957 n20035 ; n20036
g17601 and pi0625_not n20036 ; n20037
g17602 and pi0625 n19978 ; n20038
g17603 nor pi1153 n20038 ; n20039
g17604 and n20037_not n20039 ; n20040
g17605 nor pi0608 n19912 ; n20041
g17606 and n20040_not n20041 ; n20042
g17607 and pi0625_not n19978 ; n20043
g17608 and pi0625 n20036 ; n20044
g17609 and pi1153 n20043_not ; n20045
g17610 and n20044_not n20045 ; n20046
g17611 and pi0608 n19916_not ; n20047
g17612 and n20046_not n20047 ; n20048
g17613 nor n20042 n20048 ; n20049
g17614 and pi0778 n20049_not ; n20050
g17615 and pi0778_not n20036 ; n20051
g17616 nor n20050 n20051 ; n20052
g17617 nor pi0609 n20052 ; n20053
g17618 and pi0609 n19919 ; n20054
g17619 nor pi1155 n20054 ; n20055
g17620 and n20053_not n20055 ; n20056
g17621 nor pi0660 n19985 ; n20057
g17622 and n20056_not n20057 ; n20058
g17623 and pi0609_not n19919 ; n20059
g17624 and pi0609 n20052_not ; n20060
g17625 and pi1155 n20059_not ; n20061
g17626 and n20060_not n20061 ; n20062
g17627 and pi0660 n19989_not ; n20063
g17628 and n20062_not n20063 ; n20064
g17629 nor n20058 n20064 ; n20065
g17630 and pi0785 n20065_not ; n20066
g17631 nor pi0785 n20052 ; n20067
g17632 nor n20066 n20067 ; n20068
g17633 nor pi0618 n20068 ; n20069
g17634 and pi0618 n19921_not ; n20070
g17635 nor pi1154 n20070 ; n20071
g17636 and n20069_not n20071 ; n20072
g17637 nor pi0627 n19997 ; n20073
g17638 and n20072_not n20073 ; n20074
g17639 and pi0618 n20068_not ; n20075
g17640 nor pi0618 n19921 ; n20076
g17641 and pi1154 n20076_not ; n20077
g17642 and n20075_not n20077 ; n20078
g17643 and pi0627 n20001_not ; n20079
g17644 and n20078_not n20079 ; n20080
g17645 nor n20074 n20080 ; n20081
g17646 and pi0781 n20081_not ; n20082
g17647 nor pi0781 n20068 ; n20083
g17648 nor n20082 n20083 ; n20084
g17649 nor pi0619 n20084 ; n20085
g17650 and pi0619 n19924 ; n20086
g17651 nor pi1159 n20086 ; n20087
g17652 and n20085_not n20087 ; n20088
g17653 nor pi0648 n20007 ; n20089
g17654 and n20088_not n20089 ; n20090
g17655 and pi0619 n19892_not ; n20091
g17656 and pi0619_not n20004 ; n20092
g17657 nor pi1159 n20091 ; n20093
g17658 and n20092_not n20093 ; n20094
g17659 and pi0619_not n19924 ; n20095
g17660 and pi0619 n20084_not ; n20096
g17661 and pi1159 n20095_not ; n20097
g17662 and n20096_not n20097 ; n20098
g17663 and pi0648 n20094_not ; n20099
g17664 and n20098_not n20099 ; n20100
g17665 nor n20090 n20100 ; n20101
g17666 and pi0789 n20101_not ; n20102
g17667 nor pi0789 n20084 ; n20103
g17668 nor n20102 n20103 ; n20104
g17669 and pi0788_not n20104 ; n20105
g17670 and pi0626_not n20104 ; n20106
g17671 and pi0626 n19926 ; n20107
g17672 nor pi0641 n20107 ; n20108
g17673 and n20106_not n20108 ; n20109
g17674 nor pi0789 n20004 ; n20110
g17675 nor n20007 n20094 ; n20111
g17676 and pi0789 n20111_not ; n20112
g17677 nor n20110 n20112 ; n20113
g17678 and pi0626_not n20113 ; n20114
g17679 and pi0626 n19892_not ; n20115
g17680 nor pi1158 n20115 ; n20116
g17681 and n20114_not n20116 ; n20117
g17682 nor n17730 n20117 ; n20118
g17683 nor n20109 n20118 ; n20119
g17684 and pi0626 n20104 ; n20120
g17685 and pi0626_not n19926 ; n20121
g17686 and pi0641 n20121_not ; n20122
g17687 and n20120_not n20122 ; n20123
g17688 and pi0626 n20113 ; n20124
g17689 nor pi0626 n19892 ; n20125
g17690 and pi1158 n20125_not ; n20126
g17691 and n20124_not n20126 ; n20127
g17692 nor n17745 n20127 ; n20128
g17693 nor n20123 n20128 ; n20129
g17694 nor n20119 n20129 ; n20130
g17695 and pi0788 n20130_not ; n20131
g17696 nor n20105 n20131 ; n20132
g17697 and pi0628_not n20132 ; n20133
g17698 nor n20117 n20127 ; n20134
g17699 and pi0788 n20134_not ; n20135
g17700 nor pi0788 n20113 ; n20136
g17701 nor n20135 n20136 ; n20137
g17702 and pi0628 n20137 ; n20138
g17703 nor pi1156 n20138 ; n20139
g17704 and n20133_not n20139 ; n20140
g17705 nor pi0629 n19934 ; n20141
g17706 and n20140_not n20141 ; n20142
g17707 and pi0628 n20132 ; n20143
g17708 and pi0628_not n20137 ; n20144
g17709 and pi1156 n20144_not ; n20145
g17710 and n20143_not n20145 ; n20146
g17711 and pi0629 n19938_not ; n20147
g17712 and n20146_not n20147 ; n20148
g17713 nor n20142 n20148 ; n20149
g17714 and pi0792 n20149_not ; n20150
g17715 and pi0792_not n20132 ; n20151
g17716 nor n20150 n20151 ; n20152
g17717 nor pi0647 n20152 ; n20153
g17718 nor n17779 n20137 ; n20154
g17719 and n17779 n19892 ; n20155
g17720 nor n20154 n20155 ; n20156
g17721 and pi0647 n20156 ; n20157
g17722 nor pi1157 n20157 ; n20158
g17723 and n20153_not n20158 ; n20159
g17724 nor pi0630 n19946 ; n20160
g17725 and n20159_not n20160 ; n20161
g17726 and pi0647 n20152_not ; n20162
g17727 and pi0647_not n20156 ; n20163
g17728 and pi1157 n20163_not ; n20164
g17729 and n20162_not n20164 ; n20165
g17730 and pi0630 n19950_not ; n20166
g17731 and n20165_not n20166 ; n20167
g17732 nor n20161 n20167 ; n20168
g17733 and pi0787 n20168_not ; n20169
g17734 nor pi0787 n20152 ; n20170
g17735 nor n20169 n20170 ; n20171
g17736 and pi0644 n20171_not ; n20172
g17737 and pi0715 n19954_not ; n20173
g17738 and n20172_not n20173 ; n20174
g17739 and n17804 n19892_not ; n20175
g17740 and n17804_not n20156 ; n20176
g17741 nor n20175 n20176 ; n20177
g17742 and pi0644 n20177_not ; n20178
g17743 nor pi0644 n19892 ; n20179
g17744 nor pi0715 n20179 ; n20180
g17745 and n20178_not n20180 ; n20181
g17746 and pi1160 n20181_not ; n20182
g17747 and n20174_not n20182 ; n20183
g17748 nor pi0644 n20171 ; n20184
g17749 and pi0644 n19953 ; n20185
g17750 nor pi0715 n20185 ; n20186
g17751 and n20184_not n20186 ; n20187
g17752 nor pi0644 n20177 ; n20188
g17753 and pi0644 n19892_not ; n20189
g17754 and pi0715 n20189_not ; n20190
g17755 and n20188_not n20190 ; n20191
g17756 nor pi1160 n20191 ; n20192
g17757 and n20187_not n20192 ; n20193
g17758 and pi0790 n20183_not ; n20194
g17759 and n20193_not n20194 ; n20195
g17760 and pi0790_not n20171 ; n20196
g17761 and n6305 n20196_not ; n20197
g17762 and n20195_not n20197 ; n20198
g17763 nor pi0144 n6305 ; n20199
g17764 nor pi0057 n20199 ; n20200
g17765 and n20198_not n20200 ; n20201
g17766 and pi0057 pi0144 ; n20202
g17767 nor pi0832 n20202 ; n20203
g17768 and n20201_not n20203 ; n20204
g17769 and n17803 n19341 ; n20205
g17770 and pi0787 n20205_not ; n20206
g17771 and pi0144 n2926_not ; n20207
g17772 and pi0736 n16645 ; n20208
g17773 nor n20207 n20208 ; n20209
g17774 and pi0778_not n20209 ; n20210
g17775 and pi0625 n20208 ; n20211
g17776 nor n20209 n20211 ; n20212
g17777 nor pi1153 n20212 ; n20213
g17778 and pi1153 n20207_not ; n20214
g17779 and n20211_not n20214 ; n20215
g17780 nor n20213 n20215 ; n20216
g17781 and pi0778 n20216_not ; n20217
g17782 nor n20210 n20217 ; n20218
g17783 and n19151 n20218 ; n20219
g17784 and pi0628_not n20219 ; n20220
g17785 and pi0629 n20220_not ; n20221
g17786 nor pi0609 pi1155 ; n20222
g17787 and pi0609 pi1155 ; n20223
g17788 and pi0785 n20222_not ; n20224
g17789 and n20223_not n20224 ; n20225
g17790 and pi0758 n17244 ; n20226
g17791 and n20225_not n20226 ; n20227
g17792 and pi0619_not pi1159 ; n20228
g17793 and pi0619 pi1159_not ; n20229
g17794 nor n20228 n20229 ; n20230
g17795 and pi0789 n20230_not ; n20231
g17796 nor pi0618 pi1154 ; n20232
g17797 and pi0618 pi1154 ; n20233
g17798 and pi0781 n20232_not ; n20234
g17799 and n20233_not n20234 ; n20235
g17800 nor n17117 n20231 ; n20236
g17801 and n20235_not n20236 ; n20237
g17802 and n20227 n20237 ; n20238
g17803 and n17969_not n20238 ; n20239
g17804 and pi0628 n20239_not ; n20240
g17805 nor n20221 n20240 ; n20241
g17806 nor pi1156 n20241 ; n20242
g17807 and pi0628 n20219 ; n20243
g17808 nor pi0628 n20239 ; n20244
g17809 and pi0629 n20244_not ; n20245
g17810 and pi1156 n20245_not ; n20246
g17811 and n20243_not n20246 ; n20247
g17812 nor n20242 n20247 ; n20248
g17813 nor n20207 n20248 ; n20249
g17814 and pi0792 n20249 ; n20250
g17815 and n16635 n20207_not ; n20251
g17816 and n17075_not n20218 ; n20252
g17817 and n16639_not n20252 ; n20253
g17818 nor n20207 n20253 ; n20254
g17819 nor n20251 n20254 ; n20255
g17820 and n17865 n20255 ; n20256
g17821 and pi0626_not n20238 ; n20257
g17822 nor n20207 n20257 ; n20258
g17823 nor pi1158 n20258 ; n20259
g17824 and pi0641 n20259_not ; n20260
g17825 and n20256_not n20260 ; n20261
g17826 and pi0626 n20238 ; n20262
g17827 nor n20207 n20262 ; n20263
g17828 and pi1158 n20263_not ; n20264
g17829 and n17866 n20255 ; n20265
g17830 nor pi0641 n20264 ; n20266
g17831 and n20265_not n20266 ; n20267
g17832 and pi0788 n20261_not ; n20268
g17833 and n20267_not n20268 ; n20269
g17834 and pi0618 n17117_not ; n20270
g17835 and n20227 n20270 ; n20271
g17836 and pi1154 n20207_not ; n20272
g17837 and n20271_not n20272 ; n20273
g17838 nor n20207 n20252 ; n20274
g17839 and pi0618 n20274_not ; n20275
g17840 and n17291 n20226 ; n20276
g17841 and pi1155 n20207_not ; n20277
g17842 and n20276_not n20277 ; n20278
g17843 and pi0609 n20218 ; n20279
g17844 nor n20207 n20226 ; n20280
g17845 and pi0736 n17469 ; n20281
g17846 and n20280 n20281_not ; n20282
g17847 and pi0625 n20281 ; n20283
g17848 nor n20282 n20283 ; n20284
g17849 nor pi1153 n20284 ; n20285
g17850 nor pi0608 n20215 ; n20286
g17851 and n20285_not n20286 ; n20287
g17852 and pi1153 n20280 ; n20288
g17853 and n20283_not n20288 ; n20289
g17854 and pi0608 n20213_not ; n20290
g17855 and n20289_not n20290 ; n20291
g17856 nor n20287 n20291 ; n20292
g17857 and pi0778 n20292_not ; n20293
g17858 nor pi0778 n20282 ; n20294
g17859 nor n20293 n20294 ; n20295
g17860 nor pi0609 n20295 ; n20296
g17861 nor pi1155 n20279 ; n20297
g17862 and n20296_not n20297 ; n20298
g17863 nor pi0660 n20278 ; n20299
g17864 and n20298_not n20299 ; n20300
g17865 and n17296 n20226 ; n20301
g17866 nor pi1155 n20207 ; n20302
g17867 and n20301_not n20302 ; n20303
g17868 and pi0609_not n20218 ; n20304
g17869 and pi0609 n20295_not ; n20305
g17870 and pi1155 n20304_not ; n20306
g17871 and n20305_not n20306 ; n20307
g17872 and pi0660 n20303_not ; n20308
g17873 and n20307_not n20308 ; n20309
g17874 nor n20300 n20309 ; n20310
g17875 and pi0785 n20310_not ; n20311
g17876 nor pi0785 n20295 ; n20312
g17877 nor n20311 n20312 ; n20313
g17878 nor pi0618 n20313 ; n20314
g17879 nor pi1154 n20275 ; n20315
g17880 and n20314_not n20315 ; n20316
g17881 nor pi0627 n20273 ; n20317
g17882 and n20316_not n20317 ; n20318
g17883 nor pi0618 n17117 ; n20319
g17884 and n20227 n20319 ; n20320
g17885 nor pi1154 n20207 ; n20321
g17886 and n20320_not n20321 ; n20322
g17887 nor pi0618 n20274 ; n20323
g17888 and pi0618 n20313_not ; n20324
g17889 and pi1154 n20323_not ; n20325
g17890 and n20324_not n20325 ; n20326
g17891 and pi0627 n20322_not ; n20327
g17892 and n20326_not n20327 ; n20328
g17893 nor n20318 n20328 ; n20329
g17894 and pi0781 n20329_not ; n20330
g17895 nor pi0781 n20313 ; n20331
g17896 nor n20330 n20331 ; n20332
g17897 and pi0789_not n20332 ; n20333
g17898 and n20227 n20235_not ; n20334
g17899 and pi0619 n17117_not ; n20335
g17900 and n20334 n20335 ; n20336
g17901 and pi1159 n20207_not ; n20337
g17902 and n20336_not n20337 ; n20338
g17903 and pi0619 n20254_not ; n20339
g17904 nor pi0619 n20332 ; n20340
g17905 nor pi1159 n20339 ; n20341
g17906 and n20340_not n20341 ; n20342
g17907 nor pi0648 n20338 ; n20343
g17908 and n20342_not n20343 ; n20344
g17909 nor pi0619 n17117 ; n20345
g17910 and n20334 n20345 ; n20346
g17911 nor pi1159 n20207 ; n20347
g17912 and n20346_not n20347 ; n20348
g17913 nor pi0619 n20254 ; n20349
g17914 and pi0619 n20332_not ; n20350
g17915 and pi1159 n20349_not ; n20351
g17916 and n20350_not n20351 ; n20352
g17917 and pi0648 n20348_not ; n20353
g17918 and n20352_not n20353 ; n20354
g17919 and pi0789 n20344_not ; n20355
g17920 and n20354_not n20355 ; n20356
g17921 and n17970 n20333_not ; n20357
g17922 and n20356_not n20357 ; n20358
g17923 nor n20269 n20358 ; n20359
g17924 nor n20250 n20359 ; n20360
g17925 and pi0629 n19139 ; n20361
g17926 and pi0629_not n19140 ; n20362
g17927 and pi0792 n20361_not ; n20363
g17928 and n20362_not n20363 ; n20364
g17929 and n20249_not n20364 ; n20365
g17930 nor n20206 n20365 ; n20366
g17931 and n20360_not n20366 ; n20367
g17932 and n17779_not n20239 ; n20368
g17933 and pi0630_not n20368 ; n20369
g17934 and pi0647 n20369_not ; n20370
g17935 and n19142_not n20219 ; n20371
g17936 and pi0630 n20371_not ; n20372
g17937 nor n20370 n20372 ; n20373
g17938 nor pi1157 n20373 ; n20374
g17939 and pi0630 n20368 ; n20375
g17940 nor pi0630 n20371 ; n20376
g17941 and pi0647 n20376_not ; n20377
g17942 and pi1157 n20375_not ; n20378
g17943 and n20377_not n20378 ; n20379
g17944 nor n20374 n20379 ; n20380
g17945 and pi0787 n20207_not ; n20381
g17946 and n20380_not n20381 ; n20382
g17947 nor n20367 n20382 ; n20383
g17948 and pi0790_not n20383 ; n20384
g17949 and n17804_not n20368 ; n20385
g17950 and pi0644 n20385 ; n20386
g17951 nor pi0715 n20207 ; n20387
g17952 and n20386_not n20387 ; n20388
g17953 and n19342_not n20371 ; n20389
g17954 nor n20207 n20389 ; n20390
g17955 nor pi0644 n20390 ; n20391
g17956 and pi0644 n20383 ; n20392
g17957 and pi0715 n20391_not ; n20393
g17958 and n20392_not n20393 ; n20394
g17959 and pi1160 n20388_not ; n20395
g17960 and n20394_not n20395 ; n20396
g17961 and pi0644_not n20385 ; n20397
g17962 and pi0715 n20207_not ; n20398
g17963 and n20397_not n20398 ; n20399
g17964 and pi0644_not n20383 ; n20400
g17965 and pi0644 n20390_not ; n20401
g17966 nor pi0715 n20401 ; n20402
g17967 and n20400_not n20402 ; n20403
g17968 nor pi1160 n20399 ; n20404
g17969 and n20403_not n20404 ; n20405
g17970 nor n20396 n20405 ; n20406
g17971 and pi0790 n20406_not ; n20407
g17972 and pi0832 n20384_not ; n20408
g17973 and n20407_not n20408 ; n20409
g17974 nor n20204 n20409 ; po0301
g17975 and pi0145_not po1038 ; n20411
g17976 nor pi0145 n17059 ; n20412
g17977 and n16635 n20412_not ; n20413
g17978 and pi0698_not n2571 ; n20414
g17979 and n20412 n20414_not ; n20415
g17980 nor pi0145 n16641 ; n20416
g17981 and n16647 n20416_not ; n20417
g17982 and pi0145 n18076_not ; n20418
g17983 nor pi0038 n20418 ; n20419
g17984 and n2571 n20419_not ; n20420
g17985 and pi0145_not n18072 ; n20421
g17986 nor n20420 n20421 ; n20422
g17987 nor pi0698 n20417 ; n20423
g17988 and n20422_not n20423 ; n20424
g17989 nor n20415 n20424 ; n20425
g17990 and pi0778_not n20425 ; n20426
g17991 and pi0625_not n20412 ; n20427
g17992 and pi0625 n20425_not ; n20428
g17993 and pi1153 n20427_not ; n20429
g17994 and n20428_not n20429 ; n20430
g17995 and pi0625 n20412 ; n20431
g17996 nor pi0625 n20425 ; n20432
g17997 nor pi1153 n20431 ; n20433
g17998 and n20432_not n20433 ; n20434
g17999 nor n20430 n20434 ; n20435
g18000 and pi0778 n20435_not ; n20436
g18001 nor n20426 n20436 ; n20437
g18002 nor n17075 n20437 ; n20438
g18003 and n17075 n20412_not ; n20439
g18004 nor n20438 n20439 ; n20440
g18005 and n16639_not n20440 ; n20441
g18006 and n16639 n20412 ; n20442
g18007 nor n20441 n20442 ; n20443
g18008 and n16635_not n20443 ; n20444
g18009 nor n20413 n20444 ; n20445
g18010 and n16631_not n20445 ; n20446
g18011 and n16631 n20412 ; n20447
g18012 nor n20446 n20447 ; n20448
g18013 and pi0792_not n20448 ; n20449
g18014 and pi0628 n20448_not ; n20450
g18015 and pi0628_not n20412 ; n20451
g18016 and pi1156 n20451_not ; n20452
g18017 and n20450_not n20452 ; n20453
g18018 and pi0628 n20412 ; n20454
g18019 nor pi0628 n20448 ; n20455
g18020 nor pi1156 n20454 ; n20456
g18021 and n20455_not n20456 ; n20457
g18022 nor n20453 n20457 ; n20458
g18023 and pi0792 n20458_not ; n20459
g18024 nor n20449 n20459 ; n20460
g18025 nor pi0647 n20460 ; n20461
g18026 and pi0647 n20412_not ; n20462
g18027 nor n20461 n20462 ; n20463
g18028 and pi1157_not n20463 ; n20464
g18029 and pi0647 n20460_not ; n20465
g18030 nor pi0647 n20412 ; n20466
g18031 nor n20465 n20466 ; n20467
g18032 and pi1157 n20467 ; n20468
g18033 nor n20464 n20468 ; n20469
g18034 and pi0787 n20469_not ; n20470
g18035 and pi0787_not n20460 ; n20471
g18036 nor n20470 n20471 ; n20472
g18037 nor pi0644 n20472 ; n20473
g18038 and pi0715 n20473_not ; n20474
g18039 and pi0145 n2571_not ; n20475
g18040 and pi0145 n17275_not ; n20476
g18041 nor pi0145 n17048 ; n20477
g18042 and pi0767 n20477_not ; n20478
g18043 nor pi0145 pi0767 ; n20479
g18044 and n17221 n20479 ; n20480
g18045 nor n20476 n20480 ; n20481
g18046 and n20478_not n20481 ; n20482
g18047 nor pi0038 n20482 ; n20483
g18048 and pi0767_not n17280 ; n20484
g18049 and pi0038 n20416_not ; n20485
g18050 and n20484_not n20485 ; n20486
g18051 nor n20483 n20486 ; n20487
g18052 and n2571 n20487_not ; n20488
g18053 nor n20475 n20488 ; n20489
g18054 nor n17117 n20489 ; n20490
g18055 and n17117 n20412_not ; n20491
g18056 nor n20490 n20491 ; n20492
g18057 nor pi0785 n20492 ; n20493
g18058 nor n17291 n20412 ; n20494
g18059 and pi0609 n20490 ; n20495
g18060 nor n20494 n20495 ; n20496
g18061 and pi1155 n20496_not ; n20497
g18062 nor n17296 n20412 ; n20498
g18063 and pi0609_not n20490 ; n20499
g18064 nor n20498 n20499 ; n20500
g18065 nor pi1155 n20500 ; n20501
g18066 nor n20497 n20501 ; n20502
g18067 and pi0785 n20502_not ; n20503
g18068 nor n20493 n20503 ; n20504
g18069 nor pi0781 n20504 ; n20505
g18070 and pi0618_not n20412 ; n20506
g18071 and pi0618 n20504 ; n20507
g18072 and pi1154 n20506_not ; n20508
g18073 and n20507_not n20508 ; n20509
g18074 and pi0618_not n20504 ; n20510
g18075 and pi0618 n20412 ; n20511
g18076 nor pi1154 n20511 ; n20512
g18077 and n20510_not n20512 ; n20513
g18078 nor n20509 n20513 ; n20514
g18079 and pi0781 n20514_not ; n20515
g18080 nor n20505 n20515 ; n20516
g18081 nor pi0789 n20516 ; n20517
g18082 and pi0619_not n20412 ; n20518
g18083 and pi0619 n20516 ; n20519
g18084 and pi1159 n20518_not ; n20520
g18085 and n20519_not n20520 ; n20521
g18086 and pi0619_not n20516 ; n20522
g18087 and pi0619 n20412 ; n20523
g18088 nor pi1159 n20523 ; n20524
g18089 and n20522_not n20524 ; n20525
g18090 nor n20521 n20525 ; n20526
g18091 and pi0789 n20526_not ; n20527
g18092 nor n20517 n20527 ; n20528
g18093 nor pi0788 n20528 ; n20529
g18094 and pi0626_not n20412 ; n20530
g18095 and pi0626 n20528 ; n20531
g18096 and pi1158 n20530_not ; n20532
g18097 and n20531_not n20532 ; n20533
g18098 and pi0626_not n20528 ; n20534
g18099 and pi0626 n20412 ; n20535
g18100 nor pi1158 n20535 ; n20536
g18101 and n20534_not n20536 ; n20537
g18102 nor n20533 n20537 ; n20538
g18103 and pi0788 n20538_not ; n20539
g18104 nor n20529 n20539 ; n20540
g18105 and n17779_not n20540 ; n20541
g18106 and n17779 n20412 ; n20542
g18107 nor n20541 n20542 ; n20543
g18108 nor n17804 n20543 ; n20544
g18109 and n17804 n20412 ; n20545
g18110 nor n20544 n20545 ; n20546
g18111 and pi0644 n20546_not ; n20547
g18112 and pi0644_not n20412 ; n20548
g18113 nor pi0715 n20548 ; n20549
g18114 and n20547_not n20549 ; n20550
g18115 and pi1160 n20550_not ; n20551
g18116 and n20474_not n20551 ; n20552
g18117 and pi0644 n20472_not ; n20553
g18118 and n17802 n20463_not ; n20554
g18119 and pi0630 pi0647_not ; n20555
g18120 and pi1157 n20555 ; n20556
g18121 and pi0630_not pi0647 ; n20557
g18122 and pi1157_not n20557 ; n20558
g18123 nor n20556 n20558 ; n20559
g18124 and n20543 n20559_not ; n20560
g18125 and n17801 n20467_not ; n20561
g18126 nor n20554 n20561 ; n20562
g18127 and n20560_not n20562 ; n20563
g18128 and pi0787 n20563_not ; n20564
g18129 and pi0629_not n20453 ; n20565
g18130 and pi0628_not pi0629 ; n20566
g18131 and pi1156 n20566 ; n20567
g18132 and pi0628 pi0629_not ; n20568
g18133 and pi1156_not n20568 ; n20569
g18134 nor n20567 n20569 ; n20570
g18135 nor n20540 n20570 ; n20571
g18136 and pi0629 n20457 ; n20572
g18137 nor n20565 n20572 ; n20573
g18138 and n20571_not n20573 ; n20574
g18139 and pi0792 n20574_not ; n20575
g18140 and pi0609 n20437 ; n20576
g18141 and pi0145 n17625_not ; n20577
g18142 nor pi0145 n17612 ; n20578
g18143 and pi0767 n20577_not ; n20579
g18144 and n20578_not n20579 ; n20580
g18145 and pi0145_not n17629 ; n20581
g18146 and pi0145 n17631 ; n20582
g18147 nor pi0767 n20582 ; n20583
g18148 and n20581_not n20583 ; n20584
g18149 nor n20580 n20584 ; n20585
g18150 nor pi0039 n20585 ; n20586
g18151 and pi0145 n17605 ; n20587
g18152 nor pi0145 n17546 ; n20588
g18153 nor pi0767 n20588 ; n20589
g18154 and n20587_not n20589 ; n20590
g18155 and pi0145_not n17404 ; n20591
g18156 and pi0145 n17485 ; n20592
g18157 and pi0767 n20592_not ; n20593
g18158 and n20591_not n20593 ; n20594
g18159 and pi0039 n20590_not ; n20595
g18160 and n20594_not n20595 ; n20596
g18161 nor pi0038 n20586 ; n20597
g18162 and n20596_not n20597 ; n20598
g18163 nor pi0767 n17490 ; n20599
g18164 and n19471 n20599_not ; n20600
g18165 nor pi0145 n20600 ; n20601
g18166 and pi0767_not n17244 ; n20602
g18167 nor n17469 n20602 ; n20603
g18168 and pi0145 n20603_not ; n20604
g18169 and n6284 n20604 ; n20605
g18170 and pi0038 n20605_not ; n20606
g18171 and n20601_not n20606 ; n20607
g18172 nor pi0698 n20607 ; n20608
g18173 and n20598_not n20608 ; n20609
g18174 and pi0698 n20487 ; n20610
g18175 and n2571 n20609_not ; n20611
g18176 and n20610_not n20611 ; n20612
g18177 nor n20475 n20612 ; n20613
g18178 and pi0625_not n20613 ; n20614
g18179 and pi0625 n20489 ; n20615
g18180 nor pi1153 n20615 ; n20616
g18181 and n20614_not n20616 ; n20617
g18182 nor pi0608 n20430 ; n20618
g18183 and n20617_not n20618 ; n20619
g18184 and pi0625_not n20489 ; n20620
g18185 and pi0625 n20613 ; n20621
g18186 and pi1153 n20620_not ; n20622
g18187 and n20621_not n20622 ; n20623
g18188 and pi0608 n20434_not ; n20624
g18189 and n20623_not n20624 ; n20625
g18190 nor n20619 n20625 ; n20626
g18191 and pi0778 n20626_not ; n20627
g18192 and pi0778_not n20613 ; n20628
g18193 nor n20627 n20628 ; n20629
g18194 nor pi0609 n20629 ; n20630
g18195 nor pi1155 n20576 ; n20631
g18196 and n20630_not n20631 ; n20632
g18197 nor pi0660 n20497 ; n20633
g18198 and n20632_not n20633 ; n20634
g18199 and pi0609_not n20437 ; n20635
g18200 and pi0609 n20629_not ; n20636
g18201 and pi1155 n20635_not ; n20637
g18202 and n20636_not n20637 ; n20638
g18203 and pi0660 n20501_not ; n20639
g18204 and n20638_not n20639 ; n20640
g18205 nor n20634 n20640 ; n20641
g18206 and pi0785 n20641_not ; n20642
g18207 nor pi0785 n20629 ; n20643
g18208 nor n20642 n20643 ; n20644
g18209 nor pi0618 n20644 ; n20645
g18210 and pi0618 n20440 ; n20646
g18211 nor pi1154 n20646 ; n20647
g18212 and n20645_not n20647 ; n20648
g18213 nor pi0627 n20509 ; n20649
g18214 and n20648_not n20649 ; n20650
g18215 and pi0618_not n20440 ; n20651
g18216 and pi0618 n20644_not ; n20652
g18217 and pi1154 n20651_not ; n20653
g18218 and n20652_not n20653 ; n20654
g18219 and pi0627 n20513_not ; n20655
g18220 and n20654_not n20655 ; n20656
g18221 nor n20650 n20656 ; n20657
g18222 and pi0781 n20657_not ; n20658
g18223 nor pi0781 n20644 ; n20659
g18224 nor n20658 n20659 ; n20660
g18225 and pi0789_not n20660 ; n20661
g18226 and pi0619 n20443_not ; n20662
g18227 nor pi0619 n20660 ; n20663
g18228 nor pi1159 n20662 ; n20664
g18229 and n20663_not n20664 ; n20665
g18230 nor pi0648 n20521 ; n20666
g18231 and n20665_not n20666 ; n20667
g18232 and pi0619 n20660_not ; n20668
g18233 nor pi0619 n20443 ; n20669
g18234 and pi1159 n20669_not ; n20670
g18235 and n20668_not n20670 ; n20671
g18236 and pi0648 n20525_not ; n20672
g18237 and n20671_not n20672 ; n20673
g18238 and pi0789 n20667_not ; n20674
g18239 and n20673_not n20674 ; n20675
g18240 and n17970 n20661_not ; n20676
g18241 and n20675_not n20676 ; n20677
g18242 and n17871 n20445 ; n20678
g18243 and n16630_not n20538 ; n20679
g18244 nor n20678 n20679 ; n20680
g18245 and pi0788 n20680_not ; n20681
g18246 nor n20364 n20681 ; n20682
g18247 and n20677_not n20682 ; n20683
g18248 nor n20575 n20683 ; n20684
g18249 nor n20206 n20684 ; n20685
g18250 nor n20564 n20685 ; n20686
g18251 and pi0644_not n20686 ; n20687
g18252 nor pi0715 n20553 ; n20688
g18253 and n20687_not n20688 ; n20689
g18254 and pi0644 n20412 ; n20690
g18255 nor pi0644 n20546 ; n20691
g18256 and pi0715 n20690_not ; n20692
g18257 and n20691_not n20692 ; n20693
g18258 nor pi1160 n20693 ; n20694
g18259 and n20689_not n20694 ; n20695
g18260 nor n20552 n20695 ; n20696
g18261 and pi0790 n20696_not ; n20697
g18262 and pi0644 n20551 ; n20698
g18263 and pi0790 n20698_not ; n20699
g18264 and n20686 n20699_not ; n20700
g18265 nor n20697 n20700 ; n20701
g18266 nor po1038 n20701 ; n20702
g18267 nor pi0832 n20411 ; n20703
g18268 and n20702_not n20703 ; n20704
g18269 nor pi0145 n2926 ; n20705
g18270 and pi0698_not n16645 ; n20706
g18271 nor n20705 n20706 ; n20707
g18272 and pi0778_not n20707 ; n20708
g18273 and pi0625_not n20706 ; n20709
g18274 nor n20707 n20709 ; n20710
g18275 and pi1153 n20710_not ; n20711
g18276 nor pi1153 n20705 ; n20712
g18277 and n20709_not n20712 ; n20713
g18278 nor n20711 n20713 ; n20714
g18279 and pi0778 n20714_not ; n20715
g18280 nor n20708 n20715 ; n20716
g18281 and n17845_not n20716 ; n20717
g18282 and n17847_not n20717 ; n20718
g18283 and n17849_not n20718 ; n20719
g18284 and n17851_not n20719 ; n20720
g18285 and n17857_not n20720 ; n20721
g18286 and pi0647_not n20721 ; n20722
g18287 and pi0647 n20705 ; n20723
g18288 nor pi1157 n20723 ; n20724
g18289 and n20722_not n20724 ; n20725
g18290 and pi0630 n20725 ; n20726
g18291 nor n20602 n20705 ; n20727
g18292 nor n17874 n20727 ; n20728
g18293 nor pi0785 n20728 ; n20729
g18294 nor n17879 n20727 ; n20730
g18295 and pi1155 n20730_not ; n20731
g18296 and n17882_not n20728 ; n20732
g18297 nor pi1155 n20732 ; n20733
g18298 nor n20731 n20733 ; n20734
g18299 and pi0785 n20734_not ; n20735
g18300 nor n20729 n20735 ; n20736
g18301 nor pi0781 n20736 ; n20737
g18302 and n17889_not n20736 ; n20738
g18303 and pi1154 n20738_not ; n20739
g18304 and n17892_not n20736 ; n20740
g18305 nor pi1154 n20740 ; n20741
g18306 nor n20739 n20741 ; n20742
g18307 and pi0781 n20742_not ; n20743
g18308 nor n20737 n20743 ; n20744
g18309 nor pi0789 n20744 ; n20745
g18310 and pi0619_not n20705 ; n20746
g18311 and pi0619 n20744 ; n20747
g18312 and pi1159 n20746_not ; n20748
g18313 and n20747_not n20748 ; n20749
g18314 and pi0619_not n20744 ; n20750
g18315 and pi0619 n20705 ; n20751
g18316 nor pi1159 n20751 ; n20752
g18317 and n20750_not n20752 ; n20753
g18318 nor n20749 n20753 ; n20754
g18319 and pi0789 n20754_not ; n20755
g18320 nor n20745 n20755 ; n20756
g18321 nor pi0788 n20756 ; n20757
g18322 and pi0626_not n20705 ; n20758
g18323 and pi0626 n20756 ; n20759
g18324 and pi1158 n20758_not ; n20760
g18325 and n20759_not n20760 ; n20761
g18326 and pi0626_not n20756 ; n20762
g18327 and pi0626 n20705 ; n20763
g18328 nor pi1158 n20763 ; n20764
g18329 and n20762_not n20764 ; n20765
g18330 nor n20761 n20765 ; n20766
g18331 and pi0788 n20766_not ; n20767
g18332 nor n20757 n20767 ; n20768
g18333 and n17779_not n20768 ; n20769
g18334 and n17779 n20705 ; n20770
g18335 nor n20769 n20770 ; n20771
g18336 and n20559_not n20771 ; n20772
g18337 and pi0647 n20721_not ; n20773
g18338 nor pi0647 n20705 ; n20774
g18339 nor n20773 n20774 ; n20775
g18340 and n17801 n20775_not ; n20776
g18341 nor n20726 n20776 ; n20777
g18342 and n20772_not n20777 ; n20778
g18343 and pi0787 n20778_not ; n20779
g18344 and n17871 n20719 ; n20780
g18345 and n16630_not n20766 ; n20781
g18346 nor n20780 n20781 ; n20782
g18347 and pi0788 n20782_not ; n20783
g18348 and pi0618 n20717 ; n20784
g18349 and pi0609 n20716 ; n20785
g18350 nor n17168 n20707 ; n20786
g18351 and pi0625 n20786 ; n20787
g18352 and n20727 n20786_not ; n20788
g18353 nor n20787 n20788 ; n20789
g18354 and n20712 n20789_not ; n20790
g18355 nor pi0608 n20711 ; n20791
g18356 and n20790_not n20791 ; n20792
g18357 and pi1153 n20727 ; n20793
g18358 and n20787_not n20793 ; n20794
g18359 and pi0608 n20713_not ; n20795
g18360 and n20794_not n20795 ; n20796
g18361 nor n20792 n20796 ; n20797
g18362 and pi0778 n20797_not ; n20798
g18363 nor pi0778 n20788 ; n20799
g18364 nor n20798 n20799 ; n20800
g18365 nor pi0609 n20800 ; n20801
g18366 nor pi1155 n20785 ; n20802
g18367 and n20801_not n20802 ; n20803
g18368 nor pi0660 n20731 ; n20804
g18369 and n20803_not n20804 ; n20805
g18370 and pi0609_not n20716 ; n20806
g18371 and pi0609 n20800_not ; n20807
g18372 and pi1155 n20806_not ; n20808
g18373 and n20807_not n20808 ; n20809
g18374 and pi0660 n20733_not ; n20810
g18375 and n20809_not n20810 ; n20811
g18376 nor n20805 n20811 ; n20812
g18377 and pi0785 n20812_not ; n20813
g18378 nor pi0785 n20800 ; n20814
g18379 nor n20813 n20814 ; n20815
g18380 nor pi0618 n20815 ; n20816
g18381 nor pi1154 n20784 ; n20817
g18382 and n20816_not n20817 ; n20818
g18383 nor pi0627 n20739 ; n20819
g18384 and n20818_not n20819 ; n20820
g18385 and pi0618_not n20717 ; n20821
g18386 and pi0618 n20815_not ; n20822
g18387 and pi1154 n20821_not ; n20823
g18388 and n20822_not n20823 ; n20824
g18389 and pi0627 n20741_not ; n20825
g18390 and n20824_not n20825 ; n20826
g18391 nor n20820 n20826 ; n20827
g18392 and pi0781 n20827_not ; n20828
g18393 nor pi0781 n20815 ; n20829
g18394 nor n20828 n20829 ; n20830
g18395 and pi0789_not n20830 ; n20831
g18396 nor pi0619 n20830 ; n20832
g18397 and pi0619 n20718 ; n20833
g18398 nor pi1159 n20833 ; n20834
g18399 and n20832_not n20834 ; n20835
g18400 nor pi0648 n20749 ; n20836
g18401 and n20835_not n20836 ; n20837
g18402 and pi0619_not n20718 ; n20838
g18403 and pi0619 n20830_not ; n20839
g18404 and pi1159 n20838_not ; n20840
g18405 and n20839_not n20840 ; n20841
g18406 and pi0648 n20753_not ; n20842
g18407 and n20841_not n20842 ; n20843
g18408 and pi0789 n20837_not ; n20844
g18409 and n20843_not n20844 ; n20845
g18410 and n17970 n20831_not ; n20846
g18411 and n20845_not n20846 ; n20847
g18412 nor n20783 n20847 ; n20848
g18413 nor n20364 n20848 ; n20849
g18414 and n17854 n20768 ; n20850
g18415 and pi1156 n17862_not ; n20851
g18416 and n20720 n20851 ; n20852
g18417 nor n20850 n20852 ; n20853
g18418 nor pi0629 n20853 ; n20854
g18419 nor pi1156 n17997 ; n20855
g18420 and n20720 n20855 ; n20856
g18421 and n17853 n20768 ; n20857
g18422 nor n20856 n20857 ; n20858
g18423 and pi0629 n20858_not ; n20859
g18424 nor n20854 n20859 ; n20860
g18425 and pi0792 n20860_not ; n20861
g18426 nor n20206 n20861 ; n20862
g18427 and n20849_not n20862 ; n20863
g18428 nor n20779 n20863 ; n20864
g18429 and pi0790_not n20864 ; n20865
g18430 nor pi0787 n20721 ; n20866
g18431 and pi1157 n20775_not ; n20867
g18432 nor n20725 n20867 ; n20868
g18433 and pi0787 n20868_not ; n20869
g18434 nor n20866 n20869 ; n20870
g18435 and pi0644_not n20870 ; n20871
g18436 and pi0644 n20864 ; n20872
g18437 and pi0715 n20871_not ; n20873
g18438 and n20872_not n20873 ; n20874
g18439 nor n17804 n20771 ; n20875
g18440 and n17804 n20705 ; n20876
g18441 nor n20875 n20876 ; n20877
g18442 and pi0644 n20877_not ; n20878
g18443 and pi0644_not n20705 ; n20879
g18444 nor pi0715 n20879 ; n20880
g18445 and n20878_not n20880 ; n20881
g18446 and pi1160 n20881_not ; n20882
g18447 and n20874_not n20882 ; n20883
g18448 nor pi0644 n20877 ; n20884
g18449 and pi0644 n20705 ; n20885
g18450 and pi0715 n20885_not ; n20886
g18451 and n20884_not n20886 ; n20887
g18452 and pi0644 n20870 ; n20888
g18453 and pi0644_not n20864 ; n20889
g18454 nor pi0715 n20888 ; n20890
g18455 and n20889_not n20890 ; n20891
g18456 nor pi1160 n20887 ; n20892
g18457 and n20891_not n20892 ; n20893
g18458 nor n20883 n20893 ; n20894
g18459 and pi0790 n20894_not ; n20895
g18460 and pi0832 n20865_not ; n20896
g18461 and n20895_not n20896 ; n20897
g18462 nor n20704 n20897 ; po0302
g18463 nor pi0146 n10197 ; n20899
g18464 nor pi0146 n16641 ; n20900
g18465 and pi0743 pi0947 ; n20901
g18466 and pi0907 pi0947_not ; n20902
g18467 and pi0735 n20902 ; n20903
g18468 nor n20901 n20903 ; n20904
g18469 and n2926 n20904 ; n20905
g18470 and n6284 n20905 ; n20906
g18471 and pi0038 n20906_not ; n20907
g18472 and n20900_not n20907 ; n20908
g18473 nor pi0146 n16941 ; n20909
g18474 and n16941 n20904 ; n20910
g18475 and pi0299 n20909_not ; n20911
g18476 and n20910_not n20911 ; n20912
g18477 nor pi0146 n16930 ; n20913
g18478 and n16930 n20904 ; n20914
g18479 nor pi0299 n20913 ; n20915
g18480 and n20914_not n20915 ; n20916
g18481 nor pi0039 n20912 ; n20917
g18482 and n20916_not n20917 ; n20918
g18483 and n16653 n20904_not ; n20919
g18484 and pi0146 n16653_not ; n20920
g18485 nor n20919 n20920 ; n20921
g18486 and n3448 n20921_not ; n20922
g18487 and pi0907_not n6241 ; n20923
g18488 and pi0146 n17018_not ; n20924
g18489 and n20923_not n20924 ; n20925
g18490 and pi0735 pi0907 ; n20926
g18491 and n17018 n20926 ; n20927
g18492 and pi0146 n17011_not ; n20928
g18493 and n20923 n20928 ; n20929
g18494 nor pi0947 n20927 ; n20930
g18495 and n20929_not n20930 ; n20931
g18496 and pi0743 n17018 ; n20932
g18497 and pi0947 n20924_not ; n20933
g18498 and n20932_not n20933 ; n20934
g18499 nor n20931 n20934 ; n20935
g18500 nor n20925 n20935 ; n20936
g18501 nor n3448 n20936 ; n20937
g18502 nor pi0215 n20922 ; n20938
g18503 and n20937_not n20938 ; n20939
g18504 and n16970 n20904_not ; n20940
g18505 and pi0146 n17042 ; n20941
g18506 and pi0215 n20940_not ; n20942
g18507 and n20941_not n20942 ; n20943
g18508 nor n20939 n20943 ; n20944
g18509 and pi0299 n20944_not ; n20945
g18510 and pi0146 n16970_not ; n20946
g18511 nor n20940 n20946 ; n20947
g18512 nor n6205 n20947 ; n20948
g18513 nor pi0146 n16990 ; n20949
g18514 and n16990 n20904 ; n20950
g18515 and n6205 n20949_not ; n20951
g18516 and n20950_not n20951 ; n20952
g18517 nor n20948 n20952 ; n20953
g18518 and pi0223 n20953_not ; n20954
g18519 and n2603 n20921 ; n20955
g18520 and n17018 n20904_not ; n20956
g18521 nor n6205 n20924 ; n20957
g18522 and n20956_not n20957 ; n20958
g18523 and n17011 n20904_not ; n20959
g18524 and n6205 n20928_not ; n20960
g18525 and n20959_not n20960 ; n20961
g18526 nor n20958 n20961 ; n20962
g18527 nor n2603 n20962 ; n20963
g18528 nor pi0223 n20955 ; n20964
g18529 and n20963_not n20964 ; n20965
g18530 nor pi0299 n20954 ; n20966
g18531 and n20965_not n20966 ; n20967
g18532 nor n20945 n20967 ; n20968
g18533 and pi0039 n20968_not ; n20969
g18534 nor pi0038 n20918 ; n20970
g18535 and n20969_not n20970 ; n20971
g18536 and n10197 n20908_not ; n20972
g18537 and n20971_not n20972 ; n20973
g18538 nor pi0832 n20899 ; n20974
g18539 and n20973_not n20974 ; n20975
g18540 nor pi0146 n2926 ; n20976
g18541 and pi0832 n20976_not ; n20977
g18542 and n20905_not n20977 ; n20978
g18543 or n20975 n20978 ; po0303
g18544 nor pi0147 n2926 ; n20980
g18545 and pi0770_not pi0947 ; n20981
g18546 and pi0726 n20902 ; n20982
g18547 nor n20981 n20982 ; n20983
g18548 and n2926 n20983_not ; n20984
g18549 and pi0832 n20980_not ; n20985
g18550 and n20984_not n20985 ; n20986
g18551 nor pi0147 n10197 ; n20987
g18552 and pi0947_not n16958 ; n20988
g18553 nor pi0039 n20988 ; n20989
g18554 and pi0299_not n17024 ; n20990
g18555 and pi0947 n20990 ; n20991
g18556 and pi0947_not n17026 ; n20992
g18557 and n17018 n20902 ; n20993
g18558 nor n17030 n20993 ; n20994
g18559 nor n3448 n20994 ; n20995
g18560 nor pi0215 n20995 ; n20996
g18561 and n20992_not n20996 ; n20997
g18562 and pi0215 n17041_not ; n20998
g18563 and n16970 n20902 ; n20999
g18564 and n20998 n20999_not ; n21000
g18565 nor n20997 n21000 ; n21001
g18566 and pi0299 n21001_not ; n21002
g18567 nor n17025 n21002 ; n21003
g18568 and n20991_not n21003 ; n21004
g18569 and pi0039 n21004_not ; n21005
g18570 nor n20989 n21005 ; n21006
g18571 and pi0038_not n21006 ; n21007
g18572 and pi0038 pi0947_not ; n21008
g18573 and n17050 n21008 ; n21009
g18574 nor n21007 n21009 ; n21010
g18575 and pi0770_not n21010 ; n21011
g18576 and pi0770 n17052_not ; n21012
g18577 nor n21011 n21012 ; n21013
g18578 nor pi0147 n21013 ; n21014
g18579 nor n17051 n21009 ; n21015
g18580 and pi0947 n16958 ; n21016
g18581 nor pi0039 n21016 ; n21017
g18582 and pi0947 n17024 ; n21018
g18583 nor pi0299 n21018 ; n21019
g18584 and pi0215 pi0947 ; n21020
g18585 and n16970 n21020 ; n21021
g18586 and pi0299 n21021_not ; n21022
g18587 and pi0947 n17018 ; n21023
g18588 nor n3448 n21023 ; n21024
g18589 and pi0947 n16653 ; n21025
g18590 and n3448 n21025_not ; n21026
g18591 nor pi0215 n21026 ; n21027
g18592 and n21024_not n21027 ; n21028
g18593 and n21022 n21028_not ; n21029
g18594 nor n21019 n21029 ; n21030
g18595 and pi0039 n21030_not ; n21031
g18596 nor n21017 n21031 ; n21032
g18597 nor pi0038 n21032 ; n21033
g18598 and n21015 n21033_not ; n21034
g18599 and pi0147 pi0770_not ; n21035
g18600 and n21034 n21035 ; n21036
g18601 nor pi0726 n21036 ; n21037
g18602 and n21014_not n21037 ; n21038
g18603 and n6236 n17050 ; n21039
g18604 nor pi0147 n21039 ; n21040
g18605 and n6236_not n16641 ; n21041
g18606 and pi0038 n21041_not ; n21042
g18607 and n21040_not n21042 ; n21043
g18608 and pi0299 pi0947 ; n21044
g18609 and n17026 n20902_not ; n21045
g18610 nor n17030 n21023 ; n21046
g18611 nor n3448 n21046 ; n21047
g18612 nor pi0215 n21047 ; n21048
g18613 and n21045_not n21048 ; n21049
g18614 nor n20998 n21049 ; n21050
g18615 and pi0299 n21050_not ; n21051
g18616 and pi0947_not n16992 ; n21052
g18617 and pi0223 n21052_not ; n21053
g18618 and n16992 n20902_not ; n21054
g18619 and pi0223 n21054_not ; n21055
g18620 and n2521 n16654 ; n21056
g18621 nor n17021 n21056 ; n21057
g18622 and n6236 n21057_not ; n21058
g18623 nor pi0223 n21058 ; n21059
g18624 nor n21053 n21055 ; n21060
g18625 and n21059_not n21060 ; n21061
g18626 nor pi0299 n21061 ; n21062
g18627 nor n21044 n21051 ; n21063
g18628 and n21062_not n21063 ; n21064
g18629 and pi0039 n21064 ; n21065
g18630 and n6236_not n16958 ; n21066
g18631 nor pi0039 n21066 ; n21067
g18632 and n16958 n21067 ; n21068
g18633 nor n21065 n21068 ; n21069
g18634 and pi0147_not n21069 ; n21070
g18635 and n6236_not n17024 ; n21071
g18636 and pi0299_not n21071 ; n21072
g18637 and pi0215 n17037_not ; n21073
g18638 and n6236_not n16653 ; n21074
g18639 and n3448 n21074 ; n21075
g18640 nor pi0215 n21075 ; n21076
g18641 and n17033_not n21076 ; n21077
g18642 and pi0299 n21073_not ; n21078
g18643 and n21077_not n21078 ; n21079
g18644 nor n21072 n21079 ; n21080
g18645 and pi0039 n21080 ; n21081
g18646 nor n21067 n21081 ; n21082
g18647 and pi0147 n21082 ; n21083
g18648 nor pi0038 n21083 ; n21084
g18649 and n21070_not n21084 ; n21085
g18650 nor pi0770 n21043 ; n21086
g18651 and n21085_not n21086 ; n21087
g18652 nor pi0147 n16641 ; n21088
g18653 and n16641 n20902 ; n21089
g18654 and pi0038 n21089_not ; n21090
g18655 and n21088_not n21090 ; n21091
g18656 nor n21021 n21050 ; n21092
g18657 and pi0299 n21092_not ; n21093
g18658 and n20902_not n20990 ; n21094
g18659 nor n21093 n21094 ; n21095
g18660 and pi0039 n21095_not ; n21096
g18661 and n16958 n20902_not ; n21097
g18662 and pi0039_not n21097 ; n21098
g18663 nor n21096 n21098 ; n21099
g18664 and pi0147_not n21099 ; n21100
g18665 and pi0215 n20999_not ; n21101
g18666 nor n3448 n20993 ; n21102
g18667 and pi0907 n16653 ; n21103
g18668 and pi0947_not n21103 ; n21104
g18669 and n3448 n21104_not ; n21105
g18670 nor n21102 n21105 ; n21106
g18671 nor pi0215 n21106 ; n21107
g18672 nor n21101 n21107 ; n21108
g18673 and pi0299 n21108_not ; n21109
g18674 and n17024 n20902 ; n21110
g18675 nor pi0299 n21110 ; n21111
g18676 nor n21109 n21111 ; n21112
g18677 and pi0039 n21112_not ; n21113
g18678 and n16958 n20902 ; n21114
g18679 nor pi0039 n21114 ; n21115
g18680 nor n21113 n21115 ; n21116
g18681 and pi0147 n21116 ; n21117
g18682 nor pi0038 n21117 ; n21118
g18683 and n21100_not n21118 ; n21119
g18684 and pi0770 n21091_not ; n21120
g18685 and n21119_not n21120 ; n21121
g18686 and pi0726 n21087_not ; n21122
g18687 and n21121_not n21122 ; n21123
g18688 and n10197 n21123_not ; n21124
g18689 and n21038_not n21124 ; n21125
g18690 nor pi0832 n20987 ; n21126
g18691 and n21125_not n21126 ; n21127
g18692 nor n20986 n21127 ; po0304
g18693 and pi0057 pi0148 ; n21129
g18694 and n2571 n6305 ; n21130
g18695 nor pi0148 n21130 ; n21131
g18696 and pi0749_not pi0947 ; n21132
g18697 and n21041 n21132_not ; n21133
g18698 nor pi0148 n16641 ; n21134
g18699 nor n21133 n21134 ; n21135
g18700 and pi0038 n21135_not ; n21136
g18701 nor n17025 n21109 ; n21137
g18702 and pi0148 n21137_not ; n21138
g18703 nor n9737 n21095 ; n21139
g18704 nor pi0749 n21138 ; n21140
g18705 and n21139_not n21140 ; n21141
g18706 and pi0148_not n21064 ; n21142
g18707 and pi0148 n21080 ; n21143
g18708 and pi0749 n21143_not ; n21144
g18709 and n21142_not n21144 ; n21145
g18710 and pi0039 n21141_not ; n21146
g18711 and n21145_not n21146 ; n21147
g18712 nor pi0148 n16958 ; n21148
g18713 nor pi0039 n21148 ; n21149
g18714 and n21066 n21132_not ; n21150
g18715 and n21149 n21150_not ; n21151
g18716 nor pi0038 n21151 ; n21152
g18717 and n21147_not n21152 ; n21153
g18718 and pi0706 n21136_not ; n21154
g18719 and n21153_not n21154 ; n21155
g18720 and pi0749 pi0947 ; n21156
g18721 and n16958 n21156 ; n21157
g18722 and n21149 n21157_not ; n21158
g18723 nor pi0148 pi0749 ; n21159
g18724 and n17046_not n21159 ; n21160
g18725 nor pi0148 n21001 ; n21161
g18726 nor n21021 n21028 ; n21162
g18727 and pi0148 n21162_not ; n21163
g18728 and pi0299 n21163_not ; n21164
g18729 and n21161_not n21164 ; n21165
g18730 nor pi0148 n17024 ; n21166
g18731 and n21019 n21166_not ; n21167
g18732 and pi0749 n21167_not ; n21168
g18733 and n21165_not n21168 ; n21169
g18734 and pi0039 n21160_not ; n21170
g18735 and n21169_not n21170 ; n21171
g18736 nor pi0038 n21158 ; n21172
g18737 and n21171_not n21172 ; n21173
g18738 and n16641 n21156_not ; n21174
g18739 and pi0148 n17050_not ; n21175
g18740 and pi0038 n21174_not ; n21176
g18741 and n21175_not n21176 ; n21177
g18742 nor pi0706 n21177 ; n21178
g18743 and n21173_not n21178 ; n21179
g18744 and n21130 n21179_not ; n21180
g18745 and n21155_not n21180 ; n21181
g18746 nor pi0057 n21131 ; n21182
g18747 and n21181_not n21182 ; n21183
g18748 nor pi0832 n21129 ; n21184
g18749 and n21183_not n21184 ; n21185
g18750 and pi0706 n20902 ; n21186
g18751 and n2926 n21156_not ; n21187
g18752 and n21186_not n21187 ; n21188
g18753 and pi0148 n2926_not ; n21189
g18754 and pi0832 n21189_not ; n21190
g18755 and n21188_not n21190 ; n21191
g18756 or n21185 n21191 ; po0305
g18757 nor pi0149 n2926 ; n21193
g18758 and pi0755_not pi0947 ; n21194
g18759 and pi0725_not n20902 ; n21195
g18760 nor n21194 n21195 ; n21196
g18761 and n2926 n21196_not ; n21197
g18762 and pi0832 n21193_not ; n21198
g18763 and n21197_not n21198 ; n21199
g18764 nor pi0149 n10197 ; n21200
g18765 and n16641 n21194_not ; n21201
g18766 and pi0149 n17050_not ; n21202
g18767 and pi0038 n21201_not ; n21203
g18768 and n21202_not n21203 ; n21204
g18769 nor pi0149 n16958 ; n21205
g18770 and n16958 n21194 ; n21206
g18771 nor pi0039 n21205 ; n21207
g18772 and n21206_not n21207 ; n21208
g18773 nor pi0149 n17024 ; n21209
g18774 and n21019 n21209_not ; n21210
g18775 nor pi0149 n21001 ; n21211
g18776 nor n16116 n21029 ; n21212
g18777 nor n21211 n21212 ; n21213
g18778 nor pi0755 n21210 ; n21214
g18779 and n21213_not n21214 ; n21215
g18780 and pi0149_not pi0755 ; n21216
g18781 and n17046_not n21216 ; n21217
g18782 and pi0039 n21217_not ; n21218
g18783 and n21215_not n21218 ; n21219
g18784 nor pi0038 n21208 ; n21220
g18785 and n21219_not n21220 ; n21221
g18786 nor n21204 n21221 ; n21222
g18787 and pi0725 n21222_not ; n21223
g18788 and n21114_not n21208 ; n21224
g18789 and pi0149_not n21064 ; n21225
g18790 and pi0149 n21080 ; n21226
g18791 nor pi0755 n21226 ; n21227
g18792 and n21225_not n21227 ; n21228
g18793 and pi0149_not n21093 ; n21229
g18794 and pi0149 n21137_not ; n21230
g18795 and pi0755 n21094_not ; n21231
g18796 and n21230_not n21231 ; n21232
g18797 and n21229_not n21232 ; n21233
g18798 and pi0039 n21233_not ; n21234
g18799 and n21228_not n21234 ; n21235
g18800 nor n21224 n21235 ; n21236
g18801 nor pi0038 n21236 ; n21237
g18802 nor pi0149 n16641 ; n21238
g18803 and n6236_not n16667 ; n21239
g18804 and pi0755 pi0947 ; n21240
g18805 nor pi0039 n21240 ; n21241
g18806 and n21239 n21241 ; n21242
g18807 and pi0038 n21238_not ; n21243
g18808 and n21242_not n21243 ; n21244
g18809 nor pi0725 n21244 ; n21245
g18810 and n21237_not n21245 ; n21246
g18811 nor n21223 n21246 ; n21247
g18812 and n10197 n21247_not ; n21248
g18813 nor pi0832 n21200 ; n21249
g18814 and n21248_not n21249 ; n21250
g18815 nor n21199 n21250 ; po0306
g18816 nor pi0150 n10197 ; n21252
g18817 and pi0150 n17050_not ; n21253
g18818 and pi0751_not pi0947 ; n21254
g18819 and n16641 n21254_not ; n21255
g18820 nor n21253 n21255 ; n21256
g18821 and pi0038 n21256_not ; n21257
g18822 and pi0150 n16958_not ; n21258
g18823 and pi0751 n16958 ; n21259
g18824 nor n21258 n21259 ; n21260
g18825 and n20989 n21260 ; n21261
g18826 and pi0150_not n21004 ; n21262
g18827 and pi0150 n21030_not ; n21263
g18828 nor pi0751 n21263 ; n21264
g18829 and n21262_not n21264 ; n21265
g18830 and pi0150_not pi0751 ; n21266
g18831 and n17046_not n21266 ; n21267
g18832 nor n21265 n21267 ; n21268
g18833 and pi0039 n21268_not ; n21269
g18834 nor pi0038 n21261 ; n21270
g18835 and n21269_not n21270 ; n21271
g18836 and pi0701 n21257_not ; n21272
g18837 and n21271_not n21272 ; n21273
g18838 nor pi0150 n16641 ; n21274
g18839 and pi0751 pi0947 ; n21275
g18840 nor pi0039 n21275 ; n21276
g18841 and n21239 n21276 ; n21277
g18842 and pi0038 n21274_not ; n21278
g18843 and n21277_not n21278 ; n21279
g18844 and n21097 n21254_not ; n21280
g18845 nor pi0039 n21258 ; n21281
g18846 and n21280_not n21281 ; n21282
g18847 nor pi0150 n21095 ; n21283
g18848 and pi0150 n21112_not ; n21284
g18849 and pi0751 n21284_not ; n21285
g18850 and n21283_not n21285 ; n21286
g18851 and pi0150_not n21064 ; n21287
g18852 and pi0150 n21080 ; n21288
g18853 nor pi0751 n21288 ; n21289
g18854 and n21287_not n21289 ; n21290
g18855 nor n21286 n21290 ; n21291
g18856 and pi0039 n21291_not ; n21292
g18857 nor pi0038 n21282 ; n21293
g18858 and n21292_not n21293 ; n21294
g18859 nor pi0701 n21279 ; n21295
g18860 and n21294_not n21295 ; n21296
g18861 nor n21273 n21296 ; n21297
g18862 and n10197 n21297_not ; n21298
g18863 nor pi0832 n21252 ; n21299
g18864 and n21298_not n21299 ; n21300
g18865 nor pi0150 n2926 ; n21301
g18866 and pi0701_not n20902 ; n21302
g18867 nor n21254 n21302 ; n21303
g18868 and n2926 n21303_not ; n21304
g18869 and pi0832 n21301_not ; n21305
g18870 and n21304_not n21305 ; n21306
g18871 nor n21300 n21306 ; po0307
g18872 nor pi0151 n2926 ; n21308
g18873 and pi0745_not pi0947 ; n21309
g18874 and pi0723_not n20902 ; n21310
g18875 nor n21309 n21310 ; n21311
g18876 and n2926 n21311_not ; n21312
g18877 and pi0832 n21308_not ; n21313
g18878 and n21312_not n21313 ; n21314
g18879 nor pi0151 n10197 ; n21315
g18880 nor pi0151 n16641 ; n21316
g18881 and pi0745 pi0947 ; n21317
g18882 nor pi0039 n21317 ; n21318
g18883 and n21239 n21318 ; n21319
g18884 and pi0038 n21316_not ; n21320
g18885 and n21319_not n21320 ; n21321
g18886 nor pi0151 n16958 ; n21322
g18887 and pi0745_not n21016 ; n21323
g18888 nor n21322 n21323 ; n21324
g18889 and n21115 n21324 ; n21325
g18890 nor n17041 n20999 ; n21326
g18891 and pi0151_not n21326 ; n21327
g18892 nor n17037 n21327 ; n21328
g18893 and pi0215 n21328_not ; n21329
g18894 and pi0151 n3448_not ; n21330
g18895 and n17032_not n21330 ; n21331
g18896 nor n17031 n21331 ; n21332
g18897 nor pi0151 n16653 ; n21333
g18898 and n21105 n21333_not ; n21334
g18899 and n21074_not n21334 ; n21335
g18900 nor pi0215 n21335 ; n21336
g18901 and n21332 n21336 ; n21337
g18902 nor n21329 n21337 ; n21338
g18903 and pi0299 n21338_not ; n21339
g18904 and pi0151 n21071_not ; n21340
g18905 and n21062 n21340_not ; n21341
g18906 nor n21339 n21341 ; n21342
g18907 nor pi0745 n21342 ; n21343
g18908 and n21332 n21334_not ; n21344
g18909 and n21048 n21344 ; n21345
g18910 nor n21329 n21345 ; n21346
g18911 nor n21021 n21346 ; n21347
g18912 and pi0299 n21347_not ; n21348
g18913 nor pi0151 n17024 ; n21349
g18914 and n21111 n21349_not ; n21350
g18915 and pi0745 n21350_not ; n21351
g18916 and n21348_not n21351 ; n21352
g18917 and pi0039 n21352_not ; n21353
g18918 and n21343_not n21353 ; n21354
g18919 nor n21325 n21354 ; n21355
g18920 nor pi0038 n21355 ; n21356
g18921 nor pi0723 n21321 ; n21357
g18922 and n21356_not n21357 ; n21358
g18923 and pi0151 n17050_not ; n21359
g18924 and n16641 n21309_not ; n21360
g18925 nor n21359 n21360 ; n21361
g18926 and pi0038 n21361_not ; n21362
g18927 nor pi0039 n21324 ; n21363
g18928 nor pi0745 n17025 ; n21364
g18929 nor pi0151 n17046 ; n21365
g18930 and n21364_not n21365 ; n21366
g18931 and n21026 n21333_not ; n21367
g18932 and n21332 n21367_not ; n21368
g18933 and n20996 n21368 ; n21369
g18934 and n21101 n21328_not ; n21370
g18935 and pi0299 n21370_not ; n21371
g18936 and n21369_not n21371 ; n21372
g18937 nor pi0745 n21019 ; n21373
g18938 and n21372_not n21373 ; n21374
g18939 nor n21366 n21374 ; n21375
g18940 and pi0039 n21375_not ; n21376
g18941 nor pi0038 n21363 ; n21377
g18942 and n21376_not n21377 ; n21378
g18943 and pi0723 n21362_not ; n21379
g18944 and n21378_not n21379 ; n21380
g18945 nor n21358 n21380 ; n21381
g18946 and n10197 n21381_not ; n21382
g18947 nor pi0832 n21315 ; n21383
g18948 and n21382_not n21383 ; n21384
g18949 nor n21314 n21384 ; po0308
g18950 nor pi0152 n10197 ; n21386
g18951 nor pi0152 n16641 ; n21387
g18952 and pi0759 pi0947 ; n21388
g18953 nor pi0039 n21388 ; n21389
g18954 and n16667 n20902_not ; n21390
g18955 and n21389 n21390 ; n21391
g18956 and pi0038 n21387_not ; n21392
g18957 and n21391_not n21392 ; n21393
g18958 and pi0152 n16958_not ; n21394
g18959 nor n16959 n21389 ; n21395
g18960 nor n21394 n21395 ; n21396
g18961 and n21114_not n21396 ; n21397
g18962 nor pi0152 n17037 ; n21398
g18963 and n20998 n21398_not ; n21399
g18964 nor n20902 n21073 ; n21400
g18965 and n21399 n21400_not ; n21401
g18966 and pi0152 n21046 ; n21402
g18967 and n21102 n21402_not ; n21403
g18968 and pi0152 n16653_not ; n21404
g18969 nor n21074 n21404 ; n21405
g18970 and n3448 n21405 ; n21406
g18971 nor pi0215 n21406 ; n21407
g18972 and n21045_not n21407 ; n21408
g18973 and n21403_not n21408 ; n21409
g18974 and pi0299 n21401_not ; n21410
g18975 and n21409_not n21410 ; n21411
g18976 nor n21104 n21404 ; n21412
g18977 and n2603 n21412_not ; n21413
g18978 nor pi0152 n17020 ; n21414
g18979 and n17020 n20902_not ; n21415
g18980 nor n2603 n21415 ; n21416
g18981 and n21414_not n21416 ; n21417
g18982 nor n21413 n21417 ; n21418
g18983 nor pi0223 n21418 ; n21419
g18984 nor pi0152 n16992 ; n21420
g18985 and n21055 n21420_not ; n21421
g18986 nor pi0299 n21421 ; n21422
g18987 and n21419_not n21422 ; n21423
g18988 nor pi0759 n21411 ; n21424
g18989 and n21423_not n21424 ; n21425
g18990 and n17032_not n21403 ; n21426
g18991 and n21407 n21426_not ; n21427
g18992 and pi0299 n21399_not ; n21428
g18993 and n21427_not n21428 ; n21429
g18994 and n2603 n21405 ; n21430
g18995 and pi0947_not n17020 ; n21431
g18996 nor n2603 n21431 ; n21432
g18997 and n21414_not n21432 ; n21433
g18998 and n6236_not n17020 ; n21434
g18999 nor n2603 n21434 ; n21435
g19000 and n21433_not n21435 ; n21436
g19001 nor pi0223 n21430 ; n21437
g19002 and n21436_not n21437 ; n21438
g19003 and n21053 n21420_not ; n21439
g19004 nor pi0299 n21439 ; n21440
g19005 and n21421_not n21440 ; n21441
g19006 and n21438_not n21441 ; n21442
g19007 and pi0759 n21429_not ; n21443
g19008 and n21442_not n21443 ; n21444
g19009 and pi0039 n21425_not ; n21445
g19010 and n21444_not n21445 ; n21446
g19011 nor pi0038 n21397 ; n21447
g19012 and n21446_not n21447 ; n21448
g19013 and pi0696 n21393_not ; n21449
g19014 and n21448_not n21449 ; n21450
g19015 nor pi0152 n17050 ; n21451
g19016 and n16641 n21388_not ; n21452
g19017 and pi0038 n21452_not ; n21453
g19018 and n21451_not n21453 ; n21454
g19019 nor n21025 n21404 ; n21455
g19020 and n2603 n21455_not ; n21456
g19021 nor n21433 n21456 ; n21457
g19022 nor pi0223 n21457 ; n21458
g19023 and n21440 n21458_not ; n21459
g19024 and pi0152 n21000 ; n21460
g19025 and n3448 n21455 ; n21461
g19026 nor n20995 n21403 ; n21462
g19027 nor n21023 n21462 ; n21463
g19028 nor pi0215 n21461 ; n21464
g19029 and n21463_not n21464 ; n21465
g19030 and n21022 n21460_not ; n21466
g19031 and n21465_not n21466 ; n21467
g19032 and pi0759 n21459_not ; n21468
g19033 and n21467_not n21468 ; n21469
g19034 nor pi0759 n17046 ; n21470
g19035 and pi0152 n21470 ; n21471
g19036 and pi0039 n21471_not ; n21472
g19037 and n21469_not n21472 ; n21473
g19038 nor pi0038 n21396 ; n21474
g19039 and n21473_not n21474 ; n21475
g19040 nor pi0696 n21454 ; n21476
g19041 and n21475_not n21476 ; n21477
g19042 nor n21450 n21477 ; n21478
g19043 and n10197 n21478_not ; n21479
g19044 nor pi0832 n21386 ; n21480
g19045 and n21479_not n21480 ; n21481
g19046 nor pi0152 n2926 ; n21482
g19047 and pi0696 n20902 ; n21483
g19048 and n2926 n21388_not ; n21484
g19049 and n21483_not n21484 ; n21485
g19050 and pi0832 n21482_not ; n21486
g19051 and n21485_not n21486 ; n21487
g19052 or n21481 n21487 ; po0309
g19053 and pi0153 n2926_not ; n21489
g19054 and pi0766 pi0947 ; n21490
g19055 and n2926 n21490_not ; n21491
g19056 and pi0700 n20902 ; n21492
g19057 and n21491 n21492_not ; n21493
g19058 and pi0832 n21489_not ; n21494
g19059 and n21493_not n21494 ; n21495
g19060 and pi0057 pi0153 ; n21496
g19061 nor pi0153 n21130 ; n21497
g19062 nor pi0153 n16958 ; n21498
g19063 and pi0766_not n18147 ; n21499
g19064 nor n21017 n21499 ; n21500
g19065 nor n21498 n21500 ; n21501
g19066 and n21114_not n21501 ; n21502
g19067 nor pi0153 n17024 ; n21503
g19068 and n21111 n21503_not ; n21504
g19069 and pi0153 n17037_not ; n21505
g19070 and n20998 n21505_not ; n21506
g19071 and n21073 n21506_not ; n21507
g19072 and pi0153 n3448_not ; n21508
g19073 and n17032_not n21508 ; n21509
g19074 nor n17031 n21509 ; n21510
g19075 nor pi0153 n16653 ; n21511
g19076 and n21105 n21511_not ; n21512
g19077 nor n21047 n21512 ; n21513
g19078 and n21510 n21513 ; n21514
g19079 nor pi0215 n21514 ; n21515
g19080 nor n21021 n21507 ; n21516
g19081 and n21515_not n21516 ; n21517
g19082 and pi0299 n21517_not ; n21518
g19083 nor pi0766 n21504 ; n21519
g19084 and n21518_not n21519 ; n21520
g19085 and n21026 n21511_not ; n21521
g19086 and n21103_not n21521 ; n21522
g19087 nor pi0215 n21522 ; n21523
g19088 and n21510 n21523 ; n21524
g19089 nor n21506 n21524 ; n21525
g19090 and pi0299 n21525_not ; n21526
g19091 and pi0153 n21071_not ; n21527
g19092 and n21062 n21527_not ; n21528
g19093 nor n21526 n21528 ; n21529
g19094 and pi0766 n21529_not ; n21530
g19095 and pi0039 n21520_not ; n21531
g19096 and n21530_not n21531 ; n21532
g19097 nor n21502 n21532 ; n21533
g19098 nor pi0038 n21533 ; n21534
g19099 nor pi0153 n16641 ; n21535
g19100 and pi0766_not pi0947 ; n21536
g19101 nor pi0039 n21536 ; n21537
g19102 and n21239 n21537 ; n21538
g19103 and pi0038 n21535_not ; n21539
g19104 and n21538_not n21539 ; n21540
g19105 nor n21534 n21540 ; n21541
g19106 and pi0700 n21541_not ; n21542
g19107 and n6284 n21491 ; n21543
g19108 and pi0153 n17050_not ; n21544
g19109 and pi0038 n21543_not ; n21545
g19110 and n21544_not n21545 ; n21546
g19111 and n21019 n21503_not ; n21547
g19112 and n21000 n21505_not ; n21548
g19113 and n21510 n21521_not ; n21549
g19114 and n20996 n21549 ; n21550
g19115 and pi0299 n21548_not ; n21551
g19116 and n21550_not n21551 ; n21552
g19117 and pi0766 n21552_not ; n21553
g19118 and n21547_not n21553 ; n21554
g19119 nor pi0153 pi0766 ; n21555
g19120 and n17046_not n21555 ; n21556
g19121 and pi0039 n21556_not ; n21557
g19122 and n21554_not n21557 ; n21558
g19123 nor pi0038 n21501 ; n21559
g19124 and n21558_not n21559 ; n21560
g19125 nor pi0700 n21546 ; n21561
g19126 and n21560_not n21561 ; n21562
g19127 and n21130 n21562_not ; n21563
g19128 and n21542_not n21563 ; n21564
g19129 nor pi0057 n21497 ; n21565
g19130 and n21564_not n21565 ; n21566
g19131 nor pi0832 n21496 ; n21567
g19132 and n21566_not n21567 ; n21568
g19133 or n21495 n21568 ; po0310
g19134 nor pi0154 n2926 ; n21570
g19135 and pi0742_not pi0947 ; n21571
g19136 and pi0704_not n20902 ; n21572
g19137 nor n21571 n21572 ; n21573
g19138 and n2926 n21573_not ; n21574
g19139 and pi0832 n21570_not ; n21575
g19140 and n21574_not n21575 ; n21576
g19141 nor pi0154 n10197 ; n21577
g19142 nor pi0154 n16641 ; n21578
g19143 and n21090 n21578_not ; n21579
g19144 nor pi0154 n16958 ; n21580
g19145 and n21115 n21580_not ; n21581
g19146 and pi0154_not n21095 ; n21582
g19147 and pi0154 n21112 ; n21583
g19148 and pi0039 n21583_not ; n21584
g19149 and n21582_not n21584 ; n21585
g19150 nor n21581 n21585 ; n21586
g19151 nor pi0038 n21586 ; n21587
g19152 and pi0742 n21579_not ; n21588
g19153 and n21587_not n21588 ; n21589
g19154 and n21042 n21578_not ; n21590
g19155 and n21066_not n21581 ; n21591
g19156 nor pi0154 n21064 ; n21592
g19157 and pi0154 n21080_not ; n21593
g19158 and pi0039 n21593_not ; n21594
g19159 and n21592_not n21594 ; n21595
g19160 nor n21591 n21595 ; n21596
g19161 nor pi0038 n21596 ; n21597
g19162 nor pi0742 n21590 ; n21598
g19163 and n21597_not n21598 ; n21599
g19164 nor pi0704 n21589 ; n21600
g19165 and n21599_not n21600 ; n21601
g19166 nor pi0154 n17050 ; n21602
g19167 nor n21015 n21602 ; n21603
g19168 and n21017 n21580_not ; n21604
g19169 and pi0154 n21030 ; n21605
g19170 nor pi0154 n21004 ; n21606
g19171 and pi0039 n21605_not ; n21607
g19172 and n21606_not n21607 ; n21608
g19173 nor n21604 n21608 ; n21609
g19174 nor pi0038 n21609 ; n21610
g19175 nor pi0742 n21603 ; n21611
g19176 and n21610_not n21611 ; n21612
g19177 and pi0154_not pi0742 ; n21613
g19178 and n17052_not n21613 ; n21614
g19179 and pi0704 n21614_not ; n21615
g19180 and n21612_not n21615 ; n21616
g19181 and n10197 n21616_not ; n21617
g19182 and n21601_not n21617 ; n21618
g19183 nor pi0832 n21577 ; n21619
g19184 and n21618_not n21619 ; n21620
g19185 nor n21576 n21620 ; po0311
g19186 and pi0757_not n21034 ; n21622
g19187 and pi0686 n21622_not ; n21623
g19188 nor pi0038 n21082 ; n21624
g19189 nor n21042 n21624 ; n21625
g19190 and pi0757_not n21625 ; n21626
g19191 nor pi0038 n21116 ; n21627
g19192 nor n21090 n21627 ; n21628
g19193 and pi0757 n21628 ; n21629
g19194 nor pi0686 n21626 ; n21630
g19195 and n21629_not n21630 ; n21631
g19196 and n10197 n21623_not ; n21632
g19197 and n21631_not n21632 ; n21633
g19198 and pi0155 n21633_not ; n21634
g19199 nor pi0038 n21069 ; n21635
g19200 and pi0038 n21039 ; n21636
g19201 nor n21635 n21636 ; n21637
g19202 and pi0757_not n21637 ; n21638
g19203 nor pi0038 n21099 ; n21639
g19204 and n16641 n21090 ; n21640
g19205 nor n21639 n21640 ; n21641
g19206 and pi0757 n21641 ; n21642
g19207 nor pi0686 n21638 ; n21643
g19208 and n21642_not n21643 ; n21644
g19209 and pi0757_not n21010 ; n21645
g19210 and pi0757 n17052_not ; n21646
g19211 and pi0686 n21646_not ; n21647
g19212 and n21645_not n21647 ; n21648
g19213 nor n21644 n21648 ; n21649
g19214 and pi0155_not n10197 ; n21650
g19215 and n21649_not n21650 ; n21651
g19216 nor n21634 n21651 ; n21652
g19217 nor pi0832 n21652 ; n21653
g19218 nor pi0155 n2926 ; n21654
g19219 and pi0757_not pi0947 ; n21655
g19220 and pi0686_not n20902 ; n21656
g19221 nor n21655 n21656 ; n21657
g19222 and n2926 n21657_not ; n21658
g19223 and pi0832 n21654_not ; n21659
g19224 and n21658_not n21659 ; n21660
g19225 nor n21653 n21660 ; po0312
g19226 nor pi0156 n2926 ; n21662
g19227 and pi0741_not pi0947 ; n21663
g19228 and pi0724_not n20902 ; n21664
g19229 nor n21663 n21664 ; n21665
g19230 and n2926 n21665_not ; n21666
g19231 and pi0832 n21662_not ; n21667
g19232 and n21666_not n21667 ; n21668
g19233 nor pi0741 n21637 ; n21669
g19234 and pi0741 n21641_not ; n21670
g19235 nor pi0724 n21669 ; n21671
g19236 and n21670_not n21671 ; n21672
g19237 nor pi0741 n21010 ; n21673
g19238 and pi0741 n17052 ; n21674
g19239 and pi0724 n21674_not ; n21675
g19240 and n21673_not n21675 ; n21676
g19241 and n10197 n21676_not ; n21677
g19242 and n21672_not n21677 ; n21678
g19243 nor pi0156 n21678 ; n21679
g19244 nor pi0741 n21625 ; n21680
g19245 and pi0741 n21628_not ; n21681
g19246 nor pi0724 n21680 ; n21682
g19247 and n21681_not n21682 ; n21683
g19248 and pi0724 pi0741_not ; n21684
g19249 and n21034 n21684 ; n21685
g19250 nor n21683 n21685 ; n21686
g19251 and pi0156 n10197 ; n21687
g19252 and n21686_not n21687 ; n21688
g19253 nor pi0832 n21688 ; n21689
g19254 and n21679_not n21689 ; n21690
g19255 nor n21668 n21690 ; po0313
g19256 nor pi0157 n2926 ; n21692
g19257 and pi0760_not pi0947 ; n21693
g19258 and pi0688_not n20902 ; n21694
g19259 nor n21693 n21694 ; n21695
g19260 and n2926 n21695_not ; n21696
g19261 and pi0832 n21692_not ; n21697
g19262 and n21696_not n21697 ; n21698
g19263 nor pi0157 n10197 ; n21699
g19264 and n16641 n21693_not ; n21700
g19265 and pi0157 n17050_not ; n21701
g19266 and pi0038 n21700_not ; n21702
g19267 and n21701_not n21702 ; n21703
g19268 and pi0157_not pi0760 ; n21704
g19269 and n17046_not n21704 ; n21705
g19270 nor pi0157 n17024 ; n21706
g19271 and n21019 n21706_not ; n21707
g19272 nor pi0157 n21001 ; n21708
g19273 nor n13717 n21029 ; n21709
g19274 nor n21708 n21709 ; n21710
g19275 nor pi0760 n21707 ; n21711
g19276 and n21710_not n21711 ; n21712
g19277 and pi0039 n21705_not ; n21713
g19278 and n21712_not n21713 ; n21714
g19279 nor pi0157 n16958 ; n21715
g19280 and n16958 n21693 ; n21716
g19281 nor pi0039 n21715 ; n21717
g19282 and n21716_not n21717 ; n21718
g19283 nor pi0038 n21718 ; n21719
g19284 and n21714_not n21719 ; n21720
g19285 nor n21703 n21720 ; n21721
g19286 and pi0688 n21721_not ; n21722
g19287 and n21114_not n21718 ; n21723
g19288 and pi0760_not n21080 ; n21724
g19289 and pi0760 n21112_not ; n21725
g19290 and pi0157 n21724_not ; n21726
g19291 and n21725_not n21726 ; n21727
g19292 and pi0760 n21095_not ; n21728
g19293 and pi0760_not n21064 ; n21729
g19294 nor pi0157 n21728 ; n21730
g19295 and n21729_not n21730 ; n21731
g19296 and pi0039 n21727_not ; n21732
g19297 and n21731_not n21732 ; n21733
g19298 nor n21723 n21733 ; n21734
g19299 nor pi0038 n21734 ; n21735
g19300 nor pi0157 n16641 ; n21736
g19301 and pi0760 pi0947 ; n21737
g19302 nor pi0039 n21737 ; n21738
g19303 and n21239 n21738 ; n21739
g19304 and pi0038 n21736_not ; n21740
g19305 and n21739_not n21740 ; n21741
g19306 nor pi0688 n21741 ; n21742
g19307 and n21735_not n21742 ; n21743
g19308 nor n21722 n21743 ; n21744
g19309 and n10197 n21744_not ; n21745
g19310 nor pi0832 n21699 ; n21746
g19311 and n21745_not n21746 ; n21747
g19312 nor n21698 n21747 ; po0314
g19313 nor pi0158 n10197 ; n21749
g19314 and pi0158 n17050_not ; n21750
g19315 and pi0753_not pi0947 ; n21751
g19316 and n16641 n21751_not ; n21752
g19317 nor n21750 n21752 ; n21753
g19318 and pi0038 n21753_not ; n21754
g19319 and pi0158 n16958_not ; n21755
g19320 and pi0753 n16958 ; n21756
g19321 nor n21755 n21756 ; n21757
g19322 and n20989 n21757 ; n21758
g19323 and pi0158_not n21004 ; n21759
g19324 and pi0158 n21030_not ; n21760
g19325 nor pi0753 n21760 ; n21761
g19326 and n21759_not n21761 ; n21762
g19327 and pi0158_not pi0753 ; n21763
g19328 and n17046_not n21763 ; n21764
g19329 nor n21762 n21764 ; n21765
g19330 and pi0039 n21765_not ; n21766
g19331 nor pi0038 n21758 ; n21767
g19332 and n21766_not n21767 ; n21768
g19333 and pi0702 n21754_not ; n21769
g19334 and n21768_not n21769 ; n21770
g19335 nor pi0158 n16641 ; n21771
g19336 and pi0753 pi0947 ; n21772
g19337 nor pi0039 n21772 ; n21773
g19338 and n21239 n21773 ; n21774
g19339 and pi0038 n21771_not ; n21775
g19340 and n21774_not n21775 ; n21776
g19341 and n21097 n21751_not ; n21777
g19342 nor pi0039 n21755 ; n21778
g19343 and n21777_not n21778 ; n21779
g19344 nor pi0158 n21095 ; n21780
g19345 and pi0158 n21112_not ; n21781
g19346 and pi0753 n21781_not ; n21782
g19347 and n21780_not n21782 ; n21783
g19348 and pi0158_not n21064 ; n21784
g19349 and pi0158 n21080 ; n21785
g19350 nor pi0753 n21785 ; n21786
g19351 and n21784_not n21786 ; n21787
g19352 nor n21783 n21787 ; n21788
g19353 and pi0039 n21788_not ; n21789
g19354 nor pi0038 n21779 ; n21790
g19355 and n21789_not n21790 ; n21791
g19356 nor pi0702 n21776 ; n21792
g19357 and n21791_not n21792 ; n21793
g19358 nor n21770 n21793 ; n21794
g19359 and n10197 n21794_not ; n21795
g19360 nor pi0832 n21749 ; n21796
g19361 and n21795_not n21796 ; n21797
g19362 nor pi0158 n2926 ; n21798
g19363 and pi0702_not n20902 ; n21799
g19364 nor n21751 n21799 ; n21800
g19365 and n2926 n21800_not ; n21801
g19366 and pi0832 n21798_not ; n21802
g19367 and n21801_not n21802 ; n21803
g19368 nor n21797 n21803 ; po0315
g19369 nor pi0159 n10197 ; n21805
g19370 and pi0159 n17050_not ; n21806
g19371 and pi0754_not pi0947 ; n21807
g19372 and n16641 n21807_not ; n21808
g19373 nor n21806 n21808 ; n21809
g19374 and pi0038 n21809_not ; n21810
g19375 and pi0159 n16958_not ; n21811
g19376 and pi0754 n16958 ; n21812
g19377 nor n21811 n21812 ; n21813
g19378 and n20989 n21813 ; n21814
g19379 and pi0159_not n21004 ; n21815
g19380 and pi0159 n21030_not ; n21816
g19381 nor pi0754 n21816 ; n21817
g19382 and n21815_not n21817 ; n21818
g19383 and pi0159_not pi0754 ; n21819
g19384 and n17046_not n21819 ; n21820
g19385 nor n21818 n21820 ; n21821
g19386 and pi0039 n21821_not ; n21822
g19387 nor pi0038 n21814 ; n21823
g19388 and n21822_not n21823 ; n21824
g19389 and pi0709 n21810_not ; n21825
g19390 and n21824_not n21825 ; n21826
g19391 nor pi0159 n16641 ; n21827
g19392 and pi0754 pi0947 ; n21828
g19393 nor pi0039 n21828 ; n21829
g19394 and n21239 n21829 ; n21830
g19395 and pi0038 n21827_not ; n21831
g19396 and n21830_not n21831 ; n21832
g19397 and n21097 n21807_not ; n21833
g19398 nor pi0039 n21811 ; n21834
g19399 and n21833_not n21834 ; n21835
g19400 nor pi0159 n21095 ; n21836
g19401 and pi0159 n21112_not ; n21837
g19402 and pi0754 n21837_not ; n21838
g19403 and n21836_not n21838 ; n21839
g19404 and pi0159_not n21064 ; n21840
g19405 and pi0159 n21080 ; n21841
g19406 nor pi0754 n21841 ; n21842
g19407 and n21840_not n21842 ; n21843
g19408 nor n21839 n21843 ; n21844
g19409 and pi0039 n21844_not ; n21845
g19410 nor pi0038 n21835 ; n21846
g19411 and n21845_not n21846 ; n21847
g19412 nor pi0709 n21832 ; n21848
g19413 and n21847_not n21848 ; n21849
g19414 nor n21826 n21849 ; n21850
g19415 and n10197 n21850_not ; n21851
g19416 nor pi0832 n21805 ; n21852
g19417 and n21851_not n21852 ; n21853
g19418 nor pi0159 n2926 ; n21854
g19419 and pi0709_not n20902 ; n21855
g19420 nor n21807 n21855 ; n21856
g19421 and n2926 n21856_not ; n21857
g19422 and pi0832 n21854_not ; n21858
g19423 and n21857_not n21858 ; n21859
g19424 nor n21853 n21859 ; po0316
g19425 nor pi0160 n2926 ; n21861
g19426 and pi0756_not pi0947 ; n21862
g19427 and pi0734_not n20902 ; n21863
g19428 nor n21862 n21863 ; n21864
g19429 and n2926 n21864_not ; n21865
g19430 and pi0832 n21861_not ; n21866
g19431 and n21865_not n21866 ; n21867
g19432 nor pi0160 n10197 ; n21868
g19433 and n16641 n21862_not ; n21869
g19434 and pi0160 n17050_not ; n21870
g19435 and pi0038 n21869_not ; n21871
g19436 and n21870_not n21871 ; n21872
g19437 nor pi0160 n16958 ; n21873
g19438 and n16958 n21862 ; n21874
g19439 nor pi0039 n21873 ; n21875
g19440 and n21874_not n21875 ; n21876
g19441 nor pi0160 n21001 ; n21877
g19442 and pi0160 n21162_not ; n21878
g19443 and pi0299 n21878_not ; n21879
g19444 and n21877_not n21879 ; n21880
g19445 nor pi0160 n17024 ; n21881
g19446 and n21019 n21881_not ; n21882
g19447 nor pi0756 n21882 ; n21883
g19448 and n21880_not n21883 ; n21884
g19449 and pi0160_not pi0756 ; n21885
g19450 and n17046_not n21885 ; n21886
g19451 and pi0039 n21886_not ; n21887
g19452 and n21884_not n21887 ; n21888
g19453 nor pi0038 n21876 ; n21889
g19454 and n21888_not n21889 ; n21890
g19455 nor n21872 n21890 ; n21891
g19456 and pi0734 n21891_not ; n21892
g19457 and n21114_not n21876 ; n21893
g19458 and pi0160_not n21064 ; n21894
g19459 and pi0160 n21080 ; n21895
g19460 nor pi0756 n21895 ; n21896
g19461 and n21894_not n21896 ; n21897
g19462 and pi0160 n21137_not ; n21898
g19463 and pi0160_not n21093 ; n21899
g19464 and pi0756 n21094_not ; n21900
g19465 and n21898_not n21900 ; n21901
g19466 and n21899_not n21901 ; n21902
g19467 and pi0039 n21902_not ; n21903
g19468 and n21897_not n21903 ; n21904
g19469 nor n21893 n21904 ; n21905
g19470 nor pi0038 n21905 ; n21906
g19471 nor pi0160 n16641 ; n21907
g19472 and pi0756 pi0947 ; n21908
g19473 nor pi0039 n21908 ; n21909
g19474 and n21239 n21909 ; n21910
g19475 and pi0038 n21907_not ; n21911
g19476 and n21910_not n21911 ; n21912
g19477 nor pi0734 n21912 ; n21913
g19478 and n21906_not n21913 ; n21914
g19479 nor n21892 n21914 ; n21915
g19480 and n10197 n21915_not ; n21916
g19481 nor pi0832 n21868 ; n21917
g19482 and n21916_not n21917 ; n21918
g19483 nor n21867 n21918 ; po0317
g19484 nor pi0161 n10197 ; n21920
g19485 nor pi0161 n16641 ; n21921
g19486 and pi0758 pi0947 ; n21922
g19487 nor pi0039 n21922 ; n21923
g19488 and n21390 n21923 ; n21924
g19489 and pi0038 n21921_not ; n21925
g19490 and n21924_not n21925 ; n21926
g19491 and n16958 n21922 ; n21927
g19492 and pi0161 n16958_not ; n21928
g19493 nor pi0039 n21927 ; n21929
g19494 and n21928_not n21929 ; n21930
g19495 and n21114_not n21930 ; n21931
g19496 nor pi0161 n17037 ; n21932
g19497 and n20998 n21932_not ; n21933
g19498 and n21400_not n21933 ; n21934
g19499 and pi0161 n21046 ; n21935
g19500 and n21102 n21935_not ; n21936
g19501 and pi0161 n16653_not ; n21937
g19502 nor n21074 n21937 ; n21938
g19503 and n3448 n21938 ; n21939
g19504 nor pi0215 n21939 ; n21940
g19505 and n21045_not n21940 ; n21941
g19506 and n21936_not n21941 ; n21942
g19507 and pi0299 n21934_not ; n21943
g19508 and n21942_not n21943 ; n21944
g19509 nor n21104 n21937 ; n21945
g19510 and n2603 n21945_not ; n21946
g19511 nor pi0161 n17020 ; n21947
g19512 and n21416 n21947_not ; n21948
g19513 nor n21946 n21948 ; n21949
g19514 nor pi0223 n21949 ; n21950
g19515 nor pi0161 n16992 ; n21951
g19516 and n21055 n21951_not ; n21952
g19517 nor pi0299 n21952 ; n21953
g19518 and n21950_not n21953 ; n21954
g19519 nor pi0758 n21944 ; n21955
g19520 and n21954_not n21955 ; n21956
g19521 and n17032_not n21936 ; n21957
g19522 and n21940 n21957_not ; n21958
g19523 and pi0299 n21933_not ; n21959
g19524 and n21958_not n21959 ; n21960
g19525 and n2603 n21938 ; n21961
g19526 and n21432 n21947_not ; n21962
g19527 and n21435 n21962_not ; n21963
g19528 nor pi0223 n21961 ; n21964
g19529 and n21963_not n21964 ; n21965
g19530 and n21053 n21951_not ; n21966
g19531 nor pi0299 n21966 ; n21967
g19532 and n21952_not n21967 ; n21968
g19533 and n21965_not n21968 ; n21969
g19534 and pi0758 n21960_not ; n21970
g19535 and n21969_not n21970 ; n21971
g19536 and pi0039 n21956_not ; n21972
g19537 and n21971_not n21972 ; n21973
g19538 nor pi0038 n21931 ; n21974
g19539 and n21973_not n21974 ; n21975
g19540 and pi0736 n21926_not ; n21976
g19541 and n21975_not n21976 ; n21977
g19542 nor pi0161 n17050 ; n21978
g19543 and n16641 n21922_not ; n21979
g19544 and pi0038 n21979_not ; n21980
g19545 and n21978_not n21980 ; n21981
g19546 nor n21025 n21937 ; n21982
g19547 and n2603 n21982_not ; n21983
g19548 nor n21962 n21983 ; n21984
g19549 nor pi0223 n21984 ; n21985
g19550 and n21967 n21985_not ; n21986
g19551 and pi0161 n21000 ; n21987
g19552 and n3448 n21982 ; n21988
g19553 nor n20995 n21936 ; n21989
g19554 nor n21023 n21989 ; n21990
g19555 nor pi0215 n21988 ; n21991
g19556 and n21990_not n21991 ; n21992
g19557 and n21022 n21987_not ; n21993
g19558 and n21992_not n21993 ; n21994
g19559 and pi0758 n21986_not ; n21995
g19560 and n21994_not n21995 ; n21996
g19561 and pi0161 n19958 ; n21997
g19562 and pi0039 n21997_not ; n21998
g19563 and n21996_not n21998 ; n21999
g19564 nor pi0038 n21930 ; n22000
g19565 and n21999_not n22000 ; n22001
g19566 nor pi0736 n21981 ; n22002
g19567 and n22001_not n22002 ; n22003
g19568 nor n21977 n22003 ; n22004
g19569 and n10197 n22004_not ; n22005
g19570 nor pi0832 n21920 ; n22006
g19571 and n22005_not n22006 ; n22007
g19572 nor pi0161 n2926 ; n22008
g19573 and pi0736 n20902 ; n22009
g19574 and n2926 n21922_not ; n22010
g19575 and n22009_not n22010 ; n22011
g19576 and pi0832 n22008_not ; n22012
g19577 and n22011_not n22012 ; n22013
g19578 or n22007 n22013 ; po0318
g19579 nor pi0162 n10197 ; n22015
g19580 and pi0761_not pi0947 ; n22016
g19581 and n16641 n22016_not ; n22017
g19582 and pi0162 n17050_not ; n22018
g19583 and pi0038 n22017_not ; n22019
g19584 and n22018_not n22019 ; n22020
g19585 nor pi0162 n16958 ; n22021
g19586 and n16958 n22016 ; n22022
g19587 nor pi0039 n22021 ; n22023
g19588 and n22022_not n22023 ; n22024
g19589 and n14933 n21162_not ; n22025
g19590 nor n20991 n22025 ; n22026
g19591 nor pi0761 n22026 ; n22027
g19592 and pi0761_not n21003 ; n22028
g19593 and pi0761 n17046 ; n22029
g19594 nor pi0162 n22029 ; n22030
g19595 and n22028_not n22030 ; n22031
g19596 and pi0039 n22027_not ; n22032
g19597 and n22031_not n22032 ; n22033
g19598 nor pi0038 n22024 ; n22034
g19599 and n22033_not n22034 ; n22035
g19600 nor n22020 n22035 ; n22036
g19601 and pi0738 n22036_not ; n22037
g19602 and n21114_not n22024 ; n22038
g19603 and pi0162 n21137_not ; n22039
g19604 nor n14933 n21095 ; n22040
g19605 and pi0761 n22039_not ; n22041
g19606 and n22040_not n22041 ; n22042
g19607 and pi0162_not n21064 ; n22043
g19608 and pi0162 n21080 ; n22044
g19609 nor pi0761 n22044 ; n22045
g19610 and n22043_not n22045 ; n22046
g19611 and pi0039 n22042_not ; n22047
g19612 and n22046_not n22047 ; n22048
g19613 nor n22038 n22048 ; n22049
g19614 nor pi0038 n22049 ; n22050
g19615 nor pi0162 n16641 ; n22051
g19616 and pi0761 pi0947 ; n22052
g19617 nor pi0039 n22052 ; n22053
g19618 and n21239 n22053 ; n22054
g19619 and pi0038 n22051_not ; n22055
g19620 and n22054_not n22055 ; n22056
g19621 nor pi0738 n22056 ; n22057
g19622 and n22050_not n22057 ; n22058
g19623 nor n22037 n22058 ; n22059
g19624 and n10197 n22059_not ; n22060
g19625 nor pi0832 n22015 ; n22061
g19626 and n22060_not n22061 ; n22062
g19627 nor pi0162 n2926 ; n22063
g19628 and pi0738_not n20902 ; n22064
g19629 nor n22016 n22064 ; n22065
g19630 and n2926 n22065_not ; n22066
g19631 and pi0832 n22063_not ; n22067
g19632 and n22066_not n22067 ; n22068
g19633 nor n22062 n22068 ; po0319
g19634 nor pi0163 n2926 ; n22070
g19635 and pi0777_not pi0947 ; n22071
g19636 and pi0737_not n20902 ; n22072
g19637 nor n22071 n22072 ; n22073
g19638 and n2926 n22073_not ; n22074
g19639 and pi0832 n22070_not ; n22075
g19640 and n22074_not n22075 ; n22076
g19641 nor pi0163 n10197 ; n22077
g19642 and n16641 n22071_not ; n22078
g19643 and pi0163 n17050_not ; n22079
g19644 and pi0038 n22078_not ; n22080
g19645 and n22079_not n22080 ; n22081
g19646 nor pi0163 n16958 ; n22082
g19647 and n16958 n22071 ; n22083
g19648 nor pi0039 n22082 ; n22084
g19649 and n22083_not n22084 ; n22085
g19650 nor pi0163 n17024 ; n22086
g19651 and n21019 n22086_not ; n22087
g19652 nor pi0163 n21001 ; n22088
g19653 nor n14735 n21029 ; n22089
g19654 nor n22088 n22089 ; n22090
g19655 nor pi0777 n22087 ; n22091
g19656 and n22090_not n22091 ; n22092
g19657 and pi0163_not pi0777 ; n22093
g19658 and n17046_not n22093 ; n22094
g19659 and pi0039 n22094_not ; n22095
g19660 and n22092_not n22095 ; n22096
g19661 nor pi0038 n22085 ; n22097
g19662 and n22096_not n22097 ; n22098
g19663 nor n22081 n22098 ; n22099
g19664 and pi0737 n22099_not ; n22100
g19665 and n21114_not n22085 ; n22101
g19666 and pi0163_not n21064 ; n22102
g19667 and pi0163 n21080 ; n22103
g19668 nor pi0777 n22103 ; n22104
g19669 and n22102_not n22104 ; n22105
g19670 and pi0163_not n21093 ; n22106
g19671 and pi0163 n21137_not ; n22107
g19672 and pi0777 n21094_not ; n22108
g19673 and n22107_not n22108 ; n22109
g19674 and n22106_not n22109 ; n22110
g19675 and pi0039 n22110_not ; n22111
g19676 and n22105_not n22111 ; n22112
g19677 nor n22101 n22112 ; n22113
g19678 nor pi0038 n22113 ; n22114
g19679 nor pi0163 n16641 ; n22115
g19680 and pi0777 pi0947 ; n22116
g19681 nor pi0039 n22116 ; n22117
g19682 and n21239 n22117 ; n22118
g19683 and pi0038 n22115_not ; n22119
g19684 and n22118_not n22119 ; n22120
g19685 nor pi0737 n22120 ; n22121
g19686 and n22114_not n22121 ; n22122
g19687 nor n22100 n22122 ; n22123
g19688 and n10197 n22123_not ; n22124
g19689 nor pi0832 n22077 ; n22125
g19690 and n22124_not n22125 ; n22126
g19691 nor n22076 n22126 ; po0320
g19692 nor pi0164 n2926 ; n22128
g19693 and pi0752_not pi0947 ; n22129
g19694 and pi0703 n20902 ; n22130
g19695 nor n22129 n22130 ; n22131
g19696 and n2926 n22131_not ; n22132
g19697 and pi0832 n22128_not ; n22133
g19698 and n22132_not n22133 ; n22134
g19699 nor pi0164 n10197 ; n22135
g19700 nor pi0164 n21039 ; n22136
g19701 and n21042 n22136_not ; n22137
g19702 and pi0164_not n21069 ; n22138
g19703 and pi0164 n21082 ; n22139
g19704 nor pi0038 n22139 ; n22140
g19705 and n22138_not n22140 ; n22141
g19706 nor pi0752 n22137 ; n22142
g19707 and n22141_not n22142 ; n22143
g19708 nor pi0164 n16641 ; n22144
g19709 and n21090 n22144_not ; n22145
g19710 and pi0164_not n21099 ; n22146
g19711 and pi0164 n21116 ; n22147
g19712 nor pi0038 n22147 ; n22148
g19713 and n22146_not n22148 ; n22149
g19714 and pi0752 n22145_not ; n22150
g19715 and n22149_not n22150 ; n22151
g19716 nor n22143 n22151 ; n22152
g19717 and pi0703 n22152_not ; n22153
g19718 and pi0752 n17052 ; n22154
g19719 and pi0752_not n21034 ; n22155
g19720 and pi0164 n22155_not ; n22156
g19721 and pi0164 n21009_not ; n22157
g19722 nor pi0752 n22157 ; n22158
g19723 and n21010_not n22158 ; n22159
g19724 nor pi0703 n22154 ; n22160
g19725 and n22156_not n22160 ; n22161
g19726 and n22159_not n22161 ; n22162
g19727 nor n22153 n22162 ; n22163
g19728 and n10197 n22163_not ; n22164
g19729 nor pi0832 n22135 ; n22165
g19730 and n22164_not n22165 ; n22166
g19731 nor n22134 n22166 ; po0321
g19732 nor pi0165 n2926 ; n22168
g19733 and pi0774_not pi0947 ; n22169
g19734 and pi0687 n20902 ; n22170
g19735 nor n22169 n22170 ; n22171
g19736 and n2926 n22171_not ; n22172
g19737 and pi0832 n22168_not ; n22173
g19738 and n22172_not n22173 ; n22174
g19739 nor pi0165 n10197 ; n22175
g19740 nor pi0165 n21039 ; n22176
g19741 and n21042 n22176_not ; n22177
g19742 and pi0165_not n21069 ; n22178
g19743 and pi0165 n21082 ; n22179
g19744 nor pi0038 n22179 ; n22180
g19745 and n22178_not n22180 ; n22181
g19746 nor pi0774 n22177 ; n22182
g19747 and n22181_not n22182 ; n22183
g19748 nor pi0165 n16641 ; n22184
g19749 and n21090 n22184_not ; n22185
g19750 and pi0165_not n21099 ; n22186
g19751 and pi0165 n21116 ; n22187
g19752 nor pi0038 n22187 ; n22188
g19753 and n22186_not n22188 ; n22189
g19754 and pi0774 n22185_not ; n22190
g19755 and n22189_not n22190 ; n22191
g19756 nor n22183 n22191 ; n22192
g19757 and pi0687 n22192_not ; n22193
g19758 and pi0774 n17052 ; n22194
g19759 and pi0774_not n21034 ; n22195
g19760 and pi0165 n22195_not ; n22196
g19761 and pi0165 n21009_not ; n22197
g19762 nor pi0774 n22197 ; n22198
g19763 and n21010_not n22198 ; n22199
g19764 nor pi0687 n22194 ; n22200
g19765 and n22196_not n22200 ; n22201
g19766 and n22199_not n22201 ; n22202
g19767 nor n22193 n22202 ; n22203
g19768 and n10197 n22203_not ; n22204
g19769 nor pi0832 n22175 ; n22205
g19770 and n22204_not n22205 ; n22206
g19771 nor n22174 n22206 ; po0322
g19772 nor pi0166 n10197 ; n22208
g19773 nor pi0166 n17050 ; n22209
g19774 and pi0772 pi0947 ; n22210
g19775 and n16641 n22210_not ; n22211
g19776 and pi0038 n22211_not ; n22212
g19777 and n22209_not n22212 ; n22213
g19778 and pi0166 n16958_not ; n22214
g19779 nor pi0039 n22210 ; n22215
g19780 nor n16959 n22215 ; n22216
g19781 nor n22214 n22216 ; n22217
g19782 nor pi0166 n16992 ; n22218
g19783 and n21053 n22218_not ; n22219
g19784 nor pi0299 n22219 ; n22220
g19785 and pi0166 n16653_not ; n22221
g19786 nor n21025 n22221 ; n22222
g19787 and n2603 n22222_not ; n22223
g19788 nor pi0166 n17020 ; n22224
g19789 and n21432 n22224_not ; n22225
g19790 nor n22223 n22225 ; n22226
g19791 nor pi0223 n22226 ; n22227
g19792 and n22220 n22227_not ; n22228
g19793 and pi0166 n21000 ; n22229
g19794 and n3448 n22222 ; n22230
g19795 and pi0166 n21046 ; n22231
g19796 and n21102 n22231_not ; n22232
g19797 nor n20995 n22232 ; n22233
g19798 nor n21023 n22233 ; n22234
g19799 nor pi0215 n22230 ; n22235
g19800 and n22234_not n22235 ; n22236
g19801 and n21022 n22229_not ; n22237
g19802 and n22236_not n22237 ; n22238
g19803 and pi0772 n22228_not ; n22239
g19804 and n22238_not n22239 ; n22240
g19805 nor pi0772 n17046 ; n22241
g19806 and pi0166 n22241 ; n22242
g19807 and pi0039 n22242_not ; n22243
g19808 and n22240_not n22243 ; n22244
g19809 nor pi0038 n22217 ; n22245
g19810 and n22244_not n22245 ; n22246
g19811 nor pi0727 n22213 ; n22247
g19812 and n22246_not n22247 ; n22248
g19813 and n21390 n22215 ; n22249
g19814 nor pi0166 n16641 ; n22250
g19815 and pi0038 n22249_not ; n22251
g19816 and n22250_not n22251 ; n22252
g19817 and n21114_not n22217 ; n22253
g19818 and n6236_not n16992 ; n22254
g19819 nor pi0166 n22254 ; n22255
g19820 and n21055 n22255_not ; n22256
g19821 nor n21074 n22221 ; n22257
g19822 and n2603 n22257 ; n22258
g19823 nor pi0223 n22258 ; n22259
g19824 nor n21415 n22224 ; n22260
g19825 and n21435 n22260_not ; n22261
g19826 and n22259 n22261_not ; n22262
g19827 and n22220 n22256_not ; n22263
g19828 and n22262_not n22263 ; n22264
g19829 nor pi0166 n17037 ; n22265
g19830 and n20998 n22265_not ; n22266
g19831 and n3448 n22257 ; n22267
g19832 nor pi0215 n22267 ; n22268
g19833 and n17032_not n22232 ; n22269
g19834 and n22268 n22269_not ; n22270
g19835 and pi0299 n22266_not ; n22271
g19836 and n22270_not n22271 ; n22272
g19837 and pi0772 n22264_not ; n22273
g19838 and n22272_not n22273 ; n22274
g19839 nor n2603 n22260 ; n22275
g19840 and n2603 n21025 ; n22276
g19841 and n22259 n22276_not ; n22277
g19842 and n22275_not n22277 ; n22278
g19843 nor pi0299 n22256 ; n22279
g19844 and n22278_not n22279 ; n22280
g19845 and n21045_not n22268 ; n22281
g19846 and n22232_not n22281 ; n22282
g19847 and n21400_not n22266 ; n22283
g19848 and pi0299 n22283_not ; n22284
g19849 and n22282_not n22284 ; n22285
g19850 nor pi0772 n22280 ; n22286
g19851 and n22285_not n22286 ; n22287
g19852 and pi0039 n22274_not ; n22288
g19853 and n22287_not n22288 ; n22289
g19854 nor pi0038 n22253 ; n22290
g19855 and n22289_not n22290 ; n22291
g19856 and pi0727 n22252_not ; n22292
g19857 and n22291_not n22292 ; n22293
g19858 nor n22248 n22293 ; n22294
g19859 and n10197 n22294_not ; n22295
g19860 nor pi0832 n22208 ; n22296
g19861 and n22295_not n22296 ; n22297
g19862 nor pi0166 n2926 ; n22298
g19863 and pi0727 n20902 ; n22299
g19864 and n2926 n22210_not ; n22300
g19865 and n22299_not n22300 ; n22301
g19866 and pi0832 n22298_not ; n22302
g19867 and n22301_not n22302 ; n22303
g19868 or n22297 n22303 ; po0323
g19869 nor pi0167 n2926 ; n22305
g19870 and pi0768_not pi0947 ; n22306
g19871 and pi0705 n20902 ; n22307
g19872 nor n22306 n22307 ; n22308
g19873 and n2926 n22308_not ; n22309
g19874 and pi0832 n22305_not ; n22310
g19875 and n22309_not n22310 ; n22311
g19876 nor pi0167 n10197 ; n22312
g19877 and pi0768 n17052_not ; n22313
g19878 and pi0167_not n22313 ; n22314
g19879 nor pi0167 n17050 ; n22315
g19880 nor n21015 n22315 ; n22316
g19881 and pi0167 n21032 ; n22317
g19882 nor pi0167 n21006 ; n22318
g19883 nor pi0038 n22317 ; n22319
g19884 and n22318_not n22319 ; n22320
g19885 nor pi0768 n22316 ; n22321
g19886 and n22320_not n22321 ; n22322
g19887 nor pi0705 n22314 ; n22323
g19888 and n22322_not n22323 ; n22324
g19889 nor pi0167 n16641 ; n22325
g19890 and n21090 n22325_not ; n22326
g19891 and pi0167_not n21099 ; n22327
g19892 and pi0167 n21116 ; n22328
g19893 nor pi0038 n22328 ; n22329
g19894 and n22327_not n22329 ; n22330
g19895 and pi0768 n22326_not ; n22331
g19896 and n22330_not n22331 ; n22332
g19897 nor pi0167 n21039 ; n22333
g19898 and n21042 n22333_not ; n22334
g19899 and pi0167_not n21069 ; n22335
g19900 and pi0167 n21082 ; n22336
g19901 nor pi0038 n22336 ; n22337
g19902 and n22335_not n22337 ; n22338
g19903 nor pi0768 n22334 ; n22339
g19904 and n22338_not n22339 ; n22340
g19905 and pi0705 n22332_not ; n22341
g19906 and n22340_not n22341 ; n22342
g19907 and n10197 n22324_not ; n22343
g19908 and n22342_not n22343 ; n22344
g19909 nor pi0832 n22312 ; n22345
g19910 and n22344_not n22345 ; n22346
g19911 nor n22311 n22346 ; po0324
g19912 and pi0168 n2926_not ; n22348
g19913 and pi0763 pi0947 ; n22349
g19914 and n2926 n22349_not ; n22350
g19915 and pi0699 n20902 ; n22351
g19916 and n22350 n22351_not ; n22352
g19917 and pi0832 n22348_not ; n22353
g19918 and n22352_not n22353 ; n22354
g19919 and pi0057 pi0168 ; n22355
g19920 nor pi0168 n21130 ; n22356
g19921 nor pi0168 n16958 ; n22357
g19922 and pi0763_not n18147 ; n22358
g19923 nor n21017 n22358 ; n22359
g19924 nor n22357 n22359 ; n22360
g19925 and n21114_not n22360 ; n22361
g19926 nor pi0168 n17024 ; n22362
g19927 and n21111 n22362_not ; n22363
g19928 and pi0168 n17037_not ; n22364
g19929 and n20998 n22364_not ; n22365
g19930 and n21073 n22365_not ; n22366
g19931 and pi0168 n3448_not ; n22367
g19932 and n17032_not n22367 ; n22368
g19933 nor n17031 n22368 ; n22369
g19934 nor pi0168 n16653 ; n22370
g19935 and n21105 n22370_not ; n22371
g19936 nor n21047 n22371 ; n22372
g19937 and n22369 n22372 ; n22373
g19938 nor pi0215 n22373 ; n22374
g19939 nor n21021 n22366 ; n22375
g19940 and n22374_not n22375 ; n22376
g19941 and pi0299 n22376_not ; n22377
g19942 nor pi0763 n22363 ; n22378
g19943 and n22377_not n22378 ; n22379
g19944 and n21026 n22370_not ; n22380
g19945 and n21103_not n22380 ; n22381
g19946 nor pi0215 n22381 ; n22382
g19947 and n22369 n22382 ; n22383
g19948 nor n22365 n22383 ; n22384
g19949 and pi0299 n22384_not ; n22385
g19950 and pi0168 n21071_not ; n22386
g19951 and n21062 n22386_not ; n22387
g19952 nor n22385 n22387 ; n22388
g19953 and pi0763 n22388_not ; n22389
g19954 and pi0039 n22379_not ; n22390
g19955 and n22389_not n22390 ; n22391
g19956 nor n22361 n22391 ; n22392
g19957 nor pi0038 n22392 ; n22393
g19958 nor pi0168 n16641 ; n22394
g19959 and pi0763_not pi0947 ; n22395
g19960 nor pi0039 n22395 ; n22396
g19961 and n21239 n22396 ; n22397
g19962 and pi0038 n22394_not ; n22398
g19963 and n22397_not n22398 ; n22399
g19964 nor n22393 n22399 ; n22400
g19965 and pi0699 n22400_not ; n22401
g19966 and n6284 n22350 ; n22402
g19967 and pi0168 n17050_not ; n22403
g19968 and pi0038 n22402_not ; n22404
g19969 and n22403_not n22404 ; n22405
g19970 and n21019 n22362_not ; n22406
g19971 and n21000 n22364_not ; n22407
g19972 and n22369 n22380_not ; n22408
g19973 and n20996 n22408 ; n22409
g19974 and pi0299 n22407_not ; n22410
g19975 and n22409_not n22410 ; n22411
g19976 and pi0763 n22411_not ; n22412
g19977 and n22406_not n22412 ; n22413
g19978 nor pi0168 pi0763 ; n22414
g19979 and n17046_not n22414 ; n22415
g19980 and pi0039 n22415_not ; n22416
g19981 and n22413_not n22416 ; n22417
g19982 nor pi0038 n22360 ; n22418
g19983 and n22417_not n22418 ; n22419
g19984 nor pi0699 n22405 ; n22420
g19985 and n22419_not n22420 ; n22421
g19986 and n21130 n22421_not ; n22422
g19987 and n22401_not n22422 ; n22423
g19988 nor pi0057 n22356 ; n22424
g19989 and n22423_not n22424 ; n22425
g19990 nor pi0832 n22355 ; n22426
g19991 and n22425_not n22426 ; n22427
g19992 or n22354 n22427 ; po0325
g19993 and pi0169 n2926_not ; n22429
g19994 and pi0746 pi0947 ; n22430
g19995 and n2926 n22430_not ; n22431
g19996 and pi0729 n20902 ; n22432
g19997 and n22431 n22432_not ; n22433
g19998 and pi0832 n22429_not ; n22434
g19999 and n22433_not n22434 ; n22435
g20000 and pi0057 pi0169 ; n22436
g20001 nor pi0169 n21130 ; n22437
g20002 nor pi0169 n16958 ; n22438
g20003 and pi0746_not n18147 ; n22439
g20004 nor n21017 n22439 ; n22440
g20005 nor n22438 n22440 ; n22441
g20006 and n21114_not n22441 ; n22442
g20007 nor pi0169 n17024 ; n22443
g20008 and n21111 n22443_not ; n22444
g20009 and pi0169 n17037_not ; n22445
g20010 and n20998 n22445_not ; n22446
g20011 and n21073 n22446_not ; n22447
g20012 and pi0169 n3448_not ; n22448
g20013 and n17032_not n22448 ; n22449
g20014 nor n17031 n22449 ; n22450
g20015 nor pi0169 n16653 ; n22451
g20016 and n21105 n22451_not ; n22452
g20017 nor n21047 n22452 ; n22453
g20018 and n22450 n22453 ; n22454
g20019 nor pi0215 n22454 ; n22455
g20020 nor n21021 n22447 ; n22456
g20021 and n22455_not n22456 ; n22457
g20022 and pi0299 n22457_not ; n22458
g20023 nor pi0746 n22444 ; n22459
g20024 and n22458_not n22459 ; n22460
g20025 and n21026 n22451_not ; n22461
g20026 and n21103_not n22461 ; n22462
g20027 nor pi0215 n22462 ; n22463
g20028 and n22450 n22463 ; n22464
g20029 nor n22446 n22464 ; n22465
g20030 and pi0299 n22465_not ; n22466
g20031 and pi0169 n21071_not ; n22467
g20032 and n21062 n22467_not ; n22468
g20033 nor n22466 n22468 ; n22469
g20034 and pi0746 n22469_not ; n22470
g20035 and pi0039 n22460_not ; n22471
g20036 and n22470_not n22471 ; n22472
g20037 nor n22442 n22472 ; n22473
g20038 nor pi0038 n22473 ; n22474
g20039 nor pi0169 n16641 ; n22475
g20040 and pi0746_not pi0947 ; n22476
g20041 nor pi0039 n22476 ; n22477
g20042 and n21239 n22477 ; n22478
g20043 and pi0038 n22475_not ; n22479
g20044 and n22478_not n22479 ; n22480
g20045 nor n22474 n22480 ; n22481
g20046 and pi0729 n22481_not ; n22482
g20047 and n6284 n22431 ; n22483
g20048 and pi0169 n17050_not ; n22484
g20049 and pi0038 n22483_not ; n22485
g20050 and n22484_not n22485 ; n22486
g20051 and n21019 n22443_not ; n22487
g20052 and n21000 n22445_not ; n22488
g20053 and n22450 n22461_not ; n22489
g20054 and n20996 n22489 ; n22490
g20055 and pi0299 n22488_not ; n22491
g20056 and n22490_not n22491 ; n22492
g20057 and pi0746 n22492_not ; n22493
g20058 and n22487_not n22493 ; n22494
g20059 nor pi0169 pi0746 ; n22495
g20060 and n17046_not n22495 ; n22496
g20061 and pi0039 n22496_not ; n22497
g20062 and n22494_not n22497 ; n22498
g20063 nor pi0038 n22441 ; n22499
g20064 and n22498_not n22499 ; n22500
g20065 nor pi0729 n22486 ; n22501
g20066 and n22500_not n22501 ; n22502
g20067 and n21130 n22502_not ; n22503
g20068 and n22482_not n22503 ; n22504
g20069 nor pi0057 n22437 ; n22505
g20070 and n22504_not n22505 ; n22506
g20071 nor pi0832 n22436 ; n22507
g20072 and n22506_not n22507 ; n22508
g20073 or n22435 n22508 ; po0326
g20074 and pi0730 n20902 ; n22510
g20075 and pi0748 pi0947 ; n22511
g20076 and n2926 n22511_not ; n22512
g20077 and n22510_not n22512 ; n22513
g20078 and pi0170 n2926_not ; n22514
g20079 and pi0832 n22514_not ; n22515
g20080 and n22513_not n22515 ; n22516
g20081 and pi0057 pi0170 ; n22517
g20082 nor pi0170 n21130 ; n22518
g20083 nor pi0170 n16641 ; n22519
g20084 and n21090 n22519_not ; n22520
g20085 and pi0170 n17037_not ; n22521
g20086 and n20998 n22521_not ; n22522
g20087 and n21073 n22522_not ; n22523
g20088 and pi0170 n3448_not ; n22524
g20089 and n17032_not n22524 ; n22525
g20090 nor n17031 n22525 ; n22526
g20091 nor pi0170 n16653 ; n22527
g20092 and n21105 n22527_not ; n22528
g20093 nor n21047 n22528 ; n22529
g20094 and n22526 n22529 ; n22530
g20095 nor pi0215 n22530 ; n22531
g20096 nor n21021 n22523 ; n22532
g20097 and n22531_not n22532 ; n22533
g20098 and pi0299 n22533_not ; n22534
g20099 nor pi0170 n17024 ; n22535
g20100 nor pi0299 n22535 ; n22536
g20101 and n21110_not n22536 ; n22537
g20102 nor n22534 n22537 ; n22538
g20103 and pi0039 n22538_not ; n22539
g20104 nor pi0170 n16958 ; n22540
g20105 and n21115 n22540_not ; n22541
g20106 nor n22539 n22541 ; n22542
g20107 nor pi0038 n22542 ; n22543
g20108 nor pi0748 n22520 ; n22544
g20109 and n22543_not n22544 ; n22545
g20110 and n21042 n22519_not ; n22546
g20111 and n21067 n22540_not ; n22547
g20112 and n21026 n22527_not ; n22548
g20113 and n21103_not n22548 ; n22549
g20114 nor pi0215 n22549 ; n22550
g20115 and n22526 n22550 ; n22551
g20116 nor n22522 n22551 ; n22552
g20117 and pi0299 n22552_not ; n22553
g20118 and pi0170 n21071_not ; n22554
g20119 and n21062 n22554_not ; n22555
g20120 and pi0039 n22553_not ; n22556
g20121 and n22555_not n22556 ; n22557
g20122 nor n22547 n22557 ; n22558
g20123 nor pi0038 n22558 ; n22559
g20124 and pi0748 n22546_not ; n22560
g20125 and n22559_not n22560 ; n22561
g20126 and pi0730 n22561_not ; n22562
g20127 and n22545_not n22562 ; n22563
g20128 nor pi0170 n17050 ; n22564
g20129 nor n21015 n22564 ; n22565
g20130 and n21017 n22540_not ; n22566
g20131 and n21000 n22521_not ; n22567
g20132 and n22526 n22548_not ; n22568
g20133 and n20996 n22568 ; n22569
g20134 and pi0299 n22567_not ; n22570
g20135 and n22569_not n22570 ; n22571
g20136 and n21018_not n22536 ; n22572
g20137 nor n22571 n22572 ; n22573
g20138 and pi0039 n22573_not ; n22574
g20139 nor n22566 n22574 ; n22575
g20140 nor pi0038 n22575 ; n22576
g20141 and pi0748 n22565_not ; n22577
g20142 and n22576_not n22577 ; n22578
g20143 nor pi0170 pi0748 ; n22579
g20144 and n17052_not n22579 ; n22580
g20145 nor pi0730 n22580 ; n22581
g20146 and n22578_not n22581 ; n22582
g20147 and n21130 n22582_not ; n22583
g20148 and n22563_not n22583 ; n22584
g20149 nor pi0057 n22518 ; n22585
g20150 and n22584_not n22585 ; n22586
g20151 nor pi0832 n22517 ; n22587
g20152 and n22586_not n22587 ; n22588
g20153 or n22516 n22588 ; po0327
g20154 and pi0171 n2926_not ; n22590
g20155 and pi0764 pi0947 ; n22591
g20156 and n2926 n22591_not ; n22592
g20157 and pi0691 n20902 ; n22593
g20158 and n22592 n22593_not ; n22594
g20159 and pi0832 n22590_not ; n22595
g20160 and n22594_not n22595 ; n22596
g20161 and pi0057 pi0171 ; n22597
g20162 nor pi0171 n21130 ; n22598
g20163 nor pi0171 n16958 ; n22599
g20164 and pi0764_not n18147 ; n22600
g20165 nor n21017 n22600 ; n22601
g20166 nor n22599 n22601 ; n22602
g20167 and n21114_not n22602 ; n22603
g20168 nor pi0171 n17024 ; n22604
g20169 and n21111 n22604_not ; n22605
g20170 and pi0171 n17037_not ; n22606
g20171 and n20998 n22606_not ; n22607
g20172 and n21073 n22607_not ; n22608
g20173 and pi0171 n3448_not ; n22609
g20174 and n17032_not n22609 ; n22610
g20175 nor n17031 n22610 ; n22611
g20176 nor pi0171 n16653 ; n22612
g20177 and n21105 n22612_not ; n22613
g20178 nor n21047 n22613 ; n22614
g20179 and n22611 n22614 ; n22615
g20180 nor pi0215 n22615 ; n22616
g20181 nor n21021 n22608 ; n22617
g20182 and n22616_not n22617 ; n22618
g20183 and pi0299 n22618_not ; n22619
g20184 nor pi0764 n22605 ; n22620
g20185 and n22619_not n22620 ; n22621
g20186 and n21026 n22612_not ; n22622
g20187 and n21103_not n22622 ; n22623
g20188 nor pi0215 n22623 ; n22624
g20189 and n22611 n22624 ; n22625
g20190 nor n22607 n22625 ; n22626
g20191 and pi0299 n22626_not ; n22627
g20192 and pi0171 n21071_not ; n22628
g20193 and n21062 n22628_not ; n22629
g20194 nor n22627 n22629 ; n22630
g20195 and pi0764 n22630_not ; n22631
g20196 and pi0039 n22621_not ; n22632
g20197 and n22631_not n22632 ; n22633
g20198 nor n22603 n22633 ; n22634
g20199 nor pi0038 n22634 ; n22635
g20200 nor pi0171 n16641 ; n22636
g20201 and pi0764_not pi0947 ; n22637
g20202 nor pi0039 n22637 ; n22638
g20203 and n21239 n22638 ; n22639
g20204 and pi0038 n22636_not ; n22640
g20205 and n22639_not n22640 ; n22641
g20206 nor n22635 n22641 ; n22642
g20207 and pi0691 n22642_not ; n22643
g20208 and n6284 n22592 ; n22644
g20209 and pi0171 n17050_not ; n22645
g20210 and pi0038 n22644_not ; n22646
g20211 and n22645_not n22646 ; n22647
g20212 and n21019 n22604_not ; n22648
g20213 and n21000 n22606_not ; n22649
g20214 and n22611 n22622_not ; n22650
g20215 and n20996 n22650 ; n22651
g20216 and pi0299 n22649_not ; n22652
g20217 and n22651_not n22652 ; n22653
g20218 and pi0764 n22653_not ; n22654
g20219 and n22648_not n22654 ; n22655
g20220 nor pi0171 pi0764 ; n22656
g20221 and n17046_not n22656 ; n22657
g20222 and pi0039 n22657_not ; n22658
g20223 and n22655_not n22658 ; n22659
g20224 nor pi0038 n22602 ; n22660
g20225 and n22659_not n22660 ; n22661
g20226 nor pi0691 n22647 ; n22662
g20227 and n22661_not n22662 ; n22663
g20228 and n21130 n22663_not ; n22664
g20229 and n22643_not n22664 ; n22665
g20230 nor pi0057 n22598 ; n22666
g20231 and n22665_not n22666 ; n22667
g20232 nor pi0832 n22597 ; n22668
g20233 and n22667_not n22668 ; n22669
g20234 or n22596 n22669 ; po0328
g20235 and pi0172 n2926_not ; n22671
g20236 and pi0739 pi0947 ; n22672
g20237 and n2926 n22672_not ; n22673
g20238 and pi0690 n20902 ; n22674
g20239 and n22673 n22674_not ; n22675
g20240 and pi0832 n22671_not ; n22676
g20241 and n22675_not n22676 ; n22677
g20242 and pi0057 pi0172 ; n22678
g20243 nor pi0172 n21130 ; n22679
g20244 nor pi0172 n16958 ; n22680
g20245 and n16958 n22672 ; n22681
g20246 nor pi0039 n22680 ; n22682
g20247 and n22681_not n22682 ; n22683
g20248 and n21114_not n22683 ; n22684
g20249 nor pi0172 n17024 ; n22685
g20250 and n21111 n22685_not ; n22686
g20251 and pi0172 n17037_not ; n22687
g20252 and n20998 n22687_not ; n22688
g20253 and n21073 n22688_not ; n22689
g20254 and pi0172 n3448_not ; n22690
g20255 and n17032_not n22690 ; n22691
g20256 nor n17031 n22691 ; n22692
g20257 nor pi0172 n16653 ; n22693
g20258 and n21105 n22693_not ; n22694
g20259 nor n21047 n22694 ; n22695
g20260 and n22692 n22695 ; n22696
g20261 nor pi0215 n22696 ; n22697
g20262 nor n21021 n22689 ; n22698
g20263 and n22697_not n22698 ; n22699
g20264 and pi0299 n22699_not ; n22700
g20265 nor pi0739 n22686 ; n22701
g20266 and n22700_not n22701 ; n22702
g20267 and n21026 n22693_not ; n22703
g20268 and n21103_not n22703 ; n22704
g20269 nor pi0215 n22704 ; n22705
g20270 and n22692 n22705 ; n22706
g20271 nor n22688 n22706 ; n22707
g20272 and pi0299 n22707_not ; n22708
g20273 and pi0172 n21071_not ; n22709
g20274 and n21062 n22709_not ; n22710
g20275 nor n22708 n22710 ; n22711
g20276 and pi0739 n22711_not ; n22712
g20277 and pi0039 n22702_not ; n22713
g20278 and n22712_not n22713 ; n22714
g20279 nor n22684 n22714 ; n22715
g20280 nor pi0038 n22715 ; n22716
g20281 nor pi0172 n16641 ; n22717
g20282 and pi0739_not pi0947 ; n22718
g20283 nor pi0039 n22718 ; n22719
g20284 and n21239 n22719 ; n22720
g20285 and pi0038 n22717_not ; n22721
g20286 and n22720_not n22721 ; n22722
g20287 nor n22716 n22722 ; n22723
g20288 and pi0690 n22723_not ; n22724
g20289 and n6284 n22673 ; n22725
g20290 and pi0172 n17050_not ; n22726
g20291 and pi0038 n22725_not ; n22727
g20292 and n22726_not n22727 ; n22728
g20293 and n21019 n22685_not ; n22729
g20294 and n21000 n22687_not ; n22730
g20295 and n22692 n22703_not ; n22731
g20296 and n20996 n22731 ; n22732
g20297 and pi0299 n22730_not ; n22733
g20298 and n22732_not n22733 ; n22734
g20299 and pi0739 n22734_not ; n22735
g20300 and n22729_not n22735 ; n22736
g20301 nor pi0172 pi0739 ; n22737
g20302 and n17046_not n22737 ; n22738
g20303 and pi0039 n22738_not ; n22739
g20304 and n22736_not n22739 ; n22740
g20305 nor pi0038 n22683 ; n22741
g20306 and n22740_not n22741 ; n22742
g20307 nor pi0690 n22728 ; n22743
g20308 and n22742_not n22743 ; n22744
g20309 and n21130 n22744_not ; n22745
g20310 and n22724_not n22745 ; n22746
g20311 nor pi0057 n22679 ; n22747
g20312 and n22746_not n22747 ; n22748
g20313 nor pi0832 n22678 ; n22749
g20314 and n22748_not n22749 ; n22750
g20315 or n22677 n22750 ; po0329
g20316 and pi0173_not po1038 ; n22752
g20317 nor pi0173 n17059 ; n22753
g20318 and n16635 n22753_not ; n22754
g20319 and pi0723_not n2571 ; n22755
g20320 and n22753 n22755_not ; n22756
g20321 nor pi0173 n16641 ; n22757
g20322 and n16647 n22757_not ; n22758
g20323 and pi0173 n18076_not ; n22759
g20324 nor pi0038 n22759 ; n22760
g20325 and n2571 n22760_not ; n22761
g20326 and pi0173_not n18072 ; n22762
g20327 nor n22761 n22762 ; n22763
g20328 nor pi0723 n22758 ; n22764
g20329 and n22763_not n22764 ; n22765
g20330 nor n22756 n22765 ; n22766
g20331 and pi0778_not n22766 ; n22767
g20332 and pi0625_not n22753 ; n22768
g20333 and pi0625 n22766_not ; n22769
g20334 and pi1153 n22768_not ; n22770
g20335 and n22769_not n22770 ; n22771
g20336 and pi0625 n22753 ; n22772
g20337 nor pi0625 n22766 ; n22773
g20338 nor pi1153 n22772 ; n22774
g20339 and n22773_not n22774 ; n22775
g20340 nor n22771 n22775 ; n22776
g20341 and pi0778 n22776_not ; n22777
g20342 nor n22767 n22777 ; n22778
g20343 nor n17075 n22778 ; n22779
g20344 and n17075 n22753_not ; n22780
g20345 nor n22779 n22780 ; n22781
g20346 and n16639_not n22781 ; n22782
g20347 and n16639 n22753 ; n22783
g20348 nor n22782 n22783 ; n22784
g20349 and n16635_not n22784 ; n22785
g20350 nor n22754 n22785 ; n22786
g20351 and n16631_not n22786 ; n22787
g20352 and n16631 n22753 ; n22788
g20353 nor n22787 n22788 ; n22789
g20354 and pi0792_not n22789 ; n22790
g20355 and pi0628 n22789_not ; n22791
g20356 and pi0628_not n22753 ; n22792
g20357 and pi1156 n22792_not ; n22793
g20358 and n22791_not n22793 ; n22794
g20359 and pi0628 n22753 ; n22795
g20360 nor pi0628 n22789 ; n22796
g20361 nor pi1156 n22795 ; n22797
g20362 and n22796_not n22797 ; n22798
g20363 nor n22794 n22798 ; n22799
g20364 and pi0792 n22799_not ; n22800
g20365 nor n22790 n22800 ; n22801
g20366 nor pi0647 n22801 ; n22802
g20367 and pi0647 n22753_not ; n22803
g20368 nor n22802 n22803 ; n22804
g20369 and pi1157_not n22804 ; n22805
g20370 and pi0647 n22801_not ; n22806
g20371 nor pi0647 n22753 ; n22807
g20372 nor n22806 n22807 ; n22808
g20373 and pi1157 n22808 ; n22809
g20374 nor n22805 n22809 ; n22810
g20375 and pi0787 n22810_not ; n22811
g20376 and pi0787_not n22801 ; n22812
g20377 nor n22811 n22812 ; n22813
g20378 nor pi0644 n22813 ; n22814
g20379 and pi0715 n22814_not ; n22815
g20380 and pi0173 n2571_not ; n22816
g20381 and pi0173 n17275_not ; n22817
g20382 nor pi0173 n17048 ; n22818
g20383 and pi0745 n22818_not ; n22819
g20384 nor pi0173 pi0745 ; n22820
g20385 and n17221 n22820 ; n22821
g20386 nor n22817 n22821 ; n22822
g20387 and n22819_not n22822 ; n22823
g20388 nor pi0038 n22823 ; n22824
g20389 and pi0745_not n17280 ; n22825
g20390 and pi0038 n22757_not ; n22826
g20391 and n22825_not n22826 ; n22827
g20392 nor n22824 n22827 ; n22828
g20393 and n2571 n22828_not ; n22829
g20394 nor n22816 n22829 ; n22830
g20395 nor n17117 n22830 ; n22831
g20396 and n17117 n22753_not ; n22832
g20397 nor n22831 n22832 ; n22833
g20398 nor pi0785 n22833 ; n22834
g20399 nor n17291 n22753 ; n22835
g20400 and pi0609 n22831 ; n22836
g20401 nor n22835 n22836 ; n22837
g20402 and pi1155 n22837_not ; n22838
g20403 nor n17296 n22753 ; n22839
g20404 and pi0609_not n22831 ; n22840
g20405 nor n22839 n22840 ; n22841
g20406 nor pi1155 n22841 ; n22842
g20407 nor n22838 n22842 ; n22843
g20408 and pi0785 n22843_not ; n22844
g20409 nor n22834 n22844 ; n22845
g20410 nor pi0781 n22845 ; n22846
g20411 and pi0618_not n22753 ; n22847
g20412 and pi0618 n22845 ; n22848
g20413 and pi1154 n22847_not ; n22849
g20414 and n22848_not n22849 ; n22850
g20415 and pi0618_not n22845 ; n22851
g20416 and pi0618 n22753 ; n22852
g20417 nor pi1154 n22852 ; n22853
g20418 and n22851_not n22853 ; n22854
g20419 nor n22850 n22854 ; n22855
g20420 and pi0781 n22855_not ; n22856
g20421 nor n22846 n22856 ; n22857
g20422 nor pi0789 n22857 ; n22858
g20423 and pi0619_not n22753 ; n22859
g20424 and pi0619 n22857 ; n22860
g20425 and pi1159 n22859_not ; n22861
g20426 and n22860_not n22861 ; n22862
g20427 and pi0619_not n22857 ; n22863
g20428 and pi0619 n22753 ; n22864
g20429 nor pi1159 n22864 ; n22865
g20430 and n22863_not n22865 ; n22866
g20431 nor n22862 n22866 ; n22867
g20432 and pi0789 n22867_not ; n22868
g20433 nor n22858 n22868 ; n22869
g20434 nor pi0788 n22869 ; n22870
g20435 and pi0626_not n22753 ; n22871
g20436 and pi0626 n22869 ; n22872
g20437 and pi1158 n22871_not ; n22873
g20438 and n22872_not n22873 ; n22874
g20439 and pi0626_not n22869 ; n22875
g20440 and pi0626 n22753 ; n22876
g20441 nor pi1158 n22876 ; n22877
g20442 and n22875_not n22877 ; n22878
g20443 nor n22874 n22878 ; n22879
g20444 and pi0788 n22879_not ; n22880
g20445 nor n22870 n22880 ; n22881
g20446 and n17779_not n22881 ; n22882
g20447 and n17779 n22753 ; n22883
g20448 nor n22882 n22883 ; n22884
g20449 nor n17804 n22884 ; n22885
g20450 and n17804 n22753 ; n22886
g20451 nor n22885 n22886 ; n22887
g20452 and pi0644 n22887_not ; n22888
g20453 and pi0644_not n22753 ; n22889
g20454 nor pi0715 n22889 ; n22890
g20455 and n22888_not n22890 ; n22891
g20456 and pi1160 n22891_not ; n22892
g20457 and n22815_not n22892 ; n22893
g20458 and pi0644 n22813_not ; n22894
g20459 and n17802 n22804_not ; n22895
g20460 and n20559_not n22884 ; n22896
g20461 and n17801 n22808_not ; n22897
g20462 nor n22895 n22897 ; n22898
g20463 and n22896_not n22898 ; n22899
g20464 and pi0787 n22899_not ; n22900
g20465 and pi0629_not n22794 ; n22901
g20466 nor n20570 n22881 ; n22902
g20467 and pi0629 n22798 ; n22903
g20468 nor n22901 n22903 ; n22904
g20469 and n22902_not n22904 ; n22905
g20470 and pi0792 n22905_not ; n22906
g20471 and pi0609 n22778 ; n22907
g20472 and pi0173 n17625_not ; n22908
g20473 nor pi0173 n17612 ; n22909
g20474 and pi0745 n22908_not ; n22910
g20475 and n22909_not n22910 ; n22911
g20476 and pi0173_not n17629 ; n22912
g20477 and pi0173 n17631 ; n22913
g20478 nor pi0745 n22913 ; n22914
g20479 and n22912_not n22914 ; n22915
g20480 nor n22911 n22915 ; n22916
g20481 nor pi0039 n22916 ; n22917
g20482 and pi0173 n17605 ; n22918
g20483 nor pi0173 n17546 ; n22919
g20484 nor pi0745 n22919 ; n22920
g20485 and n22918_not n22920 ; n22921
g20486 and pi0173_not n17404 ; n22922
g20487 and pi0173 n17485 ; n22923
g20488 and pi0745 n22923_not ; n22924
g20489 and n22922_not n22924 ; n22925
g20490 and pi0039 n22921_not ; n22926
g20491 and n22925_not n22926 ; n22927
g20492 nor pi0038 n22917 ; n22928
g20493 and n22927_not n22928 ; n22929
g20494 nor pi0745 n17490 ; n22930
g20495 and n19471 n22930_not ; n22931
g20496 nor pi0173 n22931 ; n22932
g20497 and pi0745_not n17244 ; n22933
g20498 nor n17469 n22933 ; n22934
g20499 and pi0173 n22934_not ; n22935
g20500 and n6284 n22935 ; n22936
g20501 and pi0038 n22936_not ; n22937
g20502 and n22932_not n22937 ; n22938
g20503 nor pi0723 n22938 ; n22939
g20504 and n22929_not n22939 ; n22940
g20505 and pi0723 n22828 ; n22941
g20506 and n2571 n22940_not ; n22942
g20507 and n22941_not n22942 ; n22943
g20508 nor n22816 n22943 ; n22944
g20509 and pi0625_not n22944 ; n22945
g20510 and pi0625 n22830 ; n22946
g20511 nor pi1153 n22946 ; n22947
g20512 and n22945_not n22947 ; n22948
g20513 nor pi0608 n22771 ; n22949
g20514 and n22948_not n22949 ; n22950
g20515 and pi0625_not n22830 ; n22951
g20516 and pi0625 n22944 ; n22952
g20517 and pi1153 n22951_not ; n22953
g20518 and n22952_not n22953 ; n22954
g20519 and pi0608 n22775_not ; n22955
g20520 and n22954_not n22955 ; n22956
g20521 nor n22950 n22956 ; n22957
g20522 and pi0778 n22957_not ; n22958
g20523 and pi0778_not n22944 ; n22959
g20524 nor n22958 n22959 ; n22960
g20525 nor pi0609 n22960 ; n22961
g20526 nor pi1155 n22907 ; n22962
g20527 and n22961_not n22962 ; n22963
g20528 nor pi0660 n22838 ; n22964
g20529 and n22963_not n22964 ; n22965
g20530 and pi0609_not n22778 ; n22966
g20531 and pi0609 n22960_not ; n22967
g20532 and pi1155 n22966_not ; n22968
g20533 and n22967_not n22968 ; n22969
g20534 and pi0660 n22842_not ; n22970
g20535 and n22969_not n22970 ; n22971
g20536 nor n22965 n22971 ; n22972
g20537 and pi0785 n22972_not ; n22973
g20538 nor pi0785 n22960 ; n22974
g20539 nor n22973 n22974 ; n22975
g20540 nor pi0618 n22975 ; n22976
g20541 and pi0618 n22781 ; n22977
g20542 nor pi1154 n22977 ; n22978
g20543 and n22976_not n22978 ; n22979
g20544 nor pi0627 n22850 ; n22980
g20545 and n22979_not n22980 ; n22981
g20546 and pi0618_not n22781 ; n22982
g20547 and pi0618 n22975_not ; n22983
g20548 and pi1154 n22982_not ; n22984
g20549 and n22983_not n22984 ; n22985
g20550 and pi0627 n22854_not ; n22986
g20551 and n22985_not n22986 ; n22987
g20552 nor n22981 n22987 ; n22988
g20553 and pi0781 n22988_not ; n22989
g20554 nor pi0781 n22975 ; n22990
g20555 nor n22989 n22990 ; n22991
g20556 and pi0789_not n22991 ; n22992
g20557 and pi0619 n22784_not ; n22993
g20558 nor pi0619 n22991 ; n22994
g20559 nor pi1159 n22993 ; n22995
g20560 and n22994_not n22995 ; n22996
g20561 nor pi0648 n22862 ; n22997
g20562 and n22996_not n22997 ; n22998
g20563 and pi0619 n22991_not ; n22999
g20564 nor pi0619 n22784 ; n23000
g20565 and pi1159 n23000_not ; n23001
g20566 and n22999_not n23001 ; n23002
g20567 and pi0648 n22866_not ; n23003
g20568 and n23002_not n23003 ; n23004
g20569 and pi0789 n22998_not ; n23005
g20570 and n23004_not n23005 ; n23006
g20571 and n17970 n22992_not ; n23007
g20572 and n23006_not n23007 ; n23008
g20573 and n17871 n22786 ; n23009
g20574 and n16630_not n22879 ; n23010
g20575 nor n23009 n23010 ; n23011
g20576 and pi0788 n23011_not ; n23012
g20577 nor n20364 n23012 ; n23013
g20578 and n23008_not n23013 ; n23014
g20579 nor n22906 n23014 ; n23015
g20580 nor n20206 n23015 ; n23016
g20581 nor n22900 n23016 ; n23017
g20582 and pi0644_not n23017 ; n23018
g20583 nor pi0715 n22894 ; n23019
g20584 and n23018_not n23019 ; n23020
g20585 and pi0644 n22753 ; n23021
g20586 nor pi0644 n22887 ; n23022
g20587 and pi0715 n23021_not ; n23023
g20588 and n23022_not n23023 ; n23024
g20589 nor pi1160 n23024 ; n23025
g20590 and n23020_not n23025 ; n23026
g20591 nor n22893 n23026 ; n23027
g20592 and pi0790 n23027_not ; n23028
g20593 and pi0644 n22892 ; n23029
g20594 and pi0790 n23029_not ; n23030
g20595 and n23017 n23030_not ; n23031
g20596 nor n23028 n23031 ; n23032
g20597 nor po1038 n23032 ; n23033
g20598 nor pi0832 n22752 ; n23034
g20599 and n23033_not n23034 ; n23035
g20600 nor pi0173 n2926 ; n23036
g20601 and pi0723_not n16645 ; n23037
g20602 nor n23036 n23037 ; n23038
g20603 nor pi0778 n23038 ; n23039
g20604 and pi0625_not n23037 ; n23040
g20605 nor n23038 n23040 ; n23041
g20606 and pi1153 n23041_not ; n23042
g20607 nor pi1153 n23036 ; n23043
g20608 and n23040_not n23043 ; n23044
g20609 and pi0778 n23044_not ; n23045
g20610 and n23042_not n23045 ; n23046
g20611 nor n23039 n23046 ; n23047
g20612 nor n17845 n23047 ; n23048
g20613 and n17847_not n23048 ; n23049
g20614 and n17849_not n23049 ; n23050
g20615 and n17851_not n23050 ; n23051
g20616 and n17857_not n23051 ; n23052
g20617 and pi0647_not n23052 ; n23053
g20618 and pi0647 n23036 ; n23054
g20619 nor pi1157 n23054 ; n23055
g20620 and n23053_not n23055 ; n23056
g20621 and pi0630 n23056 ; n23057
g20622 nor n22933 n23036 ; n23058
g20623 nor n17874 n23058 ; n23059
g20624 nor pi0785 n23059 ; n23060
g20625 and n17296 n22933 ; n23061
g20626 and n23059 n23061_not ; n23062
g20627 and pi1155 n23062_not ; n23063
g20628 nor pi1155 n23036 ; n23064
g20629 and n23061_not n23064 ; n23065
g20630 nor n23063 n23065 ; n23066
g20631 and pi0785 n23066_not ; n23067
g20632 nor n23060 n23067 ; n23068
g20633 nor pi0781 n23068 ; n23069
g20634 and n17889_not n23068 ; n23070
g20635 and pi1154 n23070_not ; n23071
g20636 and n17892_not n23068 ; n23072
g20637 nor pi1154 n23072 ; n23073
g20638 nor n23071 n23073 ; n23074
g20639 and pi0781 n23074_not ; n23075
g20640 nor n23069 n23075 ; n23076
g20641 nor pi0789 n23076 ; n23077
g20642 and pi0619_not n2926 ; n23078
g20643 and n23076 n23078_not ; n23079
g20644 and pi1159 n23079_not ; n23080
g20645 and pi0619 n2926 ; n23081
g20646 and n23076 n23081_not ; n23082
g20647 nor pi1159 n23082 ; n23083
g20648 nor n23080 n23083 ; n23084
g20649 and pi0789 n23084_not ; n23085
g20650 nor n23077 n23085 ; n23086
g20651 nor pi0788 n23086 ; n23087
g20652 and pi0626_not n23036 ; n23088
g20653 and pi0626 n23086 ; n23089
g20654 and pi1158 n23088_not ; n23090
g20655 and n23089_not n23090 ; n23091
g20656 and pi0626_not n23086 ; n23092
g20657 and pi0626 n23036 ; n23093
g20658 nor pi1158 n23093 ; n23094
g20659 and n23092_not n23094 ; n23095
g20660 nor n23091 n23095 ; n23096
g20661 and pi0788 n23096_not ; n23097
g20662 nor n23087 n23097 ; n23098
g20663 and n17779_not n23098 ; n23099
g20664 and n17779 n23036 ; n23100
g20665 nor n23099 n23100 ; n23101
g20666 and n20559_not n23101 ; n23102
g20667 and pi0647 n23052_not ; n23103
g20668 nor pi0647 n23036 ; n23104
g20669 nor n23103 n23104 ; n23105
g20670 and n17801 n23105_not ; n23106
g20671 nor n23057 n23106 ; n23107
g20672 and n23102_not n23107 ; n23108
g20673 and pi0787 n23108_not ; n23109
g20674 and n17871 n23050 ; n23110
g20675 and n16630_not n23096 ; n23111
g20676 nor n23110 n23111 ; n23112
g20677 and pi0788 n23112_not ; n23113
g20678 and pi0618 n23048 ; n23114
g20679 nor n17168 n23038 ; n23115
g20680 and pi0625 n23115 ; n23116
g20681 and n23058 n23115_not ; n23117
g20682 nor n23116 n23117 ; n23118
g20683 and n23043 n23118_not ; n23119
g20684 nor pi0608 n23042 ; n23120
g20685 and n23119_not n23120 ; n23121
g20686 and pi1153 n23058 ; n23122
g20687 and n23116_not n23122 ; n23123
g20688 and pi0608 n23044_not ; n23124
g20689 and n23123_not n23124 ; n23125
g20690 nor n23121 n23125 ; n23126
g20691 and pi0778 n23126_not ; n23127
g20692 nor pi0778 n23117 ; n23128
g20693 nor n23127 n23128 ; n23129
g20694 nor pi0609 n23129 ; n23130
g20695 and pi0609 n23047_not ; n23131
g20696 nor pi1155 n23131 ; n23132
g20697 and n23130_not n23132 ; n23133
g20698 nor pi0660 n23063 ; n23134
g20699 and n23133_not n23134 ; n23135
g20700 and pi0609 n23129_not ; n23136
g20701 nor pi0609 n23047 ; n23137
g20702 and pi1155 n23137_not ; n23138
g20703 and n23136_not n23138 ; n23139
g20704 and pi0660 n23065_not ; n23140
g20705 and n23139_not n23140 ; n23141
g20706 nor n23135 n23141 ; n23142
g20707 and pi0785 n23142_not ; n23143
g20708 nor pi0785 n23129 ; n23144
g20709 nor n23143 n23144 ; n23145
g20710 nor pi0618 n23145 ; n23146
g20711 nor pi1154 n23114 ; n23147
g20712 and n23146_not n23147 ; n23148
g20713 nor pi0627 n23071 ; n23149
g20714 and n23148_not n23149 ; n23150
g20715 and pi0618_not n23048 ; n23151
g20716 and pi0618 n23145_not ; n23152
g20717 and pi1154 n23151_not ; n23153
g20718 and n23152_not n23153 ; n23154
g20719 and pi0627 n23073_not ; n23155
g20720 and n23154_not n23155 ; n23156
g20721 nor n23150 n23156 ; n23157
g20722 and pi0781 n23157_not ; n23158
g20723 nor pi0781 n23145 ; n23159
g20724 nor n23158 n23159 ; n23160
g20725 and pi0789_not n23160 ; n23161
g20726 nor pi0619 n23160 ; n23162
g20727 and pi0619 n23049 ; n23163
g20728 nor pi1159 n23163 ; n23164
g20729 and n23162_not n23164 ; n23165
g20730 nor pi0648 n23080 ; n23166
g20731 and n23165_not n23166 ; n23167
g20732 and pi0619_not n23049 ; n23168
g20733 and pi0619 n23160_not ; n23169
g20734 and pi1159 n23168_not ; n23170
g20735 and n23169_not n23170 ; n23171
g20736 and pi0648 n23083_not ; n23172
g20737 and n23171_not n23172 ; n23173
g20738 and pi0789 n23167_not ; n23174
g20739 and n23173_not n23174 ; n23175
g20740 and n17970 n23161_not ; n23176
g20741 and n23175_not n23176 ; n23177
g20742 nor n23113 n23177 ; n23178
g20743 nor n20364 n23178 ; n23179
g20744 and n17854 n23098 ; n23180
g20745 and n20851 n23051 ; n23181
g20746 nor n23180 n23181 ; n23182
g20747 nor pi0629 n23182 ; n23183
g20748 and n20855 n23051 ; n23184
g20749 and n17853 n23098 ; n23185
g20750 nor n23184 n23185 ; n23186
g20751 and pi0629 n23186_not ; n23187
g20752 nor n23183 n23187 ; n23188
g20753 and pi0792 n23188_not ; n23189
g20754 nor n20206 n23189 ; n23190
g20755 and n23179_not n23190 ; n23191
g20756 nor n23109 n23191 ; n23192
g20757 and pi0790_not n23192 ; n23193
g20758 nor pi0787 n23052 ; n23194
g20759 and pi1157 n23105_not ; n23195
g20760 nor n23056 n23195 ; n23196
g20761 and pi0787 n23196_not ; n23197
g20762 nor n23194 n23197 ; n23198
g20763 and pi0644_not n23198 ; n23199
g20764 and pi0644 n23192 ; n23200
g20765 and pi0715 n23199_not ; n23201
g20766 and n23200_not n23201 ; n23202
g20767 nor n17804 n23101 ; n23203
g20768 and n17804 n23036 ; n23204
g20769 nor n23203 n23204 ; n23205
g20770 and pi0644 n23205_not ; n23206
g20771 and pi0644_not n23036 ; n23207
g20772 nor pi0715 n23207 ; n23208
g20773 and n23206_not n23208 ; n23209
g20774 and pi1160 n23209_not ; n23210
g20775 and n23202_not n23210 ; n23211
g20776 nor pi0644 n23205 ; n23212
g20777 and pi0644 n23036 ; n23213
g20778 and pi0715 n23213_not ; n23214
g20779 and n23212_not n23214 ; n23215
g20780 and pi0644 n23198 ; n23216
g20781 and pi0644_not n23192 ; n23217
g20782 nor pi0715 n23216 ; n23218
g20783 and n23217_not n23218 ; n23219
g20784 nor pi1160 n23215 ; n23220
g20785 and n23219_not n23220 ; n23221
g20786 nor n23211 n23221 ; n23222
g20787 and pi0790 n23222_not ; n23223
g20788 and pi0832 n23193_not ; n23224
g20789 and n23223_not n23224 ; n23225
g20790 nor n23035 n23225 ; po0330
g20791 and pi0174 n17059_not ; n23227
g20792 and n16635 n23227_not ; n23228
g20793 and n17075 n23227_not ; n23229
g20794 and pi0696 n2571 ; n23230
g20795 nor n23227 n23230 ; n23231
g20796 nor pi0174 n16641 ; n23232
g20797 and n19899 n23232_not ; n23233
g20798 and pi0174_not n18076 ; n23234
g20799 and pi0174 n18072_not ; n23235
g20800 nor pi0038 n23234 ; n23236
g20801 and n23235_not n23236 ; n23237
g20802 and n23230 n23233_not ; n23238
g20803 and n23237_not n23238 ; n23239
g20804 nor n23231 n23239 ; n23240
g20805 and pi0778_not n23240 ; n23241
g20806 nor pi0625 n23227 ; n23242
g20807 and pi0625 n23240_not ; n23243
g20808 and pi1153 n23242_not ; n23244
g20809 and n23243_not n23244 ; n23245
g20810 nor pi0625 n23240 ; n23246
g20811 and pi0625 n23227_not ; n23247
g20812 nor pi1153 n23247 ; n23248
g20813 and n23246_not n23248 ; n23249
g20814 nor n23245 n23249 ; n23250
g20815 and pi0778 n23250_not ; n23251
g20816 nor n23241 n23251 ; n23252
g20817 and n17075_not n23252 ; n23253
g20818 nor n23229 n23253 ; n23254
g20819 and n16639_not n23254 ; n23255
g20820 and n16639 n23227 ; n23256
g20821 nor n23255 n23256 ; n23257
g20822 and n16635_not n23257 ; n23258
g20823 nor n23228 n23258 ; n23259
g20824 and n16631_not n23259 ; n23260
g20825 and n16631 n23227 ; n23261
g20826 nor n23260 n23261 ; n23262
g20827 nor pi0792 n23262 ; n23263
g20828 nor pi0628 n23227 ; n23264
g20829 and pi0628 n23262 ; n23265
g20830 and pi1156 n23264_not ; n23266
g20831 and n23265_not n23266 ; n23267
g20832 and pi0628 n23227_not ; n23268
g20833 and pi0628_not n23262 ; n23269
g20834 nor pi1156 n23268 ; n23270
g20835 and n23269_not n23270 ; n23271
g20836 nor n23267 n23271 ; n23272
g20837 and pi0792 n23272_not ; n23273
g20838 nor n23263 n23273 ; n23274
g20839 nor pi0787 n23274 ; n23275
g20840 nor pi0647 n23227 ; n23276
g20841 and pi0647 n23274 ; n23277
g20842 and pi1157 n23276_not ; n23278
g20843 and n23277_not n23278 ; n23279
g20844 and pi0647 n23227_not ; n23280
g20845 and pi0647_not n23274 ; n23281
g20846 nor pi1157 n23280 ; n23282
g20847 and n23281_not n23282 ; n23283
g20848 nor n23279 n23283 ; n23284
g20849 and pi0787 n23284_not ; n23285
g20850 nor n23275 n23285 ; n23286
g20851 and pi0644_not n23286 ; n23287
g20852 nor pi0619 n23227 ; n23288
g20853 and n17117 n23227_not ; n23289
g20854 and pi0174 n2571_not ; n23290
g20855 and pi0759 n17219 ; n23291
g20856 nor n21470 n23291 ; n23292
g20857 and pi0039 n23292_not ; n23293
g20858 and pi0759_not n16958 ; n23294
g20859 and pi0759 n17139 ; n23295
g20860 nor pi0039 n23294 ; n23296
g20861 and n23295_not n23296 ; n23297
g20862 nor n23293 n23297 ; n23298
g20863 and pi0174 n23298_not ; n23299
g20864 and pi0174_not pi0759 ; n23300
g20865 and n17275 n23300 ; n23301
g20866 nor n23299 n23301 ; n23302
g20867 nor pi0038 n23302 ; n23303
g20868 and pi0759 n17168 ; n23304
g20869 and n16641 n23304_not ; n23305
g20870 and pi0038 n23232_not ; n23306
g20871 and n23305_not n23306 ; n23307
g20872 nor n23303 n23307 ; n23308
g20873 and n2571 n23308_not ; n23309
g20874 nor n23290 n23309 ; n23310
g20875 and n17117_not n23310 ; n23311
g20876 nor n23289 n23311 ; n23312
g20877 and pi0785_not n23312 ; n23313
g20878 nor pi0609 n23227 ; n23314
g20879 and pi0609 n23312_not ; n23315
g20880 and pi1155 n23314_not ; n23316
g20881 and n23315_not n23316 ; n23317
g20882 nor pi0609 n23312 ; n23318
g20883 and pi0609 n23227_not ; n23319
g20884 nor pi1155 n23319 ; n23320
g20885 and n23318_not n23320 ; n23321
g20886 nor n23317 n23321 ; n23322
g20887 and pi0785 n23322_not ; n23323
g20888 nor n23313 n23323 ; n23324
g20889 nor pi0781 n23324 ; n23325
g20890 nor pi0618 n23227 ; n23326
g20891 and pi0618 n23324 ; n23327
g20892 and pi1154 n23326_not ; n23328
g20893 and n23327_not n23328 ; n23329
g20894 and pi0618 n23227_not ; n23330
g20895 and pi0618_not n23324 ; n23331
g20896 nor pi1154 n23330 ; n23332
g20897 and n23331_not n23332 ; n23333
g20898 nor n23329 n23333 ; n23334
g20899 and pi0781 n23334_not ; n23335
g20900 nor n23325 n23335 ; n23336
g20901 and pi0619 n23336 ; n23337
g20902 and pi1159 n23288_not ; n23338
g20903 and n23337_not n23338 ; n23339
g20904 and pi0696_not n23308 ; n23340
g20905 nor pi0174 n17605 ; n23341
g20906 and pi0174 n17546 ; n23342
g20907 and pi0759 n23342_not ; n23343
g20908 and n23341_not n23343 ; n23344
g20909 and pi0174 n17404_not ; n23345
g20910 nor pi0174 n17485 ; n23346
g20911 nor pi0759 n23346 ; n23347
g20912 and n23345_not n23347 ; n23348
g20913 and pi0039 n23344_not ; n23349
g20914 and n23348_not n23349 ; n23350
g20915 and pi0174_not n17631 ; n23351
g20916 and pi0174 n17629 ; n23352
g20917 and pi0759 n23351_not ; n23353
g20918 and n23352_not n23353 ; n23354
g20919 nor pi0174 n17625 ; n23355
g20920 and pi0174 n17612_not ; n23356
g20921 nor pi0759 n23355 ; n23357
g20922 and n23356_not n23357 ; n23358
g20923 nor pi0039 n23354 ; n23359
g20924 and n23358_not n23359 ; n23360
g20925 nor pi0038 n23360 ; n23361
g20926 and n23350_not n23361 ; n23362
g20927 and pi0696 n19470_not ; n23363
g20928 and n23307_not n23363 ; n23364
g20929 and n23362_not n23364 ; n23365
g20930 and n2571 n23365_not ; n23366
g20931 and n23340_not n23366 ; n23367
g20932 nor n23290 n23367 ; n23368
g20933 and pi0625_not n23368 ; n23369
g20934 and pi0625 n23310 ; n23370
g20935 nor pi1153 n23370 ; n23371
g20936 and n23369_not n23371 ; n23372
g20937 nor pi0608 n23245 ; n23373
g20938 and n23372_not n23373 ; n23374
g20939 and pi0625_not n23310 ; n23375
g20940 and pi0625 n23368 ; n23376
g20941 and pi1153 n23375_not ; n23377
g20942 and n23376_not n23377 ; n23378
g20943 and pi0608 n23249_not ; n23379
g20944 and n23378_not n23379 ; n23380
g20945 nor n23374 n23380 ; n23381
g20946 and pi0778 n23381_not ; n23382
g20947 and pi0778_not n23368 ; n23383
g20948 nor n23382 n23383 ; n23384
g20949 nor pi0609 n23384 ; n23385
g20950 and pi0609 n23252 ; n23386
g20951 nor pi1155 n23386 ; n23387
g20952 and n23385_not n23387 ; n23388
g20953 nor pi0660 n23317 ; n23389
g20954 and n23388_not n23389 ; n23390
g20955 and pi0609_not n23252 ; n23391
g20956 and pi0609 n23384_not ; n23392
g20957 and pi1155 n23391_not ; n23393
g20958 and n23392_not n23393 ; n23394
g20959 and pi0660 n23321_not ; n23395
g20960 and n23394_not n23395 ; n23396
g20961 nor n23390 n23396 ; n23397
g20962 and pi0785 n23397_not ; n23398
g20963 nor pi0785 n23384 ; n23399
g20964 nor n23398 n23399 ; n23400
g20965 nor pi0618 n23400 ; n23401
g20966 and pi0618 n23254_not ; n23402
g20967 nor pi1154 n23402 ; n23403
g20968 and n23401_not n23403 ; n23404
g20969 nor pi0627 n23329 ; n23405
g20970 and n23404_not n23405 ; n23406
g20971 and pi0618 n23400_not ; n23407
g20972 nor pi0618 n23254 ; n23408
g20973 and pi1154 n23408_not ; n23409
g20974 and n23407_not n23409 ; n23410
g20975 and pi0627 n23333_not ; n23411
g20976 and n23410_not n23411 ; n23412
g20977 nor n23406 n23412 ; n23413
g20978 and pi0781 n23413_not ; n23414
g20979 nor pi0781 n23400 ; n23415
g20980 nor n23414 n23415 ; n23416
g20981 nor pi0619 n23416 ; n23417
g20982 and pi0619 n23257 ; n23418
g20983 nor pi1159 n23418 ; n23419
g20984 and n23417_not n23419 ; n23420
g20985 nor pi0648 n23339 ; n23421
g20986 and n23420_not n23421 ; n23422
g20987 and pi0619 n23227_not ; n23423
g20988 and pi0619_not n23336 ; n23424
g20989 nor pi1159 n23423 ; n23425
g20990 and n23424_not n23425 ; n23426
g20991 and pi0619_not n23257 ; n23427
g20992 and pi0619 n23416_not ; n23428
g20993 and pi1159 n23427_not ; n23429
g20994 and n23428_not n23429 ; n23430
g20995 and pi0648 n23426_not ; n23431
g20996 and n23430_not n23431 ; n23432
g20997 nor n23422 n23432 ; n23433
g20998 and pi0789 n23433_not ; n23434
g20999 nor pi0789 n23416 ; n23435
g21000 nor n23434 n23435 ; n23436
g21001 and pi0788_not n23436 ; n23437
g21002 and pi0626_not n23436 ; n23438
g21003 and pi0626 n23259 ; n23439
g21004 nor pi0641 n23439 ; n23440
g21005 and n23438_not n23440 ; n23441
g21006 nor pi0789 n23336 ; n23442
g21007 nor n23339 n23426 ; n23443
g21008 and pi0789 n23443_not ; n23444
g21009 nor n23442 n23444 ; n23445
g21010 nor pi0626 n23445 ; n23446
g21011 and pi0626 n23227 ; n23447
g21012 and pi0641 n23447_not ; n23448
g21013 and n23446_not n23448 ; n23449
g21014 nor pi1158 n23449 ; n23450
g21015 and n23441_not n23450 ; n23451
g21016 and pi0626 n23436 ; n23452
g21017 and pi0626_not n23259 ; n23453
g21018 and pi0641 n23453_not ; n23454
g21019 and n23452_not n23454 ; n23455
g21020 and pi0626 n23445_not ; n23456
g21021 and pi0626_not n23227 ; n23457
g21022 nor pi0641 n23457 ; n23458
g21023 and n23456_not n23458 ; n23459
g21024 and pi1158 n23459_not ; n23460
g21025 and n23455_not n23460 ; n23461
g21026 nor n23451 n23461 ; n23462
g21027 and pi0788 n23462_not ; n23463
g21028 nor n23437 n23463 ; n23464
g21029 and pi0628_not n23464 ; n23465
g21030 nor n17969 n23445 ; n23466
g21031 and n17969 n23227 ; n23467
g21032 nor n23466 n23467 ; n23468
g21033 and pi0628 n23468 ; n23469
g21034 nor pi1156 n23469 ; n23470
g21035 and n23465_not n23470 ; n23471
g21036 nor pi0629 n23267 ; n23472
g21037 and n23471_not n23472 ; n23473
g21038 and pi0628 n23464 ; n23474
g21039 and pi0628_not n23468 ; n23475
g21040 and pi1156 n23475_not ; n23476
g21041 and n23474_not n23476 ; n23477
g21042 and pi0629 n23271_not ; n23478
g21043 and n23477_not n23478 ; n23479
g21044 nor n23473 n23479 ; n23480
g21045 and pi0792 n23480_not ; n23481
g21046 and pi0792_not n23464 ; n23482
g21047 nor n23481 n23482 ; n23483
g21048 nor pi0647 n23483 ; n23484
g21049 nor n17779 n23468 ; n23485
g21050 and n17779 n23227 ; n23486
g21051 nor n23485 n23486 ; n23487
g21052 and pi0647 n23487 ; n23488
g21053 nor pi1157 n23488 ; n23489
g21054 and n23484_not n23489 ; n23490
g21055 nor pi0630 n23279 ; n23491
g21056 and n23490_not n23491 ; n23492
g21057 and pi0647 n23483_not ; n23493
g21058 and pi0647_not n23487 ; n23494
g21059 and pi1157 n23494_not ; n23495
g21060 and n23493_not n23495 ; n23496
g21061 and pi0630 n23283_not ; n23497
g21062 and n23496_not n23497 ; n23498
g21063 nor n23492 n23498 ; n23499
g21064 and pi0787 n23499_not ; n23500
g21065 nor pi0787 n23483 ; n23501
g21066 nor n23500 n23501 ; n23502
g21067 and pi0644 n23502_not ; n23503
g21068 and pi0715 n23287_not ; n23504
g21069 and n23503_not n23504 ; n23505
g21070 and n17804 n23227_not ; n23506
g21071 and n17804_not n23487 ; n23507
g21072 nor n23506 n23507 ; n23508
g21073 and pi0644 n23508_not ; n23509
g21074 nor pi0644 n23227 ; n23510
g21075 nor pi0715 n23510 ; n23511
g21076 and n23509_not n23511 ; n23512
g21077 and pi1160 n23512_not ; n23513
g21078 and n23505_not n23513 ; n23514
g21079 nor pi0644 n23502 ; n23515
g21080 and pi0644 n23286 ; n23516
g21081 nor pi0715 n23516 ; n23517
g21082 and n23515_not n23517 ; n23518
g21083 nor pi0644 n23508 ; n23519
g21084 and pi0644 n23227_not ; n23520
g21085 and pi0715 n23520_not ; n23521
g21086 and n23519_not n23521 ; n23522
g21087 nor pi1160 n23522 ; n23523
g21088 and n23518_not n23523 ; n23524
g21089 and pi0790 n23514_not ; n23525
g21090 and n23524_not n23525 ; n23526
g21091 and pi0790_not n23502 ; n23527
g21092 and n6305 n23527_not ; n23528
g21093 and n23526_not n23528 ; n23529
g21094 nor pi0174 n6305 ; n23530
g21095 nor pi0057 n23530 ; n23531
g21096 and n23529_not n23531 ; n23532
g21097 and pi0057 pi0174 ; n23533
g21098 nor pi0832 n23533 ; n23534
g21099 and n23532_not n23534 ; n23535
g21100 and pi0174 n2926_not ; n23536
g21101 and pi0759 n17244 ; n23537
g21102 and n17291 n23537 ; n23538
g21103 and pi1155 n23536_not ; n23539
g21104 and n23538_not n23539 ; n23540
g21105 and pi0696 n16645 ; n23541
g21106 nor n23536 n23541 ; n23542
g21107 and pi0778_not n23542 ; n23543
g21108 and pi0625 n23541 ; n23544
g21109 nor n23542 n23544 ; n23545
g21110 nor pi1153 n23545 ; n23546
g21111 and pi1153 n23536_not ; n23547
g21112 and n23544_not n23547 ; n23548
g21113 nor n23546 n23548 ; n23549
g21114 and pi0778 n23549_not ; n23550
g21115 nor n23543 n23550 ; n23551
g21116 and pi0609 n23551 ; n23552
g21117 nor n23536 n23537 ; n23553
g21118 and pi0696 n17469 ; n23554
g21119 and n23553 n23554_not ; n23555
g21120 and pi0625 n23554 ; n23556
g21121 nor n23555 n23556 ; n23557
g21122 nor pi1153 n23557 ; n23558
g21123 nor pi0608 n23548 ; n23559
g21124 and n23558_not n23559 ; n23560
g21125 and pi1153 n23553 ; n23561
g21126 and n23556_not n23561 ; n23562
g21127 and pi0608 n23546_not ; n23563
g21128 and n23562_not n23563 ; n23564
g21129 nor n23560 n23564 ; n23565
g21130 and pi0778 n23565_not ; n23566
g21131 nor pi0778 n23555 ; n23567
g21132 nor n23566 n23567 ; n23568
g21133 nor pi0609 n23568 ; n23569
g21134 nor pi1155 n23552 ; n23570
g21135 and n23569_not n23570 ; n23571
g21136 nor pi0660 n23540 ; n23572
g21137 and n23571_not n23572 ; n23573
g21138 and n17296 n23537 ; n23574
g21139 nor pi1155 n23536 ; n23575
g21140 and n23574_not n23575 ; n23576
g21141 and pi0609_not n23551 ; n23577
g21142 and pi0609 n23568_not ; n23578
g21143 and pi1155 n23577_not ; n23579
g21144 and n23578_not n23579 ; n23580
g21145 and pi0660 n23576_not ; n23581
g21146 and n23580_not n23581 ; n23582
g21147 nor n23573 n23582 ; n23583
g21148 and pi0785 n23583_not ; n23584
g21149 nor pi0785 n23568 ; n23585
g21150 nor n23584 n23585 ; n23586
g21151 nor pi0781 n23586 ; n23587
g21152 and n20225_not n23537 ; n23588
g21153 and n20270 n23588 ; n23589
g21154 and pi1154 n23536_not ; n23590
g21155 and n23589_not n23590 ; n23591
g21156 and n17075_not n23551 ; n23592
g21157 nor n23536 n23592 ; n23593
g21158 and pi0618 n23593_not ; n23594
g21159 nor pi0618 n23586 ; n23595
g21160 nor pi1154 n23594 ; n23596
g21161 and n23595_not n23596 ; n23597
g21162 nor pi0627 n23591 ; n23598
g21163 and n23597_not n23598 ; n23599
g21164 and n20319 n23588 ; n23600
g21165 nor pi1154 n23536 ; n23601
g21166 and n23600_not n23601 ; n23602
g21167 nor pi0618 n23593 ; n23603
g21168 and pi0618 n23586_not ; n23604
g21169 and pi1154 n23603_not ; n23605
g21170 and n23604_not n23605 ; n23606
g21171 and pi0627 n23602_not ; n23607
g21172 and n23606_not n23607 ; n23608
g21173 nor n23599 n23608 ; n23609
g21174 and pi0781 n23609_not ; n23610
g21175 and pi0648 n20228 ; n23611
g21176 and pi0648_not n20229 ; n23612
g21177 nor n23611 n23612 ; n23613
g21178 and n16634 n23613 ; n23614
g21179 and pi0789 n23614_not ; n23615
g21180 nor n23587 n23615 ; n23616
g21181 and n23610_not n23616 ; n23617
g21182 and n20235_not n23588 ; n23618
g21183 and n20345 n23618 ; n23619
g21184 and n16633 n23619_not ; n23620
g21185 and n19150 n23551 ; n23621
g21186 nor n23613 n23621 ; n23622
g21187 and n20335 n23618 ; n23623
g21188 and n16632 n23623_not ; n23624
g21189 nor n23620 n23624 ; n23625
g21190 and n23622_not n23625 ; n23626
g21191 and pi0789 n23536_not ; n23627
g21192 and n23626_not n23627 ; n23628
g21193 and n17970 n23628_not ; n23629
g21194 and n23617_not n23629 ; n23630
g21195 and n20237 n23588 ; n23631
g21196 and pi0626_not n23631 ; n23632
g21197 nor n23536 n23632 ; n23633
g21198 nor pi1158 n23633 ; n23634
g21199 and n16635_not n23621 ; n23635
g21200 nor n23536 n23635 ; n23636
g21201 and n17865 n23636_not ; n23637
g21202 and pi0641 n23634_not ; n23638
g21203 and n23637_not n23638 ; n23639
g21204 and n17866 n23636_not ; n23640
g21205 and pi0626 n23631 ; n23641
g21206 nor n23536 n23641 ; n23642
g21207 and pi1158 n23642_not ; n23643
g21208 nor pi0641 n23643 ; n23644
g21209 and n23640_not n23644 ; n23645
g21210 and pi0788 n23639_not ; n23646
g21211 and n23645_not n23646 ; n23647
g21212 nor n20364 n23647 ; n23648
g21213 and n23630_not n23648 ; n23649
g21214 and n17969_not n23631 ; n23650
g21215 and pi0629_not n23650 ; n23651
g21216 and pi0628 n23651_not ; n23652
g21217 and n19151 n23551 ; n23653
g21218 and pi0629 n23653_not ; n23654
g21219 nor n23652 n23654 ; n23655
g21220 nor pi1156 n23655 ; n23656
g21221 nor pi0628 n23650 ; n23657
g21222 and pi0629 n23657_not ; n23658
g21223 and pi0628 n23653 ; n23659
g21224 and pi1156 n23658_not ; n23660
g21225 and n23659_not n23660 ; n23661
g21226 nor n23656 n23661 ; n23662
g21227 and pi0792 n23536_not ; n23663
g21228 and n23662_not n23663 ; n23664
g21229 nor n23649 n23664 ; n23665
g21230 nor n20206 n23665 ; n23666
g21231 and n17779_not n23650 ; n23667
g21232 and pi0630_not n23667 ; n23668
g21233 and pi0647 n23668_not ; n23669
g21234 and n19142_not n23653 ; n23670
g21235 and pi0630 n23670_not ; n23671
g21236 nor n23669 n23671 ; n23672
g21237 nor pi1157 n23672 ; n23673
g21238 and pi0630 n23667 ; n23674
g21239 nor pi0630 n23670 ; n23675
g21240 and pi0647 n23675_not ; n23676
g21241 and pi1157 n23674_not ; n23677
g21242 and n23676_not n23677 ; n23678
g21243 nor n23673 n23678 ; n23679
g21244 and pi0787 n23536_not ; n23680
g21245 and n23679_not n23680 ; n23681
g21246 nor n23666 n23681 ; n23682
g21247 and pi0790_not n23682 ; n23683
g21248 nor n17779 n17804 ; n23684
g21249 and n23650 n23684 ; n23685
g21250 and pi0644 n23685 ; n23686
g21251 nor pi0715 n23536 ; n23687
g21252 and n23686_not n23687 ; n23688
g21253 and n19342_not n23670 ; n23689
g21254 nor n23536 n23689 ; n23690
g21255 nor pi0644 n23690 ; n23691
g21256 and pi0644 n23682 ; n23692
g21257 and pi0715 n23691_not ; n23693
g21258 and n23692_not n23693 ; n23694
g21259 and pi1160 n23688_not ; n23695
g21260 and n23694_not n23695 ; n23696
g21261 and pi0644_not n23685 ; n23697
g21262 and pi0715 n23536_not ; n23698
g21263 and n23697_not n23698 ; n23699
g21264 and pi0644_not n23682 ; n23700
g21265 and pi0644 n23690_not ; n23701
g21266 nor pi0715 n23701 ; n23702
g21267 and n23700_not n23702 ; n23703
g21268 nor pi1160 n23699 ; n23704
g21269 and n23703_not n23704 ; n23705
g21270 nor n23696 n23705 ; n23706
g21271 and pi0790 n23706_not ; n23707
g21272 and pi0832 n23683_not ; n23708
g21273 and n23707_not n23708 ; n23709
g21274 nor n23535 n23709 ; po0331
g21275 nor pi0175 n2926 ; n23711
g21276 and pi0700 n16645 ; n23712
g21277 nor n23711 n23712 ; n23713
g21278 nor pi0778 n23713 ; n23714
g21279 and pi0625_not n23712 ; n23715
g21280 nor n23713 n23715 ; n23716
g21281 and pi1153 n23716_not ; n23717
g21282 nor pi1153 n23711 ; n23718
g21283 and n23715_not n23718 ; n23719
g21284 and pi0778 n23719_not ; n23720
g21285 and n23717_not n23720 ; n23721
g21286 nor n23714 n23721 ; n23722
g21287 nor n17845 n23722 ; n23723
g21288 and n17847_not n23723 ; n23724
g21289 and n17849_not n23724 ; n23725
g21290 and n17851_not n23725 ; n23726
g21291 and n17857_not n23726 ; n23727
g21292 and pi0647_not n23727 ; n23728
g21293 and pi0647 n23711 ; n23729
g21294 nor pi1157 n23729 ; n23730
g21295 and n23728_not n23730 ; n23731
g21296 and pi0630 n23731 ; n23732
g21297 and pi0766 n17244 ; n23733
g21298 nor n23711 n23733 ; n23734
g21299 nor n17874 n23734 ; n23735
g21300 nor pi0785 n23735 ; n23736
g21301 and n17296 n23733 ; n23737
g21302 and n23735 n23737_not ; n23738
g21303 and pi1155 n23738_not ; n23739
g21304 nor pi1155 n23711 ; n23740
g21305 and n23737_not n23740 ; n23741
g21306 nor n23739 n23741 ; n23742
g21307 and pi0785 n23742_not ; n23743
g21308 nor n23736 n23743 ; n23744
g21309 nor pi0781 n23744 ; n23745
g21310 and n17889_not n23744 ; n23746
g21311 and pi1154 n23746_not ; n23747
g21312 and n17892_not n23744 ; n23748
g21313 nor pi1154 n23748 ; n23749
g21314 nor n23747 n23749 ; n23750
g21315 and pi0781 n23750_not ; n23751
g21316 nor n23745 n23751 ; n23752
g21317 nor pi0789 n23752 ; n23753
g21318 and n23078_not n23752 ; n23754
g21319 and pi1159 n23754_not ; n23755
g21320 and n23081_not n23752 ; n23756
g21321 nor pi1159 n23756 ; n23757
g21322 nor n23755 n23757 ; n23758
g21323 and pi0789 n23758_not ; n23759
g21324 nor n23753 n23759 ; n23760
g21325 and n17969_not n23760 ; n23761
g21326 and n17969 n23711 ; n23762
g21327 nor n23761 n23762 ; n23763
g21328 nor n17779 n23763 ; n23764
g21329 and n17779 n23711 ; n23765
g21330 nor n23764 n23765 ; n23766
g21331 and n20559_not n23766 ; n23767
g21332 and pi0647 n23727_not ; n23768
g21333 nor pi0647 n23711 ; n23769
g21334 nor n23768 n23769 ; n23770
g21335 and n17801 n23770_not ; n23771
g21336 nor n23732 n23771 ; n23772
g21337 and n23767_not n23772 ; n23773
g21338 and pi0787 n23773_not ; n23774
g21339 and n17871 n23725 ; n23775
g21340 nor pi0626 n23760 ; n23776
g21341 and pi0626 n23711_not ; n23777
g21342 and n16629 n23777_not ; n23778
g21343 and n23776_not n23778 ; n23779
g21344 and pi0626 n23760_not ; n23780
g21345 nor pi0626 n23711 ; n23781
g21346 and n16628 n23781_not ; n23782
g21347 and n23780_not n23782 ; n23783
g21348 nor n23775 n23779 ; n23784
g21349 and n23783_not n23784 ; n23785
g21350 and pi0788 n23785_not ; n23786
g21351 and pi0618 n23723 ; n23787
g21352 nor n17168 n23713 ; n23788
g21353 and pi0625 n23788 ; n23789
g21354 and n23734 n23788_not ; n23790
g21355 nor n23789 n23790 ; n23791
g21356 and n23718 n23791_not ; n23792
g21357 nor pi0608 n23717 ; n23793
g21358 and n23792_not n23793 ; n23794
g21359 and pi1153 n23734 ; n23795
g21360 and n23789_not n23795 ; n23796
g21361 and pi0608 n23719_not ; n23797
g21362 and n23796_not n23797 ; n23798
g21363 nor n23794 n23798 ; n23799
g21364 and pi0778 n23799_not ; n23800
g21365 nor pi0778 n23790 ; n23801
g21366 nor n23800 n23801 ; n23802
g21367 nor pi0609 n23802 ; n23803
g21368 and pi0609 n23722_not ; n23804
g21369 nor pi1155 n23804 ; n23805
g21370 and n23803_not n23805 ; n23806
g21371 nor pi0660 n23739 ; n23807
g21372 and n23806_not n23807 ; n23808
g21373 and pi0609 n23802_not ; n23809
g21374 nor pi0609 n23722 ; n23810
g21375 and pi1155 n23810_not ; n23811
g21376 and n23809_not n23811 ; n23812
g21377 and pi0660 n23741_not ; n23813
g21378 and n23812_not n23813 ; n23814
g21379 nor n23808 n23814 ; n23815
g21380 and pi0785 n23815_not ; n23816
g21381 nor pi0785 n23802 ; n23817
g21382 nor n23816 n23817 ; n23818
g21383 nor pi0618 n23818 ; n23819
g21384 nor pi1154 n23787 ; n23820
g21385 and n23819_not n23820 ; n23821
g21386 nor pi0627 n23747 ; n23822
g21387 and n23821_not n23822 ; n23823
g21388 and pi0618_not n23723 ; n23824
g21389 and pi0618 n23818_not ; n23825
g21390 and pi1154 n23824_not ; n23826
g21391 and n23825_not n23826 ; n23827
g21392 and pi0627 n23749_not ; n23828
g21393 and n23827_not n23828 ; n23829
g21394 nor n23823 n23829 ; n23830
g21395 and pi0781 n23830_not ; n23831
g21396 nor pi0781 n23818 ; n23832
g21397 nor n23831 n23832 ; n23833
g21398 and pi0789_not n23833 ; n23834
g21399 nor pi0619 n23833 ; n23835
g21400 and pi0619 n23724 ; n23836
g21401 nor pi1159 n23836 ; n23837
g21402 and n23835_not n23837 ; n23838
g21403 nor pi0648 n23755 ; n23839
g21404 and n23838_not n23839 ; n23840
g21405 and pi0619 n23833_not ; n23841
g21406 and pi0619_not n23724 ; n23842
g21407 and pi1159 n23842_not ; n23843
g21408 and n23841_not n23843 ; n23844
g21409 and pi0648 n23757_not ; n23845
g21410 and n23844_not n23845 ; n23846
g21411 and pi0789 n23840_not ; n23847
g21412 and n23846_not n23847 ; n23848
g21413 and n17970 n23834_not ; n23849
g21414 and n23848_not n23849 ; n23850
g21415 nor n23786 n23850 ; n23851
g21416 nor n20364 n23851 ; n23852
g21417 and n17854 n23763_not ; n23853
g21418 and n20851 n23726 ; n23854
g21419 nor n23853 n23854 ; n23855
g21420 nor pi0629 n23855 ; n23856
g21421 and n20855 n23726 ; n23857
g21422 and n17853 n23763_not ; n23858
g21423 nor n23857 n23858 ; n23859
g21424 and pi0629 n23859_not ; n23860
g21425 nor n23856 n23860 ; n23861
g21426 and pi0792 n23861_not ; n23862
g21427 nor n20206 n23862 ; n23863
g21428 and n23852_not n23863 ; n23864
g21429 nor n23774 n23864 ; n23865
g21430 and pi0790_not n23865 ; n23866
g21431 nor pi0787 n23727 ; n23867
g21432 and pi1157 n23770_not ; n23868
g21433 nor n23731 n23868 ; n23869
g21434 and pi0787 n23869_not ; n23870
g21435 nor n23867 n23870 ; n23871
g21436 and pi0644_not n23871 ; n23872
g21437 and pi0644 n23865 ; n23873
g21438 and pi0715 n23872_not ; n23874
g21439 and n23873_not n23874 ; n23875
g21440 nor n17804 n23766 ; n23876
g21441 and n17804 n23711 ; n23877
g21442 nor n23876 n23877 ; n23878
g21443 and pi0644 n23878_not ; n23879
g21444 and pi0644_not n23711 ; n23880
g21445 nor pi0715 n23880 ; n23881
g21446 and n23879_not n23881 ; n23882
g21447 and pi1160 n23882_not ; n23883
g21448 and n23875_not n23883 ; n23884
g21449 nor pi0644 n23878 ; n23885
g21450 and pi0644 n23711 ; n23886
g21451 and pi0715 n23886_not ; n23887
g21452 and n23885_not n23887 ; n23888
g21453 and pi0644 n23871 ; n23889
g21454 and pi0644_not n23865 ; n23890
g21455 nor pi0715 n23889 ; n23891
g21456 and n23890_not n23891 ; n23892
g21457 nor pi1160 n23888 ; n23893
g21458 and n23892_not n23893 ; n23894
g21459 nor n23884 n23894 ; n23895
g21460 and pi0790 n23895_not ; n23896
g21461 and pi0832 n23866_not ; n23897
g21462 and n23896_not n23897 ; n23898
g21463 and pi0175_not po1038 ; n23899
g21464 nor pi0175 n17059 ; n23900
g21465 and n16635 n23900_not ; n23901
g21466 and pi0175 n2571_not ; n23902
g21467 nor pi0175 n16641 ; n23903
g21468 and n16647 n23903_not ; n23904
g21469 and pi0175_not n18072 ; n23905
g21470 and pi0175 n18076_not ; n23906
g21471 nor pi0038 n23906 ; n23907
g21472 and n23905_not n23907 ; n23908
g21473 and pi0700 n23904_not ; n23909
g21474 and n23908_not n23909 ; n23910
g21475 nor pi0175 pi0700 ; n23911
g21476 and n17052_not n23911 ; n23912
g21477 and n2571 n23912_not ; n23913
g21478 and n23910_not n23913 ; n23914
g21479 nor n23902 n23914 ; n23915
g21480 nor pi0778 n23915 ; n23916
g21481 and pi0625_not n23900 ; n23917
g21482 and pi0625 n23915 ; n23918
g21483 and pi1153 n23917_not ; n23919
g21484 and n23918_not n23919 ; n23920
g21485 and pi0625_not n23915 ; n23921
g21486 and pi0625 n23900 ; n23922
g21487 nor pi1153 n23922 ; n23923
g21488 and n23921_not n23923 ; n23924
g21489 nor n23920 n23924 ; n23925
g21490 and pi0778 n23925_not ; n23926
g21491 nor n23916 n23926 ; n23927
g21492 nor n17075 n23927 ; n23928
g21493 and n17075 n23900_not ; n23929
g21494 nor n23928 n23929 ; n23930
g21495 and n16639_not n23930 ; n23931
g21496 and n16639 n23900 ; n23932
g21497 nor n23931 n23932 ; n23933
g21498 and n16635_not n23933 ; n23934
g21499 nor n23901 n23934 ; n23935
g21500 and n16631_not n23935 ; n23936
g21501 and n16631 n23900 ; n23937
g21502 nor n23936 n23937 ; n23938
g21503 nor pi0628 n23938 ; n23939
g21504 and pi0628 n23900 ; n23940
g21505 nor n23939 n23940 ; n23941
g21506 nor pi1156 n23941 ; n23942
g21507 and pi0628 n23938_not ; n23943
g21508 and pi0628_not n23900 ; n23944
g21509 nor n23943 n23944 ; n23945
g21510 and pi1156 n23945_not ; n23946
g21511 nor n23942 n23946 ; n23947
g21512 and pi0792 n23947_not ; n23948
g21513 nor pi0792 n23938 ; n23949
g21514 nor n23948 n23949 ; n23950
g21515 nor pi0647 n23950 ; n23951
g21516 and pi0647 n23900 ; n23952
g21517 nor n23951 n23952 ; n23953
g21518 nor pi1157 n23953 ; n23954
g21519 and pi0647 n23950_not ; n23955
g21520 and pi0647_not n23900 ; n23956
g21521 nor n23955 n23956 ; n23957
g21522 and pi1157 n23957_not ; n23958
g21523 nor n23954 n23958 ; n23959
g21524 and pi0787 n23959_not ; n23960
g21525 nor pi0787 n23950 ; n23961
g21526 nor n23960 n23961 ; n23962
g21527 nor pi0644 n23962 ; n23963
g21528 and pi0715 n23963_not ; n23964
g21529 and pi0766_not n17046 ; n23965
g21530 and pi0175 n17273 ; n23966
g21531 nor n23965 n23966 ; n23967
g21532 and pi0039 n23967_not ; n23968
g21533 and pi0766 n17234_not ; n23969
g21534 and pi0175 n23969_not ; n23970
g21535 and pi0175_not pi0766 ; n23971
g21536 and n17221 n23971 ; n23972
g21537 nor n21499 n23970 ; n23973
g21538 and n23972_not n23973 ; n23974
g21539 and n23968_not n23974 ; n23975
g21540 nor pi0038 n23975 ; n23976
g21541 and pi0766 n17280 ; n23977
g21542 and pi0038 n23903_not ; n23978
g21543 and n23977_not n23978 ; n23979
g21544 nor n23976 n23979 ; n23980
g21545 and n2571 n23980_not ; n23981
g21546 nor n23902 n23981 ; n23982
g21547 nor n17117 n23982 ; n23983
g21548 and n17117 n23900_not ; n23984
g21549 nor n23983 n23984 ; n23985
g21550 nor pi0785 n23985 ; n23986
g21551 nor n17291 n23900 ; n23987
g21552 and pi0609 n23983 ; n23988
g21553 nor n23987 n23988 ; n23989
g21554 and pi1155 n23989_not ; n23990
g21555 nor n17296 n23900 ; n23991
g21556 and pi0609_not n23983 ; n23992
g21557 nor n23991 n23992 ; n23993
g21558 nor pi1155 n23993 ; n23994
g21559 nor n23990 n23994 ; n23995
g21560 and pi0785 n23995_not ; n23996
g21561 nor n23986 n23996 ; n23997
g21562 nor pi0781 n23997 ; n23998
g21563 and pi0618_not n23900 ; n23999
g21564 and pi0618 n23997 ; n24000
g21565 and pi1154 n23999_not ; n24001
g21566 and n24000_not n24001 ; n24002
g21567 and pi0618_not n23997 ; n24003
g21568 and pi0618 n23900 ; n24004
g21569 nor pi1154 n24004 ; n24005
g21570 and n24003_not n24005 ; n24006
g21571 nor n24002 n24006 ; n24007
g21572 and pi0781 n24007_not ; n24008
g21573 nor n23998 n24008 ; n24009
g21574 nor pi0789 n24009 ; n24010
g21575 and pi0619_not n23900 ; n24011
g21576 and pi0619 n24009 ; n24012
g21577 and pi1159 n24011_not ; n24013
g21578 and n24012_not n24013 ; n24014
g21579 and pi0619_not n24009 ; n24015
g21580 and pi0619 n23900 ; n24016
g21581 nor pi1159 n24016 ; n24017
g21582 and n24015_not n24017 ; n24018
g21583 nor n24014 n24018 ; n24019
g21584 and pi0789 n24019_not ; n24020
g21585 nor n24010 n24020 ; n24021
g21586 and n17969_not n24021 ; n24022
g21587 and n17969 n23900 ; n24023
g21588 nor n24022 n24023 ; n24024
g21589 nor n17779 n24024 ; n24025
g21590 and n17779 n23900 ; n24026
g21591 nor n24025 n24026 ; n24027
g21592 nor n17804 n24027 ; n24028
g21593 and n17804 n23900 ; n24029
g21594 nor n24028 n24029 ; n24030
g21595 and pi0644 n24030_not ; n24031
g21596 and pi0644_not n23900 ; n24032
g21597 nor pi0715 n24032 ; n24033
g21598 and n24031_not n24033 ; n24034
g21599 and pi1160 n24034_not ; n24035
g21600 and n23964_not n24035 ; n24036
g21601 and pi0644 n23962_not ; n24037
g21602 nor pi0715 n24037 ; n24038
g21603 nor pi0644 n24030 ; n24039
g21604 and pi0644 n23900 ; n24040
g21605 and pi0715 n24040_not ; n24041
g21606 and n24039_not n24041 ; n24042
g21607 nor pi1160 n24042 ; n24043
g21608 and n24038_not n24043 ; n24044
g21609 nor n24036 n24044 ; n24045
g21610 and pi0790 n24045_not ; n24046
g21611 and n17777 n23941 ; n24047
g21612 and n20570_not n24024 ; n24048
g21613 and n17776 n23945 ; n24049
g21614 nor n24047 n24049 ; n24050
g21615 and n24048_not n24050 ; n24051
g21616 and pi0792 n24051_not ; n24052
g21617 and pi0609 n23927 ; n24053
g21618 and pi0700_not n23980 ; n24054
g21619 and n16667 n17336_not ; n24055
g21620 and pi0766_not n24055 ; n24056
g21621 nor n17490 n24056 ; n24057
g21622 nor pi0039 n24057 ; n24058
g21623 nor pi0175 n24058 ; n24059
g21624 nor n17469 n23733 ; n24060
g21625 and pi0175 n24060_not ; n24061
g21626 and n6284 n24061 ; n24062
g21627 and pi0038 n24062_not ; n24063
g21628 and n24059_not n24063 ; n24064
g21629 nor pi0175 n17629 ; n24065
g21630 and pi0175 n17631_not ; n24066
g21631 and pi0766 n24066_not ; n24067
g21632 and n24065_not n24067 ; n24068
g21633 and pi0175_not n17612 ; n24069
g21634 and pi0175 n17625 ; n24070
g21635 nor pi0766 n24069 ; n24071
g21636 and n24070_not n24071 ; n24072
g21637 nor pi0039 n24068 ; n24073
g21638 and n24072_not n24073 ; n24074
g21639 and pi0175 n17605 ; n24075
g21640 nor pi0175 n17546 ; n24076
g21641 and pi0766 n24076_not ; n24077
g21642 and n24075_not n24077 ; n24078
g21643 and pi0175_not n17404 ; n24079
g21644 and pi0175 n17485 ; n24080
g21645 nor pi0766 n24080 ; n24081
g21646 and n24079_not n24081 ; n24082
g21647 and pi0039 n24078_not ; n24083
g21648 and n24082_not n24083 ; n24084
g21649 nor pi0038 n24074 ; n24085
g21650 and n24084_not n24085 ; n24086
g21651 and pi0700 n24064_not ; n24087
g21652 and n24086_not n24087 ; n24088
g21653 and n2571 n24088_not ; n24089
g21654 and n24054_not n24089 ; n24090
g21655 nor n23902 n24090 ; n24091
g21656 and pi0625_not n24091 ; n24092
g21657 and pi0625 n23982 ; n24093
g21658 nor pi1153 n24093 ; n24094
g21659 and n24092_not n24094 ; n24095
g21660 nor pi0608 n23920 ; n24096
g21661 and n24095_not n24096 ; n24097
g21662 and pi0625_not n23982 ; n24098
g21663 and pi0625 n24091 ; n24099
g21664 and pi1153 n24098_not ; n24100
g21665 and n24099_not n24100 ; n24101
g21666 and pi0608 n23924_not ; n24102
g21667 and n24101_not n24102 ; n24103
g21668 nor n24097 n24103 ; n24104
g21669 and pi0778 n24104_not ; n24105
g21670 and pi0778_not n24091 ; n24106
g21671 nor n24105 n24106 ; n24107
g21672 nor pi0609 n24107 ; n24108
g21673 nor pi1155 n24053 ; n24109
g21674 and n24108_not n24109 ; n24110
g21675 nor pi0660 n23990 ; n24111
g21676 and n24110_not n24111 ; n24112
g21677 and pi0609_not n23927 ; n24113
g21678 and pi0609 n24107_not ; n24114
g21679 and pi1155 n24113_not ; n24115
g21680 and n24114_not n24115 ; n24116
g21681 and pi0660 n23994_not ; n24117
g21682 and n24116_not n24117 ; n24118
g21683 nor n24112 n24118 ; n24119
g21684 and pi0785 n24119_not ; n24120
g21685 nor pi0785 n24107 ; n24121
g21686 nor n24120 n24121 ; n24122
g21687 nor pi0618 n24122 ; n24123
g21688 and pi0618 n23930 ; n24124
g21689 nor pi1154 n24124 ; n24125
g21690 and n24123_not n24125 ; n24126
g21691 nor pi0627 n24002 ; n24127
g21692 and n24126_not n24127 ; n24128
g21693 and pi0618_not n23930 ; n24129
g21694 and pi0618 n24122_not ; n24130
g21695 and pi1154 n24129_not ; n24131
g21696 and n24130_not n24131 ; n24132
g21697 and pi0627 n24006_not ; n24133
g21698 and n24132_not n24133 ; n24134
g21699 nor n24128 n24134 ; n24135
g21700 and pi0781 n24135_not ; n24136
g21701 nor pi0781 n24122 ; n24137
g21702 nor n24136 n24137 ; n24138
g21703 and pi0789_not n24138 ; n24139
g21704 and pi0619 n23933_not ; n24140
g21705 nor pi0619 n24138 ; n24141
g21706 nor pi1159 n24140 ; n24142
g21707 and n24141_not n24142 ; n24143
g21708 nor pi0648 n24014 ; n24144
g21709 and n24143_not n24144 ; n24145
g21710 nor pi0619 n23933 ; n24146
g21711 and pi0619 n24138_not ; n24147
g21712 and pi1159 n24146_not ; n24148
g21713 and n24147_not n24148 ; n24149
g21714 and pi0648 n24018_not ; n24150
g21715 and n24149_not n24150 ; n24151
g21716 and pi0789 n24145_not ; n24152
g21717 and n24151_not n24152 ; n24153
g21718 and n17970 n24139_not ; n24154
g21719 and n24153_not n24154 ; n24155
g21720 and n17871 n23935 ; n24156
g21721 nor pi0626 n24021 ; n24157
g21722 and pi0626 n23900_not ; n24158
g21723 and n16629 n24158_not ; n24159
g21724 and n24157_not n24159 ; n24160
g21725 and pi0626 n24021_not ; n24161
g21726 nor pi0626 n23900 ; n24162
g21727 and n16628 n24162_not ; n24163
g21728 and n24161_not n24163 ; n24164
g21729 nor n24156 n24160 ; n24165
g21730 and n24164_not n24165 ; n24166
g21731 and pi0788 n24166_not ; n24167
g21732 nor n20364 n24167 ; n24168
g21733 and n24155_not n24168 ; n24169
g21734 nor n24052 n24169 ; n24170
g21735 nor n20206 n24170 ; n24171
g21736 and n17802 n23953 ; n24172
g21737 and n20559_not n24027 ; n24173
g21738 and n17801 n23957 ; n24174
g21739 nor n24172 n24173 ; n24175
g21740 and n24174_not n24175 ; n24176
g21741 and pi0787 n24176_not ; n24177
g21742 and pi0644_not n24043 ; n24178
g21743 and pi0644 n24035 ; n24179
g21744 and pi0790 n24178_not ; n24180
g21745 and n24179_not n24180 ; n24181
g21746 nor n24171 n24177 ; n24182
g21747 and n24181_not n24182 ; n24183
g21748 nor n24046 n24183 ; n24184
g21749 nor po1038 n24184 ; n24185
g21750 nor pi0832 n23899 ; n24186
g21751 and n24185_not n24186 ; n24187
g21752 nor n23898 n24187 ; po0332
g21753 nor pi0176 n2926 ; n24189
g21754 and pi0704_not n16645 ; n24190
g21755 nor n24189 n24190 ; n24191
g21756 and pi0778_not n24191 ; n24192
g21757 and pi0625_not n24190 ; n24193
g21758 nor n24191 n24193 ; n24194
g21759 and pi1153 n24194_not ; n24195
g21760 nor pi1153 n24189 ; n24196
g21761 and n24193_not n24196 ; n24197
g21762 nor n24195 n24197 ; n24198
g21763 and pi0778 n24198_not ; n24199
g21764 nor n24192 n24199 ; n24200
g21765 and n17845_not n24200 ; n24201
g21766 and n17847_not n24201 ; n24202
g21767 and n17849_not n24202 ; n24203
g21768 and n17851_not n24203 ; n24204
g21769 and n17857_not n24204 ; n24205
g21770 and pi0647_not n24205 ; n24206
g21771 and pi0647 n24189 ; n24207
g21772 nor pi1157 n24207 ; n24208
g21773 and n24206_not n24208 ; n24209
g21774 and pi0630 n24209 ; n24210
g21775 and pi0742_not n17244 ; n24211
g21776 nor n24189 n24211 ; n24212
g21777 nor n17874 n24212 ; n24213
g21778 nor pi0785 n24213 ; n24214
g21779 nor n17879 n24212 ; n24215
g21780 and pi1155 n24215_not ; n24216
g21781 and n17882_not n24213 ; n24217
g21782 nor pi1155 n24217 ; n24218
g21783 nor n24216 n24218 ; n24219
g21784 and pi0785 n24219_not ; n24220
g21785 nor n24214 n24220 ; n24221
g21786 nor pi0781 n24221 ; n24222
g21787 and n17889_not n24221 ; n24223
g21788 and pi1154 n24223_not ; n24224
g21789 and n17892_not n24221 ; n24225
g21790 nor pi1154 n24225 ; n24226
g21791 nor n24224 n24226 ; n24227
g21792 and pi0781 n24227_not ; n24228
g21793 nor n24222 n24228 ; n24229
g21794 nor pi0789 n24229 ; n24230
g21795 and pi0619_not n24189 ; n24231
g21796 and pi0619 n24229 ; n24232
g21797 and pi1159 n24231_not ; n24233
g21798 and n24232_not n24233 ; n24234
g21799 and pi0619_not n24229 ; n24235
g21800 and pi0619 n24189 ; n24236
g21801 nor pi1159 n24236 ; n24237
g21802 and n24235_not n24237 ; n24238
g21803 nor n24234 n24238 ; n24239
g21804 and pi0789 n24239_not ; n24240
g21805 nor n24230 n24240 ; n24241
g21806 and n17969_not n24241 ; n24242
g21807 and n17969 n24189 ; n24243
g21808 nor n24242 n24243 ; n24244
g21809 nor n17779 n24244 ; n24245
g21810 and n17779 n24189 ; n24246
g21811 nor n24245 n24246 ; n24247
g21812 and n20559_not n24247 ; n24248
g21813 and pi0647 n24205_not ; n24249
g21814 nor pi0647 n24189 ; n24250
g21815 nor n24249 n24250 ; n24251
g21816 and n17801 n24251_not ; n24252
g21817 nor n24210 n24252 ; n24253
g21818 and n24248_not n24253 ; n24254
g21819 and pi0787 n24254_not ; n24255
g21820 and n17871 n24203 ; n24256
g21821 nor pi0626 n24241 ; n24257
g21822 and pi0626 n24189_not ; n24258
g21823 and n16629 n24258_not ; n24259
g21824 and n24257_not n24259 ; n24260
g21825 and pi0626 n24241_not ; n24261
g21826 nor pi0626 n24189 ; n24262
g21827 and n16628 n24262_not ; n24263
g21828 and n24261_not n24263 ; n24264
g21829 nor n24256 n24260 ; n24265
g21830 and n24264_not n24265 ; n24266
g21831 and pi0788 n24266_not ; n24267
g21832 and pi0618 n24201 ; n24268
g21833 and pi0609 n24200 ; n24269
g21834 nor n17168 n24191 ; n24270
g21835 and pi0625 n24270 ; n24271
g21836 and n24212 n24270_not ; n24272
g21837 nor n24271 n24272 ; n24273
g21838 and n24196 n24273_not ; n24274
g21839 nor pi0608 n24195 ; n24275
g21840 and n24274_not n24275 ; n24276
g21841 and pi1153 n24212 ; n24277
g21842 and n24271_not n24277 ; n24278
g21843 and pi0608 n24197_not ; n24279
g21844 and n24278_not n24279 ; n24280
g21845 nor n24276 n24280 ; n24281
g21846 and pi0778 n24281_not ; n24282
g21847 nor pi0778 n24272 ; n24283
g21848 nor n24282 n24283 ; n24284
g21849 nor pi0609 n24284 ; n24285
g21850 nor pi1155 n24269 ; n24286
g21851 and n24285_not n24286 ; n24287
g21852 nor pi0660 n24216 ; n24288
g21853 and n24287_not n24288 ; n24289
g21854 and pi0609_not n24200 ; n24290
g21855 and pi0609 n24284_not ; n24291
g21856 and pi1155 n24290_not ; n24292
g21857 and n24291_not n24292 ; n24293
g21858 and pi0660 n24218_not ; n24294
g21859 and n24293_not n24294 ; n24295
g21860 nor n24289 n24295 ; n24296
g21861 and pi0785 n24296_not ; n24297
g21862 nor pi0785 n24284 ; n24298
g21863 nor n24297 n24298 ; n24299
g21864 nor pi0618 n24299 ; n24300
g21865 nor pi1154 n24268 ; n24301
g21866 and n24300_not n24301 ; n24302
g21867 nor pi0627 n24224 ; n24303
g21868 and n24302_not n24303 ; n24304
g21869 and pi0618_not n24201 ; n24305
g21870 and pi0618 n24299_not ; n24306
g21871 and pi1154 n24305_not ; n24307
g21872 and n24306_not n24307 ; n24308
g21873 and pi0627 n24226_not ; n24309
g21874 and n24308_not n24309 ; n24310
g21875 nor n24304 n24310 ; n24311
g21876 and pi0781 n24311_not ; n24312
g21877 nor pi0781 n24299 ; n24313
g21878 nor n24312 n24313 ; n24314
g21879 and pi0789_not n24314 ; n24315
g21880 nor pi0619 n24314 ; n24316
g21881 and pi0619 n24202 ; n24317
g21882 nor pi1159 n24317 ; n24318
g21883 and n24316_not n24318 ; n24319
g21884 nor pi0648 n24234 ; n24320
g21885 and n24319_not n24320 ; n24321
g21886 and pi0619 n24314_not ; n24322
g21887 and pi0619_not n24202 ; n24323
g21888 and pi1159 n24323_not ; n24324
g21889 and n24322_not n24324 ; n24325
g21890 and pi0648 n24238_not ; n24326
g21891 and n24325_not n24326 ; n24327
g21892 and pi0789 n24321_not ; n24328
g21893 and n24327_not n24328 ; n24329
g21894 and n17970 n24315_not ; n24330
g21895 and n24329_not n24330 ; n24331
g21896 nor n24267 n24331 ; n24332
g21897 nor n20364 n24332 ; n24333
g21898 and n17854 n24244_not ; n24334
g21899 and n20851 n24204 ; n24335
g21900 nor n24334 n24335 ; n24336
g21901 nor pi0629 n24336 ; n24337
g21902 and n20855 n24204 ; n24338
g21903 and n17853 n24244_not ; n24339
g21904 nor n24338 n24339 ; n24340
g21905 and pi0629 n24340_not ; n24341
g21906 nor n24337 n24341 ; n24342
g21907 and pi0792 n24342_not ; n24343
g21908 nor n20206 n24343 ; n24344
g21909 and n24333_not n24344 ; n24345
g21910 nor n24255 n24345 ; n24346
g21911 and pi0790_not n24346 ; n24347
g21912 nor pi0787 n24205 ; n24348
g21913 and pi1157 n24251_not ; n24349
g21914 nor n24209 n24349 ; n24350
g21915 and pi0787 n24350_not ; n24351
g21916 nor n24348 n24351 ; n24352
g21917 and pi0644_not n24352 ; n24353
g21918 and pi0644 n24346 ; n24354
g21919 and pi0715 n24353_not ; n24355
g21920 and n24354_not n24355 ; n24356
g21921 nor n17804 n24247 ; n24357
g21922 and n17804 n24189 ; n24358
g21923 nor n24357 n24358 ; n24359
g21924 and pi0644 n24359_not ; n24360
g21925 and pi0644_not n24189 ; n24361
g21926 nor pi0715 n24361 ; n24362
g21927 and n24360_not n24362 ; n24363
g21928 and pi1160 n24363_not ; n24364
g21929 and n24356_not n24364 ; n24365
g21930 nor pi0644 n24359 ; n24366
g21931 and pi0644 n24189 ; n24367
g21932 and pi0715 n24367_not ; n24368
g21933 and n24366_not n24368 ; n24369
g21934 and pi0644 n24352 ; n24370
g21935 and pi0644_not n24346 ; n24371
g21936 nor pi0715 n24370 ; n24372
g21937 and n24371_not n24372 ; n24373
g21938 nor pi1160 n24369 ; n24374
g21939 and n24373_not n24374 ; n24375
g21940 nor n24365 n24375 ; n24376
g21941 and pi0790 n24376_not ; n24377
g21942 and pi0832 n24347_not ; n24378
g21943 and n24377_not n24378 ; n24379
g21944 and pi0176_not po1038 ; n24380
g21945 nor pi0176 n17059 ; n24381
g21946 and n16635 n24381_not ; n24382
g21947 and pi0038_not n18076 ; n24383
g21948 and n2571 n16647_not ; n24384
g21949 and n24383_not n24384 ; n24385
g21950 and pi0176 n24385_not ; n24386
g21951 and pi0038_not n18072 ; n24387
g21952 nor n19899 n24387 ; n24388
g21953 and pi0176_not n24388 ; n24389
g21954 nor pi0704 n24389 ; n24390
g21955 nor pi0176 n17052 ; n24391
g21956 and pi0704 n24391 ; n24392
g21957 and n2571 n24392_not ; n24393
g21958 and n24390_not n24393 ; n24394
g21959 nor n24386 n24394 ; n24395
g21960 nor pi0778 n24395 ; n24396
g21961 and pi0625_not n24381 ; n24397
g21962 and pi0625 n24395 ; n24398
g21963 and pi1153 n24397_not ; n24399
g21964 and n24398_not n24399 ; n24400
g21965 and pi0625_not n24395 ; n24401
g21966 and pi0625 n24381 ; n24402
g21967 nor pi1153 n24402 ; n24403
g21968 and n24401_not n24403 ; n24404
g21969 nor n24400 n24404 ; n24405
g21970 and pi0778 n24405_not ; n24406
g21971 nor n24396 n24406 ; n24407
g21972 nor n17075 n24407 ; n24408
g21973 and n17075 n24381_not ; n24409
g21974 nor n24408 n24409 ; n24410
g21975 and n16639_not n24410 ; n24411
g21976 and n16639 n24381 ; n24412
g21977 nor n24411 n24412 ; n24413
g21978 and n16635_not n24413 ; n24414
g21979 nor n24382 n24414 ; n24415
g21980 and n16631_not n24415 ; n24416
g21981 and n16631 n24381 ; n24417
g21982 nor n24416 n24417 ; n24418
g21983 nor pi0628 n24418 ; n24419
g21984 and pi0628 n24381 ; n24420
g21985 nor n24419 n24420 ; n24421
g21986 nor pi1156 n24421 ; n24422
g21987 and pi0628 n24418_not ; n24423
g21988 and pi0628_not n24381 ; n24424
g21989 nor n24423 n24424 ; n24425
g21990 and pi1156 n24425_not ; n24426
g21991 nor n24422 n24426 ; n24427
g21992 and pi0792 n24427_not ; n24428
g21993 nor pi0792 n24418 ; n24429
g21994 nor n24428 n24429 ; n24430
g21995 nor pi0647 n24430 ; n24431
g21996 and pi0647 n24381 ; n24432
g21997 nor n24431 n24432 ; n24433
g21998 nor pi1157 n24433 ; n24434
g21999 and pi0647 n24430_not ; n24435
g22000 and pi0647_not n24381 ; n24436
g22001 nor n24435 n24436 ; n24437
g22002 and pi1157 n24437_not ; n24438
g22003 nor n24434 n24438 ; n24439
g22004 and pi0787 n24439_not ; n24440
g22005 nor pi0787 n24430 ; n24441
g22006 nor n24440 n24441 ; n24442
g22007 nor pi0644 n24442 ; n24443
g22008 and pi0715 n24443_not ; n24444
g22009 and pi0176 n2571_not ; n24445
g22010 and pi0176_not n19439 ; n24446
g22011 nor n19433 n19434 ; n24447
g22012 and pi0176 n24447 ; n24448
g22013 nor n24446 n24448 ; n24449
g22014 nor pi0742 n24449 ; n24450
g22015 and pi0742 n24391_not ; n24451
g22016 nor n24450 n24451 ; n24452
g22017 and n2571 n24452_not ; n24453
g22018 nor n24445 n24453 ; n24454
g22019 nor n17117 n24454 ; n24455
g22020 and n17117 n24381_not ; n24456
g22021 nor n24455 n24456 ; n24457
g22022 nor pi0785 n24457 ; n24458
g22023 nor n17291 n24381 ; n24459
g22024 and pi0609 n24455 ; n24460
g22025 nor n24459 n24460 ; n24461
g22026 and pi1155 n24461_not ; n24462
g22027 nor n17296 n24381 ; n24463
g22028 and pi0609_not n24455 ; n24464
g22029 nor n24463 n24464 ; n24465
g22030 nor pi1155 n24465 ; n24466
g22031 nor n24462 n24466 ; n24467
g22032 and pi0785 n24467_not ; n24468
g22033 nor n24458 n24468 ; n24469
g22034 nor pi0781 n24469 ; n24470
g22035 and pi0618_not n24381 ; n24471
g22036 and pi0618 n24469 ; n24472
g22037 and pi1154 n24471_not ; n24473
g22038 and n24472_not n24473 ; n24474
g22039 and pi0618_not n24469 ; n24475
g22040 and pi0618 n24381 ; n24476
g22041 nor pi1154 n24476 ; n24477
g22042 and n24475_not n24477 ; n24478
g22043 nor n24474 n24478 ; n24479
g22044 and pi0781 n24479_not ; n24480
g22045 nor n24470 n24480 ; n24481
g22046 nor pi0789 n24481 ; n24482
g22047 and pi0619_not n24381 ; n24483
g22048 and pi0619 n24481 ; n24484
g22049 and pi1159 n24483_not ; n24485
g22050 and n24484_not n24485 ; n24486
g22051 and pi0619_not n24481 ; n24487
g22052 and pi0619 n24381 ; n24488
g22053 nor pi1159 n24488 ; n24489
g22054 and n24487_not n24489 ; n24490
g22055 nor n24486 n24490 ; n24491
g22056 and pi0789 n24491_not ; n24492
g22057 nor n24482 n24492 ; n24493
g22058 and n17969_not n24493 ; n24494
g22059 and n17969 n24381 ; n24495
g22060 nor n24494 n24495 ; n24496
g22061 nor n17779 n24496 ; n24497
g22062 and n17779 n24381 ; n24498
g22063 nor n24497 n24498 ; n24499
g22064 nor n17804 n24499 ; n24500
g22065 and n17804 n24381 ; n24501
g22066 nor n24500 n24501 ; n24502
g22067 and pi0644 n24502_not ; n24503
g22068 and pi0644_not n24381 ; n24504
g22069 nor pi0715 n24504 ; n24505
g22070 and n24503_not n24505 ; n24506
g22071 and pi1160 n24506_not ; n24507
g22072 and n24444_not n24507 ; n24508
g22073 and pi0644 n24442_not ; n24509
g22074 nor pi0715 n24509 ; n24510
g22075 nor pi0644 n24502 ; n24511
g22076 and pi0644 n24381 ; n24512
g22077 and pi0715 n24512_not ; n24513
g22078 and n24511_not n24513 ; n24514
g22079 nor pi1160 n24514 ; n24515
g22080 and n24510_not n24515 ; n24516
g22081 nor n24508 n24516 ; n24517
g22082 and pi0790 n24517_not ; n24518
g22083 and n17802 n24433 ; n24519
g22084 and n20559_not n24499 ; n24520
g22085 and n17801 n24437 ; n24521
g22086 nor n24519 n24520 ; n24522
g22087 and n24521_not n24522 ; n24523
g22088 and pi0787 n24523_not ; n24524
g22089 and n17777 n24421 ; n24525
g22090 and n20570_not n24496 ; n24526
g22091 and n17776 n24425 ; n24527
g22092 nor n24525 n24527 ; n24528
g22093 and n24526_not n24528 ; n24529
g22094 and pi0792 n24529_not ; n24530
g22095 and n17871 n24415 ; n24531
g22096 nor pi0626 n24493 ; n24532
g22097 and pi0626 n24381_not ; n24533
g22098 and n16629 n24533_not ; n24534
g22099 and n24532_not n24534 ; n24535
g22100 and pi0626 n24493_not ; n24536
g22101 nor pi0626 n24381 ; n24537
g22102 and n16628 n24537_not ; n24538
g22103 and n24536_not n24538 ; n24539
g22104 nor n24531 n24535 ; n24540
g22105 and n24539_not n24540 ; n24541
g22106 and pi0788 n24541_not ; n24542
g22107 and pi0609 n24407 ; n24543
g22108 nor pi0176 n19488 ; n24544
g22109 and pi0176 n19496 ; n24545
g22110 nor pi0742 n24544 ; n24546
g22111 and n24545_not n24546 ; n24547
g22112 and pi0176_not n19477 ; n24548
g22113 nor n19468 n19470 ; n24549
g22114 and pi0176 n24549_not ; n24550
g22115 and pi0742 n24550_not ; n24551
g22116 and n24548_not n24551 ; n24552
g22117 nor pi0704 n24547 ; n24553
g22118 and n24552_not n24553 ; n24554
g22119 and pi0704 n24452 ; n24555
g22120 and n2571 n24554_not ; n24556
g22121 and n24555_not n24556 ; n24557
g22122 nor n24445 n24557 ; n24558
g22123 and pi0625_not n24558 ; n24559
g22124 and pi0625 n24454 ; n24560
g22125 nor pi1153 n24560 ; n24561
g22126 and n24559_not n24561 ; n24562
g22127 nor pi0608 n24400 ; n24563
g22128 and n24562_not n24563 ; n24564
g22129 and pi0625_not n24454 ; n24565
g22130 and pi0625 n24558 ; n24566
g22131 and pi1153 n24565_not ; n24567
g22132 and n24566_not n24567 ; n24568
g22133 and pi0608 n24404_not ; n24569
g22134 and n24568_not n24569 ; n24570
g22135 nor n24564 n24570 ; n24571
g22136 and pi0778 n24571_not ; n24572
g22137 and pi0778_not n24558 ; n24573
g22138 nor n24572 n24573 ; n24574
g22139 nor pi0609 n24574 ; n24575
g22140 nor pi1155 n24543 ; n24576
g22141 and n24575_not n24576 ; n24577
g22142 nor pi0660 n24462 ; n24578
g22143 and n24577_not n24578 ; n24579
g22144 and pi0609_not n24407 ; n24580
g22145 and pi0609 n24574_not ; n24581
g22146 and pi1155 n24580_not ; n24582
g22147 and n24581_not n24582 ; n24583
g22148 and pi0660 n24466_not ; n24584
g22149 and n24583_not n24584 ; n24585
g22150 nor n24579 n24585 ; n24586
g22151 and pi0785 n24586_not ; n24587
g22152 nor pi0785 n24574 ; n24588
g22153 nor n24587 n24588 ; n24589
g22154 nor pi0618 n24589 ; n24590
g22155 and pi0618 n24410 ; n24591
g22156 nor pi1154 n24591 ; n24592
g22157 and n24590_not n24592 ; n24593
g22158 nor pi0627 n24474 ; n24594
g22159 and n24593_not n24594 ; n24595
g22160 and pi0618_not n24410 ; n24596
g22161 and pi0618 n24589_not ; n24597
g22162 and pi1154 n24596_not ; n24598
g22163 and n24597_not n24598 ; n24599
g22164 and pi0627 n24478_not ; n24600
g22165 and n24599_not n24600 ; n24601
g22166 nor n24595 n24601 ; n24602
g22167 and pi0781 n24602_not ; n24603
g22168 nor pi0781 n24589 ; n24604
g22169 nor n24603 n24604 ; n24605
g22170 and pi0789_not n24605 ; n24606
g22171 and pi0619 n24413_not ; n24607
g22172 nor pi0619 n24605 ; n24608
g22173 nor pi1159 n24607 ; n24609
g22174 and n24608_not n24609 ; n24610
g22175 nor pi0648 n24486 ; n24611
g22176 and n24610_not n24611 ; n24612
g22177 and pi0619 n24605_not ; n24613
g22178 nor pi0619 n24413 ; n24614
g22179 and pi1159 n24614_not ; n24615
g22180 and n24613_not n24615 ; n24616
g22181 and pi0648 n24490_not ; n24617
g22182 and n24616_not n24617 ; n24618
g22183 and pi0789 n24612_not ; n24619
g22184 and n24618_not n24619 ; n24620
g22185 and n17970 n24606_not ; n24621
g22186 and n24620_not n24621 ; n24622
g22187 nor n24542 n24622 ; n24623
g22188 nor n24530 n24623 ; n24624
g22189 and n20364 n24529 ; n24625
g22190 nor n20206 n24625 ; n24626
g22191 and n24624_not n24626 ; n24627
g22192 and pi0644_not n24515 ; n24628
g22193 and pi0644 n24507 ; n24629
g22194 and pi0790 n24628_not ; n24630
g22195 and n24629_not n24630 ; n24631
g22196 nor n24524 n24627 ; n24632
g22197 and n24631_not n24632 ; n24633
g22198 nor n24518 n24633 ; n24634
g22199 nor po1038 n24634 ; n24635
g22200 nor pi0832 n24380 ; n24636
g22201 and n24635_not n24636 ; n24637
g22202 nor n24379 n24637 ; po0333
g22203 nor pi0177 n17059 ; n24639
g22204 and n16635 n24639_not ; n24640
g22205 and pi0177 n2571_not ; n24641
g22206 and pi0177_not n18072 ; n24642
g22207 and pi0177 n18076_not ; n24643
g22208 nor pi0038 n24643 ; n24644
g22209 and n24642_not n24644 ; n24645
g22210 nor pi0177 n16641 ; n24646
g22211 and n16647 n24646_not ; n24647
g22212 nor pi0686 n24647 ; n24648
g22213 and n24645_not n24648 ; n24649
g22214 and pi0177_not pi0686 ; n24650
g22215 and n17052_not n24650 ; n24651
g22216 and n2571 n24651_not ; n24652
g22217 and n24649_not n24652 ; n24653
g22218 nor n24641 n24653 ; n24654
g22219 nor pi0778 n24654 ; n24655
g22220 and pi0625_not n24639 ; n24656
g22221 and pi0625 n24654 ; n24657
g22222 and pi1153 n24656_not ; n24658
g22223 and n24657_not n24658 ; n24659
g22224 and pi0625_not n24654 ; n24660
g22225 and pi0625 n24639 ; n24661
g22226 nor pi1153 n24661 ; n24662
g22227 and n24660_not n24662 ; n24663
g22228 nor n24659 n24663 ; n24664
g22229 and pi0778 n24664_not ; n24665
g22230 nor n24655 n24665 ; n24666
g22231 nor n17075 n24666 ; n24667
g22232 and n17075 n24639_not ; n24668
g22233 nor n24667 n24668 ; n24669
g22234 and n16639_not n24669 ; n24670
g22235 and n16639 n24639 ; n24671
g22236 nor n24670 n24671 ; n24672
g22237 and n16635_not n24672 ; n24673
g22238 nor n24640 n24673 ; n24674
g22239 and n16631_not n24674 ; n24675
g22240 and n16631 n24639 ; n24676
g22241 nor n24675 n24676 ; n24677
g22242 and pi0792_not n24677 ; n24678
g22243 and pi0628_not n24639 ; n24679
g22244 and pi0628 n24677_not ; n24680
g22245 and pi1156 n24679_not ; n24681
g22246 and n24680_not n24681 ; n24682
g22247 and pi0628 n24639 ; n24683
g22248 nor pi0628 n24677 ; n24684
g22249 nor pi1156 n24683 ; n24685
g22250 and n24684_not n24685 ; n24686
g22251 nor n24682 n24686 ; n24687
g22252 and pi0792 n24687_not ; n24688
g22253 nor n24678 n24688 ; n24689
g22254 nor pi0787 n24689 ; n24690
g22255 and pi0647_not n24639 ; n24691
g22256 and pi0647 n24689 ; n24692
g22257 and pi1157 n24691_not ; n24693
g22258 and n24692_not n24693 ; n24694
g22259 and pi0647_not n24689 ; n24695
g22260 and pi0647 n24639 ; n24696
g22261 nor pi1157 n24696 ; n24697
g22262 and n24695_not n24697 ; n24698
g22263 nor n24694 n24698 ; n24699
g22264 and pi0787 n24699_not ; n24700
g22265 nor n24690 n24700 ; n24701
g22266 and pi0644_not n24701 ; n24702
g22267 and pi0619_not n24639 ; n24703
g22268 nor pi0757 n19439 ; n24704
g22269 nor n21646 n24704 ; n24705
g22270 nor pi0177 n24705 ; n24706
g22271 nor pi0177 n19433 ; n24707
g22272 nor pi0757 n24707 ; n24708
g22273 and n24447_not n24708 ; n24709
g22274 nor n24706 n24709 ; n24710
g22275 and n2571 n24710 ; n24711
g22276 nor n24641 n24711 ; n24712
g22277 nor n17117 n24712 ; n24713
g22278 and n17117 n24639_not ; n24714
g22279 nor n24713 n24714 ; n24715
g22280 nor pi0785 n24715 ; n24716
g22281 nor n17291 n24639 ; n24717
g22282 and pi0609 n24713 ; n24718
g22283 nor n24717 n24718 ; n24719
g22284 and pi1155 n24719_not ; n24720
g22285 nor n17296 n24639 ; n24721
g22286 and pi0609_not n24713 ; n24722
g22287 nor n24721 n24722 ; n24723
g22288 nor pi1155 n24723 ; n24724
g22289 nor n24720 n24724 ; n24725
g22290 and pi0785 n24725_not ; n24726
g22291 nor n24716 n24726 ; n24727
g22292 nor pi0781 n24727 ; n24728
g22293 and pi0618_not n24639 ; n24729
g22294 and pi0618 n24727 ; n24730
g22295 and pi1154 n24729_not ; n24731
g22296 and n24730_not n24731 ; n24732
g22297 and pi0618_not n24727 ; n24733
g22298 and pi0618 n24639 ; n24734
g22299 nor pi1154 n24734 ; n24735
g22300 and n24733_not n24735 ; n24736
g22301 nor n24732 n24736 ; n24737
g22302 and pi0781 n24737_not ; n24738
g22303 nor n24728 n24738 ; n24739
g22304 and pi0619 n24739 ; n24740
g22305 and pi1159 n24703_not ; n24741
g22306 and n24740_not n24741 ; n24742
g22307 and n18176 n24646_not ; n24743
g22308 and pi0177_not n19475 ; n24744
g22309 and pi0177 n19467 ; n24745
g22310 nor pi0038 n24745 ; n24746
g22311 and n24744_not n24746 ; n24747
g22312 and pi0757 n24743_not ; n24748
g22313 and n24747_not n24748 ; n24749
g22314 nor pi0177 n19485 ; n24750
g22315 and pi0177 n19490 ; n24751
g22316 and pi0038 n24751_not ; n24752
g22317 and n24750_not n24752 ; n24753
g22318 nor n19482 n19484 ; n24754
g22319 nor pi0177 n24754 ; n24755
g22320 and pi0177 n19494 ; n24756
g22321 nor pi0038 n24755 ; n24757
g22322 and n24756_not n24757 ; n24758
g22323 nor pi0757 n24753 ; n24759
g22324 and n24758_not n24759 ; n24760
g22325 nor n24749 n24760 ; n24761
g22326 nor pi0686 n24761 ; n24762
g22327 and pi0686 n24710_not ; n24763
g22328 and n2571 n24762_not ; n24764
g22329 and n24763_not n24764 ; n24765
g22330 nor n24641 n24765 ; n24766
g22331 and pi0625_not n24766 ; n24767
g22332 and pi0625 n24712 ; n24768
g22333 nor pi1153 n24768 ; n24769
g22334 and n24767_not n24769 ; n24770
g22335 nor pi0608 n24659 ; n24771
g22336 and n24770_not n24771 ; n24772
g22337 and pi0625_not n24712 ; n24773
g22338 and pi0625 n24766 ; n24774
g22339 and pi1153 n24773_not ; n24775
g22340 and n24774_not n24775 ; n24776
g22341 and pi0608 n24663_not ; n24777
g22342 and n24776_not n24777 ; n24778
g22343 nor n24772 n24778 ; n24779
g22344 and pi0778 n24779_not ; n24780
g22345 and pi0778_not n24766 ; n24781
g22346 nor n24780 n24781 ; n24782
g22347 nor pi0609 n24782 ; n24783
g22348 and pi0609 n24666 ; n24784
g22349 nor pi1155 n24784 ; n24785
g22350 and n24783_not n24785 ; n24786
g22351 nor pi0660 n24720 ; n24787
g22352 and n24786_not n24787 ; n24788
g22353 and pi0609_not n24666 ; n24789
g22354 and pi0609 n24782_not ; n24790
g22355 and pi1155 n24789_not ; n24791
g22356 and n24790_not n24791 ; n24792
g22357 and pi0660 n24724_not ; n24793
g22358 and n24792_not n24793 ; n24794
g22359 nor n24788 n24794 ; n24795
g22360 and pi0785 n24795_not ; n24796
g22361 nor pi0785 n24782 ; n24797
g22362 nor n24796 n24797 ; n24798
g22363 nor pi0618 n24798 ; n24799
g22364 and pi0618 n24669 ; n24800
g22365 nor pi1154 n24800 ; n24801
g22366 and n24799_not n24801 ; n24802
g22367 nor pi0627 n24732 ; n24803
g22368 and n24802_not n24803 ; n24804
g22369 and pi0618_not n24669 ; n24805
g22370 and pi0618 n24798_not ; n24806
g22371 and pi1154 n24805_not ; n24807
g22372 and n24806_not n24807 ; n24808
g22373 and pi0627 n24736_not ; n24809
g22374 and n24808_not n24809 ; n24810
g22375 nor n24804 n24810 ; n24811
g22376 and pi0781 n24811_not ; n24812
g22377 nor pi0781 n24798 ; n24813
g22378 nor n24812 n24813 ; n24814
g22379 nor pi0619 n24814 ; n24815
g22380 and pi0619 n24672_not ; n24816
g22381 nor pi1159 n24816 ; n24817
g22382 and n24815_not n24817 ; n24818
g22383 nor pi0648 n24742 ; n24819
g22384 and n24818_not n24819 ; n24820
g22385 and pi0619_not n24739 ; n24821
g22386 and pi0619 n24639 ; n24822
g22387 nor pi1159 n24822 ; n24823
g22388 and n24821_not n24823 ; n24824
g22389 and pi0619 n24814_not ; n24825
g22390 nor pi0619 n24672 ; n24826
g22391 and pi1159 n24826_not ; n24827
g22392 and n24825_not n24827 ; n24828
g22393 and pi0648 n24824_not ; n24829
g22394 and n24828_not n24829 ; n24830
g22395 nor n24820 n24830 ; n24831
g22396 and pi0789 n24831_not ; n24832
g22397 nor pi0789 n24814 ; n24833
g22398 nor n24832 n24833 ; n24834
g22399 and pi0788_not n24834 ; n24835
g22400 and pi0626_not n24834 ; n24836
g22401 and pi0626 n24674_not ; n24837
g22402 nor pi0641 n24837 ; n24838
g22403 and n24836_not n24838 ; n24839
g22404 nor pi0789 n24739 ; n24840
g22405 nor n24742 n24824 ; n24841
g22406 and pi0789 n24841_not ; n24842
g22407 nor n24840 n24842 ; n24843
g22408 nor pi0626 n24843 ; n24844
g22409 and pi0626 n24639_not ; n24845
g22410 and pi0641 n24845_not ; n24846
g22411 and n24844_not n24846 ; n24847
g22412 nor pi1158 n24847 ; n24848
g22413 and n24839_not n24848 ; n24849
g22414 and pi0626 n24834 ; n24850
g22415 nor pi0626 n24674 ; n24851
g22416 and pi0641 n24851_not ; n24852
g22417 and n24850_not n24852 ; n24853
g22418 and pi0626 n24843_not ; n24854
g22419 nor pi0626 n24639 ; n24855
g22420 nor pi0641 n24855 ; n24856
g22421 and n24854_not n24856 ; n24857
g22422 and pi1158 n24857_not ; n24858
g22423 and n24853_not n24858 ; n24859
g22424 nor n24849 n24859 ; n24860
g22425 and pi0788 n24860_not ; n24861
g22426 nor n24835 n24861 ; n24862
g22427 and pi0628_not n24862 ; n24863
g22428 and n17969_not n24843 ; n24864
g22429 and n17969 n24639 ; n24865
g22430 nor n24864 n24865 ; n24866
g22431 and pi0628 n24866_not ; n24867
g22432 nor pi1156 n24867 ; n24868
g22433 and n24863_not n24868 ; n24869
g22434 nor pi0629 n24682 ; n24870
g22435 and n24869_not n24870 ; n24871
g22436 and pi0628 n24862 ; n24872
g22437 nor pi0628 n24866 ; n24873
g22438 and pi1156 n24873_not ; n24874
g22439 and n24872_not n24874 ; n24875
g22440 and pi0629 n24686_not ; n24876
g22441 and n24875_not n24876 ; n24877
g22442 nor n24871 n24877 ; n24878
g22443 and pi0792 n24878_not ; n24879
g22444 and pi0792_not n24862 ; n24880
g22445 nor n24879 n24880 ; n24881
g22446 nor pi0647 n24881 ; n24882
g22447 nor n17779 n24866 ; n24883
g22448 and n17779 n24639 ; n24884
g22449 nor n24883 n24884 ; n24885
g22450 and pi0647 n24885_not ; n24886
g22451 nor pi1157 n24886 ; n24887
g22452 and n24882_not n24887 ; n24888
g22453 nor pi0630 n24694 ; n24889
g22454 and n24888_not n24889 ; n24890
g22455 and pi0647 n24881_not ; n24891
g22456 nor pi0647 n24885 ; n24892
g22457 and pi1157 n24892_not ; n24893
g22458 and n24891_not n24893 ; n24894
g22459 and pi0630 n24698_not ; n24895
g22460 and n24894_not n24895 ; n24896
g22461 nor n24890 n24896 ; n24897
g22462 and pi0787 n24897_not ; n24898
g22463 nor pi0787 n24881 ; n24899
g22464 nor n24898 n24899 ; n24900
g22465 and pi0644 n24900_not ; n24901
g22466 and pi0715 n24702_not ; n24902
g22467 and n24901_not n24902 ; n24903
g22468 and n17804 n24639_not ; n24904
g22469 and n17804_not n24885 ; n24905
g22470 nor n24904 n24905 ; n24906
g22471 and pi0644 n24906 ; n24907
g22472 and pi0644_not n24639 ; n24908
g22473 nor pi0715 n24908 ; n24909
g22474 and n24907_not n24909 ; n24910
g22475 and pi1160 n24910_not ; n24911
g22476 and n24903_not n24911 ; n24912
g22477 nor pi0644 n24900 ; n24913
g22478 and pi0644 n24701 ; n24914
g22479 nor pi0715 n24914 ; n24915
g22480 and n24913_not n24915 ; n24916
g22481 and pi0644_not n24906 ; n24917
g22482 and pi0644 n24639 ; n24918
g22483 and pi0715 n24918_not ; n24919
g22484 and n24917_not n24919 ; n24920
g22485 nor pi1160 n24920 ; n24921
g22486 and n24916_not n24921 ; n24922
g22487 and pi0790 n24912_not ; n24923
g22488 and n24922_not n24923 ; n24924
g22489 and pi0790_not n24900 ; n24925
g22490 nor po1038 n24925 ; n24926
g22491 and n24924_not n24926 ; n24927
g22492 and pi0177_not po1038 ; n24928
g22493 nor pi0832 n24928 ; n24929
g22494 and n24927_not n24929 ; n24930
g22495 nor pi0177 n2926 ; n24931
g22496 and pi0686_not n16645 ; n24932
g22497 nor n24931 n24932 ; n24933
g22498 and pi0778_not n24933 ; n24934
g22499 and pi0625_not n24932 ; n24935
g22500 nor n24933 n24935 ; n24936
g22501 and pi1153 n24936_not ; n24937
g22502 nor pi1153 n24931 ; n24938
g22503 and n24935_not n24938 ; n24939
g22504 nor n24937 n24939 ; n24940
g22505 and pi0778 n24940_not ; n24941
g22506 nor n24934 n24941 ; n24942
g22507 and n17845_not n24942 ; n24943
g22508 and n17847_not n24943 ; n24944
g22509 and n17849_not n24944 ; n24945
g22510 and n17851_not n24945 ; n24946
g22511 and n17857_not n24946 ; n24947
g22512 and pi0647_not n24947 ; n24948
g22513 and pi0647 n24931 ; n24949
g22514 nor pi1157 n24949 ; n24950
g22515 and n24948_not n24950 ; n24951
g22516 and pi0630 n24951 ; n24952
g22517 and pi0757_not n17244 ; n24953
g22518 nor n24931 n24953 ; n24954
g22519 nor n17874 n24954 ; n24955
g22520 nor pi0785 n24955 ; n24956
g22521 nor n17879 n24954 ; n24957
g22522 and pi1155 n24957_not ; n24958
g22523 and n17882_not n24955 ; n24959
g22524 nor pi1155 n24959 ; n24960
g22525 nor n24958 n24960 ; n24961
g22526 and pi0785 n24961_not ; n24962
g22527 nor n24956 n24962 ; n24963
g22528 nor pi0781 n24963 ; n24964
g22529 and n17889_not n24963 ; n24965
g22530 and pi1154 n24965_not ; n24966
g22531 and n17892_not n24963 ; n24967
g22532 nor pi1154 n24967 ; n24968
g22533 nor n24966 n24968 ; n24969
g22534 and pi0781 n24969_not ; n24970
g22535 nor n24964 n24970 ; n24971
g22536 nor pi0789 n24971 ; n24972
g22537 and pi0619_not n24931 ; n24973
g22538 and pi0619 n24971 ; n24974
g22539 and pi1159 n24973_not ; n24975
g22540 and n24974_not n24975 ; n24976
g22541 and pi0619_not n24971 ; n24977
g22542 and pi0619 n24931 ; n24978
g22543 nor pi1159 n24978 ; n24979
g22544 and n24977_not n24979 ; n24980
g22545 nor n24976 n24980 ; n24981
g22546 and pi0789 n24981_not ; n24982
g22547 nor n24972 n24982 ; n24983
g22548 and n17969_not n24983 ; n24984
g22549 and n17969 n24931 ; n24985
g22550 nor n24984 n24985 ; n24986
g22551 nor n17779 n24986 ; n24987
g22552 and n17779 n24931 ; n24988
g22553 nor n24987 n24988 ; n24989
g22554 and n20559_not n24989 ; n24990
g22555 and pi0647 n24947_not ; n24991
g22556 nor pi0647 n24931 ; n24992
g22557 nor n24991 n24992 ; n24993
g22558 and n17801 n24993_not ; n24994
g22559 nor n24952 n24994 ; n24995
g22560 and n24990_not n24995 ; n24996
g22561 and pi0787 n24996_not ; n24997
g22562 and n17871 n24945 ; n24998
g22563 nor pi0626 n24983 ; n24999
g22564 and pi0626 n24931_not ; n25000
g22565 and n16629 n25000_not ; n25001
g22566 and n24999_not n25001 ; n25002
g22567 and pi0626 n24983_not ; n25003
g22568 nor pi0626 n24931 ; n25004
g22569 and n16628 n25004_not ; n25005
g22570 and n25003_not n25005 ; n25006
g22571 nor n24998 n25002 ; n25007
g22572 and n25006_not n25007 ; n25008
g22573 and pi0788 n25008_not ; n25009
g22574 and pi0618 n24943 ; n25010
g22575 and pi0609 n24942 ; n25011
g22576 nor n17168 n24933 ; n25012
g22577 and pi0625 n25012 ; n25013
g22578 and n24954 n25012_not ; n25014
g22579 nor n25013 n25014 ; n25015
g22580 and n24938 n25015_not ; n25016
g22581 nor pi0608 n24937 ; n25017
g22582 and n25016_not n25017 ; n25018
g22583 and pi1153 n24954 ; n25019
g22584 and n25013_not n25019 ; n25020
g22585 and pi0608 n24939_not ; n25021
g22586 and n25020_not n25021 ; n25022
g22587 nor n25018 n25022 ; n25023
g22588 and pi0778 n25023_not ; n25024
g22589 nor pi0778 n25014 ; n25025
g22590 nor n25024 n25025 ; n25026
g22591 nor pi0609 n25026 ; n25027
g22592 nor pi1155 n25011 ; n25028
g22593 and n25027_not n25028 ; n25029
g22594 nor pi0660 n24958 ; n25030
g22595 and n25029_not n25030 ; n25031
g22596 and pi0609_not n24942 ; n25032
g22597 and pi0609 n25026_not ; n25033
g22598 and pi1155 n25032_not ; n25034
g22599 and n25033_not n25034 ; n25035
g22600 and pi0660 n24960_not ; n25036
g22601 and n25035_not n25036 ; n25037
g22602 nor n25031 n25037 ; n25038
g22603 and pi0785 n25038_not ; n25039
g22604 nor pi0785 n25026 ; n25040
g22605 nor n25039 n25040 ; n25041
g22606 nor pi0618 n25041 ; n25042
g22607 nor pi1154 n25010 ; n25043
g22608 and n25042_not n25043 ; n25044
g22609 nor pi0627 n24966 ; n25045
g22610 and n25044_not n25045 ; n25046
g22611 and pi0618_not n24943 ; n25047
g22612 and pi0618 n25041_not ; n25048
g22613 and pi1154 n25047_not ; n25049
g22614 and n25048_not n25049 ; n25050
g22615 and pi0627 n24968_not ; n25051
g22616 and n25050_not n25051 ; n25052
g22617 nor n25046 n25052 ; n25053
g22618 and pi0781 n25053_not ; n25054
g22619 nor pi0781 n25041 ; n25055
g22620 nor n25054 n25055 ; n25056
g22621 and pi0789_not n25056 ; n25057
g22622 nor pi0619 n25056 ; n25058
g22623 and pi0619 n24944 ; n25059
g22624 nor pi1159 n25059 ; n25060
g22625 and n25058_not n25060 ; n25061
g22626 nor pi0648 n24976 ; n25062
g22627 and n25061_not n25062 ; n25063
g22628 and pi0619 n25056_not ; n25064
g22629 and pi0619_not n24944 ; n25065
g22630 and pi1159 n25065_not ; n25066
g22631 and n25064_not n25066 ; n25067
g22632 and pi0648 n24980_not ; n25068
g22633 and n25067_not n25068 ; n25069
g22634 and pi0789 n25063_not ; n25070
g22635 and n25069_not n25070 ; n25071
g22636 and n17970 n25057_not ; n25072
g22637 and n25071_not n25072 ; n25073
g22638 nor n25009 n25073 ; n25074
g22639 nor n20364 n25074 ; n25075
g22640 and n17854 n24986_not ; n25076
g22641 and n20851 n24946 ; n25077
g22642 nor n25076 n25077 ; n25078
g22643 nor pi0629 n25078 ; n25079
g22644 and n20855 n24946 ; n25080
g22645 and n17853 n24986_not ; n25081
g22646 nor n25080 n25081 ; n25082
g22647 and pi0629 n25082_not ; n25083
g22648 nor n25079 n25083 ; n25084
g22649 and pi0792 n25084_not ; n25085
g22650 nor n20206 n25085 ; n25086
g22651 and n25075_not n25086 ; n25087
g22652 nor n24997 n25087 ; n25088
g22653 and pi0790_not n25088 ; n25089
g22654 nor pi0787 n24947 ; n25090
g22655 and pi1157 n24993_not ; n25091
g22656 nor n24951 n25091 ; n25092
g22657 and pi0787 n25092_not ; n25093
g22658 nor n25090 n25093 ; n25094
g22659 and pi0644_not n25094 ; n25095
g22660 and pi0644 n25088 ; n25096
g22661 and pi0715 n25095_not ; n25097
g22662 and n25096_not n25097 ; n25098
g22663 nor n17804 n24989 ; n25099
g22664 and n17804 n24931 ; n25100
g22665 nor n25099 n25100 ; n25101
g22666 and pi0644 n25101_not ; n25102
g22667 and pi0644_not n24931 ; n25103
g22668 nor pi0715 n25103 ; n25104
g22669 and n25102_not n25104 ; n25105
g22670 and pi1160 n25105_not ; n25106
g22671 and n25098_not n25106 ; n25107
g22672 nor pi0644 n25101 ; n25108
g22673 and pi0644 n24931 ; n25109
g22674 and pi0715 n25109_not ; n25110
g22675 and n25108_not n25110 ; n25111
g22676 and pi0644 n25094 ; n25112
g22677 and pi0644_not n25088 ; n25113
g22678 nor pi0715 n25112 ; n25114
g22679 and n25113_not n25114 ; n25115
g22680 nor pi1160 n25111 ; n25116
g22681 and n25115_not n25116 ; n25117
g22682 nor n25107 n25117 ; n25118
g22683 and pi0790 n25118_not ; n25119
g22684 and pi0832 n25089_not ; n25120
g22685 and n25119_not n25120 ; n25121
g22686 nor n24930 n25121 ; po0334
g22687 nor pi0178 n2926 ; n25123
g22688 and pi0688_not n16645 ; n25124
g22689 nor n25123 n25124 ; n25125
g22690 nor pi0778 n25125 ; n25126
g22691 and pi0625_not n25124 ; n25127
g22692 nor n25125 n25127 ; n25128
g22693 and pi1153 n25128_not ; n25129
g22694 nor pi1153 n25123 ; n25130
g22695 and n25127_not n25130 ; n25131
g22696 and pi0778 n25131_not ; n25132
g22697 and n25129_not n25132 ; n25133
g22698 nor n25126 n25133 ; n25134
g22699 nor n17845 n25134 ; n25135
g22700 and n17847_not n25135 ; n25136
g22701 and n17849_not n25136 ; n25137
g22702 and n17851_not n25137 ; n25138
g22703 and n17857_not n25138 ; n25139
g22704 and pi0647_not n25139 ; n25140
g22705 and pi0647 n25123 ; n25141
g22706 nor pi1157 n25141 ; n25142
g22707 and n25140_not n25142 ; n25143
g22708 and pi0630 n25143 ; n25144
g22709 and pi0760_not n17244 ; n25145
g22710 nor n25123 n25145 ; n25146
g22711 nor n17874 n25146 ; n25147
g22712 nor pi0785 n25147 ; n25148
g22713 and n17296 n25145 ; n25149
g22714 and n25147 n25149_not ; n25150
g22715 and pi1155 n25150_not ; n25151
g22716 nor pi1155 n25123 ; n25152
g22717 and n25149_not n25152 ; n25153
g22718 nor n25151 n25153 ; n25154
g22719 and pi0785 n25154_not ; n25155
g22720 nor n25148 n25155 ; n25156
g22721 nor pi0781 n25156 ; n25157
g22722 and n17889_not n25156 ; n25158
g22723 and pi1154 n25158_not ; n25159
g22724 and n17892_not n25156 ; n25160
g22725 nor pi1154 n25160 ; n25161
g22726 nor n25159 n25161 ; n25162
g22727 and pi0781 n25162_not ; n25163
g22728 nor n25157 n25163 ; n25164
g22729 nor pi0789 n25164 ; n25165
g22730 and n23078_not n25164 ; n25166
g22731 and pi1159 n25166_not ; n25167
g22732 and n23081_not n25164 ; n25168
g22733 nor pi1159 n25168 ; n25169
g22734 nor n25167 n25169 ; n25170
g22735 and pi0789 n25170_not ; n25171
g22736 nor n25165 n25171 ; n25172
g22737 and n17969_not n25172 ; n25173
g22738 and n17969 n25123 ; n25174
g22739 nor n25173 n25174 ; n25175
g22740 nor n17779 n25175 ; n25176
g22741 and n17779 n25123 ; n25177
g22742 nor n25176 n25177 ; n25178
g22743 and n20559_not n25178 ; n25179
g22744 and pi0647 n25139_not ; n25180
g22745 nor pi0647 n25123 ; n25181
g22746 nor n25180 n25181 ; n25182
g22747 and n17801 n25182_not ; n25183
g22748 nor n25144 n25183 ; n25184
g22749 and n25179_not n25184 ; n25185
g22750 and pi0787 n25185_not ; n25186
g22751 and n17871 n25137 ; n25187
g22752 nor pi0626 n25172 ; n25188
g22753 and pi0626 n25123_not ; n25189
g22754 and n16629 n25189_not ; n25190
g22755 and n25188_not n25190 ; n25191
g22756 and pi0626 n25172_not ; n25192
g22757 nor pi0626 n25123 ; n25193
g22758 and n16628 n25193_not ; n25194
g22759 and n25192_not n25194 ; n25195
g22760 nor n25187 n25191 ; n25196
g22761 and n25195_not n25196 ; n25197
g22762 and pi0788 n25197_not ; n25198
g22763 and pi0618 n25135 ; n25199
g22764 nor n17168 n25125 ; n25200
g22765 and pi0625 n25200 ; n25201
g22766 and n25146 n25200_not ; n25202
g22767 nor n25201 n25202 ; n25203
g22768 and n25130 n25203_not ; n25204
g22769 nor pi0608 n25129 ; n25205
g22770 and n25204_not n25205 ; n25206
g22771 and pi1153 n25146 ; n25207
g22772 and n25201_not n25207 ; n25208
g22773 and pi0608 n25131_not ; n25209
g22774 and n25208_not n25209 ; n25210
g22775 nor n25206 n25210 ; n25211
g22776 and pi0778 n25211_not ; n25212
g22777 nor pi0778 n25202 ; n25213
g22778 nor n25212 n25213 ; n25214
g22779 nor pi0609 n25214 ; n25215
g22780 and pi0609 n25134_not ; n25216
g22781 nor pi1155 n25216 ; n25217
g22782 and n25215_not n25217 ; n25218
g22783 nor pi0660 n25151 ; n25219
g22784 and n25218_not n25219 ; n25220
g22785 and pi0609 n25214_not ; n25221
g22786 nor pi0609 n25134 ; n25222
g22787 and pi1155 n25222_not ; n25223
g22788 and n25221_not n25223 ; n25224
g22789 and pi0660 n25153_not ; n25225
g22790 and n25224_not n25225 ; n25226
g22791 nor n25220 n25226 ; n25227
g22792 and pi0785 n25227_not ; n25228
g22793 nor pi0785 n25214 ; n25229
g22794 nor n25228 n25229 ; n25230
g22795 nor pi0618 n25230 ; n25231
g22796 nor pi1154 n25199 ; n25232
g22797 and n25231_not n25232 ; n25233
g22798 nor pi0627 n25159 ; n25234
g22799 and n25233_not n25234 ; n25235
g22800 and pi0618_not n25135 ; n25236
g22801 and pi0618 n25230_not ; n25237
g22802 and pi1154 n25236_not ; n25238
g22803 and n25237_not n25238 ; n25239
g22804 and pi0627 n25161_not ; n25240
g22805 and n25239_not n25240 ; n25241
g22806 nor n25235 n25241 ; n25242
g22807 and pi0781 n25242_not ; n25243
g22808 nor pi0781 n25230 ; n25244
g22809 nor n25243 n25244 ; n25245
g22810 and pi0789_not n25245 ; n25246
g22811 nor pi0619 n25245 ; n25247
g22812 and pi0619 n25136 ; n25248
g22813 nor pi1159 n25248 ; n25249
g22814 and n25247_not n25249 ; n25250
g22815 nor pi0648 n25167 ; n25251
g22816 and n25250_not n25251 ; n25252
g22817 and pi0619 n25245_not ; n25253
g22818 and pi0619_not n25136 ; n25254
g22819 and pi1159 n25254_not ; n25255
g22820 and n25253_not n25255 ; n25256
g22821 and pi0648 n25169_not ; n25257
g22822 and n25256_not n25257 ; n25258
g22823 and pi0789 n25252_not ; n25259
g22824 and n25258_not n25259 ; n25260
g22825 and n17970 n25246_not ; n25261
g22826 and n25260_not n25261 ; n25262
g22827 nor n25198 n25262 ; n25263
g22828 nor n20364 n25263 ; n25264
g22829 and n17854 n25175_not ; n25265
g22830 and n20851 n25138 ; n25266
g22831 nor n25265 n25266 ; n25267
g22832 nor pi0629 n25267 ; n25268
g22833 and n20855 n25138 ; n25269
g22834 and n17853 n25175_not ; n25270
g22835 nor n25269 n25270 ; n25271
g22836 and pi0629 n25271_not ; n25272
g22837 nor n25268 n25272 ; n25273
g22838 and pi0792 n25273_not ; n25274
g22839 nor n20206 n25274 ; n25275
g22840 and n25264_not n25275 ; n25276
g22841 nor n25186 n25276 ; n25277
g22842 and pi0790_not n25277 ; n25278
g22843 nor pi0787 n25139 ; n25279
g22844 and pi1157 n25182_not ; n25280
g22845 nor n25143 n25280 ; n25281
g22846 and pi0787 n25281_not ; n25282
g22847 nor n25279 n25282 ; n25283
g22848 and pi0644_not n25283 ; n25284
g22849 and pi0644 n25277 ; n25285
g22850 and pi0715 n25284_not ; n25286
g22851 and n25285_not n25286 ; n25287
g22852 nor n17804 n25178 ; n25288
g22853 and n17804 n25123 ; n25289
g22854 nor n25288 n25289 ; n25290
g22855 and pi0644 n25290_not ; n25291
g22856 and pi0644_not n25123 ; n25292
g22857 nor pi0715 n25292 ; n25293
g22858 and n25291_not n25293 ; n25294
g22859 and pi1160 n25294_not ; n25295
g22860 and n25287_not n25295 ; n25296
g22861 nor pi0644 n25290 ; n25297
g22862 and pi0644 n25123 ; n25298
g22863 and pi0715 n25298_not ; n25299
g22864 and n25297_not n25299 ; n25300
g22865 and pi0644 n25283 ; n25301
g22866 and pi0644_not n25277 ; n25302
g22867 nor pi0715 n25301 ; n25303
g22868 and n25302_not n25303 ; n25304
g22869 nor pi1160 n25300 ; n25305
g22870 and n25304_not n25305 ; n25306
g22871 nor n25296 n25306 ; n25307
g22872 and pi0790 n25307_not ; n25308
g22873 and pi0832 n25278_not ; n25309
g22874 and n25308_not n25309 ; n25310
g22875 and pi0178_not po1038 ; n25311
g22876 nor pi0178 n17059 ; n25312
g22877 and n16635 n25312_not ; n25313
g22878 and pi0688_not n2571 ; n25314
g22879 and n25312 n25314_not ; n25315
g22880 nor pi0178 n16641 ; n25316
g22881 and n16647 n25316_not ; n25317
g22882 and pi0178 n18076_not ; n25318
g22883 nor pi0038 n25318 ; n25319
g22884 and n2571 n25319_not ; n25320
g22885 and pi0178_not n18072 ; n25321
g22886 nor n25320 n25321 ; n25322
g22887 nor pi0688 n25317 ; n25323
g22888 and n25322_not n25323 ; n25324
g22889 nor n25315 n25324 ; n25325
g22890 and pi0778_not n25325 ; n25326
g22891 and pi0625_not n25312 ; n25327
g22892 and pi0625 n25325_not ; n25328
g22893 and pi1153 n25327_not ; n25329
g22894 and n25328_not n25329 ; n25330
g22895 and pi0625 n25312 ; n25331
g22896 nor pi0625 n25325 ; n25332
g22897 nor pi1153 n25331 ; n25333
g22898 and n25332_not n25333 ; n25334
g22899 nor n25330 n25334 ; n25335
g22900 and pi0778 n25335_not ; n25336
g22901 nor n25326 n25336 ; n25337
g22902 nor n17075 n25337 ; n25338
g22903 and n17075 n25312_not ; n25339
g22904 nor n25338 n25339 ; n25340
g22905 and n16639_not n25340 ; n25341
g22906 and n16639 n25312 ; n25342
g22907 nor n25341 n25342 ; n25343
g22908 and n16635_not n25343 ; n25344
g22909 nor n25313 n25344 ; n25345
g22910 and n16631_not n25345 ; n25346
g22911 and n16631 n25312 ; n25347
g22912 nor n25346 n25347 ; n25348
g22913 and pi0792_not n25348 ; n25349
g22914 and pi0628 n25348_not ; n25350
g22915 and pi0628_not n25312 ; n25351
g22916 and pi1156 n25351_not ; n25352
g22917 and n25350_not n25352 ; n25353
g22918 and pi0628 n25312 ; n25354
g22919 nor pi0628 n25348 ; n25355
g22920 nor pi1156 n25354 ; n25356
g22921 and n25355_not n25356 ; n25357
g22922 nor n25353 n25357 ; n25358
g22923 and pi0792 n25358_not ; n25359
g22924 nor n25349 n25359 ; n25360
g22925 nor pi0647 n25360 ; n25361
g22926 and pi0647 n25312_not ; n25362
g22927 nor n25361 n25362 ; n25363
g22928 and pi1157_not n25363 ; n25364
g22929 and pi0647 n25360_not ; n25365
g22930 nor pi0647 n25312 ; n25366
g22931 nor n25365 n25366 ; n25367
g22932 and pi1157 n25367 ; n25368
g22933 nor n25364 n25368 ; n25369
g22934 and pi0787 n25369_not ; n25370
g22935 and pi0787_not n25360 ; n25371
g22936 nor n25370 n25371 ; n25372
g22937 nor pi0644 n25372 ; n25373
g22938 and pi0715 n25373_not ; n25374
g22939 and pi0178 n2571_not ; n25375
g22940 and pi0760_not n17280 ; n25376
g22941 nor n25316 n25376 ; n25377
g22942 and pi0038 n25377_not ; n25378
g22943 and pi0178_not n17221 ; n25379
g22944 and pi0178 n17275_not ; n25380
g22945 nor pi0760 n25380 ; n25381
g22946 and n25379_not n25381 ; n25382
g22947 and pi0178_not pi0760 ; n25383
g22948 and n17048_not n25383 ; n25384
g22949 nor n25382 n25384 ; n25385
g22950 nor pi0038 n25385 ; n25386
g22951 nor n25378 n25386 ; n25387
g22952 and n2571 n25387 ; n25388
g22953 nor n25375 n25388 ; n25389
g22954 nor n17117 n25389 ; n25390
g22955 and n17117 n25312_not ; n25391
g22956 nor n25390 n25391 ; n25392
g22957 nor pi0785 n25392 ; n25393
g22958 nor n17291 n25312 ; n25394
g22959 and pi0609 n25390 ; n25395
g22960 nor n25394 n25395 ; n25396
g22961 and pi1155 n25396_not ; n25397
g22962 nor n17296 n25312 ; n25398
g22963 and pi0609_not n25390 ; n25399
g22964 nor n25398 n25399 ; n25400
g22965 nor pi1155 n25400 ; n25401
g22966 nor n25397 n25401 ; n25402
g22967 and pi0785 n25402_not ; n25403
g22968 nor n25393 n25403 ; n25404
g22969 nor pi0781 n25404 ; n25405
g22970 and pi0618_not n25312 ; n25406
g22971 and pi0618 n25404 ; n25407
g22972 and pi1154 n25406_not ; n25408
g22973 and n25407_not n25408 ; n25409
g22974 and pi0618_not n25404 ; n25410
g22975 and pi0618 n25312 ; n25411
g22976 nor pi1154 n25411 ; n25412
g22977 and n25410_not n25412 ; n25413
g22978 nor n25409 n25413 ; n25414
g22979 and pi0781 n25414_not ; n25415
g22980 nor n25405 n25415 ; n25416
g22981 nor pi0789 n25416 ; n25417
g22982 and pi0619_not n25312 ; n25418
g22983 and pi0619 n25416 ; n25419
g22984 and pi1159 n25418_not ; n25420
g22985 and n25419_not n25420 ; n25421
g22986 and pi0619_not n25416 ; n25422
g22987 and pi0619 n25312 ; n25423
g22988 nor pi1159 n25423 ; n25424
g22989 and n25422_not n25424 ; n25425
g22990 nor n25421 n25425 ; n25426
g22991 and pi0789 n25426_not ; n25427
g22992 nor n25417 n25427 ; n25428
g22993 and n17969_not n25428 ; n25429
g22994 and n17969 n25312 ; n25430
g22995 nor n25429 n25430 ; n25431
g22996 nor n17779 n25431 ; n25432
g22997 and n17779 n25312 ; n25433
g22998 nor n25432 n25433 ; n25434
g22999 nor n17804 n25434 ; n25435
g23000 and n17804 n25312 ; n25436
g23001 nor n25435 n25436 ; n25437
g23002 and pi0644 n25437_not ; n25438
g23003 and pi0644_not n25312 ; n25439
g23004 nor pi0715 n25439 ; n25440
g23005 and n25438_not n25440 ; n25441
g23006 and pi1160 n25441_not ; n25442
g23007 and n25374_not n25442 ; n25443
g23008 and pi0644 n25372_not ; n25444
g23009 nor pi0715 n25444 ; n25445
g23010 nor pi0644 n25437 ; n25446
g23011 and pi0644 n25312 ; n25447
g23012 and pi0715 n25447_not ; n25448
g23013 and n25446_not n25448 ; n25449
g23014 nor pi1160 n25449 ; n25450
g23015 and n25445_not n25450 ; n25451
g23016 nor n25443 n25451 ; n25452
g23017 and pi0790 n25452_not ; n25453
g23018 and pi0629_not n25353 ; n25454
g23019 and n20570_not n25431 ; n25455
g23020 and pi0629 n25357 ; n25456
g23021 nor n25454 n25456 ; n25457
g23022 and n25455_not n25457 ; n25458
g23023 and pi0792 n25458_not ; n25459
g23024 and pi0609 n25337 ; n25460
g23025 and pi0178 n17625_not ; n25461
g23026 nor pi0178 n17612 ; n25462
g23027 and pi0760 n25461_not ; n25463
g23028 and n25462_not n25463 ; n25464
g23029 and pi0178_not n17629 ; n25465
g23030 and pi0178 n17631 ; n25466
g23031 nor pi0760 n25466 ; n25467
g23032 and n25465_not n25467 ; n25468
g23033 nor n25464 n25468 ; n25469
g23034 nor pi0039 n25469 ; n25470
g23035 and pi0178 n17605 ; n25471
g23036 nor pi0178 n17546 ; n25472
g23037 nor pi0760 n25472 ; n25473
g23038 and n25471_not n25473 ; n25474
g23039 and pi0178_not n17404 ; n25475
g23040 and pi0178 n17485 ; n25476
g23041 and pi0760 n25476_not ; n25477
g23042 and n25475_not n25477 ; n25478
g23043 and pi0039 n25474_not ; n25479
g23044 and n25478_not n25479 ; n25480
g23045 nor pi0038 n25470 ; n25481
g23046 and n25480_not n25481 ; n25482
g23047 nor pi0760 n17490 ; n25483
g23048 and n19471 n25483_not ; n25484
g23049 nor pi0178 n25484 ; n25485
g23050 nor n17469 n25145 ; n25486
g23051 and pi0178 n25486_not ; n25487
g23052 and n6284 n25487 ; n25488
g23053 and pi0038 n25488_not ; n25489
g23054 and n25485_not n25489 ; n25490
g23055 nor pi0688 n25490 ; n25491
g23056 and n25482_not n25491 ; n25492
g23057 and pi0688 n25387_not ; n25493
g23058 and n2571 n25492_not ; n25494
g23059 and n25493_not n25494 ; n25495
g23060 nor n25375 n25495 ; n25496
g23061 and pi0625_not n25496 ; n25497
g23062 and pi0625 n25389 ; n25498
g23063 nor pi1153 n25498 ; n25499
g23064 and n25497_not n25499 ; n25500
g23065 nor pi0608 n25330 ; n25501
g23066 and n25500_not n25501 ; n25502
g23067 and pi0625_not n25389 ; n25503
g23068 and pi0625 n25496 ; n25504
g23069 and pi1153 n25503_not ; n25505
g23070 and n25504_not n25505 ; n25506
g23071 and pi0608 n25334_not ; n25507
g23072 and n25506_not n25507 ; n25508
g23073 nor n25502 n25508 ; n25509
g23074 and pi0778 n25509_not ; n25510
g23075 and pi0778_not n25496 ; n25511
g23076 nor n25510 n25511 ; n25512
g23077 nor pi0609 n25512 ; n25513
g23078 nor pi1155 n25460 ; n25514
g23079 and n25513_not n25514 ; n25515
g23080 nor pi0660 n25397 ; n25516
g23081 and n25515_not n25516 ; n25517
g23082 and pi0609_not n25337 ; n25518
g23083 and pi0609 n25512_not ; n25519
g23084 and pi1155 n25518_not ; n25520
g23085 and n25519_not n25520 ; n25521
g23086 and pi0660 n25401_not ; n25522
g23087 and n25521_not n25522 ; n25523
g23088 nor n25517 n25523 ; n25524
g23089 and pi0785 n25524_not ; n25525
g23090 nor pi0785 n25512 ; n25526
g23091 nor n25525 n25526 ; n25527
g23092 nor pi0618 n25527 ; n25528
g23093 and pi0618 n25340 ; n25529
g23094 nor pi1154 n25529 ; n25530
g23095 and n25528_not n25530 ; n25531
g23096 nor pi0627 n25409 ; n25532
g23097 and n25531_not n25532 ; n25533
g23098 and pi0618_not n25340 ; n25534
g23099 and pi0618 n25527_not ; n25535
g23100 and pi1154 n25534_not ; n25536
g23101 and n25535_not n25536 ; n25537
g23102 and pi0627 n25413_not ; n25538
g23103 and n25537_not n25538 ; n25539
g23104 nor n25533 n25539 ; n25540
g23105 and pi0781 n25540_not ; n25541
g23106 nor pi0781 n25527 ; n25542
g23107 nor n25541 n25542 ; n25543
g23108 and pi0789_not n25543 ; n25544
g23109 and pi0619 n25343_not ; n25545
g23110 nor pi0619 n25543 ; n25546
g23111 nor pi1159 n25545 ; n25547
g23112 and n25546_not n25547 ; n25548
g23113 nor pi0648 n25421 ; n25549
g23114 and n25548_not n25549 ; n25550
g23115 nor pi0619 n25343 ; n25551
g23116 and pi0619 n25543_not ; n25552
g23117 and pi1159 n25551_not ; n25553
g23118 and n25552_not n25553 ; n25554
g23119 and pi0648 n25425_not ; n25555
g23120 and n25554_not n25555 ; n25556
g23121 and pi0789 n25550_not ; n25557
g23122 and n25556_not n25557 ; n25558
g23123 and n17970 n25544_not ; n25559
g23124 and n25558_not n25559 ; n25560
g23125 and n17871 n25345 ; n25561
g23126 nor pi0626 n25428 ; n25562
g23127 and pi0626 n25312_not ; n25563
g23128 and n16629 n25563_not ; n25564
g23129 and n25562_not n25564 ; n25565
g23130 and pi0626 n25428_not ; n25566
g23131 nor pi0626 n25312 ; n25567
g23132 and n16628 n25567_not ; n25568
g23133 and n25566_not n25568 ; n25569
g23134 nor n25561 n25565 ; n25570
g23135 and n25569_not n25570 ; n25571
g23136 and pi0788 n25571_not ; n25572
g23137 nor n20364 n25572 ; n25573
g23138 and n25560_not n25573 ; n25574
g23139 nor n25459 n25574 ; n25575
g23140 nor n20206 n25575 ; n25576
g23141 and n17802 n25363_not ; n25577
g23142 and n20559_not n25434 ; n25578
g23143 and n17801 n25367_not ; n25579
g23144 nor n25577 n25579 ; n25580
g23145 and n25578_not n25580 ; n25581
g23146 and pi0787 n25581_not ; n25582
g23147 and pi0644_not n25450 ; n25583
g23148 and pi0644 n25442 ; n25584
g23149 and pi0790 n25583_not ; n25585
g23150 and n25584_not n25585 ; n25586
g23151 nor n25576 n25582 ; n25587
g23152 and n25586_not n25587 ; n25588
g23153 nor n25453 n25588 ; n25589
g23154 nor po1038 n25589 ; n25590
g23155 nor pi0832 n25311 ; n25591
g23156 and n25590_not n25591 ; n25592
g23157 nor n25310 n25592 ; po0335
g23158 nor pi0179 n17059 ; n25594
g23159 and n16635 n25594_not ; n25595
g23160 and pi0724_not n2571 ; n25596
g23161 and n25594 n25596_not ; n25597
g23162 nor pi0179 n16641 ; n25598
g23163 and n16647 n25598_not ; n25599
g23164 and pi0179_not n18072 ; n25600
g23165 and pi0179 n18076_not ; n25601
g23166 nor pi0038 n25601 ; n25602
g23167 and n2571 n25602_not ; n25603
g23168 nor n25600 n25603 ; n25604
g23169 nor pi0724 n25599 ; n25605
g23170 and n25604_not n25605 ; n25606
g23171 nor n25597 n25606 ; n25607
g23172 and pi0778_not n25607 ; n25608
g23173 and pi0625_not n25594 ; n25609
g23174 and pi0625 n25607_not ; n25610
g23175 and pi1153 n25609_not ; n25611
g23176 and n25610_not n25611 ; n25612
g23177 and pi0625 n25594 ; n25613
g23178 nor pi0625 n25607 ; n25614
g23179 nor pi1153 n25613 ; n25615
g23180 and n25614_not n25615 ; n25616
g23181 nor n25612 n25616 ; n25617
g23182 and pi0778 n25617_not ; n25618
g23183 nor n25608 n25618 ; n25619
g23184 nor n17075 n25619 ; n25620
g23185 and n17075 n25594_not ; n25621
g23186 nor n25620 n25621 ; n25622
g23187 and n16639_not n25622 ; n25623
g23188 and n16639 n25594 ; n25624
g23189 nor n25623 n25624 ; n25625
g23190 and n16635_not n25625 ; n25626
g23191 nor n25595 n25626 ; n25627
g23192 and n16631_not n25627 ; n25628
g23193 and n16631 n25594 ; n25629
g23194 nor n25628 n25629 ; n25630
g23195 and pi0792_not n25630 ; n25631
g23196 and pi0628_not n25594 ; n25632
g23197 and pi0628 n25630_not ; n25633
g23198 and pi1156 n25632_not ; n25634
g23199 and n25633_not n25634 ; n25635
g23200 and pi0628 n25594 ; n25636
g23201 nor pi0628 n25630 ; n25637
g23202 nor pi1156 n25636 ; n25638
g23203 and n25637_not n25638 ; n25639
g23204 nor n25635 n25639 ; n25640
g23205 and pi0792 n25640_not ; n25641
g23206 nor n25631 n25641 ; n25642
g23207 nor pi0787 n25642 ; n25643
g23208 and pi0647_not n25594 ; n25644
g23209 and pi0647 n25642 ; n25645
g23210 and pi1157 n25644_not ; n25646
g23211 and n25645_not n25646 ; n25647
g23212 and pi0647_not n25642 ; n25648
g23213 and pi0647 n25594 ; n25649
g23214 nor pi1157 n25649 ; n25650
g23215 and n25648_not n25650 ; n25651
g23216 nor n25647 n25651 ; n25652
g23217 and pi0787 n25652_not ; n25653
g23218 nor n25643 n25653 ; n25654
g23219 and pi0644_not n25654 ; n25655
g23220 and pi0618_not n25594 ; n25656
g23221 and pi0179 n2571_not ; n25657
g23222 nor pi0741 n24447 ; n25658
g23223 and pi0179 n25658_not ; n25659
g23224 nor pi0179 pi0741 ; n25660
g23225 and n19433_not n25660 ; n25661
g23226 and n19439 n25661 ; n25662
g23227 nor n25659 n25662 ; n25663
g23228 and n21674_not n25663 ; n25664
g23229 and n2571 n25664_not ; n25665
g23230 nor n25657 n25665 ; n25666
g23231 nor n17117 n25666 ; n25667
g23232 and n17117 n25594_not ; n25668
g23233 nor n25667 n25668 ; n25669
g23234 nor pi0785 n25669 ; n25670
g23235 nor n17291 n25594 ; n25671
g23236 and pi0609 n25667 ; n25672
g23237 nor n25671 n25672 ; n25673
g23238 and pi1155 n25673_not ; n25674
g23239 nor n17296 n25594 ; n25675
g23240 and pi0609_not n25667 ; n25676
g23241 nor n25675 n25676 ; n25677
g23242 nor pi1155 n25677 ; n25678
g23243 nor n25674 n25678 ; n25679
g23244 and pi0785 n25679_not ; n25680
g23245 nor n25670 n25680 ; n25681
g23246 and pi0618 n25681 ; n25682
g23247 and pi1154 n25656_not ; n25683
g23248 and n25682_not n25683 ; n25684
g23249 and n18176 n25598_not ; n25685
g23250 and pi0179_not n17404 ; n25686
g23251 and pi0179 n17485 ; n25687
g23252 and pi0039 n25687_not ; n25688
g23253 and n25686_not n25688 ; n25689
g23254 and pi0179_not n17612 ; n25690
g23255 and pi0179 n17625 ; n25691
g23256 nor pi0039 n25690 ; n25692
g23257 and n25691_not n25692 ; n25693
g23258 nor n25689 n25693 ; n25694
g23259 nor pi0038 n25694 ; n25695
g23260 nor n25685 n25695 ; n25696
g23261 and pi0741 n25696_not ; n25697
g23262 nor pi0179 n19488 ; n25698
g23263 and pi0179 n19496 ; n25699
g23264 nor pi0741 n25698 ; n25700
g23265 and n25699_not n25700 ; n25701
g23266 nor pi0724 n25701 ; n25702
g23267 and n25697_not n25702 ; n25703
g23268 and pi0724 n25664 ; n25704
g23269 and n2571 n25704_not ; n25705
g23270 and n25703_not n25705 ; n25706
g23271 nor n25657 n25706 ; n25707
g23272 and pi0625_not n25707 ; n25708
g23273 and pi0625 n25666 ; n25709
g23274 nor pi1153 n25709 ; n25710
g23275 and n25708_not n25710 ; n25711
g23276 nor pi0608 n25612 ; n25712
g23277 and n25711_not n25712 ; n25713
g23278 and pi0625_not n25666 ; n25714
g23279 and pi0625 n25707 ; n25715
g23280 and pi1153 n25714_not ; n25716
g23281 and n25715_not n25716 ; n25717
g23282 and pi0608 n25616_not ; n25718
g23283 and n25717_not n25718 ; n25719
g23284 nor n25713 n25719 ; n25720
g23285 and pi0778 n25720_not ; n25721
g23286 and pi0778_not n25707 ; n25722
g23287 nor n25721 n25722 ; n25723
g23288 nor pi0609 n25723 ; n25724
g23289 and pi0609 n25619 ; n25725
g23290 nor pi1155 n25725 ; n25726
g23291 and n25724_not n25726 ; n25727
g23292 nor pi0660 n25674 ; n25728
g23293 and n25727_not n25728 ; n25729
g23294 and pi0609_not n25619 ; n25730
g23295 and pi0609 n25723_not ; n25731
g23296 and pi1155 n25730_not ; n25732
g23297 and n25731_not n25732 ; n25733
g23298 and pi0660 n25678_not ; n25734
g23299 and n25733_not n25734 ; n25735
g23300 nor n25729 n25735 ; n25736
g23301 and pi0785 n25736_not ; n25737
g23302 nor pi0785 n25723 ; n25738
g23303 nor n25737 n25738 ; n25739
g23304 nor pi0618 n25739 ; n25740
g23305 and pi0618 n25622 ; n25741
g23306 nor pi1154 n25741 ; n25742
g23307 and n25740_not n25742 ; n25743
g23308 nor pi0627 n25684 ; n25744
g23309 and n25743_not n25744 ; n25745
g23310 and pi0618_not n25681 ; n25746
g23311 and pi0618 n25594 ; n25747
g23312 nor pi1154 n25747 ; n25748
g23313 and n25746_not n25748 ; n25749
g23314 and pi0618_not n25622 ; n25750
g23315 and pi0618 n25739_not ; n25751
g23316 and pi1154 n25750_not ; n25752
g23317 and n25751_not n25752 ; n25753
g23318 and pi0627 n25749_not ; n25754
g23319 and n25753_not n25754 ; n25755
g23320 nor n25745 n25755 ; n25756
g23321 and pi0781 n25756_not ; n25757
g23322 nor pi0781 n25739 ; n25758
g23323 nor n25757 n25758 ; n25759
g23324 nor pi0619 n25759 ; n25760
g23325 and pi0619 n25625_not ; n25761
g23326 nor pi1159 n25761 ; n25762
g23327 and n25760_not n25762 ; n25763
g23328 and pi0619_not n25594 ; n25764
g23329 nor pi0781 n25681 ; n25765
g23330 nor n25684 n25749 ; n25766
g23331 and pi0781 n25766_not ; n25767
g23332 nor n25765 n25767 ; n25768
g23333 and pi0619 n25768 ; n25769
g23334 and pi1159 n25764_not ; n25770
g23335 and n25769_not n25770 ; n25771
g23336 nor pi0648 n25771 ; n25772
g23337 and n25763_not n25772 ; n25773
g23338 and pi0619 n25759_not ; n25774
g23339 nor pi0619 n25625 ; n25775
g23340 and pi1159 n25775_not ; n25776
g23341 and n25774_not n25776 ; n25777
g23342 and pi0619_not n25768 ; n25778
g23343 and pi0619 n25594 ; n25779
g23344 nor pi1159 n25779 ; n25780
g23345 and n25778_not n25780 ; n25781
g23346 and pi0648 n25781_not ; n25782
g23347 and n25777_not n25782 ; n25783
g23348 nor n25773 n25783 ; n25784
g23349 and pi0789 n25784_not ; n25785
g23350 nor pi0789 n25759 ; n25786
g23351 nor n25785 n25786 ; n25787
g23352 and pi0788_not n25787 ; n25788
g23353 and pi0626_not n25787 ; n25789
g23354 and pi0626 n25627_not ; n25790
g23355 nor pi0641 n25790 ; n25791
g23356 and n25789_not n25791 ; n25792
g23357 nor pi0789 n25768 ; n25793
g23358 nor n25771 n25781 ; n25794
g23359 and pi0789 n25794_not ; n25795
g23360 nor n25793 n25795 ; n25796
g23361 nor pi0626 n25796 ; n25797
g23362 and pi0626 n25594_not ; n25798
g23363 and pi0641 n25798_not ; n25799
g23364 and n25797_not n25799 ; n25800
g23365 nor pi1158 n25800 ; n25801
g23366 and n25792_not n25801 ; n25802
g23367 and pi0626 n25787 ; n25803
g23368 nor pi0626 n25627 ; n25804
g23369 and pi0641 n25804_not ; n25805
g23370 and n25803_not n25805 ; n25806
g23371 and pi0626 n25796_not ; n25807
g23372 nor pi0626 n25594 ; n25808
g23373 nor pi0641 n25808 ; n25809
g23374 and n25807_not n25809 ; n25810
g23375 and pi1158 n25810_not ; n25811
g23376 and n25806_not n25811 ; n25812
g23377 nor n25802 n25812 ; n25813
g23378 and pi0788 n25813_not ; n25814
g23379 nor n25788 n25814 ; n25815
g23380 and pi0628_not n25815 ; n25816
g23381 and n17969_not n25796 ; n25817
g23382 and n17969 n25594 ; n25818
g23383 nor n25817 n25818 ; n25819
g23384 and pi0628 n25819_not ; n25820
g23385 nor pi1156 n25820 ; n25821
g23386 and n25816_not n25821 ; n25822
g23387 nor pi0629 n25635 ; n25823
g23388 and n25822_not n25823 ; n25824
g23389 and pi0628 n25815 ; n25825
g23390 nor pi0628 n25819 ; n25826
g23391 and pi1156 n25826_not ; n25827
g23392 and n25825_not n25827 ; n25828
g23393 and pi0629 n25639_not ; n25829
g23394 and n25828_not n25829 ; n25830
g23395 nor n25824 n25830 ; n25831
g23396 and pi0792 n25831_not ; n25832
g23397 and pi0792_not n25815 ; n25833
g23398 nor n25832 n25833 ; n25834
g23399 nor pi0647 n25834 ; n25835
g23400 nor n17779 n25819 ; n25836
g23401 and n17779 n25594 ; n25837
g23402 nor n25836 n25837 ; n25838
g23403 and pi0647 n25838_not ; n25839
g23404 nor pi1157 n25839 ; n25840
g23405 and n25835_not n25840 ; n25841
g23406 nor pi0630 n25647 ; n25842
g23407 and n25841_not n25842 ; n25843
g23408 and pi0647 n25834_not ; n25844
g23409 nor pi0647 n25838 ; n25845
g23410 and pi1157 n25845_not ; n25846
g23411 and n25844_not n25846 ; n25847
g23412 and pi0630 n25651_not ; n25848
g23413 and n25847_not n25848 ; n25849
g23414 nor n25843 n25849 ; n25850
g23415 and pi0787 n25850_not ; n25851
g23416 nor pi0787 n25834 ; n25852
g23417 nor n25851 n25852 ; n25853
g23418 and pi0644 n25853_not ; n25854
g23419 and pi0715 n25655_not ; n25855
g23420 and n25854_not n25855 ; n25856
g23421 and n17804 n25594_not ; n25857
g23422 and n17804_not n25838 ; n25858
g23423 nor n25857 n25858 ; n25859
g23424 and pi0644 n25859 ; n25860
g23425 and pi0644_not n25594 ; n25861
g23426 nor pi0715 n25861 ; n25862
g23427 and n25860_not n25862 ; n25863
g23428 and pi1160 n25863_not ; n25864
g23429 and n25856_not n25864 ; n25865
g23430 nor pi0644 n25853 ; n25866
g23431 and pi0644 n25654 ; n25867
g23432 nor pi0715 n25867 ; n25868
g23433 and n25866_not n25868 ; n25869
g23434 and pi0644_not n25859 ; n25870
g23435 and pi0644 n25594 ; n25871
g23436 and pi0715 n25871_not ; n25872
g23437 and n25870_not n25872 ; n25873
g23438 nor pi1160 n25873 ; n25874
g23439 and n25869_not n25874 ; n25875
g23440 and pi0790 n25865_not ; n25876
g23441 and n25875_not n25876 ; n25877
g23442 and pi0790_not n25853 ; n25878
g23443 nor po1038 n25878 ; n25879
g23444 and n25877_not n25879 ; n25880
g23445 and pi0179_not po1038 ; n25881
g23446 nor pi0832 n25881 ; n25882
g23447 and n25880_not n25882 ; n25883
g23448 nor pi0179 n2926 ; n25884
g23449 and pi0724_not n16645 ; n25885
g23450 nor n25884 n25885 ; n25886
g23451 and pi0778_not n25886 ; n25887
g23452 and pi0625_not n25885 ; n25888
g23453 nor n25886 n25888 ; n25889
g23454 and pi1153 n25889_not ; n25890
g23455 nor pi1153 n25884 ; n25891
g23456 and n25888_not n25891 ; n25892
g23457 nor n25890 n25892 ; n25893
g23458 and pi0778 n25893_not ; n25894
g23459 nor n25887 n25894 ; n25895
g23460 and n17845_not n25895 ; n25896
g23461 and n17847_not n25896 ; n25897
g23462 and n17849_not n25897 ; n25898
g23463 and n17851_not n25898 ; n25899
g23464 and n17857_not n25899 ; n25900
g23465 and pi0647_not n25900 ; n25901
g23466 and pi0647 n25884 ; n25902
g23467 nor pi1157 n25902 ; n25903
g23468 and n25901_not n25903 ; n25904
g23469 and pi0630 n25904 ; n25905
g23470 and pi0741_not n17244 ; n25906
g23471 nor n25884 n25906 ; n25907
g23472 nor n17874 n25907 ; n25908
g23473 nor pi0785 n25908 ; n25909
g23474 nor n17879 n25907 ; n25910
g23475 and pi1155 n25910_not ; n25911
g23476 and n17882_not n25908 ; n25912
g23477 nor pi1155 n25912 ; n25913
g23478 nor n25911 n25913 ; n25914
g23479 and pi0785 n25914_not ; n25915
g23480 nor n25909 n25915 ; n25916
g23481 nor pi0781 n25916 ; n25917
g23482 and n17889_not n25916 ; n25918
g23483 and pi1154 n25918_not ; n25919
g23484 and n17892_not n25916 ; n25920
g23485 nor pi1154 n25920 ; n25921
g23486 nor n25919 n25921 ; n25922
g23487 and pi0781 n25922_not ; n25923
g23488 nor n25917 n25923 ; n25924
g23489 nor pi0789 n25924 ; n25925
g23490 and pi0619_not n25884 ; n25926
g23491 and pi0619 n25924 ; n25927
g23492 and pi1159 n25926_not ; n25928
g23493 and n25927_not n25928 ; n25929
g23494 and pi0619_not n25924 ; n25930
g23495 and pi0619 n25884 ; n25931
g23496 nor pi1159 n25931 ; n25932
g23497 and n25930_not n25932 ; n25933
g23498 nor n25929 n25933 ; n25934
g23499 and pi0789 n25934_not ; n25935
g23500 nor n25925 n25935 ; n25936
g23501 and n17969_not n25936 ; n25937
g23502 and n17969 n25884 ; n25938
g23503 nor n25937 n25938 ; n25939
g23504 nor n17779 n25939 ; n25940
g23505 and n17779 n25884 ; n25941
g23506 nor n25940 n25941 ; n25942
g23507 and n20559_not n25942 ; n25943
g23508 and pi0647 n25900_not ; n25944
g23509 nor pi0647 n25884 ; n25945
g23510 nor n25944 n25945 ; n25946
g23511 and n17801 n25946_not ; n25947
g23512 nor n25905 n25947 ; n25948
g23513 and n25943_not n25948 ; n25949
g23514 and pi0787 n25949_not ; n25950
g23515 and n17871 n25898 ; n25951
g23516 nor pi0626 n25936 ; n25952
g23517 and pi0626 n25884_not ; n25953
g23518 and n16629 n25953_not ; n25954
g23519 and n25952_not n25954 ; n25955
g23520 and pi0626 n25936_not ; n25956
g23521 nor pi0626 n25884 ; n25957
g23522 and n16628 n25957_not ; n25958
g23523 and n25956_not n25958 ; n25959
g23524 nor n25951 n25955 ; n25960
g23525 and n25959_not n25960 ; n25961
g23526 and pi0788 n25961_not ; n25962
g23527 and pi0618 n25896 ; n25963
g23528 and pi0609 n25895 ; n25964
g23529 nor n17168 n25886 ; n25965
g23530 and pi0625 n25965 ; n25966
g23531 and n25907 n25965_not ; n25967
g23532 nor n25966 n25967 ; n25968
g23533 and n25891 n25968_not ; n25969
g23534 nor pi0608 n25890 ; n25970
g23535 and n25969_not n25970 ; n25971
g23536 and pi1153 n25907 ; n25972
g23537 and n25966_not n25972 ; n25973
g23538 and pi0608 n25892_not ; n25974
g23539 and n25973_not n25974 ; n25975
g23540 nor n25971 n25975 ; n25976
g23541 and pi0778 n25976_not ; n25977
g23542 nor pi0778 n25967 ; n25978
g23543 nor n25977 n25978 ; n25979
g23544 nor pi0609 n25979 ; n25980
g23545 nor pi1155 n25964 ; n25981
g23546 and n25980_not n25981 ; n25982
g23547 nor pi0660 n25911 ; n25983
g23548 and n25982_not n25983 ; n25984
g23549 and pi0609_not n25895 ; n25985
g23550 and pi0609 n25979_not ; n25986
g23551 and pi1155 n25985_not ; n25987
g23552 and n25986_not n25987 ; n25988
g23553 and pi0660 n25913_not ; n25989
g23554 and n25988_not n25989 ; n25990
g23555 nor n25984 n25990 ; n25991
g23556 and pi0785 n25991_not ; n25992
g23557 nor pi0785 n25979 ; n25993
g23558 nor n25992 n25993 ; n25994
g23559 nor pi0618 n25994 ; n25995
g23560 nor pi1154 n25963 ; n25996
g23561 and n25995_not n25996 ; n25997
g23562 nor pi0627 n25919 ; n25998
g23563 and n25997_not n25998 ; n25999
g23564 and pi0618_not n25896 ; n26000
g23565 and pi0618 n25994_not ; n26001
g23566 and pi1154 n26000_not ; n26002
g23567 and n26001_not n26002 ; n26003
g23568 and pi0627 n25921_not ; n26004
g23569 and n26003_not n26004 ; n26005
g23570 nor n25999 n26005 ; n26006
g23571 and pi0781 n26006_not ; n26007
g23572 nor pi0781 n25994 ; n26008
g23573 nor n26007 n26008 ; n26009
g23574 and pi0789_not n26009 ; n26010
g23575 nor pi0619 n26009 ; n26011
g23576 and pi0619 n25897 ; n26012
g23577 nor pi1159 n26012 ; n26013
g23578 and n26011_not n26013 ; n26014
g23579 nor pi0648 n25929 ; n26015
g23580 and n26014_not n26015 ; n26016
g23581 and pi0619 n26009_not ; n26017
g23582 and pi0619_not n25897 ; n26018
g23583 and pi1159 n26018_not ; n26019
g23584 and n26017_not n26019 ; n26020
g23585 and pi0648 n25933_not ; n26021
g23586 and n26020_not n26021 ; n26022
g23587 and pi0789 n26016_not ; n26023
g23588 and n26022_not n26023 ; n26024
g23589 and n17970 n26010_not ; n26025
g23590 and n26024_not n26025 ; n26026
g23591 nor n25962 n26026 ; n26027
g23592 nor n20364 n26027 ; n26028
g23593 and n17854 n25939_not ; n26029
g23594 and n20851 n25899 ; n26030
g23595 nor n26029 n26030 ; n26031
g23596 nor pi0629 n26031 ; n26032
g23597 and n20855 n25899 ; n26033
g23598 and n17853 n25939_not ; n26034
g23599 nor n26033 n26034 ; n26035
g23600 and pi0629 n26035_not ; n26036
g23601 nor n26032 n26036 ; n26037
g23602 and pi0792 n26037_not ; n26038
g23603 nor n20206 n26038 ; n26039
g23604 and n26028_not n26039 ; n26040
g23605 nor n25950 n26040 ; n26041
g23606 and pi0790_not n26041 ; n26042
g23607 nor pi0787 n25900 ; n26043
g23608 and pi1157 n25946_not ; n26044
g23609 nor n25904 n26044 ; n26045
g23610 and pi0787 n26045_not ; n26046
g23611 nor n26043 n26046 ; n26047
g23612 and pi0644_not n26047 ; n26048
g23613 and pi0644 n26041 ; n26049
g23614 and pi0715 n26048_not ; n26050
g23615 and n26049_not n26050 ; n26051
g23616 nor n17804 n25942 ; n26052
g23617 and n17804 n25884 ; n26053
g23618 nor n26052 n26053 ; n26054
g23619 and pi0644 n26054_not ; n26055
g23620 and pi0644_not n25884 ; n26056
g23621 nor pi0715 n26056 ; n26057
g23622 and n26055_not n26057 ; n26058
g23623 and pi1160 n26058_not ; n26059
g23624 and n26051_not n26059 ; n26060
g23625 nor pi0644 n26054 ; n26061
g23626 and pi0644 n25884 ; n26062
g23627 and pi0715 n26062_not ; n26063
g23628 and n26061_not n26063 ; n26064
g23629 and pi0644 n26047 ; n26065
g23630 and pi0644_not n26041 ; n26066
g23631 nor pi0715 n26065 ; n26067
g23632 and n26066_not n26067 ; n26068
g23633 nor pi1160 n26064 ; n26069
g23634 and n26068_not n26069 ; n26070
g23635 nor n26060 n26070 ; n26071
g23636 and pi0790 n26071_not ; n26072
g23637 and pi0832 n26042_not ; n26073
g23638 and n26072_not n26073 ; n26074
g23639 nor n25883 n26074 ; po0336
g23640 nor pi0180 n2926 ; n26076
g23641 and pi0702_not n16645 ; n26077
g23642 nor n26076 n26077 ; n26078
g23643 nor pi0778 n26078 ; n26079
g23644 and pi0625_not n26077 ; n26080
g23645 nor n26078 n26080 ; n26081
g23646 and pi1153 n26081_not ; n26082
g23647 nor pi1153 n26076 ; n26083
g23648 and n26080_not n26083 ; n26084
g23649 and pi0778 n26084_not ; n26085
g23650 and n26082_not n26085 ; n26086
g23651 nor n26079 n26086 ; n26087
g23652 nor n17845 n26087 ; n26088
g23653 and n17847_not n26088 ; n26089
g23654 and n17849_not n26089 ; n26090
g23655 and n17851_not n26090 ; n26091
g23656 and n17857_not n26091 ; n26092
g23657 and pi0647_not n26092 ; n26093
g23658 and pi0647 n26076 ; n26094
g23659 nor pi1157 n26094 ; n26095
g23660 and n26093_not n26095 ; n26096
g23661 and pi0630 n26096 ; n26097
g23662 and pi0753_not n17244 ; n26098
g23663 nor n26076 n26098 ; n26099
g23664 nor n17874 n26099 ; n26100
g23665 nor pi0785 n26100 ; n26101
g23666 and n17296 n26098 ; n26102
g23667 and n26100 n26102_not ; n26103
g23668 and pi1155 n26103_not ; n26104
g23669 nor pi1155 n26076 ; n26105
g23670 and n26102_not n26105 ; n26106
g23671 nor n26104 n26106 ; n26107
g23672 and pi0785 n26107_not ; n26108
g23673 nor n26101 n26108 ; n26109
g23674 nor pi0781 n26109 ; n26110
g23675 and n17889_not n26109 ; n26111
g23676 and pi1154 n26111_not ; n26112
g23677 and n17892_not n26109 ; n26113
g23678 nor pi1154 n26113 ; n26114
g23679 nor n26112 n26114 ; n26115
g23680 and pi0781 n26115_not ; n26116
g23681 nor n26110 n26116 ; n26117
g23682 nor pi0789 n26117 ; n26118
g23683 and n23078_not n26117 ; n26119
g23684 and pi1159 n26119_not ; n26120
g23685 and n23081_not n26117 ; n26121
g23686 nor pi1159 n26121 ; n26122
g23687 nor n26120 n26122 ; n26123
g23688 and pi0789 n26123_not ; n26124
g23689 nor n26118 n26124 ; n26125
g23690 and n17969_not n26125 ; n26126
g23691 and n17969 n26076 ; n26127
g23692 nor n26126 n26127 ; n26128
g23693 nor n17779 n26128 ; n26129
g23694 and n17779 n26076 ; n26130
g23695 nor n26129 n26130 ; n26131
g23696 and n20559_not n26131 ; n26132
g23697 and pi0647 n26092_not ; n26133
g23698 nor pi0647 n26076 ; n26134
g23699 nor n26133 n26134 ; n26135
g23700 and n17801 n26135_not ; n26136
g23701 nor n26097 n26136 ; n26137
g23702 and n26132_not n26137 ; n26138
g23703 and pi0787 n26138_not ; n26139
g23704 and n17871 n26090 ; n26140
g23705 nor pi0626 n26125 ; n26141
g23706 and pi0626 n26076_not ; n26142
g23707 and n16629 n26142_not ; n26143
g23708 and n26141_not n26143 ; n26144
g23709 and pi0626 n26125_not ; n26145
g23710 nor pi0626 n26076 ; n26146
g23711 and n16628 n26146_not ; n26147
g23712 and n26145_not n26147 ; n26148
g23713 nor n26140 n26144 ; n26149
g23714 and n26148_not n26149 ; n26150
g23715 and pi0788 n26150_not ; n26151
g23716 and pi0618 n26088 ; n26152
g23717 nor n17168 n26078 ; n26153
g23718 and pi0625 n26153 ; n26154
g23719 and n26099 n26153_not ; n26155
g23720 nor n26154 n26155 ; n26156
g23721 and n26083 n26156_not ; n26157
g23722 nor pi0608 n26082 ; n26158
g23723 and n26157_not n26158 ; n26159
g23724 and pi1153 n26099 ; n26160
g23725 and n26154_not n26160 ; n26161
g23726 and pi0608 n26084_not ; n26162
g23727 and n26161_not n26162 ; n26163
g23728 nor n26159 n26163 ; n26164
g23729 and pi0778 n26164_not ; n26165
g23730 nor pi0778 n26155 ; n26166
g23731 nor n26165 n26166 ; n26167
g23732 nor pi0609 n26167 ; n26168
g23733 and pi0609 n26087_not ; n26169
g23734 nor pi1155 n26169 ; n26170
g23735 and n26168_not n26170 ; n26171
g23736 nor pi0660 n26104 ; n26172
g23737 and n26171_not n26172 ; n26173
g23738 and pi0609 n26167_not ; n26174
g23739 nor pi0609 n26087 ; n26175
g23740 and pi1155 n26175_not ; n26176
g23741 and n26174_not n26176 ; n26177
g23742 and pi0660 n26106_not ; n26178
g23743 and n26177_not n26178 ; n26179
g23744 nor n26173 n26179 ; n26180
g23745 and pi0785 n26180_not ; n26181
g23746 nor pi0785 n26167 ; n26182
g23747 nor n26181 n26182 ; n26183
g23748 nor pi0618 n26183 ; n26184
g23749 nor pi1154 n26152 ; n26185
g23750 and n26184_not n26185 ; n26186
g23751 nor pi0627 n26112 ; n26187
g23752 and n26186_not n26187 ; n26188
g23753 and pi0618_not n26088 ; n26189
g23754 and pi0618 n26183_not ; n26190
g23755 and pi1154 n26189_not ; n26191
g23756 and n26190_not n26191 ; n26192
g23757 and pi0627 n26114_not ; n26193
g23758 and n26192_not n26193 ; n26194
g23759 nor n26188 n26194 ; n26195
g23760 and pi0781 n26195_not ; n26196
g23761 nor pi0781 n26183 ; n26197
g23762 nor n26196 n26197 ; n26198
g23763 and pi0789_not n26198 ; n26199
g23764 nor pi0619 n26198 ; n26200
g23765 and pi0619 n26089 ; n26201
g23766 nor pi1159 n26201 ; n26202
g23767 and n26200_not n26202 ; n26203
g23768 nor pi0648 n26120 ; n26204
g23769 and n26203_not n26204 ; n26205
g23770 and pi0619 n26198_not ; n26206
g23771 and pi0619_not n26089 ; n26207
g23772 and pi1159 n26207_not ; n26208
g23773 and n26206_not n26208 ; n26209
g23774 and pi0648 n26122_not ; n26210
g23775 and n26209_not n26210 ; n26211
g23776 and pi0789 n26205_not ; n26212
g23777 and n26211_not n26212 ; n26213
g23778 and n17970 n26199_not ; n26214
g23779 and n26213_not n26214 ; n26215
g23780 nor n26151 n26215 ; n26216
g23781 nor n20364 n26216 ; n26217
g23782 and n17854 n26128_not ; n26218
g23783 and n20851 n26091 ; n26219
g23784 nor n26218 n26219 ; n26220
g23785 nor pi0629 n26220 ; n26221
g23786 and n20855 n26091 ; n26222
g23787 and n17853 n26128_not ; n26223
g23788 nor n26222 n26223 ; n26224
g23789 and pi0629 n26224_not ; n26225
g23790 nor n26221 n26225 ; n26226
g23791 and pi0792 n26226_not ; n26227
g23792 nor n20206 n26227 ; n26228
g23793 and n26217_not n26228 ; n26229
g23794 nor n26139 n26229 ; n26230
g23795 and pi0790_not n26230 ; n26231
g23796 nor pi0787 n26092 ; n26232
g23797 and pi1157 n26135_not ; n26233
g23798 nor n26096 n26233 ; n26234
g23799 and pi0787 n26234_not ; n26235
g23800 nor n26232 n26235 ; n26236
g23801 and pi0644_not n26236 ; n26237
g23802 and pi0644 n26230 ; n26238
g23803 and pi0715 n26237_not ; n26239
g23804 and n26238_not n26239 ; n26240
g23805 nor n17804 n26131 ; n26241
g23806 and n17804 n26076 ; n26242
g23807 nor n26241 n26242 ; n26243
g23808 and pi0644 n26243_not ; n26244
g23809 and pi0644_not n26076 ; n26245
g23810 nor pi0715 n26245 ; n26246
g23811 and n26244_not n26246 ; n26247
g23812 and pi1160 n26247_not ; n26248
g23813 and n26240_not n26248 ; n26249
g23814 nor pi0644 n26243 ; n26250
g23815 and pi0644 n26076 ; n26251
g23816 and pi0715 n26251_not ; n26252
g23817 and n26250_not n26252 ; n26253
g23818 and pi0644 n26236 ; n26254
g23819 and pi0644_not n26230 ; n26255
g23820 nor pi0715 n26254 ; n26256
g23821 and n26255_not n26256 ; n26257
g23822 nor pi1160 n26253 ; n26258
g23823 and n26257_not n26258 ; n26259
g23824 nor n26249 n26259 ; n26260
g23825 and pi0790 n26260_not ; n26261
g23826 and pi0832 n26231_not ; n26262
g23827 and n26261_not n26262 ; n26263
g23828 and pi0180_not po1038 ; n26264
g23829 nor pi0180 n17059 ; n26265
g23830 and n16635 n26265_not ; n26266
g23831 and pi0702_not n2571 ; n26267
g23832 and n26265 n26267_not ; n26268
g23833 nor pi0180 n16641 ; n26269
g23834 and n16647 n26269_not ; n26270
g23835 and pi0180 n18076_not ; n26271
g23836 nor pi0038 n26271 ; n26272
g23837 and n2571 n26272_not ; n26273
g23838 and pi0180_not n18072 ; n26274
g23839 nor n26273 n26274 ; n26275
g23840 nor pi0702 n26270 ; n26276
g23841 and n26275_not n26276 ; n26277
g23842 nor n26268 n26277 ; n26278
g23843 and pi0778_not n26278 ; n26279
g23844 and pi0625_not n26265 ; n26280
g23845 and pi0625 n26278_not ; n26281
g23846 and pi1153 n26280_not ; n26282
g23847 and n26281_not n26282 ; n26283
g23848 and pi0625 n26265 ; n26284
g23849 nor pi0625 n26278 ; n26285
g23850 nor pi1153 n26284 ; n26286
g23851 and n26285_not n26286 ; n26287
g23852 nor n26283 n26287 ; n26288
g23853 and pi0778 n26288_not ; n26289
g23854 nor n26279 n26289 ; n26290
g23855 nor n17075 n26290 ; n26291
g23856 and n17075 n26265_not ; n26292
g23857 nor n26291 n26292 ; n26293
g23858 and n16639_not n26293 ; n26294
g23859 and n16639 n26265 ; n26295
g23860 nor n26294 n26295 ; n26296
g23861 and n16635_not n26296 ; n26297
g23862 nor n26266 n26297 ; n26298
g23863 and n16631_not n26298 ; n26299
g23864 and n16631 n26265 ; n26300
g23865 nor n26299 n26300 ; n26301
g23866 and pi0792_not n26301 ; n26302
g23867 and pi0628 n26301_not ; n26303
g23868 and pi0628_not n26265 ; n26304
g23869 and pi1156 n26304_not ; n26305
g23870 and n26303_not n26305 ; n26306
g23871 and pi0628 n26265 ; n26307
g23872 nor pi0628 n26301 ; n26308
g23873 nor pi1156 n26307 ; n26309
g23874 and n26308_not n26309 ; n26310
g23875 nor n26306 n26310 ; n26311
g23876 and pi0792 n26311_not ; n26312
g23877 nor n26302 n26312 ; n26313
g23878 nor pi0647 n26313 ; n26314
g23879 and pi0647 n26265_not ; n26315
g23880 nor n26314 n26315 ; n26316
g23881 and pi1157_not n26316 ; n26317
g23882 and pi0647 n26313_not ; n26318
g23883 nor pi0647 n26265 ; n26319
g23884 nor n26318 n26319 ; n26320
g23885 and pi1157 n26320 ; n26321
g23886 nor n26317 n26321 ; n26322
g23887 and pi0787 n26322_not ; n26323
g23888 and pi0787_not n26313 ; n26324
g23889 nor n26323 n26324 ; n26325
g23890 nor pi0644 n26325 ; n26326
g23891 and pi0715 n26326_not ; n26327
g23892 and pi0180 n2571_not ; n26328
g23893 and pi0180 pi0753 ; n26329
g23894 and pi0753 n17046 ; n26330
g23895 and pi0180 n17273 ; n26331
g23896 nor n26330 n26331 ; n26332
g23897 and pi0039 n26332_not ; n26333
g23898 and pi0180 n17233_not ; n26334
g23899 nor n21756 n26334 ; n26335
g23900 nor pi0039 n26335 ; n26336
g23901 nor pi0180 pi0753 ; n26337
g23902 and n17221 n26337 ; n26338
g23903 nor n26329 n26336 ; n26339
g23904 and n26338_not n26339 ; n26340
g23905 and n26333_not n26340 ; n26341
g23906 nor pi0038 n26341 ; n26342
g23907 and pi0753_not n17280 ; n26343
g23908 and pi0038 n26269_not ; n26344
g23909 and n26343_not n26344 ; n26345
g23910 nor n26342 n26345 ; n26346
g23911 and n2571 n26346_not ; n26347
g23912 nor n26328 n26347 ; n26348
g23913 nor n17117 n26348 ; n26349
g23914 and n17117 n26265_not ; n26350
g23915 nor n26349 n26350 ; n26351
g23916 nor pi0785 n26351 ; n26352
g23917 nor n17291 n26265 ; n26353
g23918 and pi0609 n26349 ; n26354
g23919 nor n26353 n26354 ; n26355
g23920 and pi1155 n26355_not ; n26356
g23921 nor n17296 n26265 ; n26357
g23922 and pi0609_not n26349 ; n26358
g23923 nor n26357 n26358 ; n26359
g23924 nor pi1155 n26359 ; n26360
g23925 nor n26356 n26360 ; n26361
g23926 and pi0785 n26361_not ; n26362
g23927 nor n26352 n26362 ; n26363
g23928 nor pi0781 n26363 ; n26364
g23929 and pi0618_not n26265 ; n26365
g23930 and pi0618 n26363 ; n26366
g23931 and pi1154 n26365_not ; n26367
g23932 and n26366_not n26367 ; n26368
g23933 and pi0618_not n26363 ; n26369
g23934 and pi0618 n26265 ; n26370
g23935 nor pi1154 n26370 ; n26371
g23936 and n26369_not n26371 ; n26372
g23937 nor n26368 n26372 ; n26373
g23938 and pi0781 n26373_not ; n26374
g23939 nor n26364 n26374 ; n26375
g23940 nor pi0789 n26375 ; n26376
g23941 and pi0619_not n26265 ; n26377
g23942 and pi0619 n26375 ; n26378
g23943 and pi1159 n26377_not ; n26379
g23944 and n26378_not n26379 ; n26380
g23945 and pi0619_not n26375 ; n26381
g23946 and pi0619 n26265 ; n26382
g23947 nor pi1159 n26382 ; n26383
g23948 and n26381_not n26383 ; n26384
g23949 nor n26380 n26384 ; n26385
g23950 and pi0789 n26385_not ; n26386
g23951 nor n26376 n26386 ; n26387
g23952 and n17969_not n26387 ; n26388
g23953 and n17969 n26265 ; n26389
g23954 nor n26388 n26389 ; n26390
g23955 nor n17779 n26390 ; n26391
g23956 and n17779 n26265 ; n26392
g23957 nor n26391 n26392 ; n26393
g23958 nor n17804 n26393 ; n26394
g23959 and n17804 n26265 ; n26395
g23960 nor n26394 n26395 ; n26396
g23961 and pi0644 n26396_not ; n26397
g23962 and pi0644_not n26265 ; n26398
g23963 nor pi0715 n26398 ; n26399
g23964 and n26397_not n26399 ; n26400
g23965 and pi1160 n26400_not ; n26401
g23966 and n26327_not n26401 ; n26402
g23967 and pi0644 n26325_not ; n26403
g23968 nor pi0715 n26403 ; n26404
g23969 nor pi0644 n26396 ; n26405
g23970 and pi0644 n26265 ; n26406
g23971 and pi0715 n26406_not ; n26407
g23972 and n26405_not n26407 ; n26408
g23973 nor pi1160 n26408 ; n26409
g23974 and n26404_not n26409 ; n26410
g23975 nor n26402 n26410 ; n26411
g23976 and pi0790 n26411_not ; n26412
g23977 and pi0629_not n26306 ; n26413
g23978 and n20570_not n26390 ; n26414
g23979 and pi0629 n26310 ; n26415
g23980 nor n26413 n26415 ; n26416
g23981 and n26414_not n26416 ; n26417
g23982 and pi0792 n26417_not ; n26418
g23983 and pi0609 n26290 ; n26419
g23984 and pi0180 n17625_not ; n26420
g23985 nor pi0180 n17612 ; n26421
g23986 and pi0753 n26420_not ; n26422
g23987 and n26421_not n26422 ; n26423
g23988 and pi0180_not n17629 ; n26424
g23989 and pi0180 n17631 ; n26425
g23990 nor pi0753 n26425 ; n26426
g23991 and n26424_not n26426 ; n26427
g23992 nor n26423 n26427 ; n26428
g23993 nor pi0039 n26428 ; n26429
g23994 and pi0180 n17605 ; n26430
g23995 nor pi0180 n17546 ; n26431
g23996 nor pi0753 n26431 ; n26432
g23997 and n26430_not n26432 ; n26433
g23998 and pi0180_not n17404 ; n26434
g23999 and pi0180 n17485 ; n26435
g24000 and pi0753 n26435_not ; n26436
g24001 and n26434_not n26436 ; n26437
g24002 and pi0039 n26433_not ; n26438
g24003 and n26437_not n26438 ; n26439
g24004 nor pi0038 n26429 ; n26440
g24005 and n26439_not n26440 ; n26441
g24006 nor n17469 n26098 ; n26442
g24007 and pi0180 n26442_not ; n26443
g24008 and n6284 n26443 ; n26444
g24009 nor pi0753 n17490 ; n26445
g24010 and n19471 n26445_not ; n26446
g24011 nor pi0180 n26446 ; n26447
g24012 and pi0038 n26444_not ; n26448
g24013 and n26447_not n26448 ; n26449
g24014 nor pi0702 n26449 ; n26450
g24015 and n26441_not n26450 ; n26451
g24016 and pi0702 n26346 ; n26452
g24017 and n2571 n26451_not ; n26453
g24018 and n26452_not n26453 ; n26454
g24019 nor n26328 n26454 ; n26455
g24020 and pi0625_not n26455 ; n26456
g24021 and pi0625 n26348 ; n26457
g24022 nor pi1153 n26457 ; n26458
g24023 and n26456_not n26458 ; n26459
g24024 nor pi0608 n26283 ; n26460
g24025 and n26459_not n26460 ; n26461
g24026 and pi0625_not n26348 ; n26462
g24027 and pi0625 n26455 ; n26463
g24028 and pi1153 n26462_not ; n26464
g24029 and n26463_not n26464 ; n26465
g24030 and pi0608 n26287_not ; n26466
g24031 and n26465_not n26466 ; n26467
g24032 nor n26461 n26467 ; n26468
g24033 and pi0778 n26468_not ; n26469
g24034 and pi0778_not n26455 ; n26470
g24035 nor n26469 n26470 ; n26471
g24036 nor pi0609 n26471 ; n26472
g24037 nor pi1155 n26419 ; n26473
g24038 and n26472_not n26473 ; n26474
g24039 nor pi0660 n26356 ; n26475
g24040 and n26474_not n26475 ; n26476
g24041 and pi0609_not n26290 ; n26477
g24042 and pi0609 n26471_not ; n26478
g24043 and pi1155 n26477_not ; n26479
g24044 and n26478_not n26479 ; n26480
g24045 and pi0660 n26360_not ; n26481
g24046 and n26480_not n26481 ; n26482
g24047 nor n26476 n26482 ; n26483
g24048 and pi0785 n26483_not ; n26484
g24049 nor pi0785 n26471 ; n26485
g24050 nor n26484 n26485 ; n26486
g24051 nor pi0618 n26486 ; n26487
g24052 and pi0618 n26293 ; n26488
g24053 nor pi1154 n26488 ; n26489
g24054 and n26487_not n26489 ; n26490
g24055 nor pi0627 n26368 ; n26491
g24056 and n26490_not n26491 ; n26492
g24057 and pi0618_not n26293 ; n26493
g24058 and pi0618 n26486_not ; n26494
g24059 and pi1154 n26493_not ; n26495
g24060 and n26494_not n26495 ; n26496
g24061 and pi0627 n26372_not ; n26497
g24062 and n26496_not n26497 ; n26498
g24063 nor n26492 n26498 ; n26499
g24064 and pi0781 n26499_not ; n26500
g24065 nor pi0781 n26486 ; n26501
g24066 nor n26500 n26501 ; n26502
g24067 and pi0789_not n26502 ; n26503
g24068 and pi0619 n26296_not ; n26504
g24069 nor pi0619 n26502 ; n26505
g24070 nor pi1159 n26504 ; n26506
g24071 and n26505_not n26506 ; n26507
g24072 nor pi0648 n26380 ; n26508
g24073 and n26507_not n26508 ; n26509
g24074 nor pi0619 n26296 ; n26510
g24075 and pi0619 n26502_not ; n26511
g24076 and pi1159 n26510_not ; n26512
g24077 and n26511_not n26512 ; n26513
g24078 and pi0648 n26384_not ; n26514
g24079 and n26513_not n26514 ; n26515
g24080 and pi0789 n26509_not ; n26516
g24081 and n26515_not n26516 ; n26517
g24082 and n17970 n26503_not ; n26518
g24083 and n26517_not n26518 ; n26519
g24084 and n17871 n26298 ; n26520
g24085 nor pi0626 n26387 ; n26521
g24086 and pi0626 n26265_not ; n26522
g24087 and n16629 n26522_not ; n26523
g24088 and n26521_not n26523 ; n26524
g24089 and pi0626 n26387_not ; n26525
g24090 nor pi0626 n26265 ; n26526
g24091 and n16628 n26526_not ; n26527
g24092 and n26525_not n26527 ; n26528
g24093 nor n26520 n26524 ; n26529
g24094 and n26528_not n26529 ; n26530
g24095 and pi0788 n26530_not ; n26531
g24096 nor n20364 n26531 ; n26532
g24097 and n26519_not n26532 ; n26533
g24098 nor n26418 n26533 ; n26534
g24099 nor n20206 n26534 ; n26535
g24100 and n17802 n26316_not ; n26536
g24101 and n20559_not n26393 ; n26537
g24102 and n17801 n26320_not ; n26538
g24103 nor n26536 n26538 ; n26539
g24104 and n26537_not n26539 ; n26540
g24105 and pi0787 n26540_not ; n26541
g24106 and pi0644_not n26409 ; n26542
g24107 and pi0644 n26401 ; n26543
g24108 and pi0790 n26542_not ; n26544
g24109 and n26543_not n26544 ; n26545
g24110 nor n26535 n26541 ; n26546
g24111 and n26545_not n26546 ; n26547
g24112 nor n26412 n26547 ; n26548
g24113 nor po1038 n26548 ; n26549
g24114 nor pi0832 n26264 ; n26550
g24115 and n26549_not n26550 ; n26551
g24116 nor n26263 n26551 ; po0337
g24117 nor pi0181 n2926 ; n26553
g24118 and pi0709_not n16645 ; n26554
g24119 nor n26553 n26554 ; n26555
g24120 nor pi0778 n26555 ; n26556
g24121 and pi0625_not n26554 ; n26557
g24122 nor n26555 n26557 ; n26558
g24123 and pi1153 n26558_not ; n26559
g24124 nor pi1153 n26553 ; n26560
g24125 and n26557_not n26560 ; n26561
g24126 and pi0778 n26561_not ; n26562
g24127 and n26559_not n26562 ; n26563
g24128 nor n26556 n26563 ; n26564
g24129 nor n17845 n26564 ; n26565
g24130 and n17847_not n26565 ; n26566
g24131 and n17849_not n26566 ; n26567
g24132 and n17851_not n26567 ; n26568
g24133 and n17857_not n26568 ; n26569
g24134 and pi0647_not n26569 ; n26570
g24135 and pi0647 n26553 ; n26571
g24136 nor pi1157 n26571 ; n26572
g24137 and n26570_not n26572 ; n26573
g24138 and pi0630 n26573 ; n26574
g24139 and pi0754_not n17244 ; n26575
g24140 nor n26553 n26575 ; n26576
g24141 nor n17874 n26576 ; n26577
g24142 nor pi0785 n26577 ; n26578
g24143 and n17296 n26575 ; n26579
g24144 and n26577 n26579_not ; n26580
g24145 and pi1155 n26580_not ; n26581
g24146 nor pi1155 n26553 ; n26582
g24147 and n26579_not n26582 ; n26583
g24148 nor n26581 n26583 ; n26584
g24149 and pi0785 n26584_not ; n26585
g24150 nor n26578 n26585 ; n26586
g24151 nor pi0781 n26586 ; n26587
g24152 and n17889_not n26586 ; n26588
g24153 and pi1154 n26588_not ; n26589
g24154 and n17892_not n26586 ; n26590
g24155 nor pi1154 n26590 ; n26591
g24156 nor n26589 n26591 ; n26592
g24157 and pi0781 n26592_not ; n26593
g24158 nor n26587 n26593 ; n26594
g24159 nor pi0789 n26594 ; n26595
g24160 and n23078_not n26594 ; n26596
g24161 and pi1159 n26596_not ; n26597
g24162 and n23081_not n26594 ; n26598
g24163 nor pi1159 n26598 ; n26599
g24164 nor n26597 n26599 ; n26600
g24165 and pi0789 n26600_not ; n26601
g24166 nor n26595 n26601 ; n26602
g24167 and n17969_not n26602 ; n26603
g24168 and n17969 n26553 ; n26604
g24169 nor n26603 n26604 ; n26605
g24170 nor n17779 n26605 ; n26606
g24171 and n17779 n26553 ; n26607
g24172 nor n26606 n26607 ; n26608
g24173 and n20559_not n26608 ; n26609
g24174 and pi0647 n26569_not ; n26610
g24175 nor pi0647 n26553 ; n26611
g24176 nor n26610 n26611 ; n26612
g24177 and n17801 n26612_not ; n26613
g24178 nor n26574 n26613 ; n26614
g24179 and n26609_not n26614 ; n26615
g24180 and pi0787 n26615_not ; n26616
g24181 and n17871 n26567 ; n26617
g24182 nor pi0626 n26602 ; n26618
g24183 and pi0626 n26553_not ; n26619
g24184 and n16629 n26619_not ; n26620
g24185 and n26618_not n26620 ; n26621
g24186 and pi0626 n26602_not ; n26622
g24187 nor pi0626 n26553 ; n26623
g24188 and n16628 n26623_not ; n26624
g24189 and n26622_not n26624 ; n26625
g24190 nor n26617 n26621 ; n26626
g24191 and n26625_not n26626 ; n26627
g24192 and pi0788 n26627_not ; n26628
g24193 and pi0618 n26565 ; n26629
g24194 nor n17168 n26555 ; n26630
g24195 and pi0625 n26630 ; n26631
g24196 and n26576 n26630_not ; n26632
g24197 nor n26631 n26632 ; n26633
g24198 and n26560 n26633_not ; n26634
g24199 nor pi0608 n26559 ; n26635
g24200 and n26634_not n26635 ; n26636
g24201 and pi1153 n26576 ; n26637
g24202 and n26631_not n26637 ; n26638
g24203 and pi0608 n26561_not ; n26639
g24204 and n26638_not n26639 ; n26640
g24205 nor n26636 n26640 ; n26641
g24206 and pi0778 n26641_not ; n26642
g24207 nor pi0778 n26632 ; n26643
g24208 nor n26642 n26643 ; n26644
g24209 nor pi0609 n26644 ; n26645
g24210 and pi0609 n26564_not ; n26646
g24211 nor pi1155 n26646 ; n26647
g24212 and n26645_not n26647 ; n26648
g24213 nor pi0660 n26581 ; n26649
g24214 and n26648_not n26649 ; n26650
g24215 and pi0609 n26644_not ; n26651
g24216 nor pi0609 n26564 ; n26652
g24217 and pi1155 n26652_not ; n26653
g24218 and n26651_not n26653 ; n26654
g24219 and pi0660 n26583_not ; n26655
g24220 and n26654_not n26655 ; n26656
g24221 nor n26650 n26656 ; n26657
g24222 and pi0785 n26657_not ; n26658
g24223 nor pi0785 n26644 ; n26659
g24224 nor n26658 n26659 ; n26660
g24225 nor pi0618 n26660 ; n26661
g24226 nor pi1154 n26629 ; n26662
g24227 and n26661_not n26662 ; n26663
g24228 nor pi0627 n26589 ; n26664
g24229 and n26663_not n26664 ; n26665
g24230 and pi0618_not n26565 ; n26666
g24231 and pi0618 n26660_not ; n26667
g24232 and pi1154 n26666_not ; n26668
g24233 and n26667_not n26668 ; n26669
g24234 and pi0627 n26591_not ; n26670
g24235 and n26669_not n26670 ; n26671
g24236 nor n26665 n26671 ; n26672
g24237 and pi0781 n26672_not ; n26673
g24238 nor pi0781 n26660 ; n26674
g24239 nor n26673 n26674 ; n26675
g24240 and pi0789_not n26675 ; n26676
g24241 nor pi0619 n26675 ; n26677
g24242 and pi0619 n26566 ; n26678
g24243 nor pi1159 n26678 ; n26679
g24244 and n26677_not n26679 ; n26680
g24245 nor pi0648 n26597 ; n26681
g24246 and n26680_not n26681 ; n26682
g24247 and pi0619 n26675_not ; n26683
g24248 and pi0619_not n26566 ; n26684
g24249 and pi1159 n26684_not ; n26685
g24250 and n26683_not n26685 ; n26686
g24251 and pi0648 n26599_not ; n26687
g24252 and n26686_not n26687 ; n26688
g24253 and pi0789 n26682_not ; n26689
g24254 and n26688_not n26689 ; n26690
g24255 and n17970 n26676_not ; n26691
g24256 and n26690_not n26691 ; n26692
g24257 nor n26628 n26692 ; n26693
g24258 nor n20364 n26693 ; n26694
g24259 and n17854 n26605_not ; n26695
g24260 and n20851 n26568 ; n26696
g24261 nor n26695 n26696 ; n26697
g24262 nor pi0629 n26697 ; n26698
g24263 and n20855 n26568 ; n26699
g24264 and n17853 n26605_not ; n26700
g24265 nor n26699 n26700 ; n26701
g24266 and pi0629 n26701_not ; n26702
g24267 nor n26698 n26702 ; n26703
g24268 and pi0792 n26703_not ; n26704
g24269 nor n20206 n26704 ; n26705
g24270 and n26694_not n26705 ; n26706
g24271 nor n26616 n26706 ; n26707
g24272 and pi0790_not n26707 ; n26708
g24273 nor pi0787 n26569 ; n26709
g24274 and pi1157 n26612_not ; n26710
g24275 nor n26573 n26710 ; n26711
g24276 and pi0787 n26711_not ; n26712
g24277 nor n26709 n26712 ; n26713
g24278 and pi0644_not n26713 ; n26714
g24279 and pi0644 n26707 ; n26715
g24280 and pi0715 n26714_not ; n26716
g24281 and n26715_not n26716 ; n26717
g24282 nor n17804 n26608 ; n26718
g24283 and n17804 n26553 ; n26719
g24284 nor n26718 n26719 ; n26720
g24285 and pi0644 n26720_not ; n26721
g24286 and pi0644_not n26553 ; n26722
g24287 nor pi0715 n26722 ; n26723
g24288 and n26721_not n26723 ; n26724
g24289 and pi1160 n26724_not ; n26725
g24290 and n26717_not n26725 ; n26726
g24291 nor pi0644 n26720 ; n26727
g24292 and pi0644 n26553 ; n26728
g24293 and pi0715 n26728_not ; n26729
g24294 and n26727_not n26729 ; n26730
g24295 and pi0644 n26713 ; n26731
g24296 and pi0644_not n26707 ; n26732
g24297 nor pi0715 n26731 ; n26733
g24298 and n26732_not n26733 ; n26734
g24299 nor pi1160 n26730 ; n26735
g24300 and n26734_not n26735 ; n26736
g24301 nor n26726 n26736 ; n26737
g24302 and pi0790 n26737_not ; n26738
g24303 and pi0832 n26708_not ; n26739
g24304 and n26738_not n26739 ; n26740
g24305 and pi0181_not po1038 ; n26741
g24306 nor pi0181 n17059 ; n26742
g24307 and n16635 n26742_not ; n26743
g24308 and pi0709_not n2571 ; n26744
g24309 and n26742 n26744_not ; n26745
g24310 nor pi0181 n16641 ; n26746
g24311 and n16647 n26746_not ; n26747
g24312 and pi0181 n18076_not ; n26748
g24313 nor pi0038 n26748 ; n26749
g24314 and n2571 n26749_not ; n26750
g24315 and pi0181_not n18072 ; n26751
g24316 nor n26750 n26751 ; n26752
g24317 nor pi0709 n26747 ; n26753
g24318 and n26752_not n26753 ; n26754
g24319 nor n26745 n26754 ; n26755
g24320 and pi0778_not n26755 ; n26756
g24321 and pi0625_not n26742 ; n26757
g24322 and pi0625 n26755_not ; n26758
g24323 and pi1153 n26757_not ; n26759
g24324 and n26758_not n26759 ; n26760
g24325 and pi0625 n26742 ; n26761
g24326 nor pi0625 n26755 ; n26762
g24327 nor pi1153 n26761 ; n26763
g24328 and n26762_not n26763 ; n26764
g24329 nor n26760 n26764 ; n26765
g24330 and pi0778 n26765_not ; n26766
g24331 nor n26756 n26766 ; n26767
g24332 nor n17075 n26767 ; n26768
g24333 and n17075 n26742_not ; n26769
g24334 nor n26768 n26769 ; n26770
g24335 and n16639_not n26770 ; n26771
g24336 and n16639 n26742 ; n26772
g24337 nor n26771 n26772 ; n26773
g24338 and n16635_not n26773 ; n26774
g24339 nor n26743 n26774 ; n26775
g24340 and n16631_not n26775 ; n26776
g24341 and n16631 n26742 ; n26777
g24342 nor n26776 n26777 ; n26778
g24343 and pi0792_not n26778 ; n26779
g24344 and pi0628 n26778_not ; n26780
g24345 and pi0628_not n26742 ; n26781
g24346 and pi1156 n26781_not ; n26782
g24347 and n26780_not n26782 ; n26783
g24348 and pi0628 n26742 ; n26784
g24349 nor pi0628 n26778 ; n26785
g24350 nor pi1156 n26784 ; n26786
g24351 and n26785_not n26786 ; n26787
g24352 nor n26783 n26787 ; n26788
g24353 and pi0792 n26788_not ; n26789
g24354 nor n26779 n26789 ; n26790
g24355 nor pi0647 n26790 ; n26791
g24356 and pi0647 n26742_not ; n26792
g24357 nor n26791 n26792 ; n26793
g24358 and pi1157_not n26793 ; n26794
g24359 and pi0647 n26790_not ; n26795
g24360 nor pi0647 n26742 ; n26796
g24361 nor n26795 n26796 ; n26797
g24362 and pi1157 n26797 ; n26798
g24363 nor n26794 n26798 ; n26799
g24364 and pi0787 n26799_not ; n26800
g24365 and pi0787_not n26790 ; n26801
g24366 nor n26800 n26801 ; n26802
g24367 nor pi0644 n26802 ; n26803
g24368 and pi0715 n26803_not ; n26804
g24369 and pi0181 n2571_not ; n26805
g24370 and pi0181 pi0754 ; n26806
g24371 and pi0754 n17046 ; n26807
g24372 and pi0181 n17273 ; n26808
g24373 nor n26807 n26808 ; n26809
g24374 and pi0039 n26809_not ; n26810
g24375 and pi0181 n17233_not ; n26811
g24376 nor n21812 n26811 ; n26812
g24377 nor pi0039 n26812 ; n26813
g24378 nor pi0181 pi0754 ; n26814
g24379 and n17221 n26814 ; n26815
g24380 nor n26806 n26813 ; n26816
g24381 and n26815_not n26816 ; n26817
g24382 and n26810_not n26817 ; n26818
g24383 nor pi0038 n26818 ; n26819
g24384 and pi0754_not n17280 ; n26820
g24385 and pi0038 n26746_not ; n26821
g24386 and n26820_not n26821 ; n26822
g24387 nor n26819 n26822 ; n26823
g24388 and n2571 n26823_not ; n26824
g24389 nor n26805 n26824 ; n26825
g24390 nor n17117 n26825 ; n26826
g24391 and n17117 n26742_not ; n26827
g24392 nor n26826 n26827 ; n26828
g24393 nor pi0785 n26828 ; n26829
g24394 nor n17291 n26742 ; n26830
g24395 and pi0609 n26826 ; n26831
g24396 nor n26830 n26831 ; n26832
g24397 and pi1155 n26832_not ; n26833
g24398 nor n17296 n26742 ; n26834
g24399 and pi0609_not n26826 ; n26835
g24400 nor n26834 n26835 ; n26836
g24401 nor pi1155 n26836 ; n26837
g24402 nor n26833 n26837 ; n26838
g24403 and pi0785 n26838_not ; n26839
g24404 nor n26829 n26839 ; n26840
g24405 nor pi0781 n26840 ; n26841
g24406 and pi0618_not n26742 ; n26842
g24407 and pi0618 n26840 ; n26843
g24408 and pi1154 n26842_not ; n26844
g24409 and n26843_not n26844 ; n26845
g24410 and pi0618_not n26840 ; n26846
g24411 and pi0618 n26742 ; n26847
g24412 nor pi1154 n26847 ; n26848
g24413 and n26846_not n26848 ; n26849
g24414 nor n26845 n26849 ; n26850
g24415 and pi0781 n26850_not ; n26851
g24416 nor n26841 n26851 ; n26852
g24417 nor pi0789 n26852 ; n26853
g24418 and pi0619_not n26742 ; n26854
g24419 and pi0619 n26852 ; n26855
g24420 and pi1159 n26854_not ; n26856
g24421 and n26855_not n26856 ; n26857
g24422 and pi0619_not n26852 ; n26858
g24423 and pi0619 n26742 ; n26859
g24424 nor pi1159 n26859 ; n26860
g24425 and n26858_not n26860 ; n26861
g24426 nor n26857 n26861 ; n26862
g24427 and pi0789 n26862_not ; n26863
g24428 nor n26853 n26863 ; n26864
g24429 and n17969_not n26864 ; n26865
g24430 and n17969 n26742 ; n26866
g24431 nor n26865 n26866 ; n26867
g24432 nor n17779 n26867 ; n26868
g24433 and n17779 n26742 ; n26869
g24434 nor n26868 n26869 ; n26870
g24435 nor n17804 n26870 ; n26871
g24436 and n17804 n26742 ; n26872
g24437 nor n26871 n26872 ; n26873
g24438 and pi0644 n26873_not ; n26874
g24439 and pi0644_not n26742 ; n26875
g24440 nor pi0715 n26875 ; n26876
g24441 and n26874_not n26876 ; n26877
g24442 and pi1160 n26877_not ; n26878
g24443 and n26804_not n26878 ; n26879
g24444 and pi0644 n26802_not ; n26880
g24445 nor pi0715 n26880 ; n26881
g24446 nor pi0644 n26873 ; n26882
g24447 and pi0644 n26742 ; n26883
g24448 and pi0715 n26883_not ; n26884
g24449 and n26882_not n26884 ; n26885
g24450 nor pi1160 n26885 ; n26886
g24451 and n26881_not n26886 ; n26887
g24452 nor n26879 n26887 ; n26888
g24453 and pi0790 n26888_not ; n26889
g24454 and pi0629_not n26783 ; n26890
g24455 and n20570_not n26867 ; n26891
g24456 and pi0629 n26787 ; n26892
g24457 nor n26890 n26892 ; n26893
g24458 and n26891_not n26893 ; n26894
g24459 and pi0792 n26894_not ; n26895
g24460 and pi0609 n26767 ; n26896
g24461 and pi0181 n17625_not ; n26897
g24462 nor pi0181 n17612 ; n26898
g24463 and pi0754 n26897_not ; n26899
g24464 and n26898_not n26899 ; n26900
g24465 and pi0181_not n17629 ; n26901
g24466 and pi0181 n17631 ; n26902
g24467 nor pi0754 n26902 ; n26903
g24468 and n26901_not n26903 ; n26904
g24469 nor n26900 n26904 ; n26905
g24470 nor pi0039 n26905 ; n26906
g24471 and pi0181 n17605 ; n26907
g24472 nor pi0181 n17546 ; n26908
g24473 nor pi0754 n26908 ; n26909
g24474 and n26907_not n26909 ; n26910
g24475 and pi0181_not n17404 ; n26911
g24476 and pi0181 n17485 ; n26912
g24477 and pi0754 n26912_not ; n26913
g24478 and n26911_not n26913 ; n26914
g24479 and pi0039 n26910_not ; n26915
g24480 and n26914_not n26915 ; n26916
g24481 nor pi0038 n26906 ; n26917
g24482 and n26916_not n26917 ; n26918
g24483 nor n17469 n26575 ; n26919
g24484 and pi0181 n26919_not ; n26920
g24485 and n6284 n26920 ; n26921
g24486 nor pi0754 n17490 ; n26922
g24487 and n19471 n26922_not ; n26923
g24488 nor pi0181 n26923 ; n26924
g24489 and pi0038 n26921_not ; n26925
g24490 and n26924_not n26925 ; n26926
g24491 nor pi0709 n26926 ; n26927
g24492 and n26918_not n26927 ; n26928
g24493 and pi0709 n26823 ; n26929
g24494 and n2571 n26928_not ; n26930
g24495 and n26929_not n26930 ; n26931
g24496 nor n26805 n26931 ; n26932
g24497 and pi0625_not n26932 ; n26933
g24498 and pi0625 n26825 ; n26934
g24499 nor pi1153 n26934 ; n26935
g24500 and n26933_not n26935 ; n26936
g24501 nor pi0608 n26760 ; n26937
g24502 and n26936_not n26937 ; n26938
g24503 and pi0625_not n26825 ; n26939
g24504 and pi0625 n26932 ; n26940
g24505 and pi1153 n26939_not ; n26941
g24506 and n26940_not n26941 ; n26942
g24507 and pi0608 n26764_not ; n26943
g24508 and n26942_not n26943 ; n26944
g24509 nor n26938 n26944 ; n26945
g24510 and pi0778 n26945_not ; n26946
g24511 and pi0778_not n26932 ; n26947
g24512 nor n26946 n26947 ; n26948
g24513 nor pi0609 n26948 ; n26949
g24514 nor pi1155 n26896 ; n26950
g24515 and n26949_not n26950 ; n26951
g24516 nor pi0660 n26833 ; n26952
g24517 and n26951_not n26952 ; n26953
g24518 and pi0609_not n26767 ; n26954
g24519 and pi0609 n26948_not ; n26955
g24520 and pi1155 n26954_not ; n26956
g24521 and n26955_not n26956 ; n26957
g24522 and pi0660 n26837_not ; n26958
g24523 and n26957_not n26958 ; n26959
g24524 nor n26953 n26959 ; n26960
g24525 and pi0785 n26960_not ; n26961
g24526 nor pi0785 n26948 ; n26962
g24527 nor n26961 n26962 ; n26963
g24528 nor pi0618 n26963 ; n26964
g24529 and pi0618 n26770 ; n26965
g24530 nor pi1154 n26965 ; n26966
g24531 and n26964_not n26966 ; n26967
g24532 nor pi0627 n26845 ; n26968
g24533 and n26967_not n26968 ; n26969
g24534 and pi0618_not n26770 ; n26970
g24535 and pi0618 n26963_not ; n26971
g24536 and pi1154 n26970_not ; n26972
g24537 and n26971_not n26972 ; n26973
g24538 and pi0627 n26849_not ; n26974
g24539 and n26973_not n26974 ; n26975
g24540 nor n26969 n26975 ; n26976
g24541 and pi0781 n26976_not ; n26977
g24542 nor pi0781 n26963 ; n26978
g24543 nor n26977 n26978 ; n26979
g24544 and pi0789_not n26979 ; n26980
g24545 and pi0619 n26773_not ; n26981
g24546 nor pi0619 n26979 ; n26982
g24547 nor pi1159 n26981 ; n26983
g24548 and n26982_not n26983 ; n26984
g24549 nor pi0648 n26857 ; n26985
g24550 and n26984_not n26985 ; n26986
g24551 nor pi0619 n26773 ; n26987
g24552 and pi0619 n26979_not ; n26988
g24553 and pi1159 n26987_not ; n26989
g24554 and n26988_not n26989 ; n26990
g24555 and pi0648 n26861_not ; n26991
g24556 and n26990_not n26991 ; n26992
g24557 and pi0789 n26986_not ; n26993
g24558 and n26992_not n26993 ; n26994
g24559 and n17970 n26980_not ; n26995
g24560 and n26994_not n26995 ; n26996
g24561 and n17871 n26775 ; n26997
g24562 nor pi0626 n26864 ; n26998
g24563 and pi0626 n26742_not ; n26999
g24564 and n16629 n26999_not ; n27000
g24565 and n26998_not n27000 ; n27001
g24566 and pi0626 n26864_not ; n27002
g24567 nor pi0626 n26742 ; n27003
g24568 and n16628 n27003_not ; n27004
g24569 and n27002_not n27004 ; n27005
g24570 nor n26997 n27001 ; n27006
g24571 and n27005_not n27006 ; n27007
g24572 and pi0788 n27007_not ; n27008
g24573 nor n20364 n27008 ; n27009
g24574 and n26996_not n27009 ; n27010
g24575 nor n26895 n27010 ; n27011
g24576 nor n20206 n27011 ; n27012
g24577 and n17802 n26793_not ; n27013
g24578 and n20559_not n26870 ; n27014
g24579 and n17801 n26797_not ; n27015
g24580 nor n27013 n27015 ; n27016
g24581 and n27014_not n27016 ; n27017
g24582 and pi0787 n27017_not ; n27018
g24583 and pi0644_not n26886 ; n27019
g24584 and pi0644 n26878 ; n27020
g24585 and pi0790 n27019_not ; n27021
g24586 and n27020_not n27021 ; n27022
g24587 nor n27012 n27018 ; n27023
g24588 and n27022_not n27023 ; n27024
g24589 nor n26889 n27024 ; n27025
g24590 nor po1038 n27025 ; n27026
g24591 nor pi0832 n26741 ; n27027
g24592 and n27026_not n27027 ; n27028
g24593 nor n26740 n27028 ; po0338
g24594 nor pi0182 n2926 ; n27030
g24595 and pi0734_not n16645 ; n27031
g24596 nor n27030 n27031 ; n27032
g24597 nor pi0778 n27032 ; n27033
g24598 and pi0625_not n27031 ; n27034
g24599 nor n27032 n27034 ; n27035
g24600 and pi1153 n27035_not ; n27036
g24601 nor pi1153 n27030 ; n27037
g24602 and n27034_not n27037 ; n27038
g24603 and pi0778 n27038_not ; n27039
g24604 and n27036_not n27039 ; n27040
g24605 nor n27033 n27040 ; n27041
g24606 nor n17845 n27041 ; n27042
g24607 and n17847_not n27042 ; n27043
g24608 and n17849_not n27043 ; n27044
g24609 and n17851_not n27044 ; n27045
g24610 and n17857_not n27045 ; n27046
g24611 and pi0647_not n27046 ; n27047
g24612 and pi0647 n27030 ; n27048
g24613 nor pi1157 n27048 ; n27049
g24614 and n27047_not n27049 ; n27050
g24615 and pi0630 n27050 ; n27051
g24616 and pi0756_not n17244 ; n27052
g24617 nor n27030 n27052 ; n27053
g24618 nor n17874 n27053 ; n27054
g24619 nor pi0785 n27054 ; n27055
g24620 and n17296 n27052 ; n27056
g24621 and n27054 n27056_not ; n27057
g24622 and pi1155 n27057_not ; n27058
g24623 nor pi1155 n27030 ; n27059
g24624 and n27056_not n27059 ; n27060
g24625 nor n27058 n27060 ; n27061
g24626 and pi0785 n27061_not ; n27062
g24627 nor n27055 n27062 ; n27063
g24628 nor pi0781 n27063 ; n27064
g24629 and n17889_not n27063 ; n27065
g24630 and pi1154 n27065_not ; n27066
g24631 and n17892_not n27063 ; n27067
g24632 nor pi1154 n27067 ; n27068
g24633 nor n27066 n27068 ; n27069
g24634 and pi0781 n27069_not ; n27070
g24635 nor n27064 n27070 ; n27071
g24636 nor pi0789 n27071 ; n27072
g24637 and n23078_not n27071 ; n27073
g24638 and pi1159 n27073_not ; n27074
g24639 and n23081_not n27071 ; n27075
g24640 nor pi1159 n27075 ; n27076
g24641 nor n27074 n27076 ; n27077
g24642 and pi0789 n27077_not ; n27078
g24643 nor n27072 n27078 ; n27079
g24644 and n17969_not n27079 ; n27080
g24645 and n17969 n27030 ; n27081
g24646 nor n27080 n27081 ; n27082
g24647 nor n17779 n27082 ; n27083
g24648 and n17779 n27030 ; n27084
g24649 nor n27083 n27084 ; n27085
g24650 and n20559_not n27085 ; n27086
g24651 and pi0647 n27046_not ; n27087
g24652 nor pi0647 n27030 ; n27088
g24653 nor n27087 n27088 ; n27089
g24654 and n17801 n27089_not ; n27090
g24655 nor n27051 n27090 ; n27091
g24656 and n27086_not n27091 ; n27092
g24657 and pi0787 n27092_not ; n27093
g24658 and n17871 n27044 ; n27094
g24659 nor pi0626 n27079 ; n27095
g24660 and pi0626 n27030_not ; n27096
g24661 and n16629 n27096_not ; n27097
g24662 and n27095_not n27097 ; n27098
g24663 and pi0626 n27079_not ; n27099
g24664 nor pi0626 n27030 ; n27100
g24665 and n16628 n27100_not ; n27101
g24666 and n27099_not n27101 ; n27102
g24667 nor n27094 n27098 ; n27103
g24668 and n27102_not n27103 ; n27104
g24669 and pi0788 n27104_not ; n27105
g24670 and pi0618 n27042 ; n27106
g24671 nor n17168 n27032 ; n27107
g24672 and pi0625 n27107 ; n27108
g24673 and n27053 n27107_not ; n27109
g24674 nor n27108 n27109 ; n27110
g24675 and n27037 n27110_not ; n27111
g24676 nor pi0608 n27036 ; n27112
g24677 and n27111_not n27112 ; n27113
g24678 and pi1153 n27053 ; n27114
g24679 and n27108_not n27114 ; n27115
g24680 and pi0608 n27038_not ; n27116
g24681 and n27115_not n27116 ; n27117
g24682 nor n27113 n27117 ; n27118
g24683 and pi0778 n27118_not ; n27119
g24684 nor pi0778 n27109 ; n27120
g24685 nor n27119 n27120 ; n27121
g24686 nor pi0609 n27121 ; n27122
g24687 and pi0609 n27041_not ; n27123
g24688 nor pi1155 n27123 ; n27124
g24689 and n27122_not n27124 ; n27125
g24690 nor pi0660 n27058 ; n27126
g24691 and n27125_not n27126 ; n27127
g24692 and pi0609 n27121_not ; n27128
g24693 nor pi0609 n27041 ; n27129
g24694 and pi1155 n27129_not ; n27130
g24695 and n27128_not n27130 ; n27131
g24696 and pi0660 n27060_not ; n27132
g24697 and n27131_not n27132 ; n27133
g24698 nor n27127 n27133 ; n27134
g24699 and pi0785 n27134_not ; n27135
g24700 nor pi0785 n27121 ; n27136
g24701 nor n27135 n27136 ; n27137
g24702 nor pi0618 n27137 ; n27138
g24703 nor pi1154 n27106 ; n27139
g24704 and n27138_not n27139 ; n27140
g24705 nor pi0627 n27066 ; n27141
g24706 and n27140_not n27141 ; n27142
g24707 and pi0618_not n27042 ; n27143
g24708 and pi0618 n27137_not ; n27144
g24709 and pi1154 n27143_not ; n27145
g24710 and n27144_not n27145 ; n27146
g24711 and pi0627 n27068_not ; n27147
g24712 and n27146_not n27147 ; n27148
g24713 nor n27142 n27148 ; n27149
g24714 and pi0781 n27149_not ; n27150
g24715 nor pi0781 n27137 ; n27151
g24716 nor n27150 n27151 ; n27152
g24717 and pi0789_not n27152 ; n27153
g24718 nor pi0619 n27152 ; n27154
g24719 and pi0619 n27043 ; n27155
g24720 nor pi1159 n27155 ; n27156
g24721 and n27154_not n27156 ; n27157
g24722 nor pi0648 n27074 ; n27158
g24723 and n27157_not n27158 ; n27159
g24724 and pi0619 n27152_not ; n27160
g24725 and pi0619_not n27043 ; n27161
g24726 and pi1159 n27161_not ; n27162
g24727 and n27160_not n27162 ; n27163
g24728 and pi0648 n27076_not ; n27164
g24729 and n27163_not n27164 ; n27165
g24730 and pi0789 n27159_not ; n27166
g24731 and n27165_not n27166 ; n27167
g24732 and n17970 n27153_not ; n27168
g24733 and n27167_not n27168 ; n27169
g24734 nor n27105 n27169 ; n27170
g24735 nor n20364 n27170 ; n27171
g24736 and n17854 n27082_not ; n27172
g24737 and n20851 n27045 ; n27173
g24738 nor n27172 n27173 ; n27174
g24739 nor pi0629 n27174 ; n27175
g24740 and n20855 n27045 ; n27176
g24741 and n17853 n27082_not ; n27177
g24742 nor n27176 n27177 ; n27178
g24743 and pi0629 n27178_not ; n27179
g24744 nor n27175 n27179 ; n27180
g24745 and pi0792 n27180_not ; n27181
g24746 nor n20206 n27181 ; n27182
g24747 and n27171_not n27182 ; n27183
g24748 nor n27093 n27183 ; n27184
g24749 and pi0790_not n27184 ; n27185
g24750 nor pi0787 n27046 ; n27186
g24751 and pi1157 n27089_not ; n27187
g24752 nor n27050 n27187 ; n27188
g24753 and pi0787 n27188_not ; n27189
g24754 nor n27186 n27189 ; n27190
g24755 and pi0644_not n27190 ; n27191
g24756 and pi0644 n27184 ; n27192
g24757 and pi0715 n27191_not ; n27193
g24758 and n27192_not n27193 ; n27194
g24759 nor n17804 n27085 ; n27195
g24760 and n17804 n27030 ; n27196
g24761 nor n27195 n27196 ; n27197
g24762 and pi0644 n27197_not ; n27198
g24763 and pi0644_not n27030 ; n27199
g24764 nor pi0715 n27199 ; n27200
g24765 and n27198_not n27200 ; n27201
g24766 and pi1160 n27201_not ; n27202
g24767 and n27194_not n27202 ; n27203
g24768 nor pi0644 n27197 ; n27204
g24769 and pi0644 n27030 ; n27205
g24770 and pi0715 n27205_not ; n27206
g24771 and n27204_not n27206 ; n27207
g24772 and pi0644 n27190 ; n27208
g24773 and pi0644_not n27184 ; n27209
g24774 nor pi0715 n27208 ; n27210
g24775 and n27209_not n27210 ; n27211
g24776 nor pi1160 n27207 ; n27212
g24777 and n27211_not n27212 ; n27213
g24778 nor n27203 n27213 ; n27214
g24779 and pi0790 n27214_not ; n27215
g24780 and pi0832 n27185_not ; n27216
g24781 and n27215_not n27216 ; n27217
g24782 and pi0182_not po1038 ; n27218
g24783 nor pi0182 n17059 ; n27219
g24784 and n16635 n27219_not ; n27220
g24785 and pi0734_not n2571 ; n27221
g24786 and n27219 n27221_not ; n27222
g24787 nor pi0182 n16641 ; n27223
g24788 and n16647 n27223_not ; n27224
g24789 and pi0182 n18076_not ; n27225
g24790 nor pi0038 n27225 ; n27226
g24791 and n2571 n27226_not ; n27227
g24792 and pi0182_not n18072 ; n27228
g24793 nor n27227 n27228 ; n27229
g24794 nor pi0734 n27224 ; n27230
g24795 and n27229_not n27230 ; n27231
g24796 nor n27222 n27231 ; n27232
g24797 and pi0778_not n27232 ; n27233
g24798 and pi0625_not n27219 ; n27234
g24799 and pi0625 n27232_not ; n27235
g24800 and pi1153 n27234_not ; n27236
g24801 and n27235_not n27236 ; n27237
g24802 and pi0625 n27219 ; n27238
g24803 nor pi0625 n27232 ; n27239
g24804 nor pi1153 n27238 ; n27240
g24805 and n27239_not n27240 ; n27241
g24806 nor n27237 n27241 ; n27242
g24807 and pi0778 n27242_not ; n27243
g24808 nor n27233 n27243 ; n27244
g24809 nor n17075 n27244 ; n27245
g24810 and n17075 n27219_not ; n27246
g24811 nor n27245 n27246 ; n27247
g24812 and n16639_not n27247 ; n27248
g24813 and n16639 n27219 ; n27249
g24814 nor n27248 n27249 ; n27250
g24815 and n16635_not n27250 ; n27251
g24816 nor n27220 n27251 ; n27252
g24817 and n16631_not n27252 ; n27253
g24818 and n16631 n27219 ; n27254
g24819 nor n27253 n27254 ; n27255
g24820 and pi0792_not n27255 ; n27256
g24821 and pi0628 n27255_not ; n27257
g24822 and pi0628_not n27219 ; n27258
g24823 and pi1156 n27258_not ; n27259
g24824 and n27257_not n27259 ; n27260
g24825 and pi0628 n27219 ; n27261
g24826 nor pi0628 n27255 ; n27262
g24827 nor pi1156 n27261 ; n27263
g24828 and n27262_not n27263 ; n27264
g24829 nor n27260 n27264 ; n27265
g24830 and pi0792 n27265_not ; n27266
g24831 nor n27256 n27266 ; n27267
g24832 nor pi0647 n27267 ; n27268
g24833 and pi0647 n27219_not ; n27269
g24834 nor n27268 n27269 ; n27270
g24835 and pi1157_not n27270 ; n27271
g24836 and pi0647 n27267_not ; n27272
g24837 nor pi0647 n27219 ; n27273
g24838 nor n27272 n27273 ; n27274
g24839 and pi1157 n27274 ; n27275
g24840 nor n27271 n27275 ; n27276
g24841 and pi0787 n27276_not ; n27277
g24842 and pi0787_not n27267 ; n27278
g24843 nor n27277 n27278 ; n27279
g24844 nor pi0644 n27279 ; n27280
g24845 and pi0715 n27280_not ; n27281
g24846 and pi0182 n2571_not ; n27282
g24847 and pi0756_not n17280 ; n27283
g24848 nor n27223 n27283 ; n27284
g24849 and pi0038 n27284_not ; n27285
g24850 and pi0182_not n17221 ; n27286
g24851 and pi0182 n17275_not ; n27287
g24852 nor pi0756 n27287 ; n27288
g24853 and n27286_not n27288 ; n27289
g24854 and pi0182_not pi0756 ; n27290
g24855 and n17048_not n27290 ; n27291
g24856 nor n27289 n27291 ; n27292
g24857 nor pi0038 n27292 ; n27293
g24858 nor n27285 n27293 ; n27294
g24859 and n2571 n27294 ; n27295
g24860 nor n27282 n27295 ; n27296
g24861 nor n17117 n27296 ; n27297
g24862 and n17117 n27219_not ; n27298
g24863 nor n27297 n27298 ; n27299
g24864 nor pi0785 n27299 ; n27300
g24865 nor n17291 n27219 ; n27301
g24866 and pi0609 n27297 ; n27302
g24867 nor n27301 n27302 ; n27303
g24868 and pi1155 n27303_not ; n27304
g24869 nor n17296 n27219 ; n27305
g24870 and pi0609_not n27297 ; n27306
g24871 nor n27305 n27306 ; n27307
g24872 nor pi1155 n27307 ; n27308
g24873 nor n27304 n27308 ; n27309
g24874 and pi0785 n27309_not ; n27310
g24875 nor n27300 n27310 ; n27311
g24876 nor pi0781 n27311 ; n27312
g24877 and pi0618_not n27219 ; n27313
g24878 and pi0618 n27311 ; n27314
g24879 and pi1154 n27313_not ; n27315
g24880 and n27314_not n27315 ; n27316
g24881 and pi0618_not n27311 ; n27317
g24882 and pi0618 n27219 ; n27318
g24883 nor pi1154 n27318 ; n27319
g24884 and n27317_not n27319 ; n27320
g24885 nor n27316 n27320 ; n27321
g24886 and pi0781 n27321_not ; n27322
g24887 nor n27312 n27322 ; n27323
g24888 nor pi0789 n27323 ; n27324
g24889 and pi0619_not n27219 ; n27325
g24890 and pi0619 n27323 ; n27326
g24891 and pi1159 n27325_not ; n27327
g24892 and n27326_not n27327 ; n27328
g24893 and pi0619_not n27323 ; n27329
g24894 and pi0619 n27219 ; n27330
g24895 nor pi1159 n27330 ; n27331
g24896 and n27329_not n27331 ; n27332
g24897 nor n27328 n27332 ; n27333
g24898 and pi0789 n27333_not ; n27334
g24899 nor n27324 n27334 ; n27335
g24900 and n17969_not n27335 ; n27336
g24901 and n17969 n27219 ; n27337
g24902 nor n27336 n27337 ; n27338
g24903 nor n17779 n27338 ; n27339
g24904 and n17779 n27219 ; n27340
g24905 nor n27339 n27340 ; n27341
g24906 nor n17804 n27341 ; n27342
g24907 and n17804 n27219 ; n27343
g24908 nor n27342 n27343 ; n27344
g24909 and pi0644 n27344_not ; n27345
g24910 and pi0644_not n27219 ; n27346
g24911 nor pi0715 n27346 ; n27347
g24912 and n27345_not n27347 ; n27348
g24913 and pi1160 n27348_not ; n27349
g24914 and n27281_not n27349 ; n27350
g24915 and pi0644 n27279_not ; n27351
g24916 nor pi0715 n27351 ; n27352
g24917 nor pi0644 n27344 ; n27353
g24918 and pi0644 n27219 ; n27354
g24919 and pi0715 n27354_not ; n27355
g24920 and n27353_not n27355 ; n27356
g24921 nor pi1160 n27356 ; n27357
g24922 and n27352_not n27357 ; n27358
g24923 nor n27350 n27358 ; n27359
g24924 and pi0790 n27359_not ; n27360
g24925 and pi0629_not n27260 ; n27361
g24926 and n20570_not n27338 ; n27362
g24927 and pi0629 n27264 ; n27363
g24928 nor n27361 n27363 ; n27364
g24929 and n27362_not n27364 ; n27365
g24930 and pi0792 n27365_not ; n27366
g24931 and pi0609 n27244 ; n27367
g24932 and pi0182 n17625_not ; n27368
g24933 nor pi0182 n17612 ; n27369
g24934 and pi0756 n27368_not ; n27370
g24935 and n27369_not n27370 ; n27371
g24936 and pi0182_not n17629 ; n27372
g24937 and pi0182 n17631 ; n27373
g24938 nor pi0756 n27373 ; n27374
g24939 and n27372_not n27374 ; n27375
g24940 nor n27371 n27375 ; n27376
g24941 nor pi0039 n27376 ; n27377
g24942 and pi0182 n17605 ; n27378
g24943 nor pi0182 n17546 ; n27379
g24944 nor pi0756 n27379 ; n27380
g24945 and n27378_not n27380 ; n27381
g24946 and pi0182_not n17404 ; n27382
g24947 and pi0182 n17485 ; n27383
g24948 and pi0756 n27383_not ; n27384
g24949 and n27382_not n27384 ; n27385
g24950 and pi0039 n27381_not ; n27386
g24951 and n27385_not n27386 ; n27387
g24952 nor pi0038 n27377 ; n27388
g24953 and n27387_not n27388 ; n27389
g24954 nor pi0756 n17490 ; n27390
g24955 and n19471 n27390_not ; n27391
g24956 nor pi0182 n27391 ; n27392
g24957 nor n17469 n27052 ; n27393
g24958 and pi0182 n27393_not ; n27394
g24959 and n6284 n27394 ; n27395
g24960 and pi0038 n27395_not ; n27396
g24961 and n27392_not n27396 ; n27397
g24962 nor pi0734 n27397 ; n27398
g24963 and n27389_not n27398 ; n27399
g24964 and pi0734 n27294_not ; n27400
g24965 and n2571 n27399_not ; n27401
g24966 and n27400_not n27401 ; n27402
g24967 nor n27282 n27402 ; n27403
g24968 and pi0625_not n27403 ; n27404
g24969 and pi0625 n27296 ; n27405
g24970 nor pi1153 n27405 ; n27406
g24971 and n27404_not n27406 ; n27407
g24972 nor pi0608 n27237 ; n27408
g24973 and n27407_not n27408 ; n27409
g24974 and pi0625_not n27296 ; n27410
g24975 and pi0625 n27403 ; n27411
g24976 and pi1153 n27410_not ; n27412
g24977 and n27411_not n27412 ; n27413
g24978 and pi0608 n27241_not ; n27414
g24979 and n27413_not n27414 ; n27415
g24980 nor n27409 n27415 ; n27416
g24981 and pi0778 n27416_not ; n27417
g24982 and pi0778_not n27403 ; n27418
g24983 nor n27417 n27418 ; n27419
g24984 nor pi0609 n27419 ; n27420
g24985 nor pi1155 n27367 ; n27421
g24986 and n27420_not n27421 ; n27422
g24987 nor pi0660 n27304 ; n27423
g24988 and n27422_not n27423 ; n27424
g24989 and pi0609_not n27244 ; n27425
g24990 and pi0609 n27419_not ; n27426
g24991 and pi1155 n27425_not ; n27427
g24992 and n27426_not n27427 ; n27428
g24993 and pi0660 n27308_not ; n27429
g24994 and n27428_not n27429 ; n27430
g24995 nor n27424 n27430 ; n27431
g24996 and pi0785 n27431_not ; n27432
g24997 nor pi0785 n27419 ; n27433
g24998 nor n27432 n27433 ; n27434
g24999 nor pi0618 n27434 ; n27435
g25000 and pi0618 n27247 ; n27436
g25001 nor pi1154 n27436 ; n27437
g25002 and n27435_not n27437 ; n27438
g25003 nor pi0627 n27316 ; n27439
g25004 and n27438_not n27439 ; n27440
g25005 and pi0618_not n27247 ; n27441
g25006 and pi0618 n27434_not ; n27442
g25007 and pi1154 n27441_not ; n27443
g25008 and n27442_not n27443 ; n27444
g25009 and pi0627 n27320_not ; n27445
g25010 and n27444_not n27445 ; n27446
g25011 nor n27440 n27446 ; n27447
g25012 and pi0781 n27447_not ; n27448
g25013 nor pi0781 n27434 ; n27449
g25014 nor n27448 n27449 ; n27450
g25015 and pi0789_not n27450 ; n27451
g25016 and pi0619 n27250_not ; n27452
g25017 nor pi0619 n27450 ; n27453
g25018 nor pi1159 n27452 ; n27454
g25019 and n27453_not n27454 ; n27455
g25020 nor pi0648 n27328 ; n27456
g25021 and n27455_not n27456 ; n27457
g25022 nor pi0619 n27250 ; n27458
g25023 and pi0619 n27450_not ; n27459
g25024 and pi1159 n27458_not ; n27460
g25025 and n27459_not n27460 ; n27461
g25026 and pi0648 n27332_not ; n27462
g25027 and n27461_not n27462 ; n27463
g25028 and pi0789 n27457_not ; n27464
g25029 and n27463_not n27464 ; n27465
g25030 and n17970 n27451_not ; n27466
g25031 and n27465_not n27466 ; n27467
g25032 and n17871 n27252 ; n27468
g25033 nor pi0626 n27335 ; n27469
g25034 and pi0626 n27219_not ; n27470
g25035 and n16629 n27470_not ; n27471
g25036 and n27469_not n27471 ; n27472
g25037 and pi0626 n27335_not ; n27473
g25038 nor pi0626 n27219 ; n27474
g25039 and n16628 n27474_not ; n27475
g25040 and n27473_not n27475 ; n27476
g25041 nor n27468 n27472 ; n27477
g25042 and n27476_not n27477 ; n27478
g25043 and pi0788 n27478_not ; n27479
g25044 nor n20364 n27479 ; n27480
g25045 and n27467_not n27480 ; n27481
g25046 nor n27366 n27481 ; n27482
g25047 nor n20206 n27482 ; n27483
g25048 and n17802 n27270_not ; n27484
g25049 and n20559_not n27341 ; n27485
g25050 and n17801 n27274_not ; n27486
g25051 nor n27484 n27486 ; n27487
g25052 and n27485_not n27487 ; n27488
g25053 and pi0787 n27488_not ; n27489
g25054 and pi0644_not n27357 ; n27490
g25055 and pi0644 n27349 ; n27491
g25056 and pi0790 n27490_not ; n27492
g25057 and n27491_not n27492 ; n27493
g25058 nor n27483 n27489 ; n27494
g25059 and n27493_not n27494 ; n27495
g25060 nor n27360 n27495 ; n27496
g25061 nor po1038 n27496 ; n27497
g25062 nor pi0832 n27218 ; n27498
g25063 and n27497_not n27498 ; n27499
g25064 nor n27217 n27499 ; po0339
g25065 nor pi0183 n2926 ; n27501
g25066 and pi0725_not n16645 ; n27502
g25067 nor n27501 n27502 ; n27503
g25068 nor pi0778 n27503 ; n27504
g25069 and pi0625_not n27502 ; n27505
g25070 nor n27503 n27505 ; n27506
g25071 and pi1153 n27506_not ; n27507
g25072 nor pi1153 n27501 ; n27508
g25073 and n27505_not n27508 ; n27509
g25074 and pi0778 n27509_not ; n27510
g25075 and n27507_not n27510 ; n27511
g25076 nor n27504 n27511 ; n27512
g25077 nor n17845 n27512 ; n27513
g25078 and n17847_not n27513 ; n27514
g25079 and n17849_not n27514 ; n27515
g25080 and n17851_not n27515 ; n27516
g25081 and n17857_not n27516 ; n27517
g25082 and pi0647_not n27517 ; n27518
g25083 and pi0647 n27501 ; n27519
g25084 nor pi1157 n27519 ; n27520
g25085 and n27518_not n27520 ; n27521
g25086 and pi0630 n27521 ; n27522
g25087 and pi0755_not n17244 ; n27523
g25088 nor n27501 n27523 ; n27524
g25089 nor n17874 n27524 ; n27525
g25090 nor pi0785 n27525 ; n27526
g25091 and n17296 n27523 ; n27527
g25092 and n27525 n27527_not ; n27528
g25093 and pi1155 n27528_not ; n27529
g25094 nor pi1155 n27501 ; n27530
g25095 and n27527_not n27530 ; n27531
g25096 nor n27529 n27531 ; n27532
g25097 and pi0785 n27532_not ; n27533
g25098 nor n27526 n27533 ; n27534
g25099 nor pi0781 n27534 ; n27535
g25100 and n17889_not n27534 ; n27536
g25101 and pi1154 n27536_not ; n27537
g25102 and n17892_not n27534 ; n27538
g25103 nor pi1154 n27538 ; n27539
g25104 nor n27537 n27539 ; n27540
g25105 and pi0781 n27540_not ; n27541
g25106 nor n27535 n27541 ; n27542
g25107 nor pi0789 n27542 ; n27543
g25108 and n23078_not n27542 ; n27544
g25109 and pi1159 n27544_not ; n27545
g25110 and n23081_not n27542 ; n27546
g25111 nor pi1159 n27546 ; n27547
g25112 nor n27545 n27547 ; n27548
g25113 and pi0789 n27548_not ; n27549
g25114 nor n27543 n27549 ; n27550
g25115 and n17969_not n27550 ; n27551
g25116 and n17969 n27501 ; n27552
g25117 nor n27551 n27552 ; n27553
g25118 nor n17779 n27553 ; n27554
g25119 and n17779 n27501 ; n27555
g25120 nor n27554 n27555 ; n27556
g25121 and n20559_not n27556 ; n27557
g25122 and pi0647 n27517_not ; n27558
g25123 nor pi0647 n27501 ; n27559
g25124 nor n27558 n27559 ; n27560
g25125 and n17801 n27560_not ; n27561
g25126 nor n27522 n27561 ; n27562
g25127 and n27557_not n27562 ; n27563
g25128 and pi0787 n27563_not ; n27564
g25129 and n17871 n27515 ; n27565
g25130 nor pi0626 n27550 ; n27566
g25131 and pi0626 n27501_not ; n27567
g25132 and n16629 n27567_not ; n27568
g25133 and n27566_not n27568 ; n27569
g25134 and pi0626 n27550_not ; n27570
g25135 nor pi0626 n27501 ; n27571
g25136 and n16628 n27571_not ; n27572
g25137 and n27570_not n27572 ; n27573
g25138 nor n27565 n27569 ; n27574
g25139 and n27573_not n27574 ; n27575
g25140 and pi0788 n27575_not ; n27576
g25141 and pi0618 n27513 ; n27577
g25142 nor n17168 n27503 ; n27578
g25143 and pi0625 n27578 ; n27579
g25144 and n27524 n27578_not ; n27580
g25145 nor n27579 n27580 ; n27581
g25146 and n27508 n27581_not ; n27582
g25147 nor pi0608 n27507 ; n27583
g25148 and n27582_not n27583 ; n27584
g25149 and pi1153 n27524 ; n27585
g25150 and n27579_not n27585 ; n27586
g25151 and pi0608 n27509_not ; n27587
g25152 and n27586_not n27587 ; n27588
g25153 nor n27584 n27588 ; n27589
g25154 and pi0778 n27589_not ; n27590
g25155 nor pi0778 n27580 ; n27591
g25156 nor n27590 n27591 ; n27592
g25157 nor pi0609 n27592 ; n27593
g25158 and pi0609 n27512_not ; n27594
g25159 nor pi1155 n27594 ; n27595
g25160 and n27593_not n27595 ; n27596
g25161 nor pi0660 n27529 ; n27597
g25162 and n27596_not n27597 ; n27598
g25163 and pi0609 n27592_not ; n27599
g25164 nor pi0609 n27512 ; n27600
g25165 and pi1155 n27600_not ; n27601
g25166 and n27599_not n27601 ; n27602
g25167 and pi0660 n27531_not ; n27603
g25168 and n27602_not n27603 ; n27604
g25169 nor n27598 n27604 ; n27605
g25170 and pi0785 n27605_not ; n27606
g25171 nor pi0785 n27592 ; n27607
g25172 nor n27606 n27607 ; n27608
g25173 nor pi0618 n27608 ; n27609
g25174 nor pi1154 n27577 ; n27610
g25175 and n27609_not n27610 ; n27611
g25176 nor pi0627 n27537 ; n27612
g25177 and n27611_not n27612 ; n27613
g25178 and pi0618_not n27513 ; n27614
g25179 and pi0618 n27608_not ; n27615
g25180 and pi1154 n27614_not ; n27616
g25181 and n27615_not n27616 ; n27617
g25182 and pi0627 n27539_not ; n27618
g25183 and n27617_not n27618 ; n27619
g25184 nor n27613 n27619 ; n27620
g25185 and pi0781 n27620_not ; n27621
g25186 nor pi0781 n27608 ; n27622
g25187 nor n27621 n27622 ; n27623
g25188 and pi0789_not n27623 ; n27624
g25189 nor pi0619 n27623 ; n27625
g25190 and pi0619 n27514 ; n27626
g25191 nor pi1159 n27626 ; n27627
g25192 and n27625_not n27627 ; n27628
g25193 nor pi0648 n27545 ; n27629
g25194 and n27628_not n27629 ; n27630
g25195 and pi0619 n27623_not ; n27631
g25196 and pi0619_not n27514 ; n27632
g25197 and pi1159 n27632_not ; n27633
g25198 and n27631_not n27633 ; n27634
g25199 and pi0648 n27547_not ; n27635
g25200 and n27634_not n27635 ; n27636
g25201 and pi0789 n27630_not ; n27637
g25202 and n27636_not n27637 ; n27638
g25203 and n17970 n27624_not ; n27639
g25204 and n27638_not n27639 ; n27640
g25205 nor n27576 n27640 ; n27641
g25206 nor n20364 n27641 ; n27642
g25207 and n17854 n27553_not ; n27643
g25208 and n20851 n27516 ; n27644
g25209 nor n27643 n27644 ; n27645
g25210 nor pi0629 n27645 ; n27646
g25211 and n20855 n27516 ; n27647
g25212 and n17853 n27553_not ; n27648
g25213 nor n27647 n27648 ; n27649
g25214 and pi0629 n27649_not ; n27650
g25215 nor n27646 n27650 ; n27651
g25216 and pi0792 n27651_not ; n27652
g25217 nor n20206 n27652 ; n27653
g25218 and n27642_not n27653 ; n27654
g25219 nor n27564 n27654 ; n27655
g25220 and pi0790_not n27655 ; n27656
g25221 nor pi0787 n27517 ; n27657
g25222 and pi1157 n27560_not ; n27658
g25223 nor n27521 n27658 ; n27659
g25224 and pi0787 n27659_not ; n27660
g25225 nor n27657 n27660 ; n27661
g25226 and pi0644_not n27661 ; n27662
g25227 and pi0644 n27655 ; n27663
g25228 and pi0715 n27662_not ; n27664
g25229 and n27663_not n27664 ; n27665
g25230 nor n17804 n27556 ; n27666
g25231 and n17804 n27501 ; n27667
g25232 nor n27666 n27667 ; n27668
g25233 and pi0644 n27668_not ; n27669
g25234 and pi0644_not n27501 ; n27670
g25235 nor pi0715 n27670 ; n27671
g25236 and n27669_not n27671 ; n27672
g25237 and pi1160 n27672_not ; n27673
g25238 and n27665_not n27673 ; n27674
g25239 nor pi0644 n27668 ; n27675
g25240 and pi0644 n27501 ; n27676
g25241 and pi0715 n27676_not ; n27677
g25242 and n27675_not n27677 ; n27678
g25243 and pi0644 n27661 ; n27679
g25244 and pi0644_not n27655 ; n27680
g25245 nor pi0715 n27679 ; n27681
g25246 and n27680_not n27681 ; n27682
g25247 nor pi1160 n27678 ; n27683
g25248 and n27682_not n27683 ; n27684
g25249 nor n27674 n27684 ; n27685
g25250 and pi0790 n27685_not ; n27686
g25251 and pi0832 n27656_not ; n27687
g25252 and n27686_not n27687 ; n27688
g25253 and pi0183_not po1038 ; n27689
g25254 nor pi0183 n17059 ; n27690
g25255 and n16635 n27690_not ; n27691
g25256 and pi0725_not n2571 ; n27692
g25257 and n27690 n27692_not ; n27693
g25258 nor pi0183 n16641 ; n27694
g25259 and n16647 n27694_not ; n27695
g25260 and pi0183 n18076_not ; n27696
g25261 nor pi0038 n27696 ; n27697
g25262 and n2571 n27697_not ; n27698
g25263 and pi0183_not n18072 ; n27699
g25264 nor n27698 n27699 ; n27700
g25265 nor pi0725 n27695 ; n27701
g25266 and n27700_not n27701 ; n27702
g25267 nor n27693 n27702 ; n27703
g25268 and pi0778_not n27703 ; n27704
g25269 and pi0625_not n27690 ; n27705
g25270 and pi0625 n27703_not ; n27706
g25271 and pi1153 n27705_not ; n27707
g25272 and n27706_not n27707 ; n27708
g25273 and pi0625 n27690 ; n27709
g25274 nor pi0625 n27703 ; n27710
g25275 nor pi1153 n27709 ; n27711
g25276 and n27710_not n27711 ; n27712
g25277 nor n27708 n27712 ; n27713
g25278 and pi0778 n27713_not ; n27714
g25279 nor n27704 n27714 ; n27715
g25280 nor n17075 n27715 ; n27716
g25281 and n17075 n27690_not ; n27717
g25282 nor n27716 n27717 ; n27718
g25283 and n16639_not n27718 ; n27719
g25284 and n16639 n27690 ; n27720
g25285 nor n27719 n27720 ; n27721
g25286 and n16635_not n27721 ; n27722
g25287 nor n27691 n27722 ; n27723
g25288 and n16631_not n27723 ; n27724
g25289 and n16631 n27690 ; n27725
g25290 nor n27724 n27725 ; n27726
g25291 and pi0792_not n27726 ; n27727
g25292 and pi0628 n27726_not ; n27728
g25293 and pi0628_not n27690 ; n27729
g25294 and pi1156 n27729_not ; n27730
g25295 and n27728_not n27730 ; n27731
g25296 and pi0628 n27690 ; n27732
g25297 nor pi0628 n27726 ; n27733
g25298 nor pi1156 n27732 ; n27734
g25299 and n27733_not n27734 ; n27735
g25300 nor n27731 n27735 ; n27736
g25301 and pi0792 n27736_not ; n27737
g25302 nor n27727 n27737 ; n27738
g25303 nor pi0647 n27738 ; n27739
g25304 and pi0647 n27690_not ; n27740
g25305 nor n27739 n27740 ; n27741
g25306 and pi1157_not n27741 ; n27742
g25307 and pi0647 n27738_not ; n27743
g25308 nor pi0647 n27690 ; n27744
g25309 nor n27743 n27744 ; n27745
g25310 and pi1157 n27745 ; n27746
g25311 nor n27742 n27746 ; n27747
g25312 and pi0787 n27747_not ; n27748
g25313 and pi0787_not n27738 ; n27749
g25314 nor n27748 n27749 ; n27750
g25315 nor pi0644 n27750 ; n27751
g25316 and pi0715 n27751_not ; n27752
g25317 and pi0183 n2571_not ; n27753
g25318 and pi0755_not n17280 ; n27754
g25319 nor n27694 n27754 ; n27755
g25320 and pi0038 n27755_not ; n27756
g25321 and pi0183_not n17221 ; n27757
g25322 and pi0183 n17275_not ; n27758
g25323 nor pi0755 n27758 ; n27759
g25324 and n27757_not n27759 ; n27760
g25325 and pi0183_not pi0755 ; n27761
g25326 and n17048_not n27761 ; n27762
g25327 nor n27760 n27762 ; n27763
g25328 nor pi0038 n27763 ; n27764
g25329 nor n27756 n27764 ; n27765
g25330 and n2571 n27765 ; n27766
g25331 nor n27753 n27766 ; n27767
g25332 nor n17117 n27767 ; n27768
g25333 and n17117 n27690_not ; n27769
g25334 nor n27768 n27769 ; n27770
g25335 nor pi0785 n27770 ; n27771
g25336 nor n17291 n27690 ; n27772
g25337 and pi0609 n27768 ; n27773
g25338 nor n27772 n27773 ; n27774
g25339 and pi1155 n27774_not ; n27775
g25340 nor n17296 n27690 ; n27776
g25341 and pi0609_not n27768 ; n27777
g25342 nor n27776 n27777 ; n27778
g25343 nor pi1155 n27778 ; n27779
g25344 nor n27775 n27779 ; n27780
g25345 and pi0785 n27780_not ; n27781
g25346 nor n27771 n27781 ; n27782
g25347 nor pi0781 n27782 ; n27783
g25348 and pi0618_not n27690 ; n27784
g25349 and pi0618 n27782 ; n27785
g25350 and pi1154 n27784_not ; n27786
g25351 and n27785_not n27786 ; n27787
g25352 and pi0618_not n27782 ; n27788
g25353 and pi0618 n27690 ; n27789
g25354 nor pi1154 n27789 ; n27790
g25355 and n27788_not n27790 ; n27791
g25356 nor n27787 n27791 ; n27792
g25357 and pi0781 n27792_not ; n27793
g25358 nor n27783 n27793 ; n27794
g25359 nor pi0789 n27794 ; n27795
g25360 and pi0619_not n27690 ; n27796
g25361 and pi0619 n27794 ; n27797
g25362 and pi1159 n27796_not ; n27798
g25363 and n27797_not n27798 ; n27799
g25364 and pi0619_not n27794 ; n27800
g25365 and pi0619 n27690 ; n27801
g25366 nor pi1159 n27801 ; n27802
g25367 and n27800_not n27802 ; n27803
g25368 nor n27799 n27803 ; n27804
g25369 and pi0789 n27804_not ; n27805
g25370 nor n27795 n27805 ; n27806
g25371 and n17969_not n27806 ; n27807
g25372 and n17969 n27690 ; n27808
g25373 nor n27807 n27808 ; n27809
g25374 nor n17779 n27809 ; n27810
g25375 and n17779 n27690 ; n27811
g25376 nor n27810 n27811 ; n27812
g25377 nor n17804 n27812 ; n27813
g25378 and n17804 n27690 ; n27814
g25379 nor n27813 n27814 ; n27815
g25380 and pi0644 n27815_not ; n27816
g25381 and pi0644_not n27690 ; n27817
g25382 nor pi0715 n27817 ; n27818
g25383 and n27816_not n27818 ; n27819
g25384 and pi1160 n27819_not ; n27820
g25385 and n27752_not n27820 ; n27821
g25386 and pi0644 n27750_not ; n27822
g25387 nor pi0715 n27822 ; n27823
g25388 nor pi0644 n27815 ; n27824
g25389 and pi0644 n27690 ; n27825
g25390 and pi0715 n27825_not ; n27826
g25391 and n27824_not n27826 ; n27827
g25392 nor pi1160 n27827 ; n27828
g25393 and n27823_not n27828 ; n27829
g25394 nor n27821 n27829 ; n27830
g25395 and pi0790 n27830_not ; n27831
g25396 and pi0629_not n27731 ; n27832
g25397 and n20570_not n27809 ; n27833
g25398 and pi0629 n27735 ; n27834
g25399 nor n27832 n27834 ; n27835
g25400 and n27833_not n27835 ; n27836
g25401 and pi0792 n27836_not ; n27837
g25402 and pi0609 n27715 ; n27838
g25403 and pi0183 n17625_not ; n27839
g25404 nor pi0183 n17612 ; n27840
g25405 and pi0755 n27839_not ; n27841
g25406 and n27840_not n27841 ; n27842
g25407 and pi0183_not n17629 ; n27843
g25408 and pi0183 n17631 ; n27844
g25409 nor pi0755 n27844 ; n27845
g25410 and n27843_not n27845 ; n27846
g25411 nor n27842 n27846 ; n27847
g25412 nor pi0039 n27847 ; n27848
g25413 and pi0183 n17605 ; n27849
g25414 nor pi0183 n17546 ; n27850
g25415 nor pi0755 n27850 ; n27851
g25416 and n27849_not n27851 ; n27852
g25417 and pi0183_not n17404 ; n27853
g25418 and pi0183 n17485 ; n27854
g25419 and pi0755 n27854_not ; n27855
g25420 and n27853_not n27855 ; n27856
g25421 and pi0039 n27852_not ; n27857
g25422 and n27856_not n27857 ; n27858
g25423 nor pi0038 n27848 ; n27859
g25424 and n27858_not n27859 ; n27860
g25425 nor pi0755 n17490 ; n27861
g25426 and n19471 n27861_not ; n27862
g25427 nor pi0183 n27862 ; n27863
g25428 nor n17469 n27523 ; n27864
g25429 and pi0183 n27864_not ; n27865
g25430 and n6284 n27865 ; n27866
g25431 and pi0038 n27866_not ; n27867
g25432 and n27863_not n27867 ; n27868
g25433 nor pi0725 n27868 ; n27869
g25434 and n27860_not n27869 ; n27870
g25435 and pi0725 n27765_not ; n27871
g25436 and n2571 n27870_not ; n27872
g25437 and n27871_not n27872 ; n27873
g25438 nor n27753 n27873 ; n27874
g25439 and pi0625_not n27874 ; n27875
g25440 and pi0625 n27767 ; n27876
g25441 nor pi1153 n27876 ; n27877
g25442 and n27875_not n27877 ; n27878
g25443 nor pi0608 n27708 ; n27879
g25444 and n27878_not n27879 ; n27880
g25445 and pi0625_not n27767 ; n27881
g25446 and pi0625 n27874 ; n27882
g25447 and pi1153 n27881_not ; n27883
g25448 and n27882_not n27883 ; n27884
g25449 and pi0608 n27712_not ; n27885
g25450 and n27884_not n27885 ; n27886
g25451 nor n27880 n27886 ; n27887
g25452 and pi0778 n27887_not ; n27888
g25453 and pi0778_not n27874 ; n27889
g25454 nor n27888 n27889 ; n27890
g25455 nor pi0609 n27890 ; n27891
g25456 nor pi1155 n27838 ; n27892
g25457 and n27891_not n27892 ; n27893
g25458 nor pi0660 n27775 ; n27894
g25459 and n27893_not n27894 ; n27895
g25460 and pi0609_not n27715 ; n27896
g25461 and pi0609 n27890_not ; n27897
g25462 and pi1155 n27896_not ; n27898
g25463 and n27897_not n27898 ; n27899
g25464 and pi0660 n27779_not ; n27900
g25465 and n27899_not n27900 ; n27901
g25466 nor n27895 n27901 ; n27902
g25467 and pi0785 n27902_not ; n27903
g25468 nor pi0785 n27890 ; n27904
g25469 nor n27903 n27904 ; n27905
g25470 nor pi0618 n27905 ; n27906
g25471 and pi0618 n27718 ; n27907
g25472 nor pi1154 n27907 ; n27908
g25473 and n27906_not n27908 ; n27909
g25474 nor pi0627 n27787 ; n27910
g25475 and n27909_not n27910 ; n27911
g25476 and pi0618_not n27718 ; n27912
g25477 and pi0618 n27905_not ; n27913
g25478 and pi1154 n27912_not ; n27914
g25479 and n27913_not n27914 ; n27915
g25480 and pi0627 n27791_not ; n27916
g25481 and n27915_not n27916 ; n27917
g25482 nor n27911 n27917 ; n27918
g25483 and pi0781 n27918_not ; n27919
g25484 nor pi0781 n27905 ; n27920
g25485 nor n27919 n27920 ; n27921
g25486 and pi0789_not n27921 ; n27922
g25487 and pi0619 n27721_not ; n27923
g25488 nor pi0619 n27921 ; n27924
g25489 nor pi1159 n27923 ; n27925
g25490 and n27924_not n27925 ; n27926
g25491 nor pi0648 n27799 ; n27927
g25492 and n27926_not n27927 ; n27928
g25493 nor pi0619 n27721 ; n27929
g25494 and pi0619 n27921_not ; n27930
g25495 and pi1159 n27929_not ; n27931
g25496 and n27930_not n27931 ; n27932
g25497 and pi0648 n27803_not ; n27933
g25498 and n27932_not n27933 ; n27934
g25499 and pi0789 n27928_not ; n27935
g25500 and n27934_not n27935 ; n27936
g25501 and n17970 n27922_not ; n27937
g25502 and n27936_not n27937 ; n27938
g25503 and n17871 n27723 ; n27939
g25504 nor pi0626 n27806 ; n27940
g25505 and pi0626 n27690_not ; n27941
g25506 and n16629 n27941_not ; n27942
g25507 and n27940_not n27942 ; n27943
g25508 and pi0626 n27806_not ; n27944
g25509 nor pi0626 n27690 ; n27945
g25510 and n16628 n27945_not ; n27946
g25511 and n27944_not n27946 ; n27947
g25512 nor n27939 n27943 ; n27948
g25513 and n27947_not n27948 ; n27949
g25514 and pi0788 n27949_not ; n27950
g25515 nor n20364 n27950 ; n27951
g25516 and n27938_not n27951 ; n27952
g25517 nor n27837 n27952 ; n27953
g25518 nor n20206 n27953 ; n27954
g25519 and n17802 n27741_not ; n27955
g25520 and n20559_not n27812 ; n27956
g25521 and n17801 n27745_not ; n27957
g25522 nor n27955 n27957 ; n27958
g25523 and n27956_not n27958 ; n27959
g25524 and pi0787 n27959_not ; n27960
g25525 and pi0644_not n27828 ; n27961
g25526 and pi0644 n27820 ; n27962
g25527 and pi0790 n27961_not ; n27963
g25528 and n27962_not n27963 ; n27964
g25529 nor n27954 n27960 ; n27965
g25530 and n27964_not n27965 ; n27966
g25531 nor n27831 n27966 ; n27967
g25532 nor po1038 n27967 ; n27968
g25533 nor pi0832 n27689 ; n27969
g25534 and n27968_not n27969 ; n27970
g25535 nor n27688 n27970 ; po0340
g25536 nor pi0184 n2926 ; n27972
g25537 and pi0737_not n16645 ; n27973
g25538 nor n27972 n27973 ; n27974
g25539 nor pi0778 n27974 ; n27975
g25540 and pi0625_not n27973 ; n27976
g25541 nor n27974 n27976 ; n27977
g25542 and pi1153 n27977_not ; n27978
g25543 nor pi1153 n27972 ; n27979
g25544 and n27976_not n27979 ; n27980
g25545 and pi0778 n27980_not ; n27981
g25546 and n27978_not n27981 ; n27982
g25547 nor n27975 n27982 ; n27983
g25548 nor n17845 n27983 ; n27984
g25549 and n17847_not n27984 ; n27985
g25550 and n17849_not n27985 ; n27986
g25551 and n17851_not n27986 ; n27987
g25552 and n17857_not n27987 ; n27988
g25553 and pi0647_not n27988 ; n27989
g25554 and pi0647 n27972 ; n27990
g25555 nor pi1157 n27990 ; n27991
g25556 and n27989_not n27991 ; n27992
g25557 and pi0630 n27992 ; n27993
g25558 and pi0777_not n17244 ; n27994
g25559 nor n27972 n27994 ; n27995
g25560 nor n17874 n27995 ; n27996
g25561 nor pi0785 n27996 ; n27997
g25562 and n17296 n27994 ; n27998
g25563 and n27996 n27998_not ; n27999
g25564 and pi1155 n27999_not ; n28000
g25565 nor pi1155 n27972 ; n28001
g25566 and n27998_not n28001 ; n28002
g25567 nor n28000 n28002 ; n28003
g25568 and pi0785 n28003_not ; n28004
g25569 nor n27997 n28004 ; n28005
g25570 nor pi0781 n28005 ; n28006
g25571 and n17889_not n28005 ; n28007
g25572 and pi1154 n28007_not ; n28008
g25573 and n17892_not n28005 ; n28009
g25574 nor pi1154 n28009 ; n28010
g25575 nor n28008 n28010 ; n28011
g25576 and pi0781 n28011_not ; n28012
g25577 nor n28006 n28012 ; n28013
g25578 nor pi0789 n28013 ; n28014
g25579 and n23078_not n28013 ; n28015
g25580 and pi1159 n28015_not ; n28016
g25581 and n23081_not n28013 ; n28017
g25582 nor pi1159 n28017 ; n28018
g25583 nor n28016 n28018 ; n28019
g25584 and pi0789 n28019_not ; n28020
g25585 nor n28014 n28020 ; n28021
g25586 and n17969_not n28021 ; n28022
g25587 and n17969 n27972 ; n28023
g25588 nor n28022 n28023 ; n28024
g25589 nor n17779 n28024 ; n28025
g25590 and n17779 n27972 ; n28026
g25591 nor n28025 n28026 ; n28027
g25592 and n20559_not n28027 ; n28028
g25593 and pi0647 n27988_not ; n28029
g25594 nor pi0647 n27972 ; n28030
g25595 nor n28029 n28030 ; n28031
g25596 and n17801 n28031_not ; n28032
g25597 nor n27993 n28032 ; n28033
g25598 and n28028_not n28033 ; n28034
g25599 and pi0787 n28034_not ; n28035
g25600 and n17871 n27986 ; n28036
g25601 nor pi0626 n28021 ; n28037
g25602 and pi0626 n27972_not ; n28038
g25603 and n16629 n28038_not ; n28039
g25604 and n28037_not n28039 ; n28040
g25605 and pi0626 n28021_not ; n28041
g25606 nor pi0626 n27972 ; n28042
g25607 and n16628 n28042_not ; n28043
g25608 and n28041_not n28043 ; n28044
g25609 nor n28036 n28040 ; n28045
g25610 and n28044_not n28045 ; n28046
g25611 and pi0788 n28046_not ; n28047
g25612 and pi0618 n27984 ; n28048
g25613 nor n17168 n27974 ; n28049
g25614 and pi0625 n28049 ; n28050
g25615 and n27995 n28049_not ; n28051
g25616 nor n28050 n28051 ; n28052
g25617 and n27979 n28052_not ; n28053
g25618 nor pi0608 n27978 ; n28054
g25619 and n28053_not n28054 ; n28055
g25620 and pi1153 n27995 ; n28056
g25621 and n28050_not n28056 ; n28057
g25622 and pi0608 n27980_not ; n28058
g25623 and n28057_not n28058 ; n28059
g25624 nor n28055 n28059 ; n28060
g25625 and pi0778 n28060_not ; n28061
g25626 nor pi0778 n28051 ; n28062
g25627 nor n28061 n28062 ; n28063
g25628 nor pi0609 n28063 ; n28064
g25629 and pi0609 n27983_not ; n28065
g25630 nor pi1155 n28065 ; n28066
g25631 and n28064_not n28066 ; n28067
g25632 nor pi0660 n28000 ; n28068
g25633 and n28067_not n28068 ; n28069
g25634 and pi0609 n28063_not ; n28070
g25635 nor pi0609 n27983 ; n28071
g25636 and pi1155 n28071_not ; n28072
g25637 and n28070_not n28072 ; n28073
g25638 and pi0660 n28002_not ; n28074
g25639 and n28073_not n28074 ; n28075
g25640 nor n28069 n28075 ; n28076
g25641 and pi0785 n28076_not ; n28077
g25642 nor pi0785 n28063 ; n28078
g25643 nor n28077 n28078 ; n28079
g25644 nor pi0618 n28079 ; n28080
g25645 nor pi1154 n28048 ; n28081
g25646 and n28080_not n28081 ; n28082
g25647 nor pi0627 n28008 ; n28083
g25648 and n28082_not n28083 ; n28084
g25649 and pi0618_not n27984 ; n28085
g25650 and pi0618 n28079_not ; n28086
g25651 and pi1154 n28085_not ; n28087
g25652 and n28086_not n28087 ; n28088
g25653 and pi0627 n28010_not ; n28089
g25654 and n28088_not n28089 ; n28090
g25655 nor n28084 n28090 ; n28091
g25656 and pi0781 n28091_not ; n28092
g25657 nor pi0781 n28079 ; n28093
g25658 nor n28092 n28093 ; n28094
g25659 and pi0789_not n28094 ; n28095
g25660 nor pi0619 n28094 ; n28096
g25661 and pi0619 n27985 ; n28097
g25662 nor pi1159 n28097 ; n28098
g25663 and n28096_not n28098 ; n28099
g25664 nor pi0648 n28016 ; n28100
g25665 and n28099_not n28100 ; n28101
g25666 and pi0619 n28094_not ; n28102
g25667 and pi0619_not n27985 ; n28103
g25668 and pi1159 n28103_not ; n28104
g25669 and n28102_not n28104 ; n28105
g25670 and pi0648 n28018_not ; n28106
g25671 and n28105_not n28106 ; n28107
g25672 and pi0789 n28101_not ; n28108
g25673 and n28107_not n28108 ; n28109
g25674 and n17970 n28095_not ; n28110
g25675 and n28109_not n28110 ; n28111
g25676 nor n28047 n28111 ; n28112
g25677 nor n20364 n28112 ; n28113
g25678 and n17854 n28024_not ; n28114
g25679 and n20851 n27987 ; n28115
g25680 nor n28114 n28115 ; n28116
g25681 nor pi0629 n28116 ; n28117
g25682 and n20855 n27987 ; n28118
g25683 and n17853 n28024_not ; n28119
g25684 nor n28118 n28119 ; n28120
g25685 and pi0629 n28120_not ; n28121
g25686 nor n28117 n28121 ; n28122
g25687 and pi0792 n28122_not ; n28123
g25688 nor n20206 n28123 ; n28124
g25689 and n28113_not n28124 ; n28125
g25690 nor n28035 n28125 ; n28126
g25691 and pi0790_not n28126 ; n28127
g25692 nor pi0787 n27988 ; n28128
g25693 and pi1157 n28031_not ; n28129
g25694 nor n27992 n28129 ; n28130
g25695 and pi0787 n28130_not ; n28131
g25696 nor n28128 n28131 ; n28132
g25697 and pi0644_not n28132 ; n28133
g25698 and pi0644 n28126 ; n28134
g25699 and pi0715 n28133_not ; n28135
g25700 and n28134_not n28135 ; n28136
g25701 nor n17804 n28027 ; n28137
g25702 and n17804 n27972 ; n28138
g25703 nor n28137 n28138 ; n28139
g25704 and pi0644 n28139_not ; n28140
g25705 and pi0644_not n27972 ; n28141
g25706 nor pi0715 n28141 ; n28142
g25707 and n28140_not n28142 ; n28143
g25708 and pi1160 n28143_not ; n28144
g25709 and n28136_not n28144 ; n28145
g25710 nor pi0644 n28139 ; n28146
g25711 and pi0644 n27972 ; n28147
g25712 and pi0715 n28147_not ; n28148
g25713 and n28146_not n28148 ; n28149
g25714 and pi0644 n28132 ; n28150
g25715 and pi0644_not n28126 ; n28151
g25716 nor pi0715 n28150 ; n28152
g25717 and n28151_not n28152 ; n28153
g25718 nor pi1160 n28149 ; n28154
g25719 and n28153_not n28154 ; n28155
g25720 nor n28145 n28155 ; n28156
g25721 and pi0790 n28156_not ; n28157
g25722 and pi0832 n28127_not ; n28158
g25723 and n28157_not n28158 ; n28159
g25724 and pi0184_not po1038 ; n28160
g25725 nor pi0184 n17059 ; n28161
g25726 and n16635 n28161_not ; n28162
g25727 and pi0737_not n2571 ; n28163
g25728 and n28161 n28163_not ; n28164
g25729 nor pi0184 n16641 ; n28165
g25730 and n16647 n28165_not ; n28166
g25731 and pi0184 n18076_not ; n28167
g25732 nor pi0038 n28167 ; n28168
g25733 and n2571 n28168_not ; n28169
g25734 and pi0184_not n18072 ; n28170
g25735 nor n28169 n28170 ; n28171
g25736 nor pi0737 n28166 ; n28172
g25737 and n28171_not n28172 ; n28173
g25738 nor n28164 n28173 ; n28174
g25739 and pi0778_not n28174 ; n28175
g25740 and pi0625_not n28161 ; n28176
g25741 and pi0625 n28174_not ; n28177
g25742 and pi1153 n28176_not ; n28178
g25743 and n28177_not n28178 ; n28179
g25744 and pi0625 n28161 ; n28180
g25745 nor pi0625 n28174 ; n28181
g25746 nor pi1153 n28180 ; n28182
g25747 and n28181_not n28182 ; n28183
g25748 nor n28179 n28183 ; n28184
g25749 and pi0778 n28184_not ; n28185
g25750 nor n28175 n28185 ; n28186
g25751 nor n17075 n28186 ; n28187
g25752 and n17075 n28161_not ; n28188
g25753 nor n28187 n28188 ; n28189
g25754 and n16639_not n28189 ; n28190
g25755 and n16639 n28161 ; n28191
g25756 nor n28190 n28191 ; n28192
g25757 and n16635_not n28192 ; n28193
g25758 nor n28162 n28193 ; n28194
g25759 and n16631_not n28194 ; n28195
g25760 and n16631 n28161 ; n28196
g25761 nor n28195 n28196 ; n28197
g25762 and pi0792_not n28197 ; n28198
g25763 and pi0628 n28197_not ; n28199
g25764 and pi0628_not n28161 ; n28200
g25765 and pi1156 n28200_not ; n28201
g25766 and n28199_not n28201 ; n28202
g25767 and pi0628 n28161 ; n28203
g25768 nor pi0628 n28197 ; n28204
g25769 nor pi1156 n28203 ; n28205
g25770 and n28204_not n28205 ; n28206
g25771 nor n28202 n28206 ; n28207
g25772 and pi0792 n28207_not ; n28208
g25773 nor n28198 n28208 ; n28209
g25774 nor pi0647 n28209 ; n28210
g25775 and pi0647 n28161_not ; n28211
g25776 nor n28210 n28211 ; n28212
g25777 and pi1157_not n28212 ; n28213
g25778 and pi0647 n28209_not ; n28214
g25779 nor pi0647 n28161 ; n28215
g25780 nor n28214 n28215 ; n28216
g25781 and pi1157 n28216 ; n28217
g25782 nor n28213 n28217 ; n28218
g25783 and pi0787 n28218_not ; n28219
g25784 and pi0787_not n28209 ; n28220
g25785 nor n28219 n28220 ; n28221
g25786 nor pi0644 n28221 ; n28222
g25787 and pi0715 n28222_not ; n28223
g25788 and pi0184 n2571_not ; n28224
g25789 and pi0777_not n17280 ; n28225
g25790 nor n28165 n28225 ; n28226
g25791 and pi0038 n28226_not ; n28227
g25792 and pi0184_not n17221 ; n28228
g25793 and pi0184 n17275_not ; n28229
g25794 nor pi0777 n28229 ; n28230
g25795 and n28228_not n28230 ; n28231
g25796 and pi0184_not pi0777 ; n28232
g25797 and n17048_not n28232 ; n28233
g25798 nor n28231 n28233 ; n28234
g25799 nor pi0038 n28234 ; n28235
g25800 nor n28227 n28235 ; n28236
g25801 and n2571 n28236 ; n28237
g25802 nor n28224 n28237 ; n28238
g25803 nor n17117 n28238 ; n28239
g25804 and n17117 n28161_not ; n28240
g25805 nor n28239 n28240 ; n28241
g25806 nor pi0785 n28241 ; n28242
g25807 nor n17291 n28161 ; n28243
g25808 and pi0609 n28239 ; n28244
g25809 nor n28243 n28244 ; n28245
g25810 and pi1155 n28245_not ; n28246
g25811 nor n17296 n28161 ; n28247
g25812 and pi0609_not n28239 ; n28248
g25813 nor n28247 n28248 ; n28249
g25814 nor pi1155 n28249 ; n28250
g25815 nor n28246 n28250 ; n28251
g25816 and pi0785 n28251_not ; n28252
g25817 nor n28242 n28252 ; n28253
g25818 nor pi0781 n28253 ; n28254
g25819 and pi0618_not n28161 ; n28255
g25820 and pi0618 n28253 ; n28256
g25821 and pi1154 n28255_not ; n28257
g25822 and n28256_not n28257 ; n28258
g25823 and pi0618_not n28253 ; n28259
g25824 and pi0618 n28161 ; n28260
g25825 nor pi1154 n28260 ; n28261
g25826 and n28259_not n28261 ; n28262
g25827 nor n28258 n28262 ; n28263
g25828 and pi0781 n28263_not ; n28264
g25829 nor n28254 n28264 ; n28265
g25830 nor pi0789 n28265 ; n28266
g25831 and pi0619_not n28161 ; n28267
g25832 and pi0619 n28265 ; n28268
g25833 and pi1159 n28267_not ; n28269
g25834 and n28268_not n28269 ; n28270
g25835 and pi0619_not n28265 ; n28271
g25836 and pi0619 n28161 ; n28272
g25837 nor pi1159 n28272 ; n28273
g25838 and n28271_not n28273 ; n28274
g25839 nor n28270 n28274 ; n28275
g25840 and pi0789 n28275_not ; n28276
g25841 nor n28266 n28276 ; n28277
g25842 and n17969_not n28277 ; n28278
g25843 and n17969 n28161 ; n28279
g25844 nor n28278 n28279 ; n28280
g25845 nor n17779 n28280 ; n28281
g25846 and n17779 n28161 ; n28282
g25847 nor n28281 n28282 ; n28283
g25848 nor n17804 n28283 ; n28284
g25849 and n17804 n28161 ; n28285
g25850 nor n28284 n28285 ; n28286
g25851 and pi0644 n28286_not ; n28287
g25852 and pi0644_not n28161 ; n28288
g25853 nor pi0715 n28288 ; n28289
g25854 and n28287_not n28289 ; n28290
g25855 and pi1160 n28290_not ; n28291
g25856 and n28223_not n28291 ; n28292
g25857 and pi0644 n28221_not ; n28293
g25858 nor pi0715 n28293 ; n28294
g25859 nor pi0644 n28286 ; n28295
g25860 and pi0644 n28161 ; n28296
g25861 and pi0715 n28296_not ; n28297
g25862 and n28295_not n28297 ; n28298
g25863 nor pi1160 n28298 ; n28299
g25864 and n28294_not n28299 ; n28300
g25865 nor n28292 n28300 ; n28301
g25866 and pi0790 n28301_not ; n28302
g25867 and pi0629_not n28202 ; n28303
g25868 and n20570_not n28280 ; n28304
g25869 and pi0629 n28206 ; n28305
g25870 nor n28303 n28305 ; n28306
g25871 and n28304_not n28306 ; n28307
g25872 and pi0792 n28307_not ; n28308
g25873 and pi0609 n28186 ; n28309
g25874 and pi0184 n17625_not ; n28310
g25875 nor pi0184 n17612 ; n28311
g25876 and pi0777 n28310_not ; n28312
g25877 and n28311_not n28312 ; n28313
g25878 and pi0184_not n17629 ; n28314
g25879 and pi0184 n17631 ; n28315
g25880 nor pi0777 n28315 ; n28316
g25881 and n28314_not n28316 ; n28317
g25882 nor n28313 n28317 ; n28318
g25883 nor pi0039 n28318 ; n28319
g25884 and pi0184 n17605 ; n28320
g25885 nor pi0184 n17546 ; n28321
g25886 nor pi0777 n28321 ; n28322
g25887 and n28320_not n28322 ; n28323
g25888 and pi0184_not n17404 ; n28324
g25889 and pi0184 n17485 ; n28325
g25890 and pi0777 n28325_not ; n28326
g25891 and n28324_not n28326 ; n28327
g25892 and pi0039 n28323_not ; n28328
g25893 and n28327_not n28328 ; n28329
g25894 nor pi0038 n28319 ; n28330
g25895 and n28329_not n28330 ; n28331
g25896 nor pi0777 n17490 ; n28332
g25897 and n19471 n28332_not ; n28333
g25898 nor pi0184 n28333 ; n28334
g25899 nor n17469 n27994 ; n28335
g25900 and pi0184 n28335_not ; n28336
g25901 and n6284 n28336 ; n28337
g25902 and pi0038 n28337_not ; n28338
g25903 and n28334_not n28338 ; n28339
g25904 nor pi0737 n28339 ; n28340
g25905 and n28331_not n28340 ; n28341
g25906 and pi0737 n28236_not ; n28342
g25907 and n2571 n28341_not ; n28343
g25908 and n28342_not n28343 ; n28344
g25909 nor n28224 n28344 ; n28345
g25910 and pi0625_not n28345 ; n28346
g25911 and pi0625 n28238 ; n28347
g25912 nor pi1153 n28347 ; n28348
g25913 and n28346_not n28348 ; n28349
g25914 nor pi0608 n28179 ; n28350
g25915 and n28349_not n28350 ; n28351
g25916 and pi0625_not n28238 ; n28352
g25917 and pi0625 n28345 ; n28353
g25918 and pi1153 n28352_not ; n28354
g25919 and n28353_not n28354 ; n28355
g25920 and pi0608 n28183_not ; n28356
g25921 and n28355_not n28356 ; n28357
g25922 nor n28351 n28357 ; n28358
g25923 and pi0778 n28358_not ; n28359
g25924 and pi0778_not n28345 ; n28360
g25925 nor n28359 n28360 ; n28361
g25926 nor pi0609 n28361 ; n28362
g25927 nor pi1155 n28309 ; n28363
g25928 and n28362_not n28363 ; n28364
g25929 nor pi0660 n28246 ; n28365
g25930 and n28364_not n28365 ; n28366
g25931 and pi0609_not n28186 ; n28367
g25932 and pi0609 n28361_not ; n28368
g25933 and pi1155 n28367_not ; n28369
g25934 and n28368_not n28369 ; n28370
g25935 and pi0660 n28250_not ; n28371
g25936 and n28370_not n28371 ; n28372
g25937 nor n28366 n28372 ; n28373
g25938 and pi0785 n28373_not ; n28374
g25939 nor pi0785 n28361 ; n28375
g25940 nor n28374 n28375 ; n28376
g25941 nor pi0618 n28376 ; n28377
g25942 and pi0618 n28189 ; n28378
g25943 nor pi1154 n28378 ; n28379
g25944 and n28377_not n28379 ; n28380
g25945 nor pi0627 n28258 ; n28381
g25946 and n28380_not n28381 ; n28382
g25947 and pi0618_not n28189 ; n28383
g25948 and pi0618 n28376_not ; n28384
g25949 and pi1154 n28383_not ; n28385
g25950 and n28384_not n28385 ; n28386
g25951 and pi0627 n28262_not ; n28387
g25952 and n28386_not n28387 ; n28388
g25953 nor n28382 n28388 ; n28389
g25954 and pi0781 n28389_not ; n28390
g25955 nor pi0781 n28376 ; n28391
g25956 nor n28390 n28391 ; n28392
g25957 and pi0789_not n28392 ; n28393
g25958 and pi0619 n28192_not ; n28394
g25959 nor pi0619 n28392 ; n28395
g25960 nor pi1159 n28394 ; n28396
g25961 and n28395_not n28396 ; n28397
g25962 nor pi0648 n28270 ; n28398
g25963 and n28397_not n28398 ; n28399
g25964 nor pi0619 n28192 ; n28400
g25965 and pi0619 n28392_not ; n28401
g25966 and pi1159 n28400_not ; n28402
g25967 and n28401_not n28402 ; n28403
g25968 and pi0648 n28274_not ; n28404
g25969 and n28403_not n28404 ; n28405
g25970 and pi0789 n28399_not ; n28406
g25971 and n28405_not n28406 ; n28407
g25972 and n17970 n28393_not ; n28408
g25973 and n28407_not n28408 ; n28409
g25974 and n17871 n28194 ; n28410
g25975 nor pi0626 n28277 ; n28411
g25976 and pi0626 n28161_not ; n28412
g25977 and n16629 n28412_not ; n28413
g25978 and n28411_not n28413 ; n28414
g25979 and pi0626 n28277_not ; n28415
g25980 nor pi0626 n28161 ; n28416
g25981 and n16628 n28416_not ; n28417
g25982 and n28415_not n28417 ; n28418
g25983 nor n28410 n28414 ; n28419
g25984 and n28418_not n28419 ; n28420
g25985 and pi0788 n28420_not ; n28421
g25986 nor n20364 n28421 ; n28422
g25987 and n28409_not n28422 ; n28423
g25988 nor n28308 n28423 ; n28424
g25989 nor n20206 n28424 ; n28425
g25990 and n17802 n28212_not ; n28426
g25991 and n20559_not n28283 ; n28427
g25992 and n17801 n28216_not ; n28428
g25993 nor n28426 n28428 ; n28429
g25994 and n28427_not n28429 ; n28430
g25995 and pi0787 n28430_not ; n28431
g25996 and pi0644_not n28299 ; n28432
g25997 and pi0644 n28291 ; n28433
g25998 and pi0790 n28432_not ; n28434
g25999 and n28433_not n28434 ; n28435
g26000 nor n28425 n28431 ; n28436
g26001 and n28435_not n28436 ; n28437
g26002 nor n28302 n28437 ; n28438
g26003 nor po1038 n28438 ; n28439
g26004 nor pi0832 n28160 ; n28440
g26005 and n28439_not n28440 ; n28441
g26006 nor n28159 n28441 ; po0341
g26007 nor pi0185 n2926 ; n28443
g26008 and pi0701_not n16645 ; n28444
g26009 nor n28443 n28444 ; n28445
g26010 nor pi0778 n28445 ; n28446
g26011 and pi0625_not n28444 ; n28447
g26012 nor n28445 n28447 ; n28448
g26013 and pi1153 n28448_not ; n28449
g26014 nor pi1153 n28443 ; n28450
g26015 and n28447_not n28450 ; n28451
g26016 and pi0778 n28451_not ; n28452
g26017 and n28449_not n28452 ; n28453
g26018 nor n28446 n28453 ; n28454
g26019 nor n17845 n28454 ; n28455
g26020 and n17847_not n28455 ; n28456
g26021 and n17849_not n28456 ; n28457
g26022 and n17851_not n28457 ; n28458
g26023 and n17857_not n28458 ; n28459
g26024 and pi0647_not n28459 ; n28460
g26025 and pi0647 n28443 ; n28461
g26026 nor pi1157 n28461 ; n28462
g26027 and n28460_not n28462 ; n28463
g26028 and pi0630 n28463 ; n28464
g26029 and pi0751_not n17244 ; n28465
g26030 nor n28443 n28465 ; n28466
g26031 nor n17874 n28466 ; n28467
g26032 nor pi0785 n28467 ; n28468
g26033 and n17296 n28465 ; n28469
g26034 and n28467 n28469_not ; n28470
g26035 and pi1155 n28470_not ; n28471
g26036 nor pi1155 n28443 ; n28472
g26037 and n28469_not n28472 ; n28473
g26038 nor n28471 n28473 ; n28474
g26039 and pi0785 n28474_not ; n28475
g26040 nor n28468 n28475 ; n28476
g26041 nor pi0781 n28476 ; n28477
g26042 and n17889_not n28476 ; n28478
g26043 and pi1154 n28478_not ; n28479
g26044 and n17892_not n28476 ; n28480
g26045 nor pi1154 n28480 ; n28481
g26046 nor n28479 n28481 ; n28482
g26047 and pi0781 n28482_not ; n28483
g26048 nor n28477 n28483 ; n28484
g26049 nor pi0789 n28484 ; n28485
g26050 and n23078_not n28484 ; n28486
g26051 and pi1159 n28486_not ; n28487
g26052 and n23081_not n28484 ; n28488
g26053 nor pi1159 n28488 ; n28489
g26054 nor n28487 n28489 ; n28490
g26055 and pi0789 n28490_not ; n28491
g26056 nor n28485 n28491 ; n28492
g26057 and n17969_not n28492 ; n28493
g26058 and n17969 n28443 ; n28494
g26059 nor n28493 n28494 ; n28495
g26060 nor n17779 n28495 ; n28496
g26061 and n17779 n28443 ; n28497
g26062 nor n28496 n28497 ; n28498
g26063 and n20559_not n28498 ; n28499
g26064 and pi0647 n28459_not ; n28500
g26065 nor pi0647 n28443 ; n28501
g26066 nor n28500 n28501 ; n28502
g26067 and n17801 n28502_not ; n28503
g26068 nor n28464 n28503 ; n28504
g26069 and n28499_not n28504 ; n28505
g26070 and pi0787 n28505_not ; n28506
g26071 and n17871 n28457 ; n28507
g26072 nor pi0626 n28492 ; n28508
g26073 and pi0626 n28443_not ; n28509
g26074 and n16629 n28509_not ; n28510
g26075 and n28508_not n28510 ; n28511
g26076 and pi0626 n28492_not ; n28512
g26077 nor pi0626 n28443 ; n28513
g26078 and n16628 n28513_not ; n28514
g26079 and n28512_not n28514 ; n28515
g26080 nor n28507 n28511 ; n28516
g26081 and n28515_not n28516 ; n28517
g26082 and pi0788 n28517_not ; n28518
g26083 and pi0618 n28455 ; n28519
g26084 nor n17168 n28445 ; n28520
g26085 and pi0625 n28520 ; n28521
g26086 and n28466 n28520_not ; n28522
g26087 nor n28521 n28522 ; n28523
g26088 and n28450 n28523_not ; n28524
g26089 nor pi0608 n28449 ; n28525
g26090 and n28524_not n28525 ; n28526
g26091 and pi1153 n28466 ; n28527
g26092 and n28521_not n28527 ; n28528
g26093 and pi0608 n28451_not ; n28529
g26094 and n28528_not n28529 ; n28530
g26095 nor n28526 n28530 ; n28531
g26096 and pi0778 n28531_not ; n28532
g26097 nor pi0778 n28522 ; n28533
g26098 nor n28532 n28533 ; n28534
g26099 nor pi0609 n28534 ; n28535
g26100 and pi0609 n28454_not ; n28536
g26101 nor pi1155 n28536 ; n28537
g26102 and n28535_not n28537 ; n28538
g26103 nor pi0660 n28471 ; n28539
g26104 and n28538_not n28539 ; n28540
g26105 and pi0609 n28534_not ; n28541
g26106 nor pi0609 n28454 ; n28542
g26107 and pi1155 n28542_not ; n28543
g26108 and n28541_not n28543 ; n28544
g26109 and pi0660 n28473_not ; n28545
g26110 and n28544_not n28545 ; n28546
g26111 nor n28540 n28546 ; n28547
g26112 and pi0785 n28547_not ; n28548
g26113 nor pi0785 n28534 ; n28549
g26114 nor n28548 n28549 ; n28550
g26115 nor pi0618 n28550 ; n28551
g26116 nor pi1154 n28519 ; n28552
g26117 and n28551_not n28552 ; n28553
g26118 nor pi0627 n28479 ; n28554
g26119 and n28553_not n28554 ; n28555
g26120 and pi0618_not n28455 ; n28556
g26121 and pi0618 n28550_not ; n28557
g26122 and pi1154 n28556_not ; n28558
g26123 and n28557_not n28558 ; n28559
g26124 and pi0627 n28481_not ; n28560
g26125 and n28559_not n28560 ; n28561
g26126 nor n28555 n28561 ; n28562
g26127 and pi0781 n28562_not ; n28563
g26128 nor pi0781 n28550 ; n28564
g26129 nor n28563 n28564 ; n28565
g26130 and pi0789_not n28565 ; n28566
g26131 nor pi0619 n28565 ; n28567
g26132 and pi0619 n28456 ; n28568
g26133 nor pi1159 n28568 ; n28569
g26134 and n28567_not n28569 ; n28570
g26135 nor pi0648 n28487 ; n28571
g26136 and n28570_not n28571 ; n28572
g26137 and pi0619 n28565_not ; n28573
g26138 and pi0619_not n28456 ; n28574
g26139 and pi1159 n28574_not ; n28575
g26140 and n28573_not n28575 ; n28576
g26141 and pi0648 n28489_not ; n28577
g26142 and n28576_not n28577 ; n28578
g26143 and pi0789 n28572_not ; n28579
g26144 and n28578_not n28579 ; n28580
g26145 and n17970 n28566_not ; n28581
g26146 and n28580_not n28581 ; n28582
g26147 nor n28518 n28582 ; n28583
g26148 nor n20364 n28583 ; n28584
g26149 and n17854 n28495_not ; n28585
g26150 and n20851 n28458 ; n28586
g26151 nor n28585 n28586 ; n28587
g26152 nor pi0629 n28587 ; n28588
g26153 and n20855 n28458 ; n28589
g26154 and n17853 n28495_not ; n28590
g26155 nor n28589 n28590 ; n28591
g26156 and pi0629 n28591_not ; n28592
g26157 nor n28588 n28592 ; n28593
g26158 and pi0792 n28593_not ; n28594
g26159 nor n20206 n28594 ; n28595
g26160 and n28584_not n28595 ; n28596
g26161 nor n28506 n28596 ; n28597
g26162 and pi0790_not n28597 ; n28598
g26163 nor pi0787 n28459 ; n28599
g26164 and pi1157 n28502_not ; n28600
g26165 nor n28463 n28600 ; n28601
g26166 and pi0787 n28601_not ; n28602
g26167 nor n28599 n28602 ; n28603
g26168 and pi0644_not n28603 ; n28604
g26169 and pi0644 n28597 ; n28605
g26170 and pi0715 n28604_not ; n28606
g26171 and n28605_not n28606 ; n28607
g26172 nor n17804 n28498 ; n28608
g26173 and n17804 n28443 ; n28609
g26174 nor n28608 n28609 ; n28610
g26175 and pi0644 n28610_not ; n28611
g26176 and pi0644_not n28443 ; n28612
g26177 nor pi0715 n28612 ; n28613
g26178 and n28611_not n28613 ; n28614
g26179 and pi1160 n28614_not ; n28615
g26180 and n28607_not n28615 ; n28616
g26181 nor pi0644 n28610 ; n28617
g26182 and pi0644 n28443 ; n28618
g26183 and pi0715 n28618_not ; n28619
g26184 and n28617_not n28619 ; n28620
g26185 and pi0644 n28603 ; n28621
g26186 and pi0644_not n28597 ; n28622
g26187 nor pi0715 n28621 ; n28623
g26188 and n28622_not n28623 ; n28624
g26189 nor pi1160 n28620 ; n28625
g26190 and n28624_not n28625 ; n28626
g26191 nor n28616 n28626 ; n28627
g26192 and pi0790 n28627_not ; n28628
g26193 and pi0832 n28598_not ; n28629
g26194 and n28628_not n28629 ; n28630
g26195 and pi0185_not po1038 ; n28631
g26196 nor pi0185 n17059 ; n28632
g26197 and n16635 n28632_not ; n28633
g26198 and pi0701_not n2571 ; n28634
g26199 and n28632 n28634_not ; n28635
g26200 nor pi0185 n16641 ; n28636
g26201 and n16647 n28636_not ; n28637
g26202 and pi0185 n18076_not ; n28638
g26203 nor pi0038 n28638 ; n28639
g26204 and n2571 n28639_not ; n28640
g26205 and pi0185_not n18072 ; n28641
g26206 nor n28640 n28641 ; n28642
g26207 nor pi0701 n28637 ; n28643
g26208 and n28642_not n28643 ; n28644
g26209 nor n28635 n28644 ; n28645
g26210 and pi0778_not n28645 ; n28646
g26211 and pi0625_not n28632 ; n28647
g26212 and pi0625 n28645_not ; n28648
g26213 and pi1153 n28647_not ; n28649
g26214 and n28648_not n28649 ; n28650
g26215 and pi0625 n28632 ; n28651
g26216 nor pi0625 n28645 ; n28652
g26217 nor pi1153 n28651 ; n28653
g26218 and n28652_not n28653 ; n28654
g26219 nor n28650 n28654 ; n28655
g26220 and pi0778 n28655_not ; n28656
g26221 nor n28646 n28656 ; n28657
g26222 nor n17075 n28657 ; n28658
g26223 and n17075 n28632_not ; n28659
g26224 nor n28658 n28659 ; n28660
g26225 and n16639_not n28660 ; n28661
g26226 and n16639 n28632 ; n28662
g26227 nor n28661 n28662 ; n28663
g26228 and n16635_not n28663 ; n28664
g26229 nor n28633 n28664 ; n28665
g26230 and n16631_not n28665 ; n28666
g26231 and n16631 n28632 ; n28667
g26232 nor n28666 n28667 ; n28668
g26233 and pi0792_not n28668 ; n28669
g26234 and pi0628 n28668_not ; n28670
g26235 and pi0628_not n28632 ; n28671
g26236 and pi1156 n28671_not ; n28672
g26237 and n28670_not n28672 ; n28673
g26238 and pi0628 n28632 ; n28674
g26239 nor pi0628 n28668 ; n28675
g26240 nor pi1156 n28674 ; n28676
g26241 and n28675_not n28676 ; n28677
g26242 nor n28673 n28677 ; n28678
g26243 and pi0792 n28678_not ; n28679
g26244 nor n28669 n28679 ; n28680
g26245 nor pi0647 n28680 ; n28681
g26246 and pi0647 n28632_not ; n28682
g26247 nor n28681 n28682 ; n28683
g26248 and pi1157_not n28683 ; n28684
g26249 and pi0647 n28680_not ; n28685
g26250 nor pi0647 n28632 ; n28686
g26251 nor n28685 n28686 ; n28687
g26252 and pi1157 n28687 ; n28688
g26253 nor n28684 n28688 ; n28689
g26254 and pi0787 n28689_not ; n28690
g26255 and pi0787_not n28680 ; n28691
g26256 nor n28690 n28691 ; n28692
g26257 nor pi0644 n28692 ; n28693
g26258 and pi0715 n28693_not ; n28694
g26259 and pi0185 n2571_not ; n28695
g26260 and pi0185 pi0751 ; n28696
g26261 and pi0751 n17046 ; n28697
g26262 and pi0185 n17273 ; n28698
g26263 nor n28697 n28698 ; n28699
g26264 and pi0039 n28699_not ; n28700
g26265 and pi0185 n17233_not ; n28701
g26266 nor n21259 n28701 ; n28702
g26267 nor pi0039 n28702 ; n28703
g26268 nor pi0185 pi0751 ; n28704
g26269 and n17221 n28704 ; n28705
g26270 nor n28696 n28703 ; n28706
g26271 and n28705_not n28706 ; n28707
g26272 and n28700_not n28707 ; n28708
g26273 nor pi0038 n28708 ; n28709
g26274 and pi0751_not n17280 ; n28710
g26275 and pi0038 n28636_not ; n28711
g26276 and n28710_not n28711 ; n28712
g26277 nor n28709 n28712 ; n28713
g26278 and n2571 n28713_not ; n28714
g26279 nor n28695 n28714 ; n28715
g26280 nor n17117 n28715 ; n28716
g26281 and n17117 n28632_not ; n28717
g26282 nor n28716 n28717 ; n28718
g26283 nor pi0785 n28718 ; n28719
g26284 nor n17291 n28632 ; n28720
g26285 and pi0609 n28716 ; n28721
g26286 nor n28720 n28721 ; n28722
g26287 and pi1155 n28722_not ; n28723
g26288 nor n17296 n28632 ; n28724
g26289 and pi0609_not n28716 ; n28725
g26290 nor n28724 n28725 ; n28726
g26291 nor pi1155 n28726 ; n28727
g26292 nor n28723 n28727 ; n28728
g26293 and pi0785 n28728_not ; n28729
g26294 nor n28719 n28729 ; n28730
g26295 nor pi0781 n28730 ; n28731
g26296 and pi0618_not n28632 ; n28732
g26297 and pi0618 n28730 ; n28733
g26298 and pi1154 n28732_not ; n28734
g26299 and n28733_not n28734 ; n28735
g26300 and pi0618_not n28730 ; n28736
g26301 and pi0618 n28632 ; n28737
g26302 nor pi1154 n28737 ; n28738
g26303 and n28736_not n28738 ; n28739
g26304 nor n28735 n28739 ; n28740
g26305 and pi0781 n28740_not ; n28741
g26306 nor n28731 n28741 ; n28742
g26307 nor pi0789 n28742 ; n28743
g26308 and pi0619_not n28632 ; n28744
g26309 and pi0619 n28742 ; n28745
g26310 and pi1159 n28744_not ; n28746
g26311 and n28745_not n28746 ; n28747
g26312 and pi0619_not n28742 ; n28748
g26313 and pi0619 n28632 ; n28749
g26314 nor pi1159 n28749 ; n28750
g26315 and n28748_not n28750 ; n28751
g26316 nor n28747 n28751 ; n28752
g26317 and pi0789 n28752_not ; n28753
g26318 nor n28743 n28753 ; n28754
g26319 and n17969_not n28754 ; n28755
g26320 and n17969 n28632 ; n28756
g26321 nor n28755 n28756 ; n28757
g26322 nor n17779 n28757 ; n28758
g26323 and n17779 n28632 ; n28759
g26324 nor n28758 n28759 ; n28760
g26325 nor n17804 n28760 ; n28761
g26326 and n17804 n28632 ; n28762
g26327 nor n28761 n28762 ; n28763
g26328 and pi0644 n28763_not ; n28764
g26329 and pi0644_not n28632 ; n28765
g26330 nor pi0715 n28765 ; n28766
g26331 and n28764_not n28766 ; n28767
g26332 and pi1160 n28767_not ; n28768
g26333 and n28694_not n28768 ; n28769
g26334 and pi0644 n28692_not ; n28770
g26335 nor pi0715 n28770 ; n28771
g26336 nor pi0644 n28763 ; n28772
g26337 and pi0644 n28632 ; n28773
g26338 and pi0715 n28773_not ; n28774
g26339 and n28772_not n28774 ; n28775
g26340 nor pi1160 n28775 ; n28776
g26341 and n28771_not n28776 ; n28777
g26342 nor n28769 n28777 ; n28778
g26343 and pi0790 n28778_not ; n28779
g26344 and pi0629_not n28673 ; n28780
g26345 and n20570_not n28757 ; n28781
g26346 and pi0629 n28677 ; n28782
g26347 nor n28780 n28782 ; n28783
g26348 and n28781_not n28783 ; n28784
g26349 and pi0792 n28784_not ; n28785
g26350 and pi0609 n28657 ; n28786
g26351 and pi0185 n17625_not ; n28787
g26352 nor pi0185 n17612 ; n28788
g26353 and pi0751 n28787_not ; n28789
g26354 and n28788_not n28789 ; n28790
g26355 and pi0185_not n17629 ; n28791
g26356 and pi0185 n17631 ; n28792
g26357 nor pi0751 n28792 ; n28793
g26358 and n28791_not n28793 ; n28794
g26359 nor n28790 n28794 ; n28795
g26360 nor pi0039 n28795 ; n28796
g26361 and pi0185 n17605 ; n28797
g26362 nor pi0185 n17546 ; n28798
g26363 nor pi0751 n28798 ; n28799
g26364 and n28797_not n28799 ; n28800
g26365 and pi0185_not n17404 ; n28801
g26366 and pi0185 n17485 ; n28802
g26367 and pi0751 n28802_not ; n28803
g26368 and n28801_not n28803 ; n28804
g26369 and pi0039 n28800_not ; n28805
g26370 and n28804_not n28805 ; n28806
g26371 nor pi0038 n28796 ; n28807
g26372 and n28806_not n28807 ; n28808
g26373 nor n17469 n28465 ; n28809
g26374 and pi0185 n28809_not ; n28810
g26375 and n6284 n28810 ; n28811
g26376 nor pi0751 n17490 ; n28812
g26377 and n19471 n28812_not ; n28813
g26378 nor pi0185 n28813 ; n28814
g26379 and pi0038 n28811_not ; n28815
g26380 and n28814_not n28815 ; n28816
g26381 nor pi0701 n28816 ; n28817
g26382 and n28808_not n28817 ; n28818
g26383 and pi0701 n28713 ; n28819
g26384 and n2571 n28818_not ; n28820
g26385 and n28819_not n28820 ; n28821
g26386 nor n28695 n28821 ; n28822
g26387 and pi0625_not n28822 ; n28823
g26388 and pi0625 n28715 ; n28824
g26389 nor pi1153 n28824 ; n28825
g26390 and n28823_not n28825 ; n28826
g26391 nor pi0608 n28650 ; n28827
g26392 and n28826_not n28827 ; n28828
g26393 and pi0625_not n28715 ; n28829
g26394 and pi0625 n28822 ; n28830
g26395 and pi1153 n28829_not ; n28831
g26396 and n28830_not n28831 ; n28832
g26397 and pi0608 n28654_not ; n28833
g26398 and n28832_not n28833 ; n28834
g26399 nor n28828 n28834 ; n28835
g26400 and pi0778 n28835_not ; n28836
g26401 and pi0778_not n28822 ; n28837
g26402 nor n28836 n28837 ; n28838
g26403 nor pi0609 n28838 ; n28839
g26404 nor pi1155 n28786 ; n28840
g26405 and n28839_not n28840 ; n28841
g26406 nor pi0660 n28723 ; n28842
g26407 and n28841_not n28842 ; n28843
g26408 and pi0609_not n28657 ; n28844
g26409 and pi0609 n28838_not ; n28845
g26410 and pi1155 n28844_not ; n28846
g26411 and n28845_not n28846 ; n28847
g26412 and pi0660 n28727_not ; n28848
g26413 and n28847_not n28848 ; n28849
g26414 nor n28843 n28849 ; n28850
g26415 and pi0785 n28850_not ; n28851
g26416 nor pi0785 n28838 ; n28852
g26417 nor n28851 n28852 ; n28853
g26418 nor pi0618 n28853 ; n28854
g26419 and pi0618 n28660 ; n28855
g26420 nor pi1154 n28855 ; n28856
g26421 and n28854_not n28856 ; n28857
g26422 nor pi0627 n28735 ; n28858
g26423 and n28857_not n28858 ; n28859
g26424 and pi0618_not n28660 ; n28860
g26425 and pi0618 n28853_not ; n28861
g26426 and pi1154 n28860_not ; n28862
g26427 and n28861_not n28862 ; n28863
g26428 and pi0627 n28739_not ; n28864
g26429 and n28863_not n28864 ; n28865
g26430 nor n28859 n28865 ; n28866
g26431 and pi0781 n28866_not ; n28867
g26432 nor pi0781 n28853 ; n28868
g26433 nor n28867 n28868 ; n28869
g26434 and pi0789_not n28869 ; n28870
g26435 and pi0619 n28663_not ; n28871
g26436 nor pi0619 n28869 ; n28872
g26437 nor pi1159 n28871 ; n28873
g26438 and n28872_not n28873 ; n28874
g26439 nor pi0648 n28747 ; n28875
g26440 and n28874_not n28875 ; n28876
g26441 nor pi0619 n28663 ; n28877
g26442 and pi0619 n28869_not ; n28878
g26443 and pi1159 n28877_not ; n28879
g26444 and n28878_not n28879 ; n28880
g26445 and pi0648 n28751_not ; n28881
g26446 and n28880_not n28881 ; n28882
g26447 and pi0789 n28876_not ; n28883
g26448 and n28882_not n28883 ; n28884
g26449 and n17970 n28870_not ; n28885
g26450 and n28884_not n28885 ; n28886
g26451 and n17871 n28665 ; n28887
g26452 nor pi0626 n28754 ; n28888
g26453 and pi0626 n28632_not ; n28889
g26454 and n16629 n28889_not ; n28890
g26455 and n28888_not n28890 ; n28891
g26456 and pi0626 n28754_not ; n28892
g26457 nor pi0626 n28632 ; n28893
g26458 and n16628 n28893_not ; n28894
g26459 and n28892_not n28894 ; n28895
g26460 nor n28887 n28891 ; n28896
g26461 and n28895_not n28896 ; n28897
g26462 and pi0788 n28897_not ; n28898
g26463 nor n20364 n28898 ; n28899
g26464 and n28886_not n28899 ; n28900
g26465 nor n28785 n28900 ; n28901
g26466 nor n20206 n28901 ; n28902
g26467 and n17802 n28683_not ; n28903
g26468 and n20559_not n28760 ; n28904
g26469 and n17801 n28687_not ; n28905
g26470 nor n28903 n28905 ; n28906
g26471 and n28904_not n28906 ; n28907
g26472 and pi0787 n28907_not ; n28908
g26473 and pi0644_not n28776 ; n28909
g26474 and pi0644 n28768 ; n28910
g26475 and pi0790 n28909_not ; n28911
g26476 and n28910_not n28911 ; n28912
g26477 nor n28902 n28908 ; n28913
g26478 and n28912_not n28913 ; n28914
g26479 nor n28779 n28914 ; n28915
g26480 nor po1038 n28915 ; n28916
g26481 nor pi0832 n28631 ; n28917
g26482 and n28916_not n28917 ; n28918
g26483 nor n28630 n28918 ; po0342
g26484 nor pi0186 n17059 ; n28920
g26485 and n16635 n28920_not ; n28921
g26486 and pi0186 n2571_not ; n28922
g26487 nor pi0186 n17052 ; n28923
g26488 and pi0703_not n28923 ; n28924
g26489 nor pi0186 n16641 ; n28925
g26490 and n16647 n28925_not ; n28926
g26491 and pi0186_not n18072 ; n28927
g26492 and pi0186 n18076_not ; n28928
g26493 nor pi0038 n28928 ; n28929
g26494 and n28927_not n28929 ; n28930
g26495 and pi0703 n28926_not ; n28931
g26496 and n28930_not n28931 ; n28932
g26497 and n2571 n28924_not ; n28933
g26498 and n28932_not n28933 ; n28934
g26499 nor n28922 n28934 ; n28935
g26500 nor pi0778 n28935 ; n28936
g26501 and pi0625_not n28920 ; n28937
g26502 and pi0625 n28935 ; n28938
g26503 and pi1153 n28937_not ; n28939
g26504 and n28938_not n28939 ; n28940
g26505 and pi0625_not n28935 ; n28941
g26506 and pi0625 n28920 ; n28942
g26507 nor pi1153 n28942 ; n28943
g26508 and n28941_not n28943 ; n28944
g26509 nor n28940 n28944 ; n28945
g26510 and pi0778 n28945_not ; n28946
g26511 nor n28936 n28946 ; n28947
g26512 nor n17075 n28947 ; n28948
g26513 and n17075 n28920_not ; n28949
g26514 nor n28948 n28949 ; n28950
g26515 and n16639_not n28950 ; n28951
g26516 and n16639 n28920 ; n28952
g26517 nor n28951 n28952 ; n28953
g26518 and n16635_not n28953 ; n28954
g26519 nor n28921 n28954 ; n28955
g26520 and n16631_not n28955 ; n28956
g26521 and n16631 n28920 ; n28957
g26522 nor n28956 n28957 ; n28958
g26523 and pi0792_not n28958 ; n28959
g26524 and pi0628_not n28920 ; n28960
g26525 and pi0628 n28958_not ; n28961
g26526 and pi1156 n28960_not ; n28962
g26527 and n28961_not n28962 ; n28963
g26528 and pi0628 n28920 ; n28964
g26529 nor pi0628 n28958 ; n28965
g26530 nor pi1156 n28964 ; n28966
g26531 and n28965_not n28966 ; n28967
g26532 nor n28963 n28967 ; n28968
g26533 and pi0792 n28968_not ; n28969
g26534 nor n28959 n28969 ; n28970
g26535 nor pi0787 n28970 ; n28971
g26536 and pi0647_not n28920 ; n28972
g26537 and pi0647 n28970 ; n28973
g26538 and pi1157 n28972_not ; n28974
g26539 and n28973_not n28974 ; n28975
g26540 and pi0647_not n28970 ; n28976
g26541 and pi0647 n28920 ; n28977
g26542 nor pi1157 n28977 ; n28978
g26543 and n28976_not n28978 ; n28979
g26544 nor n28975 n28979 ; n28980
g26545 and pi0787 n28980_not ; n28981
g26546 nor n28971 n28981 ; n28982
g26547 and pi0644_not n28982 ; n28983
g26548 and pi0618_not n28920 ; n28984
g26549 and pi0752 n28923_not ; n28985
g26550 and pi0186 n19434_not ; n28986
g26551 nor pi0186 pi0752 ; n28987
g26552 and n19439 n28987 ; n28988
g26553 nor n28986 n28988 ; n28989
g26554 nor n19433 n28989 ; n28990
g26555 nor n28985 n28990 ; n28991
g26556 and n2571 n28991_not ; n28992
g26557 nor n28922 n28992 ; n28993
g26558 nor n17117 n28993 ; n28994
g26559 and n17117 n28920_not ; n28995
g26560 nor n28994 n28995 ; n28996
g26561 nor pi0785 n28996 ; n28997
g26562 nor n17291 n28920 ; n28998
g26563 and pi0609 n28994 ; n28999
g26564 nor n28998 n28999 ; n29000
g26565 and pi1155 n29000_not ; n29001
g26566 nor n17296 n28920 ; n29002
g26567 and pi0609_not n28994 ; n29003
g26568 nor n29002 n29003 ; n29004
g26569 nor pi1155 n29004 ; n29005
g26570 nor n29001 n29005 ; n29006
g26571 and pi0785 n29006_not ; n29007
g26572 nor n28997 n29007 ; n29008
g26573 and pi0618 n29008 ; n29009
g26574 and pi1154 n28984_not ; n29010
g26575 and n29009_not n29010 ; n29011
g26576 and pi0186 n19468 ; n29012
g26577 and pi0186_not n19477 ; n29013
g26578 and pi0752 n19470_not ; n29014
g26579 and n29012_not n29014 ; n29015
g26580 and n29013_not n29015 ; n29016
g26581 nor pi0186 n19488 ; n29017
g26582 and pi0186 n19496 ; n29018
g26583 nor pi0752 n29017 ; n29019
g26584 and n29018_not n29019 ; n29020
g26585 and pi0703 n29020_not ; n29021
g26586 and n29016_not n29021 ; n29022
g26587 and pi0703_not n28991 ; n29023
g26588 and n2571 n29022_not ; n29024
g26589 and n29023_not n29024 ; n29025
g26590 nor n28922 n29025 ; n29026
g26591 and pi0625_not n29026 ; n29027
g26592 and pi0625 n28993 ; n29028
g26593 nor pi1153 n29028 ; n29029
g26594 and n29027_not n29029 ; n29030
g26595 nor pi0608 n28940 ; n29031
g26596 and n29030_not n29031 ; n29032
g26597 and pi0625_not n28993 ; n29033
g26598 and pi0625 n29026 ; n29034
g26599 and pi1153 n29033_not ; n29035
g26600 and n29034_not n29035 ; n29036
g26601 and pi0608 n28944_not ; n29037
g26602 and n29036_not n29037 ; n29038
g26603 nor n29032 n29038 ; n29039
g26604 and pi0778 n29039_not ; n29040
g26605 and pi0778_not n29026 ; n29041
g26606 nor n29040 n29041 ; n29042
g26607 nor pi0609 n29042 ; n29043
g26608 and pi0609 n28947 ; n29044
g26609 nor pi1155 n29044 ; n29045
g26610 and n29043_not n29045 ; n29046
g26611 nor pi0660 n29001 ; n29047
g26612 and n29046_not n29047 ; n29048
g26613 and pi0609_not n28947 ; n29049
g26614 and pi0609 n29042_not ; n29050
g26615 and pi1155 n29049_not ; n29051
g26616 and n29050_not n29051 ; n29052
g26617 and pi0660 n29005_not ; n29053
g26618 and n29052_not n29053 ; n29054
g26619 nor n29048 n29054 ; n29055
g26620 and pi0785 n29055_not ; n29056
g26621 nor pi0785 n29042 ; n29057
g26622 nor n29056 n29057 ; n29058
g26623 nor pi0618 n29058 ; n29059
g26624 and pi0618 n28950 ; n29060
g26625 nor pi1154 n29060 ; n29061
g26626 and n29059_not n29061 ; n29062
g26627 nor pi0627 n29011 ; n29063
g26628 and n29062_not n29063 ; n29064
g26629 and pi0618_not n29008 ; n29065
g26630 and pi0618 n28920 ; n29066
g26631 nor pi1154 n29066 ; n29067
g26632 and n29065_not n29067 ; n29068
g26633 and pi0618_not n28950 ; n29069
g26634 and pi0618 n29058_not ; n29070
g26635 and pi1154 n29069_not ; n29071
g26636 and n29070_not n29071 ; n29072
g26637 and pi0627 n29068_not ; n29073
g26638 and n29072_not n29073 ; n29074
g26639 nor n29064 n29074 ; n29075
g26640 and pi0781 n29075_not ; n29076
g26641 nor pi0781 n29058 ; n29077
g26642 nor n29076 n29077 ; n29078
g26643 nor pi0619 n29078 ; n29079
g26644 and pi0619 n28953_not ; n29080
g26645 nor pi1159 n29080 ; n29081
g26646 and n29079_not n29081 ; n29082
g26647 and pi0619_not n28920 ; n29083
g26648 nor pi0781 n29008 ; n29084
g26649 nor n29011 n29068 ; n29085
g26650 and pi0781 n29085_not ; n29086
g26651 nor n29084 n29086 ; n29087
g26652 and pi0619 n29087 ; n29088
g26653 and pi1159 n29083_not ; n29089
g26654 and n29088_not n29089 ; n29090
g26655 nor pi0648 n29090 ; n29091
g26656 and n29082_not n29091 ; n29092
g26657 and pi0619 n29078_not ; n29093
g26658 nor pi0619 n28953 ; n29094
g26659 and pi1159 n29094_not ; n29095
g26660 and n29093_not n29095 ; n29096
g26661 and pi0619_not n29087 ; n29097
g26662 and pi0619 n28920 ; n29098
g26663 nor pi1159 n29098 ; n29099
g26664 and n29097_not n29099 ; n29100
g26665 and pi0648 n29100_not ; n29101
g26666 and n29096_not n29101 ; n29102
g26667 nor n29092 n29102 ; n29103
g26668 and pi0789 n29103_not ; n29104
g26669 nor pi0789 n29078 ; n29105
g26670 nor n29104 n29105 ; n29106
g26671 and pi0788_not n29106 ; n29107
g26672 and pi0626_not n29106 ; n29108
g26673 and pi0626 n28955_not ; n29109
g26674 nor pi0641 n29109 ; n29110
g26675 and n29108_not n29110 ; n29111
g26676 nor pi0789 n29087 ; n29112
g26677 nor n29090 n29100 ; n29113
g26678 and pi0789 n29113_not ; n29114
g26679 nor n29112 n29114 ; n29115
g26680 nor pi0626 n29115 ; n29116
g26681 and pi0626 n28920_not ; n29117
g26682 and pi0641 n29117_not ; n29118
g26683 and n29116_not n29118 ; n29119
g26684 nor pi1158 n29119 ; n29120
g26685 and n29111_not n29120 ; n29121
g26686 and pi0626 n29106 ; n29122
g26687 nor pi0626 n28955 ; n29123
g26688 and pi0641 n29123_not ; n29124
g26689 and n29122_not n29124 ; n29125
g26690 and pi0626 n29115_not ; n29126
g26691 nor pi0626 n28920 ; n29127
g26692 nor pi0641 n29127 ; n29128
g26693 and n29126_not n29128 ; n29129
g26694 and pi1158 n29129_not ; n29130
g26695 and n29125_not n29130 ; n29131
g26696 nor n29121 n29131 ; n29132
g26697 and pi0788 n29132_not ; n29133
g26698 nor n29107 n29133 ; n29134
g26699 and pi0628_not n29134 ; n29135
g26700 and n17969_not n29115 ; n29136
g26701 and n17969 n28920 ; n29137
g26702 nor n29136 n29137 ; n29138
g26703 and pi0628 n29138_not ; n29139
g26704 nor pi1156 n29139 ; n29140
g26705 and n29135_not n29140 ; n29141
g26706 nor pi0629 n28963 ; n29142
g26707 and n29141_not n29142 ; n29143
g26708 and pi0628 n29134 ; n29144
g26709 nor pi0628 n29138 ; n29145
g26710 and pi1156 n29145_not ; n29146
g26711 and n29144_not n29146 ; n29147
g26712 and pi0629 n28967_not ; n29148
g26713 and n29147_not n29148 ; n29149
g26714 nor n29143 n29149 ; n29150
g26715 and pi0792 n29150_not ; n29151
g26716 and pi0792_not n29134 ; n29152
g26717 nor n29151 n29152 ; n29153
g26718 nor pi0647 n29153 ; n29154
g26719 nor n17779 n29138 ; n29155
g26720 and n17779 n28920 ; n29156
g26721 nor n29155 n29156 ; n29157
g26722 and pi0647 n29157_not ; n29158
g26723 nor pi1157 n29158 ; n29159
g26724 and n29154_not n29159 ; n29160
g26725 nor pi0630 n28975 ; n29161
g26726 and n29160_not n29161 ; n29162
g26727 and pi0647 n29153_not ; n29163
g26728 nor pi0647 n29157 ; n29164
g26729 and pi1157 n29164_not ; n29165
g26730 and n29163_not n29165 ; n29166
g26731 and pi0630 n28979_not ; n29167
g26732 and n29166_not n29167 ; n29168
g26733 nor n29162 n29168 ; n29169
g26734 and pi0787 n29169_not ; n29170
g26735 nor pi0787 n29153 ; n29171
g26736 nor n29170 n29171 ; n29172
g26737 and pi0644 n29172_not ; n29173
g26738 and pi0715 n28983_not ; n29174
g26739 and n29173_not n29174 ; n29175
g26740 and n17804 n28920_not ; n29176
g26741 and n17804_not n29157 ; n29177
g26742 nor n29176 n29177 ; n29178
g26743 and pi0644 n29178 ; n29179
g26744 and pi0644_not n28920 ; n29180
g26745 nor pi0715 n29180 ; n29181
g26746 and n29179_not n29181 ; n29182
g26747 and pi1160 n29182_not ; n29183
g26748 and n29175_not n29183 ; n29184
g26749 nor pi0644 n29172 ; n29185
g26750 and pi0644 n28982 ; n29186
g26751 nor pi0715 n29186 ; n29187
g26752 and n29185_not n29187 ; n29188
g26753 and pi0644_not n29178 ; n29189
g26754 and pi0644 n28920 ; n29190
g26755 and pi0715 n29190_not ; n29191
g26756 and n29189_not n29191 ; n29192
g26757 nor pi1160 n29192 ; n29193
g26758 and n29188_not n29193 ; n29194
g26759 and pi0790 n29184_not ; n29195
g26760 and n29194_not n29195 ; n29196
g26761 and pi0790_not n29172 ; n29197
g26762 nor po1038 n29197 ; n29198
g26763 and n29196_not n29198 ; n29199
g26764 and pi0186_not po1038 ; n29200
g26765 nor pi0832 n29200 ; n29201
g26766 and n29199_not n29201 ; n29202
g26767 nor pi0186 n2926 ; n29203
g26768 and pi0703 n16645 ; n29204
g26769 nor n29203 n29204 ; n29205
g26770 and pi0778_not n29205 ; n29206
g26771 and pi0625_not n29204 ; n29207
g26772 nor n29205 n29207 ; n29208
g26773 and pi1153 n29208_not ; n29209
g26774 nor pi1153 n29203 ; n29210
g26775 and n29207_not n29210 ; n29211
g26776 nor n29209 n29211 ; n29212
g26777 and pi0778 n29212_not ; n29213
g26778 nor n29206 n29213 ; n29214
g26779 and n17845_not n29214 ; n29215
g26780 and n17847_not n29215 ; n29216
g26781 and n17849_not n29216 ; n29217
g26782 and n17851_not n29217 ; n29218
g26783 and n17857_not n29218 ; n29219
g26784 and pi0647_not n29219 ; n29220
g26785 and pi0647 n29203 ; n29221
g26786 nor pi1157 n29221 ; n29222
g26787 and n29220_not n29222 ; n29223
g26788 and pi0630 n29223 ; n29224
g26789 and pi0752_not n17244 ; n29225
g26790 nor n29203 n29225 ; n29226
g26791 nor n17874 n29226 ; n29227
g26792 nor pi0785 n29227 ; n29228
g26793 nor n17879 n29226 ; n29229
g26794 and pi1155 n29229_not ; n29230
g26795 and n17882_not n29227 ; n29231
g26796 nor pi1155 n29231 ; n29232
g26797 nor n29230 n29232 ; n29233
g26798 and pi0785 n29233_not ; n29234
g26799 nor n29228 n29234 ; n29235
g26800 nor pi0781 n29235 ; n29236
g26801 and n17889_not n29235 ; n29237
g26802 and pi1154 n29237_not ; n29238
g26803 and n17892_not n29235 ; n29239
g26804 nor pi1154 n29239 ; n29240
g26805 nor n29238 n29240 ; n29241
g26806 and pi0781 n29241_not ; n29242
g26807 nor n29236 n29242 ; n29243
g26808 nor pi0789 n29243 ; n29244
g26809 and pi0619_not n29203 ; n29245
g26810 and pi0619 n29243 ; n29246
g26811 and pi1159 n29245_not ; n29247
g26812 and n29246_not n29247 ; n29248
g26813 and pi0619_not n29243 ; n29249
g26814 and pi0619 n29203 ; n29250
g26815 nor pi1159 n29250 ; n29251
g26816 and n29249_not n29251 ; n29252
g26817 nor n29248 n29252 ; n29253
g26818 and pi0789 n29253_not ; n29254
g26819 nor n29244 n29254 ; n29255
g26820 and n17969_not n29255 ; n29256
g26821 and n17969 n29203 ; n29257
g26822 nor n29256 n29257 ; n29258
g26823 nor n17779 n29258 ; n29259
g26824 and n17779 n29203 ; n29260
g26825 nor n29259 n29260 ; n29261
g26826 and n20559_not n29261 ; n29262
g26827 and pi0647 n29219_not ; n29263
g26828 nor pi0647 n29203 ; n29264
g26829 nor n29263 n29264 ; n29265
g26830 and n17801 n29265_not ; n29266
g26831 nor n29224 n29266 ; n29267
g26832 and n29262_not n29267 ; n29268
g26833 and pi0787 n29268_not ; n29269
g26834 and n17871 n29217 ; n29270
g26835 nor pi0626 n29255 ; n29271
g26836 and pi0626 n29203_not ; n29272
g26837 and n16629 n29272_not ; n29273
g26838 and n29271_not n29273 ; n29274
g26839 and pi0626 n29255_not ; n29275
g26840 nor pi0626 n29203 ; n29276
g26841 and n16628 n29276_not ; n29277
g26842 and n29275_not n29277 ; n29278
g26843 nor n29270 n29274 ; n29279
g26844 and n29278_not n29279 ; n29280
g26845 and pi0788 n29280_not ; n29281
g26846 and pi0618 n29215 ; n29282
g26847 and pi0609 n29214 ; n29283
g26848 nor n17168 n29205 ; n29284
g26849 and pi0625 n29284 ; n29285
g26850 and n29226 n29284_not ; n29286
g26851 nor n29285 n29286 ; n29287
g26852 and n29210 n29287_not ; n29288
g26853 nor pi0608 n29209 ; n29289
g26854 and n29288_not n29289 ; n29290
g26855 and pi1153 n29226 ; n29291
g26856 and n29285_not n29291 ; n29292
g26857 and pi0608 n29211_not ; n29293
g26858 and n29292_not n29293 ; n29294
g26859 nor n29290 n29294 ; n29295
g26860 and pi0778 n29295_not ; n29296
g26861 nor pi0778 n29286 ; n29297
g26862 nor n29296 n29297 ; n29298
g26863 nor pi0609 n29298 ; n29299
g26864 nor pi1155 n29283 ; n29300
g26865 and n29299_not n29300 ; n29301
g26866 nor pi0660 n29230 ; n29302
g26867 and n29301_not n29302 ; n29303
g26868 and pi0609_not n29214 ; n29304
g26869 and pi0609 n29298_not ; n29305
g26870 and pi1155 n29304_not ; n29306
g26871 and n29305_not n29306 ; n29307
g26872 and pi0660 n29232_not ; n29308
g26873 and n29307_not n29308 ; n29309
g26874 nor n29303 n29309 ; n29310
g26875 and pi0785 n29310_not ; n29311
g26876 nor pi0785 n29298 ; n29312
g26877 nor n29311 n29312 ; n29313
g26878 nor pi0618 n29313 ; n29314
g26879 nor pi1154 n29282 ; n29315
g26880 and n29314_not n29315 ; n29316
g26881 nor pi0627 n29238 ; n29317
g26882 and n29316_not n29317 ; n29318
g26883 and pi0618_not n29215 ; n29319
g26884 and pi0618 n29313_not ; n29320
g26885 and pi1154 n29319_not ; n29321
g26886 and n29320_not n29321 ; n29322
g26887 and pi0627 n29240_not ; n29323
g26888 and n29322_not n29323 ; n29324
g26889 nor n29318 n29324 ; n29325
g26890 and pi0781 n29325_not ; n29326
g26891 nor pi0781 n29313 ; n29327
g26892 nor n29326 n29327 ; n29328
g26893 and pi0789_not n29328 ; n29329
g26894 nor pi0619 n29328 ; n29330
g26895 and pi0619 n29216 ; n29331
g26896 nor pi1159 n29331 ; n29332
g26897 and n29330_not n29332 ; n29333
g26898 nor pi0648 n29248 ; n29334
g26899 and n29333_not n29334 ; n29335
g26900 and pi0619 n29328_not ; n29336
g26901 and pi0619_not n29216 ; n29337
g26902 and pi1159 n29337_not ; n29338
g26903 and n29336_not n29338 ; n29339
g26904 and pi0648 n29252_not ; n29340
g26905 and n29339_not n29340 ; n29341
g26906 and pi0789 n29335_not ; n29342
g26907 and n29341_not n29342 ; n29343
g26908 and n17970 n29329_not ; n29344
g26909 and n29343_not n29344 ; n29345
g26910 nor n29281 n29345 ; n29346
g26911 nor n20364 n29346 ; n29347
g26912 and n17854 n29258_not ; n29348
g26913 and n20851 n29218 ; n29349
g26914 nor n29348 n29349 ; n29350
g26915 nor pi0629 n29350 ; n29351
g26916 and n20855 n29218 ; n29352
g26917 and n17853 n29258_not ; n29353
g26918 nor n29352 n29353 ; n29354
g26919 and pi0629 n29354_not ; n29355
g26920 nor n29351 n29355 ; n29356
g26921 and pi0792 n29356_not ; n29357
g26922 nor n20206 n29357 ; n29358
g26923 and n29347_not n29358 ; n29359
g26924 nor n29269 n29359 ; n29360
g26925 and pi0790_not n29360 ; n29361
g26926 nor pi0787 n29219 ; n29362
g26927 and pi1157 n29265_not ; n29363
g26928 nor n29223 n29363 ; n29364
g26929 and pi0787 n29364_not ; n29365
g26930 nor n29362 n29365 ; n29366
g26931 and pi0644_not n29366 ; n29367
g26932 and pi0644 n29360 ; n29368
g26933 and pi0715 n29367_not ; n29369
g26934 and n29368_not n29369 ; n29370
g26935 nor n17804 n29261 ; n29371
g26936 and n17804 n29203 ; n29372
g26937 nor n29371 n29372 ; n29373
g26938 and pi0644 n29373_not ; n29374
g26939 and pi0644_not n29203 ; n29375
g26940 nor pi0715 n29375 ; n29376
g26941 and n29374_not n29376 ; n29377
g26942 and pi1160 n29377_not ; n29378
g26943 and n29370_not n29378 ; n29379
g26944 nor pi0644 n29373 ; n29380
g26945 and pi0644 n29203 ; n29381
g26946 and pi0715 n29381_not ; n29382
g26947 and n29380_not n29382 ; n29383
g26948 and pi0644 n29366 ; n29384
g26949 and pi0644_not n29360 ; n29385
g26950 nor pi0715 n29384 ; n29386
g26951 and n29385_not n29386 ; n29387
g26952 nor pi1160 n29383 ; n29388
g26953 and n29387_not n29388 ; n29389
g26954 nor n29379 n29389 ; n29390
g26955 and pi0790 n29390_not ; n29391
g26956 and pi0832 n29361_not ; n29392
g26957 and n29391_not n29392 ; n29393
g26958 nor n29202 n29393 ; po0343
g26959 nor pi0187 n17059 ; n29395
g26960 and n16635 n29395_not ; n29396
g26961 and pi0187 n2571_not ; n29397
g26962 nor pi0187 pi0726 ; n29398
g26963 and n17052_not n29398 ; n29399
g26964 nor pi0187 n16641 ; n29400
g26965 and n16647 n29400_not ; n29401
g26966 and pi0187_not n18072 ; n29402
g26967 and pi0187 n18076_not ; n29403
g26968 nor pi0038 n29403 ; n29404
g26969 and n29402_not n29404 ; n29405
g26970 and pi0726 n29401_not ; n29406
g26971 and n29405_not n29406 ; n29407
g26972 and n2571 n29399_not ; n29408
g26973 and n29407_not n29408 ; n29409
g26974 nor n29397 n29409 ; n29410
g26975 nor pi0778 n29410 ; n29411
g26976 and pi0625_not n29395 ; n29412
g26977 and pi0625 n29410 ; n29413
g26978 and pi1153 n29412_not ; n29414
g26979 and n29413_not n29414 ; n29415
g26980 and pi0625_not n29410 ; n29416
g26981 and pi0625 n29395 ; n29417
g26982 nor pi1153 n29417 ; n29418
g26983 and n29416_not n29418 ; n29419
g26984 nor n29415 n29419 ; n29420
g26985 and pi0778 n29420_not ; n29421
g26986 nor n29411 n29421 ; n29422
g26987 nor n17075 n29422 ; n29423
g26988 and n17075 n29395_not ; n29424
g26989 nor n29423 n29424 ; n29425
g26990 and n16639_not n29425 ; n29426
g26991 and n16639 n29395 ; n29427
g26992 nor n29426 n29427 ; n29428
g26993 and n16635_not n29428 ; n29429
g26994 nor n29396 n29429 ; n29430
g26995 and n16631_not n29430 ; n29431
g26996 and n16631 n29395 ; n29432
g26997 nor n29431 n29432 ; n29433
g26998 and pi0792_not n29433 ; n29434
g26999 and pi0628_not n29395 ; n29435
g27000 and pi0628 n29433_not ; n29436
g27001 and pi1156 n29435_not ; n29437
g27002 and n29436_not n29437 ; n29438
g27003 and pi0628 n29395 ; n29439
g27004 nor pi0628 n29433 ; n29440
g27005 nor pi1156 n29439 ; n29441
g27006 and n29440_not n29441 ; n29442
g27007 nor n29438 n29442 ; n29443
g27008 and pi0792 n29443_not ; n29444
g27009 nor n29434 n29444 ; n29445
g27010 nor pi0787 n29445 ; n29446
g27011 and pi0647_not n29395 ; n29447
g27012 and pi0647 n29445 ; n29448
g27013 and pi1157 n29447_not ; n29449
g27014 and n29448_not n29449 ; n29450
g27015 and pi0647_not n29445 ; n29451
g27016 and pi0647 n29395 ; n29452
g27017 nor pi1157 n29452 ; n29453
g27018 and n29451_not n29453 ; n29454
g27019 nor n29450 n29454 ; n29455
g27020 and pi0787 n29455_not ; n29456
g27021 nor n29446 n29456 ; n29457
g27022 and pi0644_not n29457 ; n29458
g27023 and pi0618_not n29395 ; n29459
g27024 nor pi0770 n19439 ; n29460
g27025 nor n21012 n29460 ; n29461
g27026 nor pi0187 n29461 ; n29462
g27027 nor pi0187 n19433 ; n29463
g27028 nor pi0770 n29463 ; n29464
g27029 and n24447_not n29464 ; n29465
g27030 nor n29462 n29465 ; n29466
g27031 and n2571 n29466 ; n29467
g27032 nor n29397 n29467 ; n29468
g27033 nor n17117 n29468 ; n29469
g27034 and n17117 n29395_not ; n29470
g27035 nor n29469 n29470 ; n29471
g27036 nor pi0785 n29471 ; n29472
g27037 nor n17291 n29395 ; n29473
g27038 and pi0609 n29469 ; n29474
g27039 nor n29473 n29474 ; n29475
g27040 and pi1155 n29475_not ; n29476
g27041 nor n17296 n29395 ; n29477
g27042 and pi0609_not n29469 ; n29478
g27043 nor n29477 n29478 ; n29479
g27044 nor pi1155 n29479 ; n29480
g27045 nor n29476 n29480 ; n29481
g27046 and pi0785 n29481_not ; n29482
g27047 nor n29472 n29482 ; n29483
g27048 and pi0618 n29483 ; n29484
g27049 and pi1154 n29459_not ; n29485
g27050 and n29484_not n29485 ; n29486
g27051 and pi0187 n19468 ; n29487
g27052 and pi0187_not n19477 ; n29488
g27053 and pi0770 n19470_not ; n29489
g27054 and n29487_not n29489 ; n29490
g27055 and n29488_not n29490 ; n29491
g27056 nor pi0187 n19488 ; n29492
g27057 and pi0187 n19496 ; n29493
g27058 nor pi0770 n29492 ; n29494
g27059 and n29493_not n29494 ; n29495
g27060 and pi0726 n29495_not ; n29496
g27061 and n29491_not n29496 ; n29497
g27062 nor pi0726 n29466 ; n29498
g27063 and n2571 n29497_not ; n29499
g27064 and n29498_not n29499 ; n29500
g27065 nor n29397 n29500 ; n29501
g27066 and pi0625_not n29501 ; n29502
g27067 and pi0625 n29468 ; n29503
g27068 nor pi1153 n29503 ; n29504
g27069 and n29502_not n29504 ; n29505
g27070 nor pi0608 n29415 ; n29506
g27071 and n29505_not n29506 ; n29507
g27072 and pi0625_not n29468 ; n29508
g27073 and pi0625 n29501 ; n29509
g27074 and pi1153 n29508_not ; n29510
g27075 and n29509_not n29510 ; n29511
g27076 and pi0608 n29419_not ; n29512
g27077 and n29511_not n29512 ; n29513
g27078 nor n29507 n29513 ; n29514
g27079 and pi0778 n29514_not ; n29515
g27080 and pi0778_not n29501 ; n29516
g27081 nor n29515 n29516 ; n29517
g27082 nor pi0609 n29517 ; n29518
g27083 and pi0609 n29422 ; n29519
g27084 nor pi1155 n29519 ; n29520
g27085 and n29518_not n29520 ; n29521
g27086 nor pi0660 n29476 ; n29522
g27087 and n29521_not n29522 ; n29523
g27088 and pi0609_not n29422 ; n29524
g27089 and pi0609 n29517_not ; n29525
g27090 and pi1155 n29524_not ; n29526
g27091 and n29525_not n29526 ; n29527
g27092 and pi0660 n29480_not ; n29528
g27093 and n29527_not n29528 ; n29529
g27094 nor n29523 n29529 ; n29530
g27095 and pi0785 n29530_not ; n29531
g27096 nor pi0785 n29517 ; n29532
g27097 nor n29531 n29532 ; n29533
g27098 nor pi0618 n29533 ; n29534
g27099 and pi0618 n29425 ; n29535
g27100 nor pi1154 n29535 ; n29536
g27101 and n29534_not n29536 ; n29537
g27102 nor pi0627 n29486 ; n29538
g27103 and n29537_not n29538 ; n29539
g27104 and pi0618_not n29483 ; n29540
g27105 and pi0618 n29395 ; n29541
g27106 nor pi1154 n29541 ; n29542
g27107 and n29540_not n29542 ; n29543
g27108 and pi0618_not n29425 ; n29544
g27109 and pi0618 n29533_not ; n29545
g27110 and pi1154 n29544_not ; n29546
g27111 and n29545_not n29546 ; n29547
g27112 and pi0627 n29543_not ; n29548
g27113 and n29547_not n29548 ; n29549
g27114 nor n29539 n29549 ; n29550
g27115 and pi0781 n29550_not ; n29551
g27116 nor pi0781 n29533 ; n29552
g27117 nor n29551 n29552 ; n29553
g27118 nor pi0619 n29553 ; n29554
g27119 and pi0619 n29428_not ; n29555
g27120 nor pi1159 n29555 ; n29556
g27121 and n29554_not n29556 ; n29557
g27122 and pi0619_not n29395 ; n29558
g27123 nor pi0781 n29483 ; n29559
g27124 nor n29486 n29543 ; n29560
g27125 and pi0781 n29560_not ; n29561
g27126 nor n29559 n29561 ; n29562
g27127 and pi0619 n29562 ; n29563
g27128 and pi1159 n29558_not ; n29564
g27129 and n29563_not n29564 ; n29565
g27130 nor pi0648 n29565 ; n29566
g27131 and n29557_not n29566 ; n29567
g27132 and pi0619 n29553_not ; n29568
g27133 nor pi0619 n29428 ; n29569
g27134 and pi1159 n29569_not ; n29570
g27135 and n29568_not n29570 ; n29571
g27136 and pi0619_not n29562 ; n29572
g27137 and pi0619 n29395 ; n29573
g27138 nor pi1159 n29573 ; n29574
g27139 and n29572_not n29574 ; n29575
g27140 and pi0648 n29575_not ; n29576
g27141 and n29571_not n29576 ; n29577
g27142 nor n29567 n29577 ; n29578
g27143 and pi0789 n29578_not ; n29579
g27144 nor pi0789 n29553 ; n29580
g27145 nor n29579 n29580 ; n29581
g27146 and pi0788_not n29581 ; n29582
g27147 and pi0626_not n29581 ; n29583
g27148 and pi0626 n29430_not ; n29584
g27149 nor pi0641 n29584 ; n29585
g27150 and n29583_not n29585 ; n29586
g27151 nor pi0789 n29562 ; n29587
g27152 nor n29565 n29575 ; n29588
g27153 and pi0789 n29588_not ; n29589
g27154 nor n29587 n29589 ; n29590
g27155 nor pi0626 n29590 ; n29591
g27156 and pi0626 n29395_not ; n29592
g27157 and pi0641 n29592_not ; n29593
g27158 and n29591_not n29593 ; n29594
g27159 nor pi1158 n29594 ; n29595
g27160 and n29586_not n29595 ; n29596
g27161 and pi0626 n29581 ; n29597
g27162 nor pi0626 n29430 ; n29598
g27163 and pi0641 n29598_not ; n29599
g27164 and n29597_not n29599 ; n29600
g27165 and pi0626 n29590_not ; n29601
g27166 nor pi0626 n29395 ; n29602
g27167 nor pi0641 n29602 ; n29603
g27168 and n29601_not n29603 ; n29604
g27169 and pi1158 n29604_not ; n29605
g27170 and n29600_not n29605 ; n29606
g27171 nor n29596 n29606 ; n29607
g27172 and pi0788 n29607_not ; n29608
g27173 nor n29582 n29608 ; n29609
g27174 and pi0628_not n29609 ; n29610
g27175 and n17969_not n29590 ; n29611
g27176 and n17969 n29395 ; n29612
g27177 nor n29611 n29612 ; n29613
g27178 and pi0628 n29613_not ; n29614
g27179 nor pi1156 n29614 ; n29615
g27180 and n29610_not n29615 ; n29616
g27181 nor pi0629 n29438 ; n29617
g27182 and n29616_not n29617 ; n29618
g27183 and pi0628 n29609 ; n29619
g27184 nor pi0628 n29613 ; n29620
g27185 and pi1156 n29620_not ; n29621
g27186 and n29619_not n29621 ; n29622
g27187 and pi0629 n29442_not ; n29623
g27188 and n29622_not n29623 ; n29624
g27189 nor n29618 n29624 ; n29625
g27190 and pi0792 n29625_not ; n29626
g27191 and pi0792_not n29609 ; n29627
g27192 nor n29626 n29627 ; n29628
g27193 nor pi0647 n29628 ; n29629
g27194 nor n17779 n29613 ; n29630
g27195 and n17779 n29395 ; n29631
g27196 nor n29630 n29631 ; n29632
g27197 and pi0647 n29632_not ; n29633
g27198 nor pi1157 n29633 ; n29634
g27199 and n29629_not n29634 ; n29635
g27200 nor pi0630 n29450 ; n29636
g27201 and n29635_not n29636 ; n29637
g27202 and pi0647 n29628_not ; n29638
g27203 nor pi0647 n29632 ; n29639
g27204 and pi1157 n29639_not ; n29640
g27205 and n29638_not n29640 ; n29641
g27206 and pi0630 n29454_not ; n29642
g27207 and n29641_not n29642 ; n29643
g27208 nor n29637 n29643 ; n29644
g27209 and pi0787 n29644_not ; n29645
g27210 nor pi0787 n29628 ; n29646
g27211 nor n29645 n29646 ; n29647
g27212 and pi0644 n29647_not ; n29648
g27213 and pi0715 n29458_not ; n29649
g27214 and n29648_not n29649 ; n29650
g27215 and n17804 n29395_not ; n29651
g27216 and n17804_not n29632 ; n29652
g27217 nor n29651 n29652 ; n29653
g27218 and pi0644 n29653 ; n29654
g27219 and pi0644_not n29395 ; n29655
g27220 nor pi0715 n29655 ; n29656
g27221 and n29654_not n29656 ; n29657
g27222 and pi1160 n29657_not ; n29658
g27223 and n29650_not n29658 ; n29659
g27224 nor pi0644 n29647 ; n29660
g27225 and pi0644 n29457 ; n29661
g27226 nor pi0715 n29661 ; n29662
g27227 and n29660_not n29662 ; n29663
g27228 and pi0644_not n29653 ; n29664
g27229 and pi0644 n29395 ; n29665
g27230 and pi0715 n29665_not ; n29666
g27231 and n29664_not n29666 ; n29667
g27232 nor pi1160 n29667 ; n29668
g27233 and n29663_not n29668 ; n29669
g27234 and pi0790 n29659_not ; n29670
g27235 and n29669_not n29670 ; n29671
g27236 and pi0790_not n29647 ; n29672
g27237 nor po1038 n29672 ; n29673
g27238 and n29671_not n29673 ; n29674
g27239 and pi0187_not po1038 ; n29675
g27240 nor pi0832 n29675 ; n29676
g27241 and n29674_not n29676 ; n29677
g27242 nor pi0187 n2926 ; n29678
g27243 and pi0726 n16645 ; n29679
g27244 nor n29678 n29679 ; n29680
g27245 and pi0778_not n29680 ; n29681
g27246 and pi0625_not n29679 ; n29682
g27247 nor n29680 n29682 ; n29683
g27248 and pi1153 n29683_not ; n29684
g27249 nor pi1153 n29678 ; n29685
g27250 and n29682_not n29685 ; n29686
g27251 nor n29684 n29686 ; n29687
g27252 and pi0778 n29687_not ; n29688
g27253 nor n29681 n29688 ; n29689
g27254 and n17845_not n29689 ; n29690
g27255 and n17847_not n29690 ; n29691
g27256 and n17849_not n29691 ; n29692
g27257 and n17851_not n29692 ; n29693
g27258 and n17857_not n29693 ; n29694
g27259 and pi0647_not n29694 ; n29695
g27260 and pi0647 n29678 ; n29696
g27261 nor pi1157 n29696 ; n29697
g27262 and n29695_not n29697 ; n29698
g27263 and pi0630 n29698 ; n29699
g27264 and pi0770_not n17244 ; n29700
g27265 nor n29678 n29700 ; n29701
g27266 nor n17874 n29701 ; n29702
g27267 nor pi0785 n29702 ; n29703
g27268 nor n17879 n29701 ; n29704
g27269 and pi1155 n29704_not ; n29705
g27270 and n17882_not n29702 ; n29706
g27271 nor pi1155 n29706 ; n29707
g27272 nor n29705 n29707 ; n29708
g27273 and pi0785 n29708_not ; n29709
g27274 nor n29703 n29709 ; n29710
g27275 nor pi0781 n29710 ; n29711
g27276 and n17889_not n29710 ; n29712
g27277 and pi1154 n29712_not ; n29713
g27278 and n17892_not n29710 ; n29714
g27279 nor pi1154 n29714 ; n29715
g27280 nor n29713 n29715 ; n29716
g27281 and pi0781 n29716_not ; n29717
g27282 nor n29711 n29717 ; n29718
g27283 nor pi0789 n29718 ; n29719
g27284 and pi0619_not n29678 ; n29720
g27285 and pi0619 n29718 ; n29721
g27286 and pi1159 n29720_not ; n29722
g27287 and n29721_not n29722 ; n29723
g27288 and pi0619_not n29718 ; n29724
g27289 and pi0619 n29678 ; n29725
g27290 nor pi1159 n29725 ; n29726
g27291 and n29724_not n29726 ; n29727
g27292 nor n29723 n29727 ; n29728
g27293 and pi0789 n29728_not ; n29729
g27294 nor n29719 n29729 ; n29730
g27295 and n17969_not n29730 ; n29731
g27296 and n17969 n29678 ; n29732
g27297 nor n29731 n29732 ; n29733
g27298 nor n17779 n29733 ; n29734
g27299 and n17779 n29678 ; n29735
g27300 nor n29734 n29735 ; n29736
g27301 and n20559_not n29736 ; n29737
g27302 and pi0647 n29694_not ; n29738
g27303 nor pi0647 n29678 ; n29739
g27304 nor n29738 n29739 ; n29740
g27305 and n17801 n29740_not ; n29741
g27306 nor n29699 n29741 ; n29742
g27307 and n29737_not n29742 ; n29743
g27308 and pi0787 n29743_not ; n29744
g27309 and n17871 n29692 ; n29745
g27310 nor pi0626 n29730 ; n29746
g27311 and pi0626 n29678_not ; n29747
g27312 and n16629 n29747_not ; n29748
g27313 and n29746_not n29748 ; n29749
g27314 and pi0626 n29730_not ; n29750
g27315 nor pi0626 n29678 ; n29751
g27316 and n16628 n29751_not ; n29752
g27317 and n29750_not n29752 ; n29753
g27318 nor n29745 n29749 ; n29754
g27319 and n29753_not n29754 ; n29755
g27320 and pi0788 n29755_not ; n29756
g27321 and pi0618 n29690 ; n29757
g27322 and pi0609 n29689 ; n29758
g27323 nor n17168 n29680 ; n29759
g27324 and pi0625 n29759 ; n29760
g27325 and n29701 n29759_not ; n29761
g27326 nor n29760 n29761 ; n29762
g27327 and n29685 n29762_not ; n29763
g27328 nor pi0608 n29684 ; n29764
g27329 and n29763_not n29764 ; n29765
g27330 and pi1153 n29701 ; n29766
g27331 and n29760_not n29766 ; n29767
g27332 and pi0608 n29686_not ; n29768
g27333 and n29767_not n29768 ; n29769
g27334 nor n29765 n29769 ; n29770
g27335 and pi0778 n29770_not ; n29771
g27336 nor pi0778 n29761 ; n29772
g27337 nor n29771 n29772 ; n29773
g27338 nor pi0609 n29773 ; n29774
g27339 nor pi1155 n29758 ; n29775
g27340 and n29774_not n29775 ; n29776
g27341 nor pi0660 n29705 ; n29777
g27342 and n29776_not n29777 ; n29778
g27343 and pi0609_not n29689 ; n29779
g27344 and pi0609 n29773_not ; n29780
g27345 and pi1155 n29779_not ; n29781
g27346 and n29780_not n29781 ; n29782
g27347 and pi0660 n29707_not ; n29783
g27348 and n29782_not n29783 ; n29784
g27349 nor n29778 n29784 ; n29785
g27350 and pi0785 n29785_not ; n29786
g27351 nor pi0785 n29773 ; n29787
g27352 nor n29786 n29787 ; n29788
g27353 nor pi0618 n29788 ; n29789
g27354 nor pi1154 n29757 ; n29790
g27355 and n29789_not n29790 ; n29791
g27356 nor pi0627 n29713 ; n29792
g27357 and n29791_not n29792 ; n29793
g27358 and pi0618_not n29690 ; n29794
g27359 and pi0618 n29788_not ; n29795
g27360 and pi1154 n29794_not ; n29796
g27361 and n29795_not n29796 ; n29797
g27362 and pi0627 n29715_not ; n29798
g27363 and n29797_not n29798 ; n29799
g27364 nor n29793 n29799 ; n29800
g27365 and pi0781 n29800_not ; n29801
g27366 nor pi0781 n29788 ; n29802
g27367 nor n29801 n29802 ; n29803
g27368 and pi0789_not n29803 ; n29804
g27369 nor pi0619 n29803 ; n29805
g27370 and pi0619 n29691 ; n29806
g27371 nor pi1159 n29806 ; n29807
g27372 and n29805_not n29807 ; n29808
g27373 nor pi0648 n29723 ; n29809
g27374 and n29808_not n29809 ; n29810
g27375 and pi0619 n29803_not ; n29811
g27376 and pi0619_not n29691 ; n29812
g27377 and pi1159 n29812_not ; n29813
g27378 and n29811_not n29813 ; n29814
g27379 and pi0648 n29727_not ; n29815
g27380 and n29814_not n29815 ; n29816
g27381 and pi0789 n29810_not ; n29817
g27382 and n29816_not n29817 ; n29818
g27383 and n17970 n29804_not ; n29819
g27384 and n29818_not n29819 ; n29820
g27385 nor n29756 n29820 ; n29821
g27386 nor n20364 n29821 ; n29822
g27387 and n17854 n29733_not ; n29823
g27388 and n20851 n29693 ; n29824
g27389 nor n29823 n29824 ; n29825
g27390 nor pi0629 n29825 ; n29826
g27391 and n20855 n29693 ; n29827
g27392 and n17853 n29733_not ; n29828
g27393 nor n29827 n29828 ; n29829
g27394 and pi0629 n29829_not ; n29830
g27395 nor n29826 n29830 ; n29831
g27396 and pi0792 n29831_not ; n29832
g27397 nor n20206 n29832 ; n29833
g27398 and n29822_not n29833 ; n29834
g27399 nor n29744 n29834 ; n29835
g27400 and pi0790_not n29835 ; n29836
g27401 nor pi0787 n29694 ; n29837
g27402 and pi1157 n29740_not ; n29838
g27403 nor n29698 n29838 ; n29839
g27404 and pi0787 n29839_not ; n29840
g27405 nor n29837 n29840 ; n29841
g27406 and pi0644_not n29841 ; n29842
g27407 and pi0644 n29835 ; n29843
g27408 and pi0715 n29842_not ; n29844
g27409 and n29843_not n29844 ; n29845
g27410 nor n17804 n29736 ; n29846
g27411 and n17804 n29678 ; n29847
g27412 nor n29846 n29847 ; n29848
g27413 and pi0644 n29848_not ; n29849
g27414 and pi0644_not n29678 ; n29850
g27415 nor pi0715 n29850 ; n29851
g27416 and n29849_not n29851 ; n29852
g27417 and pi1160 n29852_not ; n29853
g27418 and n29845_not n29853 ; n29854
g27419 nor pi0644 n29848 ; n29855
g27420 and pi0644 n29678 ; n29856
g27421 and pi0715 n29856_not ; n29857
g27422 and n29855_not n29857 ; n29858
g27423 and pi0644 n29841 ; n29859
g27424 and pi0644_not n29835 ; n29860
g27425 nor pi0715 n29859 ; n29861
g27426 and n29860_not n29861 ; n29862
g27427 nor pi1160 n29858 ; n29863
g27428 and n29862_not n29863 ; n29864
g27429 nor n29854 n29864 ; n29865
g27430 and pi0790 n29865_not ; n29866
g27431 and pi0832 n29836_not ; n29867
g27432 and n29866_not n29867 ; n29868
g27433 nor n29677 n29868 ; po0344
g27434 nor pi0188 n17059 ; n29870
g27435 and n16635 n29870_not ; n29871
g27436 and pi0188 n2571_not ; n29872
g27437 nor pi0188 pi0705 ; n29873
g27438 and n17052_not n29873 ; n29874
g27439 nor pi0188 n16641 ; n29875
g27440 and n16647 n29875_not ; n29876
g27441 and pi0188_not n18072 ; n29877
g27442 and pi0188 n18076_not ; n29878
g27443 nor pi0038 n29878 ; n29879
g27444 and n29877_not n29879 ; n29880
g27445 and pi0705 n29876_not ; n29881
g27446 and n29880_not n29881 ; n29882
g27447 and n2571 n29874_not ; n29883
g27448 and n29882_not n29883 ; n29884
g27449 nor n29872 n29884 ; n29885
g27450 nor pi0778 n29885 ; n29886
g27451 and pi0625_not n29870 ; n29887
g27452 and pi0625 n29885 ; n29888
g27453 and pi1153 n29887_not ; n29889
g27454 and n29888_not n29889 ; n29890
g27455 and pi0625_not n29885 ; n29891
g27456 and pi0625 n29870 ; n29892
g27457 nor pi1153 n29892 ; n29893
g27458 and n29891_not n29893 ; n29894
g27459 nor n29890 n29894 ; n29895
g27460 and pi0778 n29895_not ; n29896
g27461 nor n29886 n29896 ; n29897
g27462 nor n17075 n29897 ; n29898
g27463 and n17075 n29870_not ; n29899
g27464 nor n29898 n29899 ; n29900
g27465 and n16639_not n29900 ; n29901
g27466 and n16639 n29870 ; n29902
g27467 nor n29901 n29902 ; n29903
g27468 and n16635_not n29903 ; n29904
g27469 nor n29871 n29904 ; n29905
g27470 and n16631_not n29905 ; n29906
g27471 and n16631 n29870 ; n29907
g27472 nor n29906 n29907 ; n29908
g27473 and pi0792_not n29908 ; n29909
g27474 and pi0628_not n29870 ; n29910
g27475 and pi0628 n29908_not ; n29911
g27476 and pi1156 n29910_not ; n29912
g27477 and n29911_not n29912 ; n29913
g27478 and pi0628 n29870 ; n29914
g27479 nor pi0628 n29908 ; n29915
g27480 nor pi1156 n29914 ; n29916
g27481 and n29915_not n29916 ; n29917
g27482 nor n29913 n29917 ; n29918
g27483 and pi0792 n29918_not ; n29919
g27484 nor n29909 n29919 ; n29920
g27485 nor pi0787 n29920 ; n29921
g27486 and pi0647_not n29870 ; n29922
g27487 and pi0647 n29920 ; n29923
g27488 and pi1157 n29922_not ; n29924
g27489 and n29923_not n29924 ; n29925
g27490 and pi0647_not n29920 ; n29926
g27491 and pi0647 n29870 ; n29927
g27492 nor pi1157 n29927 ; n29928
g27493 and n29926_not n29928 ; n29929
g27494 nor n29925 n29929 ; n29930
g27495 and pi0787 n29930_not ; n29931
g27496 nor n29921 n29931 ; n29932
g27497 and pi0644_not n29932 ; n29933
g27498 and pi0618_not n29870 ; n29934
g27499 nor pi0768 n19439 ; n29935
g27500 nor n22313 n29935 ; n29936
g27501 nor pi0188 n29936 ; n29937
g27502 nor pi0188 n19433 ; n29938
g27503 nor pi0768 n29938 ; n29939
g27504 and n24447_not n29939 ; n29940
g27505 nor n29937 n29940 ; n29941
g27506 and n2571 n29941 ; n29942
g27507 nor n29872 n29942 ; n29943
g27508 nor n17117 n29943 ; n29944
g27509 and n17117 n29870_not ; n29945
g27510 nor n29944 n29945 ; n29946
g27511 nor pi0785 n29946 ; n29947
g27512 nor n17291 n29870 ; n29948
g27513 and pi0609 n29944 ; n29949
g27514 nor n29948 n29949 ; n29950
g27515 and pi1155 n29950_not ; n29951
g27516 nor n17296 n29870 ; n29952
g27517 and pi0609_not n29944 ; n29953
g27518 nor n29952 n29953 ; n29954
g27519 nor pi1155 n29954 ; n29955
g27520 nor n29951 n29955 ; n29956
g27521 and pi0785 n29956_not ; n29957
g27522 nor n29947 n29957 ; n29958
g27523 and pi0618 n29958 ; n29959
g27524 and pi1154 n29934_not ; n29960
g27525 and n29959_not n29960 ; n29961
g27526 and pi0188 n19468 ; n29962
g27527 and pi0188_not n19477 ; n29963
g27528 and pi0768 n19470_not ; n29964
g27529 and n29962_not n29964 ; n29965
g27530 and n29963_not n29965 ; n29966
g27531 nor pi0188 n19488 ; n29967
g27532 and pi0188 n19496 ; n29968
g27533 nor pi0768 n29967 ; n29969
g27534 and n29968_not n29969 ; n29970
g27535 and pi0705 n29970_not ; n29971
g27536 and n29966_not n29971 ; n29972
g27537 nor pi0705 n29941 ; n29973
g27538 and n2571 n29972_not ; n29974
g27539 and n29973_not n29974 ; n29975
g27540 nor n29872 n29975 ; n29976
g27541 and pi0625_not n29976 ; n29977
g27542 and pi0625 n29943 ; n29978
g27543 nor pi1153 n29978 ; n29979
g27544 and n29977_not n29979 ; n29980
g27545 nor pi0608 n29890 ; n29981
g27546 and n29980_not n29981 ; n29982
g27547 and pi0625_not n29943 ; n29983
g27548 and pi0625 n29976 ; n29984
g27549 and pi1153 n29983_not ; n29985
g27550 and n29984_not n29985 ; n29986
g27551 and pi0608 n29894_not ; n29987
g27552 and n29986_not n29987 ; n29988
g27553 nor n29982 n29988 ; n29989
g27554 and pi0778 n29989_not ; n29990
g27555 and pi0778_not n29976 ; n29991
g27556 nor n29990 n29991 ; n29992
g27557 nor pi0609 n29992 ; n29993
g27558 and pi0609 n29897 ; n29994
g27559 nor pi1155 n29994 ; n29995
g27560 and n29993_not n29995 ; n29996
g27561 nor pi0660 n29951 ; n29997
g27562 and n29996_not n29997 ; n29998
g27563 and pi0609_not n29897 ; n29999
g27564 and pi0609 n29992_not ; n30000
g27565 and pi1155 n29999_not ; n30001
g27566 and n30000_not n30001 ; n30002
g27567 and pi0660 n29955_not ; n30003
g27568 and n30002_not n30003 ; n30004
g27569 nor n29998 n30004 ; n30005
g27570 and pi0785 n30005_not ; n30006
g27571 nor pi0785 n29992 ; n30007
g27572 nor n30006 n30007 ; n30008
g27573 nor pi0618 n30008 ; n30009
g27574 and pi0618 n29900 ; n30010
g27575 nor pi1154 n30010 ; n30011
g27576 and n30009_not n30011 ; n30012
g27577 nor pi0627 n29961 ; n30013
g27578 and n30012_not n30013 ; n30014
g27579 and pi0618_not n29958 ; n30015
g27580 and pi0618 n29870 ; n30016
g27581 nor pi1154 n30016 ; n30017
g27582 and n30015_not n30017 ; n30018
g27583 and pi0618_not n29900 ; n30019
g27584 and pi0618 n30008_not ; n30020
g27585 and pi1154 n30019_not ; n30021
g27586 and n30020_not n30021 ; n30022
g27587 and pi0627 n30018_not ; n30023
g27588 and n30022_not n30023 ; n30024
g27589 nor n30014 n30024 ; n30025
g27590 and pi0781 n30025_not ; n30026
g27591 nor pi0781 n30008 ; n30027
g27592 nor n30026 n30027 ; n30028
g27593 nor pi0619 n30028 ; n30029
g27594 and pi0619 n29903_not ; n30030
g27595 nor pi1159 n30030 ; n30031
g27596 and n30029_not n30031 ; n30032
g27597 and pi0619_not n29870 ; n30033
g27598 nor pi0781 n29958 ; n30034
g27599 nor n29961 n30018 ; n30035
g27600 and pi0781 n30035_not ; n30036
g27601 nor n30034 n30036 ; n30037
g27602 and pi0619 n30037 ; n30038
g27603 and pi1159 n30033_not ; n30039
g27604 and n30038_not n30039 ; n30040
g27605 nor pi0648 n30040 ; n30041
g27606 and n30032_not n30041 ; n30042
g27607 and pi0619 n30028_not ; n30043
g27608 nor pi0619 n29903 ; n30044
g27609 and pi1159 n30044_not ; n30045
g27610 and n30043_not n30045 ; n30046
g27611 and pi0619_not n30037 ; n30047
g27612 and pi0619 n29870 ; n30048
g27613 nor pi1159 n30048 ; n30049
g27614 and n30047_not n30049 ; n30050
g27615 and pi0648 n30050_not ; n30051
g27616 and n30046_not n30051 ; n30052
g27617 nor n30042 n30052 ; n30053
g27618 and pi0789 n30053_not ; n30054
g27619 nor pi0789 n30028 ; n30055
g27620 nor n30054 n30055 ; n30056
g27621 and pi0788_not n30056 ; n30057
g27622 and pi0626_not n30056 ; n30058
g27623 and pi0626 n29905_not ; n30059
g27624 nor pi0641 n30059 ; n30060
g27625 and n30058_not n30060 ; n30061
g27626 nor pi0789 n30037 ; n30062
g27627 nor n30040 n30050 ; n30063
g27628 and pi0789 n30063_not ; n30064
g27629 nor n30062 n30064 ; n30065
g27630 nor pi0626 n30065 ; n30066
g27631 and pi0626 n29870_not ; n30067
g27632 and pi0641 n30067_not ; n30068
g27633 and n30066_not n30068 ; n30069
g27634 nor pi1158 n30069 ; n30070
g27635 and n30061_not n30070 ; n30071
g27636 and pi0626 n30056 ; n30072
g27637 nor pi0626 n29905 ; n30073
g27638 and pi0641 n30073_not ; n30074
g27639 and n30072_not n30074 ; n30075
g27640 and pi0626 n30065_not ; n30076
g27641 nor pi0626 n29870 ; n30077
g27642 nor pi0641 n30077 ; n30078
g27643 and n30076_not n30078 ; n30079
g27644 and pi1158 n30079_not ; n30080
g27645 and n30075_not n30080 ; n30081
g27646 nor n30071 n30081 ; n30082
g27647 and pi0788 n30082_not ; n30083
g27648 nor n30057 n30083 ; n30084
g27649 and pi0628_not n30084 ; n30085
g27650 and n17969_not n30065 ; n30086
g27651 and n17969 n29870 ; n30087
g27652 nor n30086 n30087 ; n30088
g27653 and pi0628 n30088_not ; n30089
g27654 nor pi1156 n30089 ; n30090
g27655 and n30085_not n30090 ; n30091
g27656 nor pi0629 n29913 ; n30092
g27657 and n30091_not n30092 ; n30093
g27658 and pi0628 n30084 ; n30094
g27659 nor pi0628 n30088 ; n30095
g27660 and pi1156 n30095_not ; n30096
g27661 and n30094_not n30096 ; n30097
g27662 and pi0629 n29917_not ; n30098
g27663 and n30097_not n30098 ; n30099
g27664 nor n30093 n30099 ; n30100
g27665 and pi0792 n30100_not ; n30101
g27666 and pi0792_not n30084 ; n30102
g27667 nor n30101 n30102 ; n30103
g27668 nor pi0647 n30103 ; n30104
g27669 nor n17779 n30088 ; n30105
g27670 and n17779 n29870 ; n30106
g27671 nor n30105 n30106 ; n30107
g27672 and pi0647 n30107_not ; n30108
g27673 nor pi1157 n30108 ; n30109
g27674 and n30104_not n30109 ; n30110
g27675 nor pi0630 n29925 ; n30111
g27676 and n30110_not n30111 ; n30112
g27677 and pi0647 n30103_not ; n30113
g27678 nor pi0647 n30107 ; n30114
g27679 and pi1157 n30114_not ; n30115
g27680 and n30113_not n30115 ; n30116
g27681 and pi0630 n29929_not ; n30117
g27682 and n30116_not n30117 ; n30118
g27683 nor n30112 n30118 ; n30119
g27684 and pi0787 n30119_not ; n30120
g27685 nor pi0787 n30103 ; n30121
g27686 nor n30120 n30121 ; n30122
g27687 and pi0644 n30122_not ; n30123
g27688 and pi0715 n29933_not ; n30124
g27689 and n30123_not n30124 ; n30125
g27690 and n17804 n29870_not ; n30126
g27691 and n17804_not n30107 ; n30127
g27692 nor n30126 n30127 ; n30128
g27693 and pi0644 n30128 ; n30129
g27694 and pi0644_not n29870 ; n30130
g27695 nor pi0715 n30130 ; n30131
g27696 and n30129_not n30131 ; n30132
g27697 and pi1160 n30132_not ; n30133
g27698 and n30125_not n30133 ; n30134
g27699 nor pi0644 n30122 ; n30135
g27700 and pi0644 n29932 ; n30136
g27701 nor pi0715 n30136 ; n30137
g27702 and n30135_not n30137 ; n30138
g27703 and pi0644_not n30128 ; n30139
g27704 and pi0644 n29870 ; n30140
g27705 and pi0715 n30140_not ; n30141
g27706 and n30139_not n30141 ; n30142
g27707 nor pi1160 n30142 ; n30143
g27708 and n30138_not n30143 ; n30144
g27709 and pi0790 n30134_not ; n30145
g27710 and n30144_not n30145 ; n30146
g27711 and pi0790_not n30122 ; n30147
g27712 nor po1038 n30147 ; n30148
g27713 and n30146_not n30148 ; n30149
g27714 and pi0188_not po1038 ; n30150
g27715 nor pi0832 n30150 ; n30151
g27716 and n30149_not n30151 ; n30152
g27717 nor pi0188 n2926 ; n30153
g27718 and pi0705 n16645 ; n30154
g27719 nor n30153 n30154 ; n30155
g27720 and pi0778_not n30155 ; n30156
g27721 and pi0625_not n30154 ; n30157
g27722 nor n30155 n30157 ; n30158
g27723 and pi1153 n30158_not ; n30159
g27724 nor pi1153 n30153 ; n30160
g27725 and n30157_not n30160 ; n30161
g27726 nor n30159 n30161 ; n30162
g27727 and pi0778 n30162_not ; n30163
g27728 nor n30156 n30163 ; n30164
g27729 and n17845_not n30164 ; n30165
g27730 and n17847_not n30165 ; n30166
g27731 and n17849_not n30166 ; n30167
g27732 and n17851_not n30167 ; n30168
g27733 and n17857_not n30168 ; n30169
g27734 and pi0647_not n30169 ; n30170
g27735 and pi0647 n30153 ; n30171
g27736 nor pi1157 n30171 ; n30172
g27737 and n30170_not n30172 ; n30173
g27738 and pi0630 n30173 ; n30174
g27739 and pi0768_not n17244 ; n30175
g27740 nor n30153 n30175 ; n30176
g27741 nor n17874 n30176 ; n30177
g27742 nor pi0785 n30177 ; n30178
g27743 nor n17879 n30176 ; n30179
g27744 and pi1155 n30179_not ; n30180
g27745 and n17882_not n30177 ; n30181
g27746 nor pi1155 n30181 ; n30182
g27747 nor n30180 n30182 ; n30183
g27748 and pi0785 n30183_not ; n30184
g27749 nor n30178 n30184 ; n30185
g27750 nor pi0781 n30185 ; n30186
g27751 and n17889_not n30185 ; n30187
g27752 and pi1154 n30187_not ; n30188
g27753 and n17892_not n30185 ; n30189
g27754 nor pi1154 n30189 ; n30190
g27755 nor n30188 n30190 ; n30191
g27756 and pi0781 n30191_not ; n30192
g27757 nor n30186 n30192 ; n30193
g27758 nor pi0789 n30193 ; n30194
g27759 and pi0619_not n30153 ; n30195
g27760 and pi0619 n30193 ; n30196
g27761 and pi1159 n30195_not ; n30197
g27762 and n30196_not n30197 ; n30198
g27763 and pi0619_not n30193 ; n30199
g27764 and pi0619 n30153 ; n30200
g27765 nor pi1159 n30200 ; n30201
g27766 and n30199_not n30201 ; n30202
g27767 nor n30198 n30202 ; n30203
g27768 and pi0789 n30203_not ; n30204
g27769 nor n30194 n30204 ; n30205
g27770 and n17969_not n30205 ; n30206
g27771 and n17969 n30153 ; n30207
g27772 nor n30206 n30207 ; n30208
g27773 nor n17779 n30208 ; n30209
g27774 and n17779 n30153 ; n30210
g27775 nor n30209 n30210 ; n30211
g27776 and n20559_not n30211 ; n30212
g27777 and pi0647 n30169_not ; n30213
g27778 nor pi0647 n30153 ; n30214
g27779 nor n30213 n30214 ; n30215
g27780 and n17801 n30215_not ; n30216
g27781 nor n30174 n30216 ; n30217
g27782 and n30212_not n30217 ; n30218
g27783 and pi0787 n30218_not ; n30219
g27784 and n17871 n30167 ; n30220
g27785 nor pi0626 n30205 ; n30221
g27786 and pi0626 n30153_not ; n30222
g27787 and n16629 n30222_not ; n30223
g27788 and n30221_not n30223 ; n30224
g27789 and pi0626 n30205_not ; n30225
g27790 nor pi0626 n30153 ; n30226
g27791 and n16628 n30226_not ; n30227
g27792 and n30225_not n30227 ; n30228
g27793 nor n30220 n30224 ; n30229
g27794 and n30228_not n30229 ; n30230
g27795 and pi0788 n30230_not ; n30231
g27796 and pi0618 n30165 ; n30232
g27797 and pi0609 n30164 ; n30233
g27798 nor n17168 n30155 ; n30234
g27799 and pi0625 n30234 ; n30235
g27800 and n30176 n30234_not ; n30236
g27801 nor n30235 n30236 ; n30237
g27802 and n30160 n30237_not ; n30238
g27803 nor pi0608 n30159 ; n30239
g27804 and n30238_not n30239 ; n30240
g27805 and pi1153 n30176 ; n30241
g27806 and n30235_not n30241 ; n30242
g27807 and pi0608 n30161_not ; n30243
g27808 and n30242_not n30243 ; n30244
g27809 nor n30240 n30244 ; n30245
g27810 and pi0778 n30245_not ; n30246
g27811 nor pi0778 n30236 ; n30247
g27812 nor n30246 n30247 ; n30248
g27813 nor pi0609 n30248 ; n30249
g27814 nor pi1155 n30233 ; n30250
g27815 and n30249_not n30250 ; n30251
g27816 nor pi0660 n30180 ; n30252
g27817 and n30251_not n30252 ; n30253
g27818 and pi0609_not n30164 ; n30254
g27819 and pi0609 n30248_not ; n30255
g27820 and pi1155 n30254_not ; n30256
g27821 and n30255_not n30256 ; n30257
g27822 and pi0660 n30182_not ; n30258
g27823 and n30257_not n30258 ; n30259
g27824 nor n30253 n30259 ; n30260
g27825 and pi0785 n30260_not ; n30261
g27826 nor pi0785 n30248 ; n30262
g27827 nor n30261 n30262 ; n30263
g27828 nor pi0618 n30263 ; n30264
g27829 nor pi1154 n30232 ; n30265
g27830 and n30264_not n30265 ; n30266
g27831 nor pi0627 n30188 ; n30267
g27832 and n30266_not n30267 ; n30268
g27833 and pi0618_not n30165 ; n30269
g27834 and pi0618 n30263_not ; n30270
g27835 and pi1154 n30269_not ; n30271
g27836 and n30270_not n30271 ; n30272
g27837 and pi0627 n30190_not ; n30273
g27838 and n30272_not n30273 ; n30274
g27839 nor n30268 n30274 ; n30275
g27840 and pi0781 n30275_not ; n30276
g27841 nor pi0781 n30263 ; n30277
g27842 nor n30276 n30277 ; n30278
g27843 and pi0789_not n30278 ; n30279
g27844 nor pi0619 n30278 ; n30280
g27845 and pi0619 n30166 ; n30281
g27846 nor pi1159 n30281 ; n30282
g27847 and n30280_not n30282 ; n30283
g27848 nor pi0648 n30198 ; n30284
g27849 and n30283_not n30284 ; n30285
g27850 and pi0619 n30278_not ; n30286
g27851 and pi0619_not n30166 ; n30287
g27852 and pi1159 n30287_not ; n30288
g27853 and n30286_not n30288 ; n30289
g27854 and pi0648 n30202_not ; n30290
g27855 and n30289_not n30290 ; n30291
g27856 and pi0789 n30285_not ; n30292
g27857 and n30291_not n30292 ; n30293
g27858 and n17970 n30279_not ; n30294
g27859 and n30293_not n30294 ; n30295
g27860 nor n30231 n30295 ; n30296
g27861 nor n20364 n30296 ; n30297
g27862 and n17854 n30208_not ; n30298
g27863 and n20851 n30168 ; n30299
g27864 nor n30298 n30299 ; n30300
g27865 nor pi0629 n30300 ; n30301
g27866 and n20855 n30168 ; n30302
g27867 and n17853 n30208_not ; n30303
g27868 nor n30302 n30303 ; n30304
g27869 and pi0629 n30304_not ; n30305
g27870 nor n30301 n30305 ; n30306
g27871 and pi0792 n30306_not ; n30307
g27872 nor n20206 n30307 ; n30308
g27873 and n30297_not n30308 ; n30309
g27874 nor n30219 n30309 ; n30310
g27875 and pi0790_not n30310 ; n30311
g27876 nor pi0787 n30169 ; n30312
g27877 and pi1157 n30215_not ; n30313
g27878 nor n30173 n30313 ; n30314
g27879 and pi0787 n30314_not ; n30315
g27880 nor n30312 n30315 ; n30316
g27881 and pi0644_not n30316 ; n30317
g27882 and pi0644 n30310 ; n30318
g27883 and pi0715 n30317_not ; n30319
g27884 and n30318_not n30319 ; n30320
g27885 nor n17804 n30211 ; n30321
g27886 and n17804 n30153 ; n30322
g27887 nor n30321 n30322 ; n30323
g27888 and pi0644 n30323_not ; n30324
g27889 and pi0644_not n30153 ; n30325
g27890 nor pi0715 n30325 ; n30326
g27891 and n30324_not n30326 ; n30327
g27892 and pi1160 n30327_not ; n30328
g27893 and n30320_not n30328 ; n30329
g27894 nor pi0644 n30323 ; n30330
g27895 and pi0644 n30153 ; n30331
g27896 and pi0715 n30331_not ; n30332
g27897 and n30330_not n30332 ; n30333
g27898 and pi0644 n30316 ; n30334
g27899 and pi0644_not n30310 ; n30335
g27900 nor pi0715 n30334 ; n30336
g27901 and n30335_not n30336 ; n30337
g27902 nor pi1160 n30333 ; n30338
g27903 and n30337_not n30338 ; n30339
g27904 nor n30329 n30339 ; n30340
g27905 and pi0790 n30340_not ; n30341
g27906 and pi0832 n30311_not ; n30342
g27907 and n30341_not n30342 ; n30343
g27908 nor n30152 n30343 ; po0345
g27909 and pi0189 n17059_not ; n30345
g27910 and n16635 n30345_not ; n30346
g27911 and n17075 n30345_not ; n30347
g27912 and pi0727 n2571 ; n30348
g27913 nor n30345 n30348 ; n30349
g27914 nor pi0189 n16641 ; n30350
g27915 and n19899 n30350_not ; n30351
g27916 and pi0189_not n18076 ; n30352
g27917 and pi0189 n18072_not ; n30353
g27918 nor pi0038 n30352 ; n30354
g27919 and n30353_not n30354 ; n30355
g27920 and n30348 n30351_not ; n30356
g27921 and n30355_not n30356 ; n30357
g27922 nor n30349 n30357 ; n30358
g27923 and pi0778_not n30358 ; n30359
g27924 nor pi0625 n30345 ; n30360
g27925 and pi0625 n30358_not ; n30361
g27926 and pi1153 n30360_not ; n30362
g27927 and n30361_not n30362 ; n30363
g27928 nor pi0625 n30358 ; n30364
g27929 and pi0625 n30345_not ; n30365
g27930 nor pi1153 n30365 ; n30366
g27931 and n30364_not n30366 ; n30367
g27932 nor n30363 n30367 ; n30368
g27933 and pi0778 n30368_not ; n30369
g27934 nor n30359 n30369 ; n30370
g27935 and n17075_not n30370 ; n30371
g27936 nor n30347 n30371 ; n30372
g27937 and n16639_not n30372 ; n30373
g27938 and n16639 n30345 ; n30374
g27939 nor n30373 n30374 ; n30375
g27940 and n16635_not n30375 ; n30376
g27941 nor n30346 n30376 ; n30377
g27942 and n16631_not n30377 ; n30378
g27943 and n16631 n30345 ; n30379
g27944 nor n30378 n30379 ; n30380
g27945 nor pi0792 n30380 ; n30381
g27946 nor pi0628 n30345 ; n30382
g27947 and pi0628 n30380 ; n30383
g27948 and pi1156 n30382_not ; n30384
g27949 and n30383_not n30384 ; n30385
g27950 and pi0628 n30345_not ; n30386
g27951 and pi0628_not n30380 ; n30387
g27952 nor pi1156 n30386 ; n30388
g27953 and n30387_not n30388 ; n30389
g27954 nor n30385 n30389 ; n30390
g27955 and pi0792 n30390_not ; n30391
g27956 nor n30381 n30391 ; n30392
g27957 nor pi0787 n30392 ; n30393
g27958 nor pi0647 n30345 ; n30394
g27959 and pi0647 n30392 ; n30395
g27960 and pi1157 n30394_not ; n30396
g27961 and n30395_not n30396 ; n30397
g27962 and pi0647 n30345_not ; n30398
g27963 and pi0647_not n30392 ; n30399
g27964 nor pi1157 n30398 ; n30400
g27965 and n30399_not n30400 ; n30401
g27966 nor n30397 n30401 ; n30402
g27967 and pi0787 n30402_not ; n30403
g27968 nor n30393 n30403 ; n30404
g27969 and pi0644_not n30404 ; n30405
g27970 nor pi0619 n30345 ; n30406
g27971 and n17117 n30345_not ; n30407
g27972 and pi0189 n2571_not ; n30408
g27973 and pi0772 n17219 ; n30409
g27974 nor n22241 n30409 ; n30410
g27975 and pi0039 n30410_not ; n30411
g27976 and pi0772_not n16958 ; n30412
g27977 and pi0772 n17139 ; n30413
g27978 nor pi0039 n30412 ; n30414
g27979 and n30413_not n30414 ; n30415
g27980 nor n30411 n30415 ; n30416
g27981 and pi0189 n30416_not ; n30417
g27982 and pi0189_not pi0772 ; n30418
g27983 and n17275 n30418 ; n30419
g27984 nor n30417 n30419 ; n30420
g27985 nor pi0038 n30420 ; n30421
g27986 and pi0772 n17168 ; n30422
g27987 and n16641 n30422_not ; n30423
g27988 and pi0038 n30350_not ; n30424
g27989 and n30423_not n30424 ; n30425
g27990 nor n30421 n30425 ; n30426
g27991 and n2571 n30426_not ; n30427
g27992 nor n30408 n30427 ; n30428
g27993 and n17117_not n30428 ; n30429
g27994 nor n30407 n30429 ; n30430
g27995 and pi0785_not n30430 ; n30431
g27996 nor pi0609 n30345 ; n30432
g27997 and pi0609 n30430_not ; n30433
g27998 and pi1155 n30432_not ; n30434
g27999 and n30433_not n30434 ; n30435
g28000 nor pi0609 n30430 ; n30436
g28001 and pi0609 n30345_not ; n30437
g28002 nor pi1155 n30437 ; n30438
g28003 and n30436_not n30438 ; n30439
g28004 nor n30435 n30439 ; n30440
g28005 and pi0785 n30440_not ; n30441
g28006 nor n30431 n30441 ; n30442
g28007 nor pi0781 n30442 ; n30443
g28008 nor pi0618 n30345 ; n30444
g28009 and pi0618 n30442 ; n30445
g28010 and pi1154 n30444_not ; n30446
g28011 and n30445_not n30446 ; n30447
g28012 and pi0618 n30345_not ; n30448
g28013 and pi0618_not n30442 ; n30449
g28014 nor pi1154 n30448 ; n30450
g28015 and n30449_not n30450 ; n30451
g28016 nor n30447 n30451 ; n30452
g28017 and pi0781 n30452_not ; n30453
g28018 nor n30443 n30453 ; n30454
g28019 and pi0619 n30454 ; n30455
g28020 and pi1159 n30406_not ; n30456
g28021 and n30455_not n30456 ; n30457
g28022 and pi0727_not n30426 ; n30458
g28023 nor pi0189 n17605 ; n30459
g28024 and pi0189 n17546 ; n30460
g28025 and pi0772 n30460_not ; n30461
g28026 and n30459_not n30461 ; n30462
g28027 and pi0189 n17404_not ; n30463
g28028 nor pi0189 n17485 ; n30464
g28029 nor pi0772 n30464 ; n30465
g28030 and n30463_not n30465 ; n30466
g28031 and pi0039 n30462_not ; n30467
g28032 and n30466_not n30467 ; n30468
g28033 and pi0189_not n17631 ; n30469
g28034 and pi0189 n17629 ; n30470
g28035 and pi0772 n30469_not ; n30471
g28036 and n30470_not n30471 ; n30472
g28037 nor pi0189 n17625 ; n30473
g28038 and pi0189 n17612_not ; n30474
g28039 nor pi0772 n30473 ; n30475
g28040 and n30474_not n30475 ; n30476
g28041 nor pi0039 n30472 ; n30477
g28042 and n30476_not n30477 ; n30478
g28043 nor pi0038 n30478 ; n30479
g28044 and n30468_not n30479 ; n30480
g28045 and pi0727 n19470_not ; n30481
g28046 and n30425_not n30481 ; n30482
g28047 and n30480_not n30482 ; n30483
g28048 and n2571 n30483_not ; n30484
g28049 and n30458_not n30484 ; n30485
g28050 nor n30408 n30485 ; n30486
g28051 and pi0625_not n30486 ; n30487
g28052 and pi0625 n30428 ; n30488
g28053 nor pi1153 n30488 ; n30489
g28054 and n30487_not n30489 ; n30490
g28055 nor pi0608 n30363 ; n30491
g28056 and n30490_not n30491 ; n30492
g28057 and pi0625_not n30428 ; n30493
g28058 and pi0625 n30486 ; n30494
g28059 and pi1153 n30493_not ; n30495
g28060 and n30494_not n30495 ; n30496
g28061 and pi0608 n30367_not ; n30497
g28062 and n30496_not n30497 ; n30498
g28063 nor n30492 n30498 ; n30499
g28064 and pi0778 n30499_not ; n30500
g28065 and pi0778_not n30486 ; n30501
g28066 nor n30500 n30501 ; n30502
g28067 nor pi0609 n30502 ; n30503
g28068 and pi0609 n30370 ; n30504
g28069 nor pi1155 n30504 ; n30505
g28070 and n30503_not n30505 ; n30506
g28071 nor pi0660 n30435 ; n30507
g28072 and n30506_not n30507 ; n30508
g28073 and pi0609_not n30370 ; n30509
g28074 and pi0609 n30502_not ; n30510
g28075 and pi1155 n30509_not ; n30511
g28076 and n30510_not n30511 ; n30512
g28077 and pi0660 n30439_not ; n30513
g28078 and n30512_not n30513 ; n30514
g28079 nor n30508 n30514 ; n30515
g28080 and pi0785 n30515_not ; n30516
g28081 nor pi0785 n30502 ; n30517
g28082 nor n30516 n30517 ; n30518
g28083 nor pi0618 n30518 ; n30519
g28084 and pi0618 n30372_not ; n30520
g28085 nor pi1154 n30520 ; n30521
g28086 and n30519_not n30521 ; n30522
g28087 nor pi0627 n30447 ; n30523
g28088 and n30522_not n30523 ; n30524
g28089 and pi0618 n30518_not ; n30525
g28090 nor pi0618 n30372 ; n30526
g28091 and pi1154 n30526_not ; n30527
g28092 and n30525_not n30527 ; n30528
g28093 and pi0627 n30451_not ; n30529
g28094 and n30528_not n30529 ; n30530
g28095 nor n30524 n30530 ; n30531
g28096 and pi0781 n30531_not ; n30532
g28097 nor pi0781 n30518 ; n30533
g28098 nor n30532 n30533 ; n30534
g28099 nor pi0619 n30534 ; n30535
g28100 and pi0619 n30375 ; n30536
g28101 nor pi1159 n30536 ; n30537
g28102 and n30535_not n30537 ; n30538
g28103 nor pi0648 n30457 ; n30539
g28104 and n30538_not n30539 ; n30540
g28105 and pi0619 n30345_not ; n30541
g28106 and pi0619_not n30454 ; n30542
g28107 nor pi1159 n30541 ; n30543
g28108 and n30542_not n30543 ; n30544
g28109 and pi0619_not n30375 ; n30545
g28110 and pi0619 n30534_not ; n30546
g28111 and pi1159 n30545_not ; n30547
g28112 and n30546_not n30547 ; n30548
g28113 and pi0648 n30544_not ; n30549
g28114 and n30548_not n30549 ; n30550
g28115 nor n30540 n30550 ; n30551
g28116 and pi0789 n30551_not ; n30552
g28117 nor pi0789 n30534 ; n30553
g28118 nor n30552 n30553 ; n30554
g28119 and pi0788_not n30554 ; n30555
g28120 and pi0626_not n30554 ; n30556
g28121 and pi0626 n30377 ; n30557
g28122 nor pi0641 n30557 ; n30558
g28123 and n30556_not n30558 ; n30559
g28124 nor pi0789 n30454 ; n30560
g28125 nor n30457 n30544 ; n30561
g28126 and pi0789 n30561_not ; n30562
g28127 nor n30560 n30562 ; n30563
g28128 nor pi0626 n30563 ; n30564
g28129 and pi0626 n30345 ; n30565
g28130 and pi0641 n30565_not ; n30566
g28131 and n30564_not n30566 ; n30567
g28132 nor pi1158 n30567 ; n30568
g28133 and n30559_not n30568 ; n30569
g28134 and pi0626 n30554 ; n30570
g28135 and pi0626_not n30377 ; n30571
g28136 and pi0641 n30571_not ; n30572
g28137 and n30570_not n30572 ; n30573
g28138 and pi0626 n30563_not ; n30574
g28139 and pi0626_not n30345 ; n30575
g28140 nor pi0641 n30575 ; n30576
g28141 and n30574_not n30576 ; n30577
g28142 and pi1158 n30577_not ; n30578
g28143 and n30573_not n30578 ; n30579
g28144 nor n30569 n30579 ; n30580
g28145 and pi0788 n30580_not ; n30581
g28146 nor n30555 n30581 ; n30582
g28147 and pi0628_not n30582 ; n30583
g28148 nor n17969 n30563 ; n30584
g28149 and n17969 n30345 ; n30585
g28150 nor n30584 n30585 ; n30586
g28151 and pi0628 n30586 ; n30587
g28152 nor pi1156 n30587 ; n30588
g28153 and n30583_not n30588 ; n30589
g28154 nor pi0629 n30385 ; n30590
g28155 and n30589_not n30590 ; n30591
g28156 and pi0628 n30582 ; n30592
g28157 and pi0628_not n30586 ; n30593
g28158 and pi1156 n30593_not ; n30594
g28159 and n30592_not n30594 ; n30595
g28160 and pi0629 n30389_not ; n30596
g28161 and n30595_not n30596 ; n30597
g28162 nor n30591 n30597 ; n30598
g28163 and pi0792 n30598_not ; n30599
g28164 and pi0792_not n30582 ; n30600
g28165 nor n30599 n30600 ; n30601
g28166 nor pi0647 n30601 ; n30602
g28167 nor n17779 n30586 ; n30603
g28168 and n17779 n30345 ; n30604
g28169 nor n30603 n30604 ; n30605
g28170 and pi0647 n30605 ; n30606
g28171 nor pi1157 n30606 ; n30607
g28172 and n30602_not n30607 ; n30608
g28173 nor pi0630 n30397 ; n30609
g28174 and n30608_not n30609 ; n30610
g28175 and pi0647 n30601_not ; n30611
g28176 and pi0647_not n30605 ; n30612
g28177 and pi1157 n30612_not ; n30613
g28178 and n30611_not n30613 ; n30614
g28179 and pi0630 n30401_not ; n30615
g28180 and n30614_not n30615 ; n30616
g28181 nor n30610 n30616 ; n30617
g28182 and pi0787 n30617_not ; n30618
g28183 nor pi0787 n30601 ; n30619
g28184 nor n30618 n30619 ; n30620
g28185 and pi0644 n30620_not ; n30621
g28186 and pi0715 n30405_not ; n30622
g28187 and n30621_not n30622 ; n30623
g28188 and n17804 n30345_not ; n30624
g28189 and n17804_not n30605 ; n30625
g28190 nor n30624 n30625 ; n30626
g28191 and pi0644 n30626_not ; n30627
g28192 nor pi0644 n30345 ; n30628
g28193 nor pi0715 n30628 ; n30629
g28194 and n30627_not n30629 ; n30630
g28195 and pi1160 n30630_not ; n30631
g28196 and n30623_not n30631 ; n30632
g28197 nor pi0644 n30620 ; n30633
g28198 and pi0644 n30404 ; n30634
g28199 nor pi0715 n30634 ; n30635
g28200 and n30633_not n30635 ; n30636
g28201 nor pi0644 n30626 ; n30637
g28202 and pi0644 n30345_not ; n30638
g28203 and pi0715 n30638_not ; n30639
g28204 and n30637_not n30639 ; n30640
g28205 nor pi1160 n30640 ; n30641
g28206 and n30636_not n30641 ; n30642
g28207 and pi0790 n30632_not ; n30643
g28208 and n30642_not n30643 ; n30644
g28209 and pi0790_not n30620 ; n30645
g28210 and n6305 n30645_not ; n30646
g28211 and n30644_not n30646 ; n30647
g28212 nor pi0189 n6305 ; n30648
g28213 nor pi0057 n30648 ; n30649
g28214 and n30647_not n30649 ; n30650
g28215 and pi0057 pi0189 ; n30651
g28216 nor pi0832 n30651 ; n30652
g28217 and n30650_not n30652 ; n30653
g28218 and pi0189 n2926_not ; n30654
g28219 and pi0772 n17244 ; n30655
g28220 and n17291 n30655 ; n30656
g28221 and pi1155 n30654_not ; n30657
g28222 and n30656_not n30657 ; n30658
g28223 and pi0727 n16645 ; n30659
g28224 nor n30654 n30659 ; n30660
g28225 and pi0778_not n30660 ; n30661
g28226 and pi0625 n30659 ; n30662
g28227 nor n30660 n30662 ; n30663
g28228 nor pi1153 n30663 ; n30664
g28229 and pi1153 n30654_not ; n30665
g28230 and n30662_not n30665 ; n30666
g28231 nor n30664 n30666 ; n30667
g28232 and pi0778 n30667_not ; n30668
g28233 nor n30661 n30668 ; n30669
g28234 and pi0609 n30669 ; n30670
g28235 nor n30654 n30655 ; n30671
g28236 and pi0727 n17469 ; n30672
g28237 and n30671 n30672_not ; n30673
g28238 and pi0625 n30672 ; n30674
g28239 nor n30673 n30674 ; n30675
g28240 nor pi1153 n30675 ; n30676
g28241 nor pi0608 n30666 ; n30677
g28242 and n30676_not n30677 ; n30678
g28243 and pi1153 n30671 ; n30679
g28244 and n30674_not n30679 ; n30680
g28245 and pi0608 n30664_not ; n30681
g28246 and n30680_not n30681 ; n30682
g28247 nor n30678 n30682 ; n30683
g28248 and pi0778 n30683_not ; n30684
g28249 nor pi0778 n30673 ; n30685
g28250 nor n30684 n30685 ; n30686
g28251 nor pi0609 n30686 ; n30687
g28252 nor pi1155 n30670 ; n30688
g28253 and n30687_not n30688 ; n30689
g28254 nor pi0660 n30658 ; n30690
g28255 and n30689_not n30690 ; n30691
g28256 and n17296 n30655 ; n30692
g28257 nor pi1155 n30654 ; n30693
g28258 and n30692_not n30693 ; n30694
g28259 and pi0609_not n30669 ; n30695
g28260 and pi0609 n30686_not ; n30696
g28261 and pi1155 n30695_not ; n30697
g28262 and n30696_not n30697 ; n30698
g28263 and pi0660 n30694_not ; n30699
g28264 and n30698_not n30699 ; n30700
g28265 nor n30691 n30700 ; n30701
g28266 and pi0785 n30701_not ; n30702
g28267 nor pi0785 n30686 ; n30703
g28268 nor n30702 n30703 ; n30704
g28269 nor pi0781 n30704 ; n30705
g28270 and n20225_not n30655 ; n30706
g28271 and n20319 n30706 ; n30707
g28272 nor pi1154 n30654 ; n30708
g28273 and n30707_not n30708 ; n30709
g28274 and n17075_not n30669 ; n30710
g28275 nor n30654 n30710 ; n30711
g28276 nor pi0618 n30711 ; n30712
g28277 and pi0618 n30704_not ; n30713
g28278 and pi1154 n30712_not ; n30714
g28279 and n30713_not n30714 ; n30715
g28280 and pi0627 n30709_not ; n30716
g28281 and n30715_not n30716 ; n30717
g28282 and n20270 n30706 ; n30718
g28283 and pi1154 n30654_not ; n30719
g28284 and n30718_not n30719 ; n30720
g28285 and pi0618 n30711_not ; n30721
g28286 nor pi0618 n30704 ; n30722
g28287 nor pi1154 n30721 ; n30723
g28288 and n30722_not n30723 ; n30724
g28289 nor pi0627 n30720 ; n30725
g28290 and n30724_not n30725 ; n30726
g28291 nor n30717 n30726 ; n30727
g28292 and pi0781 n30727_not ; n30728
g28293 nor n23615 n30705 ; n30729
g28294 and n30728_not n30729 ; n30730
g28295 and n20235_not n30706 ; n30731
g28296 and n20345 n30731 ; n30732
g28297 and n16633 n30732_not ; n30733
g28298 and n19150 n30669 ; n30734
g28299 nor n23613 n30734 ; n30735
g28300 and n20335 n30731 ; n30736
g28301 and n16632 n30736_not ; n30737
g28302 nor n30733 n30737 ; n30738
g28303 and n30735_not n30738 ; n30739
g28304 and pi0789 n30654_not ; n30740
g28305 and n30739_not n30740 ; n30741
g28306 and n17970 n30741_not ; n30742
g28307 and n30730_not n30742 ; n30743
g28308 and n16635_not n30734 ; n30744
g28309 nor n30654 n30744 ; n30745
g28310 and n17865 n30745_not ; n30746
g28311 and n20237 n30706 ; n30747
g28312 and pi0626_not n30747 ; n30748
g28313 nor n30654 n30748 ; n30749
g28314 nor pi1158 n30749 ; n30750
g28315 and pi0641 n30750_not ; n30751
g28316 and n30746_not n30751 ; n30752
g28317 and pi0626 n30747 ; n30753
g28318 nor n30654 n30753 ; n30754
g28319 and pi1158 n30754_not ; n30755
g28320 and n17866 n30745_not ; n30756
g28321 nor pi0641 n30755 ; n30757
g28322 and n30756_not n30757 ; n30758
g28323 and pi0788 n30752_not ; n30759
g28324 and n30758_not n30759 ; n30760
g28325 nor n20364 n30760 ; n30761
g28326 and n30743_not n30761 ; n30762
g28327 and n17969_not n30747 ; n30763
g28328 and pi0629_not n30763 ; n30764
g28329 and pi0628 n30764_not ; n30765
g28330 and n19151 n30669 ; n30766
g28331 and pi0629 n30766_not ; n30767
g28332 nor n30765 n30767 ; n30768
g28333 nor pi1156 n30768 ; n30769
g28334 nor pi0628 n30763 ; n30770
g28335 and pi0629 n30770_not ; n30771
g28336 and pi0628 n30766 ; n30772
g28337 and pi1156 n30771_not ; n30773
g28338 and n30772_not n30773 ; n30774
g28339 nor n30769 n30774 ; n30775
g28340 and pi0792 n30654_not ; n30776
g28341 and n30775_not n30776 ; n30777
g28342 nor n30762 n30777 ; n30778
g28343 nor n20206 n30778 ; n30779
g28344 and n17779_not n30763 ; n30780
g28345 and pi0630_not n30780 ; n30781
g28346 and pi0647 n30781_not ; n30782
g28347 and n19142_not n30766 ; n30783
g28348 and pi0630 n30783_not ; n30784
g28349 nor n30782 n30784 ; n30785
g28350 nor pi1157 n30785 ; n30786
g28351 and pi0630 n30780 ; n30787
g28352 nor pi0630 n30783 ; n30788
g28353 and pi0647 n30788_not ; n30789
g28354 and pi1157 n30787_not ; n30790
g28355 and n30789_not n30790 ; n30791
g28356 nor n30786 n30791 ; n30792
g28357 and pi0787 n30654_not ; n30793
g28358 and n30792_not n30793 ; n30794
g28359 nor n30779 n30794 ; n30795
g28360 and pi0790_not n30795 ; n30796
g28361 and n17969_not n23684 ; n30797
g28362 and n30747 n30797 ; n30798
g28363 and pi0644 n30798 ; n30799
g28364 nor pi0715 n30654 ; n30800
g28365 and n30799_not n30800 ; n30801
g28366 and n19342_not n30783 ; n30802
g28367 nor n30654 n30802 ; n30803
g28368 nor pi0644 n30803 ; n30804
g28369 and pi0644 n30795 ; n30805
g28370 and pi0715 n30804_not ; n30806
g28371 and n30805_not n30806 ; n30807
g28372 and pi1160 n30801_not ; n30808
g28373 and n30807_not n30808 ; n30809
g28374 and pi0644_not n30798 ; n30810
g28375 and pi0715 n30654_not ; n30811
g28376 and n30810_not n30811 ; n30812
g28377 and pi0644_not n30795 ; n30813
g28378 and pi0644 n30803_not ; n30814
g28379 nor pi0715 n30814 ; n30815
g28380 and n30813_not n30815 ; n30816
g28381 nor pi1160 n30812 ; n30817
g28382 and n30816_not n30817 ; n30818
g28383 nor n30809 n30818 ; n30819
g28384 and pi0790 n30819_not ; n30820
g28385 and pi0832 n30796_not ; n30821
g28386 and n30820_not n30821 ; n30822
g28387 nor n30653 n30822 ; po0346
g28388 nor pi0190 n2926 ; n30824
g28389 and pi0699 n16645 ; n30825
g28390 nor n30824 n30825 ; n30826
g28391 nor pi0778 n30826 ; n30827
g28392 and pi0625_not n30825 ; n30828
g28393 nor n30826 n30828 ; n30829
g28394 and pi1153 n30829_not ; n30830
g28395 nor pi1153 n30824 ; n30831
g28396 and n30828_not n30831 ; n30832
g28397 and pi0778 n30832_not ; n30833
g28398 and n30830_not n30833 ; n30834
g28399 nor n30827 n30834 ; n30835
g28400 nor n17845 n30835 ; n30836
g28401 and n17847_not n30836 ; n30837
g28402 and n17849_not n30837 ; n30838
g28403 and n17851_not n30838 ; n30839
g28404 and n17857_not n30839 ; n30840
g28405 and pi0647_not n30840 ; n30841
g28406 and pi0647 n30824 ; n30842
g28407 nor pi1157 n30842 ; n30843
g28408 and n30841_not n30843 ; n30844
g28409 and pi0630 n30844 ; n30845
g28410 and pi0763 n17244 ; n30846
g28411 nor n30824 n30846 ; n30847
g28412 nor n17874 n30847 ; n30848
g28413 nor pi0785 n30848 ; n30849
g28414 and n17296 n30846 ; n30850
g28415 and n30848 n30850_not ; n30851
g28416 and pi1155 n30851_not ; n30852
g28417 nor pi1155 n30824 ; n30853
g28418 and n30850_not n30853 ; n30854
g28419 nor n30852 n30854 ; n30855
g28420 and pi0785 n30855_not ; n30856
g28421 nor n30849 n30856 ; n30857
g28422 nor pi0781 n30857 ; n30858
g28423 and n17889_not n30857 ; n30859
g28424 and pi1154 n30859_not ; n30860
g28425 and n17892_not n30857 ; n30861
g28426 nor pi1154 n30861 ; n30862
g28427 nor n30860 n30862 ; n30863
g28428 and pi0781 n30863_not ; n30864
g28429 nor n30858 n30864 ; n30865
g28430 nor pi0789 n30865 ; n30866
g28431 and n23078_not n30865 ; n30867
g28432 and pi1159 n30867_not ; n30868
g28433 and n23081_not n30865 ; n30869
g28434 nor pi1159 n30869 ; n30870
g28435 nor n30868 n30870 ; n30871
g28436 and pi0789 n30871_not ; n30872
g28437 nor n30866 n30872 ; n30873
g28438 and n17969_not n30873 ; n30874
g28439 and n17969 n30824 ; n30875
g28440 nor n30874 n30875 ; n30876
g28441 nor n17779 n30876 ; n30877
g28442 and n17779 n30824 ; n30878
g28443 nor n30877 n30878 ; n30879
g28444 and n20559_not n30879 ; n30880
g28445 and pi0647 n30840_not ; n30881
g28446 nor pi0647 n30824 ; n30882
g28447 nor n30881 n30882 ; n30883
g28448 and n17801 n30883_not ; n30884
g28449 nor n30845 n30884 ; n30885
g28450 and n30880_not n30885 ; n30886
g28451 and pi0787 n30886_not ; n30887
g28452 and n17871 n30838 ; n30888
g28453 nor pi0626 n30873 ; n30889
g28454 and pi0626 n30824_not ; n30890
g28455 and n16629 n30890_not ; n30891
g28456 and n30889_not n30891 ; n30892
g28457 and pi0626 n30873_not ; n30893
g28458 nor pi0626 n30824 ; n30894
g28459 and n16628 n30894_not ; n30895
g28460 and n30893_not n30895 ; n30896
g28461 nor n30888 n30892 ; n30897
g28462 and n30896_not n30897 ; n30898
g28463 and pi0788 n30898_not ; n30899
g28464 and pi0618 n30836 ; n30900
g28465 nor n17168 n30826 ; n30901
g28466 and pi0625 n30901 ; n30902
g28467 and n30847 n30901_not ; n30903
g28468 nor n30902 n30903 ; n30904
g28469 and n30831 n30904_not ; n30905
g28470 nor pi0608 n30830 ; n30906
g28471 and n30905_not n30906 ; n30907
g28472 and pi1153 n30847 ; n30908
g28473 and n30902_not n30908 ; n30909
g28474 and pi0608 n30832_not ; n30910
g28475 and n30909_not n30910 ; n30911
g28476 nor n30907 n30911 ; n30912
g28477 and pi0778 n30912_not ; n30913
g28478 nor pi0778 n30903 ; n30914
g28479 nor n30913 n30914 ; n30915
g28480 nor pi0609 n30915 ; n30916
g28481 and pi0609 n30835_not ; n30917
g28482 nor pi1155 n30917 ; n30918
g28483 and n30916_not n30918 ; n30919
g28484 nor pi0660 n30852 ; n30920
g28485 and n30919_not n30920 ; n30921
g28486 and pi0609 n30915_not ; n30922
g28487 nor pi0609 n30835 ; n30923
g28488 and pi1155 n30923_not ; n30924
g28489 and n30922_not n30924 ; n30925
g28490 and pi0660 n30854_not ; n30926
g28491 and n30925_not n30926 ; n30927
g28492 nor n30921 n30927 ; n30928
g28493 and pi0785 n30928_not ; n30929
g28494 nor pi0785 n30915 ; n30930
g28495 nor n30929 n30930 ; n30931
g28496 nor pi0618 n30931 ; n30932
g28497 nor pi1154 n30900 ; n30933
g28498 and n30932_not n30933 ; n30934
g28499 nor pi0627 n30860 ; n30935
g28500 and n30934_not n30935 ; n30936
g28501 and pi0618_not n30836 ; n30937
g28502 and pi0618 n30931_not ; n30938
g28503 and pi1154 n30937_not ; n30939
g28504 and n30938_not n30939 ; n30940
g28505 and pi0627 n30862_not ; n30941
g28506 and n30940_not n30941 ; n30942
g28507 nor n30936 n30942 ; n30943
g28508 and pi0781 n30943_not ; n30944
g28509 nor pi0781 n30931 ; n30945
g28510 nor n30944 n30945 ; n30946
g28511 and pi0789_not n30946 ; n30947
g28512 nor pi0619 n30946 ; n30948
g28513 and pi0619 n30837 ; n30949
g28514 nor pi1159 n30949 ; n30950
g28515 and n30948_not n30950 ; n30951
g28516 nor pi0648 n30868 ; n30952
g28517 and n30951_not n30952 ; n30953
g28518 and pi0619 n30946_not ; n30954
g28519 and pi0619_not n30837 ; n30955
g28520 and pi1159 n30955_not ; n30956
g28521 and n30954_not n30956 ; n30957
g28522 and pi0648 n30870_not ; n30958
g28523 and n30957_not n30958 ; n30959
g28524 and pi0789 n30953_not ; n30960
g28525 and n30959_not n30960 ; n30961
g28526 and n17970 n30947_not ; n30962
g28527 and n30961_not n30962 ; n30963
g28528 nor n30899 n30963 ; n30964
g28529 nor n20364 n30964 ; n30965
g28530 and n17854 n30876_not ; n30966
g28531 and n20851 n30839 ; n30967
g28532 nor n30966 n30967 ; n30968
g28533 nor pi0629 n30968 ; n30969
g28534 and n20855 n30839 ; n30970
g28535 and n17853 n30876_not ; n30971
g28536 nor n30970 n30971 ; n30972
g28537 and pi0629 n30972_not ; n30973
g28538 nor n30969 n30973 ; n30974
g28539 and pi0792 n30974_not ; n30975
g28540 nor n20206 n30975 ; n30976
g28541 and n30965_not n30976 ; n30977
g28542 nor n30887 n30977 ; n30978
g28543 and pi0790_not n30978 ; n30979
g28544 nor pi0787 n30840 ; n30980
g28545 and pi1157 n30883_not ; n30981
g28546 nor n30844 n30981 ; n30982
g28547 and pi0787 n30982_not ; n30983
g28548 nor n30980 n30983 ; n30984
g28549 and pi0644_not n30984 ; n30985
g28550 and pi0644 n30978 ; n30986
g28551 and pi0715 n30985_not ; n30987
g28552 and n30986_not n30987 ; n30988
g28553 nor n17804 n30879 ; n30989
g28554 and n17804 n30824 ; n30990
g28555 nor n30989 n30990 ; n30991
g28556 and pi0644 n30991_not ; n30992
g28557 and pi0644_not n30824 ; n30993
g28558 nor pi0715 n30993 ; n30994
g28559 and n30992_not n30994 ; n30995
g28560 and pi1160 n30995_not ; n30996
g28561 and n30988_not n30996 ; n30997
g28562 nor pi0644 n30991 ; n30998
g28563 and pi0644 n30824 ; n30999
g28564 and pi0715 n30999_not ; n31000
g28565 and n30998_not n31000 ; n31001
g28566 and pi0644 n30984 ; n31002
g28567 and pi0644_not n30978 ; n31003
g28568 nor pi0715 n31002 ; n31004
g28569 and n31003_not n31004 ; n31005
g28570 nor pi1160 n31001 ; n31006
g28571 and n31005_not n31006 ; n31007
g28572 nor n30997 n31007 ; n31008
g28573 and pi0790 n31008_not ; n31009
g28574 and pi0832 n30979_not ; n31010
g28575 and n31009_not n31010 ; n31011
g28576 and pi0190_not po1038 ; n31012
g28577 nor pi0190 n17059 ; n31013
g28578 and n16635 n31013_not ; n31014
g28579 and pi0190 n2571_not ; n31015
g28580 nor pi0190 n16641 ; n31016
g28581 and n16647 n31016_not ; n31017
g28582 and pi0190_not n18072 ; n31018
g28583 and pi0190 n18076_not ; n31019
g28584 nor pi0038 n31019 ; n31020
g28585 and n31018_not n31020 ; n31021
g28586 and pi0699 n31017_not ; n31022
g28587 and n31021_not n31022 ; n31023
g28588 nor pi0190 pi0699 ; n31024
g28589 and n17052_not n31024 ; n31025
g28590 and n2571 n31025_not ; n31026
g28591 and n31023_not n31026 ; n31027
g28592 nor n31015 n31027 ; n31028
g28593 nor pi0778 n31028 ; n31029
g28594 and pi0625_not n31013 ; n31030
g28595 and pi0625 n31028 ; n31031
g28596 and pi1153 n31030_not ; n31032
g28597 and n31031_not n31032 ; n31033
g28598 and pi0625_not n31028 ; n31034
g28599 and pi0625 n31013 ; n31035
g28600 nor pi1153 n31035 ; n31036
g28601 and n31034_not n31036 ; n31037
g28602 nor n31033 n31037 ; n31038
g28603 and pi0778 n31038_not ; n31039
g28604 nor n31029 n31039 ; n31040
g28605 nor n17075 n31040 ; n31041
g28606 and n17075 n31013_not ; n31042
g28607 nor n31041 n31042 ; n31043
g28608 and n16639_not n31043 ; n31044
g28609 and n16639 n31013 ; n31045
g28610 nor n31044 n31045 ; n31046
g28611 and n16635_not n31046 ; n31047
g28612 nor n31014 n31047 ; n31048
g28613 and n16631_not n31048 ; n31049
g28614 and n16631 n31013 ; n31050
g28615 nor n31049 n31050 ; n31051
g28616 nor pi0628 n31051 ; n31052
g28617 and pi0628 n31013 ; n31053
g28618 nor n31052 n31053 ; n31054
g28619 nor pi1156 n31054 ; n31055
g28620 and pi0628 n31051_not ; n31056
g28621 and pi0628_not n31013 ; n31057
g28622 nor n31056 n31057 ; n31058
g28623 and pi1156 n31058_not ; n31059
g28624 nor n31055 n31059 ; n31060
g28625 and pi0792 n31060_not ; n31061
g28626 nor pi0792 n31051 ; n31062
g28627 nor n31061 n31062 ; n31063
g28628 nor pi0647 n31063 ; n31064
g28629 and pi0647 n31013 ; n31065
g28630 nor n31064 n31065 ; n31066
g28631 nor pi1157 n31066 ; n31067
g28632 and pi0647 n31063_not ; n31068
g28633 and pi0647_not n31013 ; n31069
g28634 nor n31068 n31069 ; n31070
g28635 and pi1157 n31070_not ; n31071
g28636 nor n31067 n31071 ; n31072
g28637 and pi0787 n31072_not ; n31073
g28638 nor pi0787 n31063 ; n31074
g28639 nor n31073 n31074 ; n31075
g28640 nor pi0644 n31075 ; n31076
g28641 and pi0715 n31076_not ; n31077
g28642 and pi0763_not n17046 ; n31078
g28643 and pi0190 n17273 ; n31079
g28644 nor n31078 n31079 ; n31080
g28645 and pi0039 n31080_not ; n31081
g28646 and pi0763 n17234_not ; n31082
g28647 and pi0190 n31082_not ; n31083
g28648 and pi0190_not pi0763 ; n31084
g28649 and n17221 n31084 ; n31085
g28650 nor n22358 n31083 ; n31086
g28651 and n31085_not n31086 ; n31087
g28652 and n31081_not n31087 ; n31088
g28653 nor pi0038 n31088 ; n31089
g28654 and pi0763 n17280 ; n31090
g28655 and pi0038 n31016_not ; n31091
g28656 and n31090_not n31091 ; n31092
g28657 nor n31089 n31092 ; n31093
g28658 and n2571 n31093_not ; n31094
g28659 nor n31015 n31094 ; n31095
g28660 nor n17117 n31095 ; n31096
g28661 and n17117 n31013_not ; n31097
g28662 nor n31096 n31097 ; n31098
g28663 nor pi0785 n31098 ; n31099
g28664 nor n17291 n31013 ; n31100
g28665 and pi0609 n31096 ; n31101
g28666 nor n31100 n31101 ; n31102
g28667 and pi1155 n31102_not ; n31103
g28668 nor n17296 n31013 ; n31104
g28669 and pi0609_not n31096 ; n31105
g28670 nor n31104 n31105 ; n31106
g28671 nor pi1155 n31106 ; n31107
g28672 nor n31103 n31107 ; n31108
g28673 and pi0785 n31108_not ; n31109
g28674 nor n31099 n31109 ; n31110
g28675 nor pi0781 n31110 ; n31111
g28676 and pi0618_not n31013 ; n31112
g28677 and pi0618 n31110 ; n31113
g28678 and pi1154 n31112_not ; n31114
g28679 and n31113_not n31114 ; n31115
g28680 and pi0618_not n31110 ; n31116
g28681 and pi0618 n31013 ; n31117
g28682 nor pi1154 n31117 ; n31118
g28683 and n31116_not n31118 ; n31119
g28684 nor n31115 n31119 ; n31120
g28685 and pi0781 n31120_not ; n31121
g28686 nor n31111 n31121 ; n31122
g28687 nor pi0789 n31122 ; n31123
g28688 and pi0619_not n31013 ; n31124
g28689 and pi0619 n31122 ; n31125
g28690 and pi1159 n31124_not ; n31126
g28691 and n31125_not n31126 ; n31127
g28692 and pi0619_not n31122 ; n31128
g28693 and pi0619 n31013 ; n31129
g28694 nor pi1159 n31129 ; n31130
g28695 and n31128_not n31130 ; n31131
g28696 nor n31127 n31131 ; n31132
g28697 and pi0789 n31132_not ; n31133
g28698 nor n31123 n31133 ; n31134
g28699 and n17969_not n31134 ; n31135
g28700 and n17969 n31013 ; n31136
g28701 nor n31135 n31136 ; n31137
g28702 nor n17779 n31137 ; n31138
g28703 and n17779 n31013 ; n31139
g28704 nor n31138 n31139 ; n31140
g28705 nor n17804 n31140 ; n31141
g28706 and n17804 n31013 ; n31142
g28707 nor n31141 n31142 ; n31143
g28708 and pi0644 n31143_not ; n31144
g28709 and pi0644_not n31013 ; n31145
g28710 nor pi0715 n31145 ; n31146
g28711 and n31144_not n31146 ; n31147
g28712 and pi1160 n31147_not ; n31148
g28713 and n31077_not n31148 ; n31149
g28714 and pi0644 n31075_not ; n31150
g28715 nor pi0715 n31150 ; n31151
g28716 nor pi0644 n31143 ; n31152
g28717 and pi0644 n31013 ; n31153
g28718 and pi0715 n31153_not ; n31154
g28719 and n31152_not n31154 ; n31155
g28720 nor pi1160 n31155 ; n31156
g28721 and n31151_not n31156 ; n31157
g28722 nor n31149 n31157 ; n31158
g28723 and pi0790 n31158_not ; n31159
g28724 and n17777 n31054 ; n31160
g28725 and n20570_not n31137 ; n31161
g28726 and n17776 n31058 ; n31162
g28727 nor n31160 n31162 ; n31163
g28728 and n31161_not n31163 ; n31164
g28729 and pi0792 n31164_not ; n31165
g28730 and pi0609 n31040 ; n31166
g28731 and pi0699_not n31093 ; n31167
g28732 and pi0763_not n24055 ; n31168
g28733 nor n17490 n31168 ; n31169
g28734 nor pi0039 n31169 ; n31170
g28735 nor pi0190 n31170 ; n31171
g28736 nor n17469 n30846 ; n31172
g28737 and pi0190 n31172_not ; n31173
g28738 and n6284 n31173 ; n31174
g28739 and pi0038 n31174_not ; n31175
g28740 and n31171_not n31175 ; n31176
g28741 nor pi0190 n17629 ; n31177
g28742 and pi0190 n17631_not ; n31178
g28743 and pi0763 n31178_not ; n31179
g28744 and n31177_not n31179 ; n31180
g28745 and pi0190_not n17612 ; n31181
g28746 and pi0190 n17625 ; n31182
g28747 nor pi0763 n31181 ; n31183
g28748 and n31182_not n31183 ; n31184
g28749 nor pi0039 n31180 ; n31185
g28750 and n31184_not n31185 ; n31186
g28751 and pi0190 n17605 ; n31187
g28752 nor pi0190 n17546 ; n31188
g28753 and pi0763 n31188_not ; n31189
g28754 and n31187_not n31189 ; n31190
g28755 and pi0190_not n17404 ; n31191
g28756 and pi0190 n17485 ; n31192
g28757 nor pi0763 n31192 ; n31193
g28758 and n31191_not n31193 ; n31194
g28759 and pi0039 n31190_not ; n31195
g28760 and n31194_not n31195 ; n31196
g28761 nor pi0038 n31186 ; n31197
g28762 and n31196_not n31197 ; n31198
g28763 and pi0699 n31176_not ; n31199
g28764 and n31198_not n31199 ; n31200
g28765 and n2571 n31200_not ; n31201
g28766 and n31167_not n31201 ; n31202
g28767 nor n31015 n31202 ; n31203
g28768 and pi0625_not n31203 ; n31204
g28769 and pi0625 n31095 ; n31205
g28770 nor pi1153 n31205 ; n31206
g28771 and n31204_not n31206 ; n31207
g28772 nor pi0608 n31033 ; n31208
g28773 and n31207_not n31208 ; n31209
g28774 and pi0625_not n31095 ; n31210
g28775 and pi0625 n31203 ; n31211
g28776 and pi1153 n31210_not ; n31212
g28777 and n31211_not n31212 ; n31213
g28778 and pi0608 n31037_not ; n31214
g28779 and n31213_not n31214 ; n31215
g28780 nor n31209 n31215 ; n31216
g28781 and pi0778 n31216_not ; n31217
g28782 and pi0778_not n31203 ; n31218
g28783 nor n31217 n31218 ; n31219
g28784 nor pi0609 n31219 ; n31220
g28785 nor pi1155 n31166 ; n31221
g28786 and n31220_not n31221 ; n31222
g28787 nor pi0660 n31103 ; n31223
g28788 and n31222_not n31223 ; n31224
g28789 and pi0609_not n31040 ; n31225
g28790 and pi0609 n31219_not ; n31226
g28791 and pi1155 n31225_not ; n31227
g28792 and n31226_not n31227 ; n31228
g28793 and pi0660 n31107_not ; n31229
g28794 and n31228_not n31229 ; n31230
g28795 nor n31224 n31230 ; n31231
g28796 and pi0785 n31231_not ; n31232
g28797 nor pi0785 n31219 ; n31233
g28798 nor n31232 n31233 ; n31234
g28799 nor pi0618 n31234 ; n31235
g28800 and pi0618 n31043 ; n31236
g28801 nor pi1154 n31236 ; n31237
g28802 and n31235_not n31237 ; n31238
g28803 nor pi0627 n31115 ; n31239
g28804 and n31238_not n31239 ; n31240
g28805 and pi0618_not n31043 ; n31241
g28806 and pi0618 n31234_not ; n31242
g28807 and pi1154 n31241_not ; n31243
g28808 and n31242_not n31243 ; n31244
g28809 and pi0627 n31119_not ; n31245
g28810 and n31244_not n31245 ; n31246
g28811 nor n31240 n31246 ; n31247
g28812 and pi0781 n31247_not ; n31248
g28813 nor pi0781 n31234 ; n31249
g28814 nor n31248 n31249 ; n31250
g28815 and pi0789_not n31250 ; n31251
g28816 and pi0619 n31046_not ; n31252
g28817 nor pi0619 n31250 ; n31253
g28818 nor pi1159 n31252 ; n31254
g28819 and n31253_not n31254 ; n31255
g28820 nor pi0648 n31127 ; n31256
g28821 and n31255_not n31256 ; n31257
g28822 nor pi0619 n31046 ; n31258
g28823 and pi0619 n31250_not ; n31259
g28824 and pi1159 n31258_not ; n31260
g28825 and n31259_not n31260 ; n31261
g28826 and pi0648 n31131_not ; n31262
g28827 and n31261_not n31262 ; n31263
g28828 and pi0789 n31257_not ; n31264
g28829 and n31263_not n31264 ; n31265
g28830 and n17970 n31251_not ; n31266
g28831 and n31265_not n31266 ; n31267
g28832 and n17871 n31048 ; n31268
g28833 nor pi0626 n31134 ; n31269
g28834 and pi0626 n31013_not ; n31270
g28835 and n16629 n31270_not ; n31271
g28836 and n31269_not n31271 ; n31272
g28837 and pi0626 n31134_not ; n31273
g28838 nor pi0626 n31013 ; n31274
g28839 and n16628 n31274_not ; n31275
g28840 and n31273_not n31275 ; n31276
g28841 nor n31268 n31272 ; n31277
g28842 and n31276_not n31277 ; n31278
g28843 and pi0788 n31278_not ; n31279
g28844 nor n20364 n31279 ; n31280
g28845 and n31267_not n31280 ; n31281
g28846 nor n31165 n31281 ; n31282
g28847 nor n20206 n31282 ; n31283
g28848 and n17802 n31066 ; n31284
g28849 and n20559_not n31140 ; n31285
g28850 and n17801 n31070 ; n31286
g28851 nor n31284 n31285 ; n31287
g28852 and n31286_not n31287 ; n31288
g28853 and pi0787 n31288_not ; n31289
g28854 and pi0644_not n31156 ; n31290
g28855 and pi0644 n31148 ; n31291
g28856 and pi0790 n31290_not ; n31292
g28857 and n31291_not n31292 ; n31293
g28858 nor n31283 n31289 ; n31294
g28859 and n31293_not n31294 ; n31295
g28860 nor n31159 n31295 ; n31296
g28861 nor po1038 n31296 ; n31297
g28862 nor pi0832 n31012 ; n31298
g28863 and n31297_not n31298 ; n31299
g28864 nor n31011 n31299 ; po0347
g28865 nor pi0191 n2926 ; n31301
g28866 and pi0729 n16645 ; n31302
g28867 nor n31301 n31302 ; n31303
g28868 nor pi0778 n31303 ; n31304
g28869 and pi0625_not n31302 ; n31305
g28870 nor n31303 n31305 ; n31306
g28871 and pi1153 n31306_not ; n31307
g28872 nor pi1153 n31301 ; n31308
g28873 and n31305_not n31308 ; n31309
g28874 and pi0778 n31309_not ; n31310
g28875 and n31307_not n31310 ; n31311
g28876 nor n31304 n31311 ; n31312
g28877 nor n17845 n31312 ; n31313
g28878 and n17847_not n31313 ; n31314
g28879 and n17849_not n31314 ; n31315
g28880 and n17851_not n31315 ; n31316
g28881 and n17857_not n31316 ; n31317
g28882 and pi0647_not n31317 ; n31318
g28883 and pi0647 n31301 ; n31319
g28884 nor pi1157 n31319 ; n31320
g28885 and n31318_not n31320 ; n31321
g28886 and pi0630 n31321 ; n31322
g28887 and pi0746 n17244 ; n31323
g28888 nor n31301 n31323 ; n31324
g28889 nor n17874 n31324 ; n31325
g28890 nor pi0785 n31325 ; n31326
g28891 and n17296 n31323 ; n31327
g28892 and n31325 n31327_not ; n31328
g28893 and pi1155 n31328_not ; n31329
g28894 nor pi1155 n31301 ; n31330
g28895 and n31327_not n31330 ; n31331
g28896 nor n31329 n31331 ; n31332
g28897 and pi0785 n31332_not ; n31333
g28898 nor n31326 n31333 ; n31334
g28899 nor pi0781 n31334 ; n31335
g28900 and n17889_not n31334 ; n31336
g28901 and pi1154 n31336_not ; n31337
g28902 and n17892_not n31334 ; n31338
g28903 nor pi1154 n31338 ; n31339
g28904 nor n31337 n31339 ; n31340
g28905 and pi0781 n31340_not ; n31341
g28906 nor n31335 n31341 ; n31342
g28907 nor pi0789 n31342 ; n31343
g28908 and n23078_not n31342 ; n31344
g28909 and pi1159 n31344_not ; n31345
g28910 and n23081_not n31342 ; n31346
g28911 nor pi1159 n31346 ; n31347
g28912 nor n31345 n31347 ; n31348
g28913 and pi0789 n31348_not ; n31349
g28914 nor n31343 n31349 ; n31350
g28915 and n17969_not n31350 ; n31351
g28916 and n17969 n31301 ; n31352
g28917 nor n31351 n31352 ; n31353
g28918 nor n17779 n31353 ; n31354
g28919 and n17779 n31301 ; n31355
g28920 nor n31354 n31355 ; n31356
g28921 and n20559_not n31356 ; n31357
g28922 and pi0647 n31317_not ; n31358
g28923 nor pi0647 n31301 ; n31359
g28924 nor n31358 n31359 ; n31360
g28925 and n17801 n31360_not ; n31361
g28926 nor n31322 n31361 ; n31362
g28927 and n31357_not n31362 ; n31363
g28928 and pi0787 n31363_not ; n31364
g28929 and n17871 n31315 ; n31365
g28930 nor pi0626 n31350 ; n31366
g28931 and pi0626 n31301_not ; n31367
g28932 and n16629 n31367_not ; n31368
g28933 and n31366_not n31368 ; n31369
g28934 and pi0626 n31350_not ; n31370
g28935 nor pi0626 n31301 ; n31371
g28936 and n16628 n31371_not ; n31372
g28937 and n31370_not n31372 ; n31373
g28938 nor n31365 n31369 ; n31374
g28939 and n31373_not n31374 ; n31375
g28940 and pi0788 n31375_not ; n31376
g28941 and pi0618 n31313 ; n31377
g28942 nor n17168 n31303 ; n31378
g28943 and pi0625 n31378 ; n31379
g28944 and n31324 n31378_not ; n31380
g28945 nor n31379 n31380 ; n31381
g28946 and n31308 n31381_not ; n31382
g28947 nor pi0608 n31307 ; n31383
g28948 and n31382_not n31383 ; n31384
g28949 and pi1153 n31324 ; n31385
g28950 and n31379_not n31385 ; n31386
g28951 and pi0608 n31309_not ; n31387
g28952 and n31386_not n31387 ; n31388
g28953 nor n31384 n31388 ; n31389
g28954 and pi0778 n31389_not ; n31390
g28955 nor pi0778 n31380 ; n31391
g28956 nor n31390 n31391 ; n31392
g28957 nor pi0609 n31392 ; n31393
g28958 and pi0609 n31312_not ; n31394
g28959 nor pi1155 n31394 ; n31395
g28960 and n31393_not n31395 ; n31396
g28961 nor pi0660 n31329 ; n31397
g28962 and n31396_not n31397 ; n31398
g28963 and pi0609 n31392_not ; n31399
g28964 nor pi0609 n31312 ; n31400
g28965 and pi1155 n31400_not ; n31401
g28966 and n31399_not n31401 ; n31402
g28967 and pi0660 n31331_not ; n31403
g28968 and n31402_not n31403 ; n31404
g28969 nor n31398 n31404 ; n31405
g28970 and pi0785 n31405_not ; n31406
g28971 nor pi0785 n31392 ; n31407
g28972 nor n31406 n31407 ; n31408
g28973 nor pi0618 n31408 ; n31409
g28974 nor pi1154 n31377 ; n31410
g28975 and n31409_not n31410 ; n31411
g28976 nor pi0627 n31337 ; n31412
g28977 and n31411_not n31412 ; n31413
g28978 and pi0618_not n31313 ; n31414
g28979 and pi0618 n31408_not ; n31415
g28980 and pi1154 n31414_not ; n31416
g28981 and n31415_not n31416 ; n31417
g28982 and pi0627 n31339_not ; n31418
g28983 and n31417_not n31418 ; n31419
g28984 nor n31413 n31419 ; n31420
g28985 and pi0781 n31420_not ; n31421
g28986 nor pi0781 n31408 ; n31422
g28987 nor n31421 n31422 ; n31423
g28988 and pi0789_not n31423 ; n31424
g28989 nor pi0619 n31423 ; n31425
g28990 and pi0619 n31314 ; n31426
g28991 nor pi1159 n31426 ; n31427
g28992 and n31425_not n31427 ; n31428
g28993 nor pi0648 n31345 ; n31429
g28994 and n31428_not n31429 ; n31430
g28995 and pi0619 n31423_not ; n31431
g28996 and pi0619_not n31314 ; n31432
g28997 and pi1159 n31432_not ; n31433
g28998 and n31431_not n31433 ; n31434
g28999 and pi0648 n31347_not ; n31435
g29000 and n31434_not n31435 ; n31436
g29001 and pi0789 n31430_not ; n31437
g29002 and n31436_not n31437 ; n31438
g29003 and n17970 n31424_not ; n31439
g29004 and n31438_not n31439 ; n31440
g29005 nor n31376 n31440 ; n31441
g29006 nor n20364 n31441 ; n31442
g29007 and n17854 n31353_not ; n31443
g29008 and n20851 n31316 ; n31444
g29009 nor n31443 n31444 ; n31445
g29010 nor pi0629 n31445 ; n31446
g29011 and n20855 n31316 ; n31447
g29012 and n17853 n31353_not ; n31448
g29013 nor n31447 n31448 ; n31449
g29014 and pi0629 n31449_not ; n31450
g29015 nor n31446 n31450 ; n31451
g29016 and pi0792 n31451_not ; n31452
g29017 nor n20206 n31452 ; n31453
g29018 and n31442_not n31453 ; n31454
g29019 nor n31364 n31454 ; n31455
g29020 and pi0790_not n31455 ; n31456
g29021 nor pi0787 n31317 ; n31457
g29022 and pi1157 n31360_not ; n31458
g29023 nor n31321 n31458 ; n31459
g29024 and pi0787 n31459_not ; n31460
g29025 nor n31457 n31460 ; n31461
g29026 and pi0644_not n31461 ; n31462
g29027 and pi0644 n31455 ; n31463
g29028 and pi0715 n31462_not ; n31464
g29029 and n31463_not n31464 ; n31465
g29030 nor n17804 n31356 ; n31466
g29031 and n17804 n31301 ; n31467
g29032 nor n31466 n31467 ; n31468
g29033 and pi0644 n31468_not ; n31469
g29034 and pi0644_not n31301 ; n31470
g29035 nor pi0715 n31470 ; n31471
g29036 and n31469_not n31471 ; n31472
g29037 and pi1160 n31472_not ; n31473
g29038 and n31465_not n31473 ; n31474
g29039 nor pi0644 n31468 ; n31475
g29040 and pi0644 n31301 ; n31476
g29041 and pi0715 n31476_not ; n31477
g29042 and n31475_not n31477 ; n31478
g29043 and pi0644 n31461 ; n31479
g29044 and pi0644_not n31455 ; n31480
g29045 nor pi0715 n31479 ; n31481
g29046 and n31480_not n31481 ; n31482
g29047 nor pi1160 n31478 ; n31483
g29048 and n31482_not n31483 ; n31484
g29049 nor n31474 n31484 ; n31485
g29050 and pi0790 n31485_not ; n31486
g29051 and pi0832 n31456_not ; n31487
g29052 and n31486_not n31487 ; n31488
g29053 and pi0191_not po1038 ; n31489
g29054 nor pi0191 n17059 ; n31490
g29055 and n16635 n31490_not ; n31491
g29056 and pi0191 n2571_not ; n31492
g29057 nor pi0191 n16641 ; n31493
g29058 and n16647 n31493_not ; n31494
g29059 and pi0191_not n18072 ; n31495
g29060 and pi0191 n18076_not ; n31496
g29061 nor pi0038 n31496 ; n31497
g29062 and n31495_not n31497 ; n31498
g29063 and pi0729 n31494_not ; n31499
g29064 and n31498_not n31499 ; n31500
g29065 nor pi0191 pi0729 ; n31501
g29066 and n17052_not n31501 ; n31502
g29067 and n2571 n31502_not ; n31503
g29068 and n31500_not n31503 ; n31504
g29069 nor n31492 n31504 ; n31505
g29070 nor pi0778 n31505 ; n31506
g29071 and pi0625_not n31490 ; n31507
g29072 and pi0625 n31505 ; n31508
g29073 and pi1153 n31507_not ; n31509
g29074 and n31508_not n31509 ; n31510
g29075 and pi0625_not n31505 ; n31511
g29076 and pi0625 n31490 ; n31512
g29077 nor pi1153 n31512 ; n31513
g29078 and n31511_not n31513 ; n31514
g29079 nor n31510 n31514 ; n31515
g29080 and pi0778 n31515_not ; n31516
g29081 nor n31506 n31516 ; n31517
g29082 nor n17075 n31517 ; n31518
g29083 and n17075 n31490_not ; n31519
g29084 nor n31518 n31519 ; n31520
g29085 and n16639_not n31520 ; n31521
g29086 and n16639 n31490 ; n31522
g29087 nor n31521 n31522 ; n31523
g29088 and n16635_not n31523 ; n31524
g29089 nor n31491 n31524 ; n31525
g29090 and n16631_not n31525 ; n31526
g29091 and n16631 n31490 ; n31527
g29092 nor n31526 n31527 ; n31528
g29093 nor pi0628 n31528 ; n31529
g29094 and pi0628 n31490 ; n31530
g29095 nor n31529 n31530 ; n31531
g29096 nor pi1156 n31531 ; n31532
g29097 and pi0628 n31528_not ; n31533
g29098 and pi0628_not n31490 ; n31534
g29099 nor n31533 n31534 ; n31535
g29100 and pi1156 n31535_not ; n31536
g29101 nor n31532 n31536 ; n31537
g29102 and pi0792 n31537_not ; n31538
g29103 nor pi0792 n31528 ; n31539
g29104 nor n31538 n31539 ; n31540
g29105 nor pi0647 n31540 ; n31541
g29106 and pi0647 n31490 ; n31542
g29107 nor n31541 n31542 ; n31543
g29108 nor pi1157 n31543 ; n31544
g29109 and pi0647 n31540_not ; n31545
g29110 and pi0647_not n31490 ; n31546
g29111 nor n31545 n31546 ; n31547
g29112 and pi1157 n31547_not ; n31548
g29113 nor n31544 n31548 ; n31549
g29114 and pi0787 n31549_not ; n31550
g29115 nor pi0787 n31540 ; n31551
g29116 nor n31550 n31551 ; n31552
g29117 nor pi0644 n31552 ; n31553
g29118 and pi0715 n31553_not ; n31554
g29119 and pi0746_not n17046 ; n31555
g29120 and pi0191 n17273 ; n31556
g29121 nor n31555 n31556 ; n31557
g29122 and pi0039 n31557_not ; n31558
g29123 and pi0746 n17234_not ; n31559
g29124 and pi0191 n31559_not ; n31560
g29125 and pi0191_not pi0746 ; n31561
g29126 and n17221 n31561 ; n31562
g29127 nor n22439 n31560 ; n31563
g29128 and n31562_not n31563 ; n31564
g29129 and n31558_not n31564 ; n31565
g29130 nor pi0038 n31565 ; n31566
g29131 and pi0746 n17280 ; n31567
g29132 and pi0038 n31493_not ; n31568
g29133 and n31567_not n31568 ; n31569
g29134 nor n31566 n31569 ; n31570
g29135 and n2571 n31570_not ; n31571
g29136 nor n31492 n31571 ; n31572
g29137 nor n17117 n31572 ; n31573
g29138 and n17117 n31490_not ; n31574
g29139 nor n31573 n31574 ; n31575
g29140 nor pi0785 n31575 ; n31576
g29141 nor n17291 n31490 ; n31577
g29142 and pi0609 n31573 ; n31578
g29143 nor n31577 n31578 ; n31579
g29144 and pi1155 n31579_not ; n31580
g29145 nor n17296 n31490 ; n31581
g29146 and pi0609_not n31573 ; n31582
g29147 nor n31581 n31582 ; n31583
g29148 nor pi1155 n31583 ; n31584
g29149 nor n31580 n31584 ; n31585
g29150 and pi0785 n31585_not ; n31586
g29151 nor n31576 n31586 ; n31587
g29152 nor pi0781 n31587 ; n31588
g29153 and pi0618_not n31490 ; n31589
g29154 and pi0618 n31587 ; n31590
g29155 and pi1154 n31589_not ; n31591
g29156 and n31590_not n31591 ; n31592
g29157 and pi0618_not n31587 ; n31593
g29158 and pi0618 n31490 ; n31594
g29159 nor pi1154 n31594 ; n31595
g29160 and n31593_not n31595 ; n31596
g29161 nor n31592 n31596 ; n31597
g29162 and pi0781 n31597_not ; n31598
g29163 nor n31588 n31598 ; n31599
g29164 nor pi0789 n31599 ; n31600
g29165 and pi0619_not n31490 ; n31601
g29166 and pi0619 n31599 ; n31602
g29167 and pi1159 n31601_not ; n31603
g29168 and n31602_not n31603 ; n31604
g29169 and pi0619_not n31599 ; n31605
g29170 and pi0619 n31490 ; n31606
g29171 nor pi1159 n31606 ; n31607
g29172 and n31605_not n31607 ; n31608
g29173 nor n31604 n31608 ; n31609
g29174 and pi0789 n31609_not ; n31610
g29175 nor n31600 n31610 ; n31611
g29176 and n17969_not n31611 ; n31612
g29177 and n17969 n31490 ; n31613
g29178 nor n31612 n31613 ; n31614
g29179 nor n17779 n31614 ; n31615
g29180 and n17779 n31490 ; n31616
g29181 nor n31615 n31616 ; n31617
g29182 nor n17804 n31617 ; n31618
g29183 and n17804 n31490 ; n31619
g29184 nor n31618 n31619 ; n31620
g29185 and pi0644 n31620_not ; n31621
g29186 and pi0644_not n31490 ; n31622
g29187 nor pi0715 n31622 ; n31623
g29188 and n31621_not n31623 ; n31624
g29189 and pi1160 n31624_not ; n31625
g29190 and n31554_not n31625 ; n31626
g29191 and pi0644 n31552_not ; n31627
g29192 nor pi0715 n31627 ; n31628
g29193 nor pi0644 n31620 ; n31629
g29194 and pi0644 n31490 ; n31630
g29195 and pi0715 n31630_not ; n31631
g29196 and n31629_not n31631 ; n31632
g29197 nor pi1160 n31632 ; n31633
g29198 and n31628_not n31633 ; n31634
g29199 nor n31626 n31634 ; n31635
g29200 and pi0790 n31635_not ; n31636
g29201 and n17777 n31531 ; n31637
g29202 and n20570_not n31614 ; n31638
g29203 and n17776 n31535 ; n31639
g29204 nor n31637 n31639 ; n31640
g29205 and n31638_not n31640 ; n31641
g29206 and pi0792 n31641_not ; n31642
g29207 and pi0609 n31517 ; n31643
g29208 and pi0729_not n31570 ; n31644
g29209 and pi0746_not n24055 ; n31645
g29210 nor n17490 n31645 ; n31646
g29211 nor pi0039 n31646 ; n31647
g29212 nor pi0191 n31647 ; n31648
g29213 nor n17469 n31323 ; n31649
g29214 and pi0191 n31649_not ; n31650
g29215 and n6284 n31650 ; n31651
g29216 and pi0038 n31651_not ; n31652
g29217 and n31648_not n31652 ; n31653
g29218 nor pi0191 n17629 ; n31654
g29219 and pi0191 n17631_not ; n31655
g29220 and pi0746 n31655_not ; n31656
g29221 and n31654_not n31656 ; n31657
g29222 and pi0191_not n17612 ; n31658
g29223 and pi0191 n17625 ; n31659
g29224 nor pi0746 n31658 ; n31660
g29225 and n31659_not n31660 ; n31661
g29226 nor pi0039 n31657 ; n31662
g29227 and n31661_not n31662 ; n31663
g29228 and pi0191 n17605 ; n31664
g29229 nor pi0191 n17546 ; n31665
g29230 and pi0746 n31665_not ; n31666
g29231 and n31664_not n31666 ; n31667
g29232 and pi0191_not n17404 ; n31668
g29233 and pi0191 n17485 ; n31669
g29234 nor pi0746 n31669 ; n31670
g29235 and n31668_not n31670 ; n31671
g29236 and pi0039 n31667_not ; n31672
g29237 and n31671_not n31672 ; n31673
g29238 nor pi0038 n31663 ; n31674
g29239 and n31673_not n31674 ; n31675
g29240 and pi0729 n31653_not ; n31676
g29241 and n31675_not n31676 ; n31677
g29242 and n2571 n31677_not ; n31678
g29243 and n31644_not n31678 ; n31679
g29244 nor n31492 n31679 ; n31680
g29245 and pi0625_not n31680 ; n31681
g29246 and pi0625 n31572 ; n31682
g29247 nor pi1153 n31682 ; n31683
g29248 and n31681_not n31683 ; n31684
g29249 nor pi0608 n31510 ; n31685
g29250 and n31684_not n31685 ; n31686
g29251 and pi0625_not n31572 ; n31687
g29252 and pi0625 n31680 ; n31688
g29253 and pi1153 n31687_not ; n31689
g29254 and n31688_not n31689 ; n31690
g29255 and pi0608 n31514_not ; n31691
g29256 and n31690_not n31691 ; n31692
g29257 nor n31686 n31692 ; n31693
g29258 and pi0778 n31693_not ; n31694
g29259 and pi0778_not n31680 ; n31695
g29260 nor n31694 n31695 ; n31696
g29261 nor pi0609 n31696 ; n31697
g29262 nor pi1155 n31643 ; n31698
g29263 and n31697_not n31698 ; n31699
g29264 nor pi0660 n31580 ; n31700
g29265 and n31699_not n31700 ; n31701
g29266 and pi0609_not n31517 ; n31702
g29267 and pi0609 n31696_not ; n31703
g29268 and pi1155 n31702_not ; n31704
g29269 and n31703_not n31704 ; n31705
g29270 and pi0660 n31584_not ; n31706
g29271 and n31705_not n31706 ; n31707
g29272 nor n31701 n31707 ; n31708
g29273 and pi0785 n31708_not ; n31709
g29274 nor pi0785 n31696 ; n31710
g29275 nor n31709 n31710 ; n31711
g29276 nor pi0618 n31711 ; n31712
g29277 and pi0618 n31520 ; n31713
g29278 nor pi1154 n31713 ; n31714
g29279 and n31712_not n31714 ; n31715
g29280 nor pi0627 n31592 ; n31716
g29281 and n31715_not n31716 ; n31717
g29282 and pi0618_not n31520 ; n31718
g29283 and pi0618 n31711_not ; n31719
g29284 and pi1154 n31718_not ; n31720
g29285 and n31719_not n31720 ; n31721
g29286 and pi0627 n31596_not ; n31722
g29287 and n31721_not n31722 ; n31723
g29288 nor n31717 n31723 ; n31724
g29289 and pi0781 n31724_not ; n31725
g29290 nor pi0781 n31711 ; n31726
g29291 nor n31725 n31726 ; n31727
g29292 and pi0789_not n31727 ; n31728
g29293 and pi0619 n31523_not ; n31729
g29294 nor pi0619 n31727 ; n31730
g29295 nor pi1159 n31729 ; n31731
g29296 and n31730_not n31731 ; n31732
g29297 nor pi0648 n31604 ; n31733
g29298 and n31732_not n31733 ; n31734
g29299 nor pi0619 n31523 ; n31735
g29300 and pi0619 n31727_not ; n31736
g29301 and pi1159 n31735_not ; n31737
g29302 and n31736_not n31737 ; n31738
g29303 and pi0648 n31608_not ; n31739
g29304 and n31738_not n31739 ; n31740
g29305 and pi0789 n31734_not ; n31741
g29306 and n31740_not n31741 ; n31742
g29307 and n17970 n31728_not ; n31743
g29308 and n31742_not n31743 ; n31744
g29309 and n17871 n31525 ; n31745
g29310 nor pi0626 n31611 ; n31746
g29311 and pi0626 n31490_not ; n31747
g29312 and n16629 n31747_not ; n31748
g29313 and n31746_not n31748 ; n31749
g29314 and pi0626 n31611_not ; n31750
g29315 nor pi0626 n31490 ; n31751
g29316 and n16628 n31751_not ; n31752
g29317 and n31750_not n31752 ; n31753
g29318 nor n31745 n31749 ; n31754
g29319 and n31753_not n31754 ; n31755
g29320 and pi0788 n31755_not ; n31756
g29321 nor n20364 n31756 ; n31757
g29322 and n31744_not n31757 ; n31758
g29323 nor n31642 n31758 ; n31759
g29324 nor n20206 n31759 ; n31760
g29325 and n17802 n31543 ; n31761
g29326 and n20559_not n31617 ; n31762
g29327 and n17801 n31547 ; n31763
g29328 nor n31761 n31762 ; n31764
g29329 and n31763_not n31764 ; n31765
g29330 and pi0787 n31765_not ; n31766
g29331 and pi0644_not n31633 ; n31767
g29332 and pi0644 n31625 ; n31768
g29333 and pi0790 n31767_not ; n31769
g29334 and n31768_not n31769 ; n31770
g29335 nor n31760 n31766 ; n31771
g29336 and n31770_not n31771 ; n31772
g29337 nor n31636 n31772 ; n31773
g29338 nor po1038 n31773 ; n31774
g29339 nor pi0832 n31489 ; n31775
g29340 and n31774_not n31775 ; n31776
g29341 nor n31488 n31776 ; po0348
g29342 nor pi0192 n2926 ; n31778
g29343 and pi0691 n16645 ; n31779
g29344 nor n31778 n31779 ; n31780
g29345 nor pi0778 n31780 ; n31781
g29346 and pi0625_not n31779 ; n31782
g29347 nor n31780 n31782 ; n31783
g29348 and pi1153 n31783_not ; n31784
g29349 nor pi1153 n31778 ; n31785
g29350 and n31782_not n31785 ; n31786
g29351 and pi0778 n31786_not ; n31787
g29352 and n31784_not n31787 ; n31788
g29353 nor n31781 n31788 ; n31789
g29354 nor n17845 n31789 ; n31790
g29355 and n17847_not n31790 ; n31791
g29356 and n17849_not n31791 ; n31792
g29357 and n17851_not n31792 ; n31793
g29358 and n17857_not n31793 ; n31794
g29359 and pi0647_not n31794 ; n31795
g29360 and pi0647 n31778 ; n31796
g29361 nor pi1157 n31796 ; n31797
g29362 and n31795_not n31797 ; n31798
g29363 and pi0630 n31798 ; n31799
g29364 and pi0764 n17244 ; n31800
g29365 nor n31778 n31800 ; n31801
g29366 nor n17874 n31801 ; n31802
g29367 nor pi0785 n31802 ; n31803
g29368 and n17296 n31800 ; n31804
g29369 and n31802 n31804_not ; n31805
g29370 and pi1155 n31805_not ; n31806
g29371 nor pi1155 n31778 ; n31807
g29372 and n31804_not n31807 ; n31808
g29373 nor n31806 n31808 ; n31809
g29374 and pi0785 n31809_not ; n31810
g29375 nor n31803 n31810 ; n31811
g29376 nor pi0781 n31811 ; n31812
g29377 and n17889_not n31811 ; n31813
g29378 and pi1154 n31813_not ; n31814
g29379 and n17892_not n31811 ; n31815
g29380 nor pi1154 n31815 ; n31816
g29381 nor n31814 n31816 ; n31817
g29382 and pi0781 n31817_not ; n31818
g29383 nor n31812 n31818 ; n31819
g29384 nor pi0789 n31819 ; n31820
g29385 and n23078_not n31819 ; n31821
g29386 and pi1159 n31821_not ; n31822
g29387 and n23081_not n31819 ; n31823
g29388 nor pi1159 n31823 ; n31824
g29389 nor n31822 n31824 ; n31825
g29390 and pi0789 n31825_not ; n31826
g29391 nor n31820 n31826 ; n31827
g29392 and n17969_not n31827 ; n31828
g29393 and n17969 n31778 ; n31829
g29394 nor n31828 n31829 ; n31830
g29395 nor n17779 n31830 ; n31831
g29396 and n17779 n31778 ; n31832
g29397 nor n31831 n31832 ; n31833
g29398 and n20559_not n31833 ; n31834
g29399 and pi0647 n31794_not ; n31835
g29400 nor pi0647 n31778 ; n31836
g29401 nor n31835 n31836 ; n31837
g29402 and n17801 n31837_not ; n31838
g29403 nor n31799 n31838 ; n31839
g29404 and n31834_not n31839 ; n31840
g29405 and pi0787 n31840_not ; n31841
g29406 and n17871 n31792 ; n31842
g29407 nor pi0626 n31827 ; n31843
g29408 and pi0626 n31778_not ; n31844
g29409 and n16629 n31844_not ; n31845
g29410 and n31843_not n31845 ; n31846
g29411 and pi0626 n31827_not ; n31847
g29412 nor pi0626 n31778 ; n31848
g29413 and n16628 n31848_not ; n31849
g29414 and n31847_not n31849 ; n31850
g29415 nor n31842 n31846 ; n31851
g29416 and n31850_not n31851 ; n31852
g29417 and pi0788 n31852_not ; n31853
g29418 and pi0618 n31790 ; n31854
g29419 nor n17168 n31780 ; n31855
g29420 and pi0625 n31855 ; n31856
g29421 and n31801 n31855_not ; n31857
g29422 nor n31856 n31857 ; n31858
g29423 and n31785 n31858_not ; n31859
g29424 nor pi0608 n31784 ; n31860
g29425 and n31859_not n31860 ; n31861
g29426 and pi1153 n31801 ; n31862
g29427 and n31856_not n31862 ; n31863
g29428 and pi0608 n31786_not ; n31864
g29429 and n31863_not n31864 ; n31865
g29430 nor n31861 n31865 ; n31866
g29431 and pi0778 n31866_not ; n31867
g29432 nor pi0778 n31857 ; n31868
g29433 nor n31867 n31868 ; n31869
g29434 nor pi0609 n31869 ; n31870
g29435 and pi0609 n31789_not ; n31871
g29436 nor pi1155 n31871 ; n31872
g29437 and n31870_not n31872 ; n31873
g29438 nor pi0660 n31806 ; n31874
g29439 and n31873_not n31874 ; n31875
g29440 and pi0609 n31869_not ; n31876
g29441 nor pi0609 n31789 ; n31877
g29442 and pi1155 n31877_not ; n31878
g29443 and n31876_not n31878 ; n31879
g29444 and pi0660 n31808_not ; n31880
g29445 and n31879_not n31880 ; n31881
g29446 nor n31875 n31881 ; n31882
g29447 and pi0785 n31882_not ; n31883
g29448 nor pi0785 n31869 ; n31884
g29449 nor n31883 n31884 ; n31885
g29450 nor pi0618 n31885 ; n31886
g29451 nor pi1154 n31854 ; n31887
g29452 and n31886_not n31887 ; n31888
g29453 nor pi0627 n31814 ; n31889
g29454 and n31888_not n31889 ; n31890
g29455 and pi0618_not n31790 ; n31891
g29456 and pi0618 n31885_not ; n31892
g29457 and pi1154 n31891_not ; n31893
g29458 and n31892_not n31893 ; n31894
g29459 and pi0627 n31816_not ; n31895
g29460 and n31894_not n31895 ; n31896
g29461 nor n31890 n31896 ; n31897
g29462 and pi0781 n31897_not ; n31898
g29463 nor pi0781 n31885 ; n31899
g29464 nor n31898 n31899 ; n31900
g29465 and pi0789_not n31900 ; n31901
g29466 nor pi0619 n31900 ; n31902
g29467 and pi0619 n31791 ; n31903
g29468 nor pi1159 n31903 ; n31904
g29469 and n31902_not n31904 ; n31905
g29470 nor pi0648 n31822 ; n31906
g29471 and n31905_not n31906 ; n31907
g29472 and pi0619 n31900_not ; n31908
g29473 and pi0619_not n31791 ; n31909
g29474 and pi1159 n31909_not ; n31910
g29475 and n31908_not n31910 ; n31911
g29476 and pi0648 n31824_not ; n31912
g29477 and n31911_not n31912 ; n31913
g29478 and pi0789 n31907_not ; n31914
g29479 and n31913_not n31914 ; n31915
g29480 and n17970 n31901_not ; n31916
g29481 and n31915_not n31916 ; n31917
g29482 nor n31853 n31917 ; n31918
g29483 nor n20364 n31918 ; n31919
g29484 and n17854 n31830_not ; n31920
g29485 and n20851 n31793 ; n31921
g29486 nor n31920 n31921 ; n31922
g29487 nor pi0629 n31922 ; n31923
g29488 and n20855 n31793 ; n31924
g29489 and n17853 n31830_not ; n31925
g29490 nor n31924 n31925 ; n31926
g29491 and pi0629 n31926_not ; n31927
g29492 nor n31923 n31927 ; n31928
g29493 and pi0792 n31928_not ; n31929
g29494 nor n20206 n31929 ; n31930
g29495 and n31919_not n31930 ; n31931
g29496 nor n31841 n31931 ; n31932
g29497 and pi0790_not n31932 ; n31933
g29498 nor pi0787 n31794 ; n31934
g29499 and pi1157 n31837_not ; n31935
g29500 nor n31798 n31935 ; n31936
g29501 and pi0787 n31936_not ; n31937
g29502 nor n31934 n31937 ; n31938
g29503 and pi0644_not n31938 ; n31939
g29504 and pi0644 n31932 ; n31940
g29505 and pi0715 n31939_not ; n31941
g29506 and n31940_not n31941 ; n31942
g29507 nor n17804 n31833 ; n31943
g29508 and n17804 n31778 ; n31944
g29509 nor n31943 n31944 ; n31945
g29510 and pi0644 n31945_not ; n31946
g29511 and pi0644_not n31778 ; n31947
g29512 nor pi0715 n31947 ; n31948
g29513 and n31946_not n31948 ; n31949
g29514 and pi1160 n31949_not ; n31950
g29515 and n31942_not n31950 ; n31951
g29516 nor pi0644 n31945 ; n31952
g29517 and pi0644 n31778 ; n31953
g29518 and pi0715 n31953_not ; n31954
g29519 and n31952_not n31954 ; n31955
g29520 and pi0644 n31938 ; n31956
g29521 and pi0644_not n31932 ; n31957
g29522 nor pi0715 n31956 ; n31958
g29523 and n31957_not n31958 ; n31959
g29524 nor pi1160 n31955 ; n31960
g29525 and n31959_not n31960 ; n31961
g29526 nor n31951 n31961 ; n31962
g29527 and pi0790 n31962_not ; n31963
g29528 and pi0832 n31933_not ; n31964
g29529 and n31963_not n31964 ; n31965
g29530 and pi0192_not po1038 ; n31966
g29531 nor pi0192 n17059 ; n31967
g29532 and n16635 n31967_not ; n31968
g29533 and pi0192 n2571_not ; n31969
g29534 nor pi0192 n16641 ; n31970
g29535 and n16647 n31970_not ; n31971
g29536 and pi0192_not n18072 ; n31972
g29537 and pi0192 n18076_not ; n31973
g29538 nor pi0038 n31973 ; n31974
g29539 and n31972_not n31974 ; n31975
g29540 and pi0691 n31971_not ; n31976
g29541 and n31975_not n31976 ; n31977
g29542 nor pi0192 pi0691 ; n31978
g29543 and n17052_not n31978 ; n31979
g29544 and n2571 n31979_not ; n31980
g29545 and n31977_not n31980 ; n31981
g29546 nor n31969 n31981 ; n31982
g29547 nor pi0778 n31982 ; n31983
g29548 and pi0625_not n31967 ; n31984
g29549 and pi0625 n31982 ; n31985
g29550 and pi1153 n31984_not ; n31986
g29551 and n31985_not n31986 ; n31987
g29552 and pi0625_not n31982 ; n31988
g29553 and pi0625 n31967 ; n31989
g29554 nor pi1153 n31989 ; n31990
g29555 and n31988_not n31990 ; n31991
g29556 nor n31987 n31991 ; n31992
g29557 and pi0778 n31992_not ; n31993
g29558 nor n31983 n31993 ; n31994
g29559 nor n17075 n31994 ; n31995
g29560 and n17075 n31967_not ; n31996
g29561 nor n31995 n31996 ; n31997
g29562 and n16639_not n31997 ; n31998
g29563 and n16639 n31967 ; n31999
g29564 nor n31998 n31999 ; n32000
g29565 and n16635_not n32000 ; n32001
g29566 nor n31968 n32001 ; n32002
g29567 and n16631_not n32002 ; n32003
g29568 and n16631 n31967 ; n32004
g29569 nor n32003 n32004 ; n32005
g29570 nor pi0628 n32005 ; n32006
g29571 and pi0628 n31967 ; n32007
g29572 nor n32006 n32007 ; n32008
g29573 nor pi1156 n32008 ; n32009
g29574 and pi0628 n32005_not ; n32010
g29575 and pi0628_not n31967 ; n32011
g29576 nor n32010 n32011 ; n32012
g29577 and pi1156 n32012_not ; n32013
g29578 nor n32009 n32013 ; n32014
g29579 and pi0792 n32014_not ; n32015
g29580 nor pi0792 n32005 ; n32016
g29581 nor n32015 n32016 ; n32017
g29582 nor pi0647 n32017 ; n32018
g29583 and pi0647 n31967 ; n32019
g29584 nor n32018 n32019 ; n32020
g29585 nor pi1157 n32020 ; n32021
g29586 and pi0647 n32017_not ; n32022
g29587 and pi0647_not n31967 ; n32023
g29588 nor n32022 n32023 ; n32024
g29589 and pi1157 n32024_not ; n32025
g29590 nor n32021 n32025 ; n32026
g29591 and pi0787 n32026_not ; n32027
g29592 nor pi0787 n32017 ; n32028
g29593 nor n32027 n32028 ; n32029
g29594 nor pi0644 n32029 ; n32030
g29595 and pi0715 n32030_not ; n32031
g29596 and pi0764_not n17046 ; n32032
g29597 and pi0192 n17273 ; n32033
g29598 nor n32032 n32033 ; n32034
g29599 and pi0039 n32034_not ; n32035
g29600 and pi0764 n17234_not ; n32036
g29601 and pi0192 n32036_not ; n32037
g29602 and pi0192_not pi0764 ; n32038
g29603 and n17221 n32038 ; n32039
g29604 nor n22600 n32037 ; n32040
g29605 and n32039_not n32040 ; n32041
g29606 and n32035_not n32041 ; n32042
g29607 nor pi0038 n32042 ; n32043
g29608 and pi0764 n17280 ; n32044
g29609 and pi0038 n31970_not ; n32045
g29610 and n32044_not n32045 ; n32046
g29611 nor n32043 n32046 ; n32047
g29612 and n2571 n32047_not ; n32048
g29613 nor n31969 n32048 ; n32049
g29614 nor n17117 n32049 ; n32050
g29615 and n17117 n31967_not ; n32051
g29616 nor n32050 n32051 ; n32052
g29617 nor pi0785 n32052 ; n32053
g29618 nor n17291 n31967 ; n32054
g29619 and pi0609 n32050 ; n32055
g29620 nor n32054 n32055 ; n32056
g29621 and pi1155 n32056_not ; n32057
g29622 nor n17296 n31967 ; n32058
g29623 and pi0609_not n32050 ; n32059
g29624 nor n32058 n32059 ; n32060
g29625 nor pi1155 n32060 ; n32061
g29626 nor n32057 n32061 ; n32062
g29627 and pi0785 n32062_not ; n32063
g29628 nor n32053 n32063 ; n32064
g29629 nor pi0781 n32064 ; n32065
g29630 and pi0618_not n31967 ; n32066
g29631 and pi0618 n32064 ; n32067
g29632 and pi1154 n32066_not ; n32068
g29633 and n32067_not n32068 ; n32069
g29634 and pi0618_not n32064 ; n32070
g29635 and pi0618 n31967 ; n32071
g29636 nor pi1154 n32071 ; n32072
g29637 and n32070_not n32072 ; n32073
g29638 nor n32069 n32073 ; n32074
g29639 and pi0781 n32074_not ; n32075
g29640 nor n32065 n32075 ; n32076
g29641 nor pi0789 n32076 ; n32077
g29642 and pi0619_not n31967 ; n32078
g29643 and pi0619 n32076 ; n32079
g29644 and pi1159 n32078_not ; n32080
g29645 and n32079_not n32080 ; n32081
g29646 and pi0619_not n32076 ; n32082
g29647 and pi0619 n31967 ; n32083
g29648 nor pi1159 n32083 ; n32084
g29649 and n32082_not n32084 ; n32085
g29650 nor n32081 n32085 ; n32086
g29651 and pi0789 n32086_not ; n32087
g29652 nor n32077 n32087 ; n32088
g29653 and n17969_not n32088 ; n32089
g29654 and n17969 n31967 ; n32090
g29655 nor n32089 n32090 ; n32091
g29656 nor n17779 n32091 ; n32092
g29657 and n17779 n31967 ; n32093
g29658 nor n32092 n32093 ; n32094
g29659 nor n17804 n32094 ; n32095
g29660 and n17804 n31967 ; n32096
g29661 nor n32095 n32096 ; n32097
g29662 and pi0644 n32097_not ; n32098
g29663 and pi0644_not n31967 ; n32099
g29664 nor pi0715 n32099 ; n32100
g29665 and n32098_not n32100 ; n32101
g29666 and pi1160 n32101_not ; n32102
g29667 and n32031_not n32102 ; n32103
g29668 and pi0644 n32029_not ; n32104
g29669 nor pi0715 n32104 ; n32105
g29670 nor pi0644 n32097 ; n32106
g29671 and pi0644 n31967 ; n32107
g29672 and pi0715 n32107_not ; n32108
g29673 and n32106_not n32108 ; n32109
g29674 nor pi1160 n32109 ; n32110
g29675 and n32105_not n32110 ; n32111
g29676 nor n32103 n32111 ; n32112
g29677 and pi0790 n32112_not ; n32113
g29678 and n17777 n32008 ; n32114
g29679 and n20570_not n32091 ; n32115
g29680 and n17776 n32012 ; n32116
g29681 nor n32114 n32116 ; n32117
g29682 and n32115_not n32117 ; n32118
g29683 and pi0792 n32118_not ; n32119
g29684 and pi0609 n31994 ; n32120
g29685 and pi0691_not n32047 ; n32121
g29686 and pi0764_not n24055 ; n32122
g29687 nor n17490 n32122 ; n32123
g29688 nor pi0039 n32123 ; n32124
g29689 nor pi0192 n32124 ; n32125
g29690 nor n17469 n31800 ; n32126
g29691 and pi0192 n32126_not ; n32127
g29692 and n6284 n32127 ; n32128
g29693 and pi0038 n32128_not ; n32129
g29694 and n32125_not n32129 ; n32130
g29695 nor pi0192 n17629 ; n32131
g29696 and pi0192 n17631_not ; n32132
g29697 and pi0764 n32132_not ; n32133
g29698 and n32131_not n32133 ; n32134
g29699 and pi0192_not n17612 ; n32135
g29700 and pi0192 n17625 ; n32136
g29701 nor pi0764 n32135 ; n32137
g29702 and n32136_not n32137 ; n32138
g29703 nor pi0039 n32134 ; n32139
g29704 and n32138_not n32139 ; n32140
g29705 and pi0192 n17605 ; n32141
g29706 nor pi0192 n17546 ; n32142
g29707 and pi0764 n32142_not ; n32143
g29708 and n32141_not n32143 ; n32144
g29709 and pi0192_not n17404 ; n32145
g29710 and pi0192 n17485 ; n32146
g29711 nor pi0764 n32146 ; n32147
g29712 and n32145_not n32147 ; n32148
g29713 and pi0039 n32144_not ; n32149
g29714 and n32148_not n32149 ; n32150
g29715 nor pi0038 n32140 ; n32151
g29716 and n32150_not n32151 ; n32152
g29717 and pi0691 n32130_not ; n32153
g29718 and n32152_not n32153 ; n32154
g29719 and n2571 n32154_not ; n32155
g29720 and n32121_not n32155 ; n32156
g29721 nor n31969 n32156 ; n32157
g29722 and pi0625_not n32157 ; n32158
g29723 and pi0625 n32049 ; n32159
g29724 nor pi1153 n32159 ; n32160
g29725 and n32158_not n32160 ; n32161
g29726 nor pi0608 n31987 ; n32162
g29727 and n32161_not n32162 ; n32163
g29728 and pi0625_not n32049 ; n32164
g29729 and pi0625 n32157 ; n32165
g29730 and pi1153 n32164_not ; n32166
g29731 and n32165_not n32166 ; n32167
g29732 and pi0608 n31991_not ; n32168
g29733 and n32167_not n32168 ; n32169
g29734 nor n32163 n32169 ; n32170
g29735 and pi0778 n32170_not ; n32171
g29736 and pi0778_not n32157 ; n32172
g29737 nor n32171 n32172 ; n32173
g29738 nor pi0609 n32173 ; n32174
g29739 nor pi1155 n32120 ; n32175
g29740 and n32174_not n32175 ; n32176
g29741 nor pi0660 n32057 ; n32177
g29742 and n32176_not n32177 ; n32178
g29743 and pi0609_not n31994 ; n32179
g29744 and pi0609 n32173_not ; n32180
g29745 and pi1155 n32179_not ; n32181
g29746 and n32180_not n32181 ; n32182
g29747 and pi0660 n32061_not ; n32183
g29748 and n32182_not n32183 ; n32184
g29749 nor n32178 n32184 ; n32185
g29750 and pi0785 n32185_not ; n32186
g29751 nor pi0785 n32173 ; n32187
g29752 nor n32186 n32187 ; n32188
g29753 nor pi0618 n32188 ; n32189
g29754 and pi0618 n31997 ; n32190
g29755 nor pi1154 n32190 ; n32191
g29756 and n32189_not n32191 ; n32192
g29757 nor pi0627 n32069 ; n32193
g29758 and n32192_not n32193 ; n32194
g29759 and pi0618_not n31997 ; n32195
g29760 and pi0618 n32188_not ; n32196
g29761 and pi1154 n32195_not ; n32197
g29762 and n32196_not n32197 ; n32198
g29763 and pi0627 n32073_not ; n32199
g29764 and n32198_not n32199 ; n32200
g29765 nor n32194 n32200 ; n32201
g29766 and pi0781 n32201_not ; n32202
g29767 nor pi0781 n32188 ; n32203
g29768 nor n32202 n32203 ; n32204
g29769 and pi0789_not n32204 ; n32205
g29770 and pi0619 n32000_not ; n32206
g29771 nor pi0619 n32204 ; n32207
g29772 nor pi1159 n32206 ; n32208
g29773 and n32207_not n32208 ; n32209
g29774 nor pi0648 n32081 ; n32210
g29775 and n32209_not n32210 ; n32211
g29776 nor pi0619 n32000 ; n32212
g29777 and pi0619 n32204_not ; n32213
g29778 and pi1159 n32212_not ; n32214
g29779 and n32213_not n32214 ; n32215
g29780 and pi0648 n32085_not ; n32216
g29781 and n32215_not n32216 ; n32217
g29782 and pi0789 n32211_not ; n32218
g29783 and n32217_not n32218 ; n32219
g29784 and n17970 n32205_not ; n32220
g29785 and n32219_not n32220 ; n32221
g29786 and n17871 n32002 ; n32222
g29787 nor pi0626 n32088 ; n32223
g29788 and pi0626 n31967_not ; n32224
g29789 and n16629 n32224_not ; n32225
g29790 and n32223_not n32225 ; n32226
g29791 and pi0626 n32088_not ; n32227
g29792 nor pi0626 n31967 ; n32228
g29793 and n16628 n32228_not ; n32229
g29794 and n32227_not n32229 ; n32230
g29795 nor n32222 n32226 ; n32231
g29796 and n32230_not n32231 ; n32232
g29797 and pi0788 n32232_not ; n32233
g29798 nor n20364 n32233 ; n32234
g29799 and n32221_not n32234 ; n32235
g29800 nor n32119 n32235 ; n32236
g29801 nor n20206 n32236 ; n32237
g29802 and n17802 n32020 ; n32238
g29803 and n20559_not n32094 ; n32239
g29804 and n17801 n32024 ; n32240
g29805 nor n32238 n32239 ; n32241
g29806 and n32240_not n32241 ; n32242
g29807 and pi0787 n32242_not ; n32243
g29808 and pi0644_not n32110 ; n32244
g29809 and pi0644 n32102 ; n32245
g29810 and pi0790 n32244_not ; n32246
g29811 and n32245_not n32246 ; n32247
g29812 nor n32237 n32243 ; n32248
g29813 and n32247_not n32248 ; n32249
g29814 nor n32113 n32249 ; n32250
g29815 nor po1038 n32250 ; n32251
g29816 nor pi0832 n31966 ; n32252
g29817 and n32251_not n32252 ; n32253
g29818 nor n31965 n32253 ; po0349
g29819 nor pi0193 n2926 ; n32255
g29820 and pi0690 n16645 ; n32256
g29821 nor n32255 n32256 ; n32257
g29822 nor pi0778 n32257 ; n32258
g29823 and pi0625_not n32256 ; n32259
g29824 nor n32257 n32259 ; n32260
g29825 and pi1153 n32260_not ; n32261
g29826 nor pi1153 n32255 ; n32262
g29827 and n32259_not n32262 ; n32263
g29828 and pi0778 n32263_not ; n32264
g29829 and n32261_not n32264 ; n32265
g29830 nor n32258 n32265 ; n32266
g29831 nor n17845 n32266 ; n32267
g29832 and n17847_not n32267 ; n32268
g29833 and n17849_not n32268 ; n32269
g29834 and n17851_not n32269 ; n32270
g29835 and n17857_not n32270 ; n32271
g29836 and pi0647_not n32271 ; n32272
g29837 and pi0647 n32255 ; n32273
g29838 nor pi1157 n32273 ; n32274
g29839 and n32272_not n32274 ; n32275
g29840 and pi0630 n32275 ; n32276
g29841 and pi0739 n17244 ; n32277
g29842 nor n32255 n32277 ; n32278
g29843 nor n17874 n32278 ; n32279
g29844 nor pi0785 n32279 ; n32280
g29845 and n17296 n32277 ; n32281
g29846 and n32279 n32281_not ; n32282
g29847 and pi1155 n32282_not ; n32283
g29848 nor pi1155 n32255 ; n32284
g29849 and n32281_not n32284 ; n32285
g29850 nor n32283 n32285 ; n32286
g29851 and pi0785 n32286_not ; n32287
g29852 nor n32280 n32287 ; n32288
g29853 nor pi0781 n32288 ; n32289
g29854 and n17889_not n32288 ; n32290
g29855 and pi1154 n32290_not ; n32291
g29856 and n17892_not n32288 ; n32292
g29857 nor pi1154 n32292 ; n32293
g29858 nor n32291 n32293 ; n32294
g29859 and pi0781 n32294_not ; n32295
g29860 nor n32289 n32295 ; n32296
g29861 nor pi0789 n32296 ; n32297
g29862 and n23078_not n32296 ; n32298
g29863 and pi1159 n32298_not ; n32299
g29864 and n23081_not n32296 ; n32300
g29865 nor pi1159 n32300 ; n32301
g29866 nor n32299 n32301 ; n32302
g29867 and pi0789 n32302_not ; n32303
g29868 nor n32297 n32303 ; n32304
g29869 and n17969_not n32304 ; n32305
g29870 and n17969 n32255 ; n32306
g29871 nor n32305 n32306 ; n32307
g29872 nor n17779 n32307 ; n32308
g29873 and n17779 n32255 ; n32309
g29874 nor n32308 n32309 ; n32310
g29875 and n20559_not n32310 ; n32311
g29876 and pi0647 n32271_not ; n32312
g29877 nor pi0647 n32255 ; n32313
g29878 nor n32312 n32313 ; n32314
g29879 and n17801 n32314_not ; n32315
g29880 nor n32276 n32315 ; n32316
g29881 and n32311_not n32316 ; n32317
g29882 and pi0787 n32317_not ; n32318
g29883 and n17871 n32269 ; n32319
g29884 nor pi0626 n32304 ; n32320
g29885 and pi0626 n32255_not ; n32321
g29886 and n16629 n32321_not ; n32322
g29887 and n32320_not n32322 ; n32323
g29888 and pi0626 n32304_not ; n32324
g29889 nor pi0626 n32255 ; n32325
g29890 and n16628 n32325_not ; n32326
g29891 and n32324_not n32326 ; n32327
g29892 nor n32319 n32323 ; n32328
g29893 and n32327_not n32328 ; n32329
g29894 and pi0788 n32329_not ; n32330
g29895 and pi0618 n32267 ; n32331
g29896 nor n17168 n32257 ; n32332
g29897 and pi0625 n32332 ; n32333
g29898 and n32278 n32332_not ; n32334
g29899 nor n32333 n32334 ; n32335
g29900 and n32262 n32335_not ; n32336
g29901 nor pi0608 n32261 ; n32337
g29902 and n32336_not n32337 ; n32338
g29903 and pi1153 n32278 ; n32339
g29904 and n32333_not n32339 ; n32340
g29905 and pi0608 n32263_not ; n32341
g29906 and n32340_not n32341 ; n32342
g29907 nor n32338 n32342 ; n32343
g29908 and pi0778 n32343_not ; n32344
g29909 nor pi0778 n32334 ; n32345
g29910 nor n32344 n32345 ; n32346
g29911 nor pi0609 n32346 ; n32347
g29912 and pi0609 n32266_not ; n32348
g29913 nor pi1155 n32348 ; n32349
g29914 and n32347_not n32349 ; n32350
g29915 nor pi0660 n32283 ; n32351
g29916 and n32350_not n32351 ; n32352
g29917 and pi0609 n32346_not ; n32353
g29918 nor pi0609 n32266 ; n32354
g29919 and pi1155 n32354_not ; n32355
g29920 and n32353_not n32355 ; n32356
g29921 and pi0660 n32285_not ; n32357
g29922 and n32356_not n32357 ; n32358
g29923 nor n32352 n32358 ; n32359
g29924 and pi0785 n32359_not ; n32360
g29925 nor pi0785 n32346 ; n32361
g29926 nor n32360 n32361 ; n32362
g29927 nor pi0618 n32362 ; n32363
g29928 nor pi1154 n32331 ; n32364
g29929 and n32363_not n32364 ; n32365
g29930 nor pi0627 n32291 ; n32366
g29931 and n32365_not n32366 ; n32367
g29932 and pi0618_not n32267 ; n32368
g29933 and pi0618 n32362_not ; n32369
g29934 and pi1154 n32368_not ; n32370
g29935 and n32369_not n32370 ; n32371
g29936 and pi0627 n32293_not ; n32372
g29937 and n32371_not n32372 ; n32373
g29938 nor n32367 n32373 ; n32374
g29939 and pi0781 n32374_not ; n32375
g29940 nor pi0781 n32362 ; n32376
g29941 nor n32375 n32376 ; n32377
g29942 and pi0789_not n32377 ; n32378
g29943 nor pi0619 n32377 ; n32379
g29944 and pi0619 n32268 ; n32380
g29945 nor pi1159 n32380 ; n32381
g29946 and n32379_not n32381 ; n32382
g29947 nor pi0648 n32299 ; n32383
g29948 and n32382_not n32383 ; n32384
g29949 and pi0619 n32377_not ; n32385
g29950 and pi0619_not n32268 ; n32386
g29951 and pi1159 n32386_not ; n32387
g29952 and n32385_not n32387 ; n32388
g29953 and pi0648 n32301_not ; n32389
g29954 and n32388_not n32389 ; n32390
g29955 and pi0789 n32384_not ; n32391
g29956 and n32390_not n32391 ; n32392
g29957 and n17970 n32378_not ; n32393
g29958 and n32392_not n32393 ; n32394
g29959 nor n32330 n32394 ; n32395
g29960 nor n20364 n32395 ; n32396
g29961 and n17854 n32307_not ; n32397
g29962 and n20851 n32270 ; n32398
g29963 nor n32397 n32398 ; n32399
g29964 nor pi0629 n32399 ; n32400
g29965 and n20855 n32270 ; n32401
g29966 and n17853 n32307_not ; n32402
g29967 nor n32401 n32402 ; n32403
g29968 and pi0629 n32403_not ; n32404
g29969 nor n32400 n32404 ; n32405
g29970 and pi0792 n32405_not ; n32406
g29971 nor n20206 n32406 ; n32407
g29972 and n32396_not n32407 ; n32408
g29973 nor n32318 n32408 ; n32409
g29974 and pi0790_not n32409 ; n32410
g29975 nor pi0787 n32271 ; n32411
g29976 and pi1157 n32314_not ; n32412
g29977 nor n32275 n32412 ; n32413
g29978 and pi0787 n32413_not ; n32414
g29979 nor n32411 n32414 ; n32415
g29980 and pi0644_not n32415 ; n32416
g29981 and pi0644 n32409 ; n32417
g29982 and pi0715 n32416_not ; n32418
g29983 and n32417_not n32418 ; n32419
g29984 nor n17804 n32310 ; n32420
g29985 and n17804 n32255 ; n32421
g29986 nor n32420 n32421 ; n32422
g29987 and pi0644 n32422_not ; n32423
g29988 and pi0644_not n32255 ; n32424
g29989 nor pi0715 n32424 ; n32425
g29990 and n32423_not n32425 ; n32426
g29991 and pi1160 n32426_not ; n32427
g29992 and n32419_not n32427 ; n32428
g29993 nor pi0644 n32422 ; n32429
g29994 and pi0644 n32255 ; n32430
g29995 and pi0715 n32430_not ; n32431
g29996 and n32429_not n32431 ; n32432
g29997 and pi0644 n32415 ; n32433
g29998 and pi0644_not n32409 ; n32434
g29999 nor pi0715 n32433 ; n32435
g30000 and n32434_not n32435 ; n32436
g30001 nor pi1160 n32432 ; n32437
g30002 and n32436_not n32437 ; n32438
g30003 nor n32428 n32438 ; n32439
g30004 and pi0790 n32439_not ; n32440
g30005 and pi0832 n32410_not ; n32441
g30006 and n32440_not n32441 ; n32442
g30007 and pi0193_not po1038 ; n32443
g30008 nor pi0193 n17059 ; n32444
g30009 and n16635 n32444_not ; n32445
g30010 and pi0690 n2571 ; n32446
g30011 and n32444 n32446_not ; n32447
g30012 nor pi0193 n16641 ; n32448
g30013 and n16647 n32448_not ; n32449
g30014 and pi0193 n18076_not ; n32450
g30015 nor pi0038 n32450 ; n32451
g30016 and n2571 n32451_not ; n32452
g30017 and pi0193_not n18072 ; n32453
g30018 nor n32452 n32453 ; n32454
g30019 and pi0690 n32449_not ; n32455
g30020 and n32454_not n32455 ; n32456
g30021 nor n32447 n32456 ; n32457
g30022 and pi0778_not n32457 ; n32458
g30023 and pi0625_not n32444 ; n32459
g30024 and pi0625 n32457_not ; n32460
g30025 and pi1153 n32459_not ; n32461
g30026 and n32460_not n32461 ; n32462
g30027 and pi0625 n32444 ; n32463
g30028 nor pi0625 n32457 ; n32464
g30029 nor pi1153 n32463 ; n32465
g30030 and n32464_not n32465 ; n32466
g30031 nor n32462 n32466 ; n32467
g30032 and pi0778 n32467_not ; n32468
g30033 nor n32458 n32468 ; n32469
g30034 nor n17075 n32469 ; n32470
g30035 and n17075 n32444_not ; n32471
g30036 nor n32470 n32471 ; n32472
g30037 and n16639_not n32472 ; n32473
g30038 and n16639 n32444 ; n32474
g30039 nor n32473 n32474 ; n32475
g30040 and n16635_not n32475 ; n32476
g30041 nor n32445 n32476 ; n32477
g30042 and n16631_not n32477 ; n32478
g30043 and n16631 n32444 ; n32479
g30044 nor n32478 n32479 ; n32480
g30045 and pi0792_not n32480 ; n32481
g30046 and pi0628 n32480_not ; n32482
g30047 and pi0628_not n32444 ; n32483
g30048 and pi1156 n32483_not ; n32484
g30049 and n32482_not n32484 ; n32485
g30050 and pi0628 n32444 ; n32486
g30051 nor pi0628 n32480 ; n32487
g30052 nor pi1156 n32486 ; n32488
g30053 and n32487_not n32488 ; n32489
g30054 nor n32485 n32489 ; n32490
g30055 and pi0792 n32490_not ; n32491
g30056 nor n32481 n32491 ; n32492
g30057 nor pi0647 n32492 ; n32493
g30058 and pi0647 n32444_not ; n32494
g30059 nor n32493 n32494 ; n32495
g30060 and pi1157_not n32495 ; n32496
g30061 and pi0647 n32492_not ; n32497
g30062 nor pi0647 n32444 ; n32498
g30063 nor n32497 n32498 ; n32499
g30064 and pi1157 n32499 ; n32500
g30065 nor n32496 n32500 ; n32501
g30066 and pi0787 n32501_not ; n32502
g30067 and pi0787_not n32492 ; n32503
g30068 nor n32502 n32503 ; n32504
g30069 nor pi0644 n32504 ; n32505
g30070 and pi0715 n32505_not ; n32506
g30071 and pi0193 n2571_not ; n32507
g30072 and pi0739 n17280 ; n32508
g30073 nor n32448 n32508 ; n32509
g30074 and pi0038 n32509_not ; n32510
g30075 and pi0193_not n17221 ; n32511
g30076 and pi0193 n17275_not ; n32512
g30077 and pi0739 n32512_not ; n32513
g30078 and n32511_not n32513 ; n32514
g30079 nor pi0193 pi0739 ; n32515
g30080 and n17048_not n32515 ; n32516
g30081 nor n32514 n32516 ; n32517
g30082 nor pi0038 n32517 ; n32518
g30083 nor n32510 n32518 ; n32519
g30084 and n2571 n32519 ; n32520
g30085 nor n32507 n32520 ; n32521
g30086 nor n17117 n32521 ; n32522
g30087 and n17117 n32444_not ; n32523
g30088 nor n32522 n32523 ; n32524
g30089 nor pi0785 n32524 ; n32525
g30090 nor n17291 n32444 ; n32526
g30091 and pi0609 n32522 ; n32527
g30092 nor n32526 n32527 ; n32528
g30093 and pi1155 n32528_not ; n32529
g30094 nor n17296 n32444 ; n32530
g30095 and pi0609_not n32522 ; n32531
g30096 nor n32530 n32531 ; n32532
g30097 nor pi1155 n32532 ; n32533
g30098 nor n32529 n32533 ; n32534
g30099 and pi0785 n32534_not ; n32535
g30100 nor n32525 n32535 ; n32536
g30101 nor pi0781 n32536 ; n32537
g30102 and pi0618_not n32444 ; n32538
g30103 and pi0618 n32536 ; n32539
g30104 and pi1154 n32538_not ; n32540
g30105 and n32539_not n32540 ; n32541
g30106 and pi0618_not n32536 ; n32542
g30107 and pi0618 n32444 ; n32543
g30108 nor pi1154 n32543 ; n32544
g30109 and n32542_not n32544 ; n32545
g30110 nor n32541 n32545 ; n32546
g30111 and pi0781 n32546_not ; n32547
g30112 nor n32537 n32547 ; n32548
g30113 nor pi0789 n32548 ; n32549
g30114 and pi0619_not n32444 ; n32550
g30115 and pi0619 n32548 ; n32551
g30116 and pi1159 n32550_not ; n32552
g30117 and n32551_not n32552 ; n32553
g30118 and pi0619_not n32548 ; n32554
g30119 and pi0619 n32444 ; n32555
g30120 nor pi1159 n32555 ; n32556
g30121 and n32554_not n32556 ; n32557
g30122 nor n32553 n32557 ; n32558
g30123 and pi0789 n32558_not ; n32559
g30124 nor n32549 n32559 ; n32560
g30125 and n17969_not n32560 ; n32561
g30126 and n17969 n32444 ; n32562
g30127 nor n32561 n32562 ; n32563
g30128 nor n17779 n32563 ; n32564
g30129 and n17779 n32444 ; n32565
g30130 nor n32564 n32565 ; n32566
g30131 nor n17804 n32566 ; n32567
g30132 and n17804 n32444 ; n32568
g30133 nor n32567 n32568 ; n32569
g30134 and pi0644 n32569_not ; n32570
g30135 and pi0644_not n32444 ; n32571
g30136 nor pi0715 n32571 ; n32572
g30137 and n32570_not n32572 ; n32573
g30138 and pi1160 n32573_not ; n32574
g30139 and n32506_not n32574 ; n32575
g30140 and pi0644 n32504_not ; n32576
g30141 nor pi0715 n32576 ; n32577
g30142 nor pi0644 n32569 ; n32578
g30143 and pi0644 n32444 ; n32579
g30144 and pi0715 n32579_not ; n32580
g30145 and n32578_not n32580 ; n32581
g30146 nor pi1160 n32581 ; n32582
g30147 and n32577_not n32582 ; n32583
g30148 nor n32575 n32583 ; n32584
g30149 and pi0790 n32584_not ; n32585
g30150 and pi0629_not n32485 ; n32586
g30151 and n20570_not n32563 ; n32587
g30152 and pi0629 n32489 ; n32588
g30153 nor n32586 n32588 ; n32589
g30154 and n32587_not n32589 ; n32590
g30155 and pi0792 n32590_not ; n32591
g30156 and pi0609 n32469 ; n32592
g30157 nor pi0690 n32519 ; n32593
g30158 and pi0193_not n17629 ; n32594
g30159 and pi0193 n17631 ; n32595
g30160 and pi0739 n32595_not ; n32596
g30161 and n32594_not n32596 ; n32597
g30162 and pi0193 n17625_not ; n32598
g30163 nor pi0193 n17612 ; n32599
g30164 nor pi0739 n32598 ; n32600
g30165 and n32599_not n32600 ; n32601
g30166 nor n32597 n32601 ; n32602
g30167 nor pi0039 n32602 ; n32603
g30168 and pi0193 n17605 ; n32604
g30169 nor pi0193 n17546 ; n32605
g30170 and pi0739 n32605_not ; n32606
g30171 and n32604_not n32606 ; n32607
g30172 and pi0193_not n17404 ; n32608
g30173 and pi0193 n17485 ; n32609
g30174 nor pi0739 n32609 ; n32610
g30175 and n32608_not n32610 ; n32611
g30176 and pi0039 n32607_not ; n32612
g30177 and n32611_not n32612 ; n32613
g30178 nor pi0038 n32603 ; n32614
g30179 and n32613_not n32614 ; n32615
g30180 and pi0739_not n24055 ; n32616
g30181 nor n17490 n32616 ; n32617
g30182 nor pi0039 n32617 ; n32618
g30183 nor pi0193 n32618 ; n32619
g30184 nor n17469 n32277 ; n32620
g30185 and pi0193 n32620_not ; n32621
g30186 and n6284 n32621 ; n32622
g30187 and pi0038 n32622_not ; n32623
g30188 and n32619_not n32623 ; n32624
g30189 and pi0690 n32624_not ; n32625
g30190 and n32615_not n32625 ; n32626
g30191 and n2571 n32626_not ; n32627
g30192 and n32593_not n32627 ; n32628
g30193 nor n32507 n32628 ; n32629
g30194 and pi0625_not n32629 ; n32630
g30195 and pi0625 n32521 ; n32631
g30196 nor pi1153 n32631 ; n32632
g30197 and n32630_not n32632 ; n32633
g30198 nor pi0608 n32462 ; n32634
g30199 and n32633_not n32634 ; n32635
g30200 and pi0625_not n32521 ; n32636
g30201 and pi0625 n32629 ; n32637
g30202 and pi1153 n32636_not ; n32638
g30203 and n32637_not n32638 ; n32639
g30204 and pi0608 n32466_not ; n32640
g30205 and n32639_not n32640 ; n32641
g30206 nor n32635 n32641 ; n32642
g30207 and pi0778 n32642_not ; n32643
g30208 and pi0778_not n32629 ; n32644
g30209 nor n32643 n32644 ; n32645
g30210 nor pi0609 n32645 ; n32646
g30211 nor pi1155 n32592 ; n32647
g30212 and n32646_not n32647 ; n32648
g30213 nor pi0660 n32529 ; n32649
g30214 and n32648_not n32649 ; n32650
g30215 and pi0609_not n32469 ; n32651
g30216 and pi0609 n32645_not ; n32652
g30217 and pi1155 n32651_not ; n32653
g30218 and n32652_not n32653 ; n32654
g30219 and pi0660 n32533_not ; n32655
g30220 and n32654_not n32655 ; n32656
g30221 nor n32650 n32656 ; n32657
g30222 and pi0785 n32657_not ; n32658
g30223 nor pi0785 n32645 ; n32659
g30224 nor n32658 n32659 ; n32660
g30225 nor pi0618 n32660 ; n32661
g30226 and pi0618 n32472 ; n32662
g30227 nor pi1154 n32662 ; n32663
g30228 and n32661_not n32663 ; n32664
g30229 nor pi0627 n32541 ; n32665
g30230 and n32664_not n32665 ; n32666
g30231 and pi0618_not n32472 ; n32667
g30232 and pi0618 n32660_not ; n32668
g30233 and pi1154 n32667_not ; n32669
g30234 and n32668_not n32669 ; n32670
g30235 and pi0627 n32545_not ; n32671
g30236 and n32670_not n32671 ; n32672
g30237 nor n32666 n32672 ; n32673
g30238 and pi0781 n32673_not ; n32674
g30239 nor pi0781 n32660 ; n32675
g30240 nor n32674 n32675 ; n32676
g30241 and pi0789_not n32676 ; n32677
g30242 and pi0619 n32475_not ; n32678
g30243 nor pi0619 n32676 ; n32679
g30244 nor pi1159 n32678 ; n32680
g30245 and n32679_not n32680 ; n32681
g30246 nor pi0648 n32553 ; n32682
g30247 and n32681_not n32682 ; n32683
g30248 nor pi0619 n32475 ; n32684
g30249 and pi0619 n32676_not ; n32685
g30250 and pi1159 n32684_not ; n32686
g30251 and n32685_not n32686 ; n32687
g30252 and pi0648 n32557_not ; n32688
g30253 and n32687_not n32688 ; n32689
g30254 and pi0789 n32683_not ; n32690
g30255 and n32689_not n32690 ; n32691
g30256 and n17970 n32677_not ; n32692
g30257 and n32691_not n32692 ; n32693
g30258 and n17871 n32477 ; n32694
g30259 nor pi0626 n32560 ; n32695
g30260 and pi0626 n32444_not ; n32696
g30261 and n16629 n32696_not ; n32697
g30262 and n32695_not n32697 ; n32698
g30263 and pi0626 n32560_not ; n32699
g30264 nor pi0626 n32444 ; n32700
g30265 and n16628 n32700_not ; n32701
g30266 and n32699_not n32701 ; n32702
g30267 nor n32694 n32698 ; n32703
g30268 and n32702_not n32703 ; n32704
g30269 and pi0788 n32704_not ; n32705
g30270 nor n20364 n32705 ; n32706
g30271 and n32693_not n32706 ; n32707
g30272 nor n32591 n32707 ; n32708
g30273 nor n20206 n32708 ; n32709
g30274 and n17802 n32495_not ; n32710
g30275 and n20559_not n32566 ; n32711
g30276 and n17801 n32499_not ; n32712
g30277 nor n32710 n32712 ; n32713
g30278 and n32711_not n32713 ; n32714
g30279 and pi0787 n32714_not ; n32715
g30280 and pi0644_not n32582 ; n32716
g30281 and pi0644 n32574 ; n32717
g30282 and pi0790 n32716_not ; n32718
g30283 and n32717_not n32718 ; n32719
g30284 nor n32709 n32715 ; n32720
g30285 and n32719_not n32720 ; n32721
g30286 nor n32585 n32721 ; n32722
g30287 nor po1038 n32722 ; n32723
g30288 nor pi0832 n32443 ; n32724
g30289 and n32723_not n32724 ; n32725
g30290 nor n32442 n32725 ; po0350
g30291 nor pi0194 n17059 ; n32727
g30292 and n16635 n32727_not ; n32728
g30293 and pi0194 n24385_not ; n32729
g30294 and pi0194_not n24388 ; n32730
g30295 and pi0730 n32730_not ; n32731
g30296 nor pi0194 n17052 ; n32732
g30297 and pi0730_not n32732 ; n32733
g30298 and n2571 n32733_not ; n32734
g30299 and n32731_not n32734 ; n32735
g30300 nor n32729 n32735 ; n32736
g30301 nor pi0778 n32736 ; n32737
g30302 and pi0625_not n32727 ; n32738
g30303 and pi0625 n32736 ; n32739
g30304 and pi1153 n32738_not ; n32740
g30305 and n32739_not n32740 ; n32741
g30306 and pi0625_not n32736 ; n32742
g30307 and pi0625 n32727 ; n32743
g30308 nor pi1153 n32743 ; n32744
g30309 and n32742_not n32744 ; n32745
g30310 nor n32741 n32745 ; n32746
g30311 and pi0778 n32746_not ; n32747
g30312 nor n32737 n32747 ; n32748
g30313 nor n17075 n32748 ; n32749
g30314 and n17075 n32727_not ; n32750
g30315 nor n32749 n32750 ; n32751
g30316 and n16639_not n32751 ; n32752
g30317 and n16639 n32727 ; n32753
g30318 nor n32752 n32753 ; n32754
g30319 and n16635_not n32754 ; n32755
g30320 nor n32728 n32755 ; n32756
g30321 and n16631_not n32756 ; n32757
g30322 and n16631 n32727 ; n32758
g30323 nor n32757 n32758 ; n32759
g30324 and pi0792_not n32759 ; n32760
g30325 and pi0628_not n32727 ; n32761
g30326 and pi0628 n32759_not ; n32762
g30327 and pi1156 n32761_not ; n32763
g30328 and n32762_not n32763 ; n32764
g30329 and pi0628 n32727 ; n32765
g30330 nor pi0628 n32759 ; n32766
g30331 nor pi1156 n32765 ; n32767
g30332 and n32766_not n32767 ; n32768
g30333 nor n32764 n32768 ; n32769
g30334 and pi0792 n32769_not ; n32770
g30335 nor n32760 n32770 ; n32771
g30336 nor pi0787 n32771 ; n32772
g30337 and pi0647_not n32727 ; n32773
g30338 and pi0647 n32771 ; n32774
g30339 and pi1157 n32773_not ; n32775
g30340 and n32774_not n32775 ; n32776
g30341 and pi0647_not n32771 ; n32777
g30342 and pi0647 n32727 ; n32778
g30343 nor pi1157 n32778 ; n32779
g30344 and n32777_not n32779 ; n32780
g30345 nor n32776 n32780 ; n32781
g30346 and pi0787 n32781_not ; n32782
g30347 nor n32772 n32782 ; n32783
g30348 and pi0644_not n32783 ; n32784
g30349 and pi0618_not n32727 ; n32785
g30350 and pi0194 n2571_not ; n32786
g30351 and pi0194_not n19439 ; n32787
g30352 and pi0194 n24447 ; n32788
g30353 nor n32787 n32788 ; n32789
g30354 and pi0748 n32789_not ; n32790
g30355 nor pi0748 n32732 ; n32791
g30356 nor n32790 n32791 ; n32792
g30357 and n2571 n32792_not ; n32793
g30358 nor n32786 n32793 ; n32794
g30359 nor n17117 n32794 ; n32795
g30360 and n17117 n32727_not ; n32796
g30361 nor n32795 n32796 ; n32797
g30362 nor pi0785 n32797 ; n32798
g30363 nor n17291 n32727 ; n32799
g30364 and pi0609 n32795 ; n32800
g30365 nor n32799 n32800 ; n32801
g30366 and pi1155 n32801_not ; n32802
g30367 nor n17296 n32727 ; n32803
g30368 and pi0609_not n32795 ; n32804
g30369 nor n32803 n32804 ; n32805
g30370 nor pi1155 n32805 ; n32806
g30371 nor n32802 n32806 ; n32807
g30372 and pi0785 n32807_not ; n32808
g30373 nor n32798 n32808 ; n32809
g30374 and pi0618 n32809 ; n32810
g30375 and pi1154 n32785_not ; n32811
g30376 and n32810_not n32811 ; n32812
g30377 and pi0730_not n32792 ; n32813
g30378 and pi0194 n19496 ; n32814
g30379 nor pi0194 n19488 ; n32815
g30380 and pi0748 n32815_not ; n32816
g30381 and n32814_not n32816 ; n32817
g30382 and pi0194 n24549_not ; n32818
g30383 and pi0194_not n19477 ; n32819
g30384 nor pi0748 n32818 ; n32820
g30385 and n32819_not n32820 ; n32821
g30386 and pi0730 n32817_not ; n32822
g30387 and n32821_not n32822 ; n32823
g30388 and n2571 n32813_not ; n32824
g30389 and n32823_not n32824 ; n32825
g30390 nor n32786 n32825 ; n32826
g30391 and pi0625_not n32826 ; n32827
g30392 and pi0625 n32794 ; n32828
g30393 nor pi1153 n32828 ; n32829
g30394 and n32827_not n32829 ; n32830
g30395 nor pi0608 n32741 ; n32831
g30396 and n32830_not n32831 ; n32832
g30397 and pi0625_not n32794 ; n32833
g30398 and pi0625 n32826 ; n32834
g30399 and pi1153 n32833_not ; n32835
g30400 and n32834_not n32835 ; n32836
g30401 and pi0608 n32745_not ; n32837
g30402 and n32836_not n32837 ; n32838
g30403 nor n32832 n32838 ; n32839
g30404 and pi0778 n32839_not ; n32840
g30405 and pi0778_not n32826 ; n32841
g30406 nor n32840 n32841 ; n32842
g30407 nor pi0609 n32842 ; n32843
g30408 and pi0609 n32748 ; n32844
g30409 nor pi1155 n32844 ; n32845
g30410 and n32843_not n32845 ; n32846
g30411 nor pi0660 n32802 ; n32847
g30412 and n32846_not n32847 ; n32848
g30413 and pi0609_not n32748 ; n32849
g30414 and pi0609 n32842_not ; n32850
g30415 and pi1155 n32849_not ; n32851
g30416 and n32850_not n32851 ; n32852
g30417 and pi0660 n32806_not ; n32853
g30418 and n32852_not n32853 ; n32854
g30419 nor n32848 n32854 ; n32855
g30420 and pi0785 n32855_not ; n32856
g30421 nor pi0785 n32842 ; n32857
g30422 nor n32856 n32857 ; n32858
g30423 nor pi0618 n32858 ; n32859
g30424 and pi0618 n32751 ; n32860
g30425 nor pi1154 n32860 ; n32861
g30426 and n32859_not n32861 ; n32862
g30427 nor pi0627 n32812 ; n32863
g30428 and n32862_not n32863 ; n32864
g30429 and pi0618_not n32809 ; n32865
g30430 and pi0618 n32727 ; n32866
g30431 nor pi1154 n32866 ; n32867
g30432 and n32865_not n32867 ; n32868
g30433 and pi0618_not n32751 ; n32869
g30434 and pi0618 n32858_not ; n32870
g30435 and pi1154 n32869_not ; n32871
g30436 and n32870_not n32871 ; n32872
g30437 and pi0627 n32868_not ; n32873
g30438 and n32872_not n32873 ; n32874
g30439 nor n32864 n32874 ; n32875
g30440 and pi0781 n32875_not ; n32876
g30441 nor pi0781 n32858 ; n32877
g30442 nor n32876 n32877 ; n32878
g30443 nor pi0619 n32878 ; n32879
g30444 and pi0619 n32754_not ; n32880
g30445 nor pi1159 n32880 ; n32881
g30446 and n32879_not n32881 ; n32882
g30447 and pi0619_not n32727 ; n32883
g30448 nor pi0781 n32809 ; n32884
g30449 nor n32812 n32868 ; n32885
g30450 and pi0781 n32885_not ; n32886
g30451 nor n32884 n32886 ; n32887
g30452 and pi0619 n32887 ; n32888
g30453 and pi1159 n32883_not ; n32889
g30454 and n32888_not n32889 ; n32890
g30455 nor pi0648 n32890 ; n32891
g30456 and n32882_not n32891 ; n32892
g30457 and pi0619 n32878_not ; n32893
g30458 nor pi0619 n32754 ; n32894
g30459 and pi1159 n32894_not ; n32895
g30460 and n32893_not n32895 ; n32896
g30461 and pi0619_not n32887 ; n32897
g30462 and pi0619 n32727 ; n32898
g30463 nor pi1159 n32898 ; n32899
g30464 and n32897_not n32899 ; n32900
g30465 and pi0648 n32900_not ; n32901
g30466 and n32896_not n32901 ; n32902
g30467 nor n32892 n32902 ; n32903
g30468 and pi0789 n32903_not ; n32904
g30469 nor pi0789 n32878 ; n32905
g30470 nor n32904 n32905 ; n32906
g30471 and pi0788_not n32906 ; n32907
g30472 and pi0626_not n32906 ; n32908
g30473 and pi0626 n32756_not ; n32909
g30474 nor pi0641 n32909 ; n32910
g30475 and n32908_not n32910 ; n32911
g30476 nor pi0789 n32887 ; n32912
g30477 nor n32890 n32900 ; n32913
g30478 and pi0789 n32913_not ; n32914
g30479 nor n32912 n32914 ; n32915
g30480 nor pi0626 n32915 ; n32916
g30481 and pi0626 n32727_not ; n32917
g30482 and pi0641 n32917_not ; n32918
g30483 and n32916_not n32918 ; n32919
g30484 nor pi1158 n32919 ; n32920
g30485 and n32911_not n32920 ; n32921
g30486 and pi0626 n32906 ; n32922
g30487 nor pi0626 n32756 ; n32923
g30488 and pi0641 n32923_not ; n32924
g30489 and n32922_not n32924 ; n32925
g30490 and pi0626 n32915_not ; n32926
g30491 nor pi0626 n32727 ; n32927
g30492 nor pi0641 n32927 ; n32928
g30493 and n32926_not n32928 ; n32929
g30494 and pi1158 n32929_not ; n32930
g30495 and n32925_not n32930 ; n32931
g30496 nor n32921 n32931 ; n32932
g30497 and pi0788 n32932_not ; n32933
g30498 nor n32907 n32933 ; n32934
g30499 and pi0628_not n32934 ; n32935
g30500 and n17969_not n32915 ; n32936
g30501 and n17969 n32727 ; n32937
g30502 nor n32936 n32937 ; n32938
g30503 and pi0628 n32938_not ; n32939
g30504 nor pi1156 n32939 ; n32940
g30505 and n32935_not n32940 ; n32941
g30506 nor pi0629 n32764 ; n32942
g30507 and n32941_not n32942 ; n32943
g30508 and pi0628 n32934 ; n32944
g30509 nor pi0628 n32938 ; n32945
g30510 and pi1156 n32945_not ; n32946
g30511 and n32944_not n32946 ; n32947
g30512 and pi0629 n32768_not ; n32948
g30513 and n32947_not n32948 ; n32949
g30514 nor n32943 n32949 ; n32950
g30515 and pi0792 n32950_not ; n32951
g30516 and pi0792_not n32934 ; n32952
g30517 nor n32951 n32952 ; n32953
g30518 nor pi0647 n32953 ; n32954
g30519 nor n17779 n32938 ; n32955
g30520 and n17779 n32727 ; n32956
g30521 nor n32955 n32956 ; n32957
g30522 and pi0647 n32957_not ; n32958
g30523 nor pi1157 n32958 ; n32959
g30524 and n32954_not n32959 ; n32960
g30525 nor pi0630 n32776 ; n32961
g30526 and n32960_not n32961 ; n32962
g30527 and pi0647 n32953_not ; n32963
g30528 nor pi0647 n32957 ; n32964
g30529 and pi1157 n32964_not ; n32965
g30530 and n32963_not n32965 ; n32966
g30531 and pi0630 n32780_not ; n32967
g30532 and n32966_not n32967 ; n32968
g30533 nor n32962 n32968 ; n32969
g30534 and pi0787 n32969_not ; n32970
g30535 nor pi0787 n32953 ; n32971
g30536 nor n32970 n32971 ; n32972
g30537 and pi0644 n32972_not ; n32973
g30538 and pi0715 n32784_not ; n32974
g30539 and n32973_not n32974 ; n32975
g30540 and n17804 n32727_not ; n32976
g30541 and n17804_not n32957 ; n32977
g30542 nor n32976 n32977 ; n32978
g30543 and pi0644 n32978 ; n32979
g30544 and pi0644_not n32727 ; n32980
g30545 nor pi0715 n32980 ; n32981
g30546 and n32979_not n32981 ; n32982
g30547 and pi1160 n32982_not ; n32983
g30548 and n32975_not n32983 ; n32984
g30549 nor pi0644 n32972 ; n32985
g30550 and pi0644 n32783 ; n32986
g30551 nor pi0715 n32986 ; n32987
g30552 and n32985_not n32987 ; n32988
g30553 and pi0644_not n32978 ; n32989
g30554 and pi0644 n32727 ; n32990
g30555 and pi0715 n32990_not ; n32991
g30556 and n32989_not n32991 ; n32992
g30557 nor pi1160 n32992 ; n32993
g30558 and n32988_not n32993 ; n32994
g30559 and pi0790 n32984_not ; n32995
g30560 and n32994_not n32995 ; n32996
g30561 and pi0790_not n32972 ; n32997
g30562 nor po1038 n32997 ; n32998
g30563 and n32996_not n32998 ; n32999
g30564 and pi0194_not po1038 ; n33000
g30565 nor pi0832 n33000 ; n33001
g30566 and n32999_not n33001 ; n33002
g30567 nor pi0194 n2926 ; n33003
g30568 and pi0730 n16645 ; n33004
g30569 nor n33003 n33004 ; n33005
g30570 and pi0778_not n33005 ; n33006
g30571 and pi0625_not n33004 ; n33007
g30572 nor n33005 n33007 ; n33008
g30573 and pi1153 n33008_not ; n33009
g30574 nor pi1153 n33003 ; n33010
g30575 and n33007_not n33010 ; n33011
g30576 nor n33009 n33011 ; n33012
g30577 and pi0778 n33012_not ; n33013
g30578 nor n33006 n33013 ; n33014
g30579 and n17845_not n33014 ; n33015
g30580 and n17847_not n33015 ; n33016
g30581 and n17849_not n33016 ; n33017
g30582 and n17851_not n33017 ; n33018
g30583 and n17857_not n33018 ; n33019
g30584 and pi0647_not n33019 ; n33020
g30585 and pi0647 n33003 ; n33021
g30586 nor pi1157 n33021 ; n33022
g30587 and n33020_not n33022 ; n33023
g30588 and pi0630 n33023 ; n33024
g30589 and pi0748 n17244 ; n33025
g30590 nor n33003 n33025 ; n33026
g30591 nor n17874 n33026 ; n33027
g30592 nor pi0785 n33027 ; n33028
g30593 nor n17879 n33026 ; n33029
g30594 and pi1155 n33029_not ; n33030
g30595 and n17882_not n33027 ; n33031
g30596 nor pi1155 n33031 ; n33032
g30597 nor n33030 n33032 ; n33033
g30598 and pi0785 n33033_not ; n33034
g30599 nor n33028 n33034 ; n33035
g30600 nor pi0781 n33035 ; n33036
g30601 and n17889_not n33035 ; n33037
g30602 and pi1154 n33037_not ; n33038
g30603 and n17892_not n33035 ; n33039
g30604 nor pi1154 n33039 ; n33040
g30605 nor n33038 n33040 ; n33041
g30606 and pi0781 n33041_not ; n33042
g30607 nor n33036 n33042 ; n33043
g30608 nor pi0789 n33043 ; n33044
g30609 and pi0619_not n33003 ; n33045
g30610 and pi0619 n33043 ; n33046
g30611 and pi1159 n33045_not ; n33047
g30612 and n33046_not n33047 ; n33048
g30613 and pi0619_not n33043 ; n33049
g30614 and pi0619 n33003 ; n33050
g30615 nor pi1159 n33050 ; n33051
g30616 and n33049_not n33051 ; n33052
g30617 nor n33048 n33052 ; n33053
g30618 and pi0789 n33053_not ; n33054
g30619 nor n33044 n33054 ; n33055
g30620 and n17969_not n33055 ; n33056
g30621 and n17969 n33003 ; n33057
g30622 nor n33056 n33057 ; n33058
g30623 nor n17779 n33058 ; n33059
g30624 and n17779 n33003 ; n33060
g30625 nor n33059 n33060 ; n33061
g30626 and n20559_not n33061 ; n33062
g30627 and pi0647 n33019_not ; n33063
g30628 nor pi0647 n33003 ; n33064
g30629 nor n33063 n33064 ; n33065
g30630 and n17801 n33065_not ; n33066
g30631 nor n33024 n33066 ; n33067
g30632 and n33062_not n33067 ; n33068
g30633 and pi0787 n33068_not ; n33069
g30634 and n17871 n33017 ; n33070
g30635 nor pi0626 n33055 ; n33071
g30636 and pi0626 n33003_not ; n33072
g30637 and n16629 n33072_not ; n33073
g30638 and n33071_not n33073 ; n33074
g30639 and pi0626 n33055_not ; n33075
g30640 nor pi0626 n33003 ; n33076
g30641 and n16628 n33076_not ; n33077
g30642 and n33075_not n33077 ; n33078
g30643 nor n33070 n33074 ; n33079
g30644 and n33078_not n33079 ; n33080
g30645 and pi0788 n33080_not ; n33081
g30646 and pi0618 n33015 ; n33082
g30647 and pi0609 n33014 ; n33083
g30648 nor n17168 n33005 ; n33084
g30649 and pi0625 n33084 ; n33085
g30650 and n33026 n33084_not ; n33086
g30651 nor n33085 n33086 ; n33087
g30652 and n33010 n33087_not ; n33088
g30653 nor pi0608 n33009 ; n33089
g30654 and n33088_not n33089 ; n33090
g30655 and pi1153 n33026 ; n33091
g30656 and n33085_not n33091 ; n33092
g30657 and pi0608 n33011_not ; n33093
g30658 and n33092_not n33093 ; n33094
g30659 nor n33090 n33094 ; n33095
g30660 and pi0778 n33095_not ; n33096
g30661 nor pi0778 n33086 ; n33097
g30662 nor n33096 n33097 ; n33098
g30663 nor pi0609 n33098 ; n33099
g30664 nor pi1155 n33083 ; n33100
g30665 and n33099_not n33100 ; n33101
g30666 nor pi0660 n33030 ; n33102
g30667 and n33101_not n33102 ; n33103
g30668 and pi0609_not n33014 ; n33104
g30669 and pi0609 n33098_not ; n33105
g30670 and pi1155 n33104_not ; n33106
g30671 and n33105_not n33106 ; n33107
g30672 and pi0660 n33032_not ; n33108
g30673 and n33107_not n33108 ; n33109
g30674 nor n33103 n33109 ; n33110
g30675 and pi0785 n33110_not ; n33111
g30676 nor pi0785 n33098 ; n33112
g30677 nor n33111 n33112 ; n33113
g30678 nor pi0618 n33113 ; n33114
g30679 nor pi1154 n33082 ; n33115
g30680 and n33114_not n33115 ; n33116
g30681 nor pi0627 n33038 ; n33117
g30682 and n33116_not n33117 ; n33118
g30683 and pi0618_not n33015 ; n33119
g30684 and pi0618 n33113_not ; n33120
g30685 and pi1154 n33119_not ; n33121
g30686 and n33120_not n33121 ; n33122
g30687 and pi0627 n33040_not ; n33123
g30688 and n33122_not n33123 ; n33124
g30689 nor n33118 n33124 ; n33125
g30690 and pi0781 n33125_not ; n33126
g30691 nor pi0781 n33113 ; n33127
g30692 nor n33126 n33127 ; n33128
g30693 and pi0789_not n33128 ; n33129
g30694 nor pi0619 n33128 ; n33130
g30695 and pi0619 n33016 ; n33131
g30696 nor pi1159 n33131 ; n33132
g30697 and n33130_not n33132 ; n33133
g30698 nor pi0648 n33048 ; n33134
g30699 and n33133_not n33134 ; n33135
g30700 and pi0619 n33128_not ; n33136
g30701 and pi0619_not n33016 ; n33137
g30702 and pi1159 n33137_not ; n33138
g30703 and n33136_not n33138 ; n33139
g30704 and pi0648 n33052_not ; n33140
g30705 and n33139_not n33140 ; n33141
g30706 and pi0789 n33135_not ; n33142
g30707 and n33141_not n33142 ; n33143
g30708 and n17970 n33129_not ; n33144
g30709 and n33143_not n33144 ; n33145
g30710 nor n33081 n33145 ; n33146
g30711 nor n20364 n33146 ; n33147
g30712 and n17854 n33058_not ; n33148
g30713 and n20851 n33018 ; n33149
g30714 nor n33148 n33149 ; n33150
g30715 nor pi0629 n33150 ; n33151
g30716 and n20855 n33018 ; n33152
g30717 and n17853 n33058_not ; n33153
g30718 nor n33152 n33153 ; n33154
g30719 and pi0629 n33154_not ; n33155
g30720 nor n33151 n33155 ; n33156
g30721 and pi0792 n33156_not ; n33157
g30722 nor n20206 n33157 ; n33158
g30723 and n33147_not n33158 ; n33159
g30724 nor n33069 n33159 ; n33160
g30725 and pi0790_not n33160 ; n33161
g30726 nor pi0787 n33019 ; n33162
g30727 and pi1157 n33065_not ; n33163
g30728 nor n33023 n33163 ; n33164
g30729 and pi0787 n33164_not ; n33165
g30730 nor n33162 n33165 ; n33166
g30731 and pi0644_not n33166 ; n33167
g30732 and pi0644 n33160 ; n33168
g30733 and pi0715 n33167_not ; n33169
g30734 and n33168_not n33169 ; n33170
g30735 nor n17804 n33061 ; n33171
g30736 and n17804 n33003 ; n33172
g30737 nor n33171 n33172 ; n33173
g30738 and pi0644 n33173_not ; n33174
g30739 and pi0644_not n33003 ; n33175
g30740 nor pi0715 n33175 ; n33176
g30741 and n33174_not n33176 ; n33177
g30742 and pi1160 n33177_not ; n33178
g30743 and n33170_not n33178 ; n33179
g30744 nor pi0644 n33173 ; n33180
g30745 and pi0644 n33003 ; n33181
g30746 and pi0715 n33181_not ; n33182
g30747 and n33180_not n33182 ; n33183
g30748 and pi0644 n33166 ; n33184
g30749 and pi0644_not n33160 ; n33185
g30750 nor pi0715 n33184 ; n33186
g30751 and n33185_not n33186 ; n33187
g30752 nor pi1160 n33183 ; n33188
g30753 and n33187_not n33188 ; n33189
g30754 nor n33179 n33189 ; n33190
g30755 and pi0790 n33190_not ; n33191
g30756 and pi0832 n33161_not ; n33192
g30757 and n33191_not n33192 ; n33193
g30758 nor n33002 n33193 ; po0351
g30759 and pi0138_not n16565 ; n33195
g30760 and pi0196_not n33195 ; n33196
g30761 and pi0195 n33196_not ; n33197
g30762 and n11477_not n16193 ; n33198
g30763 and n6198_not n16168 ; n33199
g30764 and n16167 n16493_not ; n33200
g30765 nor n11480 n33199 ; n33201
g30766 nor n33198 n33200 ; n33202
g30767 and n33201 n33202 ; n33203
g30768 and pi0232 n33203_not ; n33204
g30769 nor n16491 n33204 ; n33205
g30770 and pi0039 n33205_not ; n33206
g30771 and n13910 n16170_not ; n33207
g30772 nor pi0039 n33207 ; n33208
g30773 and n10200 n33197_not ; n33209
g30774 and n33208_not n33209 ; n33210
g30775 and n33206_not n33210 ; n33211
g30776 and pi0171_not n9326 ; n33212
g30777 nor n16522 n33212 ; n33213
g30778 and n9036 n33213_not ; n33214
g30779 and n9291 n33214_not ; n33215
g30780 and pi0192_not n16511 ; n33216
g30781 and pi0192 n16520 ; n33217
g30782 nor n33215 n33216 ; n33218
g30783 and n33217_not n33218 ; n33219
g30784 and pi0232 n33219_not ; n33220
g30785 nor n16517 n33220 ; n33221
g30786 and pi0039 n33221_not ; n33222
g30787 and pi0192 n16539 ; n33223
g30788 nor n9605 n16162 ; n33224
g30789 and pi0171 n13737 ; n33225
g30790 nor n33224 n33225 ; n33226
g30791 and pi0299 n33226_not ; n33227
g30792 and pi0192_not n16533 ; n33228
g30793 and pi0232 n33228_not ; n33229
g30794 and n33223_not n33229 ; n33230
g30795 and n33227_not n33230 ; n33231
g30796 and n16536 n33231_not ; n33232
g30797 and n2608 n33222_not ; n33233
g30798 and n33232_not n33233 ; n33234
g30799 nor pi0087 n33234 ; n33235
g30800 and n16508 n33235_not ; n33236
g30801 nor pi0092 n33236 ; n33237
g30802 and n16507 n33237_not ; n33238
g30803 nor pi0055 n33238 ; n33239
g30804 nor n16559 n33239 ; n33240
g30805 and n2529 n33240_not ; n33241
g30806 and n9883 n33197 ; n33242
g30807 and n33241_not n33242 ; n33243
g30808 or n33211 n33243 ; po0352
g30809 and n13132 n16492 ; n33245
g30810 and pi0170_not n9039 ; n33246
g30811 nor n16492 n33246 ; n33247
g30812 and n13130 n33247_not ; n33248
g30813 and pi0232 n33245_not ; n33249
g30814 and n33248_not n33249 ; n33250
g30815 nor n16491 n33250 ; n33251
g30816 and pi0039 n33251_not ; n33252
g30817 and n13910 n16287 ; n33253
g30818 nor pi0039 n33253 ; n33254
g30819 nor pi0038 n33254 ; n33255
g30820 and n33252_not n33255 ; n33256
g30821 and pi0194 n33256_not ; n33257
g30822 and pi0299 n33251_not ; n33258
g30823 nor n11478 n33258 ; n33259
g30824 and pi0039 n33259_not ; n33260
g30825 and n13910 n16275_not ; n33261
g30826 nor pi0039 n33261 ; n33262
g30827 nor pi0038 n33262 ; n33263
g30828 and n33260_not n33263 ; n33264
g30829 nor pi0194 n33264 ; n33265
g30830 and n10197 n33257_not ; n33266
g30831 and n33265_not n33266 ; n33267
g30832 nor pi0196 n33267 ; n33268
g30833 and pi0170_not n9326 ; n33269
g30834 nor n16522 n33269 ; n33270
g30835 and n9036 n33270_not ; n33271
g30836 and n9291 n33271_not ; n33272
g30837 nor n16511 n33272 ; n33273
g30838 and pi0232 n33273_not ; n33274
g30839 nor n16517 n33274 ; n33275
g30840 and pi0232 n16520 ; n33276
g30841 and n33275 n33276_not ; n33277
g30842 and pi0039 n33277_not ; n33278
g30843 and pi0038_not pi0194 ; n33279
g30844 and n33278_not n33279 ; n33280
g30845 and pi0039 n33275_not ; n33281
g30846 nor pi0038 pi0194 ; n33282
g30847 and n33281_not n33282 ; n33283
g30848 nor n33280 n33283 ; n33284
g30849 nor n16536 n33284 ; n33285
g30850 nor n9605 n16274 ; n33286
g30851 and pi0170 n13737 ; n33287
g30852 nor n33286 n33287 ; n33288
g30853 and pi0299 n33288_not ; n33289
g30854 and n16539_not n33280 ; n33290
g30855 and n16533_not n33283 ; n33291
g30856 nor n33290 n33291 ; n33292
g30857 and pi0232 n33289_not ; n33293
g30858 and n33292_not n33293 ; n33294
g30859 nor n33285 n33294 ; n33295
g30860 nor pi0100 n33295 ; n33296
g30861 nor pi0087 n33296 ; n33297
g30862 and n16508 n33297_not ; n33298
g30863 nor pi0092 n33298 ; n33299
g30864 and n16507 n33299_not ; n33300
g30865 nor pi0055 n33300 ; n33301
g30866 nor n16559 n33301 ; n33302
g30867 and n2529 n33302_not ; n33303
g30868 and n9883 n33303_not ; n33304
g30869 and pi0196 n33304_not ; n33305
g30870 nor n33195 n33268 ; n33306
g30871 and n33305_not n33306 ; n33307
g30872 and pi0195 pi0196_not ; n33308
g30873 nor n33267 n33308 ; n33309
g30874 and n33304_not n33308 ; n33310
g30875 and n33195 n33309_not ; n33311
g30876 and n33310_not n33311 ; n33312
g30877 or n33307 n33312 ; po0353
g30878 nor pi0197 n2926 ; n33314
g30879 and pi0767_not pi0947 ; n33315
g30880 and pi0698_not n20902 ; n33316
g30881 nor n33315 n33316 ; n33317
g30882 and n2926 n33317_not ; n33318
g30883 and pi0832 n33314_not ; n33319
g30884 and n33318_not n33319 ; n33320
g30885 nor pi0197 n10197 ; n33321
g30886 and n16641 n33315_not ; n33322
g30887 and pi0197 n17050_not ; n33323
g30888 and pi0038 n33322_not ; n33324
g30889 and n33323_not n33324 ; n33325
g30890 nor pi0197 n16958 ; n33326
g30891 and n16958 n33315 ; n33327
g30892 nor pi0039 n33326 ; n33328
g30893 and n33327_not n33328 ; n33329
g30894 nor pi0197 n21001 ; n33330
g30895 and pi0197 n21162_not ; n33331
g30896 and pi0299 n33331_not ; n33332
g30897 and n33330_not n33332 ; n33333
g30898 nor pi0197 n17024 ; n33334
g30899 and n21019 n33334_not ; n33335
g30900 nor pi0767 n33335 ; n33336
g30901 and n33333_not n33336 ; n33337
g30902 and pi0197_not pi0767 ; n33338
g30903 and n17046_not n33338 ; n33339
g30904 and pi0039 n33339_not ; n33340
g30905 and n33337_not n33340 ; n33341
g30906 nor pi0038 n33329 ; n33342
g30907 and n33341_not n33342 ; n33343
g30908 nor n33325 n33343 ; n33344
g30909 and pi0698 n33344_not ; n33345
g30910 and n21114_not n33329 ; n33346
g30911 and n21111 n33334_not ; n33347
g30912 and pi0197 n21108 ; n33348
g30913 and pi0197_not n21092 ; n33349
g30914 and pi0299 n33348_not ; n33350
g30915 and n33349_not n33350 ; n33351
g30916 and pi0767 n33347_not ; n33352
g30917 and n33351_not n33352 ; n33353
g30918 and pi0197_not n21064 ; n33354
g30919 and pi0197 n21080 ; n33355
g30920 nor pi0767 n33355 ; n33356
g30921 and n33354_not n33356 ; n33357
g30922 and pi0039 n33353_not ; n33358
g30923 and n33357_not n33358 ; n33359
g30924 nor n33346 n33359 ; n33360
g30925 nor pi0038 n33360 ; n33361
g30926 nor pi0197 n16641 ; n33362
g30927 and pi0767 pi0947 ; n33363
g30928 nor pi0039 n33363 ; n33364
g30929 and n21239 n33364 ; n33365
g30930 and pi0038 n33362_not ; n33366
g30931 and n33365_not n33366 ; n33367
g30932 nor pi0698 n33367 ; n33368
g30933 and n33361_not n33368 ; n33369
g30934 nor n33345 n33369 ; n33370
g30935 and n10197 n33370_not ; n33371
g30936 nor pi0832 n33321 ; n33372
g30937 and n33371_not n33372 ; n33373
g30938 nor n33320 n33373 ; po0354
g30939 and n2530 n16958_not ; n33375
g30940 and n18591 n33375_not ; n33376
g30941 and pi0198 n33376_not ; n33377
g30942 and pi0198 n16797_not ; n33378
g30943 and pi0198 n16653_not ; n33379
g30944 nor po1101 n33379 ; n33380
g30945 and n33378 n33380_not ; n33381
g30946 and n6192 n16721_not ; n33382
g30947 nor n6192 n16723 ; n33383
g30948 and pi0198 n33382_not ; n33384
g30949 and n33383_not n33384 ; n33385
g30950 and n6242_not n33385 ; n33386
g30951 nor n33381 n33386 ; n33387
g30952 and pi0215 n33387_not ; n33388
g30953 and n3448 n33379_not ; n33389
g30954 and pi0198 n16684_not ; n33390
g30955 and po1101 n33390_not ; n33391
g30956 nor n33380 n33391 ; n33392
g30957 and n6242 n33392 ; n33393
g30958 and pi0198 n17143_not ; n33394
g30959 and n6242_not n33394 ; n33395
g30960 nor n3448 n33393 ; n33396
g30961 and n33395_not n33396 ; n33397
g30962 nor pi0215 n33389 ; n33398
g30963 and n33397_not n33398 ; n33399
g30964 and pi0299 n33388_not ; n33400
g30965 and n33399_not n33400 ; n33401
g30966 and n6205_not n33385 ; n33402
g30967 nor n33381 n33402 ; n33403
g30968 and pi0223 n33403_not ; n33404
g30969 and n2603 n33379_not ; n33405
g30970 and n6205_not n33394 ; n33406
g30971 and n6205 n33392 ; n33407
g30972 nor n2603 n33407 ; n33408
g30973 and n33406_not n33408 ; n33409
g30974 nor pi0223 n33405 ; n33410
g30975 and n33409_not n33410 ; n33411
g30976 nor pi0299 n33404 ; n33412
g30977 and n33411_not n33412 ; n33413
g30978 and n2571 n10982 ; n33414
g30979 and n33401_not n33414 ; n33415
g30980 and n33413_not n33415 ; n33416
g30981 nor n33377 n33416 ; n33417
g30982 and n19149_not n33417 ; n33418
g30983 and n16639 n33417_not ; n33419
g30984 and pi0198 n2571_not ; n33420
g30985 and pi0039 pi0198 ; n33421
g30986 and pi0038 n33421_not ; n33422
g30987 and pi0198 n16667_not ; n33423
g30988 and pi0634 n16644 ; n33424
g30989 and n16667 n33424 ; n33425
g30990 nor n33423 n33425 ; n33426
g30991 nor pi0039 n33426 ; n33427
g30992 and n33422 n33427_not ; n33428
g30993 and pi0198 n16721 ; n33429
g30994 and pi0634 n16721_not ; n33430
g30995 and n16658 n33430 ; n33431
g30996 nor n33429 n33431 ; n33432
g30997 and n6195 n33432_not ; n33433
g30998 and pi0680_not n33385 ; n33434
g30999 and n6192 n33432 ; n33435
g31000 nor n16658 n33379 ; n33436
g31001 and pi0634 n33436_not ; n33437
g31002 nor n33379 n33437 ; n33438
g31003 and n6197_not n33438 ; n33439
g31004 and n6197 n33432 ; n33440
g31005 nor n33439 n33440 ; n33441
g31006 nor n6192 n33441 ; n33442
g31007 and n17323 n33435_not ; n33443
g31008 and n33442_not n33443 ; n33444
g31009 nor n33433 n33434 ; n33445
g31010 and n33444_not n33445 ; n33446
g31011 and n6205_not n33446 ; n33447
g31012 and n33378 n33434 ; n33448
g31013 and n6197 n33438_not ; n33449
g31014 nor n6197 n33432 ; n33450
g31015 nor n33449 n33450 ; n33451
g31016 and n6192 n33451 ; n33452
g31017 and n6192_not n33438 ; n33453
g31018 and n17323 n33453_not ; n33454
g31019 and n33452_not n33454 ; n33455
g31020 and n6195 n33451_not ; n33456
g31021 nor n33448 n33456 ; n33457
g31022 and n33455_not n33457 ; n33458
g31023 and n6205 n33458 ; n33459
g31024 and pi0223 n33447_not ; n33460
g31025 and n33459_not n33460 ; n33461
g31026 and pi0680 n33437 ; n33462
g31027 nor n33379 n33462 ; n33463
g31028 and n2603 n33463 ; n33464
g31029 and pi0198 n16681 ; n33465
g31030 and pi0634 n16686 ; n33466
g31031 nor n33465 n33466 ; n33467
g31032 nor n6197 n33467 ; n33468
g31033 nor n33449 n33468 ; n33469
g31034 and n6195 n33469_not ; n33470
g31035 and n6192 n33469 ; n33471
g31036 and n33454 n33471_not ; n33472
g31037 nor n6192 n33379 ; n33473
g31038 and n6192 n33390_not ; n33474
g31039 nor pi0680 n33473 ; n33475
g31040 and n33474_not n33475 ; n33476
g31041 nor n33470 n33476 ; n33477
g31042 and n33472_not n33477 ; n33478
g31043 and n6205 n33478_not ; n33479
g31044 and pi0198 n16753 ; n33480
g31045 and n6195 n33467_not ; n33481
g31046 and n6192 n33467 ; n33482
g31047 and n6197 n33467 ; n33483
g31048 nor n33439 n33483 ; n33484
g31049 nor n6192 n33484 ; n33485
g31050 and n17323 n33482_not ; n33486
g31051 and n33485_not n33486 ; n33487
g31052 nor n33480 n33481 ; n33488
g31053 and n33487_not n33488 ; n33489
g31054 nor n6205 n33489 ; n33490
g31055 nor n2603 n33479 ; n33491
g31056 and n33490_not n33491 ; n33492
g31057 nor pi0223 n33464 ; n33493
g31058 and n33492_not n33493 ; n33494
g31059 nor pi0299 n33461 ; n33495
g31060 and n33494_not n33495 ; n33496
g31061 and n6242_not n33446 ; n33497
g31062 and n6242 n33458 ; n33498
g31063 and pi0215 n33497_not ; n33499
g31064 and n33498_not n33499 ; n33500
g31065 and n3448 n33463 ; n33501
g31066 nor n6242 n33489 ; n33502
g31067 and n6242 n33478_not ; n33503
g31068 nor n3448 n33502 ; n33504
g31069 and n33503_not n33504 ; n33505
g31070 nor pi0215 n33501 ; n33506
g31071 and n33505_not n33506 ; n33507
g31072 and pi0299 n33500_not ; n33508
g31073 and n33507_not n33508 ; n33509
g31074 nor n33496 n33509 ; n33510
g31075 and pi0039 n33510_not ; n33511
g31076 and pi0634 pi0680 ; n33512
g31077 and pi0198 n16931 ; n33513
g31078 and n16896_not n33512 ; n33514
g31079 and n33513_not n33514 ; n33515
g31080 nor n16929 n33515 ; n33516
g31081 nor pi0299 n33516 ; n33517
g31082 and pi0198_not n16923 ; n33518
g31083 and pi0198 n16944_not ; n33519
g31084 nor n33518 n33519 ; n33520
g31085 and n33512 n33520_not ; n33521
g31086 and pi0198 n16941_not ; n33522
g31087 and n33512_not n33522 ; n33523
g31088 nor n33521 n33523 ; n33524
g31089 and pi0299 n33524_not ; n33525
g31090 nor pi0039 n33517 ; n33526
g31091 and n33525_not n33526 ; n33527
g31092 nor n33511 n33527 ; n33528
g31093 nor pi0038 n33528 ; n33529
g31094 and n2571 n33428_not ; n33530
g31095 and n33529_not n33530 ; n33531
g31096 nor n33420 n33531 ; n33532
g31097 nor pi0778 n33532 ; n33533
g31098 and pi0625_not n33417 ; n33534
g31099 and pi0625 n33532 ; n33535
g31100 and pi1153 n33534_not ; n33536
g31101 and n33535_not n33536 ; n33537
g31102 and pi0625_not n33532 ; n33538
g31103 and pi0625 n33417 ; n33539
g31104 nor pi1153 n33539 ; n33540
g31105 and n33538_not n33540 ; n33541
g31106 nor n33537 n33541 ; n33542
g31107 and pi0778 n33542_not ; n33543
g31108 nor n33533 n33543 ; n33544
g31109 and n17075_not n33544 ; n33545
g31110 and n17075 n33417 ; n33546
g31111 nor n33545 n33546 ; n33547
g31112 and n16639_not n33547 ; n33548
g31113 nor n33419 n33548 ; n33549
g31114 and n16635_not n33549 ; n33550
g31115 and n16631_not n33550 ; n33551
g31116 nor n33418 n33551 ; n33552
g31117 and pi0792_not n33552 ; n33553
g31118 and pi0628 n33552_not ; n33554
g31119 and pi0628_not n33417 ; n33555
g31120 nor n33554 n33555 ; n33556
g31121 and pi1156 n33556 ; n33557
g31122 and pi0628 n33417 ; n33558
g31123 nor pi0628 n33552 ; n33559
g31124 nor pi1156 n33558 ; n33560
g31125 and n33559_not n33560 ; n33561
g31126 nor n33557 n33561 ; n33562
g31127 and pi0792 n33562_not ; n33563
g31128 nor n33553 n33563 ; n33564
g31129 and pi0647_not n33564 ; n33565
g31130 and pi0647 n33417 ; n33566
g31131 nor pi1157 n33566 ; n33567
g31132 and n33565_not n33567 ; n33568
g31133 and pi0630 n33568 ; n33569
g31134 and n17779 n33417_not ; n33570
g31135 nor n17127 n17131 ; n33571
g31136 and pi0633 n33571_not ; n33572
g31137 nor n16929 n33572 ; n33573
g31138 nor n17136 n33573 ; n33574
g31139 and pi0299_not n33574 ; n33575
g31140 and pi0603 pi0633 ; n33576
g31141 nor n33522 n33576 ; n33577
g31142 and pi0198 n17122_not ; n33578
g31143 and pi0198_not n17230 ; n33579
g31144 nor n33578 n33579 ; n33580
g31145 and n33576 n33580 ; n33581
g31146 nor n33577 n33581 ; n33582
g31147 and pi0299 n33582 ; n33583
g31148 nor pi0039 n33575 ; n33584
g31149 and n33583_not n33584 ; n33585
g31150 and pi0633 n17239 ; n33586
g31151 nor n33385 n33586 ; n33587
g31152 nor n6195 n33587 ; n33588
g31153 and pi0633 n16653 ; n33589
g31154 and n17144_not n33589 ; n33590
g31155 and n16721_not n33590 ; n33591
g31156 nor n33429 n33591 ; n33592
g31157 and n17188 n33592_not ; n33593
g31158 nor n33588 n33593 ; n33594
g31159 and n6205_not n33594 ; n33595
g31160 nor n33379 n33590 ; n33596
g31161 and pi0603 n33596_not ; n33597
g31162 and pi0603_not n33379 ; n33598
g31163 nor n33597 n33598 ; n33599
g31164 and n17167_not n33599 ; n33600
g31165 and n6197 n33596_not ; n33601
g31166 nor n33378 n33591 ; n33602
g31167 and n33601_not n33602 ; n33603
g31168 and pi0603 n33603_not ; n33604
g31169 and n17167 n33598_not ; n33605
g31170 and n33604_not n33605 ; n33606
g31171 nor n33600 n33606 ; n33607
g31172 and n6195_not n33607 ; n33608
g31173 nor n33378 n33604 ; n33609
g31174 and n6195 n33609_not ; n33610
g31175 nor n33608 n33610 ; n33611
g31176 and n6205 n33611 ; n33612
g31177 and pi0223 n33595_not ; n33613
g31178 and n33612_not n33613 ; n33614
g31179 and n2603 n33599 ; n33615
g31180 and pi0642 n33597_not ; n33616
g31181 and pi0633 n17147 ; n33617
g31182 nor n33465 n33617 ; n33618
g31183 nor n6197 n33618 ; n33619
g31184 nor n33601 n33619 ; n33620
g31185 and pi0603 n33620_not ; n33621
g31186 nor pi0642 n33621 ; n33622
g31187 and n6191 n33616_not ; n33623
g31188 and n33622_not n33623 ; n33624
g31189 and n6191_not n33597 ; n33625
g31190 nor n33598 n33625 ; n33626
g31191 and n33624_not n33626 ; n33627
g31192 and n6195_not n33627 ; n33628
g31193 and pi0603_not n33390 ; n33629
g31194 and n6195 n33629_not ; n33630
g31195 and n33621_not n33630 ; n33631
g31196 nor n33628 n33631 ; n33632
g31197 and n6205 n33632 ; n33633
g31198 and pi0603 n33618_not ; n33634
g31199 and n17167 n33634 ; n33635
g31200 and pi0198 n17149 ; n33636
g31201 and n6197 n33618 ; n33637
g31202 and n6197_not n33596 ; n33638
g31203 and pi0603 n17167_not ; n33639
g31204 and n33638_not n33639 ; n33640
g31205 and n33637_not n33640 ; n33641
g31206 nor n33635 n33636 ; n33642
g31207 and n33641_not n33642 ; n33643
g31208 and n6195_not n33643 ; n33644
g31209 and n6195 n33465_not ; n33645
g31210 and n33634_not n33645 ; n33646
g31211 nor n33644 n33646 ; n33647
g31212 and n6205_not n33647 ; n33648
g31213 nor n2603 n33648 ; n33649
g31214 and n33633_not n33649 ; n33650
g31215 nor pi0223 n33615 ; n33651
g31216 and n33650_not n33651 ; n33652
g31217 nor n33614 n33652 ; n33653
g31218 nor pi0299 n33653 ; n33654
g31219 and n6242_not n33594 ; n33655
g31220 and n6242 n33611 ; n33656
g31221 and pi0215 n33655_not ; n33657
g31222 and n33656_not n33657 ; n33658
g31223 and n3448 n33599 ; n33659
g31224 and n6242_not n33647 ; n33660
g31225 and n6242 n33632 ; n33661
g31226 nor n3448 n33660 ; n33662
g31227 and n33661_not n33662 ; n33663
g31228 nor pi0215 n33659 ; n33664
g31229 and n33663_not n33664 ; n33665
g31230 nor n33658 n33665 ; n33666
g31231 and pi0299 n33666_not ; n33667
g31232 and pi0039 n33654_not ; n33668
g31233 and n33667_not n33668 ; n33669
g31234 nor n33585 n33669 ; n33670
g31235 nor pi0038 n33670 ; n33671
g31236 and pi0633 n17168 ; n33672
g31237 and n16667 n33672 ; n33673
g31238 nor n33423 n33673 ; n33674
g31239 nor pi0039 n33674 ; n33675
g31240 and n33422 n33675_not ; n33676
g31241 and n2571 n33676_not ; n33677
g31242 and n33671_not n33677 ; n33678
g31243 nor n33420 n33678 ; n33679
g31244 nor n17117 n33679 ; n33680
g31245 and n17117 n33417_not ; n33681
g31246 nor n33680 n33681 ; n33682
g31247 nor pi0785 n33682 ; n33683
g31248 nor n17291 n33417 ; n33684
g31249 and pi0609 n33680 ; n33685
g31250 nor n33684 n33685 ; n33686
g31251 and pi1155 n33686_not ; n33687
g31252 nor n17296 n33417 ; n33688
g31253 and pi0609_not n33680 ; n33689
g31254 nor n33688 n33689 ; n33690
g31255 nor pi1155 n33690 ; n33691
g31256 nor n33687 n33691 ; n33692
g31257 and pi0785 n33692_not ; n33693
g31258 nor n33683 n33693 ; n33694
g31259 nor pi0781 n33694 ; n33695
g31260 and pi0618_not n33417 ; n33696
g31261 and pi0618 n33694 ; n33697
g31262 and pi1154 n33696_not ; n33698
g31263 and n33697_not n33698 ; n33699
g31264 and pi0618_not n33694 ; n33700
g31265 and pi0618 n33417 ; n33701
g31266 nor pi1154 n33701 ; n33702
g31267 and n33700_not n33702 ; n33703
g31268 nor n33699 n33703 ; n33704
g31269 and pi0781 n33704_not ; n33705
g31270 nor n33695 n33705 ; n33706
g31271 nor pi0789 n33706 ; n33707
g31272 and pi0619_not n33417 ; n33708
g31273 and pi0619 n33706 ; n33709
g31274 and pi1159 n33708_not ; n33710
g31275 and n33709_not n33710 ; n33711
g31276 and pi0619_not n33706 ; n33712
g31277 and pi0619 n33417 ; n33713
g31278 nor pi1159 n33713 ; n33714
g31279 and n33712_not n33714 ; n33715
g31280 nor n33711 n33715 ; n33716
g31281 and pi0789 n33716_not ; n33717
g31282 nor n33707 n33717 ; n33718
g31283 and n17969_not n33718 ; n33719
g31284 and n17969 n33417 ; n33720
g31285 nor n33719 n33720 ; n33721
g31286 and n17779_not n33721 ; n33722
g31287 nor n33570 n33722 ; n33723
g31288 nor n20559 n33723 ; n33724
g31289 and pi0647 n33564_not ; n33725
g31290 nor pi0647 n33417 ; n33726
g31291 nor n33725 n33726 ; n33727
g31292 and n17801 n33727_not ; n33728
g31293 nor n33569 n33728 ; n33729
g31294 and n33724_not n33729 ; n33730
g31295 and pi0787 n33730_not ; n33731
g31296 and pi0629 n33561 ; n33732
g31297 and n20570_not n33721 ; n33733
g31298 and n17776 n33556 ; n33734
g31299 nor n33732 n33734 ; n33735
g31300 and n33733_not n33735 ; n33736
g31301 and pi0792 n33736_not ; n33737
g31302 and n16635 n33417 ; n33738
g31303 nor n33550 n33738 ; n33739
g31304 and n17871 n33739_not ; n33740
g31305 nor pi0626 n33718 ; n33741
g31306 and pi0626 n33417_not ; n33742
g31307 and n16629 n33742_not ; n33743
g31308 and n33741_not n33743 ; n33744
g31309 and pi0626 n33718_not ; n33745
g31310 nor pi0626 n33417 ; n33746
g31311 and n16628 n33746_not ; n33747
g31312 and n33745_not n33747 ; n33748
g31313 nor n33740 n33744 ; n33749
g31314 and n33748_not n33749 ; n33750
g31315 and pi0788 n33750_not ; n33751
g31316 and pi0609 n33544 ; n33752
g31317 and pi0634 n17645 ; n33753
g31318 and n33674 n33753_not ; n33754
g31319 nor pi0039 n33754 ; n33755
g31320 and n33422 n33755_not ; n33756
g31321 and n33512_not n33582 ; n33757
g31322 nor pi0603 n33520 ; n33758
g31323 nor pi0198 pi0665 ; n33759
g31324 and n17122 n33759 ; n33760
g31325 and n17230_not n33519 ; n33761
g31326 nor pi0633 n33760 ; n33762
g31327 and n33761_not n33762 ; n33763
g31328 and pi0198 pi0665_not ; n33764
g31329 and pi0633 n33764_not ; n33765
g31330 and n33518_not n33765 ; n33766
g31331 and n33580 n33766 ; n33767
g31332 and pi0603 n33763_not ; n33768
g31333 and n33767_not n33768 ; n33769
g31334 nor n33758 n33769 ; n33770
g31335 and n33512 n33770_not ; n33771
g31336 and pi0299 n33757_not ; n33772
g31337 and n33771_not n33772 ; n33773
g31338 and pi0680_not n33574 ; n33774
g31339 and pi0603_not n33516 ; n33775
g31340 and pi0198 pi0633_not ; n33776
g31341 and pi0634 pi0665_not ; n33777
g31342 and n33776_not n33777 ; n33778
g31343 and n17126_not n33778 ; n33779
g31344 and pi0634_not n16929 ; n33780
g31345 and pi0634 n16932 ; n33781
g31346 and n17133_not n33781 ; n33782
g31347 nor n33780 n33782 ; n33783
g31348 nor pi0633 n33783 ; n33784
g31349 and pi0603 n33779_not ; n33785
g31350 and n33572_not n33785 ; n33786
g31351 and n33784_not n33786 ; n33787
g31352 and pi0680 n33775_not ; n33788
g31353 and n33787_not n33788 ; n33789
g31354 nor pi0299 n33774 ; n33790
g31355 and n33789_not n33790 ; n33791
g31356 nor n33773 n33791 ; n33792
g31357 nor pi0039 n33792 ; n33793
g31358 and n17355 n33437 ; n33794
g31359 and n33599 n33794_not ; n33795
g31360 and n2603 n33795 ; n33796
g31361 and pi0680_not n33627 ; n33797
g31362 nor pi0603 n33438 ; n33798
g31363 and n17159 n33777 ; n33799
g31364 and n33596 n33799_not ; n33800
g31365 and pi0603 n33800_not ; n33801
g31366 nor n33798 n33801 ; n33802
g31367 nor n6191 n33802 ; n33803
g31368 and n6197 n33800_not ; n33804
g31369 and pi0634 n17424 ; n33805
g31370 and n33618 n33805_not ; n33806
g31371 nor n6197 n33806 ; n33807
g31372 nor n33804 n33807 ; n33808
g31373 and pi0603 n33808_not ; n33809
g31374 and pi0642_not n33809 ; n33810
g31375 and pi0642 n33801 ; n33811
g31376 nor n33798 n33811 ; n33812
g31377 and n33810_not n33812 ; n33813
g31378 and n6191 n33813_not ; n33814
g31379 nor n16657 n33803 ; n33815
g31380 and n33814_not n33815 ; n33816
g31381 nor pi0603 n33469 ; n33817
g31382 and n16657 n33817_not ; n33818
g31383 and n33809_not n33818 ; n33819
g31384 nor n33816 n33819 ; n33820
g31385 and pi0680 n33820_not ; n33821
g31386 nor n33797 n33821 ; n33822
g31387 and n6205 n33822 ; n33823
g31388 nor pi0680 n33643 ; n33824
g31389 and pi0603_not n33484 ; n33825
g31390 and n17167_not n33801 ; n33826
g31391 nor n33640 n33826 ; n33827
g31392 and n6192_not n33827 ; n33828
g31393 nor n6197 n33827 ; n33829
g31394 and n33806 n33829_not ; n33830
g31395 nor n33828 n33830 ; n33831
g31396 nor n33825 n33831 ; n33832
g31397 and n17323 n33832_not ; n33833
g31398 nor n17168 n33467 ; n33834
g31399 nor n33634 n33834 ; n33835
g31400 and n6195 n33835_not ; n33836
g31401 nor n33824 n33836 ; n33837
g31402 and n33833_not n33837 ; n33838
g31403 nor n6205 n33838 ; n33839
g31404 nor n2603 n33839 ; n33840
g31405 and n33823_not n33840 ; n33841
g31406 nor pi0223 n33796 ; n33842
g31407 and n33841_not n33842 ; n33843
g31408 nor pi0680 n33587 ; n33844
g31409 and n17191 n33759 ; n33845
g31410 and n17144 n33764 ; n33846
g31411 nor n33429 n33846 ; n33847
g31412 and n33845_not n33847 ; n33848
g31413 and pi0634 n33848_not ; n33849
g31414 and pi0634_not n33429 ; n33850
g31415 nor n33591 n33850 ; n33851
g31416 and n33849_not n33851 ; n33852
g31417 and pi0603 n33852_not ; n33853
g31418 nor pi0603 n33432 ; n33854
g31419 nor n33853 n33854 ; n33855
g31420 and n6195 n33855_not ; n33856
g31421 and n17167 n33853 ; n33857
g31422 and pi0603_not n33441 ; n33858
g31423 nor n33827 n33852 ; n33859
g31424 nor n33829 n33858 ; n33860
g31425 nor n33857 n33859 ; n33861
g31426 and n33860 n33861 ; n33862
g31427 and n17323 n33862_not ; n33863
g31428 nor n33844 n33856 ; n33864
g31429 and n33863_not n33864 ; n33865
g31430 and n6205_not n33865 ; n33866
g31431 and pi0680_not n33607 ; n33867
g31432 nor n6197 n33852 ; n33868
g31433 nor n33804 n33868 ; n33869
g31434 and pi0603 n33869_not ; n33870
g31435 nor pi0603 n33451 ; n33871
g31436 nor n33870 n33871 ; n33872
g31437 and n6195 n33872_not ; n33873
g31438 and n17167_not n33802 ; n33874
g31439 and n17167 n33798_not ; n33875
g31440 and n33870_not n33875 ; n33876
g31441 and n17323 n33874_not ; n33877
g31442 and n33876_not n33877 ; n33878
g31443 nor n33867 n33873 ; n33879
g31444 and n33878_not n33879 ; n33880
g31445 and n6205 n33880 ; n33881
g31446 and pi0223 n33866_not ; n33882
g31447 and n33881_not n33882 ; n33883
g31448 nor n33843 n33883 ; n33884
g31449 nor pi0299 n33884 ; n33885
g31450 and n3448 n33795 ; n33886
g31451 and n6242 n33822 ; n33887
g31452 nor n6242 n33838 ; n33888
g31453 nor n3448 n33888 ; n33889
g31454 and n33887_not n33889 ; n33890
g31455 nor pi0215 n33886 ; n33891
g31456 and n33890_not n33891 ; n33892
g31457 and n6242_not n33865 ; n33893
g31458 and n6242 n33880 ; n33894
g31459 and pi0215 n33893_not ; n33895
g31460 and n33894_not n33895 ; n33896
g31461 nor n33892 n33896 ; n33897
g31462 and pi0299 n33897_not ; n33898
g31463 and pi0039 n33885_not ; n33899
g31464 and n33898_not n33899 ; n33900
g31465 nor n33793 n33900 ; n33901
g31466 nor pi0038 n33901 ; n33902
g31467 and n2571 n33756_not ; n33903
g31468 and n33902_not n33903 ; n33904
g31469 nor n33420 n33904 ; n33905
g31470 and pi0625_not n33905 ; n33906
g31471 and pi0625 n33679 ; n33907
g31472 nor pi1153 n33907 ; n33908
g31473 and n33906_not n33908 ; n33909
g31474 nor pi0608 n33537 ; n33910
g31475 and n33909_not n33910 ; n33911
g31476 and pi0625_not n33679 ; n33912
g31477 and pi0625 n33905 ; n33913
g31478 and pi1153 n33912_not ; n33914
g31479 and n33913_not n33914 ; n33915
g31480 and pi0608 n33541_not ; n33916
g31481 and n33915_not n33916 ; n33917
g31482 nor n33911 n33917 ; n33918
g31483 and pi0778 n33918_not ; n33919
g31484 and pi0778_not n33905 ; n33920
g31485 nor n33919 n33920 ; n33921
g31486 nor pi0609 n33921 ; n33922
g31487 nor pi1155 n33752 ; n33923
g31488 and n33922_not n33923 ; n33924
g31489 nor pi0660 n33687 ; n33925
g31490 and n33924_not n33925 ; n33926
g31491 and pi0609_not n33544 ; n33927
g31492 and pi0609 n33921_not ; n33928
g31493 and pi1155 n33927_not ; n33929
g31494 and n33928_not n33929 ; n33930
g31495 and pi0660 n33691_not ; n33931
g31496 and n33930_not n33931 ; n33932
g31497 nor n33926 n33932 ; n33933
g31498 and pi0785 n33933_not ; n33934
g31499 nor pi0785 n33921 ; n33935
g31500 nor n33934 n33935 ; n33936
g31501 nor pi0618 n33936 ; n33937
g31502 and pi0618 n33547_not ; n33938
g31503 nor pi1154 n33938 ; n33939
g31504 and n33937_not n33939 ; n33940
g31505 nor pi0627 n33699 ; n33941
g31506 and n33940_not n33941 ; n33942
g31507 and pi0618 n33936_not ; n33943
g31508 nor pi0618 n33547 ; n33944
g31509 and pi1154 n33944_not ; n33945
g31510 and n33943_not n33945 ; n33946
g31511 and pi0627 n33703_not ; n33947
g31512 and n33946_not n33947 ; n33948
g31513 nor n33942 n33948 ; n33949
g31514 and pi0781 n33949_not ; n33950
g31515 nor pi0781 n33936 ; n33951
g31516 nor n33950 n33951 ; n33952
g31517 and pi0789_not n33952 ; n33953
g31518 nor pi0619 n33952 ; n33954
g31519 and pi0619 n33549 ; n33955
g31520 nor pi1159 n33955 ; n33956
g31521 and n33954_not n33956 ; n33957
g31522 nor pi0648 n33711 ; n33958
g31523 and n33957_not n33958 ; n33959
g31524 and pi0619_not n33549 ; n33960
g31525 and pi0619 n33952_not ; n33961
g31526 and pi1159 n33960_not ; n33962
g31527 and n33961_not n33962 ; n33963
g31528 and pi0648 n33715_not ; n33964
g31529 and n33963_not n33964 ; n33965
g31530 and pi0789 n33959_not ; n33966
g31531 and n33965_not n33966 ; n33967
g31532 and n17970 n33953_not ; n33968
g31533 and n33967_not n33968 ; n33969
g31534 nor n33751 n33969 ; n33970
g31535 nor n33737 n33970 ; n33971
g31536 and n20364 n33736 ; n33972
g31537 nor n20206 n33972 ; n33973
g31538 and n33971_not n33973 ; n33974
g31539 nor n33731 n33974 ; n33975
g31540 nor pi0790 n33975 ; n33976
g31541 nor pi0787 n33564 ; n33977
g31542 and pi1157 n33727_not ; n33978
g31543 nor n33568 n33978 ; n33979
g31544 and pi0787 n33979_not ; n33980
g31545 nor n33977 n33980 ; n33981
g31546 and pi0644_not n33981 ; n33982
g31547 and pi0644 n33975 ; n33983
g31548 and pi0715 n33982_not ; n33984
g31549 and n33983_not n33984 ; n33985
g31550 and n17804_not n33723 ; n33986
g31551 and n17804 n33417 ; n33987
g31552 nor n33986 n33987 ; n33988
g31553 and pi0644 n33988_not ; n33989
g31554 and pi0644_not n33417 ; n33990
g31555 nor pi0715 n33990 ; n33991
g31556 and n33989_not n33991 ; n33992
g31557 and pi1160 n33992_not ; n33993
g31558 and n33985_not n33993 ; n33994
g31559 nor pi0644 n33988 ; n33995
g31560 and pi0644 n33417 ; n33996
g31561 and pi0715 n33996_not ; n33997
g31562 and n33995_not n33997 ; n33998
g31563 and pi0644 n33981 ; n33999
g31564 and pi0644_not n33975 ; n34000
g31565 nor pi0715 n33999 ; n34001
g31566 and n34000_not n34001 ; n34002
g31567 nor pi1160 n33998 ; n34003
g31568 and n34002_not n34003 ; n34004
g31569 and pi0790 n33994_not ; n34005
g31570 and n34004_not n34005 ; n34006
g31571 nor n33976 n34006 ; n34007
g31572 nor po1038 n34007 ; n34008
g31573 and pi0198 po1038 ; n34009
g31574 or n34008 n34009 ; po0355
g31575 and pi0199 n17059_not ; n34011
g31576 nor pi0619 n34011 ; n34012
g31577 nor pi0617 n34011 ; n34013
g31578 nor pi0199 n19432 ; n34014
g31579 and n19438 n34014_not ; n34015
g31580 nor pi0199 n17275 ; n34016
g31581 and pi0199 n17221 ; n34017
g31582 nor pi0038 n34016 ; n34018
g31583 and n34017_not n34018 ; n34019
g31584 nor n34015 n34019 ; n34020
g31585 and n2571 n34020_not ; n34021
g31586 and pi0199 n2571_not ; n34022
g31587 and pi0617 n34022_not ; n34023
g31588 and n34021_not n34023 ; n34024
g31589 nor n34013 n34024 ; n34025
g31590 nor n17117 n34025 ; n34026
g31591 and n17117 n34011_not ; n34027
g31592 nor n34026 n34027 ; n34028
g31593 and pi0785_not n34028 ; n34029
g31594 nor pi0609 n34011 ; n34030
g31595 and pi0609 n34028_not ; n34031
g31596 and pi1155 n34030_not ; n34032
g31597 and n34031_not n34032 ; n34033
g31598 nor pi0609 n34028 ; n34034
g31599 and pi0609 n34011_not ; n34035
g31600 nor pi1155 n34035 ; n34036
g31601 and n34034_not n34036 ; n34037
g31602 nor n34033 n34037 ; n34038
g31603 and pi0785 n34038_not ; n34039
g31604 nor n34029 n34039 ; n34040
g31605 nor pi0781 n34040 ; n34041
g31606 nor pi0618 n34011 ; n34042
g31607 and pi0618 n34040 ; n34043
g31608 and pi1154 n34042_not ; n34044
g31609 and n34043_not n34044 ; n34045
g31610 and pi0618 n34011_not ; n34046
g31611 and pi0618_not n34040 ; n34047
g31612 nor pi1154 n34046 ; n34048
g31613 and n34047_not n34048 ; n34049
g31614 nor n34045 n34049 ; n34050
g31615 and pi0781 n34050_not ; n34051
g31616 nor n34041 n34051 ; n34052
g31617 and pi0619 n34052 ; n34053
g31618 and pi1159 n34012_not ; n34054
g31619 and n34053_not n34054 ; n34055
g31620 nor pi0625 n34011 ; n34056
g31621 nor pi0637 n34011 ; n34057
g31622 nor pi0199 n16641 ; n34058
g31623 and n19899 n34058_not ; n34059
g31624 and pi0199 n16840_not ; n34060
g31625 nor pi0199 n16749 ; n34061
g31626 and pi0039 n34061_not ; n34062
g31627 and n34060_not n34062 ; n34063
g31628 and pi0199 n16948_not ; n34064
g31629 and pi0199_not n16926 ; n34065
g31630 nor pi0039 n34064 ; n34066
g31631 and n34065_not n34066 ; n34067
g31632 nor pi0038 n34067 ; n34068
g31633 and n34063_not n34068 ; n34069
g31634 nor n34059 n34069 ; n34070
g31635 and n2571 n34070_not ; n34071
g31636 and pi0637 n34022_not ; n34072
g31637 and n34071_not n34072 ; n34073
g31638 nor n34057 n34073 ; n34074
g31639 and pi0625 n34074_not ; n34075
g31640 and pi1153 n34056_not ; n34076
g31641 and n34075_not n34076 ; n34077
g31642 and pi0637_not n34025 ; n34078
g31643 and pi0199 n19476 ; n34079
g31644 and n2571 n24549_not ; n34080
g31645 nor pi0199 n34080 ; n34081
g31646 nor pi0617 n19472 ; n34082
g31647 and n34081_not n34082 ; n34083
g31648 and n34079_not n34083 ; n34084
g31649 and n2571 n19496 ; n34085
g31650 nor pi0199 n34085 ; n34086
g31651 and pi0199 n19488 ; n34087
g31652 and pi0617 n34087_not ; n34088
g31653 and n34086_not n34088 ; n34089
g31654 nor n34022 n34089 ; n34090
g31655 and n34084_not n34090 ; n34091
g31656 and pi0637 n34091_not ; n34092
g31657 nor n34078 n34092 ; n34093
g31658 and pi0625_not n34093 ; n34094
g31659 and pi0625 n34025_not ; n34095
g31660 nor pi1153 n34095 ; n34096
g31661 and n34094_not n34096 ; n34097
g31662 nor pi0608 n34077 ; n34098
g31663 and n34097_not n34098 ; n34099
g31664 nor pi0625 n34074 ; n34100
g31665 and pi0625 n34011_not ; n34101
g31666 nor pi1153 n34101 ; n34102
g31667 and n34100_not n34102 ; n34103
g31668 and pi0625 n34093 ; n34104
g31669 nor pi0625 n34025 ; n34105
g31670 and pi1153 n34105_not ; n34106
g31671 and n34104_not n34106 ; n34107
g31672 and pi0608 n34103_not ; n34108
g31673 and n34107_not n34108 ; n34109
g31674 nor n34099 n34109 ; n34110
g31675 and pi0778 n34110_not ; n34111
g31676 and pi0778_not n34093 ; n34112
g31677 nor n34111 n34112 ; n34113
g31678 nor pi0609 n34113 ; n34114
g31679 and pi0778_not n34074 ; n34115
g31680 nor n34077 n34103 ; n34116
g31681 and pi0778 n34116_not ; n34117
g31682 nor n34115 n34117 ; n34118
g31683 and pi0609 n34118 ; n34119
g31684 nor pi1155 n34119 ; n34120
g31685 and n34114_not n34120 ; n34121
g31686 nor pi0660 n34033 ; n34122
g31687 and n34121_not n34122 ; n34123
g31688 and pi0609_not n34118 ; n34124
g31689 and pi0609 n34113_not ; n34125
g31690 and pi1155 n34124_not ; n34126
g31691 and n34125_not n34126 ; n34127
g31692 and pi0660 n34037_not ; n34128
g31693 and n34127_not n34128 ; n34129
g31694 nor n34123 n34129 ; n34130
g31695 and pi0785 n34130_not ; n34131
g31696 nor pi0785 n34113 ; n34132
g31697 nor n34131 n34132 ; n34133
g31698 nor pi0618 n34133 ; n34134
g31699 and n17075 n34011_not ; n34135
g31700 and n17075_not n34118 ; n34136
g31701 nor n34135 n34136 ; n34137
g31702 and pi0618 n34137_not ; n34138
g31703 nor pi1154 n34138 ; n34139
g31704 and n34134_not n34139 ; n34140
g31705 nor pi0627 n34045 ; n34141
g31706 and n34140_not n34141 ; n34142
g31707 and pi0618 n34133_not ; n34143
g31708 nor pi0618 n34137 ; n34144
g31709 and pi1154 n34144_not ; n34145
g31710 and n34143_not n34145 ; n34146
g31711 and pi0627 n34049_not ; n34147
g31712 and n34146_not n34147 ; n34148
g31713 nor n34142 n34148 ; n34149
g31714 and pi0781 n34149_not ; n34150
g31715 nor pi0781 n34133 ; n34151
g31716 nor n34150 n34151 ; n34152
g31717 nor pi0619 n34152 ; n34153
g31718 and n16639_not n34137 ; n34154
g31719 and n16639 n34011 ; n34155
g31720 nor n34154 n34155 ; n34156
g31721 and pi0619 n34156 ; n34157
g31722 nor pi1159 n34157 ; n34158
g31723 and n34153_not n34158 ; n34159
g31724 nor pi0648 n34055 ; n34160
g31725 and n34159_not n34160 ; n34161
g31726 and pi0619 n34011_not ; n34162
g31727 and pi0619_not n34052 ; n34163
g31728 nor pi1159 n34162 ; n34164
g31729 and n34163_not n34164 ; n34165
g31730 and pi0619_not n34156 ; n34166
g31731 and pi0619 n34152_not ; n34167
g31732 and pi1159 n34166_not ; n34168
g31733 and n34167_not n34168 ; n34169
g31734 and pi0648 n34165_not ; n34170
g31735 and n34169_not n34170 ; n34171
g31736 nor n34161 n34171 ; n34172
g31737 and pi0789 n34172_not ; n34173
g31738 nor pi0789 n34152 ; n34174
g31739 nor n34173 n34174 ; n34175
g31740 and pi0788_not n34175 ; n34176
g31741 and pi0626_not n34175 ; n34177
g31742 and n16635 n34011_not ; n34178
g31743 and n16635_not n34156 ; n34179
g31744 nor n34178 n34179 ; n34180
g31745 and pi0626 n34180 ; n34181
g31746 nor pi0641 n34181 ; n34182
g31747 and n34177_not n34182 ; n34183
g31748 nor pi0789 n34052 ; n34184
g31749 nor n34055 n34165 ; n34185
g31750 and pi0789 n34185_not ; n34186
g31751 nor n34184 n34186 ; n34187
g31752 nor pi0626 n34187 ; n34188
g31753 and pi0626 n34011 ; n34189
g31754 and pi0641 n34189_not ; n34190
g31755 and n34188_not n34190 ; n34191
g31756 nor pi1158 n34191 ; n34192
g31757 and n34183_not n34192 ; n34193
g31758 and pi0626_not n34180 ; n34194
g31759 and pi0626 n34175 ; n34195
g31760 and pi0641 n34194_not ; n34196
g31761 and n34195_not n34196 ; n34197
g31762 and pi0626 n34187_not ; n34198
g31763 and pi0626_not n34011 ; n34199
g31764 nor pi0641 n34199 ; n34200
g31765 and n34198_not n34200 ; n34201
g31766 and pi1158 n34201_not ; n34202
g31767 and n34197_not n34202 ; n34203
g31768 nor n34193 n34203 ; n34204
g31769 and pi0788 n34204_not ; n34205
g31770 nor n34176 n34205 ; n34206
g31771 and pi0628_not n34206 ; n34207
g31772 nor n17969 n34187 ; n34208
g31773 and n17969 n34011 ; n34209
g31774 nor n34208 n34209 ; n34210
g31775 and pi0628 n34210 ; n34211
g31776 nor pi1156 n34211 ; n34212
g31777 and n34207_not n34212 ; n34213
g31778 nor pi0628 n34011 ; n34214
g31779 and n16631_not n34180 ; n34215
g31780 and n16631 n34011 ; n34216
g31781 nor n34215 n34216 ; n34217
g31782 and pi0628 n34217 ; n34218
g31783 and pi1156 n34214_not ; n34219
g31784 and n34218_not n34219 ; n34220
g31785 nor pi0629 n34220 ; n34221
g31786 and n34213_not n34221 ; n34222
g31787 and pi0628 n34206 ; n34223
g31788 and pi0628_not n34210 ; n34224
g31789 and pi1156 n34224_not ; n34225
g31790 and n34223_not n34225 ; n34226
g31791 and pi0628 n34011_not ; n34227
g31792 and pi0628_not n34217 ; n34228
g31793 nor pi1156 n34227 ; n34229
g31794 and n34228_not n34229 ; n34230
g31795 and pi0629 n34230_not ; n34231
g31796 and n34226_not n34231 ; n34232
g31797 nor n34222 n34232 ; n34233
g31798 and pi0792 n34233_not ; n34234
g31799 and pi0792_not n34206 ; n34235
g31800 nor n34234 n34235 ; n34236
g31801 nor pi0647 n34236 ; n34237
g31802 nor n17779 n34210 ; n34238
g31803 and n17779 n34011 ; n34239
g31804 nor n34238 n34239 ; n34240
g31805 and pi0647 n34240 ; n34241
g31806 nor pi1157 n34241 ; n34242
g31807 and n34237_not n34242 ; n34243
g31808 nor pi0647 n34011 ; n34244
g31809 nor pi0792 n34217 ; n34245
g31810 nor n34220 n34230 ; n34246
g31811 and pi0792 n34246_not ; n34247
g31812 nor n34245 n34247 ; n34248
g31813 and pi0647 n34248 ; n34249
g31814 and pi1157 n34244_not ; n34250
g31815 and n34249_not n34250 ; n34251
g31816 nor pi0630 n34251 ; n34252
g31817 and n34243_not n34252 ; n34253
g31818 and pi0647 n34236_not ; n34254
g31819 and pi0647_not n34240 ; n34255
g31820 and pi1157 n34255_not ; n34256
g31821 and n34254_not n34256 ; n34257
g31822 and pi0647 n34011_not ; n34258
g31823 and pi0647_not n34248 ; n34259
g31824 nor pi1157 n34258 ; n34260
g31825 and n34259_not n34260 ; n34261
g31826 and pi0630 n34261_not ; n34262
g31827 and n34257_not n34262 ; n34263
g31828 nor n34253 n34263 ; n34264
g31829 and pi0787 n34264_not ; n34265
g31830 nor pi0787 n34236 ; n34266
g31831 nor n34265 n34266 ; n34267
g31832 and pi0790_not n34267 ; n34268
g31833 nor pi0787 n34248 ; n34269
g31834 nor n34251 n34261 ; n34270
g31835 and pi0787 n34270_not ; n34271
g31836 nor n34269 n34271 ; n34272
g31837 and pi0644_not n34272 ; n34273
g31838 and pi0644 n34267_not ; n34274
g31839 and pi0715 n34273_not ; n34275
g31840 and n34274_not n34275 ; n34276
g31841 and n17804 n34011_not ; n34277
g31842 and n17804_not n34240 ; n34278
g31843 nor n34277 n34278 ; n34279
g31844 and pi0644 n34279_not ; n34280
g31845 nor pi0644 n34011 ; n34281
g31846 nor pi0715 n34281 ; n34282
g31847 and n34280_not n34282 ; n34283
g31848 and pi1160 n34283_not ; n34284
g31849 and n34276_not n34284 ; n34285
g31850 nor pi0644 n34267 ; n34286
g31851 and pi0644 n34272 ; n34287
g31852 nor pi0715 n34287 ; n34288
g31853 and n34286_not n34288 ; n34289
g31854 nor pi0644 n34279 ; n34290
g31855 and pi0644 n34011_not ; n34291
g31856 and pi0715 n34291_not ; n34292
g31857 and n34290_not n34292 ; n34293
g31858 nor pi1160 n34293 ; n34294
g31859 and n34289_not n34294 ; n34295
g31860 and pi0790 n34285_not ; n34296
g31861 and n34295_not n34296 ; n34297
g31862 nor n34268 n34297 ; n34298
g31863 nor po1038 n34298 ; n34299
g31864 and pi0199 po1038 ; n34300
g31865 or n34299 n34300 ; po0356
g31866 and pi0200 n17059_not ; n34302
g31867 nor pi0606 n34302 ; n34303
g31868 and pi0200 n2571_not ; n34304
g31869 nor pi0200 n19432 ; n34305
g31870 and n19438 n34305_not ; n34306
g31871 nor pi0200 n17275 ; n34307
g31872 and pi0200 n17221 ; n34308
g31873 nor pi0038 n34307 ; n34309
g31874 and n34308_not n34309 ; n34310
g31875 nor n34306 n34310 ; n34311
g31876 and n2571 n34311_not ; n34312
g31877 and pi0606 n34304_not ; n34313
g31878 and n34312_not n34313 ; n34314
g31879 nor n34303 n34314 ; n34315
g31880 nor n17117 n34315 ; n34316
g31881 and n17117 n34302_not ; n34317
g31882 nor n34316 n34317 ; n34318
g31883 and pi0785_not n34318 ; n34319
g31884 nor pi0609 n34302 ; n34320
g31885 and pi0609 n34318_not ; n34321
g31886 and pi1155 n34320_not ; n34322
g31887 and n34321_not n34322 ; n34323
g31888 nor pi0609 n34318 ; n34324
g31889 and pi0609 n34302_not ; n34325
g31890 nor pi1155 n34325 ; n34326
g31891 and n34324_not n34326 ; n34327
g31892 nor n34323 n34327 ; n34328
g31893 and pi0785 n34328_not ; n34329
g31894 nor n34319 n34329 ; n34330
g31895 nor pi0781 n34330 ; n34331
g31896 nor pi0618 n34302 ; n34332
g31897 and pi0618 n34330 ; n34333
g31898 and pi1154 n34332_not ; n34334
g31899 and n34333_not n34334 ; n34335
g31900 and pi0618 n34302_not ; n34336
g31901 and pi0618_not n34330 ; n34337
g31902 nor pi1154 n34336 ; n34338
g31903 and n34337_not n34338 ; n34339
g31904 nor n34335 n34339 ; n34340
g31905 and pi0781 n34340_not ; n34341
g31906 nor n34331 n34341 ; n34342
g31907 nor pi0789 n34342 ; n34343
g31908 nor pi0619 n34302 ; n34344
g31909 and pi0619 n34342 ; n34345
g31910 and pi1159 n34344_not ; n34346
g31911 and n34345_not n34346 ; n34347
g31912 and pi0619 n34302_not ; n34348
g31913 and pi0619_not n34342 ; n34349
g31914 nor pi1159 n34348 ; n34350
g31915 and n34349_not n34350 ; n34351
g31916 nor n34347 n34351 ; n34352
g31917 and pi0789 n34352_not ; n34353
g31918 nor n34343 n34353 ; n34354
g31919 nor n17969 n34354 ; n34355
g31920 and n17969 n34302 ; n34356
g31921 nor n34355 n34356 ; n34357
g31922 nor n17779 n34357 ; n34358
g31923 and n17779 n34302 ; n34359
g31924 nor n34358 n34359 ; n34360
g31925 nor n17804 n34360 ; n34361
g31926 and n17804 n34302 ; n34362
g31927 nor n34361 n34362 ; n34363
g31928 and pi0644_not n34363 ; n34364
g31929 and pi0644 n34302_not ; n34365
g31930 and pi0715 n34365_not ; n34366
g31931 and n34364_not n34366 ; n34367
g31932 and n16635 n34302_not ; n34368
g31933 and n17075 n34302_not ; n34369
g31934 nor pi0643 n34302 ; n34370
g31935 nor pi0200 n16641 ; n34371
g31936 and n19899 n34371_not ; n34372
g31937 and pi0200_not n16733 ; n34373
g31938 and pi0200 n16823 ; n34374
g31939 nor pi0299 n34373 ; n34375
g31940 and n34374_not n34375 ; n34376
g31941 and pi0200_not n16747 ; n34377
g31942 and pi0200 n16838 ; n34378
g31943 and pi0299 n34377_not ; n34379
g31944 and n34378_not n34379 ; n34380
g31945 nor n34376 n34380 ; n34381
g31946 and pi0039 n34381_not ; n34382
g31947 nor pi0200 n16926 ; n34383
g31948 and pi0200 n16948 ; n34384
g31949 nor pi0039 n34383 ; n34385
g31950 and n34384_not n34385 ; n34386
g31951 nor n34382 n34386 ; n34387
g31952 nor pi0038 n34387 ; n34388
g31953 nor n34372 n34388 ; n34389
g31954 and n2571 n34389_not ; n34390
g31955 and pi0643 n34304_not ; n34391
g31956 and n34390_not n34391 ; n34392
g31957 nor n34370 n34392 ; n34393
g31958 and pi0778_not n34393 ; n34394
g31959 nor pi0625 n34302 ; n34395
g31960 and pi0625 n34393_not ; n34396
g31961 and pi1153 n34395_not ; n34397
g31962 and n34396_not n34397 ; n34398
g31963 nor pi0625 n34393 ; n34399
g31964 and pi0625 n34302_not ; n34400
g31965 nor pi1153 n34400 ; n34401
g31966 and n34399_not n34401 ; n34402
g31967 nor n34398 n34402 ; n34403
g31968 and pi0778 n34403_not ; n34404
g31969 nor n34394 n34404 ; n34405
g31970 and n17075_not n34405 ; n34406
g31971 nor n34369 n34406 ; n34407
g31972 and n16639_not n34407 ; n34408
g31973 and n16639 n34302 ; n34409
g31974 nor n34408 n34409 ; n34410
g31975 and n16635_not n34410 ; n34411
g31976 nor n34368 n34411 ; n34412
g31977 and n16631_not n34412 ; n34413
g31978 and n16631 n34302 ; n34414
g31979 nor n34413 n34414 ; n34415
g31980 nor pi0792 n34415 ; n34416
g31981 and pi0628 n34302_not ; n34417
g31982 and pi0628_not n34415 ; n34418
g31983 nor pi1156 n34417 ; n34419
g31984 and n34418_not n34419 ; n34420
g31985 nor pi0628 n34302 ; n34421
g31986 and pi0628 n34415 ; n34422
g31987 and pi1156 n34421_not ; n34423
g31988 and n34422_not n34423 ; n34424
g31989 nor n34420 n34424 ; n34425
g31990 and pi0792 n34425_not ; n34426
g31991 nor n34416 n34426 ; n34427
g31992 nor pi0787 n34427 ; n34428
g31993 and pi0647 n34427_not ; n34429
g31994 and pi0647_not n34302 ; n34430
g31995 nor n34429 n34430 ; n34431
g31996 and pi1157 n34431_not ; n34432
g31997 and pi0647 n34302_not ; n34433
g31998 and pi0647_not n34427 ; n34434
g31999 nor pi1157 n34433 ; n34435
g32000 and n34434_not n34435 ; n34436
g32001 nor n34432 n34436 ; n34437
g32002 and pi0787 n34437_not ; n34438
g32003 nor n34428 n34438 ; n34439
g32004 and pi0644 n34439 ; n34440
g32005 and pi0629_not n34424 ; n34441
g32006 nor n20570 n34357 ; n34442
g32007 and pi0629 n34420 ; n34443
g32008 nor n34441 n34443 ; n34444
g32009 and n34442_not n34444 ; n34445
g32010 and pi0792 n34445_not ; n34446
g32011 and pi0609 n34405 ; n34447
g32012 and pi0643_not n34315 ; n34448
g32013 nor n19491 n19492 ; n34449
g32014 nor pi0200 n34449 ; n34450
g32015 and pi0038 pi0200 ; n34451
g32016 and n19485 n34451 ; n34452
g32017 nor pi0200 n19493 ; n34453
g32018 and pi0200 n24754_not ; n34454
g32019 nor pi0038 n34453 ; n34455
g32020 and n34454_not n34455 ; n34456
g32021 and pi0606 n2571 ; n34457
g32022 and n34452_not n34457 ; n34458
g32023 and n34450_not n34458 ; n34459
g32024 and n34456_not n34459 ; n34460
g32025 nor n16647 n17355 ; n34461
g32026 and n34372 n34461_not ; n34462
g32027 nor pi0200 n19467 ; n34463
g32028 and pi0200 n19475_not ; n34464
g32029 nor pi0038 n34463 ; n34465
g32030 and n34464_not n34465 ; n34466
g32031 nor n34462 n34466 ; n34467
g32032 and pi0606_not n2571 ; n34468
g32033 and n34467_not n34468 ; n34469
g32034 nor n34304 n34460 ; n34470
g32035 and n34469_not n34470 ; n34471
g32036 and pi0643 n34471_not ; n34472
g32037 nor n34448 n34472 ; n34473
g32038 and pi0625_not n34473 ; n34474
g32039 and pi0625 n34315_not ; n34475
g32040 nor pi1153 n34475 ; n34476
g32041 and n34474_not n34476 ; n34477
g32042 nor pi0608 n34398 ; n34478
g32043 and n34477_not n34478 ; n34479
g32044 and pi0625 n34473 ; n34480
g32045 nor pi0625 n34315 ; n34481
g32046 and pi1153 n34481_not ; n34482
g32047 and n34480_not n34482 ; n34483
g32048 and pi0608 n34402_not ; n34484
g32049 and n34483_not n34484 ; n34485
g32050 nor n34479 n34485 ; n34486
g32051 and pi0778 n34486_not ; n34487
g32052 and pi0778_not n34473 ; n34488
g32053 nor n34487 n34488 ; n34489
g32054 nor pi0609 n34489 ; n34490
g32055 nor pi1155 n34447 ; n34491
g32056 and n34490_not n34491 ; n34492
g32057 nor pi0660 n34323 ; n34493
g32058 and n34492_not n34493 ; n34494
g32059 and pi0609_not n34405 ; n34495
g32060 and pi0609 n34489_not ; n34496
g32061 and pi1155 n34495_not ; n34497
g32062 and n34496_not n34497 ; n34498
g32063 and pi0660 n34327_not ; n34499
g32064 and n34498_not n34499 ; n34500
g32065 nor n34494 n34500 ; n34501
g32066 and pi0785 n34501_not ; n34502
g32067 nor pi0785 n34489 ; n34503
g32068 nor n34502 n34503 ; n34504
g32069 nor pi0618 n34504 ; n34505
g32070 and pi0618 n34407_not ; n34506
g32071 nor pi1154 n34506 ; n34507
g32072 and n34505_not n34507 ; n34508
g32073 nor pi0627 n34335 ; n34509
g32074 and n34508_not n34509 ; n34510
g32075 and pi0618 n34504_not ; n34511
g32076 nor pi0618 n34407 ; n34512
g32077 and pi1154 n34512_not ; n34513
g32078 and n34511_not n34513 ; n34514
g32079 and pi0627 n34339_not ; n34515
g32080 and n34514_not n34515 ; n34516
g32081 nor n34510 n34516 ; n34517
g32082 and pi0781 n34517_not ; n34518
g32083 nor pi0781 n34504 ; n34519
g32084 nor n34518 n34519 ; n34520
g32085 and pi0789_not n34520 ; n34521
g32086 nor pi0619 n34520 ; n34522
g32087 and pi0619 n34410 ; n34523
g32088 nor pi1159 n34523 ; n34524
g32089 and n34522_not n34524 ; n34525
g32090 nor pi0648 n34347 ; n34526
g32091 and n34525_not n34526 ; n34527
g32092 and pi0619 n34520_not ; n34528
g32093 and pi0619_not n34410 ; n34529
g32094 and pi1159 n34529_not ; n34530
g32095 and n34528_not n34530 ; n34531
g32096 and pi0648 n34351_not ; n34532
g32097 and n34531_not n34532 ; n34533
g32098 and pi0789 n34527_not ; n34534
g32099 and n34533_not n34534 ; n34535
g32100 and n17970 n34521_not ; n34536
g32101 and n34535_not n34536 ; n34537
g32102 and n17871 n34412_not ; n34538
g32103 and pi0626 n34302 ; n34539
g32104 nor pi0626 n34354 ; n34540
g32105 and n16629 n34539_not ; n34541
g32106 and n34540_not n34541 ; n34542
g32107 and pi0626_not n34302 ; n34543
g32108 and pi0626 n34354_not ; n34544
g32109 and n16628 n34543_not ; n34545
g32110 and n34544_not n34545 ; n34546
g32111 nor n34538 n34542 ; n34547
g32112 and n34546_not n34547 ; n34548
g32113 and pi0788 n34548_not ; n34549
g32114 nor n20364 n34549 ; n34550
g32115 and n34537_not n34550 ; n34551
g32116 nor n34446 n34551 ; n34552
g32117 nor n20206 n34552 ; n34553
g32118 and pi0630 n34436 ; n34554
g32119 nor n20559 n34360 ; n34555
g32120 and n17801 n34431_not ; n34556
g32121 nor n34554 n34555 ; n34557
g32122 and n34556_not n34557 ; n34558
g32123 and pi0787 n34558_not ; n34559
g32124 nor n34553 n34559 ; n34560
g32125 and pi0644_not n34560 ; n34561
g32126 nor pi0715 n34440 ; n34562
g32127 and n34561_not n34562 ; n34563
g32128 nor pi1160 n34367 ; n34564
g32129 and n34563_not n34564 ; n34565
g32130 and pi0644_not n34439 ; n34566
g32131 and pi0644 n34560 ; n34567
g32132 and pi0715 n34566_not ; n34568
g32133 and n34567_not n34568 ; n34569
g32134 and pi0644 n34363 ; n34570
g32135 nor pi0644 n34302 ; n34571
g32136 nor pi0715 n34571 ; n34572
g32137 and n34570_not n34572 ; n34573
g32138 and pi1160 n34573_not ; n34574
g32139 and n34569_not n34574 ; n34575
g32140 nor n34565 n34575 ; n34576
g32141 and pi0790 n34576_not ; n34577
g32142 and pi0790_not n34560 ; n34578
g32143 nor n34577 n34578 ; n34579
g32144 nor po1038 n34579 ; n34580
g32145 and pi0200_not po1038 ; n34581
g32146 nor n34580 n34581 ; po0357
g32147 and pi0233 pi0237 ; n34583
g32148 and pi0057 pi0332 ; n34584
g32149 and n2572 n6573 ; n34585
g32150 and n2521 n34585 ; n34586
g32151 nor pi0332 n34586 ; n34587
g32152 and n6304 n34587_not ; n34588
g32153 and pi0332 n6304_not ; n34589
g32154 and pi0059 n34589_not ; n34590
g32155 and n34588_not n34590 ; n34591
g32156 and pi0332 n2529_not ; n34592
g32157 nor pi0059 n34592 ; n34593
g32158 and pi0055 n34587 ; n34594
g32159 and pi0074 pi0332 ; n34595
g32160 nor pi0055 n34595 ; n34596
g32161 and n2726 n11086 ; n34597
g32162 and pi0468 n6192 ; n34598
g32163 and pi0299_not pi0587 ; n34599
g32164 nor n21044 n34599 ; n34600
g32165 nor pi0468 n34600 ; n34601
g32166 nor n34598 n34601 ; n34602
g32167 and n34597 n34602_not ; n34603
g32168 nor pi0332 n34603 ; n34604
g32169 and n7363 n34604_not ; n34605
g32170 and n2521 n6585 ; n34606
g32171 nor pi0332 n34606 ; n34607
g32172 and n15625 n34607_not ; n34608
g32173 and pi0332 n2611_not ; n34609
g32174 nor n34608 n34609 ; n34610
g32175 and n34605_not n34610 ; n34611
g32176 nor pi0074 n34611 ; n34612
g32177 and n34596 n34612_not ; n34613
g32178 and n2529 n34594_not ; n34614
g32179 and n34613_not n34614 ; n34615
g32180 and n34593 n34615_not ; n34616
g32181 nor pi0057 n34591 ; n34617
g32182 and n34616_not n34617 ; n34618
g32183 nor n34584 n34618 ; n34619
g32184 nor n34583 n34619 ; n34620
g32185 nor pi0332 n6192 ; n34621
g32186 nor pi0947 n34621 ; n34622
g32187 and pi0096 pi0210 ; n34623
g32188 and pi0332 n34623 ; n34624
g32189 and pi0032_not pi0070 ; n34625
g32190 nor pi0070 pi0841 ; n34626
g32191 and pi0032 n34626 ; n34627
g32192 nor n34625 n34627 ; n34628
g32193 nor pi0210 n34628 ; n34629
g32194 nor pi0032 pi0096 ; n34630
g32195 and pi0070 n34630 ; n34631
g32196 nor pi0332 n34631 ; n34632
g32197 and n34629_not n34632 ; n34633
g32198 nor n34624 n34633 ; n34634
g32199 and n6197_not n34634 ; n34635
g32200 and n6192 n34635_not ; n34636
g32201 and n34622 n34636_not ; n34637
g32202 and n6192 n34634_not ; n34638
g32203 and pi0332 pi0468 ; n34639
g32204 nor pi0468 n34633 ; n34640
g32205 nor n34639 n34640 ; n34641
g32206 and n6192_not n34641 ; n34642
g32207 and pi0947 n34638_not ; n34643
g32208 and n34642_not n34643 ; n34644
g32209 nor n34637 n34644 ; n34645
g32210 and pi0057 n34645_not ; n34646
g32211 and n6304_not n34645 ; n34647
g32212 and n2572_not n34645 ; n34648
g32213 and pi0032 n34626_not ; n34649
g32214 and pi0095_not n2736 ; n34650
g32215 and n34649_not n34650 ; n34651
g32216 and n2706 n34651 ; n34652
g32217 and n2728 n34652 ; n34653
g32218 and n34628 n34653_not ; n34654
g32219 nor pi0210 n34654 ; n34655
g32220 and pi0095_not n2975 ; n34656
g32221 nor pi0070 n34656 ; n34657
g32222 and n34630 n34657_not ; n34658
g32223 and pi0210 n34658 ; n34659
g32224 nor pi0332 n34655 ; n34660
g32225 and n34659_not n34660 ; n34661
g32226 nor n34624 n34661 ; n34662
g32227 and n6197_not n34662 ; n34663
g32228 and n6192 n34663_not ; n34664
g32229 and n34622 n34664_not ; n34665
g32230 and n6192 n34662_not ; n34666
g32231 nor pi0468 n34661 ; n34667
g32232 nor n34639 n34667 ; n34668
g32233 and n6192_not n34668 ; n34669
g32234 and pi0947 n34666_not ; n34670
g32235 and n34669_not n34670 ; n34671
g32236 nor n34665 n34671 ; n34672
g32237 and n2572 n34672 ; n34673
g32238 nor n34648 n34673 ; n34674
g32239 and n6304 n34674_not ; n34675
g32240 and pi0059 n34647_not ; n34676
g32241 and n34675_not n34676 ; n34677
g32242 and n2529_not n34645 ; n34678
g32243 and pi0055 n34674 ; n34679
g32244 and pi0074_not n2611 ; n34680
g32245 and pi0299 n34645_not ; n34681
g32246 and pi0096 pi0198 ; n34682
g32247 and pi0332 n34682 ; n34683
g32248 nor pi0198 n34628 ; n34684
g32249 and n34632 n34684_not ; n34685
g32250 nor n34683 n34685 ; n34686
g32251 and n6192 n34686_not ; n34687
g32252 and n6583 n34685_not ; n34688
g32253 and n34621 n34688_not ; n34689
g32254 nor pi0299 n6582 ; n34690
g32255 and n34687_not n34690 ; n34691
g32256 and n34689_not n34691 ; n34692
g32257 nor n34680 n34692 ; n34693
g32258 and n34681_not n34693 ; n34694
g32259 and n2726 n2962 ; n34695
g32260 and n34651 n34695 ; n34696
g32261 and n34628 n34696_not ; n34697
g32262 nor pi0210 n34697 ; n34698
g32263 and pi0095_not n2517 ; n34699
g32264 and n34695 n34699 ; n34700
g32265 nor pi0070 n34700 ; n34701
g32266 and n34630 n34701_not ; n34702
g32267 and pi0210 n34702 ; n34703
g32268 nor pi0332 n34698 ; n34704
g32269 and n34703_not n34704 ; n34705
g32270 nor n34624 n34705 ; n34706
g32271 and n6197_not n34706 ; n34707
g32272 and n6192 n34707_not ; n34708
g32273 and n34622 n34708_not ; n34709
g32274 and n6192 n34706_not ; n34710
g32275 nor pi0468 n34705 ; n34711
g32276 nor n34639 n34711 ; n34712
g32277 and n6192_not n34712 ; n34713
g32278 and pi0947 n34710_not ; n34714
g32279 and n34713_not n34714 ; n34715
g32280 and pi0299 n34709_not ; n34716
g32281 and n34715_not n34716 ; n34717
g32282 nor pi0587 n34621 ; n34718
g32283 nor pi0198 n34697 ; n34719
g32284 and pi0198 n34702 ; n34720
g32285 nor pi0332 n34719 ; n34721
g32286 and n34720_not n34721 ; n34722
g32287 nor n34683 n34722 ; n34723
g32288 and n6197_not n34723 ; n34724
g32289 and n6192 n34724_not ; n34725
g32290 and n34718 n34725_not ; n34726
g32291 and n6192 n34723_not ; n34727
g32292 nor pi0468 n34722 ; n34728
g32293 nor n6192 n34639 ; n34729
g32294 and n34728_not n34729 ; n34730
g32295 and pi0587 n34727_not ; n34731
g32296 and n34730_not n34731 ; n34732
g32297 nor pi0299 n34726 ; n34733
g32298 and n34732_not n34733 ; n34734
g32299 nor n34717 n34734 ; n34735
g32300 and n7363 n34735_not ; n34736
g32301 and pi0299 n34672_not ; n34737
g32302 nor pi0198 n34654 ; n34738
g32303 and pi0198 n34658 ; n34739
g32304 nor pi0332 n34738 ; n34740
g32305 and n34739_not n34740 ; n34741
g32306 nor n34683 n34741 ; n34742
g32307 and n6197_not n34742 ; n34743
g32308 and n6192 n34743_not ; n34744
g32309 and n34718 n34744_not ; n34745
g32310 and n6192 n34742_not ; n34746
g32311 nor pi0468 n34741 ; n34747
g32312 and n34729 n34747_not ; n34748
g32313 and pi0587 n34746_not ; n34749
g32314 and n34748_not n34749 ; n34750
g32315 nor n34745 n34750 ; n34751
g32316 nor pi0299 n34751 ; n34752
g32317 and n15625 n34737_not ; n34753
g32318 and n34752_not n34753 ; n34754
g32319 nor n34736 n34754 ; n34755
g32320 nor pi0074 n34755 ; n34756
g32321 nor pi0055 n34694 ; n34757
g32322 and n34756_not n34757 ; n34758
g32323 and n2529 n34679_not ; n34759
g32324 and n34758_not n34759 ; n34760
g32325 nor pi0059 n34678 ; n34761
g32326 and n34760_not n34761 ; n34762
g32327 nor n34677 n34762 ; n34763
g32328 nor pi0057 n34763 ; n34764
g32329 nor n34646 n34764 ; n34765
g32330 and n34583 n34765_not ; n34766
g32331 nor n34620 n34766 ; n34767
g32332 nor pi0201 n34767 ; n34768
g32333 nor n6573 n16479 ; n34769
g32334 and n6583 n34682 ; n34770
g32335 and n16479 n34770_not ; n34771
g32336 nor n16479 n34623 ; n34772
g32337 nor n34769 n34771 ; n34773
g32338 and n34772_not n34773 ; n34774
g32339 and n34583 n34774 ; n34775
g32340 and pi0201 n34775_not ; n34776
g32341 nor n34768 n34776 ; po0358
g32342 and pi0233_not pi0237 ; n34778
g32343 nor n34619 n34778 ; n34779
g32344 and n34765_not n34778 ; n34780
g32345 nor n34779 n34780 ; n34781
g32346 nor pi0202 n34781 ; n34782
g32347 and n34774 n34778 ; n34783
g32348 and pi0202 n34783_not ; n34784
g32349 nor n34782 n34784 ; po0359
g32350 nor pi0233 pi0237 ; n34786
g32351 nor n34619 n34786 ; n34787
g32352 and n34765_not n34786 ; n34788
g32353 nor n34787 n34788 ; n34789
g32354 nor pi0203 n34789 ; n34790
g32355 and n34774 n34786 ; n34791
g32356 and pi0203 n34791_not ; n34792
g32357 nor n34790 n34792 ; po0360
g32358 and n2572 n6310 ; n34794
g32359 and n2521 n34794 ; n34795
g32360 nor pi0332 n34795 ; n34796
g32361 and n6304 n34796_not ; n34797
g32362 and n34590 n34797_not ; n34798
g32363 and pi0055 n34796 ; n34799
g32364 and pi0468_not pi0602 ; n34800
g32365 and pi0468 n6195 ; n34801
g32366 nor n34800 n34801 ; n34802
g32367 nor pi0299 n34802 ; n34803
g32368 nor n6324 n34803 ; n34804
g32369 and n2521 n34804_not ; n34805
g32370 nor pi0332 n34805 ; n34806
g32371 and n15625 n34806_not ; n34807
g32372 nor pi0299 pi0602 ; n34808
g32373 and pi0299 pi0907_not ; n34809
g32374 nor pi0468 n34808 ; n34810
g32375 and n34809_not n34810 ; n34811
g32376 nor n34801 n34811 ; n34812
g32377 and n34597 n34812_not ; n34813
g32378 nor pi0332 n34813 ; n34814
g32379 and n7363 n34814_not ; n34815
g32380 nor n34807 n34815 ; n34816
g32381 nor pi0074 n34816 ; n34817
g32382 and n34596 n34609_not ; n34818
g32383 and n34817_not n34818 ; n34819
g32384 and n2529 n34799_not ; n34820
g32385 and n34819_not n34820 ; n34821
g32386 and n34593 n34821_not ; n34822
g32387 nor pi0057 n34798 ; n34823
g32388 and n34822_not n34823 ; n34824
g32389 nor n34584 n34824 ; n34825
g32390 nor n34583 n34825 ; n34826
g32391 nor pi0332 n6195 ; n34827
g32392 nor pi0907 n34827 ; n34828
g32393 and n6195 n34635_not ; n34829
g32394 and n34828 n34829_not ; n34830
g32395 and n6195 n34634_not ; n34831
g32396 and n6195_not n34641 ; n34832
g32397 and pi0907 n34831_not ; n34833
g32398 and n34832_not n34833 ; n34834
g32399 nor n34830 n34834 ; n34835
g32400 and pi0057 n34835_not ; n34836
g32401 and n6304_not n34835 ; n34837
g32402 and n2572_not n34835 ; n34838
g32403 and n6195 n34662_not ; n34839
g32404 and n6195_not n34668 ; n34840
g32405 and pi0907 n34839_not ; n34841
g32406 and n34840_not n34841 ; n34842
g32407 and pi0332 n16657_not ; n34843
g32408 and pi0680 n34843_not ; n34844
g32409 and n34663_not n34844 ; n34845
g32410 and n34828 n34845_not ; n34846
g32411 nor n34842 n34846 ; n34847
g32412 and n2572 n34847 ; n34848
g32413 nor n34838 n34848 ; n34849
g32414 and n6304 n34849_not ; n34850
g32415 and pi0059 n34837_not ; n34851
g32416 and n34850_not n34851 ; n34852
g32417 and n2529_not n34835 ; n34853
g32418 and pi0055 n34849 ; n34854
g32419 and pi0299 n34847 ; n34855
g32420 and n6195 n34682 ; n34856
g32421 and pi0332 n34856_not ; n34857
g32422 nor pi0299 n34857 ; n34858
g32423 and n6326 n34742 ; n34859
g32424 and n34858 n34859_not ; n34860
g32425 nor n34855 n34860 ; n34861
g32426 and n15625 n34861_not ; n34862
g32427 and n6326 n34723 ; n34863
g32428 and n34858 n34863_not ; n34864
g32429 and n6195 n34707_not ; n34865
g32430 and n34828 n34865_not ; n34866
g32431 and n6195 n34706_not ; n34867
g32432 and n6195_not n34712 ; n34868
g32433 and pi0907 n34867_not ; n34869
g32434 and n34868_not n34869 ; n34870
g32435 and pi0299 n34866_not ; n34871
g32436 and n34870_not n34871 ; n34872
g32437 nor n34864 n34872 ; n34873
g32438 and n7363 n34873_not ; n34874
g32439 nor n34862 n34874 ; n34875
g32440 nor pi0074 n34875 ; n34876
g32441 and pi0299 n34835_not ; n34877
g32442 and n34686 n34802_not ; n34878
g32443 nor n34857 n34878 ; n34879
g32444 nor pi0299 n34879 ; n34880
g32445 nor n34680 n34880 ; n34881
g32446 and n34877_not n34881 ; n34882
g32447 nor pi0055 n34882 ; n34883
g32448 and n34876_not n34883 ; n34884
g32449 and n2529 n34854_not ; n34885
g32450 and n34884_not n34885 ; n34886
g32451 nor pi0059 n34853 ; n34887
g32452 and n34886_not n34887 ; n34888
g32453 nor n34852 n34888 ; n34889
g32454 nor pi0057 n34889 ; n34890
g32455 nor n34836 n34890 ; n34891
g32456 and n34583 n34891_not ; n34892
g32457 nor n34826 n34892 ; n34893
g32458 nor pi0204 n34893 ; n34894
g32459 nor n6310 n16479 ; n34895
g32460 and n6326 n34682 ; n34896
g32461 and n16479 n34896_not ; n34897
g32462 nor n34772 n34895 ; n34898
g32463 and n34897_not n34898 ; n34899
g32464 and n34583 n34899 ; n34900
g32465 and pi0204 n34900_not ; n34901
g32466 nor n34894 n34901 ; po0361
g32467 nor n34778 n34825 ; n34903
g32468 and n34778 n34891_not ; n34904
g32469 nor n34903 n34904 ; n34905
g32470 nor pi0205 n34905 ; n34906
g32471 and n34778 n34899 ; n34907
g32472 and pi0205 n34907_not ; n34908
g32473 nor n34906 n34908 ; po0362
g32474 and pi0233 pi0237_not ; n34910
g32475 nor n34825 n34910 ; n34911
g32476 and n34891_not n34910 ; n34912
g32477 nor n34911 n34912 ; n34913
g32478 nor pi0206 n34913 ; n34914
g32479 and n34899 n34910 ; n34915
g32480 and pi0206 n34915_not ; n34916
g32481 nor n34914 n34916 ; po0363
g32482 and n19146_not n24385 ; n34918
g32483 and n19151 n34918 ; n34919
g32484 and n19142_not n34919 ; n34920
g32485 and pi0207 n34920_not ; n34921
g32486 and n16635 n17059_not ; n34922
g32487 and n2571 n24388 ; n34923
g32488 nor pi0778 n34923 ; n34924
g32489 nor pi0625 n17059 ; n34925
g32490 and pi0625 n34923_not ; n34926
g32491 nor n34925 n34926 ; n34927
g32492 and pi1153 n34927_not ; n34928
g32493 and pi0625 n17059_not ; n34929
g32494 nor pi0625 n34923 ; n34930
g32495 nor n34929 n34930 ; n34931
g32496 nor pi1153 n34931 ; n34932
g32497 nor n34928 n34932 ; n34933
g32498 and pi0778 n34933_not ; n34934
g32499 nor n34924 n34934 ; n34935
g32500 nor n17075 n34935 ; n34936
g32501 and n17059_not n17075 ; n34937
g32502 nor n34936 n34937 ; n34938
g32503 and n16639_not n34938 ; n34939
g32504 and n16639 n17059 ; n34940
g32505 nor n34939 n34940 ; n34941
g32506 and n16635_not n34941 ; n34942
g32507 nor n34922 n34942 ; n34943
g32508 and n16631_not n34943 ; n34944
g32509 and n16631 n17059 ; n34945
g32510 nor n34944 n34945 ; n34946
g32511 nor n19142 n34946 ; n34947
g32512 and n17059 n17856 ; n34948
g32513 nor n34947 n34948 ; n34949
g32514 nor pi0207 n34949 ; n34950
g32515 nor n34921 n34950 ; n34951
g32516 and pi0710 n34951_not ; n34952
g32517 nor pi0207 n17059 ; n34953
g32518 nor pi0710 n34953 ; n34954
g32519 nor n34952 n34954 ; n34955
g32520 nor pi0787 n34955 ; n34956
g32521 and pi0647_not n34955 ; n34957
g32522 and pi0647 n34953 ; n34958
g32523 nor pi1157 n34958 ; n34959
g32524 and n34957_not n34959 ; n34960
g32525 and pi0647_not n34953 ; n34961
g32526 and pi0647 n34955 ; n34962
g32527 and pi1157 n34961_not ; n34963
g32528 and n34962_not n34963 ; n34964
g32529 nor n34960 n34964 ; n34965
g32530 and pi0787 n34965_not ; n34966
g32531 nor n34956 n34966 ; n34967
g32532 and pi0644_not n34967 ; n34968
g32533 and pi0630_not n34964 ; n34969
g32534 and n17059_not n17117 ; n34970
g32535 and n2571 n19439 ; n34971
g32536 nor n17117 n34971 ; n34972
g32537 nor n34970 n34972 ; n34973
g32538 nor pi0785 n34973 ; n34974
g32539 nor n17059 n17296 ; n34975
g32540 and pi0609_not n34972 ; n34976
g32541 nor n34975 n34976 ; n34977
g32542 nor pi1155 n34977 ; n34978
g32543 nor n17059 n17291 ; n34979
g32544 and pi0609 n34972 ; n34980
g32545 nor n34979 n34980 ; n34981
g32546 and pi1155 n34981_not ; n34982
g32547 nor n34978 n34982 ; n34983
g32548 and pi0785 n34983_not ; n34984
g32549 nor n34974 n34984 ; n34985
g32550 nor pi0781 n34985 ; n34986
g32551 and pi0618_not n34985 ; n34987
g32552 and pi0618 n17059 ; n34988
g32553 nor pi1154 n34988 ; n34989
g32554 and n34987_not n34989 ; n34990
g32555 and pi0618_not n17059 ; n34991
g32556 and pi0618 n34985 ; n34992
g32557 and pi1154 n34991_not ; n34993
g32558 and n34992_not n34993 ; n34994
g32559 nor n34990 n34994 ; n34995
g32560 and pi0781 n34995_not ; n34996
g32561 nor n34986 n34996 ; n34997
g32562 nor pi0789 n34997 ; n34998
g32563 and pi0619_not n34997 ; n34999
g32564 and pi0619 n17059 ; n35000
g32565 nor pi1159 n35000 ; n35001
g32566 and n34999_not n35001 ; n35002
g32567 and pi0619_not n17059 ; n35003
g32568 and pi0619 n34997 ; n35004
g32569 and pi1159 n35003_not ; n35005
g32570 and n35004_not n35005 ; n35006
g32571 nor n35002 n35006 ; n35007
g32572 and pi0789 n35007_not ; n35008
g32573 nor n34998 n35008 ; n35009
g32574 and n17969_not n35009 ; n35010
g32575 and n17059 n17969 ; n35011
g32576 nor n35010 n35011 ; n35012
g32577 nor n17779 n35012 ; n35013
g32578 and n17059 n17779 ; n35014
g32579 nor n35013 n35014 ; n35015
g32580 nor pi0207 n35015 ; n35016
g32581 and n2571 n24447_not ; n35017
g32582 and n17117_not n35017 ; n35018
g32583 and n20225_not n35018 ; n35019
g32584 and n20235_not n35019 ; n35020
g32585 and n20231_not n35020 ; n35021
g32586 and n17969_not n35021 ; n35022
g32587 and n17779_not n35022 ; n35023
g32588 and pi0207 n35023_not ; n35024
g32589 and pi0623 n35024_not ; n35025
g32590 and n35016_not n35025 ; n35026
g32591 and pi0623_not n34953 ; n35027
g32592 nor n35026 n35027 ; n35028
g32593 and n20559_not n35028 ; n35029
g32594 and pi0630 n34960 ; n35030
g32595 nor n34969 n35029 ; n35031
g32596 and n35030_not n35031 ; n35032
g32597 and pi0787 n35032_not ; n35033
g32598 nor pi0710 n35028 ; n35034
g32599 nor pi0628 n17059 ; n35035
g32600 and pi0628 n34946 ; n35036
g32601 nor n35035 n35036 ; n35037
g32602 nor pi0629 n35037 ; n35038
g32603 nor n35035 n35038 ; n35039
g32604 and pi1156 n35039_not ; n35040
g32605 and pi0628 n17059_not ; n35041
g32606 and pi1156_not n35041 ; n35042
g32607 and pi0628_not n34946 ; n35043
g32608 nor n35041 n35043 ; n35044
g32609 and n17777 n35044_not ; n35045
g32610 nor n35042 n35045 ; n35046
g32611 and n35040_not n35046 ; n35047
g32612 and pi0792 n35047_not ; n35048
g32613 and pi1159 n17059_not ; n35049
g32614 and pi0619 n34941 ; n35050
g32615 and pi1154 n17059_not ; n35051
g32616 and pi0618 n34938_not ; n35052
g32617 and pi1155 n17059_not ; n35053
g32618 and pi0609 n34935_not ; n35054
g32619 and n2571 n19477_not ; n35055
g32620 nor pi0778 n35055 ; n35056
g32621 nor pi0625 n35055 ; n35057
g32622 nor n34929 n35057 ; n35058
g32623 nor pi1153 n35058 ; n35059
g32624 nor pi0608 n34928 ; n35060
g32625 and n35059_not n35060 ; n35061
g32626 and pi0625 n35055_not ; n35062
g32627 nor n34925 n35062 ; n35063
g32628 and pi1153 n35063_not ; n35064
g32629 and pi0608 n34932_not ; n35065
g32630 and n35064_not n35065 ; n35066
g32631 and pi0778 n35061_not ; n35067
g32632 and n35066_not n35067 ; n35068
g32633 nor n35056 n35068 ; n35069
g32634 nor pi0609 n35069 ; n35070
g32635 nor n35054 n35070 ; n35071
g32636 nor pi1155 n35071 ; n35072
g32637 nor pi0660 n35053 ; n35073
g32638 and n35072_not n35073 ; n35074
g32639 nor pi1155 n17059 ; n35075
g32640 nor pi0609 n34935 ; n35076
g32641 and pi0609 n35069_not ; n35077
g32642 nor n35076 n35077 ; n35078
g32643 and pi1155 n35078_not ; n35079
g32644 and pi0660 n35075_not ; n35080
g32645 and n35079_not n35080 ; n35081
g32646 nor n35074 n35081 ; n35082
g32647 and pi0785 n35082_not ; n35083
g32648 and pi0785_not n35069 ; n35084
g32649 nor n35083 n35084 ; n35085
g32650 and pi0618_not n35085 ; n35086
g32651 nor n35052 n35086 ; n35087
g32652 nor pi1154 n35087 ; n35088
g32653 nor pi0627 n35051 ; n35089
g32654 and n35088_not n35089 ; n35090
g32655 nor pi1154 n17059 ; n35091
g32656 nor pi0618 n34938 ; n35092
g32657 and pi0618 n35085 ; n35093
g32658 nor n35092 n35093 ; n35094
g32659 and pi1154 n35094_not ; n35095
g32660 and pi0627 n35091_not ; n35096
g32661 and n35095_not n35096 ; n35097
g32662 nor n35090 n35097 ; n35098
g32663 and pi0781 n35098_not ; n35099
g32664 nor pi0781 n35085 ; n35100
g32665 nor n35099 n35100 ; n35101
g32666 and pi0619_not n35101 ; n35102
g32667 nor n35050 n35102 ; n35103
g32668 nor pi1159 n35103 ; n35104
g32669 nor pi0648 n35049 ; n35105
g32670 and n35104_not n35105 ; n35106
g32671 nor pi1159 n17059 ; n35107
g32672 and pi0619_not n34941 ; n35108
g32673 and pi0619 n35101 ; n35109
g32674 nor n35108 n35109 ; n35110
g32675 and pi1159 n35110_not ; n35111
g32676 and pi0648 n35107_not ; n35112
g32677 and n35111_not n35112 ; n35113
g32678 nor n35106 n35113 ; n35114
g32679 and pi0789 n35114_not ; n35115
g32680 nor pi0789 n35101 ; n35116
g32681 nor n35115 n35116 ; n35117
g32682 nor pi0788 n35117 ; n35118
g32683 and pi0641 n17059_not ; n35119
g32684 and pi0626 n34943 ; n35120
g32685 nor pi0626 n35117 ; n35121
g32686 nor pi0641 n35120 ; n35122
g32687 and n35121_not n35122 ; n35123
g32688 nor pi1158 n35119 ; n35124
g32689 and n35123_not n35124 ; n35125
g32690 nor pi0641 n17059 ; n35126
g32691 and pi0626_not n34943 ; n35127
g32692 and pi0626 n35117_not ; n35128
g32693 and pi0641 n35127_not ; n35129
g32694 and n35128_not n35129 ; n35130
g32695 and pi1158 n35126_not ; n35131
g32696 and n35130_not n35131 ; n35132
g32697 nor n35125 n35132 ; n35133
g32698 and pi0788 n35133_not ; n35134
g32699 nor n20364 n35118 ; n35135
g32700 and n35134_not n35135 ; n35136
g32701 nor n35048 n35136 ; n35137
g32702 nor pi0207 n35137 ; n35138
g32703 and pi0609 n34918_not ; n35139
g32704 nor pi0778 n34080 ; n35140
g32705 and pi0625_not n34080 ; n35141
g32706 nor pi1153 n35141 ; n35142
g32707 and pi0625 n24385 ; n35143
g32708 and pi1153 n35143_not ; n35144
g32709 nor pi0608 n35144 ; n35145
g32710 and n35142_not n35145 ; n35146
g32711 and pi0625 n34080 ; n35147
g32712 and pi1153 n35147_not ; n35148
g32713 and pi0625_not n24385 ; n35149
g32714 nor pi1153 n35149 ; n35150
g32715 and pi0608 n35150_not ; n35151
g32716 and n35148_not n35151 ; n35152
g32717 and pi0778 n35146_not ; n35153
g32718 and n35152_not n35153 ; n35154
g32719 nor n35140 n35154 ; n35155
g32720 nor pi0609 n35155 ; n35156
g32721 and n17073 n35139_not ; n35157
g32722 and n35156_not n35157 ; n35158
g32723 and pi0609 n35155_not ; n35159
g32724 nor pi0609 n34918 ; n35160
g32725 and n17072 n35160_not ; n35161
g32726 and n35159_not n35161 ; n35162
g32727 nor n35158 n35162 ; n35163
g32728 and pi0785 n35163_not ; n35164
g32729 and pi0785_not n35155 ; n35165
g32730 nor n35164 n35165 ; n35166
g32731 and pi0781_not n35166 ; n35167
g32732 and pi0618_not n35166 ; n35168
g32733 and n17075_not n34918 ; n35169
g32734 and pi0618 n35169_not ; n35170
g32735 and n16637 n35170_not ; n35171
g32736 and n35168_not n35171 ; n35172
g32737 nor pi0618 n35169 ; n35173
g32738 and pi0618 n35166 ; n35174
g32739 and n16636 n35173_not ; n35175
g32740 and n35174_not n35175 ; n35176
g32741 and pi0781 n35172_not ; n35177
g32742 and n35176_not n35177 ; n35178
g32743 nor n23615 n35167 ; n35179
g32744 and n35178_not n35179 ; n35180
g32745 and n19150 n34918 ; n35181
g32746 and n16634 n20231 ; n35182
g32747 and n35181 n35182 ; n35183
g32748 nor n35180 n35183 ; n35184
g32749 and pi0788_not n35184 ; n35185
g32750 and n16635_not n35181 ; n35186
g32751 and pi0626 n35186_not ; n35187
g32752 nor pi0641 n35187 ; n35188
g32753 and pi0626_not n35184 ; n35189
g32754 and pi1158_not n35188 ; n35190
g32755 and n35189_not n35190 ; n35191
g32756 and pi0626 n35184 ; n35192
g32757 nor pi0626 n35186 ; n35193
g32758 and pi0641 n35193_not ; n35194
g32759 and pi1158 n35194 ; n35195
g32760 and n35192_not n35195 ; n35196
g32761 and pi0788 n35191_not ; n35197
g32762 and n35196_not n35197 ; n35198
g32763 nor n20364 n35185 ; n35199
g32764 and n35198_not n35199 ; n35200
g32765 and n17779 n17855 ; n35201
g32766 and n34919 n35201 ; n35202
g32767 nor n35200 n35202 ; n35203
g32768 and pi0207 n35203_not ; n35204
g32769 nor pi0623 n35204 ; n35205
g32770 and n35138_not n35205 ; n35206
g32771 nor pi1156 n34919 ; n35207
g32772 and pi1156 n35022_not ; n35208
g32773 and n20566 n35207_not ; n35209
g32774 and n35208_not n35209 ; n35210
g32775 and pi1156 n34919_not ; n35211
g32776 nor pi1156 n35022 ; n35212
g32777 and n20568 n35211_not ; n35213
g32778 and n35212_not n35213 ; n35214
g32779 nor n35210 n35214 ; n35215
g32780 and pi0792 n35215_not ; n35216
g32781 and n17868 n35021 ; n35217
g32782 nor pi1159 n35020 ; n35218
g32783 and pi1159 n35181_not ; n35219
g32784 and pi0619_not pi0648 ; n35220
g32785 and n35218_not n35220 ; n35221
g32786 and n35219_not n35221 ; n35222
g32787 and pi1159 n35020_not ; n35223
g32788 nor pi1159 n35181 ; n35224
g32789 and pi0619 pi0648_not ; n35225
g32790 and n35223_not n35225 ; n35226
g32791 and n35224_not n35226 ; n35227
g32792 and pi0789 n35222_not ; n35228
g32793 and n35227_not n35228 ; n35229
g32794 and pi0789 n35229_not ; n35230
g32795 nor pi1154 n35170 ; n35231
g32796 and n20233 n35019 ; n35232
g32797 nor pi0627 n35232 ; n35233
g32798 and n35231_not n35233 ; n35234
g32799 and n20232 n35019 ; n35235
g32800 nor pi0778 n34085 ; n35236
g32801 and pi0625_not n34085 ; n35237
g32802 and pi0625 n35017 ; n35238
g32803 nor pi1153 n35238 ; n35239
g32804 and n35237_not n35239 ; n35240
g32805 and n35145 n35240_not ; n35241
g32806 and pi0625_not n35017 ; n35242
g32807 and pi0625 n34085 ; n35243
g32808 and pi1153 n35242_not ; n35244
g32809 and n35243_not n35244 ; n35245
g32810 and n35151 n35245_not ; n35246
g32811 and pi0778 n35241_not ; n35247
g32812 and n35246_not n35247 ; n35248
g32813 nor n35236 n35248 ; n35249
g32814 nor pi0785 n35249 ; n35250
g32815 and n20223 n35018 ; n35251
g32816 nor pi0609 n35249 ; n35252
g32817 nor pi1155 n35139 ; n35253
g32818 and n35252_not n35253 ; n35254
g32819 nor pi0660 n35251 ; n35255
g32820 and n35254_not n35255 ; n35256
g32821 and n20222 n35018 ; n35257
g32822 and pi0609 n35249_not ; n35258
g32823 and pi1155 n35160_not ; n35259
g32824 and n35258_not n35259 ; n35260
g32825 and pi0660 n35257_not ; n35261
g32826 and n35260_not n35261 ; n35262
g32827 nor n35256 n35262 ; n35263
g32828 and pi0785 n35263_not ; n35264
g32829 nor n35250 n35264 ; n35265
g32830 and pi0618 n35265_not ; n35266
g32831 and pi1154 n35173_not ; n35267
g32832 and n35266_not n35267 ; n35268
g32833 and pi0627 n35235_not ; n35269
g32834 and n35268_not n35269 ; n35270
g32835 nor n35234 n35270 ; n35271
g32836 and pi0781 n35271_not ; n35272
g32837 nor pi0618 pi0627 ; n35273
g32838 and pi0781 n35273_not ; n35274
g32839 nor n35265 n35274 ; n35275
g32840 and n23614_not n35229 ; n35276
g32841 nor n35275 n35276 ; n35277
g32842 and n35272_not n35277 ; n35278
g32843 nor n35230 n35278 ; n35279
g32844 and pi0626_not n35279 ; n35280
g32845 and n35188 n35280_not ; n35281
g32846 nor pi1158 n35217 ; n35282
g32847 and n35281_not n35282 ; n35283
g32848 and n17869 n35021 ; n35284
g32849 and pi0626 n35279 ; n35285
g32850 and n35194 n35285_not ; n35286
g32851 and pi1158 n35284_not ; n35287
g32852 and n35286_not n35287 ; n35288
g32853 nor n35283 n35288 ; n35289
g32854 and pi0788 n35289_not ; n35290
g32855 and pi0788_not n35279 ; n35291
g32856 nor n20364 n35291 ; n35292
g32857 and n35290_not n35292 ; n35293
g32858 nor n35216 n35293 ; n35294
g32859 and pi0207 n35294_not ; n35295
g32860 and n2571 n19488 ; n35296
g32861 nor pi0778 n35296 ; n35297
g32862 and pi0625_not n34971 ; n35298
g32863 and pi0625 n35296 ; n35299
g32864 and pi1153 n35299_not ; n35300
g32865 and n35298_not n35300 ; n35301
g32866 and n35065 n35301_not ; n35302
g32867 and pi0625_not n35296 ; n35303
g32868 and pi0625 n34971 ; n35304
g32869 nor pi1153 n35303 ; n35305
g32870 and n35304_not n35305 ; n35306
g32871 and n35060 n35306_not ; n35307
g32872 and pi0778 n35302_not ; n35308
g32873 and n35307_not n35308 ; n35309
g32874 nor n35297 n35309 ; n35310
g32875 nor pi0609 n35310 ; n35311
g32876 nor n35054 n35311 ; n35312
g32877 nor pi1155 n35312 ; n35313
g32878 nor pi0660 n34982 ; n35314
g32879 and n35313_not n35314 ; n35315
g32880 and pi0609 n35310_not ; n35316
g32881 nor n35076 n35316 ; n35317
g32882 and pi1155 n35317_not ; n35318
g32883 and pi0660 n34978_not ; n35319
g32884 and n35318_not n35319 ; n35320
g32885 nor n35315 n35320 ; n35321
g32886 and pi0785 n35321_not ; n35322
g32887 and pi0785_not n35310 ; n35323
g32888 nor n35322 n35323 ; n35324
g32889 and pi0618_not n35324 ; n35325
g32890 nor n35052 n35325 ; n35326
g32891 nor pi1154 n35326 ; n35327
g32892 nor pi0627 n34994 ; n35328
g32893 and n35327_not n35328 ; n35329
g32894 and pi0618 n35324 ; n35330
g32895 nor n35092 n35330 ; n35331
g32896 and pi1154 n35331_not ; n35332
g32897 and pi0627 n34990_not ; n35333
g32898 and n35332_not n35333 ; n35334
g32899 nor n35329 n35334 ; n35335
g32900 and pi0781 n35335_not ; n35336
g32901 nor pi0781 n35324 ; n35337
g32902 nor n35336 n35337 ; n35338
g32903 and pi0789_not n35338 ; n35339
g32904 and pi0619_not n35338 ; n35340
g32905 nor n35050 n35340 ; n35341
g32906 nor pi1159 n35341 ; n35342
g32907 nor pi0648 n35006 ; n35343
g32908 and n35342_not n35343 ; n35344
g32909 and pi0619 n35338 ; n35345
g32910 nor n35108 n35345 ; n35346
g32911 and pi1159 n35346_not ; n35347
g32912 and pi0648 n35002_not ; n35348
g32913 and n35347_not n35348 ; n35349
g32914 and pi0789 n35344_not ; n35350
g32915 and n35349_not n35350 ; n35351
g32916 and n17970 n35339_not ; n35352
g32917 and n35351_not n35352 ; n35353
g32918 and pi0641 n34943_not ; n35354
g32919 and n17865 n35126_not ; n35355
g32920 and n35354_not n35355 ; n35356
g32921 nor n16630 n17870 ; n35357
g32922 and n35009 n35357 ; n35358
g32923 nor pi0641 n34943 ; n35359
g32924 and n17866 n35119_not ; n35360
g32925 and n35359_not n35360 ; n35361
g32926 nor n35356 n35361 ; n35362
g32927 and n35358_not n35362 ; n35363
g32928 and pi0788 n35363_not ; n35364
g32929 nor n20364 n35364 ; n35365
g32930 and n35353_not n35365 ; n35366
g32931 and n20570_not n35012 ; n35367
g32932 and pi1156 n35038 ; n35368
g32933 nor n35045 n35367 ; n35369
g32934 and n35368_not n35369 ; n35370
g32935 and pi0792 n35370_not ; n35371
g32936 nor n35366 n35371 ; n35372
g32937 nor pi0207 n35372 ; n35373
g32938 and pi0623 n35295_not ; n35374
g32939 and n35373_not n35374 ; n35375
g32940 and pi0710 n35375_not ; n35376
g32941 and n35206_not n35376 ; n35377
g32942 nor n20206 n35034 ; n35378
g32943 and n35377_not n35378 ; n35379
g32944 nor n35033 n35379 ; n35380
g32945 and pi0644 n35380 ; n35381
g32946 and pi0715 n34968_not ; n35382
g32947 and n35381_not n35382 ; n35383
g32948 and n17804 n34953_not ; n35384
g32949 and n17804_not n35028 ; n35385
g32950 nor n35384 n35385 ; n35386
g32951 and pi0644 n35386 ; n35387
g32952 and pi0644_not n34953 ; n35388
g32953 nor pi0715 n35388 ; n35389
g32954 and n35387_not n35389 ; n35390
g32955 and pi1160 n35390_not ; n35391
g32956 and n35383_not n35391 ; n35392
g32957 and pi0644 n34967 ; n35393
g32958 and pi0644_not n35380 ; n35394
g32959 nor pi0715 n35393 ; n35395
g32960 and n35394_not n35395 ; n35396
g32961 and pi0644_not n35386 ; n35397
g32962 and pi0644 n34953 ; n35398
g32963 and pi0715 n35398_not ; n35399
g32964 and n35397_not n35399 ; n35400
g32965 nor pi1160 n35400 ; n35401
g32966 and n35396_not n35401 ; n35402
g32967 nor n35392 n35402 ; n35403
g32968 and pi0790 n35403_not ; n35404
g32969 and pi0790_not n35380 ; n35405
g32970 nor n35404 n35405 ; n35406
g32971 nor po1038 n35406 ; n35407
g32972 and pi0207_not po1038 ; n35408
g32973 or n35407 n35408 ; po0364
g32974 and pi0208 n34920_not ; n35410
g32975 nor pi0208 n34949 ; n35411
g32976 nor n35410 n35411 ; n35412
g32977 and pi0638 n35412_not ; n35413
g32978 nor pi0208 n17059 ; n35414
g32979 nor pi0638 n35414 ; n35415
g32980 nor n35413 n35415 ; n35416
g32981 nor pi0787 n35416 ; n35417
g32982 and pi0647_not n35416 ; n35418
g32983 and pi0647 n35414 ; n35419
g32984 nor pi1157 n35419 ; n35420
g32985 and n35418_not n35420 ; n35421
g32986 and pi0647_not n35414 ; n35422
g32987 and pi0647 n35416 ; n35423
g32988 and pi1157 n35422_not ; n35424
g32989 and n35423_not n35424 ; n35425
g32990 nor n35421 n35425 ; n35426
g32991 and pi0787 n35426_not ; n35427
g32992 nor n35417 n35427 ; n35428
g32993 and pi0644_not n35428 ; n35429
g32994 and pi0630_not n35425 ; n35430
g32995 nor pi0208 n35015 ; n35431
g32996 and pi0208 n35023_not ; n35432
g32997 and pi0607 n35432_not ; n35433
g32998 and n35431_not n35433 ; n35434
g32999 and pi0607_not n35414 ; n35435
g33000 nor n35434 n35435 ; n35436
g33001 and n20559_not n35436 ; n35437
g33002 and pi0630 n35421 ; n35438
g33003 nor n35430 n35437 ; n35439
g33004 and n35438_not n35439 ; n35440
g33005 and pi0787 n35440_not ; n35441
g33006 nor pi0638 n35436 ; n35442
g33007 nor pi0208 n35137 ; n35443
g33008 and pi0208 n35203_not ; n35444
g33009 nor pi0607 n35444 ; n35445
g33010 and n35443_not n35445 ; n35446
g33011 and pi0208 n35294_not ; n35447
g33012 nor pi0208 n35372 ; n35448
g33013 and pi0607 n35447_not ; n35449
g33014 and n35448_not n35449 ; n35450
g33015 and pi0638 n35450_not ; n35451
g33016 and n35446_not n35451 ; n35452
g33017 nor n20206 n35442 ; n35453
g33018 and n35452_not n35453 ; n35454
g33019 nor n35441 n35454 ; n35455
g33020 and pi0644 n35455 ; n35456
g33021 and pi0715 n35429_not ; n35457
g33022 and n35456_not n35457 ; n35458
g33023 and n17804 n35414_not ; n35459
g33024 and n17804_not n35436 ; n35460
g33025 nor n35459 n35460 ; n35461
g33026 and pi0644 n35461 ; n35462
g33027 and pi0644_not n35414 ; n35463
g33028 nor pi0715 n35463 ; n35464
g33029 and n35462_not n35464 ; n35465
g33030 and pi1160 n35465_not ; n35466
g33031 and n35458_not n35466 ; n35467
g33032 and pi0644 n35428 ; n35468
g33033 and pi0644_not n35455 ; n35469
g33034 nor pi0715 n35468 ; n35470
g33035 and n35469_not n35470 ; n35471
g33036 and pi0644_not n35461 ; n35472
g33037 and pi0644 n35414 ; n35473
g33038 and pi0715 n35473_not ; n35474
g33039 and n35472_not n35474 ; n35475
g33040 nor pi1160 n35475 ; n35476
g33041 and n35471_not n35476 ; n35477
g33042 nor n35467 n35477 ; n35478
g33043 and pi0790 n35478_not ; n35479
g33044 and pi0790_not n35455 ; n35480
g33045 nor n35479 n35480 ; n35481
g33046 nor po1038 n35481 ; n35482
g33047 and pi0208_not po1038 ; n35483
g33048 or n35482 n35483 ; po0365
g33049 and n10197 n17052 ; n35485
g33050 and pi0639_not n35485 ; n35486
g33051 and pi0715 n17059 ; n35487
g33052 nor n20206 n35137 ; n35488
g33053 nor pi0647 n17059 ; n35489
g33054 and pi0647 n34949 ; n35490
g33055 nor n35489 n35490 ; n35491
g33056 nor pi0630 n35491 ; n35492
g33057 nor n35489 n35492 ; n35493
g33058 and pi1157 n35493_not ; n35494
g33059 and pi0647 n17059_not ; n35495
g33060 and pi1157_not n35495 ; n35496
g33061 and pi0647_not n34949 ; n35497
g33062 nor n35495 n35497 ; n35498
g33063 and n17802 n35498_not ; n35499
g33064 nor n35496 n35499 ; n35500
g33065 and n35494_not n35500 ; n35501
g33066 and pi0787 n35501_not ; n35502
g33067 nor n35488 n35502 ; n35503
g33068 nor pi0644 n35503 ; n35504
g33069 and n19342_not n34949 ; n35505
g33070 and n17059_not n19342 ; n35506
g33071 nor n35505 n35506 ; n35507
g33072 and pi0644 n35507_not ; n35508
g33073 nor pi0715 n35508 ; n35509
g33074 and n35504_not n35509 ; n35510
g33075 nor pi1160 n35487 ; n35511
g33076 and n35510_not n35511 ; n35512
g33077 and pi0715_not n17059 ; n35513
g33078 and pi0644 n35503_not ; n35514
g33079 nor pi0644 n35507 ; n35515
g33080 and pi0715 n35515_not ; n35516
g33081 and n35514_not n35516 ; n35517
g33082 and pi1160 n35513_not ; n35518
g33083 and n35517_not n35518 ; n35519
g33084 nor n35512 n35519 ; n35520
g33085 and pi0790 n35520_not ; n35521
g33086 nor pi0790 n35503 ; n35522
g33087 nor po1038 n35522 ; n35523
g33088 and n35521_not n35523 ; n35524
g33089 and pi0639 n35524 ; n35525
g33090 nor pi0622 n35486 ; n35526
g33091 and n35525_not n35526 ; n35527
g33092 and n17059_not n17804 ; n35528
g33093 and n17804_not n35015 ; n35529
g33094 nor n35528 n35529 ; n35530
g33095 nor pi0790 n35530 ; n35531
g33096 and pi0644 n35530_not ; n35532
g33097 nor pi0644 n17059 ; n35533
g33098 nor n35532 n35533 ; n35534
g33099 and pi1160 n35534 ; n35535
g33100 nor pi0644 n35530 ; n35536
g33101 and pi0644 n17059_not ; n35537
g33102 nor n35536 n35537 ; n35538
g33103 and pi1160_not n35538 ; n35539
g33104 and pi0790 n35535_not ; n35540
g33105 and n35539_not n35540 ; n35541
g33106 nor po1038 n35531 ; n35542
g33107 and n35541_not n35542 ; n35543
g33108 and pi0639_not n35543 ; n35544
g33109 and pi0715 n35538 ; n35545
g33110 nor n20206 n35372 ; n35546
g33111 and n20559_not n35015 ; n35547
g33112 and pi1157 n35492 ; n35548
g33113 nor n35499 n35547 ; n35549
g33114 and n35548_not n35549 ; n35550
g33115 and pi0787 n35550_not ; n35551
g33116 nor n35546 n35551 ; n35552
g33117 nor pi0644 n35552 ; n35553
g33118 and n35509 n35553_not ; n35554
g33119 nor pi1160 n35545 ; n35555
g33120 and n35554_not n35555 ; n35556
g33121 and pi0715_not n35534 ; n35557
g33122 and pi0644 n35552_not ; n35558
g33123 and n35516 n35558_not ; n35559
g33124 and pi1160 n35557_not ; n35560
g33125 and n35559_not n35560 ; n35561
g33126 nor n35556 n35561 ; n35562
g33127 and pi0790 n35562_not ; n35563
g33128 nor pi0790 n35552 ; n35564
g33129 nor po1038 n35564 ; n35565
g33130 and n35563_not n35565 ; n35566
g33131 and pi0639 n35566 ; n35567
g33132 and pi0622 n35544_not ; n35568
g33133 and n35567_not n35568 ; n35569
g33134 nor n35527 n35569 ; n35570
g33135 nor pi0209 n35570 ; n35571
g33136 and pi0644_not pi1160 ; n35572
g33137 and pi0644 pi1160_not ; n35573
g33138 nor n35572 n35573 ; n35574
g33139 and pi0790 n35574_not ; n35575
g33140 and n23684 n35022 ; n35576
g33141 nor po1038 n35575 ; n35577
g33142 and n35576 n35577 ; n35578
g33143 and pi0622 n35578 ; n35579
g33144 nor pi0639 n35579 ; n35580
g33145 nor n20206 n35203 ; n35581
g33146 and n17804 n19341 ; n35582
g33147 and n34920 n35582 ; n35583
g33148 nor n35581 n35583 ; n35584
g33149 and pi0790_not n35584 ; n35585
g33150 and n19342_not n34920 ; n35586
g33151 nor pi0644 n35586 ; n35587
g33152 and pi0715 n35587_not ; n35588
g33153 and pi0644 n35584 ; n35589
g33154 and pi1160 n35588 ; n35590
g33155 and n35589_not n35590 ; n35591
g33156 and pi0644 n35586_not ; n35592
g33157 nor pi0715 n35592 ; n35593
g33158 and pi0644_not n35584 ; n35594
g33159 and pi1160_not n35593 ; n35595
g33160 and n35594_not n35595 ; n35596
g33161 and pi0790 n35591_not ; n35597
g33162 and n35596_not n35597 ; n35598
g33163 nor po1038 n35585 ; n35599
g33164 and n35598_not n35599 ; n35600
g33165 nor pi0622 n35600 ; n35601
g33166 and pi0644_not pi0715 ; n35602
g33167 and n35576 n35602 ; n35603
g33168 and pi0647 n34920 ; n35604
g33169 and pi1157 n35604_not ; n35605
g33170 and pi0647 n35023 ; n35606
g33171 nor pi0647 n35294 ; n35607
g33172 nor pi1157 n35606 ; n35608
g33173 and n35607_not n35608 ; n35609
g33174 nor pi0630 n35605 ; n35610
g33175 and n35609_not n35610 ; n35611
g33176 and pi0647_not n34920 ; n35612
g33177 nor pi1157 n35612 ; n35613
g33178 and pi0647_not n35023 ; n35614
g33179 and pi0647 n35294_not ; n35615
g33180 and pi1157 n35614_not ; n35616
g33181 and n35615_not n35616 ; n35617
g33182 and pi0630 n35613_not ; n35618
g33183 and n35617_not n35618 ; n35619
g33184 nor n35611 n35619 ; n35620
g33185 and pi0787 n35620_not ; n35621
g33186 nor pi0787 n35294 ; n35622
g33187 nor n35621 n35622 ; n35623
g33188 and pi0644_not n35623 ; n35624
g33189 and n35593 n35624_not ; n35625
g33190 nor pi1160 n35603 ; n35626
g33191 and n35625_not n35626 ; n35627
g33192 and pi0644 pi0715_not ; n35628
g33193 and n35576 n35628 ; n35629
g33194 and pi0644 n35623 ; n35630
g33195 and n35588 n35630_not ; n35631
g33196 and pi1160 n35629_not ; n35632
g33197 and n35631_not n35632 ; n35633
g33198 nor n35627 n35633 ; n35634
g33199 and pi0790 n35634_not ; n35635
g33200 and pi0790_not n35623 ; n35636
g33201 nor po1038 n35636 ; n35637
g33202 and n35635_not n35637 ; n35638
g33203 and pi0622 pi0639 ; n35639
g33204 and n35638_not n35639 ; n35640
g33205 and pi0209 n35580_not ; n35641
g33206 and n35601_not n35641 ; n35642
g33207 and n35640_not n35642 ; n35643
g33208 or n35571 n35643 ; po0366
g33209 and pi0210 n16641_not ; n35645
g33210 and pi0634 n20902 ; n35646
g33211 and pi0633 pi0947 ; n35647
g33212 nor n35646 n35647 ; n35648
g33213 and n16641 n35648_not ; n35649
g33214 and pi0038 n35645_not ; n35650
g33215 and n35649_not n35650 ; n35651
g33216 nor n16939 n35648 ; n35652
g33217 and pi0299 n35652_not ; n35653
g33218 and n16940_not n35653 ; n35654
g33219 and pi0210 n16930_not ; n35655
g33220 and n16930 n35648_not ; n35656
g33221 nor pi0299 n35655 ; n35657
g33222 and n35656_not n35657 ; n35658
g33223 nor pi0039 n35654 ; n35659
g33224 and n35658_not n35659 ; n35660
g33225 and pi0210 n16653_not ; n35661
g33226 nor n33589 n35661 ; n35662
g33227 and n6227 n35662 ; n35663
g33228 and pi0947 n35663_not ; n35664
g33229 and pi0210 n16721 ; n35665
g33230 and pi0633 n16721_not ; n35666
g33231 nor n35665 n35666 ; n35667
g33232 and n6227_not n35667 ; n35668
g33233 and n35664 n35668_not ; n35669
g33234 and pi0634 n16653 ; n35670
g33235 nor n35661 n35670 ; n35671
g33236 and n6227 n35671 ; n35672
g33237 and pi0907 n35672_not ; n35673
g33238 nor n33430 n35665 ; n35674
g33239 and n6227_not n35674 ; n35675
g33240 and n35673 n35675_not ; n35676
g33241 and n6227 n16652 ; n35677
g33242 and n2926 n35677 ; n35678
g33243 and n35665 n35678_not ; n35679
g33244 nor n35676 n35679 ; n35680
g33245 nor pi0947 n35680 ; n35681
g33246 nor n6205 n35669 ; n35682
g33247 and n35681_not n35682 ; n35683
g33248 and po1101_not n35662 ; n35684
g33249 and pi0947 n35684_not ; n35685
g33250 nor n6197 n35667 ; n35686
g33251 and po1101 n35662 ; n35687
g33252 nor n6198 n35687 ; n35688
g33253 nor n35686 n35688 ; n35689
g33254 and n35685 n35689_not ; n35690
g33255 nor n6198 n35671 ; n35691
g33256 and pi0907 n35691_not ; n35692
g33257 and n6198 n35674_not ; n35693
g33258 and n35692 n35693_not ; n35694
g33259 and po1101_not n35661 ; n35695
g33260 and pi0210 po1101 ; n35696
g33261 and n16797_not n35696 ; n35697
g33262 nor n35695 n35697 ; n35698
g33263 and pi0907_not n35698 ; n35699
g33264 nor pi0947 n35694 ; n35700
g33265 and n35699_not n35700 ; n35701
g33266 and n6205 n35690_not ; n35702
g33267 and n35701_not n35702 ; n35703
g33268 and pi0223 n35683_not ; n35704
g33269 and n35703_not n35704 ; n35705
g33270 and n16653 n35648_not ; n35706
g33271 nor n35661 n35706 ; n35707
g33272 and n2603 n35707 ; n35708
g33273 and pi0210 n16681 ; n35709
g33274 and pi0633 n16681_not ; n35710
g33275 nor n35709 n35710 ; n35711
g33276 nor n6197 n35711 ; n35712
g33277 nor n35688 n35712 ; n35713
g33278 and n35685 n35713_not ; n35714
g33279 and pi0634 n16681_not ; n35715
g33280 nor n35709 n35715 ; n35716
g33281 and n6198 n35716_not ; n35717
g33282 and n35692 n35717_not ; n35718
g33283 and n16684_not n35696 ; n35719
g33284 nor n35695 n35719 ; n35720
g33285 and pi0907_not n35720 ; n35721
g33286 nor pi0947 n35718 ; n35722
g33287 and n35721_not n35722 ; n35723
g33288 and n6205 n35714_not ; n35724
g33289 and n35723_not n35724 ; n35725
g33290 and n6227_not n35716 ; n35726
g33291 and n35673 n35726_not ; n35727
g33292 and pi0210 n17143_not ; n35728
g33293 and pi0907_not n35728 ; n35729
g33294 nor n35727 n35729 ; n35730
g33295 nor pi0947 n35730 ; n35731
g33296 and n6227_not n35711 ; n35732
g33297 and n35664 n35732_not ; n35733
g33298 nor n6205 n35733 ; n35734
g33299 and n35731_not n35734 ; n35735
g33300 nor n35725 n35735 ; n35736
g33301 nor n2603 n35736 ; n35737
g33302 nor pi0223 n35708 ; n35738
g33303 and n35737_not n35738 ; n35739
g33304 nor pi0299 n35705 ; n35740
g33305 and n35739_not n35740 ; n35741
g33306 nor n6241 n35679 ; n35742
g33307 and n6241 n35698 ; n35743
g33308 nor pi0907 n35742 ; n35744
g33309 and n35743_not n35744 ; n35745
g33310 nor n35676 n35745 ; n35746
g33311 nor pi0947 n35746 ; n35747
g33312 nor n35669 n35747 ; n35748
g33313 and pi0215 n35748_not ; n35749
g33314 and n3448 n35707 ; n35750
g33315 nor n6241 n35728 ; n35751
g33316 and n6241 n35720 ; n35752
g33317 nor pi0907 n35752 ; n35753
g33318 and n35751_not n35753 ; n35754
g33319 nor n35727 n35754 ; n35755
g33320 nor pi0947 n35755 ; n35756
g33321 nor n3448 n35733 ; n35757
g33322 and n35756_not n35757 ; n35758
g33323 nor pi0215 n35750 ; n35759
g33324 and n35758_not n35759 ; n35760
g33325 and pi0299 n35749_not ; n35761
g33326 and n35760_not n35761 ; n35762
g33327 and pi0039 n35762_not ; n35763
g33328 and n35741_not n35763 ; n35764
g33329 nor pi0038 n35660 ; n35765
g33330 and n35764_not n35765 ; n35766
g33331 nor n35651 n35766 ; n35767
g33332 and n10197 n35767_not ; n35768
g33333 nor pi0210 n10197 ; n35769
g33334 nor n35768 n35769 ; po0367
g33335 and n2571 n21641_not ; n35771
g33336 and pi0606_not n35771 ; n35772
g33337 and n2571 n21637_not ; n35773
g33338 and pi0606 n35773 ; n35774
g33339 and pi0643 n35772_not ; n35775
g33340 and n35774_not n35775 ; n35776
g33341 and pi0606_not n17059 ; n35777
g33342 and n2571 n21010_not ; n35778
g33343 and pi0606 n35778 ; n35779
g33344 nor pi0643 n35777 ; n35780
g33345 and n35779_not n35780 ; n35781
g33346 nor po1038 n35781 ; n35782
g33347 and n35776_not n35782 ; n35783
g33348 and pi0211 n35783_not ; n35784
g33349 and n2571 n21628 ; n35785
g33350 nor pi0606 n35785 ; n35786
g33351 and n2571 n21625 ; n35787
g33352 and pi0606 n35787_not ; n35788
g33353 and pi0643 n35786_not ; n35789
g33354 and n35788_not n35789 ; n35790
g33355 and n2571 n21034 ; n35791
g33356 and pi0606 pi0643_not ; n35792
g33357 and n35791 n35792 ; n35793
g33358 nor n35790 n35793 ; n35794
g33359 nor pi0211 po1038 ; n35795
g33360 and n35794_not n35795 ; n35796
g33361 or n35784 n35796 ; po0368
g33362 and pi0607_not n35771 ; n35798
g33363 and pi0607 n35773 ; n35799
g33364 and pi0638 n35798_not ; n35800
g33365 and n35799_not n35800 ; n35801
g33366 and pi0607_not n17059 ; n35802
g33367 and pi0607 n35778 ; n35803
g33368 nor pi0638 n35802 ; n35804
g33369 and n35803_not n35804 ; n35805
g33370 nor po1038 n35805 ; n35806
g33371 and n35801_not n35806 ; n35807
g33372 nor pi0212 n35807 ; n35808
g33373 and pi0607 n35787_not ; n35809
g33374 nor pi0607 n35785 ; n35810
g33375 and pi0638 n35809_not ; n35811
g33376 and n35810_not n35811 ; n35812
g33377 and pi0607 pi0638_not ; n35813
g33378 and n35791 n35813 ; n35814
g33379 nor n35812 n35814 ; n35815
g33380 and pi0212 po1038_not ; n35816
g33381 and n35815_not n35816 ; n35817
g33382 or n35808 n35817 ; po0369
g33383 and pi0213 po1038_not ; n35819
g33384 and pi0622 n35787_not ; n35820
g33385 nor pi0622 n35785 ; n35821
g33386 and pi0639 n35820_not ; n35822
g33387 and n35821_not n35822 ; n35823
g33388 and pi0622 pi0639_not ; n35824
g33389 and n35791 n35824 ; n35825
g33390 nor n35823 n35825 ; n35826
g33391 and n35819 n35826_not ; n35827
g33392 and pi0639_not n35778 ; n35828
g33393 and pi0639 n35773 ; n35829
g33394 and pi0622 n35828_not ; n35830
g33395 and n35829_not n35830 ; n35831
g33396 and pi0639_not n17059 ; n35832
g33397 and pi0639 n35771 ; n35833
g33398 nor pi0622 n35832 ; n35834
g33399 and n35833_not n35834 ; n35835
g33400 nor po1038 n35835 ; n35836
g33401 and n35831_not n35836 ; n35837
g33402 nor pi0213 n35837 ; n35838
g33403 or n35827 n35838 ; po0370
g33404 and pi0623_not n35771 ; n35840
g33405 and pi0623 n35773 ; n35841
g33406 and pi0710 n35840_not ; n35842
g33407 and n35841_not n35842 ; n35843
g33408 and pi0623_not n17059 ; n35844
g33409 and pi0623 n35778 ; n35845
g33410 nor pi0710 n35844 ; n35846
g33411 and n35845_not n35846 ; n35847
g33412 nor po1038 n35847 ; n35848
g33413 and n35843_not n35848 ; n35849
g33414 nor pi0214 n35849 ; n35850
g33415 and pi0623 n35787_not ; n35851
g33416 nor pi0623 n35785 ; n35852
g33417 and pi0710 n35851_not ; n35853
g33418 and n35852_not n35853 ; n35854
g33419 and pi0623 pi0710_not ; n35855
g33420 and n35791 n35855 ; n35856
g33421 nor n35854 n35856 ; n35857
g33422 and pi0214 po1038_not ; n35858
g33423 and n35857_not n35858 ; n35859
g33424 or n35850 n35859 ; po0371
g33425 and pi0215 n10197_not ; n35861
g33426 and pi0681 pi0907 ; n35862
g33427 and pi0947_not n35862 ; n35863
g33428 and pi0642 pi0947 ; n35864
g33429 nor n35863 n35864 ; n35865
g33430 and n16641 n35865_not ; n35866
g33431 and pi0215 n16641_not ; n35867
g33432 and pi0038 n35866_not ; n35868
g33433 and n35867_not n35868 ; n35869
g33434 and pi0215 n16941_not ; n35870
g33435 and n16941 n35865_not ; n35871
g33436 and pi0299 n35870_not ; n35872
g33437 and n35871_not n35872 ; n35873
g33438 and n16930 n35865_not ; n35874
g33439 and pi0215 n16930_not ; n35875
g33440 nor pi0299 n35874 ; n35876
g33441 and n35875_not n35876 ; n35877
g33442 nor pi0039 n35873 ; n35878
g33443 and n35877_not n35878 ; n35879
g33444 and pi0947_not n21326 ; n35880
g33445 and n16656 n16963 ; n35881
g33446 nor n6195 n16814 ; n35882
g33447 nor pi0642 n35881 ; n35883
g33448 and n35882_not n35883 ; n35884
g33449 and pi0947 n35884_not ; n35885
g33450 nor n35863 n35885 ; n35886
g33451 and n35880_not n35886 ; n35887
g33452 and pi0299 n35887_not ; n35888
g33453 and n2603 n35865_not ; n35889
g33454 and n2603 n16653_not ; n35890
g33455 and n21431 n35862_not ; n35891
g33456 and pi0642_not n17143 ; n35892
g33457 nor n6205 n35892 ; n35893
g33458 and pi0642_not n16684 ; n35894
g33459 and n6195 n35894_not ; n35895
g33460 and n16769 n17167 ; n35896
g33461 and n6191_not n16653 ; n35897
g33462 and pi0642_not n35897 ; n35898
g33463 nor n6195 n35898 ; n35899
g33464 and n35896_not n35899 ; n35900
g33465 nor n35895 n35900 ; n35901
g33466 and n6205 n35901_not ; n35902
g33467 and pi0947 n35893_not ; n35903
g33468 and n35902_not n35903 ; n35904
g33469 nor n2603 n35904 ; n35905
g33470 and n35891_not n35905 ; n35906
g33471 nor pi0223 n35889 ; n35907
g33472 and n35890_not n35907 ; n35908
g33473 and n35906_not n35908 ; n35909
g33474 nor n6205 n35884 ; n35910
g33475 and n6195 n16797_not ; n35911
g33476 nor n6195 n16803 ; n35912
g33477 nor pi0642 n35911 ; n35913
g33478 and n35912_not n35913 ; n35914
g33479 and n6205 n35914_not ; n35915
g33480 and pi0947 n35910_not ; n35916
g33481 and n35915_not n35916 ; n35917
g33482 nor n21052 n35917 ; n35918
g33483 and pi0223 n35863_not ; n35919
g33484 and n35918_not n35919 ; n35920
g33485 nor pi0299 n35920 ; n35921
g33486 and n35909_not n35921 ; n35922
g33487 nor n35888 n35922 ; n35923
g33488 and pi0215 n35923_not ; n35924
g33489 and n16653 n35889 ; n35925
g33490 and n16702 n35862 ; n35926
g33491 nor pi0947 n35926 ; n35927
g33492 and pi0642 n16657 ; n35928
g33493 and n6195_not n16699 ; n35929
g33494 nor n17142 n35929 ; n35930
g33495 and n35928 n35930 ; n35931
g33496 and pi0642 n16657_not ; n35932
g33497 and n16699_not n35932 ; n35933
g33498 and pi0947 n35933_not ; n35934
g33499 and n35931_not n35934 ; n35935
g33500 nor n35927 n35935 ; n35936
g33501 nor n6205 n35936 ; n35937
g33502 and n16653 n35932 ; n35938
g33503 and n16974_not n35928 ; n35939
g33504 and n16995_not n35939 ; n35940
g33505 nor n35938 n35940 ; n35941
g33506 and pi0947 n35941_not ; n35942
g33507 and n16776 n35863 ; n35943
g33508 and n6205 n35942_not ; n35944
g33509 and n35943_not n35944 ; n35945
g33510 nor n2603 n35937 ; n35946
g33511 and n35945_not n35946 ; n35947
g33512 nor pi0223 n35925 ; n35948
g33513 and n35947_not n35948 ; n35949
g33514 and n6205 n16803_not ; n35950
g33515 and n35862 n35950_not ; n35951
g33516 nor pi0947 n35951 ; n35952
g33517 and pi0947 n16723_not ; n35953
g33518 nor n16814 n35953 ; n35954
g33519 and n6205_not n35954 ; n35955
g33520 and n16973_not n35939 ; n35956
g33521 and pi0947 n35938_not ; n35957
g33522 and n35956_not n35957 ; n35958
g33523 nor n35955 n35958 ; n35959
g33524 and n35952_not n35959 ; n35960
g33525 and pi0223 n35960_not ; n35961
g33526 nor n35949 n35961 ; n35962
g33527 nor pi0299 n35962 ; n35963
g33528 and n17026 n35865_not ; n35964
g33529 and n3448_not n35936 ; n35965
g33530 and pi0299 n35964_not ; n35966
g33531 and n35965_not n35966 ; n35967
g33532 nor pi0215 n35967 ; n35968
g33533 and n35963_not n35968 ; n35969
g33534 nor n35924 n35969 ; n35970
g33535 and pi0039 n35970_not ; n35971
g33536 nor pi0038 n35879 ; n35972
g33537 and n35971_not n35972 ; n35973
g33538 and n10197 n35869_not ; n35974
g33539 and n35973_not n35974 ; n35975
g33540 or n35861 n35975 ; po0372
g33541 and pi0662 pi0907 ; n35977
g33542 and pi0947_not n35977 ; n35978
g33543 and pi0614 pi0947 ; n35979
g33544 nor n35978 n35979 ; n35980
g33545 and n16641 n35980_not ; n35981
g33546 and pi0216 n16641_not ; n35982
g33547 and pi0038 n35981_not ; n35983
g33548 and n35982_not n35983 ; n35984
g33549 and pi0216 n16941_not ; n35985
g33550 and n16941 n35980_not ; n35986
g33551 and pi0299 n35985_not ; n35987
g33552 and n35986_not n35987 ; n35988
g33553 and n16930 n35980_not ; n35989
g33554 and pi0216 n16930_not ; n35990
g33555 nor pi0299 n35989 ; n35991
g33556 and n35990_not n35991 ; n35992
g33557 nor pi0039 n35988 ; n35993
g33558 and n35992_not n35993 ; n35994
g33559 and n35950_not n35977 ; n35995
g33560 nor pi0947 n35995 ; n35996
g33561 and n16973_not n16997 ; n35997
g33562 and pi0947 n17000_not ; n35998
g33563 and n35997_not n35998 ; n35999
g33564 nor n35955 n35999 ; n36000
g33565 and n35996_not n36000 ; n36001
g33566 and pi0223 n36001_not ; n36002
g33567 and n2603 n35980_not ; n36003
g33568 and n16653 n36003 ; n36004
g33569 and n35930 n35979 ; n36005
g33570 and n16702 n35978 ; n36006
g33571 nor n36005 n36006 ; n36007
g33572 and n6205_not n36007 ; n36008
g33573 and n16776 n35978 ; n36009
g33574 and pi0947 n17001_not ; n36010
g33575 and n6205 n36010_not ; n36011
g33576 and n36009_not n36011 ; n36012
g33577 nor n2603 n36008 ; n36013
g33578 and n36012_not n36013 ; n36014
g33579 nor pi0223 n36004 ; n36015
g33580 and n36014_not n36015 ; n36016
g33581 nor pi0216 n36002 ; n36017
g33582 and n36016_not n36017 ; n36018
g33583 and pi0616_not n16799 ; n36019
g33584 nor n6195 n16978 ; n36020
g33585 and n36019_not n36020 ; n36021
g33586 nor pi0614 n35911 ; n36022
g33587 and n36021_not n36022 ; n36023
g33588 and n6205 n36023_not ; n36024
g33589 nor n17452 n33382 ; n36025
g33590 and n33383_not n36025 ; n36026
g33591 and n17002 n36026_not ; n36027
g33592 nor pi0614 n16721 ; n36028
g33593 and n6195 n36028 ; n36029
g33594 nor n36027 n36029 ; n36030
g33595 and n6205_not n36030 ; n36031
g33596 and pi0947 n36031_not ; n36032
g33597 and n36024_not n36032 ; n36033
g33598 nor n21052 n36033 ; n36034
g33599 and pi0223 n35978_not ; n36035
g33600 and n36034_not n36035 ; n36036
g33601 and pi0614_not n17143 ; n36037
g33602 and pi0947 n36037_not ; n36038
g33603 nor pi0947 n17018 ; n36039
g33604 nor n6205 n35978 ; n36040
g33605 and n36038_not n36040 ; n36041
g33606 and n36039_not n36041 ; n36042
g33607 and pi0947 n17008_not ; n36043
g33608 and pi0947_not n17011 ; n36044
g33609 and n35977_not n36044 ; n36045
g33610 nor n36043 n36045 ; n36046
g33611 and n6205 n36046_not ; n36047
g33612 nor n2603 n36042 ; n36048
g33613 and n36047_not n36048 ; n36049
g33614 nor pi0223 n36003 ; n36050
g33615 and n35890_not n36050 ; n36051
g33616 and n36049_not n36051 ; n36052
g33617 and pi0216 n36036_not ; n36053
g33618 and n36052_not n36053 ; n36054
g33619 nor pi0299 n36018 ; n36055
g33620 and n36054_not n36055 ; n36056
g33621 and n5777 n36007_not ; n36057
g33622 and n17026 n35980_not ; n36058
g33623 and pi0947_not n20994 ; n36059
g33624 nor n35978 n36038 ; n36060
g33625 and n36059_not n36060 ; n36061
g33626 and pi0216 n36061_not ; n36062
g33627 nor n36057 n36058 ; n36063
g33628 and n36062_not n36063 ; n36064
g33629 nor pi0215 n36064 ; n36065
g33630 and n16814 n35977 ; n36066
g33631 nor pi0947 n36066 ; n36067
g33632 and pi0947 n16723 ; n36068
g33633 nor n35999 n36068 ; n36069
g33634 and n36067_not n36069 ; n36070
g33635 nor pi0216 n36070 ; n36071
g33636 and pi0947 n36030 ; n36072
g33637 and pi0216 n35978_not ; n36073
g33638 and n36072_not n36073 ; n36074
g33639 and n35880_not n36074 ; n36075
g33640 and pi0215 n36071_not ; n36076
g33641 and n36075_not n36076 ; n36077
g33642 and pi0299 n36077_not ; n36078
g33643 and n36065_not n36078 ; n36079
g33644 and pi0039 n36056_not ; n36080
g33645 and n36079_not n36080 ; n36081
g33646 nor pi0038 n35994 ; n36082
g33647 and n36081_not n36082 ; n36083
g33648 nor n35984 n36083 ; n36084
g33649 and n10197 n36084_not ; n36085
g33650 nor pi0216 n10197 ; n36086
g33651 nor n36085 n36086 ; po0373
g33652 and pi0695_not n35600 ; n36088
g33653 and pi0217 n36088_not ; n36089
g33654 and pi0695 n35485_not ; n36090
g33655 nor pi0695 n35524 ; n36091
g33656 nor pi0217 n36090 ; n36092
g33657 and n36091_not n36092 ; n36093
g33658 nor pi0612 n36089 ; n36094
g33659 and n36093_not n36094 ; n36095
g33660 and pi0695_not n35638 ; n36096
g33661 and pi0695 n35578 ; n36097
g33662 and pi0217 n36097_not ; n36098
g33663 and n36096_not n36098 ; n36099
g33664 and pi0695 n35543_not ; n36100
g33665 nor pi0695 n35566 ; n36101
g33666 nor pi0217 n36100 ; n36102
g33667 and n36101_not n36102 ; n36103
g33668 and pi0612 n36099_not ; n36104
g33669 and n36103_not n36104 ; n36105
g33670 or n36095 n36105 ; po0374
g33671 nor n34786 n34825 ; n36107
g33672 and n34786 n34891_not ; n36108
g33673 nor n36107 n36108 ; n36109
g33674 nor pi0218 n36109 ; n36110
g33675 and n34786 n34899 ; n36111
g33676 and pi0218 n36111_not ; n36112
g33677 nor n36110 n36112 ; po0375
g33678 nor pi0219 po1038 ; n36114
g33679 and pi0617 n35787_not ; n36115
g33680 nor pi0617 n35785 ; n36116
g33681 and pi0637 n36115_not ; n36117
g33682 and n36116_not n36117 ; n36118
g33683 and pi0617 pi0637_not ; n36119
g33684 and n35791 n36119 ; n36120
g33685 nor n36118 n36120 ; n36121
g33686 and n36114 n36121_not ; n36122
g33687 and pi0617_not n35771 ; n36123
g33688 and pi0617 n35773 ; n36124
g33689 and pi0637 n36123_not ; n36125
g33690 and n36124_not n36125 ; n36126
g33691 and pi0617_not n17059 ; n36127
g33692 and pi0617 n35778 ; n36128
g33693 nor pi0637 n36127 ; n36129
g33694 and n36128_not n36129 ; n36130
g33695 nor po1038 n36130 ; n36131
g33696 and n36126_not n36131 ; n36132
g33697 and pi0219 n36132_not ; n36133
g33698 or n36122 n36133 ; po0376
g33699 nor n34619 n34910 ; n36135
g33700 and n34765_not n34910 ; n36136
g33701 nor n36135 n36136 ; n36137
g33702 nor pi0220 n36137 ; n36138
g33703 and n34774 n34910 ; n36139
g33704 and pi0220 n36139_not ; n36140
g33705 nor n36138 n36140 ; po0377
g33706 and pi0661 pi0907 ; n36142
g33707 and pi0947_not n36142 ; n36143
g33708 and pi0616 pi0947 ; n36144
g33709 nor n36143 n36144 ; n36145
g33710 and n16641 n36145_not ; n36146
g33711 and pi0221 n16641_not ; n36147
g33712 and pi0038 n36146_not ; n36148
g33713 and n36147_not n36148 ; n36149
g33714 and pi0221 n16941_not ; n36150
g33715 and n16941 n36145_not ; n36151
g33716 and pi0299 n36150_not ; n36152
g33717 and n36151_not n36152 ; n36153
g33718 and n16930 n36145_not ; n36154
g33719 and pi0221 n16930_not ; n36155
g33720 nor pi0299 n36154 ; n36156
g33721 and n36155_not n36156 ; n36157
g33722 nor pi0039 n36153 ; n36158
g33723 and n36157_not n36158 ; n36159
g33724 and pi0947 n16980_not ; n36160
g33725 nor n36143 n36160 ; n36161
g33726 and n35950 n36160_not ; n36162
g33727 nor n35955 n36161 ; n36163
g33728 and n36162_not n36163 ; n36164
g33729 and pi0223 n36164_not ; n36165
g33730 and n16653 n36145_not ; n36166
g33731 and n2603 n36166 ; n36167
g33732 nor pi0223 n36167 ; n36168
g33733 and n16976 n16995_not ; n36169
g33734 nor n16979 n36169 ; n36170
g33735 and pi0947 n36170_not ; n36171
g33736 and n16776 n36143 ; n36172
g33737 and n6205 n36171_not ; n36173
g33738 and n36172_not n36173 ; n36174
g33739 and n35930 n36144 ; n36175
g33740 and n16702 n36143 ; n36176
g33741 nor n36175 n36176 ; n36177
g33742 and n6205_not n36177 ; n36178
g33743 nor n2603 n36178 ; n36179
g33744 and n36174_not n36179 ; n36180
g33745 and n36168 n36180_not ; n36181
g33746 nor pi0221 n36165 ; n36182
g33747 and n36181_not n36182 ; n36183
g33748 nor n35892 n35931 ; n36184
g33749 and n16984 n36184_not ; n36185
g33750 and n6197_not n16774 ; n36186
g33751 nor n16697 n36186 ; n36187
g33752 and n16981 n36187_not ; n36188
g33753 and pi0947 n36185_not ; n36189
g33754 and n36188_not n36189 ; n36190
g33755 nor n36039 n36190 ; n36191
g33756 nor n6205 n36191 ; n36192
g33757 and n16774 n16981 ; n36193
g33758 and n16998_not n17008 ; n36194
g33759 and n16984 n36194_not ; n36195
g33760 nor n36193 n36195 ; n36196
g33761 and pi0947 n36196_not ; n36197
g33762 and n6205 n36044_not ; n36198
g33763 and n36197_not n36198 ; n36199
g33764 nor n36143 n36192 ; n36200
g33765 and n36199_not n36200 ; n36201
g33766 nor n2603 n36201 ; n36202
g33767 and n35890_not n36168 ; n36203
g33768 and n36202_not n36203 ; n36204
g33769 and pi0947_not n16990 ; n36205
g33770 and pi0947 n16987_not ; n36206
g33771 and n6205 n36206_not ; n36207
g33772 and n36205_not n36207 ; n36208
g33773 nor pi0947 n16970 ; n36209
g33774 nor n16723 n16800 ; n36210
g33775 nor n6195 n36210 ; n36211
g33776 nor pi0616 n35881 ; n36212
g33777 and n36211_not n36212 ; n36213
g33778 and pi0947 n36213_not ; n36214
g33779 nor n36209 n36214 ; n36215
g33780 nor n6205 n36215 ; n36216
g33781 and pi0223 n36143_not ; n36217
g33782 and n36208_not n36217 ; n36218
g33783 and n36216_not n36218 ; n36219
g33784 and pi0221 n36219_not ; n36220
g33785 and n36204_not n36220 ; n36221
g33786 nor pi0299 n36183 ; n36222
g33787 and n36221_not n36222 ; n36223
g33788 nor n20994 n36142 ; n36224
g33789 nor pi0947 n36224 ; n36225
g33790 and pi0221 n36190_not ; n36226
g33791 and n36225_not n36226 ; n36227
g33792 and pi0216 n36177_not ; n36228
g33793 and pi0216_not n36166 ; n36229
g33794 nor pi0221 n36229 ; n36230
g33795 and n36228_not n36230 ; n36231
g33796 nor pi0215 n36231 ; n36232
g33797 and n36227_not n36232 ; n36233
g33798 and pi0221 n36143_not ; n36234
g33799 and n36214_not n36234 ; n36235
g33800 and n35880_not n36235 ; n36236
g33801 nor n35954 n36161 ; n36237
g33802 nor pi0221 n36237 ; n36238
g33803 and pi0215 n36238_not ; n36239
g33804 and n36236_not n36239 ; n36240
g33805 and pi0299 n36240_not ; n36241
g33806 and n36233_not n36241 ; n36242
g33807 and pi0039 n36223_not ; n36243
g33808 and n36242_not n36243 ; n36244
g33809 nor pi0038 n36159 ; n36245
g33810 and n36244_not n36245 ; n36246
g33811 nor n36149 n36246 ; n36247
g33812 and n10197 n36247_not ; n36248
g33813 nor pi0221 n10197 ; n36249
g33814 nor n36248 n36249 ; po0378
g33815 nor pi0223 n17020 ; n36251
g33816 nor n16993 n36251 ; n36252
g33817 nor pi0299 n36252 ; n36253
g33818 and pi0039 n36253_not ; n36254
g33819 and n17045_not n36254 ; n36255
g33820 nor pi0038 n18147 ; n36256
g33821 and n36255_not n36256 ; n36257
g33822 and n18591 n36257_not ; n36258
g33823 and pi0222 n36258_not ; n36259
g33824 nor n19149 n36259 ; n36260
g33825 and pi0222 n2571_not ; n36261
g33826 and pi0222 n16641_not ; n36262
g33827 and pi0038 n36262_not ; n36263
g33828 and pi0661 n16646 ; n36264
g33829 and n36263 n36264_not ; n36265
g33830 and pi0661 pi0680 ; n36266
g33831 and n16918 n36266_not ; n36267
g33832 nor pi0222 n16918 ; n36268
g33833 and pi0222 n16935 ; n36269
g33834 nor pi0299 n36269 ; n36270
g33835 and n36267_not n36270 ; n36271
g33836 and n36268_not n36271 ; n36272
g33837 and pi0222 n16944 ; n36273
g33838 and n16923 n36266_not ; n36274
g33839 nor pi0222 n16923 ; n36275
g33840 and pi0299 n36273_not ; n36276
g33841 and n36274_not n36276 ; n36277
g33842 and n36275_not n36277 ; n36278
g33843 nor pi0039 n36272 ; n36279
g33844 and n36278_not n36279 ; n36280
g33845 nor pi0661 n17018 ; n36281
g33846 and pi0680 n16758 ; n36282
g33847 nor n16753 n36282 ; n36283
g33848 and pi0661 n36283_not ; n36284
g33849 nor n36281 n36284 ; n36285
g33850 and n6205_not n36285 ; n36286
g33851 and pi0661_not n16994 ; n36287
g33852 nor n6193 n16776 ; n36288
g33853 and pi0662_not n16995 ; n36289
g33854 nor n36288 n36289 ; n36290
g33855 and n16656 n36290_not ; n36291
g33856 and pi0661 n16786_not ; n36292
g33857 nor n36287 n36291 ; n36293
g33858 and n36292_not n36293 ; n36294
g33859 and n6205 n36294 ; n36295
g33860 and pi0222 n36286_not ; n36296
g33861 and n36295_not n36296 ; n36297
g33862 and n16690_not n36266 ; n36298
g33863 and n6205 n36298 ; n36299
g33864 and pi0661 n16703 ; n36300
g33865 and n6205_not n36300 ; n36301
g33866 and pi0224 n36299_not ; n36302
g33867 and n36301_not n36302 ; n36303
g33868 and pi0661 n16739 ; n36304
g33869 nor pi0224 n36304 ; n36305
g33870 nor pi0222 n36305 ; n36306
g33871 and n36303_not n36306 ; n36307
g33872 nor pi0223 n36307 ; n36308
g33873 and n36297_not n36308 ; n36309
g33874 and pi0222_not pi0661 ; n36310
g33875 and n16729 n36310 ; n36311
g33876 and pi0661_not n16960 ; n36312
g33877 and n16656 n16966 ; n36313
g33878 and pi0661 n16818_not ; n36314
g33879 nor n36312 n36314 ; n36315
g33880 and n36313_not n36315 ; n36316
g33881 and n6205_not n36316 ; n36317
g33882 nor pi0661 n16990 ; n36318
g33883 nor n16804 n16809 ; n36319
g33884 and pi0661 n36319_not ; n36320
g33885 nor n36318 n36320 ; n36321
g33886 and n6205 n36321 ; n36322
g33887 and pi0222 n36317_not ; n36323
g33888 and n36322_not n36323 ; n36324
g33889 and pi0223 n36311_not ; n36325
g33890 and n36324_not n36325 ; n36326
g33891 nor n36309 n36326 ; n36327
g33892 nor pi0299 n36327 ; n36328
g33893 and n16744 n36310 ; n36329
g33894 and n6242_not n36316 ; n36330
g33895 and n6242 n36321 ; n36331
g33896 and pi0222 n36330_not ; n36332
g33897 and n36331_not n36332 ; n36333
g33898 nor n36329 n36333 ; n36334
g33899 and pi0215 n36334_not ; n36335
g33900 and pi0222 n16653_not ; n36336
g33901 and n3448 n36336_not ; n36337
g33902 and n36304_not n36337 ; n36338
g33903 and n6242_not n36285 ; n36339
g33904 and n6242 n36294 ; n36340
g33905 and pi0222 n36339_not ; n36341
g33906 and n36340_not n36341 ; n36342
g33907 nor n6242 n36300 ; n36343
g33908 and n6242 n36298_not ; n36344
g33909 nor pi0222 n36343 ; n36345
g33910 and n36344_not n36345 ; n36346
g33911 nor n3448 n36346 ; n36347
g33912 and n36342_not n36347 ; n36348
g33913 nor pi0215 n36338 ; n36349
g33914 and n36348_not n36349 ; n36350
g33915 and pi0299 n36335_not ; n36351
g33916 and n36350_not n36351 ; n36352
g33917 nor n36328 n36352 ; n36353
g33918 and pi0039 n36353_not ; n36354
g33919 nor n36280 n36354 ; n36355
g33920 nor pi0038 n36355 ; n36356
g33921 and n2571 n36265_not ; n36357
g33922 and n36356_not n36357 ; n36358
g33923 nor n36261 n36358 ; n36359
g33924 nor pi0778 n36359 ; n36360
g33925 and pi0625 n36359 ; n36361
g33926 nor pi0625 n36259 ; n36362
g33927 and pi1153 n36362_not ; n36363
g33928 and n36361_not n36363 ; n36364
g33929 and pi0625_not n36359 ; n36365
g33930 and pi0625 n36259_not ; n36366
g33931 nor pi1153 n36366 ; n36367
g33932 and n36365_not n36367 ; n36368
g33933 nor n36364 n36368 ; n36369
g33934 and pi0778 n36369_not ; n36370
g33935 nor n36360 n36370 ; n36371
g33936 nor n17075 n36371 ; n36372
g33937 and n17075 n36259 ; n36373
g33938 nor n36372 n36373 ; n36374
g33939 nor n16639 n36374 ; n36375
g33940 and n16639 n36259 ; n36376
g33941 nor n36375 n36376 ; n36377
g33942 and n16635_not n36377 ; n36378
g33943 and n16631_not n36378 ; n36379
g33944 nor n36260 n36379 ; n36380
g33945 nor n19142 n36380 ; n36381
g33946 and n17856 n36259_not ; n36382
g33947 nor n36381 n36382 ; n36383
g33948 and pi0787_not n36383 ; n36384
g33949 nor pi0647 n36383 ; n36385
g33950 and pi0647 n36259_not ; n36386
g33951 nor pi1157 n36386 ; n36387
g33952 and n36385_not n36387 ; n36388
g33953 and pi0647 n36383_not ; n36389
g33954 nor pi0647 n36259 ; n36390
g33955 and pi1157 n36390_not ; n36391
g33956 and n36389_not n36391 ; n36392
g33957 nor n36388 n36392 ; n36393
g33958 and pi0787 n36393_not ; n36394
g33959 nor n36384 n36394 ; n36395
g33960 and pi0644_not n36395 ; n36396
g33961 and pi0628 n36259_not ; n36397
g33962 nor pi0628 n36380 ; n36398
g33963 and n17777 n36397_not ; n36399
g33964 and n36398_not n36399 ; n36400
g33965 and n17969 n36259_not ; n36401
g33966 and pi0616 n17280 ; n36402
g33967 and n36263 n36402_not ; n36403
g33968 and pi0616_not n17233 ; n36404
g33969 nor pi0222 n17233 ; n36405
g33970 and pi0222 n17139 ; n36406
g33971 nor pi0039 n36404 ; n36407
g33972 and n36405_not n36407 ; n36408
g33973 and n36406_not n36408 ; n36409
g33974 and n6195_not n17235 ; n36410
g33975 nor n17236 n36410 ; n36411
g33976 and pi0616 n36411_not ; n36412
g33977 and pi0222_not n36412 ; n36413
g33978 and n16743_not n36413 ; n36414
g33979 and pi0616 n17182_not ; n36415
g33980 and n16814 n36415_not ; n36416
g33981 nor n16656 n36416 ; n36417
g33982 nor n6193 n16814 ; n36418
g33983 nor n16963 n36415 ; n36419
g33984 and n36418_not n36419 ; n36420
g33985 and n16656 n36420_not ; n36421
g33986 nor n36417 n36421 ; n36422
g33987 and n6242_not n36422 ; n36423
g33988 and pi0616 n17169_not ; n36424
g33989 nor n16802 n36424 ; n36425
g33990 nor n16656 n36425 ; n36426
g33991 and pi0616 n17168 ; n36427
g33992 and n6193 n36427_not ; n36428
g33993 and n16797 n36428 ; n36429
g33994 and n6193_not n36425 ; n36430
g33995 and n16656 n36429_not ; n36431
g33996 and n36430_not n36431 ; n36432
g33997 nor n36426 n36432 ; n36433
g33998 and n6242 n36433 ; n36434
g33999 and pi0222 n36423_not ; n36435
g34000 and n36434_not n36435 ; n36436
g34001 nor n36414 n36436 ; n36437
g34002 and pi0215 n36437_not ; n36438
g34003 and n16978 n17168 ; n36439
g34004 and n36337 n36439_not ; n36440
g34005 nor n16775 n36424 ; n36441
g34006 nor n16656 n36441 ; n36442
g34007 and n16684 n36428 ; n36443
g34008 and n6193_not n36441 ; n36444
g34009 and n16656 n36443_not ; n36445
g34010 and n36444_not n36445 ; n36446
g34011 nor n36442 n36446 ; n36447
g34012 and n6242 n36447 ; n36448
g34013 and pi0616 n17154_not ; n36449
g34014 and pi0616_not n36187 ; n36450
g34015 nor n36449 n36450 ; n36451
g34016 nor n16656 n36451 ; n36452
g34017 and n17147 n36427_not ; n36453
g34018 nor n17145 n36453 ; n36454
g34019 and n6193 n36454_not ; n36455
g34020 and n6193_not n36451 ; n36456
g34021 and n16656 n36455_not ; n36457
g34022 and n36456_not n36457 ; n36458
g34023 nor n36452 n36458 ; n36459
g34024 and n6242_not n36459 ; n36460
g34025 and pi0222 n36448_not ; n36461
g34026 and n36460_not n36461 ; n36462
g34027 nor n17247 n36410 ; n36463
g34028 and pi0616 n36463_not ; n36464
g34029 and n6242 n36464_not ; n36465
g34030 and n16699_not n36427 ; n36466
g34031 nor n16656 n36466 ; n36467
g34032 and pi0616 n6193 ; n36468
g34033 and n17375 n36468 ; n36469
g34034 and n6193_not n36466 ; n36470
g34035 and n16656 n36469_not ; n36471
g34036 and n36470_not n36471 ; n36472
g34037 nor n36467 n36472 ; n36473
g34038 nor n6242 n36473 ; n36474
g34039 nor pi0222 n36465 ; n36475
g34040 and n36474_not n36475 ; n36476
g34041 nor n3448 n36476 ; n36477
g34042 and n36462_not n36477 ; n36478
g34043 nor pi0215 n36440 ; n36479
g34044 and n36478_not n36479 ; n36480
g34045 and pi0299 n36438_not ; n36481
g34046 and n36480_not n36481 ; n36482
g34047 and n6205 n36464 ; n36483
g34048 and n6205_not n36473 ; n36484
g34049 and pi0224 n36483_not ; n36485
g34050 and n36484_not n36485 ; n36486
g34051 nor pi0224 n36439 ; n36487
g34052 nor pi0222 n36487 ; n36488
g34053 and n36486_not n36488 ; n36489
g34054 and n6205 n36447 ; n36490
g34055 and n6205_not n36459 ; n36491
g34056 and pi0222 n36490_not ; n36492
g34057 and n36491_not n36492 ; n36493
g34058 nor pi0223 n36489 ; n36494
g34059 and n36493_not n36494 ; n36495
g34060 and n16724_not n36413 ; n36496
g34061 and n6205_not n36422 ; n36497
g34062 and n6205 n36433 ; n36498
g34063 and pi0222 n36497_not ; n36499
g34064 and n36498_not n36499 ; n36500
g34065 and pi0223 n36496_not ; n36501
g34066 and n36500_not n36501 ; n36502
g34067 nor n36495 n36502 ; n36503
g34068 nor pi0299 n36503 ; n36504
g34069 and pi0039 n36482_not ; n36505
g34070 and n36504_not n36505 ; n36506
g34071 nor pi0038 n36409 ; n36507
g34072 and n36506_not n36507 ; n36508
g34073 and n2571 n36403_not ; n36509
g34074 and n36508_not n36509 ; n36510
g34075 nor n36261 n36510 ; n36511
g34076 nor n17117 n36511 ; n36512
g34077 and n17117 n36259 ; n36513
g34078 nor n36512 n36513 ; n36514
g34079 nor pi0785 n36514 ; n36515
g34080 and pi0609 n36514 ; n36516
g34081 nor pi0609 n36259 ; n36517
g34082 and pi1155 n36517_not ; n36518
g34083 and n36516_not n36518 ; n36519
g34084 and pi0609_not n36514 ; n36520
g34085 and pi0609 n36259_not ; n36521
g34086 nor pi1155 n36521 ; n36522
g34087 and n36520_not n36522 ; n36523
g34088 nor n36519 n36523 ; n36524
g34089 and pi0785 n36524_not ; n36525
g34090 nor n36515 n36525 ; n36526
g34091 nor pi0781 n36526 ; n36527
g34092 and pi0618 n36526 ; n36528
g34093 nor pi0618 n36259 ; n36529
g34094 and pi1154 n36529_not ; n36530
g34095 and n36528_not n36530 ; n36531
g34096 and pi0618_not n36526 ; n36532
g34097 and pi0618 n36259_not ; n36533
g34098 nor pi1154 n36533 ; n36534
g34099 and n36532_not n36534 ; n36535
g34100 nor n36531 n36535 ; n36536
g34101 and pi0781 n36536_not ; n36537
g34102 nor n36527 n36537 ; n36538
g34103 nor pi0789 n36538 ; n36539
g34104 and pi0619 n36538 ; n36540
g34105 nor pi0619 n36259 ; n36541
g34106 and pi1159 n36541_not ; n36542
g34107 and n36540_not n36542 ; n36543
g34108 and pi0619_not n36538 ; n36544
g34109 and pi0619 n36259_not ; n36545
g34110 nor pi1159 n36545 ; n36546
g34111 and n36544_not n36546 ; n36547
g34112 nor n36543 n36547 ; n36548
g34113 and pi0789 n36548_not ; n36549
g34114 nor n36539 n36549 ; n36550
g34115 and n17969_not n36550 ; n36551
g34116 nor n36401 n36551 ; n36552
g34117 and n20570_not n36552 ; n36553
g34118 nor pi0628 n36259 ; n36554
g34119 and pi0628 n36380_not ; n36555
g34120 and n17776 n36554_not ; n36556
g34121 and n36555_not n36556 ; n36557
g34122 nor n36400 n36557 ; n36558
g34123 and n36553_not n36558 ; n36559
g34124 and pi0792 n36559_not ; n36560
g34125 and pi0609 n36371 ; n36561
g34126 and n16667 n17493 ; n36562
g34127 nor pi0222 pi0616 ; n36563
g34128 and pi0039_not pi0616 ; n36564
g34129 and n36266 n36564 ; n36565
g34130 nor n36563 n36565 ; n36566
g34131 and n36562 n36566_not ; n36567
g34132 nor n36266 n36427 ; n36568
g34133 nor pi0616 n17355 ; n36569
g34134 nor n36568 n36569 ; n36570
g34135 and n16641 n36570 ; n36571
g34136 nor n36262 n36571 ; n36572
g34137 nor n36567 n36572 ; n36573
g34138 and pi0038 n36573_not ; n36574
g34139 and pi0661_not pi0681 ; n36575
g34140 and n36425_not n36575 ; n36576
g34141 and pi0680_not n36425 ; n36577
g34142 and pi0616 n17504_not ; n36578
g34143 and pi0680 n36578_not ; n36579
g34144 and n17347_not n36579 ; n36580
g34145 and pi0661 n36577_not ; n36581
g34146 and n36580_not n36581 ; n36582
g34147 nor n36432 n36576 ; n36583
g34148 and n36582_not n36583 ; n36584
g34149 and n6242 n36584_not ; n36585
g34150 and n36416_not n36575 ; n36586
g34151 and pi0680_not n36416 ; n36587
g34152 and n17324_not n17493 ; n36588
g34153 and pi0616 n36588_not ; n36589
g34154 and pi0680 n36589_not ; n36590
g34155 and n17330 n36590 ; n36591
g34156 and pi0661 n36591_not ; n36592
g34157 and n36587_not n36592 ; n36593
g34158 nor n36421 n36586 ; n36594
g34159 and n36593_not n36594 ; n36595
g34160 nor n6242 n36595 ; n36596
g34161 and pi0222 n36585_not ; n36597
g34162 and n36596_not n36597 ; n36598
g34163 and n17444 n36266 ; n36599
g34164 nor n36412 n36599 ; n36600
g34165 and n6242 n36600_not ; n36601
g34166 and pi0616 n17237 ; n36602
g34167 nor pi0661 n36602 ; n36603
g34168 and n16721_not n36439 ; n36604
g34169 and n6195 n36604_not ; n36605
g34170 and pi0680_not n36602 ; n36606
g34171 nor n17237 n17559 ; n36607
g34172 and pi0616 n36607 ; n36608
g34173 and pi0680 n36608_not ; n36609
g34174 and n17458 n36609 ; n36610
g34175 and pi0661 n36606_not ; n36611
g34176 and n36610_not n36611 ; n36612
g34177 nor n36603 n36605 ; n36613
g34178 and n36612_not n36613 ; n36614
g34179 and n6242_not n36614 ; n36615
g34180 nor pi0222 n36601 ; n36616
g34181 and n36615_not n36616 ; n36617
g34182 and pi0215 n36617_not ; n36618
g34183 and n36598_not n36618 ; n36619
g34184 and pi0616 n17548_not ; n36620
g34185 nor pi0616 n17407 ; n36621
g34186 nor n36620 n36621 ; n36622
g34187 and n36568_not n36622 ; n36623
g34188 and n36337 n36623_not ; n36624
g34189 and n36451_not n36575 ; n36625
g34190 and pi0603 n16681 ; n36626
g34191 and n6197 n16754 ; n36627
g34192 nor n16756 n36627 ; n36628
g34193 and pi0603_not n36628 ; n36629
g34194 nor n17368 n36626 ; n36630
g34195 and n36629_not n36630 ; n36631
g34196 and pi0642_not n36631 ; n36632
g34197 and n17577_not n36628 ; n36633
g34198 and pi0642 n36633_not ; n36634
g34199 and n6191 n36632_not ; n36635
g34200 and n36634_not n36635 ; n36636
g34201 and n17452 n36633 ; n36637
g34202 and n17493 n36628_not ; n36638
g34203 and pi0616 n36638_not ; n36639
g34204 and pi0680 n36639_not ; n36640
g34205 and n36637_not n36640 ; n36641
g34206 and n36636_not n36641 ; n36642
g34207 and pi0680_not n36451 ; n36643
g34208 and pi0661 n36642_not ; n36644
g34209 and n36643_not n36644 ; n36645
g34210 nor n36458 n36625 ; n36646
g34211 and n36645_not n36646 ; n36647
g34212 nor n6242 n36647 ; n36648
g34213 and n36441_not n36575 ; n36649
g34214 and pi0680_not n36441 ; n36650
g34215 and n17363_not n36579 ; n36651
g34216 and pi0661 n36650_not ; n36652
g34217 and n36651_not n36652 ; n36653
g34218 nor n36446 n36649 ; n36654
g34219 and n36653_not n36654 ; n36655
g34220 and n6242 n36655_not ; n36656
g34221 and pi0222 n36656_not ; n36657
g34222 and n36648_not n36657 ; n36658
g34223 and n36466_not n36575 ; n36659
g34224 and pi0680_not n36466 ; n36660
g34225 and pi0616 n17578 ; n36661
g34226 and pi0680 n36661_not ; n36662
g34227 and n17433_not n36662 ; n36663
g34228 and pi0661 n36660_not ; n36664
g34229 and n36663_not n36664 ; n36665
g34230 nor n36472 n36659 ; n36666
g34231 and n36665_not n36666 ; n36667
g34232 and n6242_not n36667 ; n36668
g34233 and n6193_not n36439 ; n36669
g34234 and n17246 n36468 ; n36670
g34235 and n16656 n36669_not ; n36671
g34236 and n36670_not n36671 ; n36672
g34237 and n36439_not n36575 ; n36673
g34238 and pi0680_not n36439 ; n36674
g34239 and pi0680 n17417_not ; n36675
g34240 and n36620_not n36675 ; n36676
g34241 and pi0661 n36674_not ; n36677
g34242 and n36676_not n36677 ; n36678
g34243 nor n36672 n36673 ; n36679
g34244 and n36678_not n36679 ; n36680
g34245 and n6242 n36680 ; n36681
g34246 nor pi0222 n36681 ; n36682
g34247 and n36668_not n36682 ; n36683
g34248 nor n36658 n36683 ; n36684
g34249 nor n3448 n36684 ; n36685
g34250 nor pi0215 n36624 ; n36686
g34251 and n36685_not n36686 ; n36687
g34252 and pi0299 n36619_not ; n36688
g34253 and n36687_not n36688 ; n36689
g34254 and n36266 n36622_not ; n36690
g34255 nor n36266 n36439 ; n36691
g34256 nor pi0222 n36691 ; n36692
g34257 and n36690_not n36692 ; n36693
g34258 nor n3351 n36693 ; n36694
g34259 and n6205_not n36667 ; n36695
g34260 and n6205 n36680 ; n36696
g34261 and pi0224 n36696_not ; n36697
g34262 and n36695_not n36697 ; n36698
g34263 nor n36694 n36698 ; n36699
g34264 and n6205 n36655 ; n36700
g34265 and n6205_not n36647 ; n36701
g34266 and pi0222 n36700_not ; n36702
g34267 and n36701_not n36702 ; n36703
g34268 nor n36699 n36703 ; n36704
g34269 nor pi0223 n36704 ; n36705
g34270 and n6205 n36584_not ; n36706
g34271 nor n6205 n36595 ; n36707
g34272 and pi0222 n36706_not ; n36708
g34273 and n36707_not n36708 ; n36709
g34274 and n6205 n36600_not ; n36710
g34275 and n6205_not n36614 ; n36711
g34276 nor pi0222 n36710 ; n36712
g34277 and n36711_not n36712 ; n36713
g34278 and pi0223 n36713_not ; n36714
g34279 and n36709_not n36714 ; n36715
g34280 nor pi0299 n36715 ; n36716
g34281 and n36705_not n36716 ; n36717
g34282 and pi0039 n36717_not ; n36718
g34283 and n36689_not n36718 ; n36719
g34284 and pi0661 n17618 ; n36720
g34285 and pi0616 n17226 ; n36721
g34286 nor pi0222 n36721 ; n36722
g34287 and n36720_not n36722 ; n36723
g34288 and pi0616_not n17226 ; n36724
g34289 and n17617 n36266_not ; n36725
g34290 nor pi0603 n16935 ; n36726
g34291 nor n17367 n17614 ; n36727
g34292 and n36726_not n36727 ; n36728
g34293 nor n36724 n36728 ; n36729
g34294 and n36725_not n36729 ; n36730
g34295 and pi0222 n36730_not ; n36731
g34296 nor n36723 n36731 ; n36732
g34297 nor pi0299 n36732 ; n36733
g34298 and pi0616_not n17231 ; n36734
g34299 and n17622 n36266_not ; n36735
g34300 nor pi0603 n16944 ; n36736
g34301 nor n17123 n17367 ; n36737
g34302 and n36736_not n36737 ; n36738
g34303 nor n36734 n36738 ; n36739
g34304 and n36735_not n36739 ; n36740
g34305 and pi0222 n36740_not ; n36741
g34306 and pi0661 n17623 ; n36742
g34307 and pi0616 n17231 ; n36743
g34308 nor pi0222 n36743 ; n36744
g34309 and n36742_not n36744 ; n36745
g34310 nor n36741 n36745 ; n36746
g34311 and pi0299 n36746_not ; n36747
g34312 nor pi0039 n36733 ; n36748
g34313 and n36747_not n36748 ; n36749
g34314 nor pi0038 n36749 ; n36750
g34315 and n36719_not n36750 ; n36751
g34316 and n2571 n36574_not ; n36752
g34317 and n36751_not n36752 ; n36753
g34318 nor n36261 n36753 ; n36754
g34319 and pi0625_not n36754 ; n36755
g34320 and pi0625 n36511 ; n36756
g34321 nor pi1153 n36756 ; n36757
g34322 and n36755_not n36757 ; n36758
g34323 nor pi0608 n36364 ; n36759
g34324 and n36758_not n36759 ; n36760
g34325 and pi0625_not n36511 ; n36761
g34326 and pi0625 n36754 ; n36762
g34327 and pi1153 n36761_not ; n36763
g34328 and n36762_not n36763 ; n36764
g34329 and pi0608 n36368_not ; n36765
g34330 and n36764_not n36765 ; n36766
g34331 nor n36760 n36766 ; n36767
g34332 and pi0778 n36767_not ; n36768
g34333 and pi0778_not n36754 ; n36769
g34334 nor n36768 n36769 ; n36770
g34335 nor pi0609 n36770 ; n36771
g34336 nor pi1155 n36561 ; n36772
g34337 and n36771_not n36772 ; n36773
g34338 nor pi0660 n36519 ; n36774
g34339 and n36773_not n36774 ; n36775
g34340 and pi0609_not n36371 ; n36776
g34341 and pi0609 n36770_not ; n36777
g34342 and pi1155 n36776_not ; n36778
g34343 and n36777_not n36778 ; n36779
g34344 and pi0660 n36523_not ; n36780
g34345 and n36779_not n36780 ; n36781
g34346 nor n36775 n36781 ; n36782
g34347 and pi0785 n36782_not ; n36783
g34348 nor pi0785 n36770 ; n36784
g34349 nor n36783 n36784 ; n36785
g34350 nor pi0618 n36785 ; n36786
g34351 and pi0618 n36374 ; n36787
g34352 nor pi1154 n36787 ; n36788
g34353 and n36786_not n36788 ; n36789
g34354 nor pi0627 n36531 ; n36790
g34355 and n36789_not n36790 ; n36791
g34356 and pi0618_not n36374 ; n36792
g34357 and pi0618 n36785_not ; n36793
g34358 and pi1154 n36792_not ; n36794
g34359 and n36793_not n36794 ; n36795
g34360 and pi0627 n36535_not ; n36796
g34361 and n36795_not n36796 ; n36797
g34362 nor n36791 n36797 ; n36798
g34363 and pi0781 n36798_not ; n36799
g34364 nor pi0781 n36785 ; n36800
g34365 nor n36799 n36800 ; n36801
g34366 and pi0789_not n36801 ; n36802
g34367 and pi0626_not n36550 ; n36803
g34368 and pi0626 n36259_not ; n36804
g34369 and n16629 n36804_not ; n36805
g34370 and n36803_not n36805 ; n36806
g34371 and n16635 n36259_not ; n36807
g34372 and n17871 n36807_not ; n36808
g34373 and n36378_not n36808 ; n36809
g34374 and pi0626 n36550 ; n36810
g34375 nor pi0626 n36259 ; n36811
g34376 and n16628 n36811_not ; n36812
g34377 and n36810_not n36812 ; n36813
g34378 nor n36806 n36809 ; n36814
g34379 and n36813_not n36814 ; n36815
g34380 and pi0788 n36815_not ; n36816
g34381 nor pi0619 n36801 ; n36817
g34382 and pi0619 n36377 ; n36818
g34383 nor pi1159 n36818 ; n36819
g34384 and n36817_not n36819 ; n36820
g34385 nor pi0648 n36543 ; n36821
g34386 and n36820_not n36821 ; n36822
g34387 and pi0619 n36801_not ; n36823
g34388 and pi0619_not n36377 ; n36824
g34389 and pi1159 n36824_not ; n36825
g34390 and n36823_not n36825 ; n36826
g34391 and pi0648 n36547_not ; n36827
g34392 and n36826_not n36827 ; n36828
g34393 and pi0789 n36822_not ; n36829
g34394 and n36828_not n36829 ; n36830
g34395 nor n36802 n36816 ; n36831
g34396 and n36830_not n36831 ; n36832
g34397 and n17970_not n36815 ; n36833
g34398 nor n20364 n36833 ; n36834
g34399 and n36832_not n36834 ; n36835
g34400 nor n36560 n36835 ; n36836
g34401 nor n20206 n36836 ; n36837
g34402 and pi0630_not n36392 ; n36838
g34403 and n17779_not n36552 ; n36839
g34404 and n17779 n36259 ; n36840
g34405 nor n36839 n36840 ; n36841
g34406 nor n20559 n36841 ; n36842
g34407 and pi0630 n36388 ; n36843
g34408 nor n36838 n36843 ; n36844
g34409 and n36842_not n36844 ; n36845
g34410 and pi0787 n36845_not ; n36846
g34411 nor n36837 n36846 ; n36847
g34412 and pi0644 n36847 ; n36848
g34413 and pi0715 n36396_not ; n36849
g34414 and n36848_not n36849 ; n36850
g34415 and n17804 n36259_not ; n36851
g34416 and n17804_not n36841 ; n36852
g34417 nor n36851 n36852 ; n36853
g34418 and pi0644 n36853_not ; n36854
g34419 nor pi0644 n36259 ; n36855
g34420 nor pi0715 n36855 ; n36856
g34421 and n36854_not n36856 ; n36857
g34422 and pi1160 n36857_not ; n36858
g34423 and n36850_not n36858 ; n36859
g34424 and pi0644 n36395 ; n36860
g34425 and pi0644_not n36847 ; n36861
g34426 nor pi0715 n36860 ; n36862
g34427 and n36861_not n36862 ; n36863
g34428 nor pi0644 n36853 ; n36864
g34429 and pi0644 n36259_not ; n36865
g34430 and pi0715 n36865_not ; n36866
g34431 and n36864_not n36866 ; n36867
g34432 nor pi1160 n36867 ; n36868
g34433 and n36863_not n36868 ; n36869
g34434 nor n36859 n36869 ; n36870
g34435 and pi0790 n36870_not ; n36871
g34436 and pi0790_not n36847 ; n36872
g34437 nor n36871 n36872 ; n36873
g34438 nor po1038 n36873 ; n36874
g34439 and pi0222_not po1038 ; n36875
g34440 nor n36874 n36875 ; po0379
g34441 nor pi0299 n16992 ; n36877
g34442 and pi0039 n36877_not ; n36878
g34443 and n17045_not n36878 ; n36879
g34444 and n14873 n18147_not ; n36880
g34445 and n36879_not n36880 ; n36881
g34446 and n18591 n36881_not ; n36882
g34447 and pi0223 n36882_not ; n36883
g34448 nor n19149 n36883 ; n36884
g34449 and n17075 n36883_not ; n36885
g34450 and pi0223 n2571_not ; n36886
g34451 and pi0680 pi0681 ; n36887
g34452 and n16918 n36887_not ; n36888
g34453 nor pi0223 n16918 ; n36889
g34454 and pi0223 n16935 ; n36890
g34455 nor pi0299 n36890 ; n36891
g34456 and n36888_not n36891 ; n36892
g34457 and n36889_not n36892 ; n36893
g34458 and pi0223 n16944 ; n36894
g34459 and n16923 n36887_not ; n36895
g34460 nor pi0223 n16923 ; n36896
g34461 and pi0299 n36894_not ; n36897
g34462 and n36895_not n36897 ; n36898
g34463 and n36896_not n36898 ; n36899
g34464 nor pi0039 n36893 ; n36900
g34465 and n36899_not n36900 ; n36901
g34466 and pi0681 n16739 ; n36902
g34467 and n2603 n36902_not ; n36903
g34468 and n16690_not n36887 ; n36904
g34469 and n6205 n36904 ; n36905
g34470 and pi0681 n16703 ; n36906
g34471 and n6205_not n36906 ; n36907
g34472 nor n2603 n36905 ; n36908
g34473 and n36907_not n36908 ; n36909
g34474 nor n36903 n36909 ; n36910
g34475 nor pi0223 n36910 ; n36911
g34476 and pi0681 n36319_not ; n36912
g34477 nor n16989 n36912 ; n36913
g34478 and n6205 n36913_not ; n36914
g34479 and pi0681 n16818_not ; n36915
g34480 nor n16969 n36915 ; n36916
g34481 nor n6205 n36916 ; n36917
g34482 and pi0223 n36914_not ; n36918
g34483 and n36917_not n36918 ; n36919
g34484 nor pi0299 n36919 ; n36920
g34485 and n36911_not n36920 ; n36921
g34486 and pi0223_not pi0681 ; n36922
g34487 and n16744 n36922 ; n36923
g34488 and n6242 n36913 ; n36924
g34489 and n6242_not n36916 ; n36925
g34490 and pi0223 n36924_not ; n36926
g34491 and n36925_not n36926 ; n36927
g34492 and pi0215 n36923_not ; n36928
g34493 and n36927_not n36928 ; n36929
g34494 and pi0223 n16653_not ; n36930
g34495 and n3448 n36930_not ; n36931
g34496 and n36902_not n36931 ; n36932
g34497 and pi0681 n36283_not ; n36933
g34498 nor n6242 n17017 ; n36934
g34499 and n36933_not n36934 ; n36935
g34500 and pi0681 n16786_not ; n36936
g34501 and n6242 n17010_not ; n36937
g34502 and n36936_not n36937 ; n36938
g34503 and pi0223 n36935_not ; n36939
g34504 and n36938_not n36939 ; n36940
g34505 nor n6242 n36906 ; n36941
g34506 and n6242 n36904_not ; n36942
g34507 nor pi0223 n36941 ; n36943
g34508 and n36942_not n36943 ; n36944
g34509 nor n3448 n36944 ; n36945
g34510 and n36940_not n36945 ; n36946
g34511 nor n36932 n36946 ; n36947
g34512 nor pi0215 n36947 ; n36948
g34513 and pi0299 n36929_not ; n36949
g34514 and n36948_not n36949 ; n36950
g34515 and pi0039 n36921_not ; n36951
g34516 and n36950_not n36951 ; n36952
g34517 nor n36901 n36952 ; n36953
g34518 nor pi0038 n36953 ; n36954
g34519 and pi0681 n16646 ; n36955
g34520 and pi0223 n16641_not ; n36956
g34521 and pi0038 n36955_not ; n36957
g34522 and n36956_not n36957 ; n36958
g34523 and n2571 n36958_not ; n36959
g34524 and n36954_not n36959 ; n36960
g34525 nor n36886 n36960 ; n36961
g34526 nor pi0778 n36961 ; n36962
g34527 and pi0625 n36961 ; n36963
g34528 nor pi0625 n36883 ; n36964
g34529 and pi1153 n36964_not ; n36965
g34530 and n36963_not n36965 ; n36966
g34531 and pi0625_not n36961 ; n36967
g34532 and pi0625 n36883_not ; n36968
g34533 nor pi1153 n36968 ; n36969
g34534 and n36967_not n36969 ; n36970
g34535 nor n36966 n36970 ; n36971
g34536 and pi0778 n36971_not ; n36972
g34537 nor n36962 n36972 ; n36973
g34538 and n17075_not n36973 ; n36974
g34539 nor n36885 n36974 ; n36975
g34540 and n16639_not n36975 ; n36976
g34541 and n16639 n36883 ; n36977
g34542 nor n36976 n36977 ; n36978
g34543 and n16635_not n36978 ; n36979
g34544 and n16631_not n36979 ; n36980
g34545 nor n36884 n36980 ; n36981
g34546 nor n19142 n36981 ; n36982
g34547 and n17856 n36883_not ; n36983
g34548 nor n36982 n36983 ; n36984
g34549 and pi0787_not n36984 ; n36985
g34550 nor pi0647 n36984 ; n36986
g34551 and pi0647 n36883_not ; n36987
g34552 nor pi1157 n36987 ; n36988
g34553 and n36986_not n36988 ; n36989
g34554 and pi0647 n36984_not ; n36990
g34555 nor pi0647 n36883 ; n36991
g34556 and pi1157 n36991_not ; n36992
g34557 and n36990_not n36992 ; n36993
g34558 nor n36989 n36993 ; n36994
g34559 and pi0787 n36994_not ; n36995
g34560 nor n36985 n36995 ; n36996
g34561 and pi0644_not n36996 ; n36997
g34562 and pi0630_not n36993 ; n36998
g34563 and n17969 n36883_not ; n36999
g34564 and n17117 n36883_not ; n37000
g34565 and pi0039 pi0223 ; n37001
g34566 and pi0038 n37001_not ; n37002
g34567 and pi0642 n17168 ; n37003
g34568 and n16667 n37003_not ; n37004
g34569 nor pi0223 n16667 ; n37005
g34570 nor pi0039 n37005 ; n37006
g34571 and n37004_not n37006 ; n37007
g34572 and n37002 n37007_not ; n37008
g34573 and pi0223_not pi0642 ; n37009
g34574 and n17226 n37009 ; n37010
g34575 nor pi0299 n37010 ; n37011
g34576 and pi0642_not n17226 ; n37012
g34577 and pi0223 n37012_not ; n37013
g34578 and n17137 n37013 ; n37014
g34579 and n37011 n37014_not ; n37015
g34580 and n17231 n37009 ; n37016
g34581 and pi0299 n37016_not ; n37017
g34582 and n6190 n17230 ; n37018
g34583 and pi0223 n17124_not ; n37019
g34584 and n37018_not n37019 ; n37020
g34585 and n37017 n37020_not ; n37021
g34586 nor pi0039 n37021 ; n37022
g34587 and n37015_not n37022 ; n37023
g34588 and n35897 n37003_not ; n37024
g34589 and pi0642 n17169_not ; n37025
g34590 and n36425 n37025_not ; n37026
g34591 nor n37024 n37026 ; n37027
g34592 and pi0681 n37027 ; n37028
g34593 and n6194 n37004 ; n37029
g34594 and n16797 n37029 ; n37030
g34595 nor n6194 n37027 ; n37031
g34596 nor pi0681 n37030 ; n37032
g34597 and n37031_not n37032 ; n37033
g34598 nor n37028 n37033 ; n37034
g34599 and n6205 n37034 ; n37035
g34600 nor pi0642 n16814 ; n37036
g34601 and pi0642 n17183_not ; n37037
g34602 nor n37036 n37037 ; n37038
g34603 and n6194_not n37038 ; n37039
g34604 and pi0642 n17182_not ; n37040
g34605 and n6194 n37040_not ; n37041
g34606 and n16721_not n37041 ; n37042
g34607 nor pi0681 n37042 ; n37043
g34608 and n37039_not n37043 ; n37044
g34609 and pi0681 n37038_not ; n37045
g34610 nor n37044 n37045 ; n37046
g34611 and n6205_not n37046 ; n37047
g34612 and pi0223 n37047_not ; n37048
g34613 and n37035_not n37048 ; n37049
g34614 and pi0642 n17235 ; n37050
g34615 and n2603 n37050_not ; n37051
g34616 and n6194_not n37050 ; n37052
g34617 nor pi0681 n37052 ; n37053
g34618 and pi0642 n6194 ; n37054
g34619 and n17246 n37054 ; n37055
g34620 and n37053 n37055_not ; n37056
g34621 and pi0681 n37050_not ; n37057
g34622 nor n37056 n37057 ; n37058
g34623 and n6205 n37058 ; n37059
g34624 and n16699_not n37003 ; n37060
g34625 and pi0681 n37060_not ; n37061
g34626 and n17375 n37054 ; n37062
g34627 and n6194_not n37060 ; n37063
g34628 nor pi0681 n37062 ; n37064
g34629 and n37063_not n37064 ; n37065
g34630 nor n37061 n37065 ; n37066
g34631 and n6205_not n37066 ; n37067
g34632 nor n2603 n37059 ; n37068
g34633 and n37067_not n37068 ; n37069
g34634 nor pi0223 n37051 ; n37070
g34635 and n37069_not n37070 ; n37071
g34636 nor pi0299 n37049 ; n37072
g34637 and n37071_not n37072 ; n37073
g34638 and n17236 n37054 ; n37074
g34639 and n37053 n37074_not ; n37075
g34640 and n16723 n37043 ; n37076
g34641 nor n37075 n37076 ; n37077
g34642 and pi0642 n17237 ; n37078
g34643 and pi0681 n37078_not ; n37079
g34644 and n37077 n37079_not ; n37080
g34645 and pi0947 n37080_not ; n37081
g34646 and n6242 n37075_not ; n37082
g34647 and n37050 n37082 ; n37083
g34648 and n20923_not n37080 ; n37084
g34649 nor pi0947 n37083 ; n37085
g34650 and n37084_not n37085 ; n37086
g34651 nor pi0223 n37081 ; n37087
g34652 and n37086_not n37087 ; n37088
g34653 and n6242_not n37046 ; n37089
g34654 and n6242 n37034 ; n37090
g34655 and pi0223 n37089_not ; n37091
g34656 and n37090_not n37091 ; n37092
g34657 nor n37088 n37092 ; n37093
g34658 and pi0215 n37093_not ; n37094
g34659 and n36931 n37050_not ; n37095
g34660 and pi0947 n37066_not ; n37096
g34661 and n20923 n37058 ; n37097
g34662 and n20923_not n37066 ; n37098
g34663 nor pi0947 n37097 ; n37099
g34664 and n37098_not n37099 ; n37100
g34665 nor pi0223 n37096 ; n37101
g34666 and n37100_not n37101 ; n37102
g34667 and pi0642 n17154_not ; n37103
g34668 nor pi0642 n16702 ; n37104
g34669 nor n37103 n37104 ; n37105
g34670 and pi0681 n37105_not ; n37106
g34671 and n6194_not n37105 ; n37107
g34672 and n17014 n37003_not ; n37108
g34673 nor pi0681 n37108 ; n37109
g34674 and n37107_not n37109 ; n37110
g34675 nor n6242 n37110 ; n37111
g34676 and n37106_not n37111 ; n37112
g34677 and n6191 n37025_not ; n37113
g34678 and n16770_not n37113 ; n37114
g34679 nor n37024 n37114 ; n37115
g34680 and pi0681 n37115 ; n37116
g34681 nor n6194 n37115 ; n37117
g34682 nor n17164 n35894 ; n37118
g34683 and n6194 n37118_not ; n37119
g34684 nor pi0681 n37119 ; n37120
g34685 and n37117_not n37120 ; n37121
g34686 and n6242 n37121_not ; n37122
g34687 and n37116_not n37122 ; n37123
g34688 and pi0223 n37112_not ; n37124
g34689 and n37123_not n37124 ; n37125
g34690 nor n3448 n37102 ; n37126
g34691 and n37125_not n37126 ; n37127
g34692 nor pi0215 n37095 ; n37128
g34693 and n37127_not n37128 ; n37129
g34694 and pi0299 n37094_not ; n37130
g34695 and n37129_not n37130 ; n37131
g34696 and pi0039 n37073_not ; n37132
g34697 and n37131_not n37132 ; n37133
g34698 nor pi0038 n37023 ; n37134
g34699 and n37133_not n37134 ; n37135
g34700 and n2571 n37008_not ; n37136
g34701 and n37135_not n37136 ; n37137
g34702 nor n36886 n37137 ; n37138
g34703 and n17117_not n37138 ; n37139
g34704 nor n37000 n37139 ; n37140
g34705 and pi0785_not n37140 ; n37141
g34706 and pi0609 n37140_not ; n37142
g34707 nor pi0609 n36883 ; n37143
g34708 and pi1155 n37143_not ; n37144
g34709 and n37142_not n37144 ; n37145
g34710 nor pi0609 n37140 ; n37146
g34711 and pi0609 n36883_not ; n37147
g34712 nor pi1155 n37147 ; n37148
g34713 and n37146_not n37148 ; n37149
g34714 nor n37145 n37149 ; n37150
g34715 and pi0785 n37150_not ; n37151
g34716 nor n37141 n37151 ; n37152
g34717 nor pi0781 n37152 ; n37153
g34718 and pi0618 n37152 ; n37154
g34719 nor pi0618 n36883 ; n37155
g34720 and pi1154 n37155_not ; n37156
g34721 and n37154_not n37156 ; n37157
g34722 and pi0618_not n37152 ; n37158
g34723 and pi0618 n36883_not ; n37159
g34724 nor pi1154 n37159 ; n37160
g34725 and n37158_not n37160 ; n37161
g34726 nor n37157 n37161 ; n37162
g34727 and pi0781 n37162_not ; n37163
g34728 nor n37153 n37163 ; n37164
g34729 nor pi0789 n37164 ; n37165
g34730 and pi0619 n37164 ; n37166
g34731 nor pi0619 n36883 ; n37167
g34732 and pi1159 n37167_not ; n37168
g34733 and n37166_not n37168 ; n37169
g34734 and pi0619_not n37164 ; n37170
g34735 and pi0619 n36883_not ; n37171
g34736 nor pi1159 n37171 ; n37172
g34737 and n37170_not n37172 ; n37173
g34738 nor n37169 n37173 ; n37174
g34739 and pi0789 n37174_not ; n37175
g34740 nor n37165 n37175 ; n37176
g34741 and n17969_not n37176 ; n37177
g34742 nor n36999 n37177 ; n37178
g34743 and n17779_not n37178 ; n37179
g34744 and n17779 n36883 ; n37180
g34745 nor n37179 n37180 ; n37181
g34746 nor n20559 n37181 ; n37182
g34747 and pi0630 n36989 ; n37183
g34748 nor n36998 n37183 ; n37184
g34749 and n37182_not n37184 ; n37185
g34750 and pi0787 n37185_not ; n37186
g34751 and pi0628 n36883_not ; n37187
g34752 nor pi0628 n36981 ; n37188
g34753 and n17777 n37187_not ; n37189
g34754 and n37188_not n37189 ; n37190
g34755 and n20570_not n37178 ; n37191
g34756 nor pi0628 n36883 ; n37192
g34757 and pi0628 n36981_not ; n37193
g34758 and n17776 n37192_not ; n37194
g34759 and n37193_not n37194 ; n37195
g34760 nor n37190 n37195 ; n37196
g34761 and n37191_not n37196 ; n37197
g34762 and pi0792 n37197_not ; n37198
g34763 and n16635 n36883_not ; n37199
g34764 nor n36979 n37199 ; n37200
g34765 and n17871 n37200_not ; n37201
g34766 and pi0626_not n36883 ; n37202
g34767 and pi0626 n37176_not ; n37203
g34768 and n16628 n37202_not ; n37204
g34769 and n37203_not n37204 ; n37205
g34770 and pi0626 n36883 ; n37206
g34771 nor pi0626 n37176 ; n37207
g34772 and n16629 n37206_not ; n37208
g34773 and n37207_not n37208 ; n37209
g34774 nor n37201 n37205 ; n37210
g34775 and n37209_not n37210 ; n37211
g34776 and pi0788 n37211_not ; n37212
g34777 and pi0609 n36973 ; n37213
g34778 and n36887_not n37003 ; n37214
g34779 nor pi0642 n17336 ; n37215
g34780 and n36887 n37215_not ; n37216
g34781 and n36562_not n37216 ; n37217
g34782 nor n37214 n37217 ; n37218
g34783 and n36887_not n37004 ; n37219
g34784 and pi0642 n17493 ; n37220
g34785 nor n37215 n37220 ; n37221
g34786 and n16667 n37221_not ; n37222
g34787 and n36887 n37222 ; n37223
g34788 and pi0223 n37219_not ; n37224
g34789 and n37223_not n37224 ; n37225
g34790 and n37218 n37225_not ; n37226
g34791 and n37006 n37226_not ; n37227
g34792 and n37002 n37227_not ; n37228
g34793 and n17618 n36922 ; n37229
g34794 and n17617 n36887_not ; n37230
g34795 and n36728_not n37013 ; n37231
g34796 and n37230_not n37231 ; n37232
g34797 and n37011 n37229_not ; n37233
g34798 and n37232_not n37233 ; n37234
g34799 and n17623 n36922 ; n37235
g34800 and n17622 n36887_not ; n37236
g34801 and pi0223 n37018_not ; n37237
g34802 and n36738_not n37237 ; n37238
g34803 and n37236_not n37238 ; n37239
g34804 and n37017 n37235_not ; n37240
g34805 and n37239_not n37240 ; n37241
g34806 nor pi0039 n37234 ; n37242
g34807 and n37241_not n37242 ; n37243
g34808 nor n36887 n37028 ; n37244
g34809 and n16650_not n37222 ; n37245
g34810 nor n6191 n37245 ; n37246
g34811 and pi0680 n37246_not ; n37247
g34812 and pi0642 n17504_not ; n37248
g34813 and pi0614_not n17343 ; n37249
g34814 nor n37248 n37249 ; n37250
g34815 nor pi0616 n37250 ; n37251
g34816 and n37247 n37251_not ; n37252
g34817 nor n37244 n37252 ; n37253
g34818 nor n37033 n37253 ; n37254
g34819 and n6242 n37254_not ; n37255
g34820 and pi0680_not n37038 ; n37256
g34821 and pi0642 n36588_not ; n37257
g34822 and n6191_not n17325 ; n37258
g34823 and pi0680 n17329_not ; n37259
g34824 and n37257_not n37259 ; n37260
g34825 and n37258_not n37260 ; n37261
g34826 and pi0681 n37261_not ; n37262
g34827 and n37256_not n37262 ; n37263
g34828 nor n37044 n37263 ; n37264
g34829 nor n6242 n37264 ; n37265
g34830 and pi0223 n37265_not ; n37266
g34831 and n37255_not n37266 ; n37267
g34832 nor pi0680 n37050 ; n37268
g34833 nor n17336 n37248 ; n37269
g34834 and n35897 n37269_not ; n37270
g34835 and pi0680 n37270_not ; n37271
g34836 and pi0642 n17548_not ; n37272
g34837 and n6191 n37272_not ; n37273
g34838 and n17455_not n37273 ; n37274
g34839 and n37271 n37274_not ; n37275
g34840 nor n37268 n37275 ; n37276
g34841 and pi0681 n37276_not ; n37277
g34842 and n37082 n37277_not ; n37278
g34843 nor n36887 n37079 ; n37279
g34844 nor pi0642 n6191 ; n37280
g34845 and n17450_not n37280 ; n37281
g34846 and n17454 n17559 ; n37282
g34847 and n17167 n37282_not ; n37283
g34848 and pi0642 n36607 ; n37284
g34849 and pi0680 n37281_not ; n37285
g34850 and n37284_not n37285 ; n37286
g34851 and n37283_not n37286 ; n37287
g34852 nor n37279 n37287 ; n37288
g34853 and n6242_not n37077 ; n37289
g34854 and n37288_not n37289 ; n37290
g34855 nor pi0223 n37278 ; n37291
g34856 and n37290_not n37291 ; n37292
g34857 and pi0215 n37292_not ; n37293
g34858 and n37267_not n37293 ; n37294
g34859 nor n36887 n37116 ; n37295
g34860 nor n17359 n37248 ; n37296
g34861 and n6191 n37296_not ; n37297
g34862 and n37247 n37297_not ; n37298
g34863 nor n37295 n37298 ; n37299
g34864 and n37122 n37299_not ; n37300
g34865 nor n36887 n37106 ; n37301
g34866 and pi0642 n36638_not ; n37302
g34867 and n17167 n36631_not ; n37303
g34868 and n36633 n37280 ; n37304
g34869 and pi0680 n37302_not ; n37305
g34870 and n37303_not n37305 ; n37306
g34871 and n37304_not n37306 ; n37307
g34872 nor n37301 n37307 ; n37308
g34873 and n37111 n37308_not ; n37309
g34874 and pi0223 n37309_not ; n37310
g34875 and n37300_not n37310 ; n37311
g34876 nor pi0642 n17414 ; n37312
g34877 and n37273 n37312_not ; n37313
g34878 and n37271 n37313_not ; n37314
g34879 nor n37268 n37314 ; n37315
g34880 and pi0681 n37315_not ; n37316
g34881 nor n37056 n37316 ; n37317
g34882 and n6242 n37317_not ; n37318
g34883 nor n36887 n37061 ; n37319
g34884 and pi0642 n17578 ; n37320
g34885 and n17422_not n37280 ; n37321
g34886 and pi0680 n37320_not ; n37322
g34887 and n17430_not n37322 ; n37323
g34888 and n37321_not n37323 ; n37324
g34889 nor n37319 n37324 ; n37325
g34890 nor n37065 n37325 ; n37326
g34891 nor n6242 n37326 ; n37327
g34892 nor pi0223 n37318 ; n37328
g34893 and n37327_not n37328 ; n37329
g34894 nor n3448 n37311 ; n37330
g34895 and n37329_not n37330 ; n37331
g34896 and n16653 n37218_not ; n37332
g34897 and pi0223_not n37332 ; n37333
g34898 and n36931 n37225_not ; n37334
g34899 and n37333_not n37334 ; n37335
g34900 nor pi0215 n37335 ; n37336
g34901 and n37331_not n37336 ; n37337
g34902 and pi0299 n37294_not ; n37338
g34903 and n37337_not n37338 ; n37339
g34904 and n6205 n37254 ; n37340
g34905 and n6205_not n37264 ; n37341
g34906 and pi0223 n37341_not ; n37342
g34907 and n37340_not n37342 ; n37343
g34908 and n2603 n37332_not ; n37344
g34909 and n6205_not n37326 ; n37345
g34910 and n6205 n37317 ; n37346
g34911 nor n2603 n37345 ; n37347
g34912 and n37346_not n37347 ; n37348
g34913 nor pi0223 n37344 ; n37349
g34914 and n37348_not n37349 ; n37350
g34915 nor pi0299 n37343 ; n37351
g34916 and n37350_not n37351 ; n37352
g34917 and pi0039 n37352_not ; n37353
g34918 and n37339_not n37353 ; n37354
g34919 nor pi0038 n37243 ; n37355
g34920 and n37354_not n37355 ; n37356
g34921 and n2571 n37228_not ; n37357
g34922 and n37356_not n37357 ; n37358
g34923 nor n36886 n37358 ; n37359
g34924 and pi0625_not n37359 ; n37360
g34925 and pi0625 n37138 ; n37361
g34926 nor pi1153 n37361 ; n37362
g34927 and n37360_not n37362 ; n37363
g34928 nor pi0608 n37363 ; n37364
g34929 and n36966_not n37364 ; n37365
g34930 and pi0625_not n37138 ; n37366
g34931 and pi0625 n37359 ; n37367
g34932 and pi1153 n37366_not ; n37368
g34933 and n37367_not n37368 ; n37369
g34934 and pi0608 n37369_not ; n37370
g34935 and n36970_not n37370 ; n37371
g34936 nor n37365 n37371 ; n37372
g34937 and pi0778 n37372_not ; n37373
g34938 and pi0778_not n37359 ; n37374
g34939 nor n37373 n37374 ; n37375
g34940 nor pi0609 n37375 ; n37376
g34941 nor pi1155 n37213 ; n37377
g34942 and n37376_not n37377 ; n37378
g34943 nor pi0660 n37145 ; n37379
g34944 and n37378_not n37379 ; n37380
g34945 and pi0609_not n36973 ; n37381
g34946 and pi0609 n37375_not ; n37382
g34947 and pi1155 n37381_not ; n37383
g34948 and n37382_not n37383 ; n37384
g34949 and pi0660 n37149_not ; n37385
g34950 and n37384_not n37385 ; n37386
g34951 nor n37380 n37386 ; n37387
g34952 and pi0785 n37387_not ; n37388
g34953 nor pi0785 n37375 ; n37389
g34954 nor n37388 n37389 ; n37390
g34955 nor pi0618 n37390 ; n37391
g34956 and pi0618 n36975_not ; n37392
g34957 nor pi1154 n37392 ; n37393
g34958 and n37391_not n37393 ; n37394
g34959 nor pi0627 n37157 ; n37395
g34960 and n37394_not n37395 ; n37396
g34961 and pi0618 n37390_not ; n37397
g34962 nor pi0618 n36975 ; n37398
g34963 and pi1154 n37398_not ; n37399
g34964 and n37397_not n37399 ; n37400
g34965 and pi0627 n37161_not ; n37401
g34966 and n37400_not n37401 ; n37402
g34967 nor n37396 n37402 ; n37403
g34968 and pi0781 n37403_not ; n37404
g34969 nor pi0781 n37390 ; n37405
g34970 nor n37404 n37405 ; n37406
g34971 and pi0789_not n37406 ; n37407
g34972 nor pi0619 n37406 ; n37408
g34973 and pi0619 n36978 ; n37409
g34974 nor pi1159 n37409 ; n37410
g34975 and n37408_not n37410 ; n37411
g34976 nor pi0648 n37169 ; n37412
g34977 and n37411_not n37412 ; n37413
g34978 and pi0619_not n36978 ; n37414
g34979 and pi0619 n37406_not ; n37415
g34980 and pi1159 n37414_not ; n37416
g34981 and n37415_not n37416 ; n37417
g34982 and pi0648 n37173_not ; n37418
g34983 and n37417_not n37418 ; n37419
g34984 and pi0789 n37413_not ; n37420
g34985 and n37419_not n37420 ; n37421
g34986 and n17970 n37407_not ; n37422
g34987 and n37421_not n37422 ; n37423
g34988 nor n37212 n37423 ; n37424
g34989 nor n37198 n37424 ; n37425
g34990 and n20364 n37197 ; n37426
g34991 nor n20206 n37426 ; n37427
g34992 and n37425_not n37427 ; n37428
g34993 nor n37186 n37428 ; n37429
g34994 and pi0644 n37429 ; n37430
g34995 and pi0715 n36997_not ; n37431
g34996 and n37430_not n37431 ; n37432
g34997 and n17804 n36883_not ; n37433
g34998 and n17804_not n37181 ; n37434
g34999 nor n37433 n37434 ; n37435
g35000 and pi0644 n37435_not ; n37436
g35001 nor pi0644 n36883 ; n37437
g35002 nor pi0715 n37437 ; n37438
g35003 and n37436_not n37438 ; n37439
g35004 and pi1160 n37439_not ; n37440
g35005 and n37432_not n37440 ; n37441
g35006 and pi0644 n36996 ; n37442
g35007 and pi0644_not n37429 ; n37443
g35008 nor pi0715 n37442 ; n37444
g35009 and n37443_not n37444 ; n37445
g35010 nor pi0644 n37435 ; n37446
g35011 and pi0644 n36883_not ; n37447
g35012 and pi0715 n37447_not ; n37448
g35013 and n37446_not n37448 ; n37449
g35014 nor pi1160 n37449 ; n37450
g35015 and n37445_not n37450 ; n37451
g35016 nor n37441 n37451 ; n37452
g35017 and pi0790 n37452_not ; n37453
g35018 and pi0790_not n37429 ; n37454
g35019 nor n37453 n37454 ; n37455
g35020 nor po1038 n37455 ; n37456
g35021 and pi0223_not po1038 ; n37457
g35022 nor n37456 n37457 ; po0380
g35023 and pi0224 n36258_not ; n37459
g35024 nor n19149 n37459 ; n37460
g35025 and pi0224 n2571_not ; n37461
g35026 and pi0224 n16641_not ; n37462
g35027 and pi0038 n37462_not ; n37463
g35028 and pi0662 n16646 ; n37464
g35029 and n37463 n37464_not ; n37465
g35030 and pi0662 pi0680 ; n37466
g35031 and n16918 n37466_not ; n37467
g35032 nor pi0224 n16918 ; n37468
g35033 and pi0224 n16935 ; n37469
g35034 nor pi0299 n37469 ; n37470
g35035 and n37467_not n37470 ; n37471
g35036 and n37468_not n37471 ; n37472
g35037 and pi0224 n16944 ; n37473
g35038 and n16923 n37466_not ; n37474
g35039 nor pi0224 n16923 ; n37475
g35040 and pi0299 n37473_not ; n37476
g35041 and n37474_not n37476 ; n37477
g35042 and n37475_not n37477 ; n37478
g35043 nor pi0039 n37472 ; n37479
g35044 and n37478_not n37479 ; n37480
g35045 and pi0662 n16655 ; n37481
g35046 nor n6193 n36283 ; n37482
g35047 and n17018 n37482_not ; n37483
g35048 and n6205_not n37483 ; n37484
g35049 and pi0662 n16786_not ; n37485
g35050 nor pi0662 n17011 ; n37486
g35051 nor n37485 n37486 ; n37487
g35052 and n6205 n37487 ; n37488
g35053 and pi0224 n37484_not ; n37489
g35054 and n37488_not n37489 ; n37490
g35055 and pi0662 n16703 ; n37491
g35056 nor n6205 n37491 ; n37492
g35057 and n16690_not n37466 ; n37493
g35058 and n6205 n37493_not ; n37494
g35059 and n5810 n37492_not ; n37495
g35060 and n37494_not n37495 ; n37496
g35061 nor pi0223 n37481 ; n37497
g35062 and n37496_not n37497 ; n37498
g35063 and n37490_not n37498 ; n37499
g35064 and pi0224_not pi0662 ; n37500
g35065 and n16729 n37500 ; n37501
g35066 nor pi0662 n16990 ; n37502
g35067 and pi0662 n36319_not ; n37503
g35068 nor n37502 n37503 ; n37504
g35069 and n6205 n37504 ; n37505
g35070 nor pi0662 n16970 ; n37506
g35071 and pi0662 n16818_not ; n37507
g35072 nor n37506 n37507 ; n37508
g35073 and n6205_not n37508 ; n37509
g35074 and pi0224 n37505_not ; n37510
g35075 and n37509_not n37510 ; n37511
g35076 and pi0223 n37501_not ; n37512
g35077 and n37511_not n37512 ; n37513
g35078 nor pi0299 n37513 ; n37514
g35079 and n37499_not n37514 ; n37515
g35080 and pi0224 n16653_not ; n37516
g35081 and n3448 n37516_not ; n37517
g35082 and n16658 n37466 ; n37518
g35083 and n37517 n37518_not ; n37519
g35084 and n6242_not n37483 ; n37520
g35085 and n6242 n37487 ; n37521
g35086 and pi0224 n37520_not ; n37522
g35087 and n37521_not n37522 ; n37523
g35088 nor n6242 n37491 ; n37524
g35089 and n6242 n37493_not ; n37525
g35090 nor pi0224 n37524 ; n37526
g35091 and n37525_not n37526 ; n37527
g35092 nor n3448 n37527 ; n37528
g35093 and n37523_not n37528 ; n37529
g35094 nor n37519 n37529 ; n37530
g35095 nor pi0215 n37530 ; n37531
g35096 and n16744 n37500 ; n37532
g35097 and n6242 n37504 ; n37533
g35098 and n6242_not n37508 ; n37534
g35099 and pi0224 n37533_not ; n37535
g35100 and n37534_not n37535 ; n37536
g35101 and pi0215 n37532_not ; n37537
g35102 and n37536_not n37537 ; n37538
g35103 and pi0299 n37538_not ; n37539
g35104 and n37531_not n37539 ; n37540
g35105 and pi0039 n37515_not ; n37541
g35106 and n37540_not n37541 ; n37542
g35107 nor n37480 n37542 ; n37543
g35108 nor pi0038 n37543 ; n37544
g35109 and n2571 n37465_not ; n37545
g35110 and n37544_not n37545 ; n37546
g35111 nor n37461 n37546 ; n37547
g35112 nor pi0778 n37547 ; n37548
g35113 and pi0625 n37547 ; n37549
g35114 nor pi0625 n37459 ; n37550
g35115 and pi1153 n37550_not ; n37551
g35116 and n37549_not n37551 ; n37552
g35117 and pi0625_not n37547 ; n37553
g35118 and pi0625 n37459_not ; n37554
g35119 nor pi1153 n37554 ; n37555
g35120 and n37553_not n37555 ; n37556
g35121 nor n37552 n37556 ; n37557
g35122 and pi0778 n37557_not ; n37558
g35123 nor n37548 n37558 ; n37559
g35124 nor n17075 n37559 ; n37560
g35125 and n17075 n37459 ; n37561
g35126 nor n37560 n37561 ; n37562
g35127 nor n16639 n37562 ; n37563
g35128 and n16639 n37459 ; n37564
g35129 nor n37563 n37564 ; n37565
g35130 and n16635_not n37565 ; n37566
g35131 and n16631_not n37566 ; n37567
g35132 nor n37460 n37567 ; n37568
g35133 nor n19142 n37568 ; n37569
g35134 and n17856 n37459_not ; n37570
g35135 nor n37569 n37570 ; n37571
g35136 and pi0787_not n37571 ; n37572
g35137 nor pi0647 n37571 ; n37573
g35138 and pi0647 n37459_not ; n37574
g35139 nor pi1157 n37574 ; n37575
g35140 and n37573_not n37575 ; n37576
g35141 and pi0647 n37571_not ; n37577
g35142 nor pi0647 n37459 ; n37578
g35143 and pi1157 n37578_not ; n37579
g35144 and n37577_not n37579 ; n37580
g35145 nor n37576 n37580 ; n37581
g35146 and pi0787 n37581_not ; n37582
g35147 nor n37572 n37582 ; n37583
g35148 and pi0644_not n37583 ; n37584
g35149 and pi0628 n37459_not ; n37585
g35150 nor pi0628 n37568 ; n37586
g35151 and n17777 n37585_not ; n37587
g35152 and n37586_not n37587 ; n37588
g35153 and n17969 n37459_not ; n37589
g35154 and pi0614 n17280 ; n37590
g35155 and n37463 n37590_not ; n37591
g35156 and pi0614 n17226 ; n37592
g35157 and pi0224_not n37592 ; n37593
g35158 and pi0614_not n17226 ; n37594
g35159 and pi0224 n37594_not ; n37595
g35160 and n17137 n37595 ; n37596
g35161 nor pi0299 n37593 ; n37597
g35162 and n37596_not n37597 ; n37598
g35163 and pi0614 n17231 ; n37599
g35164 and pi0224 n17122 ; n37600
g35165 and n37599 n37600_not ; n37601
g35166 and pi0224 n16941_not ; n37602
g35167 nor n37601 n37602 ; n37603
g35168 and pi0299 n37603 ; n37604
g35169 nor pi0039 n37598 ; n37605
g35170 and n37604_not n37605 ; n37606
g35171 and pi0614 n36411_not ; n37607
g35172 and pi0224_not n37607 ; n37608
g35173 and n16743_not n37608 ; n37609
g35174 and pi0614 n17183_not ; n37610
g35175 nor n36026 n37610 ; n37611
g35176 nor pi0680 n37611 ; n37612
g35177 and pi0680 n17187_not ; n37613
g35178 and n36028_not n37613 ; n37614
g35179 nor n37612 n37614 ; n37615
g35180 and n16657 n37615_not ; n37616
g35181 nor n16657 n37611 ; n37617
g35182 nor n37616 n37617 ; n37618
g35183 and n6242_not n37618 ; n37619
g35184 and pi0614 n17168 ; n37620
g35185 and n16653 n37620_not ; n37621
g35186 nor n6192 n37621 ; n37622
g35187 nor n16802 n37622 ; n37623
g35188 nor n16657 n37623 ; n37624
g35189 nor pi0680 n37623 ; n37625
g35190 and pi0680 n37620 ; n37626
g35191 nor n16973 n37626 ; n37627
g35192 and n37625_not n37627 ; n37628
g35193 and n16657 n37628_not ; n37629
g35194 nor n37624 n37629 ; n37630
g35195 and n6242 n37630 ; n37631
g35196 and pi0224 n37619_not ; n37632
g35197 and n37631_not n37632 ; n37633
g35198 nor n37609 n37633 ; n37634
g35199 and pi0215 n37634_not ; n37635
g35200 and n16999 n17168 ; n37636
g35201 and n37517 n37636_not ; n37637
g35202 and pi0614 n17154_not ; n37638
g35203 and pi0614_not pi0616 ; n37639
g35204 and n16699 n37639 ; n37640
g35205 and n6197_not n16772 ; n37641
g35206 and n6191 n16697_not ; n37642
g35207 and n37641_not n37642 ; n37643
g35208 nor n37638 n37640 ; n37644
g35209 and n37643_not n37644 ; n37645
g35210 nor n16657 n37645 ; n37646
g35211 nor pi0680 n37645 ; n37647
g35212 and pi0614 n17375 ; n37648
g35213 and pi0680 n37648_not ; n37649
g35214 and n16681 n37649 ; n37650
g35215 nor n37626 n37650 ; n37651
g35216 and n37647_not n37651 ; n37652
g35217 and n16657 n37652_not ; n37653
g35218 nor n37646 n37653 ; n37654
g35219 and n6242_not n37654 ; n37655
g35220 nor n16775 n37622 ; n37656
g35221 nor n16657 n37656 ; n37657
g35222 nor pi0680 n37656 ; n37658
g35223 nor n16995 n37626 ; n37659
g35224 and n37658_not n37659 ; n37660
g35225 and n16657 n37660_not ; n37661
g35226 nor n37657 n37661 ; n37662
g35227 and n6242 n37662 ; n37663
g35228 and pi0224 n37655_not ; n37664
g35229 and n37663_not n37664 ; n37665
g35230 and n16699_not n37620 ; n37666
g35231 nor pi0680 n37666 ; n37667
g35232 nor n37649 n37667 ; n37668
g35233 and n16657 n37668_not ; n37669
g35234 nor n16657 n37666 ; n37670
g35235 nor n37669 n37670 ; n37671
g35236 nor n6242 n37671 ; n37672
g35237 and pi0614 n36463_not ; n37673
g35238 and n6242 n37673_not ; n37674
g35239 nor pi0224 n37674 ; n37675
g35240 and n37672_not n37675 ; n37676
g35241 nor n3448 n37676 ; n37677
g35242 and n37665_not n37677 ; n37678
g35243 nor pi0215 n37637 ; n37679
g35244 and n37678_not n37679 ; n37680
g35245 and pi0299 n37635_not ; n37681
g35246 and n37680_not n37681 ; n37682
g35247 and n16724_not n37608 ; n37683
g35248 and n6205_not n37618 ; n37684
g35249 and n6205 n37630 ; n37685
g35250 and pi0224 n37684_not ; n37686
g35251 and n37685_not n37686 ; n37687
g35252 and pi0223 n37683_not ; n37688
g35253 and n37687_not n37688 ; n37689
g35254 and pi0614 n17268 ; n37690
g35255 and n6205 n37673_not ; n37691
g35256 nor n6205 n37671 ; n37692
g35257 and n5810 n37691_not ; n37693
g35258 and n37692_not n37693 ; n37694
g35259 and n6205_not n37654 ; n37695
g35260 and n6205 n37662 ; n37696
g35261 and pi0224 n37695_not ; n37697
g35262 and n37696_not n37697 ; n37698
g35263 nor pi0223 n37690 ; n37699
g35264 and n37694_not n37699 ; n37700
g35265 and n37698_not n37700 ; n37701
g35266 nor n37689 n37701 ; n37702
g35267 nor pi0299 n37702 ; n37703
g35268 and pi0039 n37682_not ; n37704
g35269 and n37703_not n37704 ; n37705
g35270 nor pi0038 n37606 ; n37706
g35271 and n37705_not n37706 ; n37707
g35272 and n2571 n37591_not ; n37708
g35273 and n37707_not n37708 ; n37709
g35274 nor n37461 n37709 ; n37710
g35275 nor n17117 n37710 ; n37711
g35276 and n17117 n37459 ; n37712
g35277 nor n37711 n37712 ; n37713
g35278 nor pi0785 n37713 ; n37714
g35279 and pi0609 n37713 ; n37715
g35280 nor pi0609 n37459 ; n37716
g35281 and pi1155 n37716_not ; n37717
g35282 and n37715_not n37717 ; n37718
g35283 and pi0609_not n37713 ; n37719
g35284 and pi0609 n37459_not ; n37720
g35285 nor pi1155 n37720 ; n37721
g35286 and n37719_not n37721 ; n37722
g35287 nor n37718 n37722 ; n37723
g35288 and pi0785 n37723_not ; n37724
g35289 nor n37714 n37724 ; n37725
g35290 nor pi0781 n37725 ; n37726
g35291 and pi0618 n37725 ; n37727
g35292 nor pi0618 n37459 ; n37728
g35293 and pi1154 n37728_not ; n37729
g35294 and n37727_not n37729 ; n37730
g35295 and pi0618_not n37725 ; n37731
g35296 and pi0618 n37459_not ; n37732
g35297 nor pi1154 n37732 ; n37733
g35298 and n37731_not n37733 ; n37734
g35299 nor n37730 n37734 ; n37735
g35300 and pi0781 n37735_not ; n37736
g35301 nor n37726 n37736 ; n37737
g35302 nor pi0789 n37737 ; n37738
g35303 and pi0619 n37737 ; n37739
g35304 nor pi0619 n37459 ; n37740
g35305 and pi1159 n37740_not ; n37741
g35306 and n37739_not n37741 ; n37742
g35307 and pi0619_not n37737 ; n37743
g35308 and pi0619 n37459_not ; n37744
g35309 nor pi1159 n37744 ; n37745
g35310 and n37743_not n37745 ; n37746
g35311 nor n37742 n37746 ; n37747
g35312 and pi0789 n37747_not ; n37748
g35313 nor n37738 n37748 ; n37749
g35314 and n17969_not n37749 ; n37750
g35315 nor n37589 n37750 ; n37751
g35316 and n20570_not n37751 ; n37752
g35317 nor pi0628 n37459 ; n37753
g35318 and pi0628 n37568_not ; n37754
g35319 and n17776 n37753_not ; n37755
g35320 and n37754_not n37755 ; n37756
g35321 nor n37588 n37756 ; n37757
g35322 and n37752_not n37757 ; n37758
g35323 and pi0792 n37758_not ; n37759
g35324 and pi0609 n37559 ; n37760
g35325 and pi0662 n17355 ; n37761
g35326 and n16641 n37761 ; n37762
g35327 and n37591 n37762_not ; n37763
g35328 and n17617 n37466 ; n37764
g35329 nor n37592 n37764 ; n37765
g35330 nor pi0224 n37765 ; n37766
g35331 and n17617 n37466_not ; n37767
g35332 and n36728_not n37595 ; n37768
g35333 and n37767_not n37768 ; n37769
g35334 nor n37766 n37769 ; n37770
g35335 nor pi0299 n37770 ; n37771
g35336 and n37466_not n37603 ; n37772
g35337 and pi0614_not n17231 ; n37773
g35338 nor n36738 n37773 ; n37774
g35339 and pi0224 n37774_not ; n37775
g35340 nor pi0224 n17622 ; n37776
g35341 and n37599_not n37776 ; n37777
g35342 nor n37775 n37777 ; n37778
g35343 and n37466 n37778_not ; n37779
g35344 and pi0299 n37772_not ; n37780
g35345 and n37779_not n37780 ; n37781
g35346 nor n37771 n37781 ; n37782
g35347 nor pi0039 n37782 ; n37783
g35348 and n17407 n37466 ; n37784
g35349 nor n37636 n37784 ; n37785
g35350 nor pi0224 n37785 ; n37786
g35351 and pi0222_not n37786 ; n37787
g35352 and n17407_not n37639 ; n37788
g35353 nor n36620 n37788 ; n37789
g35354 and pi0680 n37789_not ; n37790
g35355 nor n36675 n37636 ; n37791
g35356 nor n37790 n37791 ; n37792
g35357 and pi0662 n37792_not ; n37793
g35358 nor pi0662 n37673 ; n37794
g35359 nor n37793 n37794 ; n37795
g35360 and n6205 n37795_not ; n37796
g35361 nor pi0662 n16656 ; n37797
g35362 and n37666_not n37797 ; n37798
g35363 and pi0614_not n17434 ; n37799
g35364 and pi0614 n17578_not ; n37800
g35365 and pi0680 n37800_not ; n37801
g35366 and n37799_not n37801 ; n37802
g35367 nor n37667 n37802 ; n37803
g35368 and pi0662 n37803_not ; n37804
g35369 nor n37669 n37798 ; n37805
g35370 and n37804_not n37805 ; n37806
g35371 nor n6205 n37806 ; n37807
g35372 and n5810 n37796_not ; n37808
g35373 and n37807_not n37808 ; n37809
g35374 and n37656_not n37797 ; n37810
g35375 nor pi0614 n24055 ; n37811
g35376 and pi0614 n36562_not ; n37812
g35377 nor n37811 n37812 ; n37813
g35378 and n16650_not n37813 ; n37814
g35379 and pi0616 n37814_not ; n37815
g35380 and pi0614 n17504_not ; n37816
g35381 nor n17361 n37816 ; n37817
g35382 nor pi0616 n37817 ; n37818
g35383 nor n37815 n37818 ; n37819
g35384 and pi0680 n37819_not ; n37820
g35385 nor n37658 n37820 ; n37821
g35386 and pi0662 n37821_not ; n37822
g35387 nor n37661 n37810 ; n37823
g35388 and n37822_not n37823 ; n37824
g35389 and n6205 n37824 ; n37825
g35390 and n37645_not n37797 ; n37826
g35391 and pi0614 n36638_not ; n37827
g35392 and n36633 n37639 ; n37828
g35393 nor n37827 n37828 ; n37829
g35394 and n36636_not n37829 ; n37830
g35395 and pi0680 n37830_not ; n37831
g35396 nor n37647 n37831 ; n37832
g35397 and pi0662 n37832_not ; n37833
g35398 nor n37653 n37826 ; n37834
g35399 and n37833_not n37834 ; n37835
g35400 and n6205_not n37835 ; n37836
g35401 and pi0224 n37836_not ; n37837
g35402 and n37825_not n37837 ; n37838
g35403 nor pi0223 n37787 ; n37839
g35404 and n37809_not n37839 ; n37840
g35405 and n37838_not n37840 ; n37841
g35406 and pi0680 n17445_not ; n37842
g35407 nor n37636 n37842 ; n37843
g35408 nor n37790 n37843 ; n37844
g35409 and pi0662 n37844_not ; n37845
g35410 nor pi0662 n37607 ; n37846
g35411 nor n37845 n37846 ; n37847
g35412 nor pi0224 n37847 ; n37848
g35413 and n37623_not n37797 ; n37849
g35414 nor n17345 n37816 ; n37850
g35415 nor pi0616 n37850 ; n37851
g35416 nor n37815 n37851 ; n37852
g35417 and pi0680 n37852_not ; n37853
g35418 nor n37625 n37853 ; n37854
g35419 and pi0662 n37854_not ; n37855
g35420 nor n37629 n37849 ; n37856
g35421 and n37855_not n37856 ; n37857
g35422 and pi0224 n37857 ; n37858
g35423 and n6205 n37848_not ; n37859
g35424 and n37858_not n37859 ; n37860
g35425 and n37611_not n37797 ; n37861
g35426 and pi0614 n36588_not ; n37862
g35427 and n17330 n37862_not ; n37863
g35428 and pi0680 n37863_not ; n37864
g35429 nor n37612 n37864 ; n37865
g35430 and pi0662 n37865_not ; n37866
g35431 nor n37616 n37861 ; n37867
g35432 and n37866_not n37867 ; n37868
g35433 and pi0224 n37868 ; n37869
g35434 and n16723_not n37607 ; n37870
g35435 nor pi0662 n37870 ; n37871
g35436 and pi0614 pi0680_not ; n37872
g35437 and n17237 n37872 ; n37873
g35438 and pi0614 n36607 ; n37874
g35439 and pi0614_not n17451 ; n37875
g35440 and pi0680 n37874_not ; n37876
g35441 and n37875_not n37876 ; n37877
g35442 and n17457_not n37877 ; n37878
g35443 and pi0662 n37873_not ; n37879
g35444 and n37878_not n37879 ; n37880
g35445 nor n37871 n37880 ; n37881
g35446 nor pi0224 n37881 ; n37882
g35447 nor n6205 n37882 ; n37883
g35448 and n37869_not n37883 ; n37884
g35449 and pi0223 n37884_not ; n37885
g35450 and n37860_not n37885 ; n37886
g35451 nor n37841 n37886 ; n37887
g35452 nor pi0299 n37887 ; n37888
g35453 nor n6242 n37868 ; n37889
g35454 and n6242 n37857_not ; n37890
g35455 and pi0224 n37889_not ; n37891
g35456 and n37890_not n37891 ; n37892
g35457 and n6242 n37847 ; n37893
g35458 and n6242_not n37881 ; n37894
g35459 nor pi0224 n37894 ; n37895
g35460 and n37893_not n37895 ; n37896
g35461 and pi0215 n37896_not ; n37897
g35462 and n37892_not n37897 ; n37898
g35463 and n37466 n37813 ; n37899
g35464 nor n37466 n37620 ; n37900
g35465 and n16667 n37900 ; n37901
g35466 and pi0224 n37901_not ; n37902
g35467 and n37899_not n37902 ; n37903
g35468 and n37517 n37903_not ; n37904
g35469 and n37786_not n37904 ; n37905
g35470 nor pi0224 n37795 ; n37906
g35471 and pi0224 n37824 ; n37907
g35472 and n6242 n37906_not ; n37908
g35473 and n37907_not n37908 ; n37909
g35474 nor pi0224 n37806 ; n37910
g35475 and pi0224 n37835 ; n37911
g35476 nor n6242 n37910 ; n37912
g35477 and n37911_not n37912 ; n37913
g35478 nor n3448 n37909 ; n37914
g35479 and n37913_not n37914 ; n37915
g35480 nor pi0215 n37905 ; n37916
g35481 and n37915_not n37916 ; n37917
g35482 and pi0299 n37898_not ; n37918
g35483 and n37917_not n37918 ; n37919
g35484 and pi0039 n37888_not ; n37920
g35485 and n37919_not n37920 ; n37921
g35486 nor pi0038 n37783 ; n37922
g35487 and n37921_not n37922 ; n37923
g35488 and n2571 n37763_not ; n37924
g35489 and n37923_not n37924 ; n37925
g35490 nor n37461 n37925 ; n37926
g35491 and pi0625_not n37926 ; n37927
g35492 and pi0625 n37710 ; n37928
g35493 nor pi1153 n37928 ; n37929
g35494 and n37927_not n37929 ; n37930
g35495 nor pi0608 n37552 ; n37931
g35496 and n37930_not n37931 ; n37932
g35497 and pi0625_not n37710 ; n37933
g35498 and pi0625 n37926 ; n37934
g35499 and pi1153 n37933_not ; n37935
g35500 and n37934_not n37935 ; n37936
g35501 and pi0608 n37556_not ; n37937
g35502 and n37936_not n37937 ; n37938
g35503 nor n37932 n37938 ; n37939
g35504 and pi0778 n37939_not ; n37940
g35505 and pi0778_not n37926 ; n37941
g35506 nor n37940 n37941 ; n37942
g35507 nor pi0609 n37942 ; n37943
g35508 nor pi1155 n37760 ; n37944
g35509 and n37943_not n37944 ; n37945
g35510 nor pi0660 n37718 ; n37946
g35511 and n37945_not n37946 ; n37947
g35512 and pi0609_not n37559 ; n37948
g35513 and pi0609 n37942_not ; n37949
g35514 and pi1155 n37948_not ; n37950
g35515 and n37949_not n37950 ; n37951
g35516 and pi0660 n37722_not ; n37952
g35517 and n37951_not n37952 ; n37953
g35518 nor n37947 n37953 ; n37954
g35519 and pi0785 n37954_not ; n37955
g35520 nor pi0785 n37942 ; n37956
g35521 nor n37955 n37956 ; n37957
g35522 nor pi0618 n37957 ; n37958
g35523 and pi0618 n37562 ; n37959
g35524 nor pi1154 n37959 ; n37960
g35525 and n37958_not n37960 ; n37961
g35526 nor pi0627 n37730 ; n37962
g35527 and n37961_not n37962 ; n37963
g35528 and pi0618_not n37562 ; n37964
g35529 and pi0618 n37957_not ; n37965
g35530 and pi1154 n37964_not ; n37966
g35531 and n37965_not n37966 ; n37967
g35532 and pi0627 n37734_not ; n37968
g35533 and n37967_not n37968 ; n37969
g35534 nor n37963 n37969 ; n37970
g35535 and pi0781 n37970_not ; n37971
g35536 nor pi0781 n37957 ; n37972
g35537 nor n37971 n37972 ; n37973
g35538 and pi0789_not n37973 ; n37974
g35539 nor pi0619 n37973 ; n37975
g35540 and pi0619 n37565 ; n37976
g35541 nor pi1159 n37976 ; n37977
g35542 and n37975_not n37977 ; n37978
g35543 nor pi0648 n37742 ; n37979
g35544 and n37978_not n37979 ; n37980
g35545 and pi0619 n37973_not ; n37981
g35546 and pi0619_not n37565 ; n37982
g35547 and pi1159 n37982_not ; n37983
g35548 and n37981_not n37983 ; n37984
g35549 and pi0648 n37746_not ; n37985
g35550 and n37984_not n37985 ; n37986
g35551 and pi0789 n37980_not ; n37987
g35552 and n37986_not n37987 ; n37988
g35553 and n17970 n37974_not ; n37989
g35554 and n37988_not n37989 ; n37990
g35555 and n16635 n37459_not ; n37991
g35556 nor n37566 n37991 ; n37992
g35557 and n17871 n37992_not ; n37993
g35558 and pi0626_not n37459 ; n37994
g35559 and pi0626 n37749_not ; n37995
g35560 and n16628 n37994_not ; n37996
g35561 and n37995_not n37996 ; n37997
g35562 and pi0626 n37459 ; n37998
g35563 nor pi0626 n37749 ; n37999
g35564 and n16629 n37998_not ; n38000
g35565 and n37999_not n38000 ; n38001
g35566 nor n37993 n37997 ; n38002
g35567 and n38001_not n38002 ; n38003
g35568 and pi0788 n38003_not ; n38004
g35569 nor n20364 n38004 ; n38005
g35570 and n37990_not n38005 ; n38006
g35571 nor n37759 n38006 ; n38007
g35572 nor n20206 n38007 ; n38008
g35573 and pi0630_not n37580 ; n38009
g35574 and n17779_not n37751 ; n38010
g35575 and n17779 n37459 ; n38011
g35576 nor n38010 n38011 ; n38012
g35577 nor n20559 n38012 ; n38013
g35578 and pi0630 n37576 ; n38014
g35579 nor n38009 n38014 ; n38015
g35580 and n38013_not n38015 ; n38016
g35581 and pi0787 n38016_not ; n38017
g35582 nor n38008 n38017 ; n38018
g35583 and pi0644 n38018 ; n38019
g35584 and pi0715 n37584_not ; n38020
g35585 and n38019_not n38020 ; n38021
g35586 and n17804 n37459_not ; n38022
g35587 and n17804_not n38012 ; n38023
g35588 nor n38022 n38023 ; n38024
g35589 and pi0644 n38024_not ; n38025
g35590 nor pi0644 n37459 ; n38026
g35591 nor pi0715 n38026 ; n38027
g35592 and n38025_not n38027 ; n38028
g35593 and pi1160 n38028_not ; n38029
g35594 and n38021_not n38029 ; n38030
g35595 and pi0644 n37583 ; n38031
g35596 and pi0644_not n38018 ; n38032
g35597 nor pi0715 n38031 ; n38033
g35598 and n38032_not n38033 ; n38034
g35599 nor pi0644 n38024 ; n38035
g35600 and pi0644 n37459_not ; n38036
g35601 and pi0715 n38036_not ; n38037
g35602 and n38035_not n38037 ; n38038
g35603 nor pi1160 n38038 ; n38039
g35604 and n38034_not n38039 ; n38040
g35605 nor n38030 n38040 ; n38041
g35606 and pi0790 n38041_not ; n38042
g35607 and pi0790_not n38018 ; n38043
g35608 nor n38042 n38043 ; n38044
g35609 nor po1038 n38044 ; n38045
g35610 and pi0224_not po1038 ; n38046
g35611 nor n38045 n38046 ; po0381
g35612 and n2547 n2625 ; n38048
g35613 and n3330 n38048 ; n38049
g35614 and pi0062_not n38049 ; n38050
g35615 nor n3328 n38050 ; n38051
g35616 and pi0062 n38049 ; n38052
g35617 and n2534 n38048 ; n38053
g35618 and pi0054 n38053_not ; n38054
g35619 and pi0092 n2533 ; n38055
g35620 and n38048 n38055 ; n38056
g35621 and n6169_not n6263 ; n38057
g35622 nor pi0137 n38057 ; n38058
g35623 and n7301 n38058_not ; n38059
g35624 and pi0075 n38059_not ; n38060
g35625 and pi0087 n38048 ; n38061
g35626 and n6286 n38058_not ; n38062
g35627 and pi0038 pi0137_not ; n38063
g35628 and pi0039 n2547 ; n38064
g35629 nor n2741 n2979 ; n38065
g35630 and pi0137 n38065_not ; n38066
g35631 nor n2740 n38066 ; n38067
g35632 nor pi0332 n38067 ; n38068
g35633 and n2517 n11417 ; n38069
g35634 and n2738 n38069_not ; n38070
g35635 and pi0137_not n2713 ; n38071
g35636 and n38070_not n38071 ; n38072
g35637 and n3168 n11417_not ; n38073
g35638 and n2903_not n38073 ; n38074
g35639 and n2746 n38074_not ; n38075
g35640 and n2744 n38075_not ; n38076
g35641 nor n2712 n38076 ; n38077
g35642 nor pi0095 n38077 ; n38078
g35643 and n3088 n38078_not ; n38079
g35644 and pi0332 n38072_not ; n38080
g35645 and n38079_not n38080 ; n38081
g35646 nor n38068 n38081 ; n38082
g35647 and pi0210 n38082_not ; n38083
g35648 and n2922 n38070_not ; n38084
g35649 and pi1093 n38084_not ; n38085
g35650 and n2922 n2933 ; n38086
g35651 and n2517 n7455_not ; n38087
g35652 and n2960_not n38087 ; n38088
g35653 nor pi0032 n38088 ; n38089
g35654 and n38086 n38089_not ; n38090
g35655 nor pi1093 n38090 ; n38091
g35656 and n2933_not n38084 ; n38092
g35657 and n11416 n38087 ; n38093
g35658 and n38086 n38093 ; n38094
g35659 nor n38092 n38094 ; n38095
g35660 and n38091 n38095 ; n38096
g35661 nor n38085 n38096 ; n38097
g35662 and n11549 n38097_not ; n38098
g35663 nor n2921 n38076 ; n38099
g35664 nor pi0095 n38099 ; n38100
g35665 nor n2741 n38100 ; n38101
g35666 and pi0137 n38101_not ; n38102
g35667 and n2933_not n3023 ; n38103
g35668 and n38091 n38103_not ; n38104
g35669 and n2997_not n38087 ; n38105
g35670 nor pi0032 n38105 ; n38106
g35671 and n38086 n38106_not ; n38107
g35672 and pi1093 n38103_not ; n38108
g35673 and n38107_not n38108 ; n38109
g35674 nor n38104 n38109 ; n38110
g35675 and n11517 n38110_not ; n38111
g35676 and n38095 n38111 ; n38112
g35677 nor n38098 n38112 ; n38113
g35678 and n38102_not n38113 ; n38114
g35679 and pi0332 n38114_not ; n38115
g35680 nor n2741 n2986 ; n38116
g35681 and pi0137 n38116_not ; n38117
g35682 and pi1093 n3023_not ; n38118
g35683 nor n38104 n38118 ; n38119
g35684 and n11549 n38119_not ; n38120
g35685 nor n38111 n38120 ; n38121
g35686 and n38117_not n38121 ; n38122
g35687 nor pi0332 n38122 ; n38123
g35688 nor n38115 n38123 ; n38124
g35689 and n2640_not n38124 ; n38125
g35690 nor pi0137 n38084 ; n38126
g35691 nor n38102 n38126 ; n38127
g35692 and pi0332 n38127_not ; n38128
g35693 nor n3024 n38117 ; n38129
g35694 nor pi0332 n38129 ; n38130
g35695 nor n38128 n38130 ; n38131
g35696 and n2640 n38131 ; n38132
g35697 nor pi0210 n38125 ; n38133
g35698 and n38132_not n38133 ; n38134
g35699 and pi0299 n38083_not ; n38135
g35700 and n38134_not n38135 ; n38136
g35701 and pi0198 n38082_not ; n38137
g35702 and n6260 n38131 ; n38138
g35703 and n6260_not n38124 ; n38139
g35704 nor pi0198 n38138 ; n38140
g35705 and n38139_not n38140 ; n38141
g35706 nor pi0299 n38137 ; n38142
g35707 and n38141_not n38142 ; n38143
g35708 nor n38136 n38143 ; n38144
g35709 nor pi0039 n38144 ; n38145
g35710 nor pi0038 n38064 ; n38146
g35711 and n38145_not n38146 ; n38147
g35712 and n6137 n38063_not ; n38148
g35713 and n38147_not n38148 ; n38149
g35714 nor n38062 n38149 ; n38150
g35715 nor pi0087 n38150 ; n38151
g35716 nor pi0075 n38061 ; n38152
g35717 and n38151_not n38152 ; n38153
g35718 nor pi0092 n38060 ; n38154
g35719 and n38153_not n38154 ; n38155
g35720 nor pi0054 n38056 ; n38156
g35721 and n38155_not n38156 ; n38157
g35722 nor pi0074 n38054 ; n38158
g35723 and n38157_not n38158 ; n38159
g35724 and pi0074 n6128 ; n38160
g35725 and n38048 n38160 ; n38161
g35726 nor pi0055 n38161 ; n38162
g35727 and n38159_not n38162 ; n38163
g35728 and n7348 n38163_not ; n38164
g35729 and pi0056 n2536 ; n38165
g35730 and n38048 n38165 ; n38166
g35731 nor n38164 n38166 ; n38167
g35732 nor pi0062 n38167 ; n38168
g35733 and n3328 n38052_not ; n38169
g35734 and n38168_not n38169 ; n38170
g35735 nor n6120 n38051 ; n38171
g35736 and n38170_not n38171 ; po0382
g35737 and pi0228 pi0231 ; n38173
g35738 nor n7360 n38173 ; n38174
g35739 and pi0056 n38174_not ; n38175
g35740 and pi0055 n38173_not ; n38176
g35741 nor n7364 n38173 ; n38177
g35742 and pi0074 n38177_not ; n38178
g35743 and pi0054 n38173_not ; n38179
g35744 nor n13971 n38173 ; n38180
g35745 and pi0075 n38180_not ; n38181
g35746 and pi0087 n38173_not ; n38182
g35747 and n7356_not n38182 ; n38183
g35748 nor n13975 n38173 ; n38184
g35749 and pi0100 n38184_not ; n38185
g35750 nor n2730 n3123 ; n38186
g35751 nor pi0070 n38186 ; n38187
g35752 nor pi0051 n38187 ; n38188
g35753 and n2748 n38188_not ; n38189
g35754 and n3168 n38189_not ; n38190
g35755 and n2746 n38190_not ; n38191
g35756 and n2744 n38191_not ; n38192
g35757 nor n6176 n38192 ; n38193
g35758 nor pi0095 n38193 ; n38194
g35759 and n2742 n38194_not ; n38195
g35760 nor pi0039 n38195 ; n38196
g35761 nor pi0038 n3402 ; n38197
g35762 and n38196_not n38197 ; n38198
g35763 and pi0228_not n38198 ; n38199
g35764 nor n38173 n38199 ; n38200
g35765 nor pi0100 n38200 ; n38201
g35766 nor pi0087 n38185 ; n38202
g35767 and n38201_not n38202 ; n38203
g35768 nor pi0075 n38183 ; n38204
g35769 and n38203_not n38204 ; n38205
g35770 nor pi0092 n38181 ; n38206
g35771 and n38205_not n38206 ; n38207
g35772 and pi0092 n38173_not ; n38208
g35773 and n7369_not n38208 ; n38209
g35774 nor n38207 n38209 ; n38210
g35775 nor pi0054 n38210 ; n38211
g35776 nor pi0074 n38179 ; n38212
g35777 and n38211_not n38212 ; n38213
g35778 nor pi0055 n38178 ; n38214
g35779 and n38213_not n38214 ; n38215
g35780 nor pi0056 n38176 ; n38216
g35781 and n38215_not n38216 ; n38217
g35782 nor pi0062 n38175 ; n38218
g35783 and n38217_not n38218 ; n38219
g35784 and pi0062 n38173_not ; n38220
g35785 and n7357_not n38220 ; n38221
g35786 nor n38219 n38221 ; n38222
g35787 and n3328 n38222_not ; n38223
g35788 nor n3328 n38173 ; n38224
g35789 nor n38223 n38224 ; po0383
g35790 and n13080 n13116_not ; n38226
g35791 and n6480 n38226 ; n38227
g35792 nor n6395 n38227 ; n38228
g35793 and pi1093 n38228_not ; n38229
g35794 and n2708 n6420 ; n38230
g35795 nor pi0091 n2761 ; n38231
g35796 and n38230 n38231_not ; n38232
g35797 nor pi0072 n38232 ; n38233
g35798 and n11022 n38230 ; n38234
g35799 and n7417_not n38234 ; n38235
g35800 and n8903_not n38233 ; n38236
g35801 and n38235_not n38236 ; n38237
g35802 and n6480 n38237_not ; n38238
g35803 nor n38229 n38238 ; n38239
g35804 and n38233 n38234_not ; n38240
g35805 and n6480 n38240_not ; n38241
g35806 and n10074 n38241_not ; n38242
g35807 and n2932_not n11022 ; n38243
g35808 and n2754 n11031 ; n38244
g35809 and n11029 n38244 ; n38245
g35810 and n38231 n38243_not ; n38246
g35811 and n38245_not n38246 ; n38247
g35812 and n38230 n38247_not ; n38248
g35813 nor pi0072 n38248 ; n38249
g35814 and n6480 n38249_not ; n38250
g35815 and pi0829 n6215_not ; n38251
g35816 and n38250_not n38251 ; n38252
g35817 nor n38239 n38242 ; n38253
g35818 and n38252_not n38253 ; n38254
g35819 nor pi0039 n38254 ; n38255
g35820 nand n11471 n38255_not ; po0384
g35821 and pi0039_not pi0228 ; n38257
g35822 nor n11420 n11425 ; n38258
g35823 and pi0039 n38258_not ; n38259
g35824 and n6391 n38259 ; n38260
g35825 nor n2930 n8904 ; n38261
g35826 and pi0032_not n10235 ; n38262
g35827 and n38261_not n38262 ; n38263
g35828 and n2967 n38263 ; n38264
g35829 and n11487_not n38264 ; n38265
g35830 nor n38260 n38265 ; n38266
g35831 and n10200 n38266_not ; n38267
g35832 or n38257 n38267 ; po0385
g35833 and n6136_not n10197 ; n38269
g35834 and pi0120 n6218 ; n38270
g35835 and n16652 n38270_not ; n38271
g35836 nor n35677 n38271 ; n38272
g35837 nor n6205 n38272 ; n38273
g35838 and n6198_not n16652 ; n38274
g35839 nor n38271 n38274 ; n38275
g35840 and n6205 n38275_not ; n38276
g35841 and pi0223 n38273_not ; n38277
g35842 and n38276_not n38277 ; n38278
g35843 and n2603 n16652 ; n38279
g35844 and n6213_not n7517 ; n38280
g35845 and n16661 n38280 ; n38281
g35846 and n16649 n38280_not ; n38282
g35847 and pi1091 n38281_not ; n38283
g35848 and n38282_not n38283 ; n38284
g35849 and n6383 n16661 ; n38285
g35850 and n6383_not n16649 ; n38286
g35851 nor pi1091 n38285 ; n38287
g35852 and n38286_not n38287 ; n38288
g35853 nor n38284 n38288 ; n38289
g35854 nor pi0120 n38289 ; n38290
g35855 nor n16651 n38290 ; n38291
g35856 and n6227_not n38291 ; n38292
g35857 nor n35677 n38292 ; n38293
g35858 and n6205_not n38293 ; n38294
g35859 and n6198 n38291 ; n38295
g35860 nor n38274 n38295 ; n38296
g35861 and n6205 n38296 ; n38297
g35862 nor n2603 n38294 ; n38298
g35863 and n38297_not n38298 ; n38299
g35864 nor pi0223 n38279 ; n38300
g35865 and n38299_not n38300 ; n38301
g35866 nor pi0299 n38278 ; n38302
g35867 and n38301_not n38302 ; n38303
g35868 nor n6242 n38272 ; n38304
g35869 and n6242 n38275_not ; n38305
g35870 and pi0215 n38304_not ; n38306
g35871 and n38305_not n38306 ; n38307
g35872 and n6242_not n38293 ; n38308
g35873 and n6242 n38296 ; n38309
g35874 nor n3448 n38308 ; n38310
g35875 and n38309_not n38310 ; n38311
g35876 nor pi0215 n16825 ; n38312
g35877 and n38311_not n38312 ; n38313
g35878 and pi0299 n38307_not ; n38314
g35879 and n38313_not n38314 ; n38315
g35880 nor n38303 n38315 ; n38316
g35881 and pi0039 n38316_not ; n38317
g35882 and n6170 n16854 ; n38318
g35883 and n16856_not n38318 ; n38319
g35884 nor pi0040 n38319 ; n38320
g35885 and n10289 n38320_not ; n38321
g35886 and pi0252 n38321_not ; n38322
g35887 and n6277 n16853_not ; n38323
g35888 and n38322_not n38323 ; n38324
g35889 and n6277_not n16866 ; n38325
g35890 nor pi1093 n38324 ; n38326
g35891 and n38325_not n38326 ; n38327
g35892 nor n6169 n6387 ; n38328
g35893 and n7417_not n16866 ; n38329
g35894 nor n16883 n38329 ; n38330
g35895 and n38328 n38330_not ; n38331
g35896 and pi0829 pi1091 ; n38332
g35897 and n16907 n38332 ; n38333
g35898 nor pi0824 n38333 ; n38334
g35899 and pi0824 n16902_not ; n38335
g35900 nor n6387 n38334 ; n38336
g35901 and n38335_not n38336 ; n38337
g35902 nor n16866 n38337 ; n38338
g35903 and n38332 n38334 ; n38339
g35904 nor n38335 n38339 ; n38340
g35905 and n2932 n6387_not ; n38341
g35906 and n38340_not n38341 ; n38342
g35907 nor n38328 n38338 ; n38343
g35908 and n38342_not n38343 ; n38344
g35909 and pi1093 n38331_not ; n38345
g35910 and n38344_not n38345 ; n38346
g35911 nor pi0039 n38327 ; n38347
g35912 and n38346_not n38347 ; n38348
g35913 nor pi0038 n38317 ; n38349
g35914 and n38348_not n38349 ; n38350
g35915 and n38269 n38350_not ; po0387
g35916 nor pi0081 n2865 ; n38352
g35917 and n6443 n38352_not ; n38353
g35918 and n2462 n38353_not ; n38354
g35919 and n2873 n38354_not ; n38355
g35920 and n2785 n38355_not ; n38356
g35921 and n2877 n38356_not ; n38357
g35922 and n2719 n38357_not ; n38358
g35923 nor n2722 n38358 ; n38359
g35924 nor pi0086 n38359 ; n38360
g35925 and n2783 n38360_not ; n38361
g35926 and n2781 n38361_not ; n38362
g35927 nor n2776 n38362 ; n38363
g35928 nor pi0108 n38363 ; n38364
g35929 and n2775 n38364_not ; n38365
g35930 and n2889 n38365_not ; n38366
g35931 nor n2766 n38366 ; n38367
g35932 and n2765 n38367_not ; n38368
g35933 and n2764 n38368_not ; n38369
g35934 and n2757 n38369_not ; n38370
g35935 and n3108 n38370_not ; n38371
g35936 and n2504 n38371_not ; n38372
g35937 and n15635 n38372_not ; n38373
g35938 nor pi0070 n38373 ; n38374
g35939 nor n3099 n38374 ; n38375
g35940 nor pi0051 n38375 ; n38376
g35941 and n2748 n38376_not ; n38377
g35942 and n3168 n38377_not ; n38378
g35943 and n2746 n38378_not ; n38379
g35944 and pi1082_not n2743 ; n38380
g35945 nor pi0032 n38380 ; n38381
g35946 and n38379_not n38381 ; n38382
g35947 nor n3412 n38382 ; n38383
g35948 nor pi0095 n38383 ; n38384
g35949 nor n2741 n38384 ; n38385
g35950 nor pi0039 n38385 ; n38386
g35951 nor n7307 n7309 ; n38387
g35952 nand n2932 n6217 ; po0950
g35953 and n6381 po0950_not ; n38389
g35954 and n38387_not n38389 ; n38390
g35955 and n6185 n11369 ; n38391
g35956 and n38390_not n38391 ; n38392
g35957 nor n3402 n38392 ; n38393
g35958 and n38386_not n38393 ; n38394
g35959 nor pi0038 n38394 ; n38395
g35960 and n6137 n38395_not ; n38396
g35961 nor pi0087 n6286 ; n38397
g35962 and n38396_not n38397 ; n38398
g35963 nor n6132 n38398 ; n38399
g35964 and n2569 n38399_not ; n38400
g35965 and n7306 n38400_not ; n38401
g35966 nor pi0054 n38401 ; n38402
g35967 nor n7341 n38402 ; n38403
g35968 and n8879 n38403_not ; n38404
g35969 and n15712 n38404_not ; n38405
g35970 nor pi0056 n38405 ; n38406
g35971 nor n6127 n38406 ; n38407
g35972 nor pi0062 n38407 ; n38408
g35973 nor n6299 n38408 ; n38409
g35974 and n3328 n38409_not ; n38410
g35975 and n6123 n38410_not ; po0389
g35976 nor pi0230 pi0233 ; n38412
g35977 nor pi0212 pi0214 ; n38413
g35978 nor pi0211 n38413 ; n38414
g35979 and pi0219 n38414_not ; n38415
g35980 and po1038 n38415_not ; n38416
g35981 and pi1142 n10486_not ; n38417
g35982 and pi0211 pi1143 ; n38418
g35983 and pi0211_not pi1144 ; n38419
g35984 nor n38418 n38419 ; n38420
g35985 and pi0212_not pi0214 ; n38421
g35986 and pi0212 pi0214_not ; n38422
g35987 nor n38421 n38422 ; n38423
g35988 nor n38420 n38423 ; n38424
g35989 and pi0211_not pi1143 ; n38425
g35990 and n10843 n38425 ; n38426
g35991 nor n38424 n38426 ; n38427
g35992 nor pi0219 n38427 ; n38428
g35993 nor n38417 n38428 ; n38429
g35994 and n38416 n38429_not ; n38430
g35995 and pi0299 n38420_not ; n38431
g35996 and pi0199 pi1142 ; n38432
g35997 nor pi0200 n38432 ; n38433
g35998 and pi0199_not pi1144 ; n38434
g35999 and n38433 n38434_not ; n38435
g36000 and pi0199_not pi1143 ; n38436
g36001 and pi0200 n38436_not ; n38437
g36002 nor n38435 n38437 ; n38438
g36003 nor pi0299 n38438 ; n38439
g36004 nor pi0207 n38439 ; n38440
g36005 and pi0207 pi0299_not ; n38441
g36006 and n38433 n38436_not ; n38442
g36007 and pi0199_not pi1142 ; n38443
g36008 and pi0200 n38443_not ; n38444
g36009 and n38441 n38444_not ; n38445
g36010 and n38442_not n38445 ; n38446
g36011 nor n38440 n38446 ; n38447
g36012 and pi0208 n38447_not ; n38448
g36013 and pi0207 pi0208_not ; n38449
g36014 and n38438 n38449 ; n38450
g36015 nor n38448 n38450 ; n38451
g36016 nor pi0299 n38451 ; n38452
g36017 nor pi0214 n38452 ; n38453
g36018 and n38431_not n38453 ; n38454
g36019 and pi0211 pi1142 ; n38455
g36020 nor n38425 n38455 ; n38456
g36021 and pi0299 n38456_not ; n38457
g36022 and pi0214 n38457_not ; n38458
g36023 and n38452_not n38458 ; n38459
g36024 and pi0212 n38459_not ; n38460
g36025 and n38454_not n38460 ; n38461
g36026 nor n38431 n38452 ; n38462
g36027 nor pi0212 n38453 ; n38463
g36028 and n38462_not n38463 ; n38464
g36029 nor pi0219 n38461 ; n38465
g36030 and n38464_not n38465 ; n38466
g36031 and n38414_not n38452 ; n38467
g36032 and pi0299_not n38451 ; n38468
g36033 and pi0299 pi1142_not ; n38469
g36034 and n38414 n38469_not ; n38470
g36035 and n38468_not n38470 ; n38471
g36036 and pi0219 n38467_not ; n38472
g36037 and n38471_not n38472 ; n38473
g36038 nor po1038 n38473 ; n38474
g36039 and n38466_not n38474 ; n38475
g36040 nor n38430 n38475 ; n38476
g36041 and pi0213 n38476 ; n38477
g36042 and pi0211_not pi1157 ; n38478
g36043 and pi0211 pi1156 ; n38479
g36044 nor n38478 n38479 ; n38480
g36045 and pi0214 n38480_not ; n38481
g36046 nor pi0212 n38481 ; n38482
g36047 and pi0211_not pi1156 ; n38483
g36048 and pi0211 pi1155 ; n38484
g36049 nor n38483 n38484 ; n38485
g36050 nor pi0214 n38485 ; n38486
g36051 and pi0211_not pi1155 ; n38487
g36052 and pi0211 pi1154 ; n38488
g36053 nor n38487 n38488 ; n38489
g36054 and pi0214 n38489_not ; n38490
g36055 nor n38486 n38490 ; n38491
g36056 and pi0212 n38491 ; n38492
g36057 nor n38482 n38492 ; n38493
g36058 nor pi0219 n38493 ; n38494
g36059 and pi0211_not pi1154 ; n38495
g36060 nor pi0214 n38495 ; n38496
g36061 and pi0211_not pi1153 ; n38497
g36062 and n10843 n38497_not ; n38498
g36063 and pi0211_not pi0214 ; n38499
g36064 and pi1155 n38499 ; n38500
g36065 nor pi0212 n38500 ; n38501
g36066 nor n38496 n38498 ; n38502
g36067 and n38501_not n38502 ; n38503
g36068 and pi0219 n38503_not ; n38504
g36069 and po1038 n38504_not ; n38505
g36070 and n38494_not n38505 ; n38506
g36071 nor pi0213 n38506 ; n38507
g36072 and pi0219_not pi0299 ; n38508
g36073 and n38493 n38508 ; n38509
g36074 and pi0299 pi1155 ; n38510
g36075 and n38421 n38510 ; n38511
g36076 and pi0299 pi1153 ; n38512
g36077 and pi0214 n38512_not ; n38513
g36078 and pi0299 pi1154 ; n38514
g36079 nor pi0214 n38514 ; n38515
g36080 and pi0212 n38513_not ; n38516
g36081 and n38515_not n38516 ; n38517
g36082 nor n38511 n38517 ; n38518
g36083 and pi0211_not pi0219 ; n38519
g36084 and n38518_not n38519 ; n38520
g36085 nor n38509 n38520 ; n38521
g36086 and n38452_not n38521 ; n38522
g36087 nor po1038 n38522 ; n38523
g36088 and n38507 n38523_not ; n38524
g36089 and pi0209 n38524_not ; n38525
g36090 and n38477_not n38525 ; n38526
g36091 and pi0211_not n10843 ; n38527
g36092 and pi0299 pi1143_not ; n38528
g36093 and pi0200_not pi1155 ; n38529
g36094 and pi0199 n38529 ; n38530
g36095 and pi0299_not n38530 ; n38531
g36096 nor pi1156 n38531 ; n38532
g36097 nor pi0299 n11444 ; n38533
g36098 and pi1156 n38530_not ; n38534
g36099 and n38533 n38534 ; n38535
g36100 nor n38532 n38535 ; n38536
g36101 and pi0207 n38536 ; n38537
g36102 nor pi0299 n38537 ; n38538
g36103 nor pi0208 n38538 ; n38539
g36104 and pi1157_not n38539 ; n38540
g36105 and n38528_not n38540 ; n38541
g36106 and pi0208_not pi1157 ; n38542
g36107 and pi0299 pi1143 ; n38543
g36108 nor pi1155 n10810 ; n38544
g36109 and pi0200 pi0299_not ; n38545
g36110 and pi1155 n38545_not ; n38546
g36111 nor n38544 n38546 ; n38547
g36112 and pi0199 pi1155_not ; n38548
g36113 and pi0199 pi0200 ; n38549
g36114 nor pi0299 n38549 ; n38550
g36115 and pi1156 n38548_not ; n38551
g36116 and n38550 n38551 ; n38552
g36117 and n38547 n38552_not ; n38553
g36118 and pi0207 n38528_not ; n38554
g36119 and n38553_not n38554 ; n38555
g36120 nor n38543 n38555 ; n38556
g36121 and n38542 n38556_not ; n38557
g36122 and pi1153 n38550_not ; n38558
g36123 and pi1154 n38558_not ; n38559
g36124 and n11384 n38529 ; n38560
g36125 nor n10809 n38549 ; n38561
g36126 nor pi1153 n11384 ; n38562
g36127 and pi1154 n38561 ; n38563
g36128 and n38562_not n38563 ; n38564
g36129 nor n38560 n38564 ; n38565
g36130 and n38559 n38565_not ; n38566
g36131 nor pi0199 pi1155 ; n38567
g36132 nor pi0200 pi0299 ; n38568
g36133 and pi0199 pi1153_not ; n38569
g36134 and n38568 n38569_not ; n38570
g36135 nor pi1154 n38567 ; n38571
g36136 and n38570 n38571 ; n38572
g36137 nor n38566 n38572 ; n38573
g36138 and pi0207 n38573 ; n38574
g36139 and n38543_not n38574 ; n38575
g36140 and pi0199_not pi1155 ; n38576
g36141 and n38545 n38576 ; n38577
g36142 nor pi1154 n38577 ; n38578
g36143 and n38543_not n38578 ; n38579
g36144 and pi1155_not n38543 ; n38580
g36145 nor pi0299 n38561 ; n38581
g36146 and pi1155 n38581_not ; n38582
g36147 and n38528_not n38582 ; n38583
g36148 nor pi0200 pi1155 ; n38584
g36149 and n11373 n38584 ; n38585
g36150 and pi1154 n38585_not ; n38586
g36151 and n38580_not n38586 ; n38587
g36152 and n38583_not n38587 ; n38588
g36153 nor pi1156 n38579 ; n38589
g36154 and n38588_not n38589 ; n38590
g36155 and pi0200 n38576_not ; n38591
g36156 nor pi0299 n38591 ; n38592
g36157 and pi1154 n38592_not ; n38593
g36158 and n38543_not n38593 ; n38594
g36159 and pi1155 n11373_not ; n38595
g36160 nor n38544 n38595 ; n38596
g36161 nor n38528 n38596 ; n38597
g36162 nor pi1154 n38597 ; n38598
g36163 and pi1156 n38594_not ; n38599
g36164 and n38598_not n38599 ; n38600
g36165 nor n38590 n38600 ; n38601
g36166 and pi0207_not n38601 ; n38602
g36167 and pi0208 n38575_not ; n38603
g36168 and n38602_not n38603 ; n38604
g36169 nor n38541 n38557 ; n38605
g36170 and n38604_not n38605 ; n38606
g36171 and n38527 n38606 ; n38607
g36172 nor n10843 n38413 ; n38608
g36173 and pi0211 n38606_not ; n38609
g36174 and pi0299 pi1144_not ; n38610
g36175 and n38540 n38610_not ; n38611
g36176 and pi0299 pi1144 ; n38612
g36177 and pi0207 n38610_not ; n38613
g36178 and n38553_not n38613 ; n38614
g36179 nor n38612 n38614 ; n38615
g36180 and n38542 n38615_not ; n38616
g36181 and n38574 n38612_not ; n38617
g36182 and n38578 n38612_not ; n38618
g36183 and pi1155_not n38612 ; n38619
g36184 and n38582 n38610_not ; n38620
g36185 and n38586 n38619_not ; n38621
g36186 and n38620_not n38621 ; n38622
g36187 nor pi1156 n38618 ; n38623
g36188 and n38622_not n38623 ; n38624
g36189 and n38593 n38612_not ; n38625
g36190 nor n38596 n38610 ; n38626
g36191 nor pi1154 n38626 ; n38627
g36192 and pi1156 n38625_not ; n38628
g36193 and n38627_not n38628 ; n38629
g36194 nor n38624 n38629 ; n38630
g36195 and pi0207_not n38630 ; n38631
g36196 and pi0208 n38617_not ; n38632
g36197 and n38631_not n38632 ; n38633
g36198 nor n38611 n38616 ; n38634
g36199 and n38633_not n38634 ; n38635
g36200 nor pi0211 n38635 ; n38636
g36201 and n38608 n38609_not ; n38637
g36202 and n38636_not n38637 ; n38638
g36203 nor n38607 n38638 ; n38639
g36204 nor pi0219 n38639 ; n38640
g36205 and pi0299_not n38561 ; n38641
g36206 and n38584_not n38641 ; n38642
g36207 and n38532_not n38642 ; n38643
g36208 and pi0207 n38643 ; n38644
g36209 nor pi0208 n38644 ; n38645
g36210 and n10810 n38591_not ; n38646
g36211 and n38578_not n38646 ; n38647
g36212 and pi0200 pi1155_not ; n38648
g36213 and n11384 n38648_not ; n38649
g36214 and pi1156 n38649 ; n38650
g36215 nor n38647 n38650 ; n38651
g36216 and pi0207_not n38651 ; n38652
g36217 nor n38574 n38652 ; n38653
g36218 and pi0208 n38653_not ; n38654
g36219 nor n38645 n38654 ; n38655
g36220 nor pi1157 n38655 ; n38656
g36221 nor pi1156 n38548 ; n38657
g36222 and n38568 n38657 ; n38658
g36223 nor n38552 n38658 ; n38659
g36224 and pi0207 n38659_not ; n38660
g36225 nor pi0208 n38660 ; n38661
g36226 nor n38654 n38661 ; n38662
g36227 and pi1157 n38662_not ; n38663
g36228 nor n38656 n38663 ; n38664
g36229 nor pi0219 n38413 ; n38665
g36230 nor n38414 n38665 ; n38666
g36231 and n38664_not n38666 ; n38667
g36232 nor pi1157 n38539 ; n38668
g36233 nor pi1156 n38547 ; n38669
g36234 and n11373 n38529_not ; n38670
g36235 and pi1156 n38670_not ; n38671
g36236 nor n38669 n38671 ; n38672
g36237 and pi0207 n38672 ; n38673
g36238 nor pi0207 pi0299 ; n38674
g36239 nor pi0208 n38674 ; n38675
g36240 and n38673_not n38675 ; n38676
g36241 and pi1157 n38676_not ; n38677
g36242 nor n38469 n38668 ; n38678
g36243 and n38677_not n38678 ; n38679
g36244 and pi0299 pi1142 ; n38680
g36245 and pi1153 n38585 ; n38681
g36246 and pi1153 n38545_not ; n38682
g36247 nor pi1153 n10810 ; n38683
g36248 nor n38682 n38683 ; n38684
g36249 and pi1155 n38684_not ; n38685
g36250 nor n38681 n38685 ; n38686
g36251 nor pi1154 n38686 ; n38687
g36252 and n38569_not n38641 ; n38688
g36253 nor n38595 n38688 ; n38689
g36254 and pi1154 n38689_not ; n38690
g36255 nor n38687 n38690 ; n38691
g36256 nor pi0299 n38691 ; n38692
g36257 and pi0207 n38680_not ; n38693
g36258 and n38692_not n38693 ; n38694
g36259 nor n38577 n38680 ; n38695
g36260 nor pi1154 pi1156 ; n38696
g36261 and n38695_not n38696 ; n38697
g36262 and pi1156 n38596_not ; n38698
g36263 and pi0199 pi0200_not ; n38699
g36264 nor pi0299 n38699 ; n38700
g36265 nor pi1155 n38700 ; n38701
g36266 nor n38582 n38701 ; n38702
g36267 and pi1154 n38702_not ; n38703
g36268 nor n38698 n38703 ; n38704
g36269 nor n38469 n38704 ; n38705
g36270 nor pi0207 n38697 ; n38706
g36271 and n38705_not n38706 ; n38707
g36272 and pi0208 n38707_not ; n38708
g36273 and n38694_not n38708 ; n38709
g36274 nor n10486 n38666 ; n38710
g36275 and n38679_not n38710 ; n38711
g36276 and n38709_not n38711 ; n38712
g36277 nor po1038 n38712 ; n38713
g36278 and n38667_not n38713 ; n38714
g36279 and n38640_not n38714 ; n38715
g36280 and pi0213 n38430_not ; n38716
g36281 and n38715_not n38716 ; n38717
g36282 and pi0211 n38664_not ; n38718
g36283 nor pi0214 n38664 ; n38719
g36284 nor pi0212 n38719 ; n38720
g36285 nor pi0207 n38510 ; n38721
g36286 nor pi0208 n38721 ; n38722
g36287 nor n11384 n38546 ; n38723
g36288 and pi1156 n38723_not ; n38724
g36289 nor pi1156 n38545 ; n38725
g36290 and n38701_not n38725 ; n38726
g36291 nor n38724 n38726 ; n38727
g36292 and pi0207 n38727 ; n38728
g36293 and pi1157 n38722 ; n38729
g36294 and n38728_not n38729 ; n38730
g36295 nor pi1155 n11384 ; n38731
g36296 and pi0299_not n38532 ; n38732
g36297 nor n38581 n38731 ; n38733
g36298 and n38732_not n38733 ; n38734
g36299 and n38722 n38734 ; n38735
g36300 and pi0207 n38691 ; n38736
g36301 and n38651 n38721 ; n38737
g36302 and pi0208 n38737_not ; n38738
g36303 and n38736_not n38738 ; n38739
g36304 nor n38730 n38735 ; n38740
g36305 and n38739_not n38740 ; n38741
g36306 and n38499 n38741 ; n38742
g36307 and n38720 n38742_not ; n38743
g36308 nor pi0211 pi0214 ; n38744
g36309 and pi0299 pi1154_not ; n38745
g36310 and pi1157 n38745_not ; n38746
g36311 and n38676 n38746 ; n38747
g36312 and n38651 n38703_not ; n38748
g36313 nor pi0207 n38748 ; n38749
g36314 and pi0299_not n38689 ; n38750
g36315 and pi1154 n38750_not ; n38751
g36316 nor n38572 n38751 ; n38752
g36317 and pi0207 n38752_not ; n38753
g36318 nor n38749 n38753 ; n38754
g36319 and pi0208 n38754_not ; n38755
g36320 nor n38514 n38644 ; n38756
g36321 nor pi0208 n38756 ; n38757
g36322 and pi1157_not n38757 ; n38758
g36323 nor n38747 n38758 ; n38759
g36324 and n38755_not n38759 ; n38760
g36325 and n38744 n38760 ; n38761
g36326 and pi1153 n38700_not ; n38762
g36327 and n38565 n38762_not ; n38763
g36328 and pi0207 n38763_not ; n38764
g36329 and pi0299 pi1155_not ; n38765
g36330 and pi1155 n38533_not ; n38766
g36331 nor n38765 n38766 ; n38767
g36332 and n38704 n38767 ; n38768
g36333 and pi0299 pi1153_not ; n38769
g36334 nor pi0207 n38769 ; n38770
g36335 and n38768_not n38770 ; n38771
g36336 nor n38764 n38771 ; n38772
g36337 and pi0208 n38772_not ; n38773
g36338 nor n38668 n38769 ; n38774
g36339 and n38677_not n38774 ; n38775
g36340 and n38499 n38773_not ; n38776
g36341 and n38775_not n38776 ; n38777
g36342 and pi0212 n38761_not ; n38778
g36343 and n38777_not n38778 ; n38779
g36344 nor n38743 n38779 ; n38780
g36345 nor n38718 n38780 ; n38781
g36346 and pi0219 n38781_not ; n38782
g36347 nor n10484 n38744 ; n38783
g36348 and n38741_not n38783 ; n38784
g36349 and n10484 n38760_not ; n38785
g36350 and n38532_not n38539 ; n38786
g36351 and pi0299 pi1156 ; n38787
g36352 nor n38660 n38787 ; n38788
g36353 and n38542 n38788_not ; n38789
g36354 and pi0207 n38573_not ; n38790
g36355 nor n38647 n38698 ; n38791
g36356 nor pi0207 n38791 ; n38792
g36357 and pi0207 n38787 ; n38793
g36358 nor n38792 n38793 ; n38794
g36359 and n38790_not n38794 ; n38795
g36360 and pi0208 n38795_not ; n38796
g36361 nor n38786 n38789 ; n38797
g36362 and n38796_not n38797 ; n38798
g36363 and n38744 n38798_not ; n38799
g36364 nor n38784 n38799 ; n38800
g36365 and n38785_not n38800 ; n38801
g36366 and pi0212 n38801_not ; n38802
g36367 and pi0211 n38798_not ; n38803
g36368 and pi0207_not n38768 ; n38804
g36369 and n38441 n38763 ; n38805
g36370 and pi0208 n38805_not ; n38806
g36371 and n38804_not n38806 ; n38807
g36372 and n38677 n38807_not ; n38808
g36373 nor pi0211 n38808 ; n38809
g36374 and n38656_not n38809 ; n38810
g36375 and pi0214 n38803_not ; n38811
g36376 and n38810_not n38811 ; n38812
g36377 and n38720 n38812_not ; n38813
g36378 nor pi0219 n38802 ; n38814
g36379 and n38813_not n38814 ; n38815
g36380 nor po1038 n38815 ; n38816
g36381 and n38782_not n38816 ; n38817
g36382 and n38507 n38817_not ; n38818
g36383 nor pi0209 n38717 ; n38819
g36384 and n38818_not n38819 ; n38820
g36385 nor n38526 n38820 ; n38821
g36386 and pi0230 n38821_not ; n38822
g36387 or n38412 n38822 ; po0390
g36388 and n10487_not n38651 ; n38824
g36389 nor pi0207 pi0208 ; n38825
g36390 nor n10487 n38825 ; n38826
g36391 and pi0199_not n38584 ; n38827
g36392 nor pi1154 n38560 ; n38828
g36393 and n38550 n38827_not ; n38829
g36394 and n38828_not n38829 ; n38830
g36395 and pi0207 n38830 ; n38831
g36396 nor n38826 n38831 ; n38832
g36397 nor n38824 n38832 ; n38833
g36398 and n38414_not n38833 ; n38834
g36399 and pi0219 n38834_not ; n38835
g36400 and pi0207_not n38514 ; n38836
g36401 and pi0207 n38748_not ; n38837
g36402 nor n38836 n38837 ; n38838
g36403 nor pi0208 n38838 ; n38839
g36404 and pi1155_not n10809 ; n38840
g36405 nor n38549 n38840 ; n38841
g36406 nor pi0299 n38841 ; n38842
g36407 nor n38828 n38842 ; n38843
g36408 and pi0207 n38843 ; n38844
g36409 nor n38749 n38844 ; n38845
g36410 and pi0208 n38845_not ; n38846
g36411 nor n38839 n38846 ; n38847
g36412 nor pi0211 n38847 ; n38848
g36413 and n38413_not n38848 ; n38849
g36414 and n38835 n38849_not ; n38850
g36415 nor pi0214 n38833 ; n38851
g36416 nor pi0212 n38851 ; n38852
g36417 and pi0207 n38791_not ; n38853
g36418 nor n38787 n38853 ; n38854
g36419 nor pi0208 n38854 ; n38855
g36420 and n38794 n38831_not ; n38856
g36421 and pi0208 n38856_not ; n38857
g36422 nor n38855 n38857 ; n38858
g36423 nor pi0211 n38858 ; n38859
g36424 and n38510_not n38651 ; n38860
g36425 and n38722 n38860_not ; n38861
g36426 and pi0207 n38510_not ; n38862
g36427 and n38830_not n38862 ; n38863
g36428 and pi0208 n38863_not ; n38864
g36429 and n38737_not n38864 ; n38865
g36430 nor n38861 n38865 ; n38866
g36431 and pi0211 n38866_not ; n38867
g36432 nor n38859 n38867 ; n38868
g36433 and pi0214 n38868 ; n38869
g36434 and n38852 n38869_not ; n38870
g36435 and pi0211 n38847_not ; n38871
g36436 nor pi0211 n38866 ; n38872
g36437 and pi0214 n38872_not ; n38873
g36438 and n38871_not n38873 ; n38874
g36439 and pi0214_not n38868 ; n38875
g36440 and pi0212 n38874_not ; n38876
g36441 and n38875_not n38876 ; n38877
g36442 nor pi0219 n38870 ; n38878
g36443 and n38877_not n38878 ; n38879
g36444 and n35819 n38850_not ; n38880
g36445 and n38879_not n38880 ; n38881
g36446 and pi0211 pi1153 ; n38882
g36447 nor n38495 n38882 ; n38883
g36448 and n10843_not n38883 ; n38884
g36449 and n38665 n38884_not ; n38885
g36450 and n38498_not n38885 ; n38886
g36451 and po1038 n38886 ; n38887
g36452 nor pi1152 n38887 ; n38888
g36453 and pi0207 n38767 ; n38889
g36454 and n38704 n38889 ; n38890
g36455 and n38675 n38890_not ; n38891
g36456 and n38441 n38843_not ; n38892
g36457 and pi0208 n38892_not ; n38893
g36458 and n38804_not n38893 ; n38894
g36459 nor n38891 n38894 ; n38895
g36460 nor n38769 n38895 ; n38896
g36461 and pi0211 n38896 ; n38897
g36462 nor n38848 n38897 ; n38898
g36463 and pi0214 n38898 ; n38899
g36464 and n38852 n38899_not ; n38900
g36465 nor pi0219 n38900 ; n38901
g36466 nor pi0214 n38898 ; n38902
g36467 nor pi0211 n38896 ; n38903
g36468 and pi0214 n38903_not ; n38904
g36469 and pi0211 n38833_not ; n38905
g36470 and n38904 n38905_not ; n38906
g36471 nor n38902 n38906 ; n38907
g36472 and pi0212 n38907_not ; n38908
g36473 and n38901 n38908_not ; n38909
g36474 and pi0219 n38833_not ; n38910
g36475 nor po1038 n38910 ; n38911
g36476 and n38909_not n38911 ; n38912
g36477 and n38888 n38912_not ; n38913
g36478 and pi1153 n38744_not ; n38914
g36479 nor n38496 n38499 ; n38915
g36480 nor n38914 n38915 ; n38916
g36481 and pi0212 n38916_not ; n38917
g36482 and n38421 n38883_not ; n38918
g36483 nor pi0219 n38918 ; n38919
g36484 and n38917_not n38919 ; n38920
g36485 and n38416 n38920_not ; n38921
g36486 and pi1152 n38921_not ; n38922
g36487 and n38895_not n38904 ; n38923
g36488 nor n38902 n38923 ; n38924
g36489 and pi0212 n38924_not ; n38925
g36490 and n38901 n38925_not ; n38926
g36491 and n38414 n38895_not ; n38927
g36492 and n38835 n38927_not ; n38928
g36493 nor po1038 n38928 ; n38929
g36494 and n38926_not n38929 ; n38930
g36495 and n38922 n38930_not ; n38931
g36496 nor pi0213 n38913 ; n38932
g36497 and n38931_not n38932 ; n38933
g36498 and pi0209 n38881_not ; n38934
g36499 and n38933_not n38934 ; n38935
g36500 and pi0199_not pi1153 ; n38936
g36501 and pi0200 n38936 ; n38937
g36502 and pi0299_not n38937 ; n38938
g36503 nor pi1154 n38938 ; n38939
g36504 and pi1154 n38545 ; n38940
g36505 and n38936_not n38940 ; n38941
g36506 nor n38939 n38941 ; n38942
g36507 and n38700 n38942_not ; n38943
g36508 and n38675 n38943_not ; n38944
g36509 nor pi0200 pi1153 ; n38945
g36510 nor pi0199 n38945 ; n38946
g36511 nor pi0299 n38946 ; n38947
g36512 and n38699_not n38947 ; n38948
g36513 and pi0207 n38948 ; n38949
g36514 and pi0207_not n38943 ; n38950
g36515 and pi0208 n38949_not ; n38951
g36516 and n38950_not n38951 ; n38952
g36517 nor n38944 n38952 ; n38953
g36518 and pi0211_not n38953 ; n38954
g36519 and pi0299_not n10809 ; n38955
g36520 nor pi1153 n38955 ; n38956
g36521 and n38559 n38956_not ; n38957
g36522 nor pi0199 pi1153 ; n38958
g36523 and n38641 n38958_not ; n38959
g36524 nor n38957 n38959 ; n38960
g36525 and n10487_not n38960 ; n38961
g36526 and pi1153_not n10809 ; n38962
g36527 and n38550 n38962_not ; n38963
g36528 and n10487 n38963_not ; n38964
g36529 nor n38825 n38964 ; n38965
g36530 and n38961_not n38965 ; n38966
g36531 and pi0211 n38966_not ; n38967
g36532 nor n38954 n38967 ; n38968
g36533 and n38413_not n38968 ; n38969
g36534 and pi0219 n38413_not ; n38970
g36535 and pi0219 n38966_not ; n38971
g36536 nor n38970 n38971 ; n38972
g36537 nor n38969 n38972 ; n38973
g36538 nor po1038 n38973 ; n38974
g36539 and pi0207_not n38512 ; n38975
g36540 nor pi1153 n38568 ; n38976
g36541 nor n38581 n38976 ; n38977
g36542 and pi1154 n11373_not ; n38978
g36543 and n38976_not n38978 ; n38979
g36544 nor n38977 n38979 ; n38980
g36545 and pi0207 n38980_not ; n38981
g36546 nor n38975 n38981 ; n38982
g36547 nor pi0208 n38982 ; n38983
g36548 nor pi0207 n38980 ; n38984
g36549 and pi0299_not n38549 ; n38985
g36550 and pi0207 n38985_not ; n38986
g36551 and n38683_not n38986 ; n38987
g36552 nor n38984 n38987 ; n38988
g36553 and pi0208 n38988_not ; n38989
g36554 nor n38983 n38989 ; n38990
g36555 nor pi0211 n38990 ; n38991
g36556 and pi0211 n38953_not ; n38992
g36557 and pi0214 n38991_not ; n38993
g36558 and n38992_not n38993 ; n38994
g36559 and pi0207 n38960_not ; n38995
g36560 nor n38514 n38995 ; n38996
g36561 nor pi0208 n38996 ; n38997
g36562 and pi0207 n38948_not ; n38998
g36563 and n38745_not n38998 ; n38999
g36564 and pi1154 n10810_not ; n39000
g36565 nor n38957 n39000 ; n39001
g36566 and n38959_not n39001 ; n39002
g36567 nor pi0207 n39002 ; n39003
g36568 nor n38999 n39003 ; n39004
g36569 and pi0208 n39004_not ; n39005
g36570 nor n38997 n39005 ; n39006
g36571 nor pi0211 n39006 ; n39007
g36572 and pi0211 n38990_not ; n39008
g36573 nor n39007 n39008 ; n39009
g36574 and pi0214_not n39009 ; n39010
g36575 and pi0212 n38994_not ; n39011
g36576 and n39010_not n39011 ; n39012
g36577 nor pi0214 n38966 ; n39013
g36578 nor pi0212 n39013 ; n39014
g36579 and pi0214 n39009 ; n39015
g36580 and n39014 n39015_not ; n39016
g36581 nor pi0219 n39012 ; n39017
g36582 and n39016_not n39017 ; n39018
g36583 and n38974 n39018_not ; n39019
g36584 and n38922 n39019_not ; n39020
g36585 and pi0200 pi1153_not ; n39021
g36586 and n11384 n39021_not ; n39022
g36587 and pi1154 n39022_not ; n39023
g36588 nor n38939 n39023 ; n39024
g36589 and n38826 n39024 ; n39025
g36590 and pi0208 n38441 ; n39026
g36591 and pi1153 n10810_not ; n39027
g36592 and n39026 n39027 ; n39028
g36593 nor n39025 n39028 ; n39029
g36594 and pi0219 n39029 ; n39030
g36595 nor po1038 n39030 ; n39031
g36596 and pi1153 pi1154_not ; n39032
g36597 and n38533_not n39032 ; n39033
g36598 nor n38979 n39033 ; n39034
g36599 and pi0207 n39034_not ; n39035
g36600 nor n38975 n39035 ; n39036
g36601 nor pi0208 n39036 ; n39037
g36602 nor pi0207 n39034 ; n39038
g36603 and pi0207 n10810_not ; n39039
g36604 and pi1153 n39039 ; n39040
g36605 nor n39038 n39040 ; n39041
g36606 and pi0208 n39041_not ; n39042
g36607 nor n39037 n39042 ; n39043
g36608 and n38527 n39043 ; n39044
g36609 and pi1153 n11373_not ; n39045
g36610 nor n38683 n39045 ; n39046
g36611 and pi1154 n39046_not ; n39047
g36612 nor n38938 n39047 ; n39048
g36613 and pi0207 n39048_not ; n39049
g36614 nor n38836 n39049 ; n39050
g36615 nor pi0208 n39050 ; n39051
g36616 nor pi0299 pi1153 ; n39052
g36617 nor n10810 n39052 ; n39053
g36618 and n38745_not n39053 ; n39054
g36619 and pi0207 n39054_not ; n39055
g36620 and pi0207_not n39048 ; n39056
g36621 and pi0208 n39055_not ; n39057
g36622 and n39056_not n39057 ; n39058
g36623 nor n39051 n39058 ; n39059
g36624 and pi0211_not n39059 ; n39060
g36625 and pi0211 n39043 ; n39061
g36626 nor n39060 n39061 ; n39062
g36627 and n38608 n39062_not ; n39063
g36628 nor n39044 n39063 ; n39064
g36629 nor pi0219 n39064 ; n39065
g36630 nor n38499 n38608 ; n39066
g36631 and n39029 n39066 ; n39067
g36632 and n39031 n39067_not ; n39068
g36633 and n39065_not n39068 ; n39069
g36634 and n38888 n39069_not ; n39070
g36635 nor n39020 n39070 ; n39071
g36636 and pi0213_not n39071 ; n39072
g36637 nor pi1152 po1038 ; n39073
g36638 and n38413 n39029_not ; n39074
g36639 nor pi0299 n38937 ; n39075
g36640 nor pi1154 n39075 ; n39076
g36641 and n38765_not n39076 ; n39077
g36642 and n38731_not n39047 ; n39078
g36643 nor n39077 n39078 ; n39079
g36644 and pi0207 n39079 ; n39080
g36645 and n38722 n39080_not ; n39081
g36646 and pi0207_not n39079 ; n39082
g36647 and n38765_not n39053 ; n39083
g36648 and pi0207 n39083_not ; n39084
g36649 and pi0208 n39084_not ; n39085
g36650 and n39082_not n39085 ; n39086
g36651 nor n39081 n39086 ; n39087
g36652 and pi0211_not n39087 ; n39088
g36653 and pi0211 n39059 ; n39089
g36654 and n10843 n39088_not ; n39090
g36655 and n39089_not n39090 ; n39091
g36656 nor pi0211 n38787 ; n39092
g36657 and n39029 n39092 ; n39093
g36658 and pi0211 n39087 ; n39094
g36659 nor n38423 n39093 ; n39095
g36660 and n39094_not n39095 ; n39096
g36661 nor n39091 n39096 ; n39097
g36662 nor pi0219 n39097 ; n39098
g36663 and pi0211 n39029 ; n39099
g36664 and n38970 n39099_not ; n39100
g36665 and n39060_not n39100 ; n39101
g36666 nor n39074 n39101 ; n39102
g36667 and n39098_not n39102 ; n39103
g36668 and n39073 n39103_not ; n39104
g36669 and n38414_not n38966 ; n39105
g36670 and n38413_not n39007 ; n39106
g36671 nor n39105 n39106 ; n39107
g36672 and pi0219 n39107_not ; n39108
g36673 and pi0212_not n39013 ; n39109
g36674 and pi0211 n39006_not ; n39110
g36675 nor pi0199 pi1154 ; n39111
g36676 and pi0200_not n39111 ; n39112
g36677 and n38674 n39112 ; n39113
g36678 and n38722 n38943_not ; n39114
g36679 nor n38952 n39114 ; n39115
g36680 nor n38765 n39113 ; n39116
g36681 and n39115_not n39116 ; n39117
g36682 and pi0211_not n39117 ; n39118
g36683 and n10843 n39118_not ; n39119
g36684 and n39110_not n39119 ; n39120
g36685 nor pi0208 n38787 ; n39121
g36686 and n38995_not n39121 ; n39122
g36687 and pi0299 pi1156_not ; n39123
g36688 and n38998 n39123_not ; n39124
g36689 and n38787_not n38960 ; n39125
g36690 nor pi0207 n39125 ; n39126
g36691 and pi0208 n39124_not ; n39127
g36692 and n39126_not n39127 ; n39128
g36693 nor pi0211 n39122 ; n39129
g36694 and n39128_not n39129 ; n39130
g36695 and pi0211 n39117 ; n39131
g36696 nor n38423 n39130 ; n39132
g36697 and n39131_not n39132 ; n39133
g36698 nor pi0219 n39109 ; n39134
g36699 and n39133_not n39134 ; n39135
g36700 and n39120_not n39135 ; n39136
g36701 nor n39108 n39136 ; n39137
g36702 and pi1152 po1038_not ; n39138
g36703 and n39137_not n39138 ; n39139
g36704 nor n39104 n39139 ; n39140
g36705 and pi0213 n39140_not ; n39141
g36706 nor pi0209 n39141 ; n39142
g36707 and n39072_not n39142 ; n39143
g36708 nor n38935 n39143 ; n39144
g36709 and pi0219 n38495_not ; n39145
g36710 and pi0212 n38491_not ; n39146
g36711 and pi0214 n38485_not ; n39147
g36712 and pi0212_not n39147 ; n39148
g36713 nor pi0219 n39148 ; n39149
g36714 and n39146_not n39149 ; n39150
g36715 and pi0213 n39145_not ; n39151
g36716 and n38416 n39151 ; n39152
g36717 and n39150_not n39152 ; n39153
g36718 nor n39144 n39153 ; n39154
g36719 and pi0230 n39154_not ; n39155
g36720 and pi0230_not pi0234 ; n39156
g36721 or n39155 n39156 ; po0391
g36722 and pi0219 n38487_not ; n39158
g36723 and pi0219 n38608_not ; n39159
g36724 and pi0212_not n38481 ; n39160
g36725 nor pi0214 n38480 ; n39161
g36726 nor n39147 n39161 ; n39162
g36727 and pi0212 n39162_not ; n39163
g36728 nor pi0219 n39163 ; n39164
g36729 and n39160_not n39164 ; n39165
g36730 nor n39158 n39159 ; n39166
g36731 and po1038 n39166 ; n39167
g36732 and n39165_not n39167 ; n39168
g36733 and pi0208 pi1157 ; n39169
g36734 nor n38650 n38766 ; n39170
g36735 and pi0207 n39170_not ; n39171
g36736 nor pi0207 n38727 ; n39172
g36737 nor n39171 n39172 ; n39173
g36738 and n39169 n39173_not ; n39174
g36739 and pi0207_not n38734 ; n39175
g36740 nor n39171 n39175 ; n39176
g36741 and pi0208 n39176_not ; n39177
g36742 nor n38735 n39177 ; n39178
g36743 nor pi1157 n39178 ; n39179
g36744 nor n38730 n39174 ; n39180
g36745 and n39179_not n39180 ; n39181
g36746 and pi0211 n39181_not ; n39182
g36747 and pi1156_not n38577 ; n39183
g36748 nor n38698 n39183 ; n39184
g36749 and pi0207 n39184_not ; n39185
g36750 nor n38658 n38671 ; n39186
g36751 nor pi0207 n39186 ; n39187
g36752 nor n39185 n39187 ; n39188
g36753 and n39169 n39188_not ; n39189
g36754 and pi0207_not n38536 ; n39190
g36755 nor n39185 n39190 ; n39191
g36756 and pi0208 n39191_not ; n39192
g36757 nor n38786 n39192 ; n39193
g36758 nor pi1157 n39193 ; n39194
g36759 nor n38789 n39189 ; n39195
g36760 and n39194_not n39195 ; n39196
g36761 nor pi0211 n39196 ; n39197
g36762 and n10843 n39182_not ; n39198
g36763 and n39197_not n39198 ; n39199
g36764 and n10487 n38650_not ; n39200
g36765 and n39183_not n39200 ; n39201
g36766 nor pi0207 n38643 ; n39202
g36767 nor n39201 n39202 ; n39203
g36768 and n38645_not n39203 ; n39204
g36769 nor pi1157 n39204 ; n39205
g36770 and pi0207_not n38659 ; n39206
g36771 nor n39201 n39206 ; n39207
g36772 and n38661_not n39207 ; n39208
g36773 and pi1157 n39208_not ; n39209
g36774 nor n39205 n39209 ; n39210
g36775 and n38413 n39210_not ; n39211
g36776 and pi0211 n39196_not ; n39212
g36777 and pi0207_not n38672 ; n39213
g36778 and pi0208 n39213_not ; n39214
g36779 and n38698_not n38889 ; n39215
g36780 and n39214 n39215_not ; n39216
g36781 nor n38676 n39216 ; n39217
g36782 and pi1157 n39217 ; n39218
g36783 nor pi0211 n39205 ; n39219
g36784 and n39218_not n39219 ; n39220
g36785 and n38608 n39220_not ; n39221
g36786 and n39212_not n39221 ; n39222
g36787 nor n39211 n39222 ; n39223
g36788 and n39199_not n39223 ; n39224
g36789 nor pi0219 n39224 ; n39225
g36790 and pi0211_not n39181 ; n39226
g36791 and pi0211 n39210_not ; n39227
g36792 nor n38423 n39227 ; n39228
g36793 and n39226_not n39228 ; n39229
g36794 and n38423 n39210 ; n39230
g36795 and pi0219 n39230_not ; n39231
g36796 and n39229_not n39231 ; n39232
g36797 and pi0209 n39232_not ; n39233
g36798 and n39225_not n39233 ; n39234
g36799 and n38691_not n38722 ; n39235
g36800 and pi0207_not n38691 ; n39236
g36801 and pi0208 n39080_not ; n39237
g36802 and n39236_not n39237 ; n39238
g36803 nor n39235 n39238 ; n39239
g36804 and pi0211 n39239_not ; n39240
g36805 and n10487 n39024_not ; n39241
g36806 nor n38573 n38825 ; n39242
g36807 nor n10487 n39242 ; n39243
g36808 nor n39241 n39243 ; n39244
g36809 nor n38787 n39244 ; n39245
g36810 nor pi0211 n39245 ; n39246
g36811 and n10843 n39240_not ; n39247
g36812 and n39246_not n39247 ; n39248
g36813 and n38413 n39244_not ; n39249
g36814 and n38675 n38805_not ; n39250
g36815 and n38674 n38763 ; n39251
g36816 nor n39047 n39076 ; n39252
g36817 and pi0207 n39252 ; n39253
g36818 and pi0208 n39251_not ; n39254
g36819 and n39253_not n39254 ; n39255
g36820 nor n39250 n39255 ; n39256
g36821 and pi1157 n39256_not ; n39257
g36822 and pi1157_not n39244 ; n39258
g36823 nor pi0211 n39257 ; n39259
g36824 and n39258_not n39259 ; n39260
g36825 and pi0211 n39245 ; n39261
g36826 nor n39260 n39261 ; n39262
g36827 and n38608 n39262_not ; n39263
g36828 nor n39248 n39249 ; n39264
g36829 and n39263_not n39264 ; n39265
g36830 nor pi0219 n39265 ; n39266
g36831 and pi0211_not n39239 ; n39267
g36832 and pi0211 n39244_not ; n39268
g36833 nor n38423 n39268 ; n39269
g36834 and n39267_not n39269 ; n39270
g36835 and n38423 n39244 ; n39271
g36836 and pi0219 n39271_not ; n39272
g36837 and n39270_not n39272 ; n39273
g36838 nor pi0209 n39273 ; n39274
g36839 and n39266_not n39274 ; n39275
g36840 nor n39234 n39275 ; n39276
g36841 nor po1038 n39276 ; n39277
g36842 and pi0213 n39168_not ; n39278
g36843 and n39277_not n39278 ; n39279
g36844 and pi0219 n38497_not ; n39280
g36845 and po1038 n39280_not ; n39281
g36846 and n38489_not n38608 ; n39282
g36847 and n10843 n38883_not ; n39283
g36848 nor pi0219 n39282 ; n39284
g36849 and n39283_not n39284 ; n39285
g36850 and n39159_not n39281 ; n39286
g36851 and n39285_not n39286 ; n39287
g36852 and pi1157 n39217_not ; n39288
g36853 and pi0299 pi1157_not ; n39289
g36854 nor n39194 n39289 ; n39290
g36855 and n39288_not n39290 ; n39291
g36856 nor n38769 n39291 ; n39292
g36857 nor pi0211 n39292 ; n39293
g36858 and n39228 n39293_not ; n39294
g36859 and n39231 n39294_not ; n39295
g36860 nor n38578 n38767 ; n39296
g36861 nor n38650 n39296 ; n39297
g36862 and pi0207 n39297_not ; n39298
g36863 and pi1154 n38535_not ; n39299
g36864 nor n38642 n39299 ; n39300
g36865 nor pi0207 n38732 ; n39301
g36866 and n39300_not n39301 ; n39302
g36867 nor n39298 n39302 ; n39303
g36868 and pi0208 n39303_not ; n39304
g36869 nor n38757 n39304 ; n39305
g36870 nor pi1157 n39305 ; n39306
g36871 and n38746 n39217_not ; n39307
g36872 nor n39306 n39307 ; n39308
g36873 nor pi0211 n39308 ; n39309
g36874 and pi0211 n39292 ; n39310
g36875 and n10843 n39309_not ; n39311
g36876 and n39310_not n39311 ; n39312
g36877 and pi0211 n39308 ; n39313
g36878 nor n39226 n39313 ; n39314
g36879 and n38608 n39314_not ; n39315
g36880 nor n39211 n39315 ; n39316
g36881 and n39312_not n39316 ; n39317
g36882 nor pi0219 n39317 ; n39318
g36883 nor n39295 n39318 ; n39319
g36884 and pi0209 n39319_not ; n39320
g36885 nor n38764 n38975 ; n39321
g36886 nor pi0208 n39321 ; n39322
g36887 nor pi0207 n38763 ; n39323
g36888 nor n39035 n39323 ; n39324
g36889 and pi0208 n39324_not ; n39325
g36890 nor n39322 n39325 ; n39326
g36891 and pi0211_not n39326 ; n39327
g36892 and n39269 n39327_not ; n39328
g36893 and n39272 n39328_not ; n39329
g36894 nor n38753 n38836 ; n39330
g36895 nor pi0208 n39330 ; n39331
g36896 nor pi0207 n38752 ; n39332
g36897 nor n39049 n39332 ; n39333
g36898 and pi0208 n39333_not ; n39334
g36899 nor n39331 n39334 ; n39335
g36900 and pi0211 n39335 ; n39336
g36901 nor n39267 n39336 ; n39337
g36902 nor n38423 n39337 ; n39338
g36903 nor pi0211 n39335 ; n39339
g36904 and pi0211 n39326_not ; n39340
g36905 and n10843 n39340_not ; n39341
g36906 and n39339_not n39341 ; n39342
g36907 nor n39249 n39342 ; n39343
g36908 and n39338_not n39343 ; n39344
g36909 nor pi0219 n39344 ; n39345
g36910 nor n39329 n39345 ; n39346
g36911 nor pi0209 n39346 ; n39347
g36912 nor po1038 n39347 ; n39348
g36913 and n39320_not n39348 ; n39349
g36914 nor pi0213 n39287 ; n39350
g36915 and n39349_not n39350 ; n39351
g36916 nor n39279 n39351 ; n39352
g36917 and pi0230 n39352_not ; n39353
g36918 nor pi0230 pi0235 ; n39354
g36919 nor n39353 n39354 ; po0392
g36920 and pi0100_not n38198 ; n39356
g36921 and n38397 n39356_not ; n39357
g36922 nor n6132 n39357 ; n39358
g36923 nor pi0075 n39358 ; n39359
g36924 nor n7302 n39359 ; n39360
g36925 nor pi0092 n39360 ; n39361
g36926 and n13654 n39361_not ; n39362
g36927 nor pi0074 n39362 ; n39363
g36928 and n6131 n39363_not ; n39364
g36929 nor pi0056 n39364 ; n39365
g36930 nor n6127 n39365 ; n39366
g36931 nor pi0062 n39366 ; n39367
g36932 and n13662 n39367_not ; po0393
g36933 and pi0211 pi1157 ; n39369
g36934 and pi0211_not pi1158 ; n39370
g36935 nor n39369 n39370 ; n39371
g36936 and n38421 n39371_not ; n39372
g36937 and n39164 n39372_not ; n39373
g36938 and pi0219_not po1038 ; n39374
g36939 and n38421 n38483 ; n39375
g36940 and po1038 n39375 ; n39376
g36941 nor n39374 n39376 ; n39377
g36942 and pi0214 n38495 ; n39378
g36943 and pi1155 n38744 ; n39379
g36944 nor n39378 n39379 ; n39380
g36945 and pi0212 n39380_not ; n39381
g36946 and po1038 n39381 ; n39382
g36947 and n39377 n39382_not ; n39383
g36948 nor n39373 n39383 ; n39384
g36949 nor pi0213 n39384 ; n39385
g36950 and n38508 n39373_not ; n39386
g36951 and pi0199 pi1143 ; n39387
g36952 nor pi0200 n39387 ; n39388
g36953 and n38434_not n39388 ; n39389
g36954 and n38437_not n39026 ; n39390
g36955 and n39389_not n39390 ; n39391
g36956 and pi0200 n38434_not ; n39392
g36957 and pi0199_not pi1145 ; n39393
g36958 and n39388 n39393_not ; n39394
g36959 and n38826 n39392_not ; n39395
g36960 and n39394_not n39395 ; n39396
g36961 nor n39391 n39396 ; n39397
g36962 nor pi0299 n39397 ; n39398
g36963 and n38421 n38787 ; n39399
g36964 and pi0214 n38514_not ; n39400
g36965 nor pi0214 n38510 ; n39401
g36966 and pi0212 n39400_not ; n39402
g36967 and n39401_not n39402 ; n39403
g36968 nor n39399 n39403 ; n39404
g36969 and n38519 n39404_not ; n39405
g36970 nor n39398 n39405 ; n39406
g36971 and n39386_not n39406 ; n39407
g36972 nor po1038 n39407 ; n39408
g36973 and n39385 n39408_not ; n39409
g36974 and pi0219 n38425_not ; n39410
g36975 and n10843 n38420 ; n39411
g36976 and pi0211_not pi1145 ; n39412
g36977 and pi0211 pi1144 ; n39413
g36978 nor n39412 n39413 ; n39414
g36979 and n10843_not n39414 ; n39415
g36980 nor n38413 n39411 ; n39416
g36981 and n39415_not n39416 ; n39417
g36982 nor pi0219 n39417 ; n39418
g36983 and n38416 n39410_not ; n39419
g36984 and n39418_not n39419 ; n39420
g36985 and n38508 n39417 ; n39421
g36986 and pi0299 n38970 ; n39422
g36987 and n38425 n39422 ; n39423
g36988 nor n39398 n39423 ; n39424
g36989 and n39421_not n39424 ; n39425
g36990 nor po1038 n39425 ; n39426
g36991 nor n39420 n39426 ; n39427
g36992 and pi0213 n39427 ; n39428
g36993 and pi0209 n39409_not ; n39429
g36994 and n39428_not n39429 ; n39430
g36995 and n38449 n38568 ; n39431
g36996 and pi1158 n38955 ; n39432
g36997 nor pi0199 pi1158 ; n39433
g36998 and pi1156 n39433_not ; n39434
g36999 nor n39432 n39434 ; n39435
g37000 and n39431 n39435_not ; n39436
g37001 and pi0207 n38651 ; n39437
g37002 and pi0208 n39202_not ; n39438
g37003 and n39437_not n39438 ; n39439
g37004 nor n39436 n39439 ; n39440
g37005 nor pi1157 n39440 ; n39441
g37006 and pi1156 n38699 ; n39442
g37007 nor pi0200 pi1158 ; n39443
g37008 nor pi0199 n39443 ; n39444
g37009 nor n39442 n39444 ; n39445
g37010 and n38441 n39445_not ; n39446
g37011 and pi0208_not n39446 ; n39447
g37012 and pi0208 n39206_not ; n39448
g37013 and n39437_not n39448 ; n39449
g37014 nor n39447 n39449 ; n39450
g37015 and pi1157 n39450_not ; n39451
g37016 nor n39441 n39451 ; n39452
g37017 and n38414_not n39452 ; n39453
g37018 and pi0200_not pi0207 ; n39454
g37019 and n39435_not n39454 ; n39455
g37020 nor pi1157 n39455 ; n39456
g37021 and pi1156 n38985_not ; n39457
g37022 nor pi1158 n38641 ; n39458
g37023 and n39457 n39458_not ; n39459
g37024 nor n39444 n39459 ; n39460
g37025 and n38441 n39460_not ; n39461
g37026 nor pi0208 n39456 ; n39462
g37027 and n39461 n39462 ; n39463
g37028 nor pi0208 n39463 ; n39464
g37029 and n38543_not n39464 ; n39465
g37030 nor pi0299 n38536 ; n39466
g37031 and pi0200_not pi1157 ; n39467
g37032 and pi0199_not n39467 ; n39468
g37033 and n39466 n39468_not ; n39469
g37034 nor pi0207 n38528 ; n39470
g37035 and n39469_not n39470 ; n39471
g37036 and pi0207 n38601_not ; n39472
g37037 and pi0208 n39471_not ; n39473
g37038 and n39472_not n39473 ; n39474
g37039 nor n39465 n39474 ; n39475
g37040 and n38414 n39475_not ; n39476
g37041 nor n39453 n39476 ; n39477
g37042 and pi0219 n39477_not ; n39478
g37043 and pi0214_not n39452 ; n39479
g37044 nor pi0212 n39479 ; n39480
g37045 and pi0299 pi1145_not ; n39481
g37046 nor pi0207 n39481 ; n39482
g37047 and n39469_not n39482 ; n39483
g37048 and pi0299 pi1145 ; n39484
g37049 and n38578 n39484_not ; n39485
g37050 nor n38702 n39481 ; n39486
g37051 and pi1154 n39486_not ; n39487
g37052 nor pi1156 n39485 ; n39488
g37053 and n39487_not n39488 ; n39489
g37054 and n38593 n39484_not ; n39490
g37055 nor n38596 n39481 ; n39491
g37056 nor pi1154 n39491 ; n39492
g37057 and pi1156 n39490_not ; n39493
g37058 and n39492_not n39493 ; n39494
g37059 nor n39489 n39494 ; n39495
g37060 and pi0207 n39495_not ; n39496
g37061 and pi0208 n39483_not ; n39497
g37062 and n39496_not n39497 ; n39498
g37063 and n38641 n38725_not ; n39499
g37064 and pi1157 n39432_not ; n39500
g37065 and n39499_not n39500 ; n39501
g37066 and pi0207 n39501_not ; n39502
g37067 and pi0299_not n39442 ; n39503
g37068 nor pi1157 n39432 ; n39504
g37069 and n39503_not n39504 ; n39505
g37070 and n39502 n39505_not ; n39506
g37071 nor pi0208 n39484 ; n39507
g37072 and n39506_not n39507 ; n39508
g37073 nor n39498 n39508 ; n39509
g37074 nor pi0211 n39509 ; n39510
g37075 and n38612_not n39464 ; n39511
g37076 nor pi0207 n38610 ; n39512
g37077 and n39469_not n39512 ; n39513
g37078 and pi0207 n38630_not ; n39514
g37079 and pi0208 n39513_not ; n39515
g37080 and n39514_not n39515 ; n39516
g37081 nor n39511 n39516 ; n39517
g37082 and pi0211 n39517_not ; n39518
g37083 nor n39510 n39518 ; n39519
g37084 and pi0214 n39519_not ; n39520
g37085 and n39480 n39520_not ; n39521
g37086 and pi0211_not n39517 ; n39522
g37087 and pi0211 n39475 ; n39523
g37088 and pi0214 n39522_not ; n39524
g37089 and n39523_not n39524 ; n39525
g37090 nor pi0214 n39519 ; n39526
g37091 and pi0212 n39525_not ; n39527
g37092 and n39526_not n39527 ; n39528
g37093 nor pi0219 n39521 ; n39529
g37094 and n39528_not n39529 ; n39530
g37095 nor po1038 n39478 ; n39531
g37096 and n39530_not n39531 ; n39532
g37097 and pi0213 n39420_not ; n39533
g37098 and n39532_not n39533 ; n39534
g37099 nor n38853 n39187 ; n39535
g37100 and n39169 n39535_not ; n39536
g37101 nor n38787 n39446 ; n39537
g37102 and n38542 n39537_not ; n39538
g37103 and n39121 n39455_not ; n39539
g37104 and pi0208 n39190_not ; n39540
g37105 and n38853_not n39540 ; n39541
g37106 nor pi1157 n39539 ; n39542
g37107 and n39541_not n39542 ; n39543
g37108 nor n39536 n39538 ; n39544
g37109 and n39543_not n39544 ; n39545
g37110 and n38421 n39545 ; n39546
g37111 and pi0207 n38860_not ; n39547
g37112 nor n39172 n39547 ; n39548
g37113 and n39169 n39548_not ; n39549
g37114 nor n38510 n39461 ; n39550
g37115 and n38542 n39550_not ; n39551
g37116 nor n39175 n39547 ; n39552
g37117 and pi0208 n39552_not ; n39553
g37118 and pi0208_not n38510 ; n39554
g37119 nor n39436 n39554 ; n39555
g37120 and n39553_not n39555 ; n39556
g37121 nor pi1157 n39556 ; n39557
g37122 nor n39549 n39551 ; n39558
g37123 and n39557_not n39558 ; n39559
g37124 nor pi0214 n39559 ; n39560
g37125 nor pi0207 n38672 ; n39561
g37126 and n38745_not n39561 ; n39562
g37127 and pi1157 n39562_not ; n39563
g37128 nor pi1157 n39436 ; n39564
g37129 and n39302_not n39564 ; n39565
g37130 nor n39563 n39565 ; n39566
g37131 and pi0208 n38837_not ; n39567
g37132 and n39566_not n39567 ; n39568
g37133 and n39461 n39564_not ; n39569
g37134 nor pi0208 n38514 ; n39570
g37135 and n39569_not n39570 ; n39571
g37136 and pi0214 n39571_not ; n39572
g37137 and n39568_not n39572 ; n39573
g37138 and pi0212 n39573_not ; n39574
g37139 and n39560_not n39574 ; n39575
g37140 nor n39546 n39575 ; n39576
g37141 nor pi0211 n39576 ; n39577
g37142 nor n39453 n39577 ; n39578
g37143 and pi0219 n39578_not ; n39579
g37144 and pi0299_not n39445 ; n39580
g37145 and n38675 n39580_not ; n39581
g37146 and n38890_not n39214 ; n39582
g37147 nor n39581 n39582 ; n39583
g37148 and pi1157 n39583_not ; n39584
g37149 nor n39441 n39584 ; n39585
g37150 and pi0211 n39585 ; n39586
g37151 and n38441 n39442 ; n39587
g37152 nor pi0299 n39039 ; n39588
g37153 and pi1158 n39588_not ; n39589
g37154 nor pi0208 n39587 ; n39590
g37155 and n39589_not n39590 ; n39591
g37156 and pi1158_not n38651 ; n39592
g37157 and pi1158 n38768 ; n39593
g37158 and pi0207 n39592_not ; n39594
g37159 and n39593_not n39594 ; n39595
g37160 and pi0299 pi1158_not ; n39596
g37161 nor pi0207 n39596 ; n39597
g37162 and n39466_not n39597 ; n39598
g37163 and pi0208 n39598_not ; n39599
g37164 and n39595_not n39599 ; n39600
g37165 nor pi1157 n39591 ; n39601
g37166 and n39600_not n39601 ; n39602
g37167 and n39561 n39596_not ; n39603
g37168 nor n39595 n39603 ; n39604
g37169 and n39169 n39604_not ; n39605
g37170 nor n39502 n39589 ; n39606
g37171 and n38542 n39606_not ; n39607
g37172 nor pi0211 n39607 ; n39608
g37173 and n39602_not n39608 ; n39609
g37174 and n39605_not n39609 ; n39610
g37175 nor n39586 n39610 ; n39611
g37176 and pi0214 n39611_not ; n39612
g37177 and n39480 n39612_not ; n39613
g37178 and n38783 n39545_not ; n39614
g37179 and n10484 n39559_not ; n39615
g37180 and n38744 n39585_not ; n39616
g37181 nor n39614 n39615 ; n39617
g37182 and n39616_not n39617 ; n39618
g37183 and pi0212 n39618_not ; n39619
g37184 nor pi0219 n39619 ; n39620
g37185 and n39613_not n39620 ; n39621
g37186 nor po1038 n39579 ; n39622
g37187 and n39621_not n39622 ; n39623
g37188 and n39385 n39623_not ; n39624
g37189 nor pi0209 n39534 ; n39625
g37190 and n39624_not n39625 ; n39626
g37191 nor n39430 n39626 ; n39627
g37192 and pi0230 n39627_not ; n39628
g37193 nor pi0230 pi0237 ; n39629
g37194 or n39628 n39629 ; po0394
g37195 nor pi0211 pi1153 ; n39631
g37196 and pi0219 n39631 ; n39632
g37197 and n38416 n39632_not ; n39633
g37198 and n39285_not n39633 ; n39634
g37199 nor pi1151 po1038 ; n39635
g37200 and n10809 n38826 ; n39636
g37201 nor pi0299 n39636 ; n39637
g37202 nor n13061 n39637 ; n39638
g37203 and n38826 n38955 ; n39639
g37204 nor pi0214 n39639 ; n39640
g37205 and pi0212_not n39640 ; n39641
g37206 and n39638 n39641_not ; n39642
g37207 and pi1153 n39642 ; n39643
g37208 nor n38665 n39643 ; n39644
g37209 and n38882 n39637_not ; n39645
g37210 and pi1153 n39639 ; n39646
g37211 nor n38514 n39646 ; n39647
g37212 nor pi0211 n39647 ; n39648
g37213 and n10843 n39645_not ; n39649
g37214 and n39648_not n39649 ; n39650
g37215 and pi0299 n38489_not ; n39651
g37216 nor n38423 n39651 ; n39652
g37217 and n39646_not n39652 ; n39653
g37218 nor n39650 n39653 ; n39654
g37219 nor pi0219 n39654 ; n39655
g37220 and n39635 n39644_not ; n39656
g37221 and n39655_not n39656 ; n39657
g37222 and n10487_not n38568 ; n39658
g37223 and n38825_not n39658 ; n39659
g37224 and n38561 n39026 ; n39660
g37225 nor n39659 n39660 ; n39661
g37226 nor n38962 n39661 ; n39662
g37227 nor pi0214 n39662 ; n39663
g37228 nor pi0212 n39663 ; n39664
g37229 and n38568 n38958_not ; n39665
g37230 nor pi1153 n38700 ; n39666
g37231 nor n38682 n39666 ; n39667
g37232 and pi1155 n39667_not ; n39668
g37233 nor n39665 n39668 ; n39669
g37234 and n38441 n38561_not ; n39670
g37235 and pi0208 n39670_not ; n39671
g37236 nor n38722 n39671 ; n39672
g37237 nor n39669 n39672 ; n39673
g37238 nor n39660 n39673 ; n39674
g37239 nor pi0299 n39674 ; n39675
g37240 and pi0214 n39651_not ; n39676
g37241 and n39675_not n39676 ; n39677
g37242 and n39664 n39677_not ; n39678
g37243 and n38514_not n38783 ; n39679
g37244 and n39662_not n39679 ; n39680
g37245 and n38744 n39674 ; n39681
g37246 nor pi0299 n39454 ; n39682
g37247 nor pi0208 n39682 ; n39683
g37248 and pi0200 n38674 ; n39684
g37249 and n39671 n39684_not ; n39685
g37250 nor n39683 n39685 ; n39686
g37251 nor n38683 n39686 ; n39687
g37252 and n10484 n39687_not ; n39688
g37253 and pi0212 n39680_not ; n39689
g37254 and n39688_not n39689 ; n39690
g37255 and n39681_not n39690 ; n39691
g37256 nor pi0219 n39691 ; n39692
g37257 and n39678_not n39692 ; n39693
g37258 and pi1151 po1038_not ; n39694
g37259 nor pi0211 n39686 ; n39695
g37260 and pi0211 n39661_not ; n39696
g37261 nor n39695 n39696 ; n39697
g37262 nor n38683 n39697 ; n39698
g37263 and n38413 n39662_not ; n39699
g37264 and n39698 n39699_not ; n39700
g37265 and pi0219 n39700_not ; n39701
g37266 and n39694 n39701_not ; n39702
g37267 and n39693_not n39702 ; n39703
g37268 nor pi1152 n39657 ; n39704
g37269 and n39703_not n39704 ; n39705
g37270 nor n11445 n39045 ; n39706
g37271 and pi0207 n39706_not ; n39707
g37272 nor n38975 n39707 ; n39708
g37273 nor pi0208 n39708 ; n39709
g37274 and pi0200 pi0207 ; n39710
g37275 nor pi0199 n39710 ; n39711
g37276 nor pi0299 n39711 ; n39712
g37277 and pi0208 n39712_not ; n39713
g37278 and pi0207_not n10809 ; n39714
g37279 nor pi0299 n39714 ; n39715
g37280 nor pi1153 n39715 ; n39716
g37281 and n39713 n39716_not ; n39717
g37282 nor n39709 n39717 ; n39718
g37283 and pi0211 n39718_not ; n39719
g37284 nor pi0207 n38947 ; n39720
g37285 nor n39039 n39720 ; n39721
g37286 and pi0208 n39721_not ; n39722
g37287 and n38675 n38947_not ; n39723
g37288 nor n39722 n39723 ; n39724
g37289 nor pi0211 n38745 ; n39725
g37290 and n39724_not n39725 ; n39726
g37291 nor n39719 n39726 ; n39727
g37292 and n10843 n39727_not ; n39728
g37293 and pi0299 n38489 ; n39729
g37294 nor n38423 n39724 ; n39730
g37295 and n39729_not n39730 ; n39731
g37296 nor n39728 n39731 ; n39732
g37297 nor pi0219 n39732 ; n39733
g37298 and n10487_not n38945 ; n39734
g37299 nor n38826 n39454 ; n39735
g37300 and n11384 n39735_not ; n39736
g37301 and n39734_not n39736 ; n39737
g37302 and pi0211_not n38512 ; n39738
g37303 and n38413_not n39738 ; n39739
g37304 nor n39737 n39739 ; n39740
g37305 nor n38665 n39740 ; n39741
g37306 nor n39733 n39741 ; n39742
g37307 and n39635 n39742_not ; n39743
g37308 and n38441 n38561 ; n39744
g37309 and pi0208 n38550 ; n39745
g37310 and n39714_not n39745 ; n39746
g37311 nor n39744 n39746 ; n39747
g37312 and pi0214_not n39747 ; n39748
g37313 and n39646_not n39748 ; n39749
g37314 nor pi0212 n39749 ; n39750
g37315 and pi0214_not n39750 ; n39751
g37316 and n38948 n38986_not ; n39752
g37317 and pi0208 n39752_not ; n39753
g37318 and n38675 n38949_not ; n39754
g37319 nor n39753 n39754 ; n39755
g37320 nor pi0211 n39755 ; n39756
g37321 and n38765_not n39756 ; n39757
g37322 and pi0211 n39755_not ; n39758
g37323 and n38745_not n39758 ; n39759
g37324 nor n39757 n39759 ; n39760
g37325 nor n38423 n39760 ; n39761
g37326 and n39645_not n39747 ; n39762
g37327 and n39726_not n39762 ; n39763
g37328 and n10843 n39763_not ; n39764
g37329 nor pi0219 n39751 ; n39765
g37330 and n39764_not n39765 ; n39766
g37331 and n39761_not n39766 ; n39767
g37332 and pi0219 n39747 ; n39768
g37333 and n39643_not n39768 ; n39769
g37334 and n39694 n39769_not ; n39770
g37335 and n39767_not n39770 ; n39771
g37336 and pi1152 n39771_not ; n39772
g37337 and n39743_not n39772 ; n39773
g37338 nor n39705 n39773 ; n39774
g37339 nor pi0209 n39774 ; n39775
g37340 and n38641 n39032 ; n39776
g37341 and n10487 n39776_not ; n39777
g37342 and n38957_not n39777 ; n39778
g37343 nor n39243 n39778 ; n39779
g37344 nor pi0214 n39779 ; n39780
g37345 and pi0212_not n39780 ; n39781
g37346 and pi0211 n39779 ; n39782
g37347 and pi1153 n38581_not ; n39783
g37348 nor n38957 n39783 ; n39784
g37349 and pi0207 n39784_not ; n39785
g37350 nor n39323 n39785 ; n39786
g37351 and pi0208 n39786_not ; n39787
g37352 nor n39322 n39787 ; n39788
g37353 nor pi0211 n39788 ; n39789
g37354 nor n39782 n39789 ; n39790
g37355 and n38970 n39790 ; n39791
g37356 and n38550_not n39084 ; n39792
g37357 nor pi1154 n39052 ; n39793
g37358 and n38581_not n39793 ; n39794
g37359 and pi0207 n39794_not ; n39795
g37360 and n39001 n39795 ; n39796
g37361 and pi0208 n39796_not ; n39797
g37362 and n39792_not n39797 ; n39798
g37363 and n39236_not n39798 ; n39799
g37364 nor n39235 n39799 ; n39800
g37365 nor pi0211 n39800 ; n39801
g37366 and n39001 n39776_not ; n39802
g37367 and pi0207 n39802_not ; n39803
g37368 nor n39332 n39803 ; n39804
g37369 and pi0208 n39804_not ; n39805
g37370 nor n39331 n39805 ; n39806
g37371 and pi0211 n39806_not ; n39807
g37372 and n38421 n39801_not ; n39808
g37373 and n39807_not n39808 ; n39809
g37374 and n10484 n39788_not ; n39810
g37375 and n38744 n39800_not ; n39811
g37376 and n38783 n39806_not ; n39812
g37377 and pi0212 n39810_not ; n39813
g37378 and n39811_not n39813 ; n39814
g37379 and n39812_not n39814 ; n39815
g37380 nor n39809 n39815 ; n39816
g37381 nor pi0219 n39816 ; n39817
g37382 nor po1038 n39781 ; n39818
g37383 and n39791_not n39818 ; n39819
g37384 and n39817_not n39819 ; n39820
g37385 and pi0209 n39820_not ; n39821
g37386 nor n39775 n39821 ; n39822
g37387 nor n39634 n39822 ; n39823
g37388 and pi0213 n39823_not ; n39824
g37389 and pi0211_not n38608 ; n39825
g37390 and pi1153 n39825 ; n39826
g37391 and n39374 n39826 ; n39827
g37392 nor pi1151 n39827 ; n39828
g37393 and pi0219 n39639_not ; n39829
g37394 nor po1038 n39829 ; n39830
g37395 nor n13061 n39646 ; n39831
g37396 and pi0212 n39640_not ; n39832
g37397 and n39831_not n39832 ; n39833
g37398 nor pi0219 n39833 ; n39834
g37399 and n39640 n39643 ; n39835
g37400 and n38421 n39738 ; n39836
g37401 nor n39639 n39836 ; n39837
g37402 and n39834 n39837 ; n39838
g37403 and n39835_not n39838 ; n39839
g37404 and n39643 n39830 ; n39840
g37405 and n39839_not n39840 ; n39841
g37406 and n39828 n39841_not ; n39842
g37407 and n10486 n39826_not ; n39843
g37408 and n38416 n39843_not ; n39844
g37409 and pi1151 n39844_not ; n39845
g37410 and pi0214_not n39698 ; n39846
g37411 and n39662_not n39831 ; n39847
g37412 and pi0214 n39847_not ; n39848
g37413 and pi0212 n39848_not ; n39849
g37414 and n39846_not n39849 ; n39850
g37415 nor pi0212 n39700 ; n39851
g37416 nor n39850 n39851 ; n39852
g37417 nor pi0219 n39852 ; n39853
g37418 and pi0211_not pi0299 ; n39854
g37419 nor n39646 n39854 ; n39855
g37420 and n39662_not n39855 ; n39856
g37421 nor n39699 n39856 ; n39857
g37422 and pi0219 n39857_not ; n39858
g37423 nor po1038 n39858 ; n39859
g37424 and n39853_not n39859 ; n39860
g37425 and n39845 n39860_not ; n39861
g37426 nor pi1152 n39842 ; n39862
g37427 and n39861_not n39862 ; n39863
g37428 and n10485_not n38665 ; n39864
g37429 and po1038 n39864 ; n39865
g37430 nor n10843 n39631 ; n39866
g37431 nor n38527 n39866 ; n39867
g37432 and n39865 n39867_not ; n39868
g37433 and n10486_not n38416 ; n39869
g37434 and pi1151 n39869_not ; n39870
g37435 and n39868_not n39870 ; n39871
g37436 and n39646_not n39747 ; n39872
g37437 and n39756_not n39872 ; n39873
g37438 and pi0214 n39873 ; n39874
g37439 nor n39749 n39874 ; n39875
g37440 nor pi0212 n39875 ; n39876
g37441 nor n39873 n39876 ; n39877
g37442 and pi0219 n39877_not ; n39878
g37443 nor po1038 n39878 ; n39879
g37444 and pi1153 n39637_not ; n39880
g37445 nor n39758 n39880 ; n39881
g37446 and pi0214 n39747 ; n39882
g37447 and n39881 n39882 ; n39883
g37448 and n39750 n39883_not ; n39884
g37449 and pi0214 n39755 ; n39885
g37450 and n39748 n39881 ; n39886
g37451 and pi0212 n39885_not ; n39887
g37452 and n39886_not n39887 ; n39888
g37453 nor pi0219 n39884 ; n39889
g37454 and n39888_not n39889 ; n39890
g37455 and n39879 n39890_not ; n39891
g37456 and n39871 n39891_not ; n39892
g37457 nor pi1151 n39868 ; n39893
g37458 and pi0219 n39737_not ; n39894
g37459 nor po1038 n39894 ; n39895
g37460 and pi0211_not n39718 ; n39896
g37461 and n39730 n39896_not ; n39897
g37462 and n38608_not n39737 ; n39898
g37463 and pi0299 n38527 ; n39899
g37464 nor pi0219 n39899 ; n39900
g37465 and n39898_not n39900 ; n39901
g37466 and n39897_not n39901 ; n39902
g37467 and n39895 n39902_not ; n39903
g37468 and n39893 n39903_not ; n39904
g37469 and pi1152 n39904_not ; n39905
g37470 and n39892_not n39905 ; n39906
g37471 nor n39863 n39906 ; n39907
g37472 and pi0209_not n39907 ; n39908
g37473 and pi0219_not n38608 ; n39909
g37474 nor n39779 n39909 ; n39910
g37475 and n39790 n39909 ; n39911
g37476 nor po1038 n39910 ; n39912
g37477 and n39911_not n39912 ; n39913
g37478 and n39828 n39913_not ; n39914
g37479 and n39251_not n39797 ; n39915
g37480 nor n39250 n39915 ; n39916
g37481 nor pi0211 n39916 ; n39917
g37482 nor n39782 n39917 ; n39918
g37483 and n38413_not n39918 ; n39919
g37484 nor n39781 n39919 ; n39920
g37485 and pi0219 n39920_not ; n39921
g37486 nor po1038 n39921 ; n39922
g37487 and pi0214 n39790 ; n39923
g37488 nor n39780 n39923 ; n39924
g37489 nor pi0212 n39924 ; n39925
g37490 nor pi0214 n39790 ; n39926
g37491 and pi0211 n39916_not ; n39927
g37492 and pi0211_not n39779 ; n39928
g37493 nor n39927 n39928 ; n39929
g37494 and pi0214 n39929_not ; n39930
g37495 and pi0212 n39926_not ; n39931
g37496 and n39930_not n39931 ; n39932
g37497 nor n39925 n39932 ; n39933
g37498 nor pi0219 n39933 ; n39934
g37499 and n39922 n39934_not ; n39935
g37500 and n39845 n39935_not ; n39936
g37501 nor pi1152 n39914 ; n39937
g37502 and n39936_not n39937 ; n39938
g37503 nor n39789 n39927 ; n39939
g37504 nor pi0214 n39939 ; n39940
g37505 and pi0214 n39918_not ; n39941
g37506 nor n39940 n39941 ; n39942
g37507 and pi0212 n39942_not ; n39943
g37508 and pi0214 n39939 ; n39944
g37509 nor pi0212 n39780 ; n39945
g37510 and n39944_not n39945 ; n39946
g37511 nor pi0219 n39946 ; n39947
g37512 and n39943_not n39947 ; n39948
g37513 and pi0219 n39779_not ; n39949
g37514 nor po1038 n39949 ; n39950
g37515 and n39948_not n39950 ; n39951
g37516 and n39893 n39951_not ; n39952
g37517 and pi0214 n39916_not ; n39953
g37518 nor n39940 n39953 ; n39954
g37519 and pi0212 n39954_not ; n39955
g37520 and n39947 n39955_not ; n39956
g37521 and n39922 n39956_not ; n39957
g37522 and n39871 n39957_not ; n39958
g37523 and pi1152 n39952_not ; n39959
g37524 and n39958_not n39959 ; n39960
g37525 and pi0209 n39938_not ; n39961
g37526 and n39960_not n39961 ; n39962
g37527 nor pi0213 n39908 ; n39963
g37528 and n39962_not n39963 ; n39964
g37529 nor n39824 n39964 ; n39965
g37530 and pi0230 n39965_not ; n39966
g37531 and pi0230_not pi0238 ; n39967
g37532 or n39966 n39967 ; po0395
g37533 and n38449 n38651_not ; n39969
g37534 and pi0212 n39969_not ; n39970
g37535 nor po1038 n39970 ; n39971
g37536 and pi0214_not n39969 ; n39972
g37537 nor pi0212 n39972 ; n39973
g37538 and pi0219_not n39973 ; n39974
g37539 and pi0299 pi1158 ; n39975
g37540 and n38449_not n39975 ; n39976
g37541 and pi0208_not n39595 ; n39977
g37542 nor n39976 n39977 ; n39978
g37543 nor pi0211 n39978 ; n39979
g37544 nor pi1157 n39969 ; n39980
g37545 and pi0208 pi0299 ; n39981
g37546 and pi1157 n39981_not ; n39982
g37547 and n38891_not n39982 ; n39983
g37548 and pi0211 n39980_not ; n39984
g37549 and n39983_not n39984 ; n39985
g37550 nor n39979 n39985 ; n39986
g37551 and pi0214 n39986_not ; n39987
g37552 and n39974 n39987_not ; n39988
g37553 and pi0219 n39973 ; n39989
g37554 and pi0211 n39969_not ; n39990
g37555 and pi0214 n39990_not ; n39991
g37556 and n38855_not n39092 ; n39992
g37557 and n39991 n39992_not ; n39993
g37558 and n39989 n39993_not ; n39994
g37559 and pi0209_not n39971 ; n39995
g37560 and n39994_not n39995 ; n39996
g37561 and n39988_not n39996 ; n39997
g37562 nor pi0219 n39372 ; n39998
g37563 nor n39377 n39998 ; n39999
g37564 and n39447 n39564_not ; n40000
g37565 and pi0214_not n40000 ; n40001
g37566 nor pi0212 n40001 ; n40002
g37567 and pi0219_not n40002 ; n40003
g37568 and n39581_not n39982 ; n40004
g37569 nor n39564 n40004 ; n40005
g37570 and pi0211 n40005_not ; n40006
g37571 and pi0208 n39975_not ; n40007
g37572 nor n38542 n40007 ; n40008
g37573 and n39591_not n40008 ; n40009
g37574 and n39608 n40009_not ; n40010
g37575 and pi0214 n40006_not ; n40011
g37576 and n40010_not n40011 ; n40012
g37577 and n40003 n40012_not ; n40013
g37578 and pi0212 n40000_not ; n40014
g37579 nor po1038 n40014 ; n40015
g37580 and pi0219 n40002 ; n40016
g37581 and pi0211 n40000_not ; n40017
g37582 and n39092 n40000_not ; n40018
g37583 and pi0214 n40018_not ; n40019
g37584 and n40017_not n40019 ; n40020
g37585 and n40016 n40020_not ; n40021
g37586 and pi0209 n40015 ; n40022
g37587 and n40021_not n40022 ; n40023
g37588 and n40013_not n40023 ; n40024
g37589 and pi0213 n39999_not ; n40025
g37590 and n40024_not n40025 ; n40026
g37591 and n39997_not n40026 ; n40027
g37592 and po1038 n39145_not ; n40028
g37593 and n38421 n39149_not ; n40029
g37594 and n40028 n40029 ; n40030
g37595 and pi0211 n38510_not ; n40031
g37596 and n39463_not n40031 ; n40032
g37597 and n40019 n40032_not ; n40033
g37598 and n40003 n40033_not ; n40034
g37599 nor pi0211 n38514 ; n40035
g37600 and n39463_not n40035 ; n40036
g37601 and pi0214 n40017_not ; n40037
g37602 and n40036_not n40037 ; n40038
g37603 and n40016 n40038_not ; n40039
g37604 and n40015 n40034_not ; n40040
g37605 and n40039_not n40040 ; n40041
g37606 and pi0209 n40041_not ; n40042
g37607 nor n38514 n38839 ; n40043
g37608 and n39991 n40043_not ; n40044
g37609 and n39989 n40044_not ; n40045
g37610 and n38861_not n40031 ; n40046
g37611 and pi0214 n40046_not ; n40047
g37612 and n39992_not n40047 ; n40048
g37613 and n39974 n40048_not ; n40049
g37614 and n39971 n40049_not ; n40050
g37615 and n40045_not n40050 ; n40051
g37616 nor pi0209 n40051 ; n40052
g37617 nor n40042 n40052 ; n40053
g37618 nor pi0213 n40030 ; n40054
g37619 and n40053_not n40054 ; n40055
g37620 nor n40027 n40055 ; n40056
g37621 and pi0230 n40056_not ; n40057
g37622 nor pi0230 pi0239 ; n40058
g37623 nor n40057 n40058 ; po0396
g37624 and po1038_not n39736 ; n40060
g37625 nor n39830 n40060 ; n40061
g37626 nor pi0214 n39736 ; n40062
g37627 nor pi0212 n40062 ; n40063
g37628 and n11384 n38449 ; n40064
g37629 nor pi0299 n40064 ; n40065
g37630 and n39713_not n40065 ; n40066
g37631 and pi0214 n40066 ; n40067
g37632 and n40063 n40067_not ; n40068
g37633 nor pi0219 n40068 ; n40069
g37634 and pi0211 n39736 ; n40070
g37635 nor pi0211 n40066 ; n40071
g37636 and pi0214 n40070_not ; n40072
g37637 and n40071_not n40072 ; n40073
g37638 and pi0212 n40073_not ; n40074
g37639 and n40066_not n40074 ; n40075
g37640 and n40069 n40075_not ; n40076
g37641 nor n40061 n40076 ; n40077
g37642 nor n39865 n40077 ; n40078
g37643 and pi1147_not n40078 ; n40079
g37644 and pi0211_not po1038 ; n40080
g37645 nor n39374 n40080 ; n40081
g37646 nor n38413 n40081 ; n40082
g37647 and pi0299 n38413_not ; n40083
g37648 nor po1038 n38415 ; n40084
g37649 and n40083 n40084 ; n40085
g37650 and n38550 n38825_not ; n40086
g37651 and po1038_not n40086 ; n40087
g37652 nor n40085 n40087 ; n40088
g37653 and n40082_not n40088 ; n40089
g37654 and pi1147 n40089 ; n40090
g37655 and pi1149 n40090_not ; n40091
g37656 and n40079_not n40091 ; n40092
g37657 and pi0211 n38421 ; n40093
g37658 and pi0212 n38783 ; n40094
g37659 nor n40093 n40094 ; n40095
g37660 and n39374 n40095_not ; n40096
g37661 nor n38826 n39039 ; n40097
g37662 and n10487_not n38533 ; n40098
g37663 nor n40097 n40098 ; n40099
g37664 and n39715 n40099 ; n40100
g37665 and pi0299 n10484 ; n40101
g37666 nor n40100 n40101 ; n40102
g37667 nor pi0212 n40102 ; n40103
g37668 nor pi0219 n40103 ; n40104
g37669 nor pi0299 n40099 ; n40105
g37670 and pi0214 n40105_not ; n40106
g37671 and pi0214_not n40100 ; n40107
g37672 nor pi0212 n40107 ; n40108
g37673 and n40106_not n40108 ; n40109
g37674 nor pi0211 n40105 ; n40110
g37675 nor n40100 n40110 ; n40111
g37676 and pi0214 n40111_not ; n40112
g37677 and pi0212 n40112_not ; n40113
g37678 nor pi0214 n40105 ; n40114
g37679 and n40113 n40114_not ; n40115
g37680 nor n40109 n40115 ; n40116
g37681 nor n13061 n40100 ; n40117
g37682 and n40106_not n40117 ; n40118
g37683 and pi0212 n40118_not ; n40119
g37684 and n40116 n40119 ; n40120
g37685 and n40104 n40120_not ; n40121
g37686 and pi0219 n40100_not ; n40122
g37687 nor po1038 n40122 ; n40123
g37688 and n40121_not n40123 ; n40124
g37689 nor n40096 n40124 ; n40125
g37690 and pi1147_not n40125 ; n40126
g37691 nor po1038 n39747 ; n40127
g37692 and pi0212 n38744_not ; n40128
g37693 nor pi0219 n40093 ; n40129
g37694 and n40128_not n40129 ; n40130
g37695 and n38416 n40130_not ; n40131
g37696 and n40085 n40130_not ; n40132
g37697 nor n40127 n40131 ; n40133
g37698 and n40132_not n40133 ; n40134
g37699 and pi1147 n40134 ; n40135
g37700 nor pi1149 n40135 ; n40136
g37701 and n40126_not n40136 ; n40137
g37702 nor n40092 n40137 ; n40138
g37703 and pi1148 n40138_not ; n40139
g37704 and n16479 n39636 ; n40140
g37705 nor pi0219 n16479 ; n40141
g37706 and n39825 n40141 ; n40142
g37707 nor n40140 n40142 ; n40143
g37708 and pi1147_not n40143 ; n40144
g37709 and n10486 n39825_not ; n40145
g37710 and n38416 n40145_not ; n40146
g37711 nor pi0211 n39661 ; n40147
g37712 and pi0211 n39686_not ; n40148
g37713 and pi0214 n40148_not ; n40149
g37714 and n40147_not n40149 ; n40150
g37715 and n10843 n40150_not ; n40151
g37716 and pi0214_not n39661 ; n40152
g37717 nor pi0212 n40152 ; n40153
g37718 and pi0214 n39697 ; n40154
g37719 and n40153 n40154_not ; n40155
g37720 nor pi0219 n40155 ; n40156
g37721 and pi0212 n40150_not ; n40157
g37722 and n39697_not n40157 ; n40158
g37723 and n40156 n40158_not ; n40159
g37724 and n40151_not n40159 ; n40160
g37725 and pi0212 n39697_not ; n40161
g37726 and pi0219 n40161_not ; n40162
g37727 and n40155_not n40162 ; n40163
g37728 nor po1038 n40163 ; n40164
g37729 and n40160_not n40164 ; n40165
g37730 nor n40146 n40165 ; n40166
g37731 and pi1147 n40166 ; n40167
g37732 and pi1149 n40144_not ; n40168
g37733 and n40167_not n40168 ; n40169
g37734 nor pi0212 n40101 ; n40170
g37735 and n39747 n40170 ; n40171
g37736 and n39747 n39854_not ; n40172
g37737 nor n39748 n40172 ; n40173
g37738 and pi0214_not n13061 ; n40174
g37739 and pi0212 n40174_not ; n40175
g37740 and n40173_not n40175 ; n40176
g37741 nor n40171 n40176 ; n40177
g37742 nor pi0219 n40177 ; n40178
g37743 and n38700 n39710_not ; n40179
g37744 and pi0208 n40179_not ; n40180
g37745 nor pi0199 n40180 ; n40181
g37746 nor n39747 n40181 ; n40182
g37747 nor pi0299 n40182 ; n40183
g37748 and pi0219_not n40183 ; n40184
g37749 nor n40178 n40184 ; n40185
g37750 nor pi0211 n40185 ; n40186
g37751 and n13061_not n39882 ; n40187
g37752 and pi0214_not n40172 ; n40188
g37753 and pi0212 n40188_not ; n40189
g37754 and n40187_not n40189 ; n40190
g37755 and pi0212_not n40173 ; n40191
g37756 nor pi0219 n40191 ; n40192
g37757 and n40190_not n40192 ; n40193
g37758 and pi0219 n39854_not ; n40194
g37759 and n40084 n40194_not ; n40195
g37760 nor n40127 n40195 ; n40196
g37761 nor n40193 n40196 ; n40197
g37762 and n40183_not n40197 ; n40198
g37763 and n40186_not n40198 ; n40199
g37764 nor n39869 n40199 ; n40200
g37765 and pi1147 pi1149_not ; n40201
g37766 and n40200_not n40201 ; n40202
g37767 nor n40169 n40202 ; n40203
g37768 nor pi1148 n40203 ; n40204
g37769 nor n40139 n40204 ; n40205
g37770 and pi0213 n40205_not ; n40206
g37771 and n10846 n38665 ; n40207
g37772 and po1038 n40207 ; n40208
g37773 and pi0211_not pi1146 ; n40209
g37774 and pi0211 pi1145 ; n40210
g37775 nor n40209 n40210 ; n40211
g37776 and pi0214 n40211_not ; n40212
g37777 and pi0211 pi1146 ; n40213
g37778 and pi0214_not n40213 ; n40214
g37779 nor n40212 n40214 ; n40215
g37780 and pi0212 n40215_not ; n40216
g37781 and n38421 n40213 ; n40217
g37782 nor n40216 n40217 ; n40218
g37783 and n38970_not n40218 ; n40219
g37784 and po1038 n39412 ; n40220
g37785 nor n39374 n40220 ; n40221
g37786 nor n40219 n40221 ; n40222
g37787 and pi1147 n40208_not ; n40223
g37788 and n40222_not n40223 ; n40224
g37789 and pi0211_not n39484 ; n40225
g37790 and pi0219 n40225_not ; n40226
g37791 and n40084 n40226_not ; n40227
g37792 nor n40127 n40227 ; n40228
g37793 and n38413 n39747_not ; n40229
g37794 nor pi0219 n40229 ; n40230
g37795 and pi0299 n40211_not ; n40231
g37796 and n39747 n40231_not ; n40232
g37797 and n10843 n40232_not ; n40233
g37798 and pi0299 pi1146 ; n40234
g37799 and pi0211 n40234 ; n40235
g37800 nor n39854 n40235 ; n40236
g37801 and n39747 n40236 ; n40237
g37802 and n38608 n40237_not ; n40238
g37803 and n40230 n40233_not ; n40239
g37804 and n40238_not n40239 ; n40240
g37805 nor n40228 n40240 ; n40241
g37806 and n40224 n40241_not ; n40242
g37807 and po1038_not n40100 ; n40243
g37808 nor pi1147 n40222 ; n40244
g37809 and pi0219 n40227 ; n40245
g37810 and pi0299 n40218_not ; n40246
g37811 and n36114 n40246 ; n40247
g37812 nor n40245 n40247 ; n40248
g37813 and n40244 n40248 ; n40249
g37814 and n40243_not n40249 ; n40250
g37815 and pi1148 n40242_not ; n40251
g37816 and n40250_not n40251 ; n40252
g37817 and n39412 n39422 ; n40253
g37818 and n38665_not n40182 ; n40254
g37819 and pi1146_not n13061 ; n40255
g37820 and n38608 n40255_not ; n40256
g37821 nor n40233 n40256 ; n40257
g37822 nor pi0219 n40183 ; n40258
g37823 and n40257_not n40258 ; n40259
g37824 nor n40253 n40254 ; n40260
g37825 and n40259_not n40260 ; n40261
g37826 nor po1038 n40261 ; n40262
g37827 and n40224 n40262_not ; n40263
g37828 nor pi1148 n40249 ; n40264
g37829 and n40263_not n40264 ; n40265
g37830 nor n40252 n40265 ; n40266
g37831 nor pi1149 n40266 ; n40267
g37832 and pi0219 n39661 ; n40268
g37833 nor po1038 n40268 ; n40269
g37834 nor n40227 n40269 ; n40270
g37835 and pi0299_not n39685 ; n40271
g37836 nor n39431 n40271 ; n40272
g37837 and n40234_not n40272 ; n40273
g37838 and pi0211 n40273_not ; n40274
g37839 nor n39695 n40274 ; n40275
g37840 and pi0214 n40275 ; n40276
g37841 and n40153 n40276_not ; n40277
g37842 and pi0214 n40231_not ; n40278
g37843 and n40272 n40278 ; n40279
g37844 and pi0214_not n40275 ; n40280
g37845 and pi0212 n40279_not ; n40281
g37846 and n40280_not n40281 ; n40282
g37847 nor pi0219 n40277 ; n40283
g37848 and n40282_not n40283 ; n40284
g37849 nor n40270 n40284 ; n40285
g37850 and n40224 n40285_not ; n40286
g37851 and n40140_not n40249 ; n40287
g37852 nor pi1148 n40287 ; n40288
g37853 and n40286_not n40288 ; n40289
g37854 and pi0219 n40086_not ; n40290
g37855 nor po1038 n40290 ; n40291
g37856 and pi0211 n40086_not ; n40292
g37857 and pi0214 pi0299 ; n40293
g37858 nor n40086 n40293 ; n40294
g37859 nor pi0212 n40294 ; n40295
g37860 and n40292_not n40295 ; n40296
g37861 nor pi0299 n40086 ; n40297
g37862 and pi0212 n40297_not ; n40298
g37863 and pi0299 n40128 ; n40299
g37864 and n40298 n40299_not ; n40300
g37865 nor pi0219 n40296 ; n40301
g37866 and n40300_not n40301 ; n40302
g37867 and n40291 n40302_not ; n40303
g37868 and n40224 n40248 ; n40304
g37869 and n40303_not n40304 ; n40305
g37870 and n38414_not n39736 ; n40306
g37871 and n38413_not n40071 ; n40307
g37872 and pi0219 n40306_not ; n40308
g37873 and n40307_not n40308 ; n40309
g37874 nor po1038 n40309 ; n40310
g37875 and n11384 n40310 ; n40311
g37876 nor n40227 n40311 ; n40312
g37877 nor n39736 n40235 ; n40313
g37878 and n40063 n40313_not ; n40314
g37879 and pi0212 n40066_not ; n40315
g37880 and n39736_not n40215 ; n40316
g37881 and n40315 n40316_not ; n40317
g37882 nor pi0219 n40314 ; n40318
g37883 and n40317_not n40318 ; n40319
g37884 nor n40312 n40319 ; n40320
g37885 and n40244 n40320_not ; n40321
g37886 and pi1148 n40305_not ; n40322
g37887 and n40321_not n40322 ; n40323
g37888 nor n40289 n40323 ; n40324
g37889 and pi1149 n40324_not ; n40325
g37890 nor n40267 n40325 ; n40326
g37891 nor pi0213 n40326 ; n40327
g37892 and pi0209 n40327_not ; n40328
g37893 and n40206_not n40328 ; n40329
g37894 and pi0200 n39393_not ; n40330
g37895 and pi0199 pi1145 ; n40331
g37896 nor pi0200 n40331 ; n40332
g37897 and pi0199_not pi1146 ; n40333
g37898 and n40332 n40333_not ; n40334
g37899 and n38441 n40330_not ; n40335
g37900 and n40334_not n40335 ; n40336
g37901 nor n38826 n40336 ; n40337
g37902 and pi0200 n40333_not ; n40338
g37903 nor pi0299 n40338 ; n40339
g37904 and n40332_not n40339 ; n40340
g37905 nor n10487 n40340 ; n40341
g37906 nor n40337 n40341 ; n40342
g37907 and n38413 n40342 ; n40343
g37908 and pi0219 n40343_not ; n40344
g37909 and n38413_not n40342 ; n40345
g37910 nor n38414 n40345 ; n40346
g37911 and n38699 n40331_not ; n40347
g37912 and n40339 n40347_not ; n40348
g37913 and pi0207_not n40348 ; n40349
g37914 and n40332 n40349 ; n40350
g37915 nor n40234 n40336 ; n40351
g37916 and n40349_not n40351 ; n40352
g37917 and pi0208 n40352_not ; n40353
g37918 and n40350_not n40353 ; n40354
g37919 and n38449 n40340 ; n40355
g37920 nor n40354 n40355 ; n40356
g37921 nor pi0299 n40356 ; n40357
g37922 nor pi0211 n39484 ; n40358
g37923 and n40357_not n40358 ; n40359
g37924 nor n40346 n40359 ; n40360
g37925 and n40344 n40360_not ; n40361
g37926 nor n40235 n40342 ; n40362
g37927 nor pi0214 n40342 ; n40363
g37928 nor pi0212 n40363 ; n40364
g37929 and n40362_not n40364 ; n40365
g37930 nor pi0219 n40365 ; n40366
g37931 and n40278 n40357_not ; n40367
g37932 and pi0214_not n40362 ; n40368
g37933 and pi0212 n40368_not ; n40369
g37934 and n40367_not n40369 ; n40370
g37935 and n40366 n40370_not ; n40371
g37936 nor po1038 n40361 ; n40372
g37937 and n40371_not n40372 ; n40373
g37938 and n40244 n40373_not ; n40374
g37939 nor n10487 n40348 ; n40375
g37940 nor n40337 n40375 ; n40376
g37941 and n38414_not n40376 ; n40377
g37942 and pi0219 n40377_not ; n40378
g37943 and n38449 n40348 ; n40379
g37944 nor n40353 n40379 ; n40380
g37945 and pi0299_not n40380 ; n40381
g37946 nor pi0211 n40381 ; n40382
g37947 and n39481_not n40382 ; n40383
g37948 and n38413_not n40383 ; n40384
g37949 and n40378 n40384_not ; n40385
g37950 nor n40376 n40382 ; n40386
g37951 nor pi0214 n40376 ; n40387
g37952 nor pi0212 n40387 ; n40388
g37953 and n40386_not n40388 ; n40389
g37954 and pi0211 n40381_not ; n40390
g37955 and n39481_not n40390 ; n40391
g37956 and n40278 n40380 ; n40392
g37957 and n10484 n40381_not ; n40393
g37958 nor n40392 n40393 ; n40394
g37959 nor n40391 n40394 ; n40395
g37960 and pi0214_not n40236 ; n40396
g37961 and n40380 n40396 ; n40397
g37962 and pi0212 n40397_not ; n40398
g37963 and n40395_not n40398 ; n40399
g37964 and n40366 n40389_not ; n40400
g37965 and n40399_not n40400 ; n40401
g37966 nor po1038 n40385 ; n40402
g37967 and n40401_not n40402 ; n40403
g37968 and n40224 n40403_not ; n40404
g37969 nor n40374 n40404 ; n40405
g37970 and pi0213_not n40405 ; n40406
g37971 and pi1147 n40131_not ; n40407
g37972 and n38413_not n40382 ; n40408
g37973 and n40378 n40408_not ; n40409
g37974 nor po1038 n40409 ; n40410
g37975 and pi0299_not n40356 ; n40411
g37976 and pi0214 n40411_not ; n40412
g37977 nor n40390 n40412 ; n40413
g37978 and pi0212 n40413_not ; n40414
g37979 nor pi0219 n40376 ; n40415
g37980 and n40393_not n40415 ; n40416
g37981 and n40414_not n40416 ; n40417
g37982 and n40410 n40417_not ; n40418
g37983 and n40407 n40418_not ; n40419
g37984 and n40343_not n40417 ; n40420
g37985 and pi0219 n40342_not ; n40421
g37986 and pi0214 n40386 ; n40422
g37987 nor n40411 n40422 ; n40423
g37988 and pi0212 n40423_not ; n40424
g37989 and pi0214_not n40342 ; n40425
g37990 nor pi0212 n40425 ; n40426
g37991 and n40412_not n40426 ; n40427
g37992 nor n40424 n40427 ; n40428
g37993 nor pi0219 n40428 ; n40429
g37994 nor po1038 n40421 ; n40430
g37995 and n40429_not n40430 ; n40431
g37996 and n40420_not n40431 ; n40432
g37997 nor pi1147 n40096 ; n40433
g37998 and n40432_not n40433 ; n40434
g37999 nor pi1149 n40419 ; n40435
g38000 and n40434_not n40435 ; n40436
g38001 and n40083_not n40415 ; n40437
g38002 and n40410 n40437_not ; n40438
g38003 and pi1147 n40082_not ; n40439
g38004 and n40438_not n40439 ; n40440
g38005 nor pi1147 n39865 ; n40441
g38006 and n40431_not n40441 ; n40442
g38007 and pi1149 n40440_not ; n40443
g38008 and n40442_not n40443 ; n40444
g38009 and pi1148 n40444_not ; n40445
g38010 and n40436_not n40445 ; n40446
g38011 nor pi1147 po1038 ; n40447
g38012 and n40342 n40447 ; n40448
g38013 and pi0214 n40376_not ; n40449
g38014 and n40390_not n40449 ; n40450
g38015 and n40382_not n40387 ; n40451
g38016 and pi0212 n40450_not ; n40452
g38017 and n40451_not n40452 ; n40453
g38018 nor pi0219 n40389 ; n40454
g38019 and n40453_not n40454 ; n40455
g38020 and n40418 n40455_not ; n40456
g38021 nor n39869 n40456 ; n40457
g38022 and pi1147 n40457_not ; n40458
g38023 nor n40448 n40458 ; n40459
g38024 nor pi1149 n40459 ; n40460
g38025 and n40410 n40455_not ; n40461
g38026 nor n40146 n40461 ; n40462
g38027 and pi1147 n40462_not ; n40463
g38028 and pi1147_not n40207 ; n40464
g38029 nor n40448 n40464 ; n40465
g38030 and n16479 n40207 ; n40466
g38031 and n40356 n40466 ; n40467
g38032 nor n40465 n40467 ; n40468
g38033 nor n40463 n40468 ; n40469
g38034 and pi1149 n40469_not ; n40470
g38035 nor pi1148 n40470 ; n40471
g38036 and n40460_not n40471 ; n40472
g38037 and pi0213 n40446_not ; n40473
g38038 and n40472_not n40473 ; n40474
g38039 nor pi0209 n40406 ; n40475
g38040 and n40474_not n40475 ; n40476
g38041 nor n40329 n40476 ; n40477
g38042 and pi0230 n40477_not ; n40478
g38043 nor pi0230 pi0240 ; n40479
g38044 nor n40478 n40479 ; po0397
g38045 and pi0213 n39907_not ; n40481
g38046 and n39635 n39646 ; n40482
g38047 and n38508 n39825 ; n40483
g38048 nor n39662 n40483 ; n40484
g38049 and po1038 n40207_not ; n40485
g38050 and pi1151 n40485_not ; n40486
g38051 and n40484_not n40486 ; n40487
g38052 nor n40482 n40487 ; n40488
g38053 nor pi1152 n40488 ; n40489
g38054 and n39755_not n40207 ; n40490
g38055 and n39872 n40490_not ; n40491
g38056 and pi1152 n40491_not ; n40492
g38057 nor po1038 n40492 ; n40493
g38058 and n40486 n40493_not ; n40494
g38059 and pi1152 n39635 ; n40495
g38060 and n39737 n40495 ; n40496
g38061 nor n40489 n40496 ; n40497
g38062 and n40494_not n40497 ; n40498
g38063 nor pi1150 n40498 ; n40499
g38064 and pi1151 n39865_not ; n40500
g38065 and pi0219 n39646_not ; n40501
g38066 nor po1038 n40501 ; n40502
g38067 nor n40127 n40502 ; n40503
g38068 and n39750 n39885_not ; n40504
g38069 nor pi0219 n40504 ; n40505
g38070 and pi0214_not n39755 ; n40506
g38071 and pi0212 n40506_not ; n40507
g38072 and n39874_not n40507 ; n40508
g38073 and n40505 n40508_not ; n40509
g38074 and pi1152 n40509_not ; n40510
g38075 nor pi0299 n39687 ; n40511
g38076 and pi0214_not n39686 ; n40512
g38077 and pi0212 n40512_not ; n40513
g38078 and n40154_not n40513 ; n40514
g38079 nor n39664 n40514 ; n40515
g38080 nor n40511 n40515 ; n40516
g38081 nor pi0219 n40516 ; n40517
g38082 nor pi1152 n40268 ; n40518
g38083 and n40517_not n40518 ; n40519
g38084 nor n40510 n40519 ; n40520
g38085 nor n40503 n40520 ; n40521
g38086 and n40500 n40521_not ; n40522
g38087 nor pi1151 n40096 ; n40523
g38088 nor pi0212 n39637 ; n40524
g38089 and n39640_not n40524 ; n40525
g38090 and n39854_not n40525 ; n40526
g38091 nor pi0219 n40526 ; n40527
g38092 and pi0214 n39638_not ; n40528
g38093 and pi0211_not n39640 ; n40529
g38094 and pi0212 n39637_not ; n40530
g38095 and n40529_not n40530 ; n40531
g38096 and n40528_not n40531 ; n40532
g38097 and n40527 n40532_not ; n40533
g38098 and n39646_not n39834 ; n40534
g38099 and pi0299_not n40534 ; n40535
g38100 nor n40533 n40535 ; n40536
g38101 and n40502 n40536 ; n40537
g38102 nor pi1152 n40537 ; n40538
g38103 nor n39737 n40536 ; n40539
g38104 and n39895 n40539_not ; n40540
g38105 and pi1152 n40540_not ; n40541
g38106 nor n40538 n40541 ; n40542
g38107 and n40523 n40542_not ; n40543
g38108 and pi1150 n40543_not ; n40544
g38109 and n40522_not n40544 ; n40545
g38110 nor n40499 n40545 ; n40546
g38111 nor pi1149 n40546 ; n40547
g38112 and pi1151 n40146_not ; n40548
g38113 nor pi0214 n39856 ; n40549
g38114 and n39849 n40549_not ; n40550
g38115 nor pi0212 n39857 ; n40551
g38116 nor n40550 n40551 ; n40552
g38117 nor pi0219 n40552 ; n40553
g38118 and pi1152_not n39859 ; n40554
g38119 and n40553_not n40554 ; n40555
g38120 nor n38783 n39755 ; n40556
g38121 and pi0212 n39872 ; n40557
g38122 and n40556_not n40557 ; n40558
g38123 nor n39876 n40558 ; n40559
g38124 nor pi0219 n40559 ; n40560
g38125 and pi1152 n40560_not ; n40561
g38126 and n39879 n40561 ; n40562
g38127 and n40548 n40555_not ; n40563
g38128 and n40562_not n40563 ; n40564
g38129 nor pi1151 n39869 ; n40565
g38130 nor n40195 n40502 ; n40566
g38131 nor n40534 n40566 ; n40567
g38132 and pi1152_not n40567 ; n40568
g38133 and n39895_not n40566 ; n40569
g38134 and n39737_not n39834 ; n40570
g38135 and pi1152 n40569_not ; n40571
g38136 and n40570_not n40571 ; n40572
g38137 and n40565 n40568_not ; n40573
g38138 and n40572_not n40573 ; n40574
g38139 nor pi1150 n40574 ; n40575
g38140 and n40564_not n40575 ; n40576
g38141 nor pi1151 n40131 ; n40577
g38142 and n10843 n39724 ; n40578
g38143 nor n39641 n39831 ; n40579
g38144 nor n10843 n39737 ; n40580
g38145 and n40579_not n40580 ; n40581
g38146 nor n40578 n40581 ; n40582
g38147 nor pi0219 n40582 ; n40583
g38148 nor n40569 n40583 ; n40584
g38149 and pi1152 n40584_not ; n40585
g38150 and n40538 n40567_not ; n40586
g38151 nor n40585 n40586 ; n40587
g38152 and n40577 n40587_not ; n40588
g38153 and pi0212 n39755_not ; n40589
g38154 and n40505 n40589_not ; n40590
g38155 and pi1152 n40590_not ; n40591
g38156 and n39879 n40591 ; n40592
g38157 and pi1151 n40082_not ; n40593
g38158 nor n39699 n40511 ; n40594
g38159 nor pi0219 n40594 ; n40595
g38160 and n40554 n40595_not ; n40596
g38161 and n40593 n40596_not ; n40597
g38162 and n40592_not n40597 ; n40598
g38163 and pi1150 n40588_not ; n40599
g38164 and n40598_not n40599 ; n40600
g38165 nor n40576 n40600 ; n40601
g38166 and pi1149 n40601_not ; n40602
g38167 nor n40547 n40602 ; n40603
g38168 nor pi0213 n40603 ; n40604
g38169 and pi0209 n40481_not ; n40605
g38170 and n40604_not n40605 ; n40606
g38171 and pi1150_not pi1151 ; n40607
g38172 and n40143_not n40607 ; n40608
g38173 and n40124_not n40523 ; n40609
g38174 and n40077_not n40500 ; n40610
g38175 and pi1150 n40610_not ; n40611
g38176 and n40609_not n40611 ; n40612
g38177 nor pi1149 n40608 ; n40613
g38178 and n40612_not n40613 ; n40614
g38179 and n40088 n40593 ; n40615
g38180 and pi1151_not n40134 ; n40616
g38181 and pi1150 n40615_not ; n40617
g38182 and n40616_not n40617 ; n40618
g38183 and n40199_not n40565 ; n40619
g38184 and n40165_not n40548 ; n40620
g38185 nor pi1150 n40619 ; n40621
g38186 and n40620_not n40621 ; n40622
g38187 and pi1149 n40618_not ; n40623
g38188 and n40622_not n40623 ; n40624
g38189 nor n40614 n40624 ; n40625
g38190 and pi0213_not n40625 ; n40626
g38191 nor n40153 n40157 ; n40627
g38192 and n38769_not n39695 ; n40628
g38193 nor n39696 n40628 ; n40629
g38194 and n40151_not n40629 ; n40630
g38195 nor n40627 n40630 ; n40631
g38196 nor pi0219 n40631 ; n40632
g38197 and n40164 n40632_not ; n40633
g38198 and n39845 n40633_not ; n40634
g38199 and pi0299 n39631 ; n40635
g38200 nor n40182 n40483 ; n40636
g38201 nor po1038 n40636 ; n40637
g38202 and n40635_not n40637 ; n40638
g38203 and n39828 n40638_not ; n40639
g38204 nor pi1152 n40639 ; n40640
g38205 and n40634_not n40640 ; n40641
g38206 nor n40150 n40152 ; n40642
g38207 nor pi0219 n40299 ; n40643
g38208 and n39700_not n40643 ; n40644
g38209 and n40642_not n40644 ; n40645
g38210 and n40164 n40645_not ; n40646
g38211 and n39871 n40646_not ; n40647
g38212 nor n40083 n40182 ; n40648
g38213 and n38641_not n39867 ; n40649
g38214 nor n40648 n40649 ; n40650
g38215 nor pi0219 n40650 ; n40651
g38216 and pi0219 n40182_not ; n40652
g38217 nor po1038 n40652 ; n40653
g38218 and n40651_not n40653 ; n40654
g38219 and n39893 n40654_not ; n40655
g38220 and pi1152 n40655_not ; n40656
g38221 and n40647_not n40656 ; n40657
g38222 nor pi1150 n40657 ; n40658
g38223 and n40641_not n40658 ; n40659
g38224 nor pi0219 n40086 ; n40660
g38225 and n40299_not n40660 ; n40661
g38226 and pi1153_not n40661 ; n40662
g38227 and pi0299 n10485 ; n40663
g38228 nor pi0219 n40663 ; n40664
g38229 and n40195 n40664_not ; n40665
g38230 nor n40303 n40665 ; n40666
g38231 nor n40662 n40666 ; n40667
g38232 and n39845 n40667_not ; n40668
g38233 and pi1153 n40483 ; n40669
g38234 and n39828 n40669_not ; n40670
g38235 nor pi1152 n40670 ; n40671
g38236 nor pi1151 n40127 ; n40672
g38237 nor pi1152 n40672 ; n40673
g38238 nor n40671 n40673 ; n40674
g38239 nor n40668 n40674 ; n40675
g38240 and pi0211_not n40661 ; n40676
g38241 nor n40088 n40676 ; n40677
g38242 and n39871 n40677_not ; n40678
g38243 and n40667_not n40678 ; n40679
g38244 nor po1038 n39768 ; n40680
g38245 and n10843 n40172_not ; n40681
g38246 and pi0299_not n39747 ; n40682
g38247 nor n38423 n40635 ; n40683
g38248 and n40682_not n40683 ; n40684
g38249 and n40230 n40681_not ; n40685
g38250 and n40684_not n40685 ; n40686
g38251 and n40680 n40686_not ; n40687
g38252 and n39893 n40687_not ; n40688
g38253 and pi1152 n40688_not ; n40689
g38254 and n40679_not n40689 ; n40690
g38255 and pi1150 n40675_not ; n40691
g38256 and n40690_not n40691 ; n40692
g38257 and pi1149 n40692_not ; n40693
g38258 and n40659_not n40693 ; n40694
g38259 and pi0219 n39642_not ; n40695
g38260 nor po1038 n40695 ; n40696
g38261 and n39839_not n40696 ; n40697
g38262 and n39845 n40697_not ; n40698
g38263 and n40671 n40698_not ; n40699
g38264 and pi0299 n39864 ; n40700
g38265 and n39867_not n40700 ; n40701
g38266 and n39893 n40701_not ; n40702
g38267 and n40527 n40531_not ; n40703
g38268 and n40696 n40703_not ; n40704
g38269 and n39871 n40697_not ; n40705
g38270 and n40704_not n40705 ; n40706
g38271 and pi1152 n40702_not ; n40707
g38272 and n40706_not n40707 ; n40708
g38273 nor pi1150 n40699 ; n40709
g38274 and n40708_not n40709 ; n40710
g38275 and n39909_not n40100 ; n40711
g38276 nor n38769 n40105 ; n40712
g38277 nor pi0211 n40712 ; n40713
g38278 and n39909 n40111_not ; n40714
g38279 and n40713_not n40714 ; n40715
g38280 nor n40711 n40715 ; n40716
g38281 nor po1038 n40716 ; n40717
g38282 and n39828 n40717_not ; n40718
g38283 and pi0211 n40066_not ; n40719
g38284 and n11373_not n38675 ; n40720
g38285 nor n39713 n40720 ; n40721
g38286 nor pi0211 n38769 ; n40722
g38287 and n40721_not n40722 ; n40723
g38288 nor n40719 n40723 ; n40724
g38289 nor n39736 n40719 ; n40725
g38290 and pi0214 n40725 ; n40726
g38291 and n40062 n40071_not ; n40727
g38292 and pi0212 n40727_not ; n40728
g38293 and n40726_not n40728 ; n40729
g38294 and n40724_not n40729 ; n40730
g38295 nor n40070 n40723 ; n40731
g38296 and n40063 n40731_not ; n40732
g38297 nor pi0219 n40732 ; n40733
g38298 and n40730_not n40733 ; n40734
g38299 and n40310 n40734_not ; n40735
g38300 and n39845 n40735_not ; n40736
g38301 nor pi1152 n40718 ; n40737
g38302 and n40736_not n40737 ; n40738
g38303 and pi0214 n40724 ; n40739
g38304 and n40063 n40739_not ; n40740
g38305 and pi0214_not n40724 ; n40741
g38306 and n40315 n40741_not ; n40742
g38307 nor pi0219 n40740 ; n40743
g38308 and n40742_not n40743 ; n40744
g38309 and n40310 n40744_not ; n40745
g38310 and n39871 n40745_not ; n40746
g38311 nor n40105 n40635 ; n40747
g38312 and pi0214 n40747 ; n40748
g38313 and n40108 n40748_not ; n40749
g38314 and pi0214_not n40747 ; n40750
g38315 and n40113 n40750_not ; n40751
g38316 nor n40749 n40751 ; n40752
g38317 nor pi0219 n40752 ; n40753
g38318 and n40123 n40753_not ; n40754
g38319 and n39893 n40754_not ; n40755
g38320 and pi1152 n40746_not ; n40756
g38321 and n40755_not n40756 ; n40757
g38322 and pi1150 n40738_not ; n40758
g38323 and n40757_not n40758 ; n40759
g38324 nor pi1149 n40710 ; n40760
g38325 and n40759_not n40760 ; n40761
g38326 nor n40694 n40761 ; n40762
g38327 and pi0213 n40762_not ; n40763
g38328 nor pi0209 n40626 ; n40764
g38329 and n40763_not n40764 ; n40765
g38330 nor n40606 n40765 ; n40766
g38331 and pi0230 n40766_not ; n40767
g38332 nor pi0230 pi0241 ; n40768
g38333 nor n40767 n40768 ; po0398
g38334 nor pi0230 pi0242 ; n40770
g38335 and pi0219 n38419_not ; n40771
g38336 and pi0214 n39414_not ; n40772
g38337 nor pi0214 n40211 ; n40773
g38338 nor n40772 n40773 ; n40774
g38339 and pi0212 n40774_not ; n40775
g38340 and pi0212_not n40212 ; n40776
g38341 nor pi0219 n40776 ; n40777
g38342 and n40775_not n40777 ; n40778
g38343 and n38416 n40771_not ; n40779
g38344 and n40778_not n40779 ; n40780
g38345 and pi0199 pi1144 ; n40781
g38346 nor pi0200 n40781 ; n40782
g38347 and n40333_not n40782 ; n40783
g38348 nor pi0299 n40330 ; n40784
g38349 and n40783_not n40784 ; n40785
g38350 and n38826 n40785 ; n40786
g38351 nor pi0207 n40785 ; n40787
g38352 nor pi0299 n39392 ; n40788
g38353 and n39393_not n40782 ; n40789
g38354 and n40788 n40789_not ; n40790
g38355 and pi0207 n40790_not ; n40791
g38356 and pi0208 n40787_not ; n40792
g38357 and n40791_not n40792 ; n40793
g38358 nor n40786 n40793 ; n40794
g38359 and pi0214_not n40794 ; n40795
g38360 nor pi0212 n40795 ; n40796
g38361 and n38449 n40785 ; n40797
g38362 nor n40234 n40797 ; n40798
g38363 and n40793_not n40798 ; n40799
g38364 nor pi0211 n40799 ; n40800
g38365 nor n39484 n40797 ; n40801
g38366 and n40793_not n40801 ; n40802
g38367 and pi0211 n40802_not ; n40803
g38368 nor n40800 n40803 ; n40804
g38369 and pi0214 n40804 ; n40805
g38370 and n40796 n40805_not ; n40806
g38371 nor pi0211 n40802 ; n40807
g38372 nor n38612 n40797 ; n40808
g38373 and n40793_not n40808 ; n40809
g38374 and pi0211 n40809_not ; n40810
g38375 and pi0214 n40807_not ; n40811
g38376 and n40810_not n40811 ; n40812
g38377 and pi0214_not n40804 ; n40813
g38378 and pi0212 n40812_not ; n40814
g38379 and n40813_not n40814 ; n40815
g38380 nor pi0219 n40806 ; n40816
g38381 and n40815_not n40816 ; n40817
g38382 nor n38414 n40794 ; n40818
g38383 and pi0219 n40818_not ; n40819
g38384 and n38414 n40809_not ; n40820
g38385 and n40819 n40820_not ; n40821
g38386 nor po1038 n40821 ; n40822
g38387 and n40817_not n40822 ; n40823
g38388 nor n40780 n40823 ; n40824
g38389 and pi0213 n40824 ; n40825
g38390 and n38413 n40786_not ; n40826
g38391 and pi0211 n40786_not ; n40827
g38392 and n38414 n38680_not ; n40828
g38393 and n40797_not n40828 ; n40829
g38394 nor n40827 n40829 ; n40830
g38395 and pi0219 n40830_not ; n40831
g38396 and n10843 n38457_not ; n40832
g38397 and n38431_not n38608 ; n40833
g38398 nor n40832 n40833 ; n40834
g38399 nor pi0219 n40797 ; n40835
g38400 and n40834_not n40835 ; n40836
g38401 nor n40826 n40836 ; n40837
g38402 and n40831_not n40837 ; n40838
g38403 nor n40793 n40838 ; n40839
g38404 nor po1038 n40839 ; n40840
g38405 nor pi0213 n38430 ; n40841
g38406 and n40840_not n40841 ; n40842
g38407 nor n40825 n40842 ; n40843
g38408 and pi0209 n40843_not ; n40844
g38409 nor pi0213 n38476 ; n40845
g38410 and pi0219 n38413 ; n40846
g38411 nor n40771 n40846 ; n40847
g38412 and n40778_not n40847 ; n40848
g38413 and pi0299 n40848_not ; n40849
g38414 nor po1038 n40849 ; n40850
g38415 and n38468_not n40850 ; n40851
g38416 nor n40780 n40851 ; n40852
g38417 and pi0213 n40852_not ; n40853
g38418 nor pi0209 n40853 ; n40854
g38419 and n40845_not n40854 ; n40855
g38420 nor n40844 n40855 ; n40856
g38421 and pi0230 n40856_not ; n40857
g38422 nor n40770 n40857 ; po0399
g38423 and pi0253 pi0254 ; n40859
g38424 and pi0267 n40859 ; n40860
g38425 and pi0263_not n40860 ; n40861
g38426 nor pi0083 pi0085 ; n40862
g38427 and pi0314 n40862_not ; n40863
g38428 and pi0802 n40863 ; n40864
g38429 and pi0276 n40864 ; n40865
g38430 and pi1091_not n40865 ; n40866
g38431 and pi0271 n40866 ; n40867
g38432 and pi0273 n40867 ; n40868
g38433 and pi0243 n40868 ; n40869
g38434 nor pi1091 n40865 ; n40870
g38435 and pi0271 n40870_not ; n40871
g38436 nor pi1091 n40871 ; n40872
g38437 and pi0273 n40872_not ; n40873
g38438 nor pi1091 n40873 ; n40874
g38439 and pi0243_not n40874 ; n40875
g38440 and pi0243 pi1091_not ; n40876
g38441 and n38478 n40876_not ; n40877
g38442 and n40866_not n40877 ; n40878
g38443 nor n40869 n40878 ; n40879
g38444 and n40875_not n40879 ; n40880
g38445 and pi0219 n40880_not ; n40881
g38446 nor n38479 n38487 ; n40882
g38447 and pi1091 n40882 ; n40883
g38448 and pi0081_not n40862 ; n40884
g38449 and pi0314 n40884_not ; n40885
g38450 and pi0802 n40885 ; n40886
g38451 and pi0276 n40886 ; n40887
g38452 and pi1091_not n40887 ; n40888
g38453 and pi0271 n40888 ; n40889
g38454 and pi0273 n40889 ; n40890
g38455 nor n40873 n40890 ; n40891
g38456 and n40876 n40891 ; n40892
g38457 and pi0243_not n40890 ; n40893
g38458 nor pi0219 n40883 ; n40894
g38459 and n40893_not n40894 ; n40895
g38460 and n40892_not n40895 ; n40896
g38461 nor n40881 n40896 ; n40897
g38462 and n40861 n40897_not ; n40898
g38463 nor pi0243 pi1091 ; n40899
g38464 nor pi0219 n40882 ; n40900
g38465 and pi1157 n38519 ; n40901
g38466 nor n40900 n40901 ; n40902
g38467 and pi1091 n40902_not ; n40903
g38468 nor n40899 n40903 ; n40904
g38469 nor n40861 n40904 ; n40905
g38470 and po1038 n40905_not ; n40906
g38471 and n40898_not n40906 ; n40907
g38472 and pi0272 pi0283 ; n40908
g38473 and pi0275 n40908 ; n40909
g38474 and pi0268 n40909 ; n40910
g38475 and pi0299_not pi1091 ; n40911
g38476 and n38841 n40911 ; n40912
g38477 nor n40899 n40912 ; n40913
g38478 and pi1156 n40913_not ; n40914
g38479 and pi1091 n38955_not ; n40915
g38480 and n39457 n40915 ; n40916
g38481 nor n40914 n40916 ; n40917
g38482 and pi0299_not n38699 ; n40918
g38483 and pi1091 n40918_not ; n40919
g38484 nor n40876 n40919 ; n40920
g38485 nor pi1155 n40899 ; n40921
g38486 nor n40876 n40921 ; n40922
g38487 and n38568 n40922 ; n40923
g38488 nor n40920 n40923 ; n40924
g38489 nor pi1156 n40924 ; n40925
g38490 and n40917 n40925_not ; n40926
g38491 and pi1157 n40926_not ; n40927
g38492 and n40915_not n40922 ; n40928
g38493 nor pi1156 n40928 ; n40929
g38494 and pi1155 n40876_not ; n40930
g38495 and pi0199 pi1091 ; n40931
g38496 and pi0299_not n40931 ; n40932
g38497 and n40930 n40932_not ; n40933
g38498 and pi1156 n40933_not ; n40934
g38499 nor pi1155 n40876 ; n40935
g38500 and n11444_not n40911 ; n40936
g38501 and n40935 n40936_not ; n40937
g38502 and n40934 n40937_not ; n40938
g38503 nor pi1157 n40929 ; n40939
g38504 and n40938_not n40939 ; n40940
g38505 nor n40927 n40940 ; n40941
g38506 and pi0211 n40941_not ; n40942
g38507 and pi1091 n11445_not ; n40943
g38508 and n40935 n40943_not ; n40944
g38509 nor n40933 n40944 ; n40945
g38510 and pi0200 pi1156_not ; n40946
g38511 and n40911 n40946 ; n40947
g38512 nor n40945 n40947 ; n40948
g38513 nor pi1157 n40948 ; n40949
g38514 and n40913 n40934 ; n40950
g38515 and pi0200 pi1091 ; n40951
g38516 and pi0299_not n40951 ; n40952
g38517 and n40930 n40952_not ; n40953
g38518 and pi1155_not n40920 ; n40954
g38519 nor pi1156 n40953 ; n40955
g38520 and n40954_not n40955 ; n40956
g38521 nor n40950 n40956 ; n40957
g38522 and pi1157 n40957_not ; n40958
g38523 nor pi0211 n40949 ; n40959
g38524 and n40958_not n40959 ; n40960
g38525 nor n40942 n40960 ; n40961
g38526 nor pi0219 n40961 ; n40962
g38527 and n39369 n40914_not ; n40963
g38528 and n40925_not n40963 ; n40964
g38529 and pi0299 pi1091 ; n40965
g38530 and n40948 n40965_not ; n40966
g38531 nor pi1157 n40966 ; n40967
g38532 and pi1091 n38700 ; n40968
g38533 and n40935 n40968_not ; n40969
g38534 nor n40953 n40969 ; n40970
g38535 nor pi1156 n40970 ; n40971
g38536 and n38478 n40971_not ; n40972
g38537 and n40917 n40972 ; n40973
g38538 and pi0219 n40964_not ; n40974
g38539 nor n40967 n40973 ; n40975
g38540 and n40974 n40975 ; n40976
g38541 nor n40962 n40976 ; n40977
g38542 nor n40861 n40977 ; n40978
g38543 and pi0199 n40874_not ; n40979
g38544 and pi1091_not n40891 ; n40980
g38545 nor pi0199 n40980 ; n40981
g38546 nor n40979 n40981 ; n40982
g38547 nor pi0200 n40888 ; n40983
g38548 nor n40982 n40983 ; n40984
g38549 nor pi0299 n40984 ; n40985
g38550 and pi0299 n40874 ; n40986
g38551 and n40890_not n40986 ; n40987
g38552 nor n40985 n40987 ; n40988
g38553 nor pi0243 n40988 ; n40989
g38554 nor pi0200 n40874 ; n40990
g38555 and n40888 n40982_not ; n40991
g38556 nor pi0299 n40991 ; n40992
g38557 and n40990_not n40992 ; n40993
g38558 and pi0299 n40868_not ; n40994
g38559 nor n40993 n40994 ; n40995
g38560 and pi0243 n40995 ; n40996
g38561 nor n40989 n40996 ; n40997
g38562 and pi1155 n40997_not ; n40998
g38563 and n40981_not n40985 ; n40999
g38564 nor n40986 n40999 ; n41000
g38565 nor pi0243 n41000 ; n41001
g38566 and n40979_not n40992 ; n41002
g38567 and n40995 n41002_not ; n41003
g38568 and pi0243 n41003 ; n41004
g38569 nor n41001 n41004 ; n41005
g38570 and n40998_not n41005 ; n41006
g38571 nor pi1156 n41006 ; n41007
g38572 and n40990_not n41002 ; n41008
g38573 nor n40986 n41008 ; n41009
g38574 and pi0243_not n41009 ; n41010
g38575 and n40979_not n40985 ; n41011
g38576 and n40981_not n40993 ; n41012
g38577 nor n40994 n41012 ; n41013
g38578 and n41011_not n41013 ; n41014
g38579 and pi0243 n41014_not ; n41015
g38580 nor n41010 n41015 ; n41016
g38581 nor pi1155 n41001 ; n41017
g38582 and pi1155 n40989_not ; n41018
g38583 and pi0243 n41013 ; n41019
g38584 and n41018 n41019_not ; n41020
g38585 nor n41017 n41020 ; n41021
g38586 nor n41016 n41021 ; n41022
g38587 and pi1156 n41022_not ; n41023
g38588 and n39369 n41007_not ; n41024
g38589 and n41023_not n41024 ; n41025
g38590 and n40981_not n40992 ; n41026
g38591 and n40996 n41026_not ; n41027
g38592 nor n40986 n41011 ; n41028
g38593 nor pi0243 n41028 ; n41029
g38594 and pi1155 n41029_not ; n41030
g38595 and n41027_not n41030 ; n41031
g38596 nor n40992 n40994 ; n41032
g38597 and n40899 n41032_not ; n41033
g38598 nor pi1155 n41033 ; n41034
g38599 and pi0243 n41032 ; n41035
g38600 and n41034 n41035_not ; n41036
g38601 nor pi1156 n41036 ; n41037
g38602 and n41031_not n41037 ; n41038
g38603 nor n40994 n41026 ; n41039
g38604 and pi1155 n41039 ; n41040
g38605 and n40985_not n41039 ; n41041
g38606 nor n41040 n41041 ; n41042
g38607 and pi0243 n41042_not ; n41043
g38608 and pi0299 n40890_not ; n41044
g38609 nor n40993 n41044 ; n41045
g38610 and pi1155_not n41045 ; n41046
g38611 and n40888_not n41046 ; n41047
g38612 nor n40986 n41002 ; n41048
g38613 nor pi0243 n41048 ; n41049
g38614 and n41047_not n41049 ; n41050
g38615 nor n41043 n41050 ; n41051
g38616 and pi1156 n41051_not ; n41052
g38617 nor pi1157 n41038 ; n41053
g38618 and n41052_not n41053 ; n41054
g38619 nor n40986 n40993 ; n41055
g38620 and pi0243 n41055_not ; n41056
g38621 nor n40994 n40999 ; n41057
g38622 nor pi0243 n41057 ; n41058
g38623 and pi0243 n41002_not ; n41059
g38624 nor pi1155 n41059 ; n41060
g38625 and n41058_not n41060 ; n41061
g38626 nor n40985 n40994 ; n41062
g38627 and pi0243_not pi1155 ; n41063
g38628 and n41062 n41063 ; n41064
g38629 nor pi1156 n41064 ; n41065
g38630 and n41056_not n41065 ; n41066
g38631 and n41061_not n41066 ; n41067
g38632 and n41014_not n41056 ; n41068
g38633 and pi1155 n41068_not ; n41069
g38634 and n41010 n41062 ; n41070
g38635 and n41069 n41070_not ; n41071
g38636 nor n41008 n41044 ; n41072
g38637 nor n40876 n41072 ; n41073
g38638 nor n41001 n41073 ; n41074
g38639 and n41016_not n41074 ; n41075
g38640 nor pi1155 n41075 ; n41076
g38641 nor n41071 n41076 ; n41077
g38642 and pi1156 n41077_not ; n41078
g38643 and n38478 n41067_not ; n41079
g38644 and n41078_not n41079 ; n41080
g38645 nor n41025 n41054 ; n41081
g38646 and n41080_not n41081 ; n41082
g38647 and pi0219 n41082_not ; n41083
g38648 nor n40992 n41044 ; n41084
g38649 and pi1155_not n41084 ; n41085
g38650 nor n41017 n41085 ; n41086
g38651 and pi0243 n41045 ; n41087
g38652 and n41002_not n41087 ; n41088
g38653 nor n41086 n41088 ; n41089
g38654 nor pi1156 n41089 ; n41090
g38655 nor n40985 n41044 ; n41091
g38656 and pi0243_not n41091 ; n41092
g38657 nor n40987 n40993 ; n41093
g38658 and pi0243 n41093_not ; n41094
g38659 nor n41092 n41094 ; n41095
g38660 and n41090 n41095 ; n41096
g38661 nor n40987 n41012 ; n41097
g38662 and pi1155 n41097 ; n41098
g38663 nor n41069 n41098 ; n41099
g38664 and n41008_not n41092 ; n41100
g38665 nor n41099 n41100 ; n41101
g38666 nor n40999 n41008 ; n41102
g38667 and n40987_not n41102 ; n41103
g38668 nor pi0243 n41103 ; n41104
g38669 nor n41011 n41044 ; n41105
g38670 and pi0243 n41012_not ; n41106
g38671 and n41105 n41106 ; n41107
g38672 nor n41104 n41107 ; n41108
g38673 nor pi1155 n41108 ; n41109
g38674 nor n41101 n41109 ; n41110
g38675 and pi1156 n41110_not ; n41111
g38676 and pi1157 n41096_not ; n41112
g38677 and n41111_not n41112 ; n41113
g38678 and pi1155_not n41093 ; n41114
g38679 and n41091_not n41114 ; n41115
g38680 nor n40987 n41026 ; n41116
g38681 and pi0243 n41116_not ; n41117
g38682 nor n41002 n41044 ; n41118
g38683 and pi0243_not n41118 ; n41119
g38684 nor n41117 n41119 ; n41120
g38685 and pi1156 n41047_not ; n41121
g38686 and n41120 n41121 ; n41122
g38687 and n41115_not n41122 ; n41123
g38688 and pi0243 n41084 ; n41124
g38689 nor n41034 n41085 ; n41125
g38690 nor n41124 n41125 ; n41126
g38691 nor pi1156 n41126 ; n41127
g38692 and n41095 n41120 ; n41128
g38693 and pi1155 n41128_not ; n41129
g38694 and n41127 n41129_not ; n41130
g38695 nor pi1157 n41123 ; n41131
g38696 and n41130_not n41131 ; n41132
g38697 nor pi0211 n41132 ; n41133
g38698 and n41113_not n41133 ; n41134
g38699 and n41018 n41087_not ; n41135
g38700 and n40930 n40979 ; n41136
g38701 nor n41135 n41136 ; n41137
g38702 and n41127 n41137 ; n41138
g38703 nor pi1157 n41122 ; n41139
g38704 and n41138_not n41139 ; n41140
g38705 and n41090 n41135_not ; n41141
g38706 and n41073_not n41110 ; n41142
g38707 and pi1156 n41142_not ; n41143
g38708 and pi1157 n41141_not ; n41144
g38709 and n41143_not n41144 ; n41145
g38710 and pi0211 n41140_not ; n41146
g38711 and n41145_not n41146 ; n41147
g38712 nor pi0219 n41134 ; n41148
g38713 and n41147_not n41148 ; n41149
g38714 and n40861 n41083_not ; n41150
g38715 and n41149_not n41150 ; n41151
g38716 nor po1038 n40978 ; n41152
g38717 and n41151_not n41152 ; n41153
g38718 and n40907_not n40910 ; n41154
g38719 and n41153_not n41154 ; n41155
g38720 and po1038_not n40977 ; n41156
g38721 and po1038 n40904 ; n41157
g38722 nor n40910 n41157 ; n41158
g38723 and n41156_not n41158 ; n41159
g38724 nor pi0230 n41159 ; n41160
g38725 and n41155_not n41160 ; n41161
g38726 nor n16479 n40902 ; n41162
g38727 and pi0199 n39467_not ; n41163
g38728 nor n38840 n40946 ; n41164
g38729 and n41163_not n41164 ; n41165
g38730 and n16479 n41165 ; n41166
g38731 and pi0230 n41162_not ; n41167
g38732 and n41166_not n41167 ; n41168
g38733 nor n41161 n41168 ; po0400
g38734 nor pi0230 pi0244 ; n41170
g38735 and pi0213 n40405_not ; n41171
g38736 nor pi0211 n38543 ; n41172
g38737 and n40357_not n41172 ; n41173
g38738 nor n40346 n41173 ; n41174
g38739 and n40344 n41174_not ; n41175
g38740 and n38610_not n40390 ; n41176
g38741 nor n40383 n41176 ; n41177
g38742 nor n40411 n41177 ; n41178
g38743 and pi0214 n41178_not ; n41179
g38744 and n40364 n41179_not ; n41180
g38745 and n38420 n40293 ; n41181
g38746 and pi0214_not n41177 ; n41182
g38747 and pi0212 n41181_not ; n41183
g38748 and n41182_not n41183 ; n41184
g38749 and n40411_not n41184 ; n41185
g38750 nor pi0219 n41180 ; n41186
g38751 and n41185_not n41186 ; n41187
g38752 and n40447 n41175_not ; n41188
g38753 and n41187_not n41188 ; n41189
g38754 and pi0299 n39410 ; n41190
g38755 and pi0214 n41177 ; n41191
g38756 and n40388 n41191_not ; n41192
g38757 and n40381_not n41184 ; n41193
g38758 nor pi0219 n41192 ; n41194
g38759 and n41193_not n41194 ; n41195
g38760 and pi1147 n41190_not ; n41196
g38761 and n40410 n41196 ; n41197
g38762 and n41195_not n41197 ; n41198
g38763 nor pi0213 n39420 ; n41199
g38764 and n41198_not n41199 ; n41200
g38765 and n41189_not n41200 ; n41201
g38766 nor n41171 n41201 ; n41202
g38767 and pi0209 n41202_not ; n41203
g38768 nor pi0213 n39427 ; n41204
g38769 and n40244 n40247_not ; n41205
g38770 nor n40224 n41205 ; n41206
g38771 and n10843_not n40236 ; n41207
g38772 and n10843 n40231_not ; n41208
g38773 and n40244 n40246_not ; n41209
g38774 and n38665 n41207_not ; n41210
g38775 and n41208_not n41210 ; n41211
g38776 and n41209_not n41211 ; n41212
g38777 nor n39398 n40253 ; n41213
g38778 and n41212_not n41213 ; n41214
g38779 nor po1038 n41214 ; n41215
g38780 nor n41206 n41215 ; n41216
g38781 and pi0213 n41216_not ; n41217
g38782 nor pi0209 n41204 ; n41218
g38783 and n41217_not n41218 ; n41219
g38784 nor n41203 n41219 ; n41220
g38785 and pi0230 n41220_not ; n41221
g38786 nor n41170 n41221 ; po0401
g38787 nor pi0213 n40824 ; n41223
g38788 and pi1146 n39869 ; n41224
g38789 nor pi1147 n41224 ; n41225
g38790 and n39865 n40145_not ; n41226
g38791 and n41225 n41226_not ; n41227
g38792 and n38413_not n40800 ; n41228
g38793 and n40819 n41228_not ; n41229
g38794 nor po1038 n41229 ; n41230
g38795 and pi0214 n40235_not ; n41231
g38796 nor pi0299 n40804 ; n41232
g38797 and n41231 n41232_not ; n41233
g38798 and pi0212 n41233_not ; n41234
g38799 and pi0299_not n40802 ; n41235
g38800 nor pi0211 n41235 ; n41236
g38801 and n40794 n41236_not ; n41237
g38802 and pi0214_not n41237 ; n41238
g38803 and n41234 n41238_not ; n41239
g38804 and n40796 n41237_not ; n41240
g38805 nor pi0219 n41240 ; n41241
g38806 and n41239_not n41241 ; n41242
g38807 and n41230 n41242_not ; n41243
g38808 and n41227 n41243_not ; n41244
g38809 and pi1147 n39865_not ; n41245
g38810 and n41224_not n41245 ; n41246
g38811 and pi0211 n40799_not ; n41247
g38812 nor n41236 n41247 ; n41248
g38813 and pi0214 n41248_not ; n41249
g38814 nor pi0214 n41235 ; n41250
g38815 nor n41249 n41250 ; n41251
g38816 and pi0212 n41251_not ; n41252
g38817 and n40796 n41235_not ; n41253
g38818 nor pi0219 n41253 ; n41254
g38819 and n41252_not n41254 ; n41255
g38820 and n41230 n41255_not ; n41256
g38821 and n41246 n41256_not ; n41257
g38822 and pi1148 n41244_not ; n41258
g38823 and n41257_not n41258 ; n41259
g38824 nor n40407 n41246 ; n41260
g38825 and n13061_not n40794 ; n41261
g38826 nor pi0214 n41261 ; n41262
g38827 nor n41249 n41262 ; n41263
g38828 and pi0212 n41263_not ; n41264
g38829 and n40796 n41261_not ; n41265
g38830 nor pi0219 n41265 ; n41266
g38831 and n41264_not n41266 ; n41267
g38832 and n41230 n41267_not ; n41268
g38833 nor n41260 n41268 ; n41269
g38834 and n40795_not n41234 ; n41270
g38835 nor pi0212 n40794 ; n41271
g38836 nor pi0219 n41271 ; n41272
g38837 and n41270_not n41272 ; n41273
g38838 and n41230 n41273_not ; n41274
g38839 and n41225 n41274_not ; n41275
g38840 nor pi1148 n41269 ; n41276
g38841 and n41275_not n41276 ; n41277
g38842 nor n41259 n41277 ; n41278
g38843 and pi0213 n41278_not ; n41279
g38844 nor pi0209 n41223 ; n41280
g38845 and n41279_not n41280 ; n41281
g38846 and pi0199 pi1146 ; n41282
g38847 and n38699 n41282_not ; n41283
g38848 and n38550 n41283_not ; n41284
g38849 nor n10487 n41284 ; n41285
g38850 and n40339 n41283_not ; n41286
g38851 and pi0207 n41286 ; n41287
g38852 nor n38826 n41287 ; n41288
g38853 nor n41285 n41288 ; n41289
g38854 and n38414_not n41289 ; n41290
g38855 and pi0219 n41290_not ; n41291
g38856 and n38449 n41284 ; n41292
g38857 and pi0208 n41286 ; n41293
g38858 nor pi0200 n41282 ; n41294
g38859 and n38550 n41294_not ; n41295
g38860 and pi0207_not n41295 ; n41296
g38861 nor n40234 n41296 ; n41297
g38862 and n41287_not n41297 ; n41298
g38863 and pi0208 n41298_not ; n41299
g38864 and pi0299_not n41299 ; n41300
g38865 nor n41292 n41293 ; n41301
g38866 and n41300_not n41301 ; n41302
g38867 and n40234_not n41302 ; n41303
g38868 and n38414 n41303_not ; n41304
g38869 and n41291 n41304_not ; n41305
g38870 nor pi0214 n41289 ; n41306
g38871 nor pi0212 n41306 ; n41307
g38872 and pi0299_not n41302 ; n41308
g38873 and n41307 n41308_not ; n41309
g38874 nor pi0219 n41309 ; n41310
g38875 and pi0212 n41308_not ; n41311
g38876 and n10484 n41303 ; n41312
g38877 and n41311 n41312_not ; n41313
g38878 and n41310 n41313_not ; n41314
g38879 nor po1038 n41305 ; n41315
g38880 and n41314_not n41315 ; n41316
g38881 and n41246 n41316_not ; n41317
g38882 and pi0208_not n40234 ; n41318
g38883 and n40339 n41294_not ; n41319
g38884 and pi0207 n41319 ; n41320
g38885 and pi1146 n38700_not ; n41321
g38886 nor n41320 n41321 ; n41322
g38887 and pi0208 n41322_not ; n41323
g38888 nor pi0207 n41293 ; n41324
g38889 and n39658 n41283_not ; n41325
g38890 and n41324_not n41325 ; n41326
g38891 nor n41318 n41323 ; n41327
g38892 and n41326_not n41327 ; n41328
g38893 nor pi0299 n41328 ; n41329
g38894 nor pi0214 n41329 ; n41330
g38895 nor pi0212 n41330 ; n41331
g38896 nor n10487 n39659 ; n41332
g38897 and n41319 n41332_not ; n41333
g38898 and pi0211 n41333_not ; n41334
g38899 nor pi0299 n41319 ; n41335
g38900 nor n41328 n41335 ; n41336
g38901 nor pi0299 n41336 ; n41337
g38902 and pi0211_not n41337 ; n41338
g38903 nor n41334 n41338 ; n41339
g38904 nor n41329 n41339 ; n41340
g38905 and n41331 n41340_not ; n41341
g38906 nor pi0219 n41341 ; n41342
g38907 and n41231 n41329_not ; n41343
g38908 and pi0214_not n41340 ; n41344
g38909 and pi0212 n41344_not ; n41345
g38910 and n41343_not n41345 ; n41346
g38911 and n41342 n41346_not ; n41347
g38912 and n38414_not n41329 ; n41348
g38913 and pi0219 n41348_not ; n41349
g38914 and n38414 n41328_not ; n41350
g38915 and n41349 n41350_not ; n41351
g38916 nor po1038 n41351 ; n41352
g38917 and n41347_not n41352 ; n41353
g38918 and n41227 n41353_not ; n41354
g38919 and pi1148 n41317_not ; n41355
g38920 and n41354_not n41355 ; n41356
g38921 nor n40663 n41329 ; n41357
g38922 nor n41322 n41357 ; n41358
g38923 nor pi0219 n41358 ; n41359
g38924 and pi0219 n41333_not ; n41360
g38925 nor n38970 n41360 ; n41361
g38926 nor n38413 n41334 ; n41362
g38927 and n41336 n41362 ; n41363
g38928 nor n41361 n41363 ; n41364
g38929 nor po1038 n41364 ; n41365
g38930 and n41359_not n41365 ; n41366
g38931 and n41225 n41366_not ; n41367
g38932 nor n10487 n41295 ; n41368
g38933 nor n41288 n41368 ; n41369
g38934 nor n13061 n41369 ; n41370
g38935 and pi0214 n41370_not ; n41371
g38936 and pi0214_not n41369 ; n41372
g38937 nor pi0212 n41372 ; n41373
g38938 and n41371_not n41373 ; n41374
g38939 nor pi0214 n41370 ; n41375
g38940 and n38449 n41295 ; n41376
g38941 nor n41318 n41376 ; n41377
g38942 and n41299_not n41377 ; n41378
g38943 and pi0299_not n41378 ; n41379
g38944 and pi0214 n41379_not ; n41380
g38945 nor pi0211 n41308 ; n41381
g38946 nor n41289 n41381 ; n41382
g38947 and n41380 n41382_not ; n41383
g38948 and pi0212 n41383_not ; n41384
g38949 and n41375_not n41384 ; n41385
g38950 nor n41374 n41385 ; n41386
g38951 nor pi0219 n41386 ; n41387
g38952 nor pi1146 n38783 ; n41388
g38953 and n40299 n41388_not ; n41389
g38954 and n41387 n41389_not ; n41390
g38955 and n38413_not n41369 ; n41391
g38956 nor n38414 n41391 ; n41392
g38957 nor n41378 n41392 ; n41393
g38958 and pi0212_not n41372 ; n41394
g38959 and pi0219 n41394_not ; n41395
g38960 and n41393_not n41395 ; n41396
g38961 nor po1038 n41396 ; n41397
g38962 and n41390_not n41397 ; n41398
g38963 nor n41260 n41398 ; n41399
g38964 nor pi1148 n41367 ; n41400
g38965 and n41399_not n41400 ; n41401
g38966 nor n41356 n41401 ; n41402
g38967 and pi0213 n41402_not ; n41403
g38968 and pi1147 po1038_not ; n41404
g38969 and n38612_not n41302 ; n41405
g38970 and n38414 n41405_not ; n41406
g38971 and n41291 n41406_not ; n41407
g38972 and n40231_not n41302 ; n41408
g38973 and pi0214 n41408 ; n41409
g38974 and n41307 n41409_not ; n41410
g38975 and pi0299 n40774_not ; n41411
g38976 and n41302 n41411_not ; n41412
g38977 and pi0212 n41412_not ; n41413
g38978 nor pi0219 n41413 ; n41414
g38979 and n41410_not n41414 ; n41415
g38980 and n41404 n41407_not ; n41416
g38981 and n41415_not n41416 ; n41417
g38982 and pi0299_not n41328 ; n41418
g38983 and n38414 n41418_not ; n41419
g38984 and n38610_not n41419 ; n41420
g38985 and n41349 n41420_not ; n41421
g38986 nor n40231 n41329 ; n41422
g38987 and n41331 n41422_not ; n41423
g38988 nor n41329 n41411 ; n41424
g38989 and pi0212 n41424_not ; n41425
g38990 nor pi0219 n41425 ; n41426
g38991 and n41423_not n41426 ; n41427
g38992 and n40447 n41421_not ; n41428
g38993 and n41427_not n41428 ; n41429
g38994 and pi1148 n40780_not ; n41430
g38995 and n41417_not n41430 ; n41431
g38996 and n41429_not n41431 ; n41432
g38997 and n41379_not n41413 ; n41433
g38998 and n41380 n41408_not ; n41434
g38999 nor n41372 n41434 ; n41435
g39000 nor pi0212 n41435 ; n41436
g39001 nor pi0219 n41433 ; n41437
g39002 and n41436_not n41437 ; n41438
g39003 nor n41379 n41405 ; n41439
g39004 nor pi0211 n41439 ; n41440
g39005 nor n41392 n41440 ; n41441
g39006 and n41395 n41441_not ; n41442
g39007 and n41404 n41438_not ; n41443
g39008 and n41442_not n41443 ; n41444
g39009 and n41335_not n41425 ; n41445
g39010 and pi0214_not n41333 ; n41446
g39011 and pi0214 n41337_not ; n41447
g39012 and n41422_not n41447 ; n41448
g39013 nor n41446 n41448 ; n41449
g39014 nor pi0212 n41449 ; n41450
g39015 nor pi0219 n41445 ; n41451
g39016 and n41450_not n41451 ; n41452
g39017 nor n38610 n41337 ; n41453
g39018 nor pi0211 n41453 ; n41454
g39019 and n41362 n41454_not ; n41455
g39020 nor n41361 n41455 ; n41456
g39021 and n40447 n41456_not ; n41457
g39022 and n41452_not n41457 ; n41458
g39023 nor pi1148 n40780 ; n41459
g39024 and n41444_not n41459 ; n41460
g39025 and n41458_not n41460 ; n41461
g39026 nor pi0213 n41432 ; n41462
g39027 and n41461_not n41462 ; n41463
g39028 and pi0209 n41463_not ; n41464
g39029 and n41403_not n41464 ; n41465
g39030 nor n41281 n41465 ; n41466
g39031 and pi0230 n41466_not ; n41467
g39032 nor pi0230 pi0245 ; n41468
g39033 nor n41467 n41468 ; po0402
g39034 and pi1150_not n40134 ; n41470
g39035 and pi1150 n40089 ; n41471
g39036 and pi1149 n41470_not ; n41472
g39037 and n41471_not n41472 ; n41473
g39038 and pi1150_not n40200 ; n41474
g39039 and pi1150 n40166 ; n41475
g39040 nor pi1149 n41474 ; n41476
g39041 and n41475_not n41476 ; n41477
g39042 nor n41473 n41477 ; n41478
g39043 and pi1148 n41478_not ; n41479
g39044 and pi1150_not n40125 ; n41480
g39045 and pi1150 n40078 ; n41481
g39046 and pi1149 n41481_not ; n41482
g39047 and n41480_not n41482 ; n41483
g39048 and pi1149_not pi1150 ; n41484
g39049 and n40143_not n41484 ; n41485
g39050 nor n41483 n41485 ; n41486
g39051 nor pi1148 n41486 ; n41487
g39052 nor n41479 n41487 ; n41488
g39053 and pi0213 n41488_not ; n41489
g39054 nor n40184 n40193 ; n41490
g39055 and n41227 n41490_not ; n41491
g39056 nor n41227 n41246 ; n41492
g39057 and pi0219 n40234_not ; n41493
g39058 and n40084 n41493_not ; n41494
g39059 and n40127 n40181_not ; n41495
g39060 nor n41494 n41495 ; n41496
g39061 nor n40183 n40255 ; n41497
g39062 and n38423 n41497_not ; n41498
g39063 nor n40648 n41498 ; n41499
g39064 nor pi0219 n41499 ; n41500
g39065 nor n41496 n41500 ; n41501
g39066 nor n41492 n41501 ; n41502
g39067 nor pi1150 n41491 ; n41503
g39068 and n41502_not n41503 ; n41504
g39069 nor n40269 n41494 ; n41505
g39070 and pi0214_not n39697 ; n41506
g39071 and pi0214 n40147_not ; n41507
g39072 and n40274_not n41507 ; n41508
g39073 and pi0212 n41506_not ; n41509
g39074 and n41508_not n41509 ; n41510
g39075 and n40156 n41510_not ; n41511
g39076 nor n41505 n41511 ; n41512
g39077 and n41227 n41512_not ; n41513
g39078 and n40276_not n40513 ; n41514
g39079 nor pi0212 n39661 ; n41515
g39080 nor pi0219 n41515 ; n41516
g39081 and n40525_not n41516 ; n41517
g39082 and n41514_not n41517 ; n41518
g39083 nor n41505 n41518 ; n41519
g39084 and n41246 n41519_not ; n41520
g39085 and pi1150 n41513_not ; n41521
g39086 and n41520_not n41521 ; n41522
g39087 nor n41504 n41522 ; n41523
g39088 and pi1148 n41523_not ; n41524
g39089 and pi1150 n39639 ; n41525
g39090 and pi0299 n40093 ; n41526
g39091 nor pi0219 n41526 ; n41527
g39092 and n41389_not n41527 ; n41528
g39093 and n41525_not n41528 ; n41529
g39094 and n41260_not n41529 ; n41530
g39095 nor pi0219 n40213 ; n41531
g39096 nor n40664 n41531 ; n41532
g39097 and n41494 n41532 ; n41533
g39098 and n41225 n41533_not ; n41534
g39099 nor n41260 n41494 ; n41535
g39100 nor n41534 n41535 ; n41536
g39101 and pi1150 n40140 ; n41537
g39102 nor n41536 n41537 ; n41538
g39103 nor pi1148 n41530 ; n41539
g39104 and n41538_not n41539 ; n41540
g39105 nor n41524 n41540 ; n41541
g39106 nor pi1149 n41541 ; n41542
g39107 and pi1146_not n40122 ; n41543
g39108 and n40084 n40105_not ; n41544
g39109 nor n40123 n41544 ; n41545
g39110 and n40213 n40293 ; n41546
g39111 nor n40100 n41546 ; n41547
g39112 and n40121 n41547 ; n41548
g39113 nor n41543 n41545 ; n41549
g39114 and n41548_not n41549 ; n41550
g39115 nor n41260 n41550 ; n41551
g39116 nor n40102 n40524 ; n41552
g39117 nor pi0219 n41552 ; n41553
g39118 nor n41545 n41553 ; n41554
g39119 nor pi1146 n40100 ; n41555
g39120 and n41554 n41555_not ; n41556
g39121 and n41225 n41556_not ; n41557
g39122 nor pi1150 n41557 ; n41558
g39123 and n41551_not n41558 ; n41559
g39124 nor n40311 n41494 ; n41560
g39125 nor n40062 n40725 ; n41561
g39126 and pi0214_not n40725 ; n41562
g39127 and n40074 n41562_not ; n41563
g39128 nor pi0219 n41563 ; n41564
g39129 and n41561_not n41564 ; n41565
g39130 and pi0212_not n41561 ; n41566
g39131 and n41564 n41566_not ; n41567
g39132 and pi0299_not n39713 ; n41568
g39133 nor n40064 n40234 ; n41569
g39134 and n41568_not n41569 ; n41570
g39135 and n41567 n41570 ; n41571
g39136 nor n41560 n41565 ; n41572
g39137 and n41571_not n41572 ; n41573
g39138 nor n40060 n41573 ; n41574
g39139 and n40063 n40073_not ; n41575
g39140 nor pi0219 n41575 ; n41576
g39141 and n40729_not n41576 ; n41577
g39142 and n40310 n41577_not ; n41578
g39143 and n41574_not n41578 ; n41579
g39144 and n41225 n41579_not ; n41580
g39145 nor n41260 n41573 ; n41581
g39146 and pi1150 n41581_not ; n41582
g39147 and n41580_not n41582 ; n41583
g39148 nor pi1148 n41583 ; n41584
g39149 and n41559_not n41584 ; n41585
g39150 nor n40127 n41494 ; n41586
g39151 and n39747 n41231 ; n41587
g39152 and n40189 n41587_not ; n41588
g39153 and n40172_not n40190 ; n41589
g39154 nor n40177 n41589 ; n41590
g39155 nor n41227 n41590 ; n41591
g39156 and n40192 n41588_not ; n41592
g39157 and n41591_not n41592 ; n41593
g39158 nor n41586 n41593 ; n41594
g39159 nor n41492 n41594 ; n41595
g39160 nor pi1150 n41595 ; n41596
g39161 nor n40303 n41533 ; n41597
g39162 and n41227 n41597 ; n41598
g39163 and pi0214 n40292 ; n41599
g39164 and n40298 n41599_not ; n41600
g39165 nor pi0219 n40295 ; n41601
g39166 and n41600_not n41601 ; n41602
g39167 and n40291 n41602_not ; n41603
g39168 and pi1146 n40085 ; n41604
g39169 and n41246 n41604_not ; n41605
g39170 and n41603_not n41605 ; n41606
g39171 and pi1150 n41606_not ; n41607
g39172 and n41598_not n41607 ; n41608
g39173 and pi1148 n41608_not ; n41609
g39174 and n41596_not n41609 ; n41610
g39175 and pi1149 n41610_not ; n41611
g39176 and n41585_not n41611 ; n41612
g39177 nor n41542 n41612 ; n41613
g39178 nor pi0213 n41613 ; n41614
g39179 and pi0209 n41489_not ; n41615
g39180 and n41614_not n41615 ; n41616
g39181 nor pi0213 n41402 ; n41617
g39182 and pi0219 n41369_not ; n41618
g39183 and n41404 n41618_not ; n41619
g39184 and n41387_not n41619 ; n41620
g39185 nor pi0212 n41446 ; n41621
g39186 nor n13061 n41333 ; n41622
g39187 and pi0214 n41622_not ; n41623
g39188 and n41621 n41623_not ; n41624
g39189 nor pi0214 n41622 ; n41625
g39190 and pi0214 n41339 ; n41626
g39191 and pi0212 n41626_not ; n41627
g39192 and n41625_not n41627 ; n41628
g39193 nor n41624 n41628 ; n41629
g39194 nor pi0219 n41629 ; n41630
g39195 and n40447 n41360_not ; n41631
g39196 and n41630_not n41631 ; n41632
g39197 nor pi1150 n40096 ; n41633
g39198 and n41620_not n41633 ; n41634
g39199 and n41632_not n41634 ; n41635
g39200 and n41373 n41380_not ; n41636
g39201 nor pi0214 n41379 ; n41637
g39202 and n41384 n41637_not ; n41638
g39203 nor n41636 n41638 ; n41639
g39204 nor pi0219 n41639 ; n41640
g39205 nor n41618 n41640 ; n41641
g39206 and pi1147 n41641_not ; n41642
g39207 and n41447_not n41621 ; n41643
g39208 nor pi0214 n41337 ; n41644
g39209 and n41627 n41644_not ; n41645
g39210 nor n41643 n41645 ; n41646
g39211 nor pi0219 n41646 ; n41647
g39212 nor n41360 n41647 ; n41648
g39213 nor pi1147 n41648 ; n41649
g39214 nor po1038 n41642 ; n41650
g39215 and n41649_not n41650 ; n41651
g39216 and pi1150 n39865_not ; n41652
g39217 and n41651_not n41652 ; n41653
g39218 nor n41635 n41653 ; n41654
g39219 and pi1149 n41654_not ; n41655
g39220 and pi1150 n40207 ; n41656
g39221 and n41333 n41656_not ; n41657
g39222 nor pi1147 n41657 ; n41658
g39223 and pi1147 n41369_not ; n41659
g39224 nor po1038 n41658 ; n41660
g39225 and n41659_not n41660 ; n41661
g39226 and pi1147_not n41336 ; n41662
g39227 and n16479 n41662_not ; n41663
g39228 and n41656 n41663_not ; n41664
g39229 nor pi1149 n41661 ; n41665
g39230 and n41664_not n41665 ; n41666
g39231 nor n41655 n41666 ; n41667
g39232 nor pi1148 n41667 ; n41668
g39233 and n38413_not n41381 ; n41669
g39234 and n41291 n41669_not ; n41670
g39235 and n41404 n41670_not ; n41671
g39236 and pi0214 n13061_not ; n41672
g39237 and n41302 n41672 ; n41673
g39238 and pi0212 n41673_not ; n41674
g39239 and n41306_not n41674 ; n41675
g39240 and pi0212_not n41289 ; n41676
g39241 nor pi0219 n41676 ; n41677
g39242 and n41675_not n41677 ; n41678
g39243 and n41671 n41678_not ; n41679
g39244 and n41349 n41419_not ; n41680
g39245 and n40447 n41680_not ; n41681
g39246 and pi0219_not n41357 ; n41682
g39247 and n41681 n41682_not ; n41683
g39248 nor pi1150 n39869 ; n41684
g39249 and n41679_not n41684 ; n41685
g39250 and n41683_not n41685 ; n41686
g39251 and n41329_not n41622 ; n41687
g39252 and pi0214 n41687 ; n41688
g39253 and n41345 n41688_not ; n41689
g39254 and n41342 n41689_not ; n41690
g39255 and n41681 n41690_not ; n41691
g39256 and pi0214_not n41382 ; n41692
g39257 and n41674 n41692_not ; n41693
g39258 and n41307 n41382_not ; n41694
g39259 nor pi0219 n41694 ; n41695
g39260 and n41693_not n41695 ; n41696
g39261 and n41671 n41696_not ; n41697
g39262 and pi1150 n40146_not ; n41698
g39263 and n41697_not n41698 ; n41699
g39264 and n41691_not n41699 ; n41700
g39265 nor pi1149 n41686 ; n41701
g39266 and n41700_not n41701 ; n41702
g39267 and pi0057 n38666 ; n41703
g39268 nor n6305 n38666 ; n41704
g39269 and n41310 n41311_not ; n41705
g39270 nor n41670 n41705 ; n41706
g39271 and n6305 n41706 ; n41707
g39272 and pi0057_not pi1147 ; n41708
g39273 and n41704_not n41708 ; n41709
g39274 and n41707_not n41709 ; n41710
g39275 and n6305 n38665_not ; n41711
g39276 and n41348 n41711 ; n41712
g39277 nor n38666 n41418 ; n41713
g39278 nor pi0057 pi1147 ; n41714
g39279 and n41704_not n41714 ; n41715
g39280 and n41713_not n41715 ; n41716
g39281 and n41712_not n41716 ; n41717
g39282 nor n41703 n41717 ; n41718
g39283 and n41710_not n41718 ; n41719
g39284 and pi1150 n41719_not ; n41720
g39285 and n41331 n41688_not ; n41721
g39286 and n41447_not n41687 ; n41722
g39287 and pi0212 n41722_not ; n41723
g39288 nor pi0219 n41721 ; n41724
g39289 and n41723_not n41724 ; n41725
g39290 and n41681 n41725_not ; n41726
g39291 and n40676_not n41404 ; n41727
g39292 and n41706 n41727 ; n41728
g39293 nor pi1150 n40131 ; n41729
g39294 and n41728_not n41729 ; n41730
g39295 and n41726_not n41730 ; n41731
g39296 and pi1149 n41731_not ; n41732
g39297 and n41720_not n41732 ; n41733
g39298 and pi1148 n41733_not ; n41734
g39299 and n41702_not n41734 ; n41735
g39300 and pi0213 n41735_not ; n41736
g39301 and n41668_not n41736 ; n41737
g39302 nor pi0209 n41617 ; n41738
g39303 and n41737_not n41738 ; n41739
g39304 nor n41616 n41739 ; n41740
g39305 and pi0230 n41740_not ; n41741
g39306 nor pi0230 pi0246 ; n41742
g39307 nor n41741 n41742 ; po0403
g39308 and pi0213 n40625 ; n41744
g39309 and pi1151 n40131_not ; n41745
g39310 and n40310 n41565_not ; n41746
g39311 and n41745 n41746_not ; n41747
g39312 and n40104 n40119_not ; n41748
g39313 nor n41545 n41748 ; n41749
g39314 nor n40131 n41749 ; n41750
g39315 and pi1151_not n41750 ; n41751
g39316 and pi1147 n41747_not ; n41752
g39317 and n41751_not n41752 ; n41753
g39318 nor pi1147 n40609 ; n41754
g39319 and pi1151 n40096_not ; n41755
g39320 nor n40061 n41567 ; n41756
g39321 and n41755 n41756_not ; n41757
g39322 and n41754 n41757_not ; n41758
g39323 nor pi1149 n41753 ; n41759
g39324 and n41758_not n41759 ; n41760
g39325 and pi1147 n40615_not ; n41761
g39326 nor n40082 n40085 ; n41762
g39327 and n40672 n41762 ; n41763
g39328 and n41761 n41763_not ; n41764
g39329 nor pi1151 n39865 ; n41765
g39330 and n40192 n41589_not ; n41766
g39331 and n40680 n41766_not ; n41767
g39332 and n40178_not n40680 ; n41768
g39333 nor n41767 n41768 ; n41769
g39334 and n41765 n41769 ; n41770
g39335 and n40500 n41603_not ; n41771
g39336 nor pi1147 n41771 ; n41772
g39337 and n41770_not n41772 ; n41773
g39338 and pi1149 n41764_not ; n41774
g39339 and n41773_not n41774 ; n41775
g39340 and pi1150 n41775_not ; n41776
g39341 and n41760_not n41776 ; n41777
g39342 and n40095_not n40141 ; n41778
g39343 nor pi1151 n41778 ; n41779
g39344 nor pi1147 n41779 ; n41780
g39345 and n39830 n40533_not ; n41781
g39346 and n41755 n41781_not ; n41782
g39347 and n41780 n41782_not ; n41783
g39348 and n40704_not n41745 ; n41784
g39349 and n40132_not n40577 ; n41785
g39350 and pi1147 n41785_not ; n41786
g39351 and n41784_not n41786 ; n41787
g39352 nor pi1149 n41783 ; n41788
g39353 and n41787_not n41788 ; n41789
g39354 and pi0212 n39686_not ; n41790
g39355 and n41517 n41790_not ; n41791
g39356 and n40164 n41791_not ; n41792
g39357 and n40593 n41792_not ; n41793
g39358 and pi1147 n41793_not ; n41794
g39359 and n38423 n40173_not ; n41795
g39360 and n40183_not n40653 ; n41796
g39361 and n41795_not n41796 ; n41797
g39362 nor pi1151 n40082 ; n41798
g39363 and n41797_not n41798 ; n41799
g39364 and n40198_not n41799 ; n41800
g39365 and n41794 n41800_not ; n41801
g39366 and n41765 n41797_not ; n41802
g39367 and n40514_not n41517 ; n41803
g39368 and n40269 n41803_not ; n41804
g39369 nor n39865 n41804 ; n41805
g39370 and pi1151 n41805 ; n41806
g39371 nor pi1147 n41802 ; n41807
g39372 and n41806_not n41807 ; n41808
g39373 and pi1149 n41808_not ; n41809
g39374 and n41801_not n41809 ; n41810
g39375 nor pi1150 n41789 ; n41811
g39376 and n41810_not n41811 ; n41812
g39377 nor n41777 n41812 ; n41813
g39378 and pi1148 n41813_not ; n41814
g39379 nor pi1151 n40243 ; n41815
g39380 nor pi1147 n41815 ; n41816
g39381 and pi1151 n40060_not ; n41817
g39382 and n41816 n41817_not ; n41818
g39383 and n41577_not n41746 ; n41819
g39384 and n39870 n41819_not ; n41820
g39385 nor n39869 n41554 ; n41821
g39386 and pi1151_not n41821 ; n41822
g39387 and pi1147 n41822_not ; n41823
g39388 and n41820_not n41823 ; n41824
g39389 and pi1150 n41818_not ; n41825
g39390 and n41824_not n41825 ; n41826
g39391 and pi1147_not pi1151 ; n41827
g39392 and n40140 n41827 ; n41828
g39393 and n39639_not n40664 ; n41829
g39394 and n40696 n41829_not ; n41830
g39395 and n39870 n41830_not ; n41831
g39396 and n40565 n40665_not ; n41832
g39397 and pi1147 n41832_not ; n41833
g39398 and n41831_not n41833 ; n41834
g39399 nor pi1150 n41828 ; n41835
g39400 and n41834_not n41835 ; n41836
g39401 nor n41826 n41836 ; n41837
g39402 nor pi1149 n41837 ; n41838
g39403 nor pi1151 n40208 ; n41839
g39404 and n40637_not n41839 ; n41840
g39405 and n40159_not n40269 ; n41841
g39406 nor n40208 n41841 ; n41842
g39407 and pi1151 n41842 ; n41843
g39408 nor pi1147 n41840 ; n41844
g39409 and n41843_not n41844 ; n41845
g39410 and pi1147 n40620_not ; n41846
g39411 nor pi1151 n40146 ; n41847
g39412 and n40198_not n41847 ; n41848
g39413 and n41846 n41848_not ; n41849
g39414 nor pi1150 n41845 ; n41850
g39415 and n41849_not n41850 ; n41851
g39416 and n40548 n40666 ; n41852
g39417 and pi1147 n41852_not ; n41853
g39418 nor n40146 n40197 ; n41854
g39419 and pi1151_not n41854 ; n41855
g39420 and n41853 n41855_not ; n41856
g39421 and n41767_not n41839 ; n41857
g39422 and pi1151 n40208_not ; n41858
g39423 and n40303_not n41858 ; n41859
g39424 nor pi1147 n41859 ; n41860
g39425 and n41857_not n41860 ; n41861
g39426 and pi1150 n41856_not ; n41862
g39427 and n41861_not n41862 ; n41863
g39428 nor n41851 n41863 ; n41864
g39429 and pi1149 n41864_not ; n41865
g39430 nor pi1148 n41838 ; n41866
g39431 and n41865_not n41866 ; n41867
g39432 nor n41814 n41867 ; n41868
g39433 nor pi0213 n41868 ; n41869
g39434 and pi0209 n41744_not ; n41870
g39435 and n41869_not n41870 ; n41871
g39436 nor pi0213 n40205 ; n41872
g39437 and n41767_not n41858 ; n41873
g39438 and pi1147 n40672_not ; n41874
g39439 and n41873_not n41874 ; n41875
g39440 nor po1038 n40711 ; n41876
g39441 and n40714_not n41876 ; n41877
g39442 nor n40485 n41877 ; n41878
g39443 and n41816 n41878 ; n41879
g39444 nor pi1150 n41879 ; n41880
g39445 and n41875_not n41880 ; n41881
g39446 and n40500 n41769 ; n41882
g39447 and n40523 n41768_not ; n41883
g39448 and pi1147 n41883_not ; n41884
g39449 and n41882_not n41884 ; n41885
g39450 and n40116 n40123 ; n41886
g39451 and n40500 n41886_not ; n41887
g39452 and n41754 n41887_not ; n41888
g39453 and pi1150 n41885_not ; n41889
g39454 and n41888_not n41889 ; n41890
g39455 nor n41881 n41890 ; n41891
g39456 nor pi1149 n41891 ; n41892
g39457 and n40565 n41819_not ; n41893
g39458 nor n40146 n41578 ; n41894
g39459 and pi1151 n41894 ; n41895
g39460 nor pi1147 n41895 ; n41896
g39461 and n41893_not n41896 ; n41897
g39462 and n40087_not n41832 ; n41898
g39463 and n41853 n41898_not ; n41899
g39464 nor pi1150 n41899 ; n41900
g39465 and n41897_not n41900 ; n41901
g39466 nor n40131 n40677 ; n41902
g39467 and pi1151_not n41902 ; n41903
g39468 and n41761 n41903_not ; n41904
g39469 and n40577 n41746_not ; n41905
g39470 and n40069 n40315_not ; n41906
g39471 and n40310 n41906_not ; n41907
g39472 and n40593 n41907_not ; n41908
g39473 nor pi1147 n41908 ; n41909
g39474 and n41905_not n41909 ; n41910
g39475 and pi1150 n41904_not ; n41911
g39476 and n41910_not n41911 ; n41912
g39477 nor n41901 n41912 ; n41913
g39478 and pi1149 n41913_not ; n41914
g39479 and pi1148 n41914_not ; n41915
g39480 and n41892_not n41915 ; n41916
g39481 and n16479_not n39864 ; n41917
g39482 and pi1151 n41917_not ; n41918
g39483 and n41780 n41918_not ; n41919
g39484 and n40500 n41797_not ; n41920
g39485 and n40185 n40653 ; n41921
g39486 nor n40096 n41921 ; n41922
g39487 and pi1151_not n41922 ; n41923
g39488 and pi1147 n41920_not ; n41924
g39489 and n41923_not n41924 ; n41925
g39490 and pi1150 n41919_not ; n41926
g39491 and n41925_not n41926 ; n41927
g39492 and n40142 n41827 ; n41928
g39493 nor n40208 n40637 ; n41929
g39494 nor pi1151 n41495 ; n41930
g39495 and pi1147 n41930_not ; n41931
g39496 and n41929_not n41931 ; n41932
g39497 nor pi1150 n41928 ; n41933
g39498 and n41932_not n41933 ; n41934
g39499 nor n41927 n41934 ; n41935
g39500 nor pi1149 n41935 ; n41936
g39501 and n39642 n39830 ; n41937
g39502 and n10843_not n41937 ; n41938
g39503 nor n41830 n41938 ; n41939
g39504 and n40548 n41939 ; n41940
g39505 and n40565 n41830_not ; n41941
g39506 nor pi1147 n41941 ; n41942
g39507 and n41940_not n41942 ; n41943
g39508 nor pi0219 n40531 ; n41944
g39509 and n40642_not n41944 ; n41945
g39510 and n40164 n41945_not ; n41946
g39511 and n40160_not n41946 ; n41947
g39512 and n40565 n41947_not ; n41948
g39513 and n41846 n41948_not ; n41949
g39514 nor pi1150 n41943 ; n41950
g39515 and n41949_not n41950 ; n41951
g39516 and n40593 n41937_not ; n41952
g39517 and n40704_not n41952 ; n41953
g39518 and n40577 n40704_not ; n41954
g39519 nor pi1147 n41953 ; n41955
g39520 and n41954_not n41955 ; n41956
g39521 nor n40131 n41946 ; n41957
g39522 and pi1151_not n41957 ; n41958
g39523 and n41794 n41958_not ; n41959
g39524 and pi1150 n41956_not ; n41960
g39525 and n41959_not n41960 ; n41961
g39526 nor n41951 n41961 ; n41962
g39527 and pi1149 n41962_not ; n41963
g39528 nor pi1148 n41936 ; n41964
g39529 and n41963_not n41964 ; n41965
g39530 nor n41916 n41965 ; n41966
g39531 and pi0213 n41966_not ; n41967
g39532 nor pi0209 n41872 ; n41968
g39533 and n41967_not n41968 ; n41969
g39534 nor n41871 n41969 ; n41970
g39535 and pi0230 n41970_not ; n41971
g39536 nor pi0230 pi0247 ; n41972
g39537 nor n41971 n41972 ; po0404
g39538 nor pi1151 n40142 ; n41974
g39539 and n40140_not n41974 ; n41975
g39540 and pi1152 n41975_not ; n41976
g39541 and n40610_not n41976 ; n41977
g39542 and pi1151 pi1152_not ; n41978
g39543 and n40125_not n41978 ; n41979
g39544 nor pi1150 n41977 ; n41980
g39545 and n41979_not n41980 ; n41981
g39546 and pi1151 n40134 ; n41982
g39547 nor pi1152 n41982 ; n41983
g39548 and n40619_not n41983 ; n41984
g39549 and pi1152 n40615_not ; n41985
g39550 and n40165_not n41847 ; n41986
g39551 and n41985 n41986_not ; n41987
g39552 and pi1150 n41984_not ; n41988
g39553 and n41987_not n41988 ; n41989
g39554 nor n41981 n41989 ; n41990
g39555 and pi0213 n41990 ; n41991
g39556 and pi1152 n41954_not ; n41992
g39557 and n41747_not n41992 ; n41993
g39558 and pi1151 n41750 ; n41994
g39559 nor pi1152 n41785 ; n41995
g39560 and n41994_not n41995 ; n41996
g39561 nor pi1150 n41993 ; n41997
g39562 and n41996_not n41997 ; n41998
g39563 and n41792_not n41798 ; n41999
g39564 and n41985 n41999_not ; n42000
g39565 and pi1151 n40127_not ; n42001
g39566 and n41762 n42001 ; n42002
g39567 nor pi1152 n42002 ; n42003
g39568 and n41800_not n42003 ; n42004
g39569 and pi1150 n42004_not ; n42005
g39570 and n42000_not n42005 ; n42006
g39571 and pi1148 n41998_not ; n42007
g39572 and n42006_not n42007 ; n42008
g39573 and n40124_not n41755 ; n42009
g39574 nor pi1152 n42009 ; n42010
g39575 and n41779_not n42010 ; n42011
g39576 and n40523 n41781_not ; n42012
g39577 and pi1152 n42012_not ; n42013
g39578 and n41757_not n42013 ; n42014
g39579 nor pi1150 n42014 ; n42015
g39580 and n42011_not n42015 ; n42016
g39581 and pi1151_not n41805 ; n42017
g39582 and pi1152 n41771_not ; n42018
g39583 and n42017_not n42018 ; n42019
g39584 nor pi1152 n41802 ; n42020
g39585 and n41882_not n42020 ; n42021
g39586 and pi1150 n42019_not ; n42022
g39587 and n42021_not n42022 ; n42023
g39588 nor pi1148 n42023 ; n42024
g39589 and n42016_not n42024 ; n42025
g39590 nor n42008 n42025 ; n42026
g39591 and pi1149 n42026_not ; n42027
g39592 nor pi1152 n41840 ; n42028
g39593 and n41873_not n42028 ; n42029
g39594 and pi1151_not n41842 ; n42030
g39595 and pi1152 n41859_not ; n42031
g39596 and n42030_not n42031 ; n42032
g39597 and pi1150 n42029_not ; n42033
g39598 and n42032_not n42033 ; n42034
g39599 and n40243 n41978 ; n42035
g39600 nor pi1151 n40140 ; n42036
g39601 and pi1152 n41817_not ; n42037
g39602 and n42036_not n42037 ; n42038
g39603 nor pi1150 n42035 ; n42039
g39604 and n42038_not n42039 ; n42040
g39605 nor n42034 n42040 ; n42041
g39606 nor pi1148 n42041 ; n42042
g39607 and pi1152 n41986_not ; n42043
g39608 and n41852_not n42043 ; n42044
g39609 and pi1151 n41854 ; n42045
g39610 nor pi1152 n41848 ; n42046
g39611 and n42045_not n42046 ; n42047
g39612 nor n42044 n42047 ; n42048
g39613 and pi1150 n42048_not ; n42049
g39614 and pi1151 n41821 ; n42050
g39615 nor n41832 n42050 ; n42051
g39616 nor pi1152 n42051 ; n42052
g39617 nor n41820 n41941 ; n42053
g39618 and pi1152 n42053_not ; n42054
g39619 nor pi1150 n42052 ; n42055
g39620 and n42054_not n42055 ; n42056
g39621 and pi1148 n42056_not ; n42057
g39622 and n42049_not n42057 ; n42058
g39623 nor pi1149 n42042 ; n42059
g39624 and n42058_not n42059 ; n42060
g39625 nor n42027 n42060 ; n42061
g39626 nor pi0213 n42061 ; n42062
g39627 and pi0209 n41991_not ; n42063
g39628 and n42062_not n42063 ; n42064
g39629 nor pi0213 n41488 ; n42065
g39630 and n41778 n41978 ; n42066
g39631 and pi1152 n41918_not ; n42067
g39632 and n41974_not n42067 ; n42068
g39633 nor pi1150 n42066 ; n42069
g39634 and n42068_not n42069 ; n42070
g39635 nor pi1152 n41941 ; n42071
g39636 and n41784_not n42071 ; n42072
g39637 and n41847 n41939 ; n42073
g39638 and pi1152 n41953_not ; n42074
g39639 and n42073_not n42074 ; n42075
g39640 and pi1150 n42072_not ; n42076
g39641 and n42075_not n42076 ; n42077
g39642 nor pi1149 n42070 ; n42078
g39643 and n42077_not n42078 ; n42079
g39644 and pi1151_not n41894 ; n42080
g39645 and pi1152 n41908_not ; n42081
g39646 and n42080_not n42081 ; n42082
g39647 nor pi1152 n41747 ; n42083
g39648 and n41893_not n42083 ; n42084
g39649 and pi1150 n42082_not ; n42085
g39650 and n42084_not n42085 ; n42086
g39651 and n41815_not n42010 ; n42087
g39652 nor pi1151 n41878 ; n42088
g39653 and pi1152 n42088_not ; n42089
g39654 and n41887_not n42089 ; n42090
g39655 nor pi1150 n42090 ; n42091
g39656 and n42087_not n42091 ; n42092
g39657 and pi1149 n42086_not ; n42093
g39658 and n42092_not n42093 ; n42094
g39659 nor pi1148 n42079 ; n42095
g39660 and n42094_not n42095 ; n42096
g39661 and n41755 n41768_not ; n42097
g39662 and n40673 n42097_not ; n42098
g39663 and pi1152 n41857_not ; n42099
g39664 and n41882_not n42099 ; n42100
g39665 nor pi1150 n42098 ; n42101
g39666 and n42100_not n42101 ; n42102
g39667 and pi1151 n41902 ; n42103
g39668 nor pi1152 n41898 ; n42104
g39669 and n42103_not n42104 ; n42105
g39670 and n40666 n41847 ; n42106
g39671 and n41985 n42106_not ; n42107
g39672 and pi1150 n42105_not ; n42108
g39673 and n42107_not n42108 ; n42109
g39674 and pi1149 n42109_not ; n42110
g39675 and n42102_not n42110 ; n42111
g39676 and pi1151 n41922 ; n42112
g39677 nor pi1152 n41930 ; n42113
g39678 and n42112_not n42113 ; n42114
g39679 and pi1152 n41840_not ; n42115
g39680 and n41920_not n42115 ; n42116
g39681 nor pi1150 n42116 ; n42117
g39682 and n42114_not n42117 ; n42118
g39683 and n41793_not n42043 ; n42119
g39684 and pi1151 n41957 ; n42120
g39685 nor pi1152 n41948 ; n42121
g39686 and n42120_not n42121 ; n42122
g39687 and pi1150 n42119_not ; n42123
g39688 and n42122_not n42123 ; n42124
g39689 nor pi1149 n42118 ; n42125
g39690 and n42124_not n42125 ; n42126
g39691 and pi1148 n42111_not ; n42127
g39692 and n42126_not n42127 ; n42128
g39693 and pi0213 n42096_not ; n42129
g39694 and n42128_not n42129 ; n42130
g39695 nor pi0209 n42065 ; n42131
g39696 and n42130_not n42131 ; n42132
g39697 nor n42064 n42132 ; n42133
g39698 and pi0230 n42133_not ; n42134
g39699 nor pi0230 pi0248 ; n42135
g39700 nor n42134 n42135 ; po0405
g39701 and pi0213_not n41990 ; n42137
g39702 and pi0057 n38886_not ; n42138
g39703 and n6305_not n38886 ; n42139
g39704 and n39738_not n39882 ; n42140
g39705 and pi0299 n38883 ; n42141
g39706 nor n40682 n42141 ; n42142
g39707 nor pi0214 n42142 ; n42143
g39708 and pi0212 n42140_not ; n42144
g39709 and n42143_not n42144 ; n42145
g39710 and pi0214 n42142_not ; n42146
g39711 nor pi0212 n39748 ; n42147
g39712 and n42146_not n42147 ; n42148
g39713 nor pi0219 n42145 ; n42149
g39714 and n42148_not n42149 ; n42150
g39715 and n6305 n39768_not ; n42151
g39716 and n42150_not n42151 ; n42152
g39717 and pi0057_not pi1151 ; n42153
g39718 and n42139_not n42153 ; n42154
g39719 and n42152_not n42154 ; n42155
g39720 nor n40183 n42141 ; n42156
g39721 and n39748_not n42156 ; n42157
g39722 nor pi0212 n42157 ; n42158
g39723 and pi0214_not n42156 ; n42159
g39724 nor n39854 n40182 ; n42160
g39725 and pi0214 n40635_not ; n42161
g39726 and n42160_not n42161 ; n42162
g39727 and pi0212 n42162_not ; n42163
g39728 and n42159_not n42163 ; n42164
g39729 nor n42158 n42164 ; n42165
g39730 nor pi0219 n42165 ; n42166
g39731 and n6305 n40652_not ; n42167
g39732 and n42166_not n42167 ; n42168
g39733 nor pi0057 pi1151 ; n42169
g39734 and n42139_not n42169 ; n42170
g39735 and n42168_not n42170 ; n42171
g39736 nor n42138 n42155 ; n42172
g39737 and n42171_not n42172 ; n42173
g39738 nor pi1152 n42173 ; n42174
g39739 and pi0299 n38883_not ; n42175
g39740 and n10843_not n42175 ; n42176
g39741 nor n38917 n42176 ; n42177
g39742 and n40083 n42177_not ; n42178
g39743 and n40660 n42178_not ; n42179
g39744 nor n40195 n40291 ; n42180
g39745 and pi1151 n42180_not ; n42181
g39746 and n42179_not n42181 ; n42182
g39747 and n40525 n42141_not ; n42183
g39748 nor n39686 n42141 ; n42184
g39749 nor pi0214 n42184 ; n42185
g39750 and n40149 n40628_not ; n42186
g39751 and pi0212 n42185_not ; n42187
g39752 and n42186_not n42187 ; n42188
g39753 and n41516 n42183_not ; n42189
g39754 and n42188_not n42189 ; n42190
g39755 nor pi1151 n42190 ; n42191
g39756 and n40164 n42191 ; n42192
g39757 and n38922 n42182_not ; n42193
g39758 and n42192_not n42193 ; n42194
g39759 and pi1150 n42194_not ; n42195
g39760 and n42174_not n42195 ; n42196
g39761 and pi0212_not n39736 ; n42197
g39762 and n40062 n42175_not ; n42198
g39763 and pi0212 n42198_not ; n42199
g39764 and n40739_not n42199 ; n42200
g39765 nor pi0219 n42197 ; n42201
g39766 and n42183_not n42201 ; n42202
g39767 and n42200_not n42202 ; n42203
g39768 and n39694 n40309_not ; n42204
g39769 and n42203_not n42204 ; n42205
g39770 and pi1151_not n41830 ; n42206
g39771 nor n39738 n42176 ; n42207
g39772 and n38885 n39635 ; n42208
g39773 and n42207_not n42208 ; n42209
g39774 and n38922 n42209_not ; n42210
g39775 and n42206_not n42210 ; n42211
g39776 and n42205_not n42211 ; n42212
g39777 and n10843 n40713 ; n42213
g39778 and n39066 n40100_not ; n42214
g39779 and n38745_not n40110 ; n42215
g39780 and pi0211 n40712 ; n42216
g39781 and n38608 n42215_not ; n42217
g39782 and n42216_not n42217 ; n42218
g39783 nor n42213 n42214 ; n42219
g39784 and n42218_not n42219 ; n42220
g39785 nor pi0219 n42220 ; n42221
g39786 and pi1151 n40123 ; n42222
g39787 and n42221_not n42222 ; n42223
g39788 and n38888 n42209_not ; n42224
g39789 and n42223_not n42224 ; n42225
g39790 nor pi1150 n42212 ; n42226
g39791 and n42225_not n42226 ; n42227
g39792 nor n42196 n42227 ; n42228
g39793 and pi0213 n42228_not ; n42229
g39794 nor pi0209 n42229 ; n42230
g39795 and n42137_not n42230 ; n42231
g39796 and pi0213 n39071 ; n42232
g39797 nor n10484 n39029 ; n42233
g39798 and n38675 n39253_not ; n42234
g39799 and pi0207 n38769_not ; n42235
g39800 and n39027_not n42235 ; n42236
g39801 and pi0207_not n39252 ; n42237
g39802 and pi0208 n42236_not ; n42238
g39803 and n42237_not n42238 ; n42239
g39804 nor n42234 n42239 ; n42240
g39805 and pi0211 n42240_not ; n42241
g39806 and pi0214 n42241 ; n42242
g39807 nor n42233 n42242 ; n42243
g39808 nor pi0212 n42243 ; n42244
g39809 nor pi0219 n42244 ; n42245
g39810 and pi0211_not n42240 ; n42246
g39811 nor n39099 n42246 ; n42247
g39812 and pi0214 n42247_not ; n42248
g39813 nor pi0211 n39029 ; n42249
g39814 nor pi0214 n42249 ; n42250
g39815 and n42241_not n42250 ; n42251
g39816 and pi0212 n42251_not ; n42252
g39817 and n42248_not n42252 ; n42253
g39818 and n42245 n42253_not ; n42254
g39819 and n39031 n42254_not ; n42255
g39820 and n41755 n42255_not ; n42256
g39821 and n39029_not n39073 ; n42257
g39822 nor n41978 n42257 ; n42258
g39823 nor n42256 n42258 ; n42259
g39824 nor n38966 n39909 ; n42260
g39825 and n38968_not n39909 ; n42261
g39826 nor po1038 n42260 ; n42262
g39827 and n42261_not n42262 ; n42263
g39828 and n41839 n42263_not ; n42264
g39829 and pi0214 n38953 ; n42265
g39830 and n39014 n42265_not ; n42266
g39831 nor pi0219 n42266 ; n42267
g39832 and pi0214 n38968_not ; n42268
g39833 and pi0214_not n38953 ; n42269
g39834 and pi0212 n42269_not ; n42270
g39835 and n42268_not n42270 ; n42271
g39836 and n42267 n42271_not ; n42272
g39837 nor po1038 n38971 ; n42273
g39838 and n42272_not n42273 ; n42274
g39839 and n40500 n42274_not ; n42275
g39840 and pi1152 n42264_not ; n42276
g39841 and n42275_not n42276 ; n42277
g39842 nor n42259 n42277 ; n42278
g39843 nor pi1150 n42278 ; n42279
g39844 and n38413_not n42247 ; n42280
g39845 and pi0219 n39074_not ; n42281
g39846 and n42280_not n42281 ; n42282
g39847 nor po1038 n42282 ; n42283
g39848 and pi0212 n42243_not ; n42284
g39849 nor pi0212 n39029 ; n42285
g39850 nor pi0219 n42285 ; n42286
g39851 and n42284_not n42286 ; n42287
g39852 and n42283 n42287_not ; n42288
g39853 and n40565 n42288_not ; n42289
g39854 and pi0214 n42240 ; n42290
g39855 and n42252 n42290_not ; n42291
g39856 and n42245 n42291_not ; n42292
g39857 and n42283 n42292_not ; n42293
g39858 and n41745 n42293_not ; n42294
g39859 nor pi1152 n42289 ; n42295
g39860 and n42294_not n42295 ; n42296
g39861 and pi0212 n38953_not ; n42297
g39862 and n42267 n42297_not ; n42298
g39863 and n38974 n42298_not ; n42299
g39864 and n40593 n42299_not ; n42300
g39865 nor n39013 n42268 ; n42301
g39866 nor pi0212 n42301 ; n42302
g39867 and pi0211_not n38966 ; n42303
g39868 nor n38992 n42303 ; n42304
g39869 and pi0214 n42304_not ; n42305
g39870 and pi0214_not n38968 ; n42306
g39871 and pi0212 n42305_not ; n42307
g39872 and n42306_not n42307 ; n42308
g39873 nor n42302 n42308 ; n42309
g39874 nor pi0219 n42309 ; n42310
g39875 and n38974 n42310_not ; n42311
g39876 and n41847 n42311_not ; n42312
g39877 and pi1152 n42300_not ; n42313
g39878 and n42312_not n42313 ; n42314
g39879 nor n42296 n42314 ; n42315
g39880 and pi1150 n42315_not ; n42316
g39881 nor n42279 n42316 ; n42317
g39882 nor pi0213 n42317 ; n42318
g39883 and pi0209 n42232_not ; n42319
g39884 and n42318_not n42319 ; n42320
g39885 nor n42231 n42320 ; n42321
g39886 and pi0230 n42321_not ; n42322
g39887 nor pi0230 pi0249 ; n42323
g39888 nor n42322 n42323 ; po0406
g39889 and n2531 n11513 ; n42325
g39890 nor n6286 n42325 ; n42326
g39891 nor pi0075 n42326 ; n42327
g39892 and n7333 n8966 ; n42328
g39893 nor n42327 n42328 ; n42329
g39894 nor pi0087 pi0250 ; n42330
g39895 and n8881 n42330 ; n42331
g39896 and n42329_not n42331 ; po0407
g39897 and pi0897 n10809 ; n42333
g39898 and pi0476_not n11444 ; n42334
g39899 nor n42333 n42334 ; n42335
g39900 and pi0200_not pi1053 ; n42336
g39901 and pi0200 pi1039 ; n42337
g39902 nor pi0199 n42336 ; n42338
g39903 and n42337_not n42338 ; n42339
g39904 nor n42335 n42339 ; n42340
g39905 and pi0251 n42335 ; n42341
g39906 or n42340 n42341 ; po0408
g39907 and n10983_not n11552 ; n42343
g39908 and n6198_not n11552 ; n42344
g39909 nor pi0979 pi0984 ; n42345
g39910 and pi1001 n42345 ; n42346
g39911 and n6186 n42346 ; n42347
g39912 and n6213_not n42347 ; n42348
g39913 and n6380 n42348 ; n42349
g39914 nor pi0252 n42349 ; n42350
g39915 and pi1092 pi1093_not ; n42351
g39916 and n42350_not n42351 ; n42352
g39917 and n6392 n42352_not ; n42353
g39918 and n6391 n42352 ; n42354
g39919 nor n42353 n42354 ; n42355
g39920 and n6198 n42355 ; n42356
g39921 nor n42344 n42356 ; n42357
g39922 and n6242 n42357_not ; n42358
g39923 and n6227_not n42355 ; n42359
g39924 and n6227 n11552 ; n42360
g39925 nor n42359 n42360 ; n42361
g39926 nor n6242 n42361 ; n42362
g39927 and pi0299 n42358_not ; n42363
g39928 and n42362_not n42363 ; n42364
g39929 and n6205 n42357_not ; n42365
g39930 nor n6205 n42361 ; n42366
g39931 nor pi0299 n42365 ; n42367
g39932 and n42366_not n42367 ; n42368
g39933 and n10983 n42364_not ; n42369
g39934 and n42368_not n42369 ; n42370
g39935 nor n7643 n42343 ; n42371
g39936 and n42370_not n42371 ; n42372
g39937 and pi0057 n11551 ; n42373
g39938 and n10982 n42347 ; n42374
g39939 and n21130 n42374 ; n42375
g39940 and n6217 n42375 ; n42376
g39941 and n38387_not n42376 ; n42377
g39942 and n6380 n42377 ; n42378
g39943 nor pi0252 n42378 ; n42379
g39944 and pi0057_not pi1092 ; n42380
g39945 and n42379_not n42380 ; n42381
g39946 and n7643 n42373_not ; n42382
g39947 and n42381_not n42382 ; n42383
g39948 nor n42372 n42383 ; po0409
g39949 nor n13061 n38508 ; n42385
g39950 and n38700_not n42385 ; n42386
g39951 and po1038_not n42386 ; n42387
g39952 and pi0219 n40080 ; n42388
g39953 nor n42387 n42388 ; n42389
g39954 and pi1153 n42389_not ; n42390
g39955 nor pi1151 n42390 ; n42391
g39956 and n10844 n38684 ; n42392
g39957 and pi0211 n38570_not ; n42393
g39958 nor n42392 n42393 ; n42394
g39959 nor n38545 n38562 ; n42395
g39960 and n38519 n42395_not ; n42396
g39961 nor po1038 n42396 ; n42397
g39962 and n42394 n42397 ; n42398
g39963 and n11446_not n39281 ; n42399
g39964 and pi1151 n42399_not ; n42400
g39965 and n42398_not n42400 ; n42401
g39966 nor n42391 n42401 ; n42402
g39967 nor pi1152 n42402 ; n42403
g39968 and n38519 n39783 ; n42404
g39969 nor pi1151 n11447 ; n42405
g39970 and n38688_not n42405 ; n42406
g39971 and n42404_not n42406 ; n42407
g39972 nor n11384 n38508 ; n42408
g39973 nor n38568 n39854 ; n42409
g39974 and pi1153 n42409_not ; n42410
g39975 and pi1151 n42408 ; n42411
g39976 and n42410_not n42411 ; n42412
g39977 nor po1038 n42412 ; n42413
g39978 and n42407_not n42413 ; n42414
g39979 and pi1151_not n10844 ; n42415
g39980 nor n39280 n42415 ; n42416
g39981 and po1038 n42416 ; n42417
g39982 and pi1152 n42417_not ; n42418
g39983 and n42414_not n42418 ; n42419
g39984 nor n42403 n42419 ; n42420
g39985 and pi0230 n42420_not ; n42421
g39986 nor pi0253 pi1091 ; n42422
g39987 and po1038 n42422_not ; n42423
g39988 and pi0211 pi1091 ; n42424
g39989 and pi1091 pi1153_not ; n42425
g39990 and pi0219 n42425 ; n42426
g39991 nor n42424 n42426 ; n42427
g39992 and n42423 n42427 ; n42428
g39993 and pi1091 n42394_not ; n42429
g39994 nor pi1153 n40915 ; n42430
g39995 and pi1153 n40952_not ; n42431
g39996 and n38519 n42431_not ; n42432
g39997 and n42430_not n42432 ; n42433
g39998 nor n42429 n42433 ; n42434
g39999 and pi0253 n42434_not ; n42435
g40000 nor n13064 n42410 ; n42436
g40001 and pi1091 n42436_not ; n42437
g40002 nor pi0253 n42437 ; n42438
g40003 nor po1038 n42438 ; n42439
g40004 and n42435_not n42439 ; n42440
g40005 and pi1151 n42428_not ; n42441
g40006 and n42440_not n42441 ; n42442
g40007 and pi0253 pi1091_not ; n42443
g40008 and pi0219 pi1091 ; n42444
g40009 and n38497_not n42444 ; n42445
g40010 and n42423 n42445_not ; n42446
g40011 and pi0219 n42446 ; n42447
g40012 and pi1091 pi1153 ; n42448
g40013 and n42387 n42448 ; n42449
g40014 nor pi1151 n42443 ; n42450
g40015 and n42449_not n42450 ; n42451
g40016 and n42447_not n42451 ; n42452
g40017 nor n42442 n42452 ; n42453
g40018 nor pi1152 n42453 ; n42454
g40019 and pi0211_not pi1091 ; n42455
g40020 and pi0219_not n42455 ; n42456
g40021 and n42446 n42456_not ; n42457
g40022 and n11446 n40911 ; n42458
g40023 and n38688_not n42458 ; n42459
g40024 nor pi1153 n40943 ; n42460
g40025 and n38561_not n40911 ; n42461
g40026 and pi1153 n42461_not ; n42462
g40027 and n38519 n42462_not ; n42463
g40028 and n42460_not n42463 ; n42464
g40029 and pi0253 n42459_not ; n42465
g40030 and n42464_not n42465 ; n42466
g40031 and pi1091 n39783 ; n42467
g40032 and pi1091 n38545 ; n42468
g40033 and n38958 n42468 ; n42469
g40034 and n38519 n42469_not ; n42470
g40035 and n42467_not n42470 ; n42471
g40036 and pi1091 n38688 ; n42472
g40037 and pi0211 n40965_not ; n42473
g40038 and n42472_not n42473 ; n42474
g40039 nor pi0253 n42471 ; n42475
g40040 and n42474_not n42475 ; n42476
g40041 nor n42466 n42476 ; n42477
g40042 nor n11446 n38519 ; n42478
g40043 and n42443_not n42478 ; n42479
g40044 and n42472_not n42479 ; n42480
g40045 and n39635 n42480_not ; n42481
g40046 and n42477_not n42481 ; n42482
g40047 and n42409 n42443_not ; n42483
g40048 nor n42425 n42483 ; n42484
g40049 and n42408 n42484_not ; n42485
g40050 nor po1038 n42422 ; n42486
g40051 and n42485_not n42486 ; n42487
g40052 nor n42446 n42487 ; n42488
g40053 and pi1151 n42488_not ; n42489
g40054 and pi1152 n42457_not ; n42490
g40055 and n42489_not n42490 ; n42491
g40056 and n42482_not n42491 ; n42492
g40057 nor n40910 n42492 ; n42493
g40058 and n42454_not n42493 ; n42494
g40059 and n40988 n41072 ; n42495
g40060 and pi1153 n42495_not ; n42496
g40061 nor pi1153 n41118 ; n42497
g40062 nor pi0219 n42497 ; n42498
g40063 and n42496_not n42498 ; n42499
g40064 nor pi1153 n41048 ; n42500
g40065 nor n40987 n41011 ; n42501
g40066 and pi0211_not n41044 ; n42502
g40067 and n42501 n42502_not ; n42503
g40068 and n41000 n41008_not ; n42504
g40069 and n42503 n42504 ; n42505
g40070 and pi1153 n42505_not ; n42506
g40071 and pi0219 n42500_not ; n42507
g40072 and n42506_not n42507 ; n42508
g40073 and pi0253 n42499_not ; n42509
g40074 and n42508_not n42509 ; n42510
g40075 and n40993_not n41048 ; n42511
g40076 and pi0211_not n42511 ; n42512
g40077 nor n41013 n42512 ; n42513
g40078 and pi1153 n42513_not ; n42514
g40079 nor n41039 n42514 ; n42515
g40080 and pi0219 n42515 ; n42516
g40081 and pi1153_not n41116 ; n42517
g40082 and pi1153 n41097 ; n42518
g40083 nor pi0219 n42517 ; n42519
g40084 and n42518_not n42519 ; n42520
g40085 nor pi0253 n42520 ; n42521
g40086 and n42516_not n42521 ; n42522
g40087 nor n42510 n42522 ; n42523
g40088 nor po1038 n42523 ; n42524
g40089 nor pi0219 n40980 ; n42525
g40090 nor pi0211 n40890 ; n42526
g40091 and n42525 n42526_not ; n42527
g40092 nor pi0219 n42527 ; n42528
g40093 and po1038 n42528 ; n42529
g40094 and n40874_not n42529 ; n42530
g40095 nor n40868 n42445 ; n42531
g40096 and n42525_not n42531 ; n42532
g40097 and pi0253 n42532_not ; n42533
g40098 nor pi0219 n40890 ; n42534
g40099 and pi0211 n40868 ; n42535
g40100 nor pi0211 n40874 ; n42536
g40101 and pi0219 n42535_not ; n42537
g40102 and n42536_not n42537 ; n42538
g40103 nor n42445 n42534 ; n42539
g40104 and n42538_not n42539 ; n42540
g40105 nor pi0253 n42540 ; n42541
g40106 and po1038 n42533_not ; n42542
g40107 and n42541_not n42542 ; n42543
g40108 and pi1151 n42530_not ; n42544
g40109 and n42543_not n42544 ; n42545
g40110 and n42524_not n42545 ; n42546
g40111 nor n41072 n42512 ; n42547
g40112 and n42525 n42547_not ; n42548
g40113 nor n40987 n40999 ; n42549
g40114 nor pi1153 n42549 ; n42550
g40115 nor n41102 n42550 ; n42551
g40116 and n42548 n42551_not ; n42552
g40117 and pi0219 n41009 ; n42553
g40118 and n41057_not n42506 ; n42554
g40119 and n42553 n42554_not ; n42555
g40120 nor n42552 n42555 ; n42556
g40121 and pi0253 n42556_not ; n42557
g40122 and n41012_not n42503 ; n42558
g40123 and n42550_not n42558 ; n42559
g40124 nor pi0219 n42559 ; n42560
g40125 and pi0219 n41011 ; n42561
g40126 nor n42560 n42561 ; n42562
g40127 and n42516_not n42562 ; n42563
g40128 nor pi0253 n42563 ; n42564
g40129 nor po1038 n42557 ; n42565
g40130 and n42564_not n42565 ; n42566
g40131 nor pi1151 n42566 ; n42567
g40132 nor n42546 n42567 ; n42568
g40133 and n42534 n42536_not ; n42569
g40134 and n42525 n42569_not ; n42570
g40135 and pi0219 n40874_not ; n42571
g40136 and po1038 n42571_not ; n42572
g40137 and n42570_not n42572 ; n42573
g40138 and n40874_not n42573 ; n42574
g40139 nor n42543 n42574 ; n42575
g40140 and n42568_not n42575 ; n42576
g40141 and pi1152 n42576_not ; n42577
g40142 and pi0219 n42515_not ; n42578
g40143 and n42520_not n42548 ; n42579
g40144 nor n42578 n42579 ; n42580
g40145 nor n40993 n42580 ; n42581
g40146 nor pi0253 n42581 ; n42582
g40147 and pi1153 n40988_not ; n42583
g40148 and n42503 n42525 ; n42584
g40149 and n42583_not n42584 ; n42585
g40150 nor pi1153 n41028 ; n42586
g40151 nor n41062 n42505 ; n42587
g40152 and pi1153 n42587 ; n42588
g40153 and pi0219 n42586_not ; n42589
g40154 and n42588_not n42589 ; n42590
g40155 nor n42585 n42590 ; n42591
g40156 and pi0253 n42591_not ; n42592
g40157 nor po1038 n42592 ; n42593
g40158 and n42582_not n42593 ; n42594
g40159 and n42545 n42594_not ; n42595
g40160 nor pi1091 n41039 ; n42596
g40161 nor pi1153 n42596 ; n42597
g40162 nor n41057 n42505 ; n42598
g40163 and pi0219_not n42549 ; n42599
g40164 nor n42597 n42599 ; n42600
g40165 and n42598 n42600 ; n42601
g40166 and pi0253 n42601_not ; n42602
g40167 and n41002_not n42578 ; n42603
g40168 nor pi1153 n41084 ; n42604
g40169 nor n40993 n42604 ; n42605
g40170 and pi0219_not n41118 ; n42606
g40171 and n42605 n42606 ; n42607
g40172 nor pi0253 n42607 ; n42608
g40173 and n42603_not n42608 ; n42609
g40174 nor po1038 n42602 ; n42610
g40175 and n42609_not n42610 ; n42611
g40176 nor pi1151 n42543 ; n42612
g40177 and n42611_not n42612 ; n42613
g40178 nor pi1152 n42613 ; n42614
g40179 and n42595_not n42614 ; n42615
g40180 nor n42577 n42615 ; n42616
g40181 and n40910 n42616_not ; n42617
g40182 nor pi0230 n42494 ; n42618
g40183 and n42617_not n42618 ; n42619
g40184 nor n42421 n42619 ; po0410
g40185 nor pi0219 n38882 ; n42621
g40186 nor n39145 n42621 ; n42622
g40187 and po1038 n42622 ; n42623
g40188 and pi1154 n38977 ; n42624
g40189 nor n39033 n42624 ; n42625
g40190 and n11446 n42625_not ; n42626
g40191 and pi0299 n38519 ; n42627
g40192 and n11446_not n38959 ; n42628
g40193 nor n42627 n42628 ; n42629
g40194 nor n38939 n42629 ; n42630
g40195 nor n42626 n42630 ; n42631
g40196 nor po1038 n42631 ; n42632
g40197 nor pi1152 n42623 ; n42633
g40198 and n42632_not n42633 ; n42634
g40199 and n11446 n38882_not ; n42635
g40200 and n40028 n42635_not ; n42636
g40201 and pi0200_not pi1154 ; n42637
g40202 and n11373 n42637_not ; n42638
g40203 and n38976 n39854_not ; n42639
g40204 nor n42638 n42639 ; n42640
g40205 nor pi0219 n42640 ; n42641
g40206 nor n38558 n38976 ; n42642
g40207 and n38488 n42642_not ; n42643
g40208 nor pi1154 n39022 ; n42644
g40209 nor n38941 n42644 ; n42645
g40210 and n42643_not n42645 ; n42646
g40211 and pi0219 n42646_not ; n42647
g40212 nor po1038 n42641 ; n42648
g40213 and n42647_not n42648 ; n42649
g40214 and pi1152 n42636_not ; n42650
g40215 and n42649_not n42650 ; n42651
g40216 nor n42634 n42651 ; n42652
g40217 and pi0230 n42652_not ; n42653
g40218 nor pi0254 pi1091 ; n42654
g40219 and pi1091 n42622_not ; n42655
g40220 and po1038 n42654_not ; n42656
g40221 and n42655_not n42656 ; n42657
g40222 and po1038 n42456 ; n42658
g40223 nor n42657 n42658 ; n42659
g40224 and pi1153 n40932_not ; n42660
g40225 nor pi1154 n42660 ; n42661
g40226 and pi0211_not n38683 ; n42662
g40227 and n42430_not n42661 ; n42663
g40228 and n42662_not n42663 ; n42664
g40229 and pi1091 n38488 ; n42665
g40230 and n38568_not n42665 ; n42666
g40231 and n39045_not n42666 ; n42667
g40232 nor n42664 n42667 ; n42668
g40233 nor pi0219 n42668 ; n42669
g40234 and pi1154 n42455 ; n42670
g40235 nor n42444 n42670 ; n42671
g40236 nor n42646 n42671 ; n42672
g40237 nor n42669 n42672 ; n42673
g40238 and pi0254 n42673_not ; n42674
g40239 and pi1154 n42409_not ; n42675
g40240 and pi0219 n39022_not ; n42676
g40241 and n42675_not n42676 ; n42677
g40242 nor n42641 n42677 ; n42678
g40243 nor pi0254 n42678 ; n42679
g40244 nor n42654 n42679 ; n42680
g40245 and n42674_not n42680 ; n42681
g40246 and po1038_not n42681 ; n42682
g40247 and pi1152 n42659 ; n42683
g40248 and n42682_not n42683 ; n42684
g40249 and n40918 n42425 ; n42685
g40250 nor n42467 n42685 ; n42686
g40251 and pi0211 n42661_not ; n42687
g40252 and n42686_not n42687 ; n42688
g40253 and n11445 n42448 ; n42689
g40254 nor pi1154 n42689 ; n42690
g40255 and pi1091 n38959 ; n42691
g40256 and pi1154 n42691_not ; n42692
g40257 nor pi0211 n42690 ; n42693
g40258 and n42692_not n42693 ; n42694
g40259 nor n42688 n42694 ; n42695
g40260 nor pi0219 n42695 ; n42696
g40261 and pi0211 n42692 ; n42697
g40262 and pi1091 n39666 ; n42698
g40263 and n38495 n42698_not ; n42699
g40264 and n42467_not n42699 ; n42700
g40265 and pi0219 n42690_not ; n42701
g40266 and n42700_not n42701 ; n42702
g40267 and n42697_not n42702 ; n42703
g40268 nor n42696 n42703 ; n42704
g40269 nor pi0254 n42704 ; n42705
g40270 nor pi1153 n40919 ; n42706
g40271 nor n42462 n42706 ; n42707
g40272 and pi1091 pi1154_not ; n42708
g40273 and n38533 n42708 ; n42709
g40274 nor n42707 n42709 ; n42710
g40275 and n11446 n42710_not ; n42711
g40276 and pi1091 n11446_not ; n42712
g40277 and n38938_not n42712 ; n42713
g40278 nor pi1154 n42713 ; n42714
g40279 and n40968 n42463 ; n42715
g40280 and pi1091 n38641_not ; n42716
g40281 nor n42707 n42716 ; n42717
g40282 and n42478 n42717_not ; n42718
g40283 and pi1154 n42715_not ; n42719
g40284 and n42718_not n42719 ; n42720
g40285 nor n42714 n42720 ; n42721
g40286 and pi0254 n42711_not ; n42722
g40287 and n42721_not n42722 ; n42723
g40288 nor n42705 n42723 ; n42724
g40289 nor po1038 n42724 ; n42725
g40290 nor pi1152 n42657 ; n42726
g40291 and n42725_not n42726 ; n42727
g40292 nor n40910 n42684 ; n42728
g40293 and n42727_not n42728 ; n42729
g40294 and pi1091 n39145 ; n42730
g40295 nor pi0211 n40866 ; n42731
g40296 and n42571 n42731_not ; n42732
g40297 and pi0219_not n40890 ; n42733
g40298 nor n42732 n42733 ; n42734
g40299 and n11446 n42425 ; n42735
g40300 and pi0254 n42735_not ; n42736
g40301 and n42730_not n42736 ; n42737
g40302 and n42734 n42737 ; n42738
g40303 and n42448_not n42569 ; n42739
g40304 nor pi0254 n42730 ; n42740
g40305 and n42538_not n42740 ; n42741
g40306 and n42739_not n42741 ; n42742
g40307 and pi0253 n42738_not ; n42743
g40308 and n42742_not n42743 ; n42744
g40309 and pi0253 po1038 ; n42745
g40310 and n42659 n42745_not ; n42746
g40311 nor n42744 n42746 ; n42747
g40312 nor pi0253 n42681 ; n42748
g40313 and pi1154 n40985_not ; n42749
g40314 and n42503 n42749 ; n42750
g40315 and n42496_not n42750 ; n42751
g40316 and pi1153_not n42559 ; n42752
g40317 nor n41118 n42752 ; n42753
g40318 nor pi1154 n42753 ; n42754
g40319 and pi0254 n42751_not ; n42755
g40320 and n42754_not n42755 ; n42756
g40321 and pi0211 n41044 ; n42757
g40322 nor n40993 n42757 ; n42758
g40323 nor pi1153 n42758 ; n42759
g40324 and n41012_not n41028 ; n42760
g40325 and pi1154 n42760 ; n42761
g40326 nor n41116 n42761 ; n42762
g40327 nor pi0254 n42759 ; n42763
g40328 and n42762_not n42763 ; n42764
g40329 nor n42756 n42764 ; n42765
g40330 nor pi0219 n42765 ; n42766
g40331 and pi1154 n42506_not ; n42767
g40332 and n42587_not n42767 ; n42768
g40333 and pi1153 n41048_not ; n42769
g40334 nor pi1154 n42586 ; n42770
g40335 and n42769_not n42770 ; n42771
g40336 and pi0254 n42771_not ; n42772
g40337 and n42768_not n42772 ; n42773
g40338 and n42500_not n42760 ; n42774
g40339 and n38495 n42774_not ; n42775
g40340 and n40990_not n42775 ; n42776
g40341 nor pi1153 n41032 ; n42777
g40342 and n41041 n42777_not ; n42778
g40343 nor pi1154 n42778 ; n42779
g40344 and n40993_not n41039 ; n42780
g40345 and n42779 n42780_not ; n42781
g40346 and pi1153 n41013 ; n42782
g40347 and n38488 n40995_not ; n42783
g40348 and n42782_not n42783 ; n42784
g40349 nor pi0254 n42784 ; n42785
g40350 and n42776_not n42785 ; n42786
g40351 and n42781_not n42786 ; n42787
g40352 nor n42773 n42787 ; n42788
g40353 and pi0219 n42788_not ; n42789
g40354 and pi0253 n42789_not ; n42790
g40355 and n42766_not n42790 ; n42791
g40356 nor po1038 n42748 ; n42792
g40357 and n42791_not n42792 ; n42793
g40358 and pi1152 n42747_not ; n42794
g40359 and n42793_not n42794 ; n42795
g40360 nor n42657 n42745 ; n42796
g40361 and n42570_not n42738 ; n42797
g40362 and n42528_not n42742 ; n42798
g40363 and pi0253 n42797_not ; n42799
g40364 and n42798_not n42799 ; n42800
g40365 nor n42796 n42800 ; n42801
g40366 and pi0253_not n42724 ; n42802
g40367 and n38495 n41057_not ; n42803
g40368 and pi1153_not n41000 ; n42804
g40369 nor pi1154 n41003 ; n42805
g40370 nor pi1154 n42805 ; n42806
g40371 nor n42504 n42804 ; n42807
g40372 and n42806_not n42807 ; n42808
g40373 and pi0219 n42803_not ; n42809
g40374 and n42808_not n42809 ; n42810
g40375 and pi1154 n40999 ; n42811
g40376 and n42547 n42804_not ; n42812
g40377 nor pi0219 n42811 ; n42813
g40378 and n42812_not n42813 ; n42814
g40379 nor n42810 n42814 ; n42815
g40380 and pi0254 n42815_not ; n42816
g40381 and n41014 n42500_not ; n42817
g40382 and n38488 n42817_not ; n42818
g40383 and pi0219 n42775_not ; n42819
g40384 and n42779_not n42819 ; n42820
g40385 and n42818_not n42820 ; n42821
g40386 and pi1154 n41011 ; n42822
g40387 nor n41044 n42822 ; n42823
g40388 nor pi0211 n42823 ; n42824
g40389 and n40985_not n41116 ; n42825
g40390 and n42604_not n42825 ; n42826
g40391 nor pi1154 n42826 ; n42827
g40392 and n40993_not n41118 ; n42828
g40393 and pi1154 n42828_not ; n42829
g40394 and n42826_not n42829 ; n42830
g40395 nor pi0219 n42824 ; n42831
g40396 and n42827_not n42831 ; n42832
g40397 and n42830_not n42832 ; n42833
g40398 nor pi0254 n42833 ; n42834
g40399 and n42821_not n42834 ; n42835
g40400 nor n42816 n42835 ; n42836
g40401 and pi0253 n42836_not ; n42837
g40402 nor po1038 n42802 ; n42838
g40403 and n42837_not n42838 ; n42839
g40404 nor pi1152 n42801 ; n42840
g40405 and n42839_not n42840 ; n42841
g40406 and n40910 n42841_not ; n42842
g40407 and n42795_not n42842 ; n42843
g40408 nor pi0230 n42729 ; n42844
g40409 and n42843_not n42844 ; n42845
g40410 nor n42653 n42845 ; po0411
g40411 and pi0200_not pi1049 ; n42847
g40412 and pi0200 pi1036 ; n42848
g40413 nor n42847 n42848 ; n42849
g40414 and n42335_not n42849 ; n42850
g40415 and pi0255_not n42335 ; n42851
g40416 nor n42850 n42851 ; po0412
g40417 and pi0200_not pi1048 ; n42853
g40418 and pi0200 pi1070 ; n42854
g40419 nor n42853 n42854 ; n42855
g40420 and n42335_not n42855 ; n42856
g40421 and pi0256_not n42335 ; n42857
g40422 nor n42856 n42857 ; po0413
g40423 and pi0200_not pi1084 ; n42859
g40424 and pi0200 pi1065 ; n42860
g40425 nor n42859 n42860 ; n42861
g40426 and n42335_not n42861 ; n42862
g40427 and pi0257_not n42335 ; n42863
g40428 nor n42862 n42863 ; po0414
g40429 and pi0200_not pi1072 ; n42865
g40430 and pi0200 pi1062 ; n42866
g40431 nor n42865 n42866 ; n42867
g40432 and n42335_not n42867 ; n42868
g40433 and pi0258_not n42335 ; n42869
g40434 nor n42868 n42869 ; po0415
g40435 and pi0200_not pi1059 ; n42871
g40436 and pi0200 pi1069 ; n42872
g40437 nor n42871 n42872 ; n42873
g40438 and n42335_not n42873 ; n42874
g40439 and pi0259_not n42335 ; n42875
g40440 nor n42874 n42875 ; po0416
g40441 and pi0200_not pi1044 ; n42877
g40442 and pi0200 pi1067 ; n42878
g40443 nor pi0199 n42877 ; n42879
g40444 and n42878_not n42879 ; n42880
g40445 nor n42335 n42880 ; n42881
g40446 and pi0260 n42335 ; n42882
g40447 or n42881 n42882 ; po0417
g40448 and pi0200_not pi1037 ; n42884
g40449 and pi0200 pi1040 ; n42885
g40450 nor pi0199 n42884 ; n42886
g40451 and n42885_not n42886 ; n42887
g40452 nor n42335 n42887 ; n42888
g40453 and pi0261 n42335 ; n42889
g40454 or n42888 n42889 ; po0418
g40455 and pi1093 pi1142 ; n42891
g40456 nor pi0262 pi1093 ; n42892
g40457 nor n42891 n42892 ; n42893
g40458 nor pi0228 n42893 ; n42894
g40459 nor pi0123 pi1142 ; n42895
g40460 and pi0123 pi0262 ; n42896
g40461 and pi0228 n42895_not ; n42897
g40462 and n42896_not n42897 ; n42898
g40463 nor n42894 n42898 ; n42899
g40464 nor pi0228 pi1093 ; n42900
g40465 and pi0123 pi0228 ; n42901
g40466 nor n42900 n42901 ; n42902
g40467 nor pi0262 n42902 ; n42903
g40468 nor n40700 n42903 ; n42904
g40469 and pi0199 n42902 ; n42905
g40470 and n38441 n42905_not ; n42906
g40471 and n42904 n42906_not ; n42907
g40472 nor n42899 n42907 ; n42908
g40473 and pi0207_not n42903 ; n42909
g40474 nor pi0208 n42909 ; n42910
g40475 nor n40700 n42910 ; n42911
g40476 nor n42908 n42911 ; n42912
g40477 and n39711_not n42902 ; n42913
g40478 nor pi0299 n42913 ; n42914
g40479 and n42899_not n42914 ; n42915
g40480 and pi0299 n42904_not ; n42916
g40481 and pi0208 n42915_not ; n42917
g40482 and n42916_not n42917 ; n42918
g40483 nor po1038 n42918 ; n42919
g40484 and n42912_not n42919 ; n42920
g40485 and n39864_not n42902 ; n42921
g40486 and po1038 n42899_not ; n42922
g40487 and n42921_not n42922 ; n42923
g40488 or n42920 n42923 ; po0419
g40489 nor n40915 n42708 ; n42925
g40490 nor pi1156 n38577 ; n42926
g40491 and n42925_not n42926 ; n42927
g40492 and pi1155 n38985_not ; n42928
g40493 and n40952 n42928_not ; n42929
g40494 and pi1154_not n42716 ; n42930
g40495 nor n42929 n42930 ; n42931
g40496 and n40965_not n42931 ; n42932
g40497 and n38479 n42932_not ; n42933
g40498 nor pi1154 n38702 ; n42934
g40499 and n38545 n38576_not ; n42935
g40500 and pi1154 n42935_not ; n42936
g40501 and pi1091 n38483 ; n42937
g40502 and n42936_not n42937 ; n42938
g40503 and n42934_not n42938 ; n42939
g40504 and pi0219 n42927_not ; n42940
g40505 and n42939_not n42940 ; n42941
g40506 and n42933_not n42941 ; n42942
g40507 nor pi0211 n42931 ; n42943
g40508 and n38568 n39111_not ; n42944
g40509 and n42424 n42944_not ; n42945
g40510 and n38766_not n42945 ; n42946
g40511 nor n42943 n42946 ; n42947
g40512 and pi1156 n42947_not ; n42948
g40513 nor n38766 n42925 ; n42949
g40514 and pi0211 n42949 ; n42950
g40515 nor n38577 n39000 ; n42951
g40516 and n42455 n42951 ; n42952
g40517 nor n42950 n42952 ; n42953
g40518 nor pi1156 n42953 ; n42954
g40519 nor pi0219 n42954 ; n42955
g40520 and n42948_not n42955 ; n42956
g40521 nor n42942 n42956 ; n42957
g40522 nor pi0263 n42957 ; n42958
g40523 and pi1154_not n38646 ; n42959
g40524 and pi1154 n38591_not ; n42960
g40525 and pi1156 n42960_not ; n42961
g40526 nor pi0299 n42961 ; n42962
g40527 nor n39854 n42959 ; n42963
g40528 and n42962_not n42963 ; n42964
g40529 and pi1156 n42964_not ; n42965
g40530 and n42951_not n42962 ; n42966
g40531 and pi0219 n42966_not ; n42967
g40532 and n42965_not n42967 ; n42968
g40533 and n38648_not n39499 ; n42969
g40534 nor n39000 n42969 ; n42970
g40535 nor pi0211 n42970 ; n42971
g40536 and pi1156_not n42949 ; n42972
g40537 nor n38568 n38595 ; n42973
g40538 and pi1154 n42973_not ; n42974
g40539 and n38544_not n42934 ; n42975
g40540 and pi1156 n42974_not ; n42976
g40541 and n42975_not n42976 ; n42977
g40542 and pi0211 n42972_not ; n42978
g40543 and n42977_not n42978 ; n42979
g40544 nor pi0219 n42971 ; n42980
g40545 and n42979_not n42980 ; n42981
g40546 and pi0263 pi1091 ; n42982
g40547 and n42968_not n42982 ; n42983
g40548 and n42981_not n42983 ; n42984
g40549 nor n42958 n42984 ; n42985
g40550 and po1038_not n42985 ; n42986
g40551 and pi0219 n38483_not ; n42987
g40552 nor pi0219 n38484 ; n42988
g40553 and n38495_not n42988 ; n42989
g40554 nor n42987 n42989 ; n42990
g40555 and pi1091 n42990_not ; n42991
g40556 and pi0263 pi1091_not ; n42992
g40557 nor n42991 n42992 ; n42993
g40558 and po1038 n42993_not ; n42994
g40559 nor n40910 n42994 ; n42995
g40560 and n42986_not n42995 ; n42996
g40561 and pi1091 n42987 ; n42997
g40562 and pi0211 n40874 ; n42998
g40563 nor pi0211 n42708 ; n42999
g40564 nor n38484 n42999 ; n43000
g40565 and n42998_not n43000 ; n43001
g40566 nor n40890 n43001 ; n43002
g40567 nor pi0219 n43002 ; n43003
g40568 nor pi0263 n42732 ; n43004
g40569 and n43003_not n43004 ; n43005
g40570 nor n38484 n42670 ; n43006
g40571 nor n42998 n43006 ; n43007
g40572 and n42534 n43007_not ; n43008
g40573 and pi0263 n42538_not ; n43009
g40574 and n43008_not n43009 ; n43010
g40575 nor n43005 n43010 ; n43011
g40576 and n40860 n42997_not ; n43012
g40577 and n43011_not n43012 ; n43013
g40578 and n40860_not n42993 ; n43014
g40579 and po1038 n43014_not ; n43015
g40580 and n43013_not n43015 ; n43016
g40581 nor n40860 n42985 ; n43017
g40582 and pi1155 n41118_not ; n43018
g40583 and pi1154 n43018_not ; n43019
g40584 and n41105 n43019 ; n43020
g40585 and pi1155_not n42596 ; n43021
g40586 and pi1155 n41009_not ; n43022
g40587 nor pi1154 n43022 ; n43023
g40588 and n43021_not n43023 ; n43024
g40589 and n41116_not n43021 ; n43025
g40590 and pi1155 n41072_not ; n43026
g40591 nor pi1154 n43026 ; n43027
g40592 and n43025_not n43027 ; n43028
g40593 nor pi1156 n43028 ; n43029
g40594 nor n43020 n43024 ; n43030
g40595 and n43029 n43030 ; n43031
g40596 and pi1155_not n41000 ; n43032
g40597 and n41044_not n41102 ; n43033
g40598 nor n43032 n43033 ; n43034
g40599 nor pi1154 n43034 ; n43035
g40600 and pi1156 n43035_not ; n43036
g40601 and n41000 n43023 ; n43037
g40602 and n40983_not n43020 ; n43038
g40603 nor n43037 n43038 ; n43039
g40604 and n43036 n43039 ; n43040
g40605 nor pi0211 n43031 ; n43041
g40606 and n43040_not n43041 ; n43042
g40607 and n40988 n43019 ; n43043
g40608 and n43036 n43043_not ; n43044
g40609 and n42501 n43019 ; n43045
g40610 and n43029 n43045_not ; n43046
g40611 and pi0211 n43044_not ; n43047
g40612 and n43046_not n43047 ; n43048
g40613 nor pi0219 n43042 ; n43049
g40614 and n43048_not n43049 ; n43050
g40615 and pi1155 n41008 ; n43051
g40616 and pi1154 n41028 ; n43052
g40617 and n43051_not n43052 ; n43053
g40618 and n40985_not n43053 ; n43054
g40619 nor n43037 n43054 ; n43055
g40620 and n38479 n43055_not ; n43056
g40621 nor n43024 n43053 ; n43057
g40622 nor pi1156 n43057 ; n43058
g40623 and pi1154_not n41039 ; n43059
g40624 nor n41062 n43059 ; n43060
g40625 and n38483 n43051_not ; n43061
g40626 and n43060_not n43061 ; n43062
g40627 and pi0219 n43062_not ; n43063
g40628 and n43056_not n43063 ; n43064
g40629 and n43058_not n43064 ; n43065
g40630 nor pi0263 n43065 ; n43066
g40631 and n43050_not n43066 ; n43067
g40632 nor n41040 n41055 ; n43068
g40633 and pi1154 n43068_not ; n43069
g40634 and pi1155 n42760_not ; n43070
g40635 nor pi1155 n42511 ; n43071
g40636 nor pi1154 n43070 ; n43072
g40637 and n43071_not n43072 ; n43073
g40638 and n38483 n43069_not ; n43074
g40639 and n43073_not n43074 ; n43075
g40640 nor n41014 n42822 ; n43076
g40641 nor n43068 n43076 ; n43077
g40642 and n38479 n43077_not ; n43078
g40643 and n41026_not n43077 ; n43079
g40644 nor pi1156 n43079 ; n43080
g40645 and pi0219 n43075_not ; n43081
g40646 and n43078_not n43081 ; n43082
g40647 and n43080_not n43082 ; n43083
g40648 and pi1154 n41098_not ; n43084
g40649 and n41046_not n43084 ; n43085
g40650 nor pi1154 n41085 ; n43086
g40651 and pi1155 n42825 ; n43087
g40652 and n43086 n43087_not ; n43088
g40653 and n41114_not n43084 ; n43089
g40654 nor pi1156 n42811 ; n43090
g40655 and n43089_not n43090 ; n43091
g40656 nor pi1156 n43091 ; n43092
g40657 nor n43088 n43092 ; n43093
g40658 and pi1156 n42828 ; n43094
g40659 nor n43093 n43094 ; n43095
g40660 nor n43085 n43095 ; n43096
g40661 and pi0211 n43096_not ; n43097
g40662 and n41026_not n41091 ; n43098
g40663 and pi1155 n43098 ; n43099
g40664 and n43086 n43099_not ; n43100
g40665 and n42828_not n43100 ; n43101
g40666 and pi1156 n43101_not ; n43102
g40667 and n43089_not n43102 ; n43103
g40668 and n43091 n43100_not ; n43104
g40669 nor pi0211 n43103 ; n43105
g40670 and n43104_not n43105 ; n43106
g40671 nor pi0219 n43106 ; n43107
g40672 and n43097_not n43107 ; n43108
g40673 and pi0263 n43083_not ; n43109
g40674 and n43108_not n43109 ; n43110
g40675 and n40860 n43067_not ; n43111
g40676 and n43110_not n43111 ; n43112
g40677 nor po1038 n43017 ; n43113
g40678 and n43112_not n43113 ; n43114
g40679 and n40910 n43016_not ; n43115
g40680 and n43114_not n43115 ; n43116
g40681 nor pi0230 n42996 ; n43117
g40682 and n43116_not n43117 ; n43118
g40683 and po1038 n42990 ; n43119
g40684 and n38578_not n38649 ; n43120
g40685 nor pi1156 n43120 ; n43121
g40686 and n38592 n39112_not ; n43122
g40687 and n43121_not n43122 ; n43123
g40688 and pi1156 n39854 ; n43124
g40689 and pi0219 n43124_not ; n43125
g40690 and n43123_not n43125 ; n43126
g40691 nor n38510 n43123 ; n43127
g40692 and pi0211 n43127_not ; n43128
g40693 and n42980 n43128_not ; n43129
g40694 nor po1038 n43126 ; n43130
g40695 and n43129_not n43130 ; n43131
g40696 and pi0230 n43119_not ; n43132
g40697 and n43131_not n43132 ; n43133
g40698 nor n43118 n43133 ; po0420
g40699 and pi1091 pi1143 ; n43135
g40700 and pi0200_not n43135 ; n43136
g40701 and pi0796_not n40863 ; n43137
g40702 and pi0264 n40863_not ; n43138
g40703 nor pi1091 n43137 ; n43139
g40704 and n43138_not n43139 ; n43140
g40705 and pi0199 n43136_not ; n43141
g40706 and n43140_not n43141 ; n43142
g40707 and pi1091 pi1141 ; n43143
g40708 and pi0796_not n40885 ; n43144
g40709 and pi0264 n40885_not ; n43145
g40710 nor pi1091 n43144 ; n43146
g40711 and n43145_not n43146 ; n43147
g40712 nor n43143 n43147 ; n43148
g40713 nor pi0200 n43148 ; n43149
g40714 and pi1091 pi1142 ; n43150
g40715 nor n43147 n43150 ; n43151
g40716 and pi0200 n43151_not ; n43152
g40717 nor pi0199 n43149 ; n43153
g40718 and n43152_not n43153 ; n43154
g40719 and n16479 n43142_not ; n43155
g40720 and n43154_not n43155 ; n43156
g40721 and pi0219 n42455_not ; n43157
g40722 nor n39410 n43157 ; n43158
g40723 nor n43140 n43158 ; n43159
g40724 nor pi0211 n43148 ; n43160
g40725 and pi0211 n43151_not ; n43161
g40726 nor pi0219 n43160 ; n43162
g40727 and n43161_not n43162 ; n43163
g40728 nor n16479 n43159 ; n43164
g40729 and n43163_not n43164 ; n43165
g40730 nor n43156 n43165 ; n43166
g40731 nor pi0230 n43166 ; n43167
g40732 and pi0211_not pi1141 ; n43168
g40733 nor pi0219 n38455 ; n43169
g40734 and n43168_not n43169 ; n43170
g40735 nor n39410 n43170 ; n43171
g40736 nor n16479 n43171 ; n43172
g40737 and pi0199_not pi1141 ; n43173
g40738 and n39388 n43173_not ; n43174
g40739 nor n38444 n43174 ; n43175
g40740 and n16479 n43175_not ; n43176
g40741 and pi0230 n43172_not ; n43177
g40742 and n43176_not n43177 ; n43178
g40743 or n43167 n43178 ; po0421
g40744 and pi1091 pi1144 ; n43180
g40745 and pi0200_not n43180 ; n43181
g40746 and pi0819_not n40863 ; n43182
g40747 and pi0265 n40863_not ; n43183
g40748 nor pi1091 n43182 ; n43184
g40749 and n43183_not n43184 ; n43185
g40750 and pi0199 n43181_not ; n43186
g40751 and n43185_not n43186 ; n43187
g40752 and pi0819_not n40885 ; n43188
g40753 and pi0265 n40885_not ; n43189
g40754 nor pi1091 n43188 ; n43190
g40755 and n43189_not n43190 ; n43191
g40756 nor n43150 n43191 ; n43192
g40757 nor pi0200 n43192 ; n43193
g40758 nor n43135 n43191 ; n43194
g40759 and pi0200 n43194_not ; n43195
g40760 nor pi0199 n43193 ; n43196
g40761 and n43195_not n43196 ; n43197
g40762 and n16479 n43187_not ; n43198
g40763 and n43197_not n43198 ; n43199
g40764 nor n40771 n43157 ; n43200
g40765 nor n43185 n43200 ; n43201
g40766 nor pi0211 n43192 ; n43202
g40767 and pi0211 n43194_not ; n43203
g40768 nor pi0219 n43202 ; n43204
g40769 and n43203_not n43204 ; n43205
g40770 nor n16479 n43201 ; n43206
g40771 and n43205_not n43206 ; n43207
g40772 nor n43199 n43207 ; n43208
g40773 nor pi0230 n43208 ; n43209
g40774 and pi0211_not pi1142 ; n43210
g40775 nor pi0219 n38418 ; n43211
g40776 and n43210_not n43211 ; n43212
g40777 nor n40771 n43212 ; n43213
g40778 nor n16479 n43213 ; n43214
g40779 and n38443_not n40782 ; n43215
g40780 nor n38437 n43215 ; n43216
g40781 and n16479 n43216_not ; n43217
g40782 and pi0230 n43214_not ; n43218
g40783 and n43217_not n43218 ; n43219
g40784 or n43209 n43219 ; po0422
g40785 and pi0211_not pi1136 ; n43221
g40786 and pi0219 n43221_not ; n43222
g40787 and pi0211 pi1135_not ; n43223
g40788 nor n43222 n43223 ; n43224
g40789 and n10844_not n43224 ; n43225
g40790 and po1038 n43225 ; n43226
g40791 and pi0299 n43225 ; n43227
g40792 and pi0199_not pi1135 ; n43228
g40793 and pi0200 n43228_not ; n43229
g40794 and pi0199 pi1136 ; n43230
g40795 nor pi0200 n43230 ; n43231
g40796 nor pi0299 n43229 ; n43232
g40797 and n43231_not n43232 ; n43233
g40798 nor n43227 n43233 ; n43234
g40799 nor po1038 n43234 ; n43235
g40800 and pi0230 n43226_not ; n43236
g40801 and n43235_not n43236 ; n43237
g40802 nor n43157 n43222 ; n43238
g40803 nor pi0266 n40863 ; n43239
g40804 and pi0948_not n40863 ; n43240
g40805 nor pi1091 n43239 ; n43241
g40806 and n43240_not n43241 ; n43242
g40807 nor n43238 n43242 ; n43243
g40808 nor n16479 n43243 ; n43244
g40809 nor pi0266 n40885 ; n43245
g40810 and pi0948_not n40885 ; n43246
g40811 nor pi1091 n43245 ; n43247
g40812 and n43246_not n43247 ; n43248
g40813 nor pi0219 n43248 ; n43249
g40814 and pi1135 n42424 ; n43250
g40815 and n43249 n43250_not ; n43251
g40816 and n43244 n43251_not ; n43252
g40817 nor pi0199 n43248 ; n43253
g40818 and pi1091 pi1136 ; n43254
g40819 and pi0199 n43242_not ; n43255
g40820 and n43254_not n43255 ; n43256
g40821 nor n43253 n43256 ; n43257
g40822 and pi0200_not n43257 ; n43258
g40823 and pi1091 pi1135 ; n43259
g40824 and n43253 n43259_not ; n43260
g40825 and pi0200 n43255_not ; n43261
g40826 and n43260_not n43261 ; n43262
g40827 nor n43258 n43262 ; n43263
g40828 and n16479 n43263_not ; n43264
g40829 nor pi0230 n43252 ; n43265
g40830 and n43264_not n43265 ; n43266
g40831 nor n43237 n43266 ; n43267
g40832 nor pi1134 n43267 ; n43268
g40833 and n38699 n43230_not ; n43269
g40834 nor n43229 n43269 ; n43270
g40835 and n16479 n43270 ; n43271
g40836 and n16479_not n43224 ; n43272
g40837 and pi0230 n43271_not ; n43273
g40838 and n43272_not n43273 ; n43274
g40839 and pi1091 n43223_not ; n43275
g40840 and n43249 n43275_not ; n43276
g40841 and n43244 n43276_not ; n43277
g40842 and pi0199_not pi1091 ; n43278
g40843 nor n43257 n43278 ; n43279
g40844 nor pi0200 n43279 ; n43280
g40845 nor n43262 n43280 ; n43281
g40846 and n16479 n43281_not ; n43282
g40847 nor pi0230 n43277 ; n43283
g40848 and n43282_not n43283 ; n43284
g40849 nor n43274 n43284 ; n43285
g40850 and pi1134 n43285_not ; n43286
g40851 nor n43268 n43286 ; po0423
g40852 and pi1155 n42431_not ; n43288
g40853 and n42706_not n43288 ; n43289
g40854 nor pi1155 n39027 ; n43290
g40855 and pi1091 n43290 ; n43291
g40856 nor n43289 n43291 ; n43292
g40857 nor pi1154 n43292 ; n43293
g40858 and n42716 n43288 ; n43294
g40859 nor pi1155 n42660 ; n43295
g40860 and n42460_not n43295 ; n43296
g40861 nor n43294 n43296 ; n43297
g40862 and pi1154 n43297_not ; n43298
g40863 nor pi0219 n43293 ; n43299
g40864 and n43298_not n43299 ; n43300
g40865 and pi1153 n38955 ; n43301
g40866 and n42708 n43301_not ; n43302
g40867 and n39668_not n43302 ; n43303
g40868 and pi1091 n42928 ; n43304
g40869 and n42430_not n43304 ; n43305
g40870 and pi1154 n43305_not ; n43306
g40871 and pi0299_not n38946 ; n43307
g40872 and pi1091 n43307_not ; n43308
g40873 and n43306 n43308 ; n43309
g40874 and pi0219 n43303_not ; n43310
g40875 and n43309_not n43310 ; n43311
g40876 nor n43300 n43311 ; n43312
g40877 nor pi0211 n43312 ; n43313
g40878 and pi1155 n38963 ; n43314
g40879 and pi1154 n43314_not ; n43315
g40880 nor pi1155 n38947 ; n43316
g40881 nor n38582 n43316 ; n43317
g40882 nor n13062 n43317 ; n43318
g40883 and pi1091 n43315 ; n43319
g40884 and n43318_not n43319 ; n43320
g40885 nor n38701 n40919 ; n43321
g40886 and n43302 n43321_not ; n43322
g40887 and pi0211 n43322_not ; n43323
g40888 and n43320_not n43323 ; n43324
g40889 nor n43313 n43324 ; n43325
g40890 and pi0267 n43325_not ; n43326
g40891 and n38568 n42448 ; n43327
g40892 nor n42685 n43327 ; n43328
g40893 nor n43290 n43328 ; n43329
g40894 and pi0211 pi1154_not ; n43330
g40895 and n43329_not n43330 ; n43331
g40896 and pi1091 pi1155_not ; n43332
g40897 and n38947_not n43332 ; n43333
g40898 and n38488 n43333_not ; n43334
g40899 and n43305_not n43334 ; n43335
g40900 and pi1154_not n38545 ; n43336
g40901 nor n38670 n43336 ; n43337
g40902 and n38683_not n43337 ; n43338
g40903 and pi1091 n43338 ; n43339
g40904 nor pi0211 n43339 ; n43340
g40905 nor pi0219 n43335 ; n43341
g40906 and n43340_not n43341 ; n43342
g40907 and n43307 n43332 ; n43343
g40908 and n43306 n43343_not ; n43344
g40909 and n42928 n43315 ; n43345
g40910 nor n43344 n43345 ; n43346
g40911 and pi0211 n43346_not ; n43347
g40912 and pi1154 n43344_not ; n43348
g40913 and n38701_not n42708 ; n43349
g40914 and n39667_not n43349 ; n43350
g40915 nor pi0211 n43350 ; n43351
g40916 and n43348_not n43351 ; n43352
g40917 and pi0219 n43347_not ; n43353
g40918 and n43352_not n43353 ; n43354
g40919 nor n43342 n43354 ; n43355
g40920 nor pi0267 n43331 ; n43356
g40921 and n43355_not n43356 ; n43357
g40922 nor n43326 n43357 ; n43358
g40923 and po1038_not n43358 ; n43359
g40924 nor pi0219 n38488 ; n43360
g40925 and n38497_not n43360 ; n43361
g40926 nor n39158 n43361 ; n43362
g40927 and pi1091 n43362_not ; n43363
g40928 nor pi0267 pi1091 ; n43364
g40929 nor n43363 n43364 ; n43365
g40930 and po1038 n43365_not ; n43366
g40931 nor n40910 n43366 ; n43367
g40932 and n43359_not n43367 ; n43368
g40933 nor pi0267 n40980 ; n43369
g40934 and n42538_not n43369 ; n43370
g40935 and pi0267 n42734 ; n43371
g40936 and n40859 n43370_not ; n43372
g40937 and n43371_not n43372 ; n43373
g40938 and n40859_not n43364 ; n43374
g40939 nor n43363 n43374 ; n43375
g40940 and n43373_not n43375 ; n43376
g40941 and po1038 n43376_not ; n43377
g40942 nor n40859 n43358 ; n43378
g40943 and n42777_not n42780 ; n43379
g40944 and n42805 n43379_not ; n43380
g40945 and pi1154 pi1155 ; n43381
g40946 and n41014_not n43381 ; n43382
g40947 and n42782_not n43382 ; n43383
g40948 nor n43380 n43383 ; n43384
g40949 and pi0211 n43384_not ; n43385
g40950 and pi1153 n41055 ; n43386
g40951 and n38487 n42511_not ; n43387
g40952 and n43386_not n43387 ; n43388
g40953 and n42761_not n43388 ; n43389
g40954 and n41039 n42749 ; n43390
g40955 nor pi1155 n43390 ; n43391
g40956 and n43379_not n43391 ; n43392
g40957 nor pi0267 n43392 ; n43393
g40958 and n43389_not n43393 ; n43394
g40959 and n43385_not n43394 ; n43395
g40960 and pi1155 n42583_not ; n43396
g40961 and n41008 n43059_not ; n43397
g40962 and n43396 n43397_not ; n43398
g40963 and n42598_not n43398 ; n43399
g40964 nor n42501 n42517 ; n43400
g40965 and n41009 n43400_not ; n43401
g40966 and pi1154 n43401_not ; n43402
g40967 nor pi1154 n41028 ; n43403
g40968 and n42597_not n43403 ; n43404
g40969 nor pi1155 n43404 ; n43405
g40970 and n43402_not n43405 ; n43406
g40971 and pi0267 n43399_not ; n43407
g40972 and n43406_not n43407 ; n43408
g40973 nor n43395 n43408 ; n43409
g40974 and pi0219 n43409_not ; n43410
g40975 nor pi1155 n42825 ; n43411
g40976 and n43379_not n43411 ; n43412
g40977 and n41072 n43401_not ; n43413
g40978 and n43070 n43413_not ; n43414
g40979 and pi1154 n43414_not ; n43415
g40980 nor pi1154 n42497 ; n43416
g40981 and pi1155 n43416_not ; n43417
g40982 and n41045 n43417_not ; n43418
g40983 nor n43415 n43418 ; n43419
g40984 and pi0211 n43412_not ; n43420
g40985 and n43419_not n43420 ; n43421
g40986 nor n42828 n43386 ; n43422
g40987 and pi1155 n43422_not ; n43423
g40988 and pi1153 n41116_not ; n43424
g40989 nor pi1155 n43424 ; n43425
g40990 and n42605 n43425 ; n43426
g40991 nor pi1154 n43423 ; n43427
g40992 and n43426_not n43427 ; n43428
g40993 nor pi1153 n43098 ; n43429
g40994 and n43425 n43429_not ; n43430
g40995 and pi1154 n43099_not ; n43431
g40996 and n43423_not n43431 ; n43432
g40997 and n43430_not n43432 ; n43433
g40998 nor pi0211 n43428 ; n43434
g40999 and n43433_not n43434 ; n43435
g41000 nor pi0267 n43435 ; n43436
g41001 and n43421_not n43436 ; n43437
g41002 and pi1153_not n41093 ; n43438
g41003 nor n41118 n43438 ; n43439
g41004 and pi1155_not n41072 ; n43440
g41005 and n43439_not n43440 ; n43441
g41006 and n43033 n43396 ; n43442
g41007 and pi1154 n43441_not ; n43443
g41008 and n43442_not n43443 ; n43444
g41009 nor pi1154 n42517 ; n43445
g41010 and n41105_not n43445 ; n43446
g41011 nor pi1155 n43446 ; n43447
g41012 and n40988_not n43445 ; n43448
g41013 and n43447_not n43448 ; n43449
g41014 nor n43444 n43449 ; n43450
g41015 and pi0211 n43450_not ; n43451
g41016 and pi1154 n43439 ; n43452
g41017 and n43447 n43452_not ; n43453
g41018 and pi1154 n41008 ; n43454
g41019 nor n41091 n42804 ; n43455
g41020 and pi1155 n43454_not ; n43456
g41021 and n43455_not n43456 ; n43457
g41022 nor pi0211 n43457 ; n43458
g41023 and n43453_not n43458 ; n43459
g41024 and pi0267 n43459_not ; n43460
g41025 and n43451_not n43460 ; n43461
g41026 nor pi0219 n43461 ; n43462
g41027 and n43437_not n43462 ; n43463
g41028 nor n43410 n43463 ; n43464
g41029 and n40859 n43464_not ; n43465
g41030 nor po1038 n43378 ; n43466
g41031 and n43465_not n43466 ; n43467
g41032 and n40910 n43377_not ; n43468
g41033 and n43467_not n43468 ; n43469
g41034 nor pi0230 n43368 ; n43470
g41035 and n43469_not n43470 ; n43471
g41036 and pi0219 n38963_not ; n43472
g41037 and pi1155_not n43301 ; n43473
g41038 nor pi1154 n43473 ; n43474
g41039 nor n38947 n43474 ; n43475
g41040 and pi1155 n39665 ; n43476
g41041 nor n43475 n43476 ; n43477
g41042 nor n43472 n43477 ; n43478
g41043 and pi0211 n43478_not ; n43479
g41044 and pi0199_not pi1154 ; n43480
g41045 and pi0200 n43480_not ; n43481
g41046 nor n38731 n38962 ; n43482
g41047 and n43481_not n43482 ; n43483
g41048 nor n38510 n43483 ; n43484
g41049 and pi0219 n43484_not ; n43485
g41050 and pi0219_not n43338 ; n43486
g41051 nor pi0211 n43486 ; n43487
g41052 and n43485_not n43487 ; n43488
g41053 nor po1038 n43488 ; n43489
g41054 and n43479_not n43489 ; n43490
g41055 and po1038 n43362 ; n43491
g41056 and pi0230 n43491_not ; n43492
g41057 and n43490_not n43492 ; n43493
g41058 nor n43471 n43493 ; po0424
g41059 and pi0268 pi1152 ; n43495
g41060 nor pi0211 n16479 ; n43496
g41061 and po1038_not n38568 ; n43497
g41062 nor n43496 n43497 ; n43498
g41063 and pi1151_not n43498 ; n43499
g41064 and pi0199_not n16479 ; n43500
g41065 nor n40141 n43500 ; n43501
g41066 and pi1152 n43498_not ; n43502
g41067 and n43501 n43502_not ; n43503
g41068 and pi1150 n43499_not ; n43504
g41069 and n43503_not n43504 ; n43505
g41070 and n43495_not n43505 ; n43506
g41071 and pi1151_not n42389 ; n43507
g41072 nor po1038 n11448 ; n43508
g41073 and po1038 n11446 ; n43509
g41074 nor n43508 n43509 ; n43510
g41075 and pi1151 n43510_not ; n43511
g41076 nor pi1152 n43511 ; n43512
g41077 and n16479_not n42478 ; n43513
g41078 and po1038_not n38581 ; n43514
g41079 nor n43513 n43514 ; n43515
g41080 and pi1151 n43515_not ; n43516
g41081 and pi1152 n43516 ; n43517
g41082 nor pi1150 n43507 ; n43518
g41083 and n43512_not n43518 ; n43519
g41084 and n43517_not n43519 ; n43520
g41085 nor n43506 n43520 ; n43521
g41086 and pi1091 n43521_not ; n43522
g41087 and pi1152 n43505 ; n43523
g41088 and pi1091 n43523_not ; n43524
g41089 and pi0268 n43524_not ; n43525
g41090 nor n43522 n43525 ; n43526
g41091 nor n40909 n43526 ; n43527
g41092 and n42527_not n42572 ; n43528
g41093 and n41012_not n42584 ; n43529
g41094 and pi0219 n42513_not ; n43530
g41095 and n41011_not n43530 ; n43531
g41096 nor n43529 n43531 ; n43532
g41097 nor po1038 n42505 ; n43533
g41098 and n43532 n43533 ; n43534
g41099 nor n43528 n43534 ; n43535
g41100 nor pi1151 n43535 ; n43536
g41101 nor po1038 n42606 ; n43537
g41102 and pi0219 n41048 ; n43538
g41103 and n43537 n43538_not ; n43539
g41104 and n42572 n42733_not ; n43540
g41105 nor n43539 n43540 ; n43541
g41106 and pi1151 n43541_not ; n43542
g41107 nor n43536 n43542 ; n43543
g41108 and pi0268 n43543_not ; n43544
g41109 and po1038 n42538_not ; n43545
g41110 and n42569_not n43545 ; n43546
g41111 and po1038 n42732_not ; n43547
g41112 and n42525_not n43547 ; n43548
g41113 and n43546 n43548_not ; n43549
g41114 and pi0219 n40994_not ; n43550
g41115 nor n42548 n43550 ; n43551
g41116 nor n40993 n43551 ; n43552
g41117 nor po1038 n41026 ; n43553
g41118 and n43552 n43553 ; n43554
g41119 nor n43549 n43554 ; n43555
g41120 and pi1151_not n43555 ; n43556
g41121 nor n40874 n43541 ; n43557
g41122 and pi0219 po1038 ; n43558
g41123 and n40868_not n43558 ; n43559
g41124 and n41032_not n43537 ; n43560
g41125 nor n42534 n43559 ; n43561
g41126 and n43560_not n43561 ; n43562
g41127 nor n43557 n43562 ; n43563
g41128 and pi1151 n43563 ; n43564
g41129 nor pi0268 n43564 ; n43565
g41130 and n43556_not n43565 ; n43566
g41131 nor n43544 n43566 ; n43567
g41132 nor pi1152 n43567 ; n43568
g41133 and n42527_not n43547 ; n43569
g41134 nor n41062 n42599 ; n43570
g41135 nor n43532 n43570 ; n43571
g41136 nor po1038 n43571 ; n43572
g41137 nor n40868 n42587 ; n43573
g41138 and n43572 n43573_not ; n43574
g41139 nor n43569 n43574 ; n43575
g41140 nor pi1151 n43575 ; n43576
g41141 and n40870_not n43533 ; n43577
g41142 and n42733_not n43547 ; n43578
g41143 nor n43539 n43578 ; n43579
g41144 and n43577_not n43579 ; n43580
g41145 and pi1151 n43580_not ; n43581
g41146 and pi0268 n43581_not ; n43582
g41147 and n43576_not n43582 ; n43583
g41148 nor n42512 n43552 ; n43584
g41149 nor po1038 n43584 ; n43585
g41150 nor n43546 n43585 ; n43586
g41151 nor pi1151 n43586 ; n43587
g41152 and n42528_not n43545 ; n43588
g41153 and pi0219_not n41097 ; n43589
g41154 nor n43530 n43589 ; n43590
g41155 nor po1038 n43590 ; n43591
g41156 nor n43549 n43588 ; n43592
g41157 and n43591_not n43592 ; n43593
g41158 and pi1151 n43593_not ; n43594
g41159 nor pi0268 n43594 ; n43595
g41160 and n43587_not n43595 ; n43596
g41161 and pi1152 n43596_not ; n43597
g41162 and n43583_not n43597 ; n43598
g41163 nor n43568 n43598 ; n43599
g41164 and pi1150 n43599_not ; n43600
g41165 and n42534_not n43545 ; n43601
g41166 nor pi0219 n41045 ; n43602
g41167 nor n41002 n43602 ; n43603
g41168 and n43591 n43603 ; n43604
g41169 nor n43601 n43604 ; n43605
g41170 nor pi1151 n43605 ; n43606
g41171 nor po1038 n43532 ; n43607
g41172 nor n43588 n43607 ; n43608
g41173 and pi1151 n43608_not ; n43609
g41174 and pi1152 n43606_not ; n43610
g41175 and n43609_not n43610 ; n43611
g41176 and pi1151_not n43562 ; n43612
g41177 nor n42529 n43559 ; n43613
g41178 and n43572_not n43613 ; n43614
g41179 and pi1151 n43614 ; n43615
g41180 nor pi1152 n43612 ; n43616
g41181 and n43615_not n43616 ; n43617
g41182 nor n43611 n43617 ; n43618
g41183 nor pi0268 n43618 ; n43619
g41184 and pi0219 n42598_not ; n43620
g41185 nor po1038 n42599 ; n43621
g41186 and n43620_not n43621 ; n43622
g41187 nor n43548 n43622 ; n43623
g41188 and pi1151_not n43623 ; n43624
g41189 and n42570_not n43547 ; n43625
g41190 nor n42548 n43620 ; n43626
g41191 and n41102 n43626_not ; n43627
g41192 nor po1038 n43627 ; n43628
g41193 nor n43625 n43628 ; n43629
g41194 and pi1151 n43629 ; n43630
g41195 and pi1152 n43624_not ; n43631
g41196 and n43630_not n43631 ; n43632
g41197 and n40874 n43541_not ; n43633
g41198 nor pi1151 n43633 ; n43634
g41199 nor po1038 n42553 ; n43635
g41200 and n42548_not n43635 ; n43636
g41201 nor n42573 n43636 ; n43637
g41202 and pi1151 n43637 ; n43638
g41203 nor pi1152 n43634 ; n43639
g41204 and n43638_not n43639 ; n43640
g41205 and pi0268 n43640_not ; n43641
g41206 and n43632_not n43641 ; n43642
g41207 nor pi1150 n43642 ; n43643
g41208 and n43619_not n43643 ; n43644
g41209 nor n43600 n43644 ; n43645
g41210 and n40909 n43645_not ; n43646
g41211 nor pi0230 n43527 ; n43647
g41212 and n43646_not n43647 ; n43648
g41213 and pi0230 n43505_not ; n43649
g41214 and n43520_not n43649 ; n43650
g41215 nor n43648 n43650 ; po0425
g41216 and pi0199_not pi1137 ; n43652
g41217 and pi0200 n43652_not ; n43653
g41218 and pi0199 pi1138 ; n43654
g41219 and pi0199_not pi1136 ; n43655
g41220 nor pi0200 n43654 ; n43656
g41221 and n43655_not n43656 ; n43657
g41222 nor n43653 n43657 ; n43658
g41223 and n16479 n43658_not ; n43659
g41224 and pi0211_not pi1138 ; n43660
g41225 and pi0219 n43660 ; n43661
g41226 and pi0211 pi1137 ; n43662
g41227 nor n43221 n43662 ; n43663
g41228 nor pi0219 n43663 ; n43664
g41229 nor n43661 n43664 ; n43665
g41230 and n16479_not n43665 ; n43666
g41231 nor n43659 n43666 ; n43667
g41232 and pi0230 n43667_not ; n43668
g41233 and pi0200_not n43254 ; n43669
g41234 and pi1137 n40951 ; n43670
g41235 nor n43669 n43670 ; n43671
g41236 and n43500 n43671 ; n43672
g41237 and pi1091 n43663_not ; n43673
g41238 and n40141 n43673_not ; n43674
g41239 nor n43672 n43674 ; n43675
g41240 and pi0817_not n40885 ; n43676
g41241 and pi0269 n40885_not ; n43677
g41242 nor pi1091 n43676 ; n43678
g41243 and n43677_not n43678 ; n43679
g41244 nor n43675 n43679 ; n43680
g41245 and pi0817_not n40863 ; n43681
g41246 and pi0269 n40863_not ; n43682
g41247 nor pi1091 n43681 ; n43683
g41248 and n43682_not n43683 ; n43684
g41249 and pi1138 n42455 ; n43685
g41250 and pi0219 n16479_not ; n43686
g41251 and n43685_not n43686 ; n43687
g41252 and pi0200_not pi1091 ; n43688
g41253 and pi1138 n43688 ; n43689
g41254 and pi0199 n43689_not ; n43690
g41255 and n16479 n43690 ; n43691
g41256 nor n43687 n43691 ; n43692
g41257 nor n43684 n43692 ; n43693
g41258 nor n43680 n43693 ; n43694
g41259 nor pi0230 n43694 ; n43695
g41260 nor n43668 n43695 ; po0426
g41261 and pi0805_not n40863 ; n43697
g41262 and pi0270 n40863_not ; n43698
g41263 nor pi1091 n43697 ; n43699
g41264 and n43698_not n43699 ; n43700
g41265 and n42455 n43168 ; n43701
g41266 and n43686 n43701_not ; n43702
g41267 and pi0200_not n43143 ; n43703
g41268 and pi0199 n43703_not ; n43704
g41269 and n16479 n43704 ; n43705
g41270 nor n43702 n43705 ; n43706
g41271 nor n43700 n43706 ; n43707
g41272 and pi0805_not n40885 ; n43708
g41273 and pi0270 n40885_not ; n43709
g41274 nor pi1091 n43708 ; n43710
g41275 and n43709_not n43710 ; n43711
g41276 and pi0211_not pi1139 ; n43712
g41277 and pi0211 pi1140 ; n43713
g41278 nor n43712 n43713 ; n43714
g41279 and pi1091 n43714_not ; n43715
g41280 and n40141 n43715_not ; n43716
g41281 and pi1091 pi1140 ; n43717
g41282 and pi0200 n43717 ; n43718
g41283 and pi1139 n43688 ; n43719
g41284 nor n43718 n43719 ; n43720
g41285 and n43500 n43720 ; n43721
g41286 nor n43716 n43721 ; n43722
g41287 nor n43711 n43722 ; n43723
g41288 nor pi0230 n43707 ; n43724
g41289 and n43723_not n43724 ; n43725
g41290 and pi0219 n43168_not ; n43726
g41291 and pi0219_not n43714 ; n43727
g41292 nor n43726 n43727 ; n43728
g41293 nor n16479 n43728 ; n43729
g41294 and pi0199_not pi1140 ; n43730
g41295 and pi0200 n43730_not ; n43731
g41296 and pi0199 pi1141 ; n43732
g41297 and pi0199_not pi1139 ; n43733
g41298 nor pi0200 n43732 ; n43734
g41299 and n43733_not n43734 ; n43735
g41300 nor n43731 n43735 ; n43736
g41301 and n16479 n43736_not ; n43737
g41302 and pi0230 n43729_not ; n43738
g41303 and n43737_not n43738 ; n43739
g41304 or n43725 n43739 ; po0427
g41305 and pi0211_not pi1147 ; n43741
g41306 and n42444 n43741 ; n43742
g41307 nor pi0271 n40866 ; n43743
g41308 nor n40871 n43743 ; n43744
g41309 and pi0219 n43744_not ; n43745
g41310 nor pi1091 n40887 ; n43746
g41311 and pi0271 n43746_not ; n43747
g41312 nor pi0271 n40888 ; n43748
g41313 nor n43747 n43748 ; n43749
g41314 and pi1091 pi1146 ; n43750
g41315 nor n43749 n43750 ; n43751
g41316 and pi0211_not n43750 ; n43752
g41317 nor n43751 n43752 ; n43753
g41318 and pi1091 n39412 ; n43754
g41319 nor pi0219 n43754 ; n43755
g41320 and n43753_not n43755 ; n43756
g41321 nor n43745 n43756 ; n43757
g41322 nor n16479 n43742 ; n43758
g41323 and n43757_not n43758 ; n43759
g41324 and pi0199 n43744_not ; n43760
g41325 and pi0199_not n43751 ; n43761
g41326 nor n43760 n43761 ; n43762
g41327 and pi0200 n43762_not ; n43763
g41328 and pi1147 n40931 ; n43764
g41329 and pi1091 pi1145 ; n43765
g41330 nor pi0199 n43765 ; n43766
g41331 and n43749_not n43766 ; n43767
g41332 nor n43760 n43767 ; n43768
g41333 nor pi0200 n43764 ; n43769
g41334 and n43768_not n43769 ; n43770
g41335 nor n43763 n43770 ; n43771
g41336 and n16479 n43771_not ; n43772
g41337 nor n43759 n43772 ; n43773
g41338 nor pi0230 n43773 ; n43774
g41339 and pi1147 n42386 ; n43775
g41340 nor n40225 n40235 ; n43776
g41341 nor pi0219 n43776 ; n43777
g41342 nor pi0200 n39393 ; n43778
g41343 and n40339 n43778_not ; n43779
g41344 nor n43775 n43777 ; n43780
g41345 and n43779_not n43780 ; n43781
g41346 nor po1038 n43781 ; n43782
g41347 and pi0219 n43741_not ; n43783
g41348 and n39412_not n41531 ; n43784
g41349 nor n43783 n43784 ; n43785
g41350 and po1038 n43785 ; n43786
g41351 and pi0230 n43786_not ; n43787
g41352 and n43782_not n43787 ; n43788
g41353 nor n43774 n43788 ; po0428
g41354 and po1038 n10844 ; n43790
g41355 nor n13065 n43790 ; n43791
g41356 and pi1150_not n43791 ; n43792
g41357 nor n43498 n43792 ; n43793
g41358 nor pi1149 n43793 ; n43794
g41359 and pi1149 pi1150_not ; n43795
g41360 nor n43498 n43795 ; n43796
g41361 and n43501 n43796_not ; n43797
g41362 nor n43794 n43797 ; n43798
g41363 and pi1091 n43798_not ; n43799
g41364 and pi1148 n43799_not ; n43800
g41365 and pi1150 n42389_not ; n43801
g41366 nor pi1149 n43801 ; n43802
g41367 and pi1091 n43802 ; n43803
g41368 and n16479_not n42712 ; n43804
g41369 and po1038_not n40936 ; n43805
g41370 nor n43804 n43805 ; n43806
g41371 and pi1150_not n43806 ; n43807
g41372 and pi1091 n43515_not ; n43808
g41373 and pi1150 n43808_not ; n43809
g41374 and pi1149 n43807_not ; n43810
g41375 and n43809_not n43810 ; n43811
g41376 nor pi1148 n43803 ; n43812
g41377 and n43811_not n43812 ; n43813
g41378 nor pi0283 n43800 ; n43814
g41379 and n43813_not n43814 ; n43815
g41380 nor pi1150 n43633 ; n43816
g41381 and pi1150 n43623 ; n43817
g41382 nor pi1149 n43816 ; n43818
g41383 and n43817_not n43818 ; n43819
g41384 and pi1150 n43629 ; n43820
g41385 and pi1150_not n43637 ; n43821
g41386 and pi1149 n43821_not ; n43822
g41387 and n43820_not n43822 ; n43823
g41388 nor n43819 n43823 ; n43824
g41389 nor pi1148 n43824 ; n43825
g41390 and pi1150_not n43541 ; n43826
g41391 and pi1150 n43580 ; n43827
g41392 and pi1149 n43826_not ; n43828
g41393 and n43827_not n43828 ; n43829
g41394 and pi1150_not n43535 ; n43830
g41395 and pi1150 n43575 ; n43831
g41396 nor pi1149 n43830 ; n43832
g41397 and n43831_not n43832 ; n43833
g41398 nor n43829 n43833 ; n43834
g41399 and pi1148 n43834_not ; n43835
g41400 and pi0283 n43825_not ; n43836
g41401 and n43835_not n43836 ; n43837
g41402 and pi0272 n43815_not ; n43838
g41403 and n43837_not n43838 ; n43839
g41404 nor pi1150 n43563 ; n43840
g41405 and pi1150 n43593_not ; n43841
g41406 and pi1149 n43840_not ; n43842
g41407 and n43841_not n43842 ; n43843
g41408 and pi1150 n43586_not ; n43844
g41409 nor pi1150 n43555 ; n43845
g41410 nor pi1149 n43845 ; n43846
g41411 and n43844_not n43846 ; n43847
g41412 nor n43843 n43847 ; n43848
g41413 and pi1148 n43848_not ; n43849
g41414 and pi1150 n43605 ; n43850
g41415 nor pi1150 n43562 ; n43851
g41416 nor pi1149 n43851 ; n43852
g41417 and n43850_not n43852 ; n43853
g41418 nor pi1150 n43614 ; n43854
g41419 and pi1150 n43608 ; n43855
g41420 and pi1149 n43855_not ; n43856
g41421 and n43854_not n43856 ; n43857
g41422 nor pi1148 n43853 ; n43858
g41423 and n43857_not n43858 ; n43859
g41424 nor n43849 n43859 ; n43860
g41425 and pi0283 n43860_not ; n43861
g41426 and po1038_not n38550 ; n43862
g41427 nor n40141 n43862 ; n43863
g41428 and n43496_not n43863 ; n43864
g41429 and pi1150 n43864_not ; n43865
g41430 and pi1149 n43865_not ; n43866
g41431 and n43501 n43866 ; n43867
g41432 and pi1148 n43794_not ; n43868
g41433 and n43867_not n43868 ; n43869
g41434 and pi1091 n43869 ; n43870
g41435 nor pi1148 n43802 ; n43871
g41436 nor pi1150 n43510 ; n43872
g41437 and pi1150 n43515 ; n43873
g41438 and pi1149 n43872_not ; n43874
g41439 and n43873_not n43874 ; n43875
g41440 and pi1091 n43875_not ; n43876
g41441 and n43871 n43876 ; n43877
g41442 nor pi0283 n43877 ; n43878
g41443 and n43870_not n43878 ; n43879
g41444 nor pi0272 n43879 ; n43880
g41445 and n43861_not n43880 ; n43881
g41446 nor pi0230 n43839 ; n43882
g41447 and n43881_not n43882 ; n43883
g41448 and pi1149 n43515_not ; n43884
g41449 nor n43866 n43884 ; n43885
g41450 nor n43872 n43885 ; n43886
g41451 and n43871 n43886_not ; n43887
g41452 and pi0230 n43869_not ; n43888
g41453 and n43887_not n43888 ; n43889
g41454 nor n43883 n43889 ; po0429
g41455 nor pi0273 n40867 ; n43891
g41456 nor n40873 n43891 ; n43892
g41457 and pi0219 n43892_not ; n43893
g41458 nor pi0273 n40889 ; n43894
g41459 and n40891 n43894_not ; n43895
g41460 nor pi0219 n43752 ; n43896
g41461 and n43895_not n43896 ; n43897
g41462 nor n43893 n43897 ; n43898
g41463 and po1038 n43898 ; n43899
g41464 and pi0299 n43898 ; n43900
g41465 and pi0199 n43892_not ; n43901
g41466 and pi0200_not n43750 ; n43902
g41467 nor pi0199 n43902 ; n43903
g41468 and n43895_not n43903 ; n43904
g41469 nor pi0299 n43901 ; n43905
g41470 and n43904_not n43905 ; n43906
g41471 nor n43900 n43906 ; n43907
g41472 nor n11447 n41041 ; n43908
g41473 and pi1091 n43908_not ; n43909
g41474 and n43907 n43909_not ; n43910
g41475 nor po1038 n43910 ; n43911
g41476 and pi1091 n42573 ; n43912
g41477 nor n43911 n43912 ; n43913
g41478 and pi1147 n43913_not ; n43914
g41479 and n40447 n43907_not ; n43915
g41480 nor pi1148 n43915 ; n43916
g41481 and pi1091 n38519 ; n43917
g41482 nor n43898 n43917 ; n43918
g41483 and pi0299 n43918_not ; n43919
g41484 and n40932 n43763_not ; n43920
g41485 nor n43906 n43920 ; n43921
g41486 and n43919_not n43921 ; n43922
g41487 nor po1038 n43922 ; n43923
g41488 and n40080 n42444 ; n43924
g41489 and pi1148 n43924_not ; n43925
g41490 and n43923_not n43925 ; n43926
g41491 nor n43916 n43926 ; n43927
g41492 nor n43899 n43927 ; n43928
g41493 and n43914_not n43928 ; n43929
g41494 nor pi0230 n43929 ; n43930
g41495 and pi1146 n41404_not ; n43931
g41496 and n43791_not n43931 ; n43932
g41497 nor pi0211 n40234 ; n43933
g41498 and n40141 n43933_not ; n43934
g41499 and pi1146_not n10809 ; n43935
g41500 and n43500 n43935_not ; n43936
g41501 nor n43934 n43936 ; n43937
g41502 and pi1147 n43937_not ; n43938
g41503 nor pi1148 n43932 ; n43939
g41504 and n43938_not n43939 ; n43940
g41505 and pi0199_not pi1147 ; n43941
g41506 and pi0200 n43941_not ; n43942
g41507 nor n43935 n43942 ; n43943
g41508 and n16479 n43943 ; n43944
g41509 and pi1146_not n10844 ; n43945
g41510 and pi1147 n40141 ; n43946
g41511 nor n43496 n43946 ; n43947
g41512 nor n43945 n43947 ; n43948
g41513 and pi1148 n43944_not ; n43949
g41514 and n43948_not n43949 ; n43950
g41515 and pi0230 n43940_not ; n43951
g41516 and n43950_not n43951 ; n43952
g41517 or n43930 n43952 ; po0430
g41518 and pi0200_not n43765 ; n43954
g41519 and pi0659_not n40863 ; n43955
g41520 and pi0274 n40863_not ; n43956
g41521 nor pi1091 n43955 ; n43957
g41522 and n43956_not n43957 ; n43958
g41523 and pi0199 n43954_not ; n43959
g41524 and n43958_not n43959 ; n43960
g41525 and pi0659_not n40885 ; n43961
g41526 and pi0274 n40885_not ; n43962
g41527 nor pi1091 n43961 ; n43963
g41528 and n43962_not n43963 ; n43964
g41529 nor n43180 n43964 ; n43965
g41530 and pi0200 n43965_not ; n43966
g41531 nor n43135 n43964 ; n43967
g41532 nor pi0200 n43967 ; n43968
g41533 nor pi0199 n43966 ; n43969
g41534 and n43968_not n43969 ; n43970
g41535 and n16479 n43960_not ; n43971
g41536 and n43970_not n43971 ; n43972
g41537 and pi0211 n43965_not ; n43973
g41538 nor pi0211 n43967 ; n43974
g41539 nor pi0219 n43973 ; n43975
g41540 and n43974_not n43975 ; n43976
g41541 and pi0219 n43754_not ; n43977
g41542 and n43958_not n43977 ; n43978
g41543 nor n16479 n43978 ; n43979
g41544 and n43976_not n43979 ; n43980
g41545 nor pi0230 n43972 ; n43981
g41546 and n43980_not n43981 ; n43982
g41547 nor n38508 n40225 ; n43983
g41548 nor pi0219 n38425 ; n43984
g41549 and n39413_not n43984 ; n43985
g41550 nor n43983 n43985 ; n43986
g41551 and n38436_not n40332 ; n43987
g41552 and n40788 n43987_not ; n43988
g41553 nor n43986 n43988 ; n43989
g41554 nor po1038 n43989 ; n43990
g41555 nor n40221 n43985 ; n43991
g41556 and pi0230 n43990_not ; n43992
g41557 and n43991_not n43992 ; n43993
g41558 nor n43982 n43993 ; po0431
g41559 and pi1151 n43498_not ; n43995
g41560 and pi1149 n43501 ; n43996
g41561 and n43995_not n43996 ; n43997
g41562 and pi1149_not n43516 ; n43998
g41563 nor n43997 n43998 ; n43999
g41564 and pi1150 n43999_not ; n44000
g41565 and pi1151_not n43791 ; n44001
g41566 and pi1149 n43498_not ; n44002
g41567 and n44001_not n44002 ; n44003
g41568 and pi1149_not pi1151 ; n44004
g41569 and n42389_not n44004 ; n44005
g41570 nor pi1150 n44005 ; n44006
g41571 and n44003_not n44006 ; n44007
g41572 nor n44000 n44007 ; n44008
g41573 and pi1091 n44008_not ; n44009
g41574 and pi1151_not n41484 ; n44010
g41575 and n43806_not n44010 ; n44011
g41576 nor n44009 n44011 ; n44012
g41577 and pi0275 n44012_not ; n44013
g41578 and n43498 n43795 ; n44014
g41579 and n40607 n42389_not ; n44015
g41580 and pi1151_not n43510 ; n44016
g41581 and pi1150 n44016_not ; n44017
g41582 and n43516_not n44017 ; n44018
g41583 nor pi1149 n44015 ; n44019
g41584 and n44018_not n44019 ; n44020
g41585 nor n43997 n44014 ; n44021
g41586 and n44020_not n44021 ; n44022
g41587 and pi1091 n44022 ; n44023
g41588 nor pi0275 n44023 ; n44024
g41589 nor n40908 n44024 ; n44025
g41590 and n44013_not n44025 ; n44026
g41591 and pi1150_not n43605 ; n44027
g41592 and pi1151 n43855_not ; n44028
g41593 and n44027_not n44028 ; n44029
g41594 and pi1150 n43614_not ; n44030
g41595 nor pi1151 n43851 ; n44031
g41596 and n44030_not n44031 ; n44032
g41597 nor n44029 n44032 ; n44033
g41598 nor pi0275 n44033 ; n44034
g41599 and pi1150 n43637 ; n44035
g41600 nor n43816 n44035 ; n44036
g41601 nor pi1151 n44036 ; n44037
g41602 and pi1150_not n43623 ; n44038
g41603 nor n43820 n44038 ; n44039
g41604 and pi1151 n44039_not ; n44040
g41605 and pi0275 n44037_not ; n44041
g41606 and n44040_not n44041 ; n44042
g41607 nor pi1149 n44042 ; n44043
g41608 and n44034_not n44043 ; n44044
g41609 and pi1150 n43563_not ; n44045
g41610 nor pi1151 n44045 ; n44046
g41611 and n43845_not n44046 ; n44047
g41612 nor pi1150 n43586 ; n44048
g41613 and pi1151 n43841_not ; n44049
g41614 and n44048_not n44049 ; n44050
g41615 nor pi0275 n44047 ; n44051
g41616 and n44050_not n44051 ; n44052
g41617 and pi1151 n43575_not ; n44053
g41618 nor pi1150 n43536 ; n44054
g41619 and n44053_not n44054 ; n44055
g41620 nor pi1151 n43541 ; n44056
g41621 and pi1150 n44056_not ; n44057
g41622 and n43581_not n44057 ; n44058
g41623 and pi0275 n44058_not ; n44059
g41624 and n44055_not n44059 ; n44060
g41625 and pi1149 n44052_not ; n44061
g41626 and n44060_not n44061 ; n44062
g41627 and n40908 n44044_not ; n44063
g41628 and n44062_not n44063 ; n44064
g41629 nor n44026 n44064 ; n44065
g41630 nor pi0230 n44065 ; n44066
g41631 and pi0230 n44022 ; n44067
g41632 or n44066 n44067 ; po0432
g41633 nor pi0276 n40886 ; n44069
g41634 and n43746 n44069_not ; n44070
g41635 nor n38419 n40210 ; n44071
g41636 and pi1091 n44071_not ; n44072
g41637 and n40141 n44072_not ; n44073
g41638 and pi1145 n40951 ; n44074
g41639 nor n43181 n44074 ; n44075
g41640 and n43500 n44075 ; n44076
g41641 nor n44073 n44076 ; n44077
g41642 nor n44070 n44077 ; n44078
g41643 nor pi0276 n40864 ; n44079
g41644 and n40870 n44079_not ; n44080
g41645 and n43686 n43752_not ; n44081
g41646 and pi0199 n43902_not ; n44082
g41647 and n16479 n44082 ; n44083
g41648 nor n44081 n44083 ; n44084
g41649 nor n44080 n44084 ; n44085
g41650 nor pi0230 n44078 ; n44086
g41651 and n44085_not n44086 ; n44087
g41652 and n38434_not n41294 ; n44088
g41653 nor n40330 n44088 ; n44089
g41654 and n16479 n44089_not ; n44090
g41655 nor pi0219 n44071 ; n44091
g41656 and pi1146 n38519 ; n44092
g41657 nor n44091 n44092 ; n44093
g41658 and n16479_not n44093 ; n44094
g41659 and pi0230 n44090_not ; n44095
g41660 and n44094_not n44095 ; n44096
g41661 or n44087 n44096 ; po0433
g41662 and pi0200_not n43150 ; n44098
g41663 and pi0820_not n40863 ; n44099
g41664 and pi0277 n40863_not ; n44100
g41665 nor pi1091 n44099 ; n44101
g41666 and n44100_not n44101 ; n44102
g41667 and pi0199 n44098_not ; n44103
g41668 and n44102_not n44103 ; n44104
g41669 and pi0820_not n40885 ; n44105
g41670 and pi0277 n40885_not ; n44106
g41671 nor pi1091 n44105 ; n44107
g41672 and n44106_not n44107 ; n44108
g41673 nor n43717 n44108 ; n44109
g41674 nor pi0200 n44109 ; n44110
g41675 nor n43143 n44108 ; n44111
g41676 and pi0200 n44111_not ; n44112
g41677 nor pi0199 n44110 ; n44113
g41678 and n44112_not n44113 ; n44114
g41679 and n16479 n44104_not ; n44115
g41680 and n44114_not n44115 ; n44116
g41681 and pi0219 n43210_not ; n44117
g41682 nor n43157 n44117 ; n44118
g41683 nor n44102 n44118 ; n44119
g41684 nor pi0211 n44109 ; n44120
g41685 and pi0211 n44111_not ; n44121
g41686 nor pi0219 n44120 ; n44122
g41687 and n44121_not n44122 ; n44123
g41688 nor n16479 n44119 ; n44124
g41689 and n44123_not n44124 ; n44125
g41690 nor n44116 n44125 ; n44126
g41691 nor pi0230 n44126 ; n44127
g41692 and pi0211 pi1141 ; n44128
g41693 and pi0211_not pi1140 ; n44129
g41694 nor pi0219 n44128 ; n44130
g41695 and n44129_not n44130 ; n44131
g41696 nor n44117 n44131 ; n44132
g41697 nor n16479 n44132 ; n44133
g41698 and n38433 n43730_not ; n44134
g41699 and pi0200 n43173_not ; n44135
g41700 nor n44134 n44135 ; n44136
g41701 and n16479 n44136_not ; n44137
g41702 and pi0230 n44133_not ; n44138
g41703 and n44137_not n44138 ; n44139
g41704 or n44127 n44139 ; po0434
g41705 nor pi0278 n40863 ; n44141
g41706 and pi0976_not n40863 ; n44142
g41707 nor pi1091 n44141 ; n44143
g41708 and n44142_not n44143 ; n44144
g41709 and pi0199 n44144_not ; n44145
g41710 and pi1091 pi1132_not ; n44146
g41711 and pi0976 n40885 ; n44147
g41712 and pi0278 n40885_not ; n44148
g41713 nor pi1091 n44147 ; n44149
g41714 and n44148_not n44149 ; n44150
g41715 nor n44146 n44150 ; n44151
g41716 nor pi0199 n44151 ; n44152
g41717 nor n44145 n44152 ; n44153
g41718 nor pi0200 n44153 ; n44154
g41719 and pi1091 pi1133_not ; n44155
g41720 nor n44150 n44155 ; n44156
g41721 nor pi0199 n44156 ; n44157
g41722 nor n44145 n44157 ; n44158
g41723 and pi0200 n44158_not ; n44159
g41724 nor pi0299 n44159 ; n44160
g41725 and n44154_not n44160 ; n44161
g41726 and pi0219 n44144_not ; n44162
g41727 and pi0211 pi1133_not ; n44163
g41728 nor pi0211 pi1132 ; n44164
g41729 nor n44163 n44164 ; n44165
g41730 and pi1091 n44165_not ; n44166
g41731 nor n44150 n44166 ; n44167
g41732 nor pi0219 n44167 ; n44168
g41733 nor n44162 n44168 ; n44169
g41734 and pi0299 n44169 ; n44170
g41735 nor n44161 n44170 ; n44171
g41736 nor po1038 n44171 ; n44172
g41737 and po1038 n44169 ; n44173
g41738 nor pi0230 n44173 ; n44174
g41739 and n44172_not n44174 ; n44175
g41740 and n39374 n44165 ; n44176
g41741 and pi0199_not pi1132 ; n44177
g41742 nor pi0200 n44177 ; n44178
g41743 and pi0199_not pi1133 ; n44179
g41744 and pi0200 n44179_not ; n44180
g41745 nor pi0299 n44180 ; n44181
g41746 and n44178_not n44181 ; n44182
g41747 and n38508 n44165 ; n44183
g41748 nor n44182 n44183 ; n44184
g41749 nor po1038 n44184 ; n44185
g41750 and pi0230 n44176_not ; n44186
g41751 and n44185_not n44186 ; n44187
g41752 nor n44175 n44187 ; n44188
g41753 nor pi1134 n44188 ; n44189
g41754 and n10809 n44177_not ; n44190
g41755 and n44181 n44190_not ; n44191
g41756 nor n42627 n44183 ; n44192
g41757 and n44191_not n44192 ; n44193
g41758 nor po1038 n44193 ; n44194
g41759 nor pi0219 n44165 ; n44195
g41760 nor n40081 n44195 ; n44196
g41761 and pi0230 n44194_not ; n44197
g41762 and n44196_not n44197 ; n44198
g41763 and n40931_not n44154 ; n44199
g41764 and n44160 n44199_not ; n44200
g41765 and n13062 n42455 ; n44201
g41766 nor n44170 n44201 ; n44202
g41767 and n44200_not n44202 ; n44203
g41768 nor po1038 n44203 ; n44204
g41769 and n43924_not n44174 ; n44205
g41770 and n44204_not n44205 ; n44206
g41771 nor n44198 n44206 ; n44207
g41772 and pi1134 n44207_not ; n44208
g41773 nor n44189 n44208 ; po0435
g41774 nor pi0279 n40863 ; n44210
g41775 and pi0958_not n40863 ; n44211
g41776 nor pi1091 n44210 ; n44212
g41777 and n44211_not n44212 ; n44213
g41778 and pi1135 n43688 ; n44214
g41779 nor n44213 n44214 ; n44215
g41780 and pi0199 n44215_not ; n44216
g41781 and pi0958 n40885 ; n44217
g41782 and pi0279 n40885_not ; n44218
g41783 nor pi1091 n44217 ; n44219
g41784 and n44218_not n44219 ; n44220
g41785 and pi1133_not n43688 ; n44221
g41786 nor pi0199 n44221 ; n44222
g41787 and n44220_not n44222 ; n44223
g41788 nor n44216 n44223 ; n44224
g41789 and n16479 n44224_not ; n44225
g41790 and n40951_not n44225 ; n44226
g41791 nor n42424 n44155 ; n44227
g41792 and n44220_not n44227 ; n44228
g41793 nor pi0219 n44228 ; n44229
g41794 and pi1135 n42455 ; n44230
g41795 and pi0219 n44230_not ; n44231
g41796 and n44213_not n44231 ; n44232
g41797 nor n16479 n44232 ; n44233
g41798 and n44229_not n44233 ; n44234
g41799 nor pi0230 n44234 ; n44235
g41800 and n44226_not n44235 ; n44236
g41801 and pi1135 n38519 ; n44237
g41802 nor pi0211 pi1133 ; n44238
g41803 nor pi0219 n44238 ; n44239
g41804 and pi0211_not n44239 ; n44240
g41805 nor n44237 n44240 ; n44241
g41806 and po1038 n44241_not ; n44242
g41807 and pi0199 pi1135 ; n44243
g41808 nor n44179 n44243 ; n44244
g41809 and n38568 n44244_not ; n44245
g41810 and pi0299 n44241_not ; n44246
g41811 nor n44245 n44246 ; n44247
g41812 nor po1038 n44247 ; n44248
g41813 and pi0230 n44242_not ; n44249
g41814 and n44248_not n44249 ; n44250
g41815 nor n44236 n44250 ; n44251
g41816 nor pi1134 n44251 ; n44252
g41817 and pi1133_not n10809 ; n44253
g41818 and pi0200_not pi1135 ; n44254
g41819 and pi0199 n44254_not ; n44255
g41820 nor n44253 n44255 ; n44256
g41821 and n16479 n44256_not ; n44257
g41822 nor n44237 n44239 ; n44258
g41823 and n16479_not n44258 ; n44259
g41824 nor n44257 n44259 ; n44260
g41825 and pi0230 n44260_not ; n44261
g41826 and pi1091 n44238_not ; n44262
g41827 and n40141 n44262 ; n44263
g41828 nor n44225 n44263 ; n44264
g41829 and n44235 n44264 ; n44265
g41830 nor n44261 n44265 ; n44266
g41831 and pi1134 n44266_not ; n44267
g41832 nor n44252 n44267 ; po0436
g41833 and pi0211_not pi1135 ; n44269
g41834 and pi0211 pi1136 ; n44270
g41835 nor n44269 n44270 ; n44271
g41836 and pi1091 n44271 ; n44272
g41837 nor pi0280 n40885 ; n44273
g41838 and pi0914 n40885 ; n44274
g41839 nor pi1091 n44273 ; n44275
g41840 and n44274_not n44275 ; n44276
g41841 nor n44272 n44276 ; n44277
g41842 nor pi0219 n44277 ; n44278
g41843 and pi0211_not pi1137 ; n44279
g41844 and pi0219 n44279_not ; n44280
g41845 nor n43157 n44280 ; n44281
g41846 and pi0914_not n40863 ; n44282
g41847 and pi0280 n40863_not ; n44283
g41848 nor pi1091 n44282 ; n44284
g41849 and n44283_not n44284 ; n44285
g41850 nor n44281 n44285 ; n44286
g41851 nor n44278 n44286 ; n44287
g41852 nor n16479 n44287 ; n44288
g41853 and pi1137 n43688 ; n44289
g41854 nor n44285 n44289 ; n44290
g41855 and pi0199 n44290_not ; n44291
g41856 and pi0200 pi1136 ; n44292
g41857 and pi1091 n44254_not ; n44293
g41858 and n44292_not n44293 ; n44294
g41859 nor pi0199 n44294 ; n44295
g41860 and n44276_not n44295 ; n44296
g41861 and n16479 n44291_not ; n44297
g41862 and n44296_not n44297 ; n44298
g41863 nor n44288 n44298 ; n44299
g41864 nor pi0230 n44299 ; n44300
g41865 and pi0200 n43655_not ; n44301
g41866 and pi0199 pi1137 ; n44302
g41867 nor pi0200 n43228 ; n44303
g41868 and n44302_not n44303 ; n44304
g41869 nor n44301 n44304 ; n44305
g41870 and n16479 n44305 ; n44306
g41871 and pi0219_not n44271 ; n44307
g41872 nor n44280 n44307 ; n44308
g41873 and n16479_not n44308 ; n44309
g41874 and pi0230 n44306_not ; n44310
g41875 and n44309_not n44310 ; n44311
g41876 nor n44300 n44311 ; po0437
g41877 and pi0199_not pi1138 ; n44313
g41878 and pi0200 n44313_not ; n44314
g41879 and pi0199 pi1139 ; n44315
g41880 nor pi0200 n43652 ; n44316
g41881 and n44315_not n44316 ; n44317
g41882 nor n44314 n44317 ; n44318
g41883 and n16479 n44318_not ; n44319
g41884 and pi0219 n43712 ; n44320
g41885 and pi0211 pi1138 ; n44321
g41886 nor n44279 n44321 ; n44322
g41887 nor pi0219 n44322 ; n44323
g41888 nor n44320 n44323 ; n44324
g41889 and n16479_not n44324 ; n44325
g41890 nor n44319 n44325 ; n44326
g41891 and pi0230 n44326_not ; n44327
g41892 and pi0830_not n40885 ; n44328
g41893 and pi0281 n40885_not ; n44329
g41894 nor pi1091 n44328 ; n44330
g41895 and n44329_not n44330 ; n44331
g41896 and pi1091 n44322_not ; n44332
g41897 and n40141 n44332_not ; n44333
g41898 and pi1138 n40951 ; n44334
g41899 nor n44289 n44334 ; n44335
g41900 and n43500 n44335 ; n44336
g41901 nor n44333 n44336 ; n44337
g41902 nor n44331 n44337 ; n44338
g41903 and pi0830_not n40863 ; n44339
g41904 and pi0281 n40863_not ; n44340
g41905 nor pi1091 n44339 ; n44341
g41906 and n44340_not n44341 ; n44342
g41907 and pi1139 n42455 ; n44343
g41908 and n43686 n44343_not ; n44344
g41909 and pi0199 n43719_not ; n44345
g41910 and n16479 n44345 ; n44346
g41911 nor n44344 n44346 ; n44347
g41912 nor n44342 n44347 ; n44348
g41913 nor n44338 n44348 ; n44349
g41914 nor pi0230 n44349 ; n44350
g41915 nor n44327 n44350 ; po0438
g41916 and pi0200 n43733_not ; n44352
g41917 and pi0199 pi1140 ; n44353
g41918 nor pi0200 n44313 ; n44354
g41919 and n44353_not n44354 ; n44355
g41920 nor n44352 n44355 ; n44356
g41921 and n16479 n44356_not ; n44357
g41922 and pi0219 n44129 ; n44358
g41923 and pi0211 pi1139 ; n44359
g41924 nor n43660 n44359 ; n44360
g41925 nor pi0219 n44360 ; n44361
g41926 nor n44358 n44361 ; n44362
g41927 and n16479_not n44362 ; n44363
g41928 nor n44357 n44363 ; n44364
g41929 and pi0230 n44364_not ; n44365
g41930 and pi0836_not n40885 ; n44366
g41931 and pi0282 n40885_not ; n44367
g41932 nor pi1091 n44366 ; n44368
g41933 and n44367_not n44368 ; n44369
g41934 and pi1091 n44360_not ; n44370
g41935 and n40141 n44370_not ; n44371
g41936 and pi1139 n40951 ; n44372
g41937 nor n43689 n44372 ; n44373
g41938 and n43500 n44373 ; n44374
g41939 nor n44371 n44374 ; n44375
g41940 nor n44369 n44375 ; n44376
g41941 and pi0836_not n40863 ; n44377
g41942 and pi0282 n40863_not ; n44378
g41943 nor pi1091 n44377 ; n44379
g41944 and n44378_not n44379 ; n44380
g41945 and pi1140 n42455 ; n44381
g41946 and n43686 n44381_not ; n44382
g41947 and pi0200_not n43717 ; n44383
g41948 and pi0199 n44383_not ; n44384
g41949 and n16479 n44384 ; n44385
g41950 nor n44382 n44385 ; n44386
g41951 nor n44380 n44386 ; n44387
g41952 nor n44376 n44387 ; n44388
g41953 nor pi0230 n44388 ; n44389
g41954 nor n44365 n44389 ; po0439
g41955 and pi1147 n43791_not ; n44391
g41956 and pi1149 n42389_not ; n44392
g41957 nor n44391 n44392 ; n44393
g41958 nor pi1148 n44393 ; n44394
g41959 and n43884 n44391_not ; n44395
g41960 and pi1147 n43501_not ; n44396
g41961 and pi1149_not n43510 ; n44397
g41962 and n44396_not n44397 ; n44398
g41963 and pi1148 n44395_not ; n44399
g41964 and n44398_not n44399 ; n44400
g41965 and pi0230 n44394_not ; n44401
g41966 and n44400_not n44401 ; n44402
g41967 and pi1147_not n43637 ; n44403
g41968 and pi1147 n43541 ; n44404
g41969 and pi1148 n44404_not ; n44405
g41970 and n44403_not n44405 ; n44406
g41971 and pi1147 n43535 ; n44407
g41972 nor pi1147 n43633 ; n44408
g41973 nor pi1148 n44408 ; n44409
g41974 and n44407_not n44409 ; n44410
g41975 nor pi1149 n44406 ; n44411
g41976 and n44410_not n44411 ; n44412
g41977 and pi1147_not n43629 ; n44413
g41978 and pi1147 n43580 ; n44414
g41979 and pi1148 n44414_not ; n44415
g41980 and n44413_not n44415 ; n44416
g41981 and pi1147_not n43623 ; n44417
g41982 and pi1147 n43575 ; n44418
g41983 nor pi1148 n44417 ; n44419
g41984 and n44418_not n44419 ; n44420
g41985 and pi1149 n44416_not ; n44421
g41986 and n44420_not n44421 ; n44422
g41987 and pi0283 n44412_not ; n44423
g41988 and n44422_not n44423 ; n44424
g41989 and pi1147_not n43605 ; n44425
g41990 and pi1147 n43586 ; n44426
g41991 and pi1149 n44425_not ; n44427
g41992 and n44426_not n44427 ; n44428
g41993 nor pi1147 n43562 ; n44429
g41994 and pi1147 n43555 ; n44430
g41995 nor pi1149 n44429 ; n44431
g41996 and n44430_not n44431 ; n44432
g41997 nor pi1148 n44432 ; n44433
g41998 and n44428_not n44433 ; n44434
g41999 and pi1147_not n43608 ; n44435
g42000 and pi1147 n43593 ; n44436
g42001 and pi1149 n44436_not ; n44437
g42002 and n44435_not n44437 ; n44438
g42003 and pi1147 n43563 ; n44439
g42004 nor pi1147 n43614 ; n44440
g42005 nor pi1149 n44439 ; n44441
g42006 and n44440_not n44441 ; n44442
g42007 and pi1148 n44438_not ; n44443
g42008 and n44442_not n44443 ; n44444
g42009 nor pi0283 n44434 ; n44445
g42010 and n44444_not n44445 ; n44446
g42011 nor pi0230 n44424 ; n44447
g42012 and n44446_not n44447 ; n44448
g42013 nor n44402 n44448 ; po0440
g42014 nor pi0284 n42902 ; n44450
g42015 and pi1143 n42902 ; n44451
g42016 and n40143_not n44451 ; n44452
g42017 or n44450 n44452 ; po0441
g42018 and n2572 n10399_not ; n44454
g42019 and n7420_not n44454 ; n44455
g42020 and pi0286 n44455 ; n44456
g42021 and pi0288 pi0289 ; n44457
g42022 and n44456 n44457 ; n44458
g42023 and pi0285 n44458 ; n44459
g42024 and pi0285 n44454 ; n44460
g42025 nor n44458 n44460 ; n44461
g42026 nor po1038 n44459 ; n44462
g42027 and n44461_not n44462 ; n44463
g42028 and po1038_not n44458 ; n44464
g42029 and pi0286_not n7420 ; n44465
g42030 and pi0288_not n44465 ; n44466
g42031 and pi0289_not n44466 ; n44467
g42032 and pi0285 n44467_not ; n44468
g42033 and n44464_not n44468 ; n44469
g42034 nor n44463 n44469 ; n44470
g42035 nor pi0793 n44470 ; po0442
g42036 nor pi0288 n7424 ; n44472
g42037 and n7420 n44472 ; n44473
g42038 and pi0286 n44473_not ; n44474
g42039 and pi0286_not n44473 ; n44475
g42040 and po1038 n44474_not ; n44476
g42041 and n44475_not n44476 ; n44477
g42042 and n7420 n44454_not ; n44478
g42043 and pi0286 n44478_not ; n44479
g42044 and n44454_not n44465 ; n44480
g42045 nor n44479 n44480 ; n44481
g42046 and n44472 n44481_not ; n44482
g42047 nor pi0286 n44455 ; n44483
g42048 and pi0288 n44456_not ; n44484
g42049 and n44483_not n44484 ; n44485
g42050 nor po1038 n44482 ; n44486
g42051 and n44485_not n44486 ; n44487
g42052 nor pi0793 n44477 ; n44488
g42053 and n44487_not n44488 ; po0443
g42054 and pi0287_not pi0457 ; n44490
g42055 nor pi0332 n44490 ; po0444
g42056 and pi0288 n7420_not ; n44492
g42057 nor n44473 n44492 ; n44493
g42058 and po1038_not n44454 ; po0637
g42059 and n44493_not po0637 ; n44495
g42060 and n44493 po0637_not ; n44496
g42061 nor pi0793 n44495 ; n44497
g42062 and n44496_not n44497 ; po0445
g42063 and pi0289 n44466_not ; n44499
g42064 and pi0285 pi0289_not ; n44500
g42065 and n44466 n44500 ; n44501
g42066 and po1038 n44499_not ; n44502
g42067 and n44501_not n44502 ; n44503
g42068 and pi0289_not n44484 ; n44504
g42069 and n44480 n44500 ; n44505
g42070 and pi0289 n44480_not ; n44506
g42071 nor pi0288 n44505 ; n44507
g42072 and n44506_not n44507 ; n44508
g42073 nor n44458 n44504 ; n44509
g42074 and n44508_not n44509 ; n44510
g42075 nor po1038 n44510 ; n44511
g42076 nor pi0793 n44503 ; n44512
g42077 and n44511_not n44512 ; po0446
g42078 and pi0290_not pi0476 ; n44514
g42079 nor pi0476 pi1048 ; n44515
g42080 nor n44514 n44515 ; po0447
g42081 and pi0291_not pi0476 ; n44517
g42082 nor pi0476 pi1049 ; n44518
g42083 nor n44517 n44518 ; po0448
g42084 and pi0292_not pi0476 ; n44520
g42085 nor pi0476 pi1084 ; n44521
g42086 nor n44520 n44521 ; po0449
g42087 and pi0293_not pi0476 ; n44523
g42088 nor pi0476 pi1059 ; n44524
g42089 nor n44523 n44524 ; po0450
g42090 and pi0294_not pi0476 ; n44526
g42091 nor pi0476 pi1072 ; n44527
g42092 nor n44526 n44527 ; po0451
g42093 and pi0295_not pi0476 ; n44529
g42094 nor pi0476 pi1053 ; n44530
g42095 nor n44529 n44530 ; po0452
g42096 and pi0296_not pi0476 ; n44532
g42097 nor pi0476 pi1037 ; n44533
g42098 nor n44532 n44533 ; po0453
g42099 and pi0297_not pi0476 ; n44535
g42100 nor pi0476 pi1044 ; n44536
g42101 nor n44535 n44536 ; po0454
g42102 and pi0478_not pi1044 ; n44538
g42103 and pi0298 pi0478 ; n44539
g42104 or n44538 n44539 ; po0455
g42105 and pi0054 n2521 ; n44541
g42106 and pi0054_not n13153 ; n44542
g42107 and n13411 n44542 ; n44543
g42108 nor n44541 n44543 ; n44544
g42109 and n2621 n8880 ; n44545
g42110 and n44544_not n44545 ; n44546
g42111 nor pi0039 n44546 ; n44547
g42112 nor n11263 n44547 ; po0456
g42113 and pi0057 pi0059_not ; n44549
g42114 and n10068 n44549 ; n44550
g42115 and pi0312_not n44550 ; n44551
g42116 and pi0300 n44551_not ; n44552
g42117 and pi0300_not n44551 ; n44553
g42118 nor pi0055 n44553 ; n44554
g42119 nand n44552_not n44554 ; po0457
g42120 and pi0301_not n44554 ; n44556
g42121 and pi0055_not pi0301 ; n44557
g42122 and n44553 n44557 ; n44558
g42123 or n44556 n44558 ; po0458
g42124 and n5836 po1038_not ; n44560
g42125 nor pi0222 pi0223 ; n44561
g42126 and pi0937 n44561_not ; n44562
g42127 and pi0273 n3351 ; n44563
g42128 nor n44562 n44563 ; n44564
g42129 and n44560 n44564 ; n44565
g42130 and n2603_not n44565 ; n44566
g42131 and n3449 n16479_not ; n44567
g42132 nor n44565 n44567 ; n44568
g42133 and pi0237 n44568_not ; n44569
g42134 and n5780 n16479_not ; n44570
g42135 nor n44560 n44570 ; n44571
g42136 and pi1148_not n44571 ; n44572
g42137 and pi0215_not n3310 ; n44573
g42138 and pi0273_not n44573 ; n44574
g42139 and pi0833 n7570 ; n44575
g42140 and pi0937_not n44575 ; n44576
g42141 nor n44574 n44576 ; n44577
g42142 nor n16479 n44577 ; n44578
g42143 nor n44566 n44578 ; n44579
g42144 and n44569_not n44579 ; n44580
g42145 and n44572_not n44580 ; po0459
g42146 and pi0478_not pi1049 ; n44582
g42147 and pi0303 pi0478 ; n44583
g42148 or n44582 n44583 ; po0460
g42149 and pi0478_not pi1048 ; n44585
g42150 and pi0304 pi0478 ; n44586
g42151 or n44585 n44586 ; po0461
g42152 and pi0478_not pi1084 ; n44588
g42153 and pi0305 pi0478 ; n44589
g42154 or n44588 n44589 ; po0462
g42155 and pi0478_not pi1059 ; n44591
g42156 and pi0306 pi0478 ; n44592
g42157 or n44591 n44592 ; po0463
g42158 and pi0478_not pi1053 ; n44594
g42159 and pi0307 pi0478 ; n44595
g42160 or n44594 n44595 ; po0464
g42161 and pi0478_not pi1037 ; n44597
g42162 and pi0308 pi0478 ; n44598
g42163 or n44597 n44598 ; po0465
g42164 and pi0478_not pi1072 ; n44600
g42165 and pi0309 pi0478 ; n44601
g42166 or n44600 n44601 ; po0466
g42167 and pi1147 n44571 ; n44603
g42168 and pi0222 pi0934_not ; n44604
g42169 and pi0271_not n3351 ; n44605
g42170 nor n44604 n44605 ; n44606
g42171 and n44560 n44606 ; n44607
g42172 and n3448_not n44570 ; n44608
g42173 and pi0934 n2526_not ; n44609
g42174 and pi0271 n3310 ; n44610
g42175 nor n44609 n44610 ; n44611
g42176 and n44608 n44611_not ; n44612
g42177 nor n44567 n44607 ; n44613
g42178 and n44612_not n44613 ; n44614
g42179 and n44603_not n44614 ; n44615
g42180 nor pi0233 n44615 ; n44616
g42181 and n2604 n16479 ; n44617
g42182 and n44560 n44606_not ; n44618
g42183 and n44570 n44611 ; n44619
g42184 and pi1147 n44617_not ; n44620
g42185 and n44618_not n44620 ; n44621
g42186 and n44619_not n44621 ; n44622
g42187 and n2603_not n44560 ; n44623
g42188 nor n44608 n44623 ; n44624
g42189 nor pi1147 n44624 ; n44625
g42190 and n44614_not n44625 ; n44626
g42191 nor n44622 n44626 ; n44627
g42192 and pi0233 n44627_not ; n44628
g42193 or n44616 n44628 ; po0467
g42194 nor pi0055 pi0311 ; n44630
g42195 nor n44558 n44630 ; n44631
g42196 and pi0311_not n44558 ; n44632
g42197 nor n44631 n44632 ; po0468
g42198 and pi0312 n44550_not ; n44634
g42199 nor n44551 n44634 ; n44635
g42200 nor pi0055 n44635 ; po0469
g42201 nor n10388 n13446 ; n44637
g42202 and po0740 n13453_not ; n44638
g42203 and n10166 n44638_not ; n44639
g42204 nand n44637_not n44639 ; po0634
g42205 and pi0954_not po0634 ; n44641
g42206 and pi0313 pi0954 ; n44642
g42207 nor n44641 n44642 ; po0470
g42208 and n6323 n8880 ; n44644
g42209 and n14440 n44644_not ; n44645
g42210 and pi0039 n15297_not ; n44646
g42211 nor pi0039 n14514 ; n44647
g42212 and n2608 n44646_not ; n44648
g42213 and n44647_not n44648 ; n44649
g42214 nor n15333 n44649 ; n44650
g42215 and n2534 n10163 ; n44651
g42216 and n44650_not n44651 ; n44652
g42217 nor n44645 n44652 ; n44653
g42218 and n14432 n14433 ; n44654
g42219 and n44653_not n44654 ; po0471
g42220 and pi0340_not n44454 ; n44656
g42221 and po1038_not n44656 ; n44657
g42222 and pi0315 n44657_not ; n44658
g42223 and pi1080 n44657 ; n44659
g42224 or n44658 n44659 ; po0472
g42225 and pi0316 n44657_not ; n44661
g42226 and pi1047 n44657 ; n44662
g42227 or n44661 n44662 ; po0473
g42228 and pi0330_not po0637 ; n44664
g42229 and pi0317 n44664_not ; n44665
g42230 and pi1078 n44664 ; n44666
g42231 or n44665 n44666 ; po0474
g42232 and pi0341_not n44454 ; n44668
g42233 and po1038_not n44668 ; n44669
g42234 and pi0318 n44669_not ; n44670
g42235 and pi1074 n44669 ; n44671
g42236 or n44670 n44671 ; po0475
g42237 and pi0319 n44669_not ; n44673
g42238 and pi1072 n44669 ; n44674
g42239 or n44673 n44674 ; po0476
g42240 and pi0320 n44657_not ; n44676
g42241 and pi1048 n44657 ; n44677
g42242 or n44676 n44677 ; po0477
g42243 and pi0321 n44657_not ; n44679
g42244 and pi1058 n44657 ; n44680
g42245 or n44679 n44680 ; po0478
g42246 and pi0322 n44657_not ; n44682
g42247 and pi1051 n44657 ; n44683
g42248 or n44682 n44683 ; po0479
g42249 and pi0323 n44657_not ; n44685
g42250 and pi1065 n44657 ; n44686
g42251 or n44685 n44686 ; po0480
g42252 and pi0324 n44669_not ; n44688
g42253 and pi1086 n44669 ; n44689
g42254 or n44688 n44689 ; po0481
g42255 and pi0325 n44669_not ; n44691
g42256 and pi1063 n44669 ; n44692
g42257 or n44691 n44692 ; po0482
g42258 and pi0326 n44669_not ; n44694
g42259 and pi1057 n44669 ; n44695
g42260 or n44694 n44695 ; po0483
g42261 and pi0327 n44657_not ; n44697
g42262 and pi1040 n44657 ; n44698
g42263 or n44697 n44698 ; po0484
g42264 and pi0328 n44669_not ; n44700
g42265 and pi1058 n44669 ; n44701
g42266 or n44700 n44701 ; po0485
g42267 and pi0329 n44669_not ; n44703
g42268 and pi1043 n44669 ; n44704
g42269 or n44703 n44704 ; po0486
g42270 and pi1092 n2930_not ; n44706
g42271 and po1038 n44706 ; n44707
g42272 and pi0330_not n44707 ; n44708
g42273 and po1038_not n44706 ; n44709
g42274 nor pi0330 n44454 ; n44710
g42275 nor n44656 n44710 ; n44711
g42276 and n44709 n44711_not ; n44712
g42277 or n44708 n44712 ; po0487
g42278 and pi0331_not n44707 ; n44714
g42279 nor pi0331 n44454 ; n44715
g42280 nor n44668 n44715 ; n44716
g42281 and n44709 n44716_not ; n44717
g42282 or n44714 n44717 ; po0488
g42283 and n11002 n13166 ; n44719
g42284 nor n11002 n13102 ; n44720
g42285 and n7445 n44720_not ; n44721
g42286 nor pi0070 n44721 ; n44722
g42287 and pi0332 n9117 ; n44723
g42288 and n44722_not n44723 ; n44724
g42289 nor n44719 n44724 ; n44725
g42290 nor pi0039 n44725 ; n44726
g42291 and pi0039 n10368 ; n44727
g42292 nor pi0038 n44727 ; n44728
g42293 and n44726_not n44728 ; n44729
g42294 and n38269 n44729_not ; po0489
g42295 and pi0333 n44669_not ; n44731
g42296 and pi1040 n44669 ; n44732
g42297 or n44731 n44732 ; po0490
g42298 and pi0334 n44669_not ; n44734
g42299 and pi1065 n44669 ; n44735
g42300 or n44734 n44735 ; po0491
g42301 and pi0335 n44669_not ; n44737
g42302 and pi1069 n44669 ; n44738
g42303 or n44737 n44738 ; po0492
g42304 and pi0336 n44664_not ; n44740
g42305 and pi1070 n44664 ; n44741
g42306 or n44740 n44741 ; po0493
g42307 and pi0337 n44664_not ; n44743
g42308 and pi1044 n44664 ; n44744
g42309 or n44743 n44744 ; po0494
g42310 and pi0338 n44664_not ; n44746
g42311 and pi1072 n44664 ; n44747
g42312 or n44746 n44747 ; po0495
g42313 and pi0339 n44664_not ; n44749
g42314 and pi1086 n44664 ; n44750
g42315 or n44749 n44750 ; po0496
g42316 and pi0340 n44707 ; n44752
g42317 nor pi0340 n44454 ; n44753
g42318 and pi0331_not n44454 ; n44754
g42319 and n44709 n44753_not ; n44755
g42320 and n44754_not n44755 ; n44756
g42321 nor n44752 n44756 ; po0497
g42322 nor pi0341 po0637 ; n44758
g42323 nor n44664 n44758 ; n44759
g42324 and n44706 n44759_not ; po0498
g42325 and pi0342 n44657_not ; n44761
g42326 and pi1049 n44657 ; n44762
g42327 or n44761 n44762 ; po0499
g42328 and pi0343 n44657_not ; n44764
g42329 and pi1062 n44657 ; n44765
g42330 or n44764 n44765 ; po0500
g42331 and pi0344 n44657_not ; n44767
g42332 and pi1069 n44657 ; n44768
g42333 or n44767 n44768 ; po0501
g42334 and pi0345 n44657_not ; n44770
g42335 and pi1039 n44657 ; n44771
g42336 or n44770 n44771 ; po0502
g42337 and pi0346 n44657_not ; n44773
g42338 and pi1067 n44657 ; n44774
g42339 or n44773 n44774 ; po0503
g42340 and pi0347 n44657_not ; n44776
g42341 and pi1055 n44657 ; n44777
g42342 or n44776 n44777 ; po0504
g42343 and pi0348 n44657_not ; n44779
g42344 and pi1087 n44657 ; n44780
g42345 or n44779 n44780 ; po0505
g42346 and pi0349 n44657_not ; n44782
g42347 and pi1043 n44657 ; n44783
g42348 or n44782 n44783 ; po0506
g42349 and pi0350 n44657_not ; n44785
g42350 and pi1035 n44657 ; n44786
g42351 or n44785 n44786 ; po0507
g42352 and pi0351 n44657_not ; n44788
g42353 and pi1079 n44657 ; n44789
g42354 or n44788 n44789 ; po0508
g42355 and pi0352 n44657_not ; n44791
g42356 and pi1078 n44657 ; n44792
g42357 or n44791 n44792 ; po0509
g42358 and pi0353 n44657_not ; n44794
g42359 and pi1063 n44657 ; n44795
g42360 or n44794 n44795 ; po0510
g42361 and pi0354 n44657_not ; n44797
g42362 and pi1045 n44657 ; n44798
g42363 or n44797 n44798 ; po0511
g42364 and pi0355 n44657_not ; n44800
g42365 and pi1084 n44657 ; n44801
g42366 or n44800 n44801 ; po0512
g42367 and pi0356 n44657_not ; n44803
g42368 and pi1081 n44657 ; n44804
g42369 or n44803 n44804 ; po0513
g42370 and pi0357 n44657_not ; n44806
g42371 and pi1076 n44657 ; n44807
g42372 or n44806 n44807 ; po0514
g42373 and pi0358 n44657_not ; n44809
g42374 and pi1071 n44657 ; n44810
g42375 or n44809 n44810 ; po0515
g42376 and pi0359 n44657_not ; n44812
g42377 and pi1068 n44657 ; n44813
g42378 or n44812 n44813 ; po0516
g42379 and pi0360 n44657_not ; n44815
g42380 and pi1042 n44657 ; n44816
g42381 or n44815 n44816 ; po0517
g42382 and pi0361 n44657_not ; n44818
g42383 and pi1059 n44657 ; n44819
g42384 or n44818 n44819 ; po0518
g42385 and pi0362 n44657_not ; n44821
g42386 and pi1070 n44657 ; n44822
g42387 or n44821 n44822 ; po0519
g42388 and pi0363 n44664_not ; n44824
g42389 and pi1049 n44664 ; n44825
g42390 or n44824 n44825 ; po0520
g42391 and pi0364 n44664_not ; n44827
g42392 and pi1062 n44664 ; n44828
g42393 or n44827 n44828 ; po0521
g42394 and pi0365 n44664_not ; n44830
g42395 and pi1065 n44664 ; n44831
g42396 or n44830 n44831 ; po0522
g42397 and pi0366 n44664_not ; n44833
g42398 and pi1069 n44664 ; n44834
g42399 or n44833 n44834 ; po0523
g42400 and pi0367 n44664_not ; n44836
g42401 and pi1039 n44664 ; n44837
g42402 or n44836 n44837 ; po0524
g42403 and pi0368 n44664_not ; n44839
g42404 and pi1067 n44664 ; n44840
g42405 or n44839 n44840 ; po0525
g42406 and pi0369 n44664_not ; n44842
g42407 and pi1080 n44664 ; n44843
g42408 or n44842 n44843 ; po0526
g42409 and pi0370 n44664_not ; n44845
g42410 and pi1055 n44664 ; n44846
g42411 or n44845 n44846 ; po0527
g42412 and pi0371 n44664_not ; n44848
g42413 and pi1051 n44664 ; n44849
g42414 or n44848 n44849 ; po0528
g42415 and pi0372 n44664_not ; n44851
g42416 and pi1048 n44664 ; n44852
g42417 or n44851 n44852 ; po0529
g42418 and pi0373 n44664_not ; n44854
g42419 and pi1087 n44664 ; n44855
g42420 or n44854 n44855 ; po0530
g42421 and pi0374 n44664_not ; n44857
g42422 and pi1035 n44664 ; n44858
g42423 or n44857 n44858 ; po0531
g42424 and pi0375 n44664_not ; n44860
g42425 and pi1047 n44664 ; n44861
g42426 or n44860 n44861 ; po0532
g42427 and pi0376 n44664_not ; n44863
g42428 and pi1079 n44664 ; n44864
g42429 or n44863 n44864 ; po0533
g42430 and pi0377 n44664_not ; n44866
g42431 and pi1074 n44664 ; n44867
g42432 or n44866 n44867 ; po0534
g42433 and pi0378 n44664_not ; n44869
g42434 and pi1063 n44664 ; n44870
g42435 or n44869 n44870 ; po0535
g42436 and pi0379 n44664_not ; n44872
g42437 and pi1045 n44664 ; n44873
g42438 or n44872 n44873 ; po0536
g42439 and pi0380 n44664_not ; n44875
g42440 and pi1084 n44664 ; n44876
g42441 or n44875 n44876 ; po0537
g42442 and pi0381 n44664_not ; n44878
g42443 and pi1081 n44664 ; n44879
g42444 or n44878 n44879 ; po0538
g42445 and pi0382 n44664_not ; n44881
g42446 and pi1076 n44664 ; n44882
g42447 or n44881 n44882 ; po0539
g42448 and pi0383 n44664_not ; n44884
g42449 and pi1071 n44664 ; n44885
g42450 or n44884 n44885 ; po0540
g42451 and pi0384 n44664_not ; n44887
g42452 and pi1068 n44664 ; n44888
g42453 or n44887 n44888 ; po0541
g42454 and pi0385 n44664_not ; n44890
g42455 and pi1042 n44664 ; n44891
g42456 or n44890 n44891 ; po0542
g42457 and pi0386 n44664_not ; n44893
g42458 and pi1059 n44664 ; n44894
g42459 or n44893 n44894 ; po0543
g42460 and pi0387 n44664_not ; n44896
g42461 and pi1053 n44664 ; n44897
g42462 or n44896 n44897 ; po0544
g42463 and pi0388 n44664_not ; n44899
g42464 and pi1037 n44664 ; n44900
g42465 or n44899 n44900 ; po0545
g42466 and pi0389 n44664_not ; n44902
g42467 and pi1036 n44664 ; n44903
g42468 or n44902 n44903 ; po0546
g42469 and pi0390 n44669_not ; n44905
g42470 and pi1049 n44669 ; n44906
g42471 or n44905 n44906 ; po0547
g42472 and pi0391 n44669_not ; n44908
g42473 and pi1062 n44669 ; n44909
g42474 or n44908 n44909 ; po0548
g42475 and pi0392 n44669_not ; n44911
g42476 and pi1039 n44669 ; n44912
g42477 or n44911 n44912 ; po0549
g42478 and pi0393 n44669_not ; n44914
g42479 and pi1067 n44669 ; n44915
g42480 or n44914 n44915 ; po0550
g42481 and pi0394 n44669_not ; n44917
g42482 and pi1080 n44669 ; n44918
g42483 or n44917 n44918 ; po0551
g42484 and pi0395 n44669_not ; n44920
g42485 and pi1055 n44669 ; n44921
g42486 or n44920 n44921 ; po0552
g42487 and pi0396 n44669_not ; n44923
g42488 and pi1051 n44669 ; n44924
g42489 or n44923 n44924 ; po0553
g42490 and pi0397 n44669_not ; n44926
g42491 and pi1048 n44669 ; n44927
g42492 or n44926 n44927 ; po0554
g42493 and pi0398 n44669_not ; n44929
g42494 and pi1087 n44669 ; n44930
g42495 or n44929 n44930 ; po0555
g42496 and pi0399 n44669_not ; n44932
g42497 and pi1047 n44669 ; n44933
g42498 or n44932 n44933 ; po0556
g42499 and pi0400 n44669_not ; n44935
g42500 and pi1035 n44669 ; n44936
g42501 or n44935 n44936 ; po0557
g42502 and pi0401 n44669_not ; n44938
g42503 and pi1079 n44669 ; n44939
g42504 or n44938 n44939 ; po0558
g42505 and pi0402 n44669_not ; n44941
g42506 and pi1078 n44669 ; n44942
g42507 or n44941 n44942 ; po0559
g42508 and pi0403 n44669_not ; n44944
g42509 and pi1045 n44669 ; n44945
g42510 or n44944 n44945 ; po0560
g42511 and pi0404 n44669_not ; n44947
g42512 and pi1084 n44669 ; n44948
g42513 or n44947 n44948 ; po0561
g42514 and pi0405 n44669_not ; n44950
g42515 and pi1081 n44669 ; n44951
g42516 or n44950 n44951 ; po0562
g42517 and pi0406 n44669_not ; n44953
g42518 and pi1076 n44669 ; n44954
g42519 or n44953 n44954 ; po0563
g42520 and pi0407 n44669_not ; n44956
g42521 and pi1071 n44669 ; n44957
g42522 or n44956 n44957 ; po0564
g42523 and pi0408 n44669_not ; n44959
g42524 and pi1068 n44669 ; n44960
g42525 or n44959 n44960 ; po0565
g42526 and pi0409 n44669_not ; n44962
g42527 and pi1042 n44669 ; n44963
g42528 or n44962 n44963 ; po0566
g42529 and pi0410 n44669_not ; n44965
g42530 and pi1059 n44669 ; n44966
g42531 or n44965 n44966 ; po0567
g42532 and pi0411 n44669_not ; n44968
g42533 and pi1053 n44669 ; n44969
g42534 or n44968 n44969 ; po0568
g42535 and pi0412 n44669_not ; n44971
g42536 and pi1037 n44669 ; n44972
g42537 or n44971 n44972 ; po0569
g42538 and pi0413 n44669_not ; n44974
g42539 and pi1036 n44669 ; n44975
g42540 or n44974 n44975 ; po0570
g42541 and po1038_not n44754 ; n44977
g42542 and pi0414 n44977_not ; n44978
g42543 and pi1049 n44977 ; n44979
g42544 or n44978 n44979 ; po0571
g42545 and pi0415 n44977_not ; n44981
g42546 and pi1062 n44977 ; n44982
g42547 or n44981 n44982 ; po0572
g42548 and pi0416 n44977_not ; n44984
g42549 and pi1069 n44977 ; n44985
g42550 or n44984 n44985 ; po0573
g42551 and pi0417 n44977_not ; n44987
g42552 and pi1039 n44977 ; n44988
g42553 or n44987 n44988 ; po0574
g42554 and pi0418 n44977_not ; n44990
g42555 and pi1067 n44977 ; n44991
g42556 or n44990 n44991 ; po0575
g42557 and pi0419 n44977_not ; n44993
g42558 and pi1080 n44977 ; n44994
g42559 or n44993 n44994 ; po0576
g42560 and pi0420 n44977_not ; n44996
g42561 and pi1055 n44977 ; n44997
g42562 or n44996 n44997 ; po0577
g42563 and pi0421 n44977_not ; n44999
g42564 and pi1051 n44977 ; n45000
g42565 or n44999 n45000 ; po0578
g42566 and pi0422 n44977_not ; n45002
g42567 and pi1048 n44977 ; n45003
g42568 or n45002 n45003 ; po0579
g42569 and pi0423 n44977_not ; n45005
g42570 and pi1087 n44977 ; n45006
g42571 or n45005 n45006 ; po0580
g42572 and pi0424 n44977_not ; n45008
g42573 and pi1047 n44977 ; n45009
g42574 or n45008 n45009 ; po0581
g42575 and pi0425 n44977_not ; n45011
g42576 and pi1035 n44977 ; n45012
g42577 or n45011 n45012 ; po0582
g42578 and pi0426 n44977_not ; n45014
g42579 and pi1079 n44977 ; n45015
g42580 or n45014 n45015 ; po0583
g42581 and pi0427 n44977_not ; n45017
g42582 and pi1078 n44977 ; n45018
g42583 or n45017 n45018 ; po0584
g42584 and pi0428 n44977_not ; n45020
g42585 and pi1045 n44977 ; n45021
g42586 or n45020 n45021 ; po0585
g42587 and pi0429 n44977_not ; n45023
g42588 and pi1084 n44977 ; n45024
g42589 or n45023 n45024 ; po0586
g42590 and pi0430 n44977_not ; n45026
g42591 and pi1076 n44977 ; n45027
g42592 or n45026 n45027 ; po0587
g42593 and pi0431 n44977_not ; n45029
g42594 and pi1071 n44977 ; n45030
g42595 or n45029 n45030 ; po0588
g42596 and pi0432 n44977_not ; n45032
g42597 and pi1068 n44977 ; n45033
g42598 or n45032 n45033 ; po0589
g42599 and pi0433 n44977_not ; n45035
g42600 and pi1042 n44977 ; n45036
g42601 or n45035 n45036 ; po0590
g42602 and pi0434 n44977_not ; n45038
g42603 and pi1059 n44977 ; n45039
g42604 or n45038 n45039 ; po0591
g42605 and pi0435 n44977_not ; n45041
g42606 and pi1053 n44977 ; n45042
g42607 or n45041 n45042 ; po0592
g42608 and pi0436 n44977_not ; n45044
g42609 and pi1037 n44977 ; n45045
g42610 or n45044 n45045 ; po0593
g42611 and pi0437 n44977_not ; n45047
g42612 and pi1070 n44977 ; n45048
g42613 or n45047 n45048 ; po0594
g42614 and pi0438 n44977_not ; n45050
g42615 and pi1036 n44977 ; n45051
g42616 or n45050 n45051 ; po0595
g42617 and pi0439 n44664_not ; n45053
g42618 and pi1057 n44664 ; n45054
g42619 or n45053 n45054 ; po0596
g42620 and pi0440 n44664_not ; n45056
g42621 and pi1043 n44664 ; n45057
g42622 or n45056 n45057 ; po0597
g42623 and pi0441 n44657_not ; n45059
g42624 and pi1044 n44657 ; n45060
g42625 or n45059 n45060 ; po0598
g42626 and pi0442 n44664_not ; n45062
g42627 and pi1058 n44664 ; n45063
g42628 or n45062 n45063 ; po0599
g42629 and pi0443 n44977_not ; n45065
g42630 and pi1044 n44977 ; n45066
g42631 or n45065 n45066 ; po0600
g42632 and pi0444 n44977_not ; n45068
g42633 and pi1072 n44977 ; n45069
g42634 or n45068 n45069 ; po0601
g42635 and pi0445 n44977_not ; n45071
g42636 and pi1081 n44977 ; n45072
g42637 or n45071 n45072 ; po0602
g42638 and pi0446 n44977_not ; n45074
g42639 and pi1086 n44977 ; n45075
g42640 or n45074 n45075 ; po0603
g42641 and pi0447 n44664_not ; n45077
g42642 and pi1040 n44664 ; n45078
g42643 or n45077 n45078 ; po0604
g42644 and pi0448 n44977_not ; n45080
g42645 and pi1074 n44977 ; n45081
g42646 or n45080 n45081 ; po0605
g42647 and pi0449 n44977_not ; n45083
g42648 and pi1057 n44977 ; n45084
g42649 or n45083 n45084 ; po0606
g42650 and pi0450 n44657_not ; n45086
g42651 and pi1036 n44657 ; n45087
g42652 or n45086 n45087 ; po0607
g42653 and pi0451 n44977_not ; n45089
g42654 and pi1063 n44977 ; n45090
g42655 or n45089 n45090 ; po0608
g42656 and pi0452 n44657_not ; n45092
g42657 and pi1053 n44657 ; n45093
g42658 or n45092 n45093 ; po0609
g42659 and pi0453 n44977_not ; n45095
g42660 and pi1040 n44977 ; n45096
g42661 or n45095 n45096 ; po0610
g42662 and pi0454 n44977_not ; n45098
g42663 and pi1043 n44977 ; n45099
g42664 or n45098 n45099 ; po0611
g42665 and pi0455 n44657_not ; n45101
g42666 and pi1037 n44657 ; n45102
g42667 or n45101 n45102 ; po0612
g42668 and pi0456 n44669_not ; n45104
g42669 and pi1044 n44669 ; n45105
g42670 or n45104 n45105 ; po0613
g42671 and pi0594 pi0600 ; n45107
g42672 and pi0597 n45107 ; n45108
g42673 and pi0601 n45108 ; n45109
g42674 nor pi0804 pi0810 ; n45110
g42675 and pi0595_not n45110 ; n45111
g42676 and pi0599_not pi0810 ; n45112
g42677 and pi0596 n45112_not ; n45113
g42678 and pi0804 n45113_not ; n45114
g42679 and pi0595 pi0815 ; n45115
g42680 and n45114_not n45115 ; n45116
g42681 nor n45111 n45116 ; n45117
g42682 and n45109 n45117_not ; n45118
g42683 and pi0600 pi0810_not ; n45119
g42684 and pi0804 n45119_not ; n45120
g42685 nor pi0601 n45110 ; n45121
g42686 nor pi0815 n45120 ; n45122
g42687 and n45121_not n45122 ; n45123
g42688 nor n45118 n45123 ; n45124
g42689 and pi0605 n45124_not ; n45125
g42690 and pi0990 n45107 ; n45126
g42691 and pi0815_not n45120 ; n45127
g42692 and n45126 n45127 ; n45128
g42693 nor n45125 n45128 ; n45129
g42694 and pi0821 n45129_not ; po0614
g42695 and pi0458 n44657_not ; n45131
g42696 and pi1072 n44657 ; n45132
g42697 or n45131 n45132 ; po0615
g42698 and pi0459 n44977_not ; n45134
g42699 and pi1058 n44977 ; n45135
g42700 or n45134 n45135 ; po0616
g42701 and pi0460 n44657_not ; n45137
g42702 and pi1086 n44657 ; n45138
g42703 or n45137 n45138 ; po0617
g42704 and pi0461 n44657_not ; n45140
g42705 and pi1057 n44657 ; n45141
g42706 or n45140 n45141 ; po0618
g42707 and pi0462 n44657_not ; n45143
g42708 and pi1074 n44657 ; n45144
g42709 or n45143 n45144 ; po0619
g42710 and pi0463 n44669_not ; n45146
g42711 and pi1070 n44669 ; n45147
g42712 or n45146 n45147 ; po0620
g42713 and pi0464 n44977_not ; n45149
g42714 and pi1065 n44977 ; n45150
g42715 or n45149 n45150 ; po0621
g42716 and pi0299_not n44561 ; n45152
g42717 nor n11423 n45152 ; n45153
g42718 nor n11396 n11399 ; n45154
g42719 nor pi0243 n45154 ; n45155
g42720 and pi0243_not pi1157 ; n45156
g42721 nor n45153 n45156 ; n45157
g42722 and n45155_not n45157 ; n45158
g42723 nor n3471 n11424 ; n45159
g42724 and pi0926 n45156 ; n45160
g42725 and n45159_not n45160 ; n45161
g42726 nor n5836 n5854 ; n45162
g42727 and pi0926 n45162_not ; n45163
g42728 and pi1157 n45162 ; n45164
g42729 nor n45155 n45163 ; n45165
g42730 and n45164_not n45165 ; n45166
g42731 nor n45158 n45161 ; n45167
g42732 and n45166_not n45167 ; n45168
g42733 nor po1038 n45168 ; n45169
g42734 and pi0243_not n44573 ; n45170
g42735 and pi0926 n44575 ; n45171
g42736 and pi1157 n5780_not ; n45172
g42737 and po1038 n45170_not ; n45173
g42738 nor n45171 n45172 ; n45174
g42739 and n45173 n45174 ; n45175
g42740 nor n45169 n45175 ; po0622
g42741 and po1038 n44573_not ; n45177
g42742 and po1038_not n45154 ; n45178
g42743 nor n45177 n45178 ; n45179
g42744 nor pi0943 n45179 ; n45180
g42745 and n44571_not n45180 ; n45181
g42746 and pi0943 n44624 ; n45182
g42747 nor n45180 n45182 ; n45183
g42748 nor pi1151 n45183 ; n45184
g42749 nor po1038 n45153 ; n45185
g42750 and n2526 po1038 ; n45186
g42751 nor n45185 n45186 ; n45187
g42752 nor pi0275 n45187 ; n45188
g42753 nor n44567 n44617 ; n45189
g42754 and pi0943 pi1151 ; n45190
g42755 and n45189_not n45190 ; n45191
g42756 nor n45181 n45188 ; n45192
g42757 and n45191_not n45192 ; n45193
g42758 and n45184_not n45193 ; po0623
g42759 and pi0040 pi0287_not ; n45195
g42760 and n42346 n45195 ; n45196
g42761 and po0950 n45196 ; n45197
g42762 nor n10165 n45197 ; n45198
g42763 nor pi0102 n13381 ; n45199
g42764 and n8897 n10162 ; n45200
g42765 and n16847 n45200 ; n45201
g42766 and n45199_not n45201 ; n45202
g42767 and n16845 n45202 ; n45203
g42768 and n45196 n45203_not ; n45204
g42769 and n45196_not n45203 ; n45205
g42770 nor n45204 n45205 ; n45206
g42771 and n7490 n45206_not ; n45207
g42772 nor n6277 n45206 ; n45208
g42773 and n6277 n45203 ; n45209
g42774 nor n45208 n45209 ; n45210
g42775 nor n7490 n45210 ; n45211
g42776 and pi1091 n45207_not ; n45212
g42777 and n45211_not n45212 ; n45213
g42778 nor pi1093 n45210 ; n45214
g42779 nor n7417 n45206 ; n45215
g42780 and n7417 n45203 ; n45216
g42781 nor n45215 n45216 ; n45217
g42782 and pi1093 n45217_not ; n45218
g42783 nor pi1091 n45214 ; n45219
g42784 and n45218_not n45219 ; n45220
g42785 nor n45213 n45220 ; n45221
g42786 and n2610 n44644 ; n45222
g42787 and n45221_not n45222 ; n45223
g42788 nor n45198 n45223 ; po0624
g42789 and n10200 n11337 ; n45225
g42790 and pi0038 pi0039_not ; n45226
g42791 and n10197 n45226 ; n45227
g42792 and n8962 n45227 ; n45228
g42793 and pi0468 n45228_not ; n45229
g42794 or n45225 n45229 ; po0625
g42795 nor pi0263 n45154 ; n45231
g42796 and pi0263_not pi1156 ; n45232
g42797 nor n45153 n45232 ; n45233
g42798 and n45231_not n45233 ; n45234
g42799 and pi0942 n45232 ; n45235
g42800 and n45159_not n45235 ; n45236
g42801 and pi0942 n45162_not ; n45237
g42802 and pi1156 n45162 ; n45238
g42803 nor n45231 n45237 ; n45239
g42804 and n45238_not n45239 ; n45240
g42805 nor n45234 n45236 ; n45241
g42806 and n45240_not n45241 ; n45242
g42807 nor po1038 n45242 ; n45243
g42808 and pi1156 n5780_not ; n45244
g42809 and pi0942 n44575 ; n45245
g42810 and pi0263_not n44573 ; n45246
g42811 and po1038 n45246_not ; n45247
g42812 nor n45244 n45245 ; n45248
g42813 and n45247 n45248 ; n45249
g42814 nor n45243 n45249 ; po0626
g42815 and pi0267 n45154_not ; n45251
g42816 and pi0267 pi1155 ; n45252
g42817 nor n45153 n45252 ; n45253
g42818 and n45251_not n45253 ; n45254
g42819 and pi0925 n45252 ; n45255
g42820 and n45159_not n45255 ; n45256
g42821 and pi0925 n45162_not ; n45257
g42822 and pi1155 n45162 ; n45258
g42823 nor n45251 n45257 ; n45259
g42824 and n45258_not n45259 ; n45260
g42825 nor n45254 n45256 ; n45261
g42826 and n45260_not n45261 ; n45262
g42827 nor po1038 n45262 ; n45263
g42828 and pi1155 n5780_not ; n45264
g42829 and pi0925 n44575 ; n45265
g42830 and pi0267 n44573 ; n45266
g42831 and po1038 n45266_not ; n45267
g42832 nor n45264 n45265 ; n45268
g42833 and n45267 n45268 ; n45269
g42834 nor n45263 n45269 ; po0627
g42835 and pi0253 n45154_not ; n45271
g42836 and pi0253 pi1153 ; n45272
g42837 nor n45153 n45272 ; n45273
g42838 and n45271_not n45273 ; n45274
g42839 and pi0941 n45272 ; n45275
g42840 and n45159_not n45275 ; n45276
g42841 and pi0941 n45162_not ; n45277
g42842 and pi1153 n45162 ; n45278
g42843 nor n45271 n45277 ; n45279
g42844 and n45278_not n45279 ; n45280
g42845 nor n45274 n45276 ; n45281
g42846 and n45280_not n45281 ; n45282
g42847 nor po1038 n45282 ; n45283
g42848 and pi1153 n5780_not ; n45284
g42849 and pi0941 n44575 ; n45285
g42850 and pi0253 n44573 ; n45286
g42851 and po1038 n45286_not ; n45287
g42852 nor n45284 n45285 ; n45288
g42853 and n45287 n45288 ; n45289
g42854 nor n45283 n45289 ; po0628
g42855 and pi0254 n45154_not ; n45291
g42856 and pi0254 pi1154 ; n45292
g42857 nor n45153 n45292 ; n45293
g42858 and n45291_not n45293 ; n45294
g42859 and pi0923 n45292 ; n45295
g42860 and n45159_not n45295 ; n45296
g42861 and pi0923 n45162_not ; n45297
g42862 and pi1154 n45162 ; n45298
g42863 nor n45291 n45297 ; n45299
g42864 and n45298_not n45299 ; n45300
g42865 nor n45294 n45296 ; n45301
g42866 and n45300_not n45301 ; n45302
g42867 nor po1038 n45302 ; n45303
g42868 and pi1154 n5780_not ; n45304
g42869 and pi0923 n44575 ; n45305
g42870 and pi0254 n44573 ; n45306
g42871 and po1038 n45306_not ; n45307
g42872 nor n45304 n45305 ; n45308
g42873 and n45307 n45308 ; n45309
g42874 nor n45303 n45309 ; po0629
g42875 nor pi0922 n45179 ; n45311
g42876 and n44571_not n45311 ; n45312
g42877 and pi0922 n44624 ; n45313
g42878 nor n45311 n45313 ; n45314
g42879 nor pi1152 n45314 ; n45315
g42880 nor pi0268 n45187 ; n45316
g42881 and pi0922 pi1152 ; n45317
g42882 and n45189_not n45317 ; n45318
g42883 nor n45312 n45316 ; n45319
g42884 and n45318_not n45319 ; n45320
g42885 and n45315_not n45320 ; po0630
g42886 nor pi0931 n45179 ; n45322
g42887 and n44571_not n45322 ; n45323
g42888 and pi0931 n44624 ; n45324
g42889 nor n45322 n45324 ; n45325
g42890 nor pi1150 n45325 ; n45326
g42891 nor pi0272 n45187 ; n45327
g42892 and pi0931 pi1150 ; n45328
g42893 and n45189_not n45328 ; n45329
g42894 nor n45323 n45327 ; n45330
g42895 and n45329_not n45330 ; n45331
g42896 and n45326_not n45331 ; po0631
g42897 nor pi0936 n45179 ; n45333
g42898 and n44571_not n45333 ; n45334
g42899 and pi0936 n44624 ; n45335
g42900 nor n45333 n45335 ; n45336
g42901 nor pi1149 n45336 ; n45337
g42902 nor pi0283 n45187 ; n45338
g42903 and pi0936 pi1149 ; n45339
g42904 and n45189_not n45339 ; n45340
g42905 nor n45334 n45338 ; n45341
g42906 and n45340_not n45341 ; n45342
g42907 and n45337_not n45342 ; po0632
g42908 and pi0071 n43509 ; n45344
g42909 and pi0071 n11448_not ; n45345
g42910 and n11448 n13052 ; n45346
g42911 and n10150 n11448_not ; n45347
g42912 and n10147 n45347 ; n45348
g42913 nor n45346 n45348 ; n45349
g42914 and n2572 n10162 ; n45350
g42915 and n45349_not n45350 ; n45351
g42916 and n13050 n45351 ; n45352
g42917 nor n45345 n45352 ; n45353
g42918 nor po1038 n45353 ; n45354
g42919 or n45344 n45354 ; po0633
g42920 and pi0071 n43791_not ; po0635
g42921 and pi0481 n34775_not ; n45357
g42922 and pi0248 n34775 ; n45358
g42923 or n45357 n45358 ; po0638
g42924 and pi0482 n34791_not ; n45360
g42925 and pi0249 n34791 ; n45361
g42926 or n45360 n45361 ; po0639
g42927 and pi0483 n34915_not ; n45363
g42928 and pi0242 n34915 ; n45364
g42929 or n45363 n45364 ; po0640
g42930 and pi0484 n34915_not ; n45366
g42931 and pi0249 n34915 ; n45367
g42932 or n45366 n45367 ; po0641
g42933 and pi0485 n36111_not ; n45369
g42934 and pi0234 n36111 ; n45370
g42935 or n45369 n45370 ; po0642
g42936 and pi0486 n36111_not ; n45372
g42937 and pi0244 n36111 ; n45373
g42938 or n45372 n45373 ; po0643
g42939 and pi0487 n34775_not ; n45375
g42940 and pi0246 n34775 ; n45376
g42941 or n45375 n45376 ; po0644
g42942 and pi0488 n34775_not ; n45378
g42943 and pi0239_not n34775 ; n45379
g42944 nor n45378 n45379 ; po0645
g42945 and pi0489 n36111_not ; n45381
g42946 and pi0242 n36111 ; n45382
g42947 or n45381 n45382 ; po0646
g42948 and pi0490 n34915_not ; n45384
g42949 and pi0241 n34915 ; n45385
g42950 or n45384 n45385 ; po0647
g42951 and pi0491 n34915_not ; n45387
g42952 and pi0238 n34915 ; n45388
g42953 or n45387 n45388 ; po0648
g42954 and pi0492 n34915_not ; n45390
g42955 and pi0240 n34915 ; n45391
g42956 or n45390 n45391 ; po0649
g42957 and pi0493 n34915_not ; n45393
g42958 and pi0244 n34915 ; n45394
g42959 or n45393 n45394 ; po0650
g42960 and pi0494 n34915_not ; n45396
g42961 and pi0239_not n34915 ; n45397
g42962 nor n45396 n45397 ; po0651
g42963 and pi0495 n34915_not ; n45399
g42964 and pi0235 n34915 ; n45400
g42965 or n45399 n45400 ; po0652
g42966 and pi0496 n34907_not ; n45402
g42967 and pi0249 n34907 ; n45403
g42968 or n45402 n45403 ; po0653
g42969 and pi0497 n34907_not ; n45405
g42970 and pi0239_not n34907 ; n45406
g42971 nor n45405 n45406 ; po0654
g42972 and pi0498 n34791_not ; n45408
g42973 and pi0238 n34791 ; n45409
g42974 or n45408 n45409 ; po0655
g42975 and pi0499 n34907_not ; n45411
g42976 and pi0246 n34907 ; n45412
g42977 or n45411 n45412 ; po0656
g42978 and pi0500 n34907_not ; n45414
g42979 and pi0241 n34907 ; n45415
g42980 or n45414 n45415 ; po0657
g42981 and pi0501 n34907_not ; n45417
g42982 and pi0248 n34907 ; n45418
g42983 or n45417 n45418 ; po0658
g42984 and pi0502 n34907_not ; n45420
g42985 and pi0247 n34907 ; n45421
g42986 or n45420 n45421 ; po0659
g42987 and pi0503 n34907_not ; n45423
g42988 and pi0245 n34907 ; n45424
g42989 or n45423 n45424 ; po0660
g42990 and pi0504 n34900_not ; n45426
g42991 and pi0242 n34900 ; n45427
g42992 or n45426 n45427 ; po0661
g42993 and n6326_not n16479 ; n45429
g42994 nor n34895 n45429 ; n45430
g42995 and pi0234_not n45430 ; n45431
g42996 and n34907 n45431 ; n45432
g42997 and pi0505 n45432_not ; n45433
g42998 and pi0234 n34899 ; n45434
g42999 and pi0505_not n34778 ; n45435
g43000 and n45434 n45435 ; n45436
g43001 or n45433 n45436 ; po0662
g43002 and pi0506 n34900_not ; n45438
g43003 and pi0241 n34900 ; n45439
g43004 or n45438 n45439 ; po0663
g43005 and pi0507 n34900_not ; n45441
g43006 and pi0238 n34900 ; n45442
g43007 or n45441 n45442 ; po0664
g43008 and pi0508 n34900_not ; n45444
g43009 and pi0247 n34900 ; n45445
g43010 or n45444 n45445 ; po0665
g43011 and pi0509 n34900_not ; n45447
g43012 and pi0245 n34900 ; n45448
g43013 or n45447 n45448 ; po0666
g43014 and pi0510 n34775_not ; n45450
g43015 and pi0242 n34775 ; n45451
g43016 or n45450 n45451 ; po0667
g43017 and n6584 po1038_not ; n45453
g43018 nor n34769 n45453 ; n45454
g43019 and pi0234_not n45454 ; n45455
g43020 and n34775 n45455_not ; n45456
g43021 and pi0511 n34775_not ; n45457
g43022 or n45456 n45457 ; po0668
g43023 and pi0512 n34775_not ; n45459
g43024 and pi0235 n34775 ; n45460
g43025 or n45459 n45460 ; po0669
g43026 and pi0513 n34775_not ; n45462
g43027 and pi0244 n34775 ; n45463
g43028 or n45462 n45463 ; po0670
g43029 and pi0514 n34775_not ; n45465
g43030 and pi0245 n34775 ; n45466
g43031 or n45465 n45466 ; po0671
g43032 and pi0515 n34775_not ; n45468
g43033 and pi0240 n34775 ; n45469
g43034 or n45468 n45469 ; po0672
g43035 and pi0516 n34775_not ; n45471
g43036 and pi0247 n34775 ; n45472
g43037 or n45471 n45472 ; po0673
g43038 and pi0517 n34775_not ; n45474
g43039 and pi0238 n34775 ; n45475
g43040 or n45474 n45475 ; po0674
g43041 and n34783 n45455 ; n45477
g43042 and pi0518 n45477_not ; n45478
g43043 and pi0234 n34774 ; n45479
g43044 and pi0518_not n34778 ; n45480
g43045 and n45479 n45480 ; n45481
g43046 or n45478 n45481 ; po0675
g43047 and pi0519 n34783_not ; n45483
g43048 and pi0239_not n34783 ; n45484
g43049 nor n45483 n45484 ; po0676
g43050 and pi0520 n34783_not ; n45486
g43051 and pi0246 n34783 ; n45487
g43052 or n45486 n45487 ; po0677
g43053 and pi0521 n34783_not ; n45489
g43054 and pi0248 n34783 ; n45490
g43055 or n45489 n45490 ; po0678
g43056 and pi0522 n34783_not ; n45492
g43057 and pi0238 n34783 ; n45493
g43058 or n45492 n45493 ; po0679
g43059 and n36139 n45455 ; n45495
g43060 and pi0523 n45495_not ; n45496
g43061 and pi0523_not n34910 ; n45497
g43062 and n45479 n45497 ; n45498
g43063 or n45496 n45498 ; po0680
g43064 and pi0524 n36139_not ; n45500
g43065 and pi0239_not n36139 ; n45501
g43066 nor n45500 n45501 ; po0681
g43067 and pi0525 n36139_not ; n45503
g43068 and pi0245 n36139 ; n45504
g43069 or n45503 n45504 ; po0682
g43070 and pi0526 n36139_not ; n45506
g43071 and pi0246 n36139 ; n45507
g43072 or n45506 n45507 ; po0683
g43073 and pi0527 n36139_not ; n45509
g43074 and pi0247 n36139 ; n45510
g43075 or n45509 n45510 ; po0684
g43076 and pi0528 n36139_not ; n45512
g43077 and pi0249 n36139 ; n45513
g43078 or n45512 n45513 ; po0685
g43079 and pi0529 n36139_not ; n45515
g43080 and pi0238 n36139 ; n45516
g43081 or n45515 n45516 ; po0686
g43082 and pi0530 n36139_not ; n45518
g43083 and pi0240 n36139 ; n45519
g43084 or n45518 n45519 ; po0687
g43085 and pi0531 n34791_not ; n45521
g43086 and pi0235 n34791 ; n45522
g43087 or n45521 n45522 ; po0688
g43088 and pi0532 n34791_not ; n45524
g43089 and pi0247 n34791 ; n45525
g43090 or n45524 n45525 ; po0689
g43091 and pi0533 n34900_not ; n45527
g43092 and pi0235 n34900 ; n45528
g43093 or n45527 n45528 ; po0690
g43094 and pi0534 n34900_not ; n45530
g43095 and pi0239_not n34900 ; n45531
g43096 nor n45530 n45531 ; po0691
g43097 and pi0535 n34900_not ; n45533
g43098 and pi0240 n34900 ; n45534
g43099 or n45533 n45534 ; po0692
g43100 and pi0536 n34900_not ; n45536
g43101 and pi0246 n34900 ; n45537
g43102 or n45536 n45537 ; po0693
g43103 and pi0537 n34900_not ; n45539
g43104 and pi0248 n34900 ; n45540
g43105 or n45539 n45540 ; po0694
g43106 and pi0538 n34900_not ; n45542
g43107 and pi0249 n34900 ; n45543
g43108 or n45542 n45543 ; po0695
g43109 and pi0539 n34907_not ; n45545
g43110 and pi0242 n34907 ; n45546
g43111 or n45545 n45546 ; po0696
g43112 and pi0540 n34907_not ; n45548
g43113 and pi0235 n34907 ; n45549
g43114 or n45548 n45549 ; po0697
g43115 and pi0541 n34907_not ; n45551
g43116 and pi0244 n34907 ; n45552
g43117 or n45551 n45552 ; po0698
g43118 and pi0542 n34907_not ; n45554
g43119 and pi0240 n34907 ; n45555
g43120 or n45554 n45555 ; po0699
g43121 and pi0543 n34907_not ; n45557
g43122 and pi0238 n34907 ; n45558
g43123 or n45557 n45558 ; po0700
g43124 and n34915 n45431 ; n45560
g43125 and pi0544 n45560_not ; n45561
g43126 and pi0544_not n34910 ; n45562
g43127 and n45434 n45562 ; n45563
g43128 or n45561 n45563 ; po0701
g43129 and pi0545 n34915_not ; n45565
g43130 and pi0245 n34915 ; n45566
g43131 or n45565 n45566 ; po0702
g43132 and pi0546 n34915_not ; n45568
g43133 and pi0246 n34915 ; n45569
g43134 or n45568 n45569 ; po0703
g43135 and pi0547 n34915_not ; n45571
g43136 and pi0247 n34915 ; n45572
g43137 or n45571 n45572 ; po0704
g43138 and pi0548 n34915_not ; n45574
g43139 and pi0248 n34915 ; n45575
g43140 or n45574 n45575 ; po0705
g43141 and pi0549 n36111_not ; n45577
g43142 and pi0235 n36111 ; n45578
g43143 or n45577 n45578 ; po0706
g43144 and pi0550 n36111_not ; n45580
g43145 and pi0239_not n36111 ; n45581
g43146 nor n45580 n45581 ; po0707
g43147 and pi0551 n36111_not ; n45583
g43148 and pi0240 n36111 ; n45584
g43149 or n45583 n45584 ; po0708
g43150 and pi0552 n36111_not ; n45586
g43151 and pi0247 n36111 ; n45587
g43152 or n45586 n45587 ; po0709
g43153 and pi0553 n36111_not ; n45589
g43154 and pi0241 n36111 ; n45590
g43155 or n45589 n45590 ; po0710
g43156 and pi0554 n36111_not ; n45592
g43157 and pi0248 n36111 ; n45593
g43158 or n45592 n45593 ; po0711
g43159 and pi0555 n36111_not ; n45595
g43160 and pi0249 n36111 ; n45596
g43161 or n45595 n45596 ; po0712
g43162 and pi0556 n34791_not ; n45598
g43163 and pi0242 n34791 ; n45599
g43164 or n45598 n45599 ; po0713
g43165 and n34900 n45431 ; n45601
g43166 and pi0557 n45601_not ; n45602
g43167 and pi0557_not n34583 ; n45603
g43168 and n45434 n45603 ; n45604
g43169 or n45602 n45604 ; po0714
g43170 and pi0558 n34900_not ; n45606
g43171 and pi0244 n34900 ; n45607
g43172 or n45606 n45607 ; po0715
g43173 and pi0559 n34775_not ; n45609
g43174 and pi0241 n34775 ; n45610
g43175 or n45609 n45610 ; po0716
g43176 and pi0560 n34791_not ; n45612
g43177 and pi0240 n34791 ; n45613
g43178 or n45612 n45613 ; po0717
g43179 and pi0561 n34783_not ; n45615
g43180 and pi0247 n34783 ; n45616
g43181 or n45615 n45616 ; po0718
g43182 and pi0562 n34791_not ; n45618
g43183 and pi0241 n34791 ; n45619
g43184 or n45618 n45619 ; po0719
g43185 and pi0563 n36111_not ; n45621
g43186 and pi0246 n36111 ; n45622
g43187 or n45621 n45622 ; po0720
g43188 and pi0564 n34791_not ; n45624
g43189 and pi0246 n34791 ; n45625
g43190 or n45624 n45625 ; po0721
g43191 and pi0565 n34791_not ; n45627
g43192 and pi0248 n34791 ; n45628
g43193 or n45627 n45628 ; po0722
g43194 and pi0566 n34791_not ; n45630
g43195 and pi0244 n34791 ; n45631
g43196 or n45630 n45631 ; po0723
g43197 and pi0567_not pi1092 ; n45633
g43198 and pi1093_not n45633 ; n45634
g43199 and pi0603 n17117_not ; n45635
g43200 and n17182 n20225_not ; n45636
g43201 and n20235_not n45636 ; n45637
g43202 and n45635 n45637 ; n45638
g43203 nor pi0789 n45634 ; n45639
g43204 and n45638_not n45639 ; n45640
g43205 and pi0619_not n45638 ; n45641
g43206 nor n45634 n45641 ; n45642
g43207 nor pi1159 n45642 ; n45643
g43208 and pi0619 n45638 ; n45644
g43209 nor n45634 n45644 ; n45645
g43210 and pi1159 n45645_not ; n45646
g43211 and pi0789 n45643_not ; n45647
g43212 and n45646_not n45647 ; n45648
g43213 nor n45640 n45648 ; n45649
g43214 and pi0680 n16826 ; n45650
g43215 and n19146_not n45650 ; n45651
g43216 nor n45634 n45651 ; n45652
g43217 and n19150 n45652_not ; n45653
g43218 and n16634_not n45648 ; n45654
g43219 and n45653 n45654_not ; n45655
g43220 nor n45649 n45655 ; n45656
g43221 and n17970 n45656_not ; n45657
g43222 and n35357 n45649 ; n45658
g43223 and n16635_not n45653 ; n45659
g43224 and pi0641 n45659 ; n45660
g43225 nor n45634 n45660 ; n45661
g43226 and n17865 n45661_not ; n45662
g43227 and pi0641_not n45659 ; n45663
g43228 nor n45634 n45663 ; n45664
g43229 and n17866 n45664_not ; n45665
g43230 nor n45662 n45665 ; n45666
g43231 and n45658_not n45666 ; n45667
g43232 and pi0788 n45667_not ; n45668
g43233 nor n45657 n45668 ; n45669
g43234 nor n20364 n45669 ; n45670
g43235 and n19151 n45652_not ; n45671
g43236 and pi0628 n45671 ; n45672
g43237 nor n45634 n45672 ; n45673
g43238 and pi1156 n45673_not ; n45674
g43239 and n17969_not n45649 ; n45675
g43240 and n17969 n45634 ; n45676
g43241 nor n45675 n45676 ; n45677
g43242 and n17854 n45677_not ; n45678
g43243 nor pi0629 n45674 ; n45679
g43244 and n45678_not n45679 ; n45680
g43245 and pi0628_not n45671 ; n45681
g43246 nor n45634 n45681 ; n45682
g43247 nor pi1156 n45682 ; n45683
g43248 and n17853 n45677_not ; n45684
g43249 and pi0629 n45683_not ; n45685
g43250 and n45684_not n45685 ; n45686
g43251 and pi0792 n45680_not ; n45687
g43252 and n45686_not n45687 ; n45688
g43253 nor n45670 n45688 ; n45689
g43254 nor pi0647 n45689 ; n45690
g43255 nor n17779 n45677 ; n45691
g43256 and n17779 n45634 ; n45692
g43257 nor n45691 n45692 ; n45693
g43258 and pi0647 n45693_not ; n45694
g43259 nor pi1157 n45694 ; n45695
g43260 and n45690_not n45695 ; n45696
g43261 and n19142_not n45671 ; n45697
g43262 and pi0647 n45697 ; n45698
g43263 and pi1157 n45634_not ; n45699
g43264 and n45698_not n45699 ; n45700
g43265 nor pi0630 n45700 ; n45701
g43266 and n45696_not n45701 ; n45702
g43267 and pi0647 n45689_not ; n45703
g43268 nor pi0647 n45693 ; n45704
g43269 and pi1157 n45704_not ; n45705
g43270 and n45703_not n45705 ; n45706
g43271 and pi0647_not n45697 ; n45707
g43272 nor pi1157 n45634 ; n45708
g43273 and n45707_not n45708 ; n45709
g43274 and pi0630 n45709_not ; n45710
g43275 and n45706_not n45710 ; n45711
g43276 nor n45702 n45711 ; n45712
g43277 and pi0787 n45712_not ; n45713
g43278 nor pi0787 n45689 ; n45714
g43279 nor n45713 n45714 ; n45715
g43280 nor pi0790 n45715 ; n45716
g43281 and n19342_not n45697 ; n45717
g43282 nor n45634 n45717 ; n45718
g43283 and pi0644 n45718_not ; n45719
g43284 nor pi0644 n45715 ; n45720
g43285 nor pi0715 n45719 ; n45721
g43286 and n45720_not n45721 ; n45722
g43287 and n17804_not n45691 ; n45723
g43288 and pi0644_not n45723 ; n45724
g43289 and pi0715 n45634_not ; n45725
g43290 and n45724_not n45725 ; n45726
g43291 nor n45722 n45726 ; n45727
g43292 nor pi1160 n45727 ; n45728
g43293 and pi0644 n45723 ; n45729
g43294 nor n45634 n45729 ; n45730
g43295 nor pi0715 n45730 ; n45731
g43296 and pi0644_not n45718 ; n45732
g43297 and pi0644 n45715 ; n45733
g43298 and pi0715 n45732_not ; n45734
g43299 and n45733_not n45734 ; n45735
g43300 and pi1160 n45731_not ; n45736
g43301 and n45735_not n45736 ; n45737
g43302 and pi0790 n45737_not ; n45738
g43303 and n45728_not n45738 ; n45739
g43304 nor n45716 n45739 ; n45740
g43305 and pi0230 n45740_not ; n45741
g43306 and pi0230_not n45633 ; n45742
g43307 or n45741 n45742 ; po0724
g43308 and pi0568 n34791_not ; n45744
g43309 and pi0245 n34791 ; n45745
g43310 or n45744 n45745 ; po0725
g43311 and pi0569 n34791_not ; n45747
g43312 and pi0239_not n34791 ; n45748
g43313 nor n45747 n45748 ; po0726
g43314 and n34791 n45455 ; n45750
g43315 and pi0570 n45750_not ; n45751
g43316 and pi0570_not n34786 ; n45752
g43317 and n45479 n45752 ; n45753
g43318 or n45751 n45753 ; po0727
g43319 and pi0571 n36139_not ; n45755
g43320 and pi0241 n36139 ; n45756
g43321 or n45755 n45756 ; po0728
g43322 and pi0572 n36139_not ; n45758
g43323 and pi0244 n36139 ; n45759
g43324 or n45758 n45759 ; po0729
g43325 and pi0573 n36139_not ; n45761
g43326 and pi0242 n36139 ; n45762
g43327 or n45761 n45762 ; po0730
g43328 and pi0574 n34783_not ; n45764
g43329 and pi0241 n34783 ; n45765
g43330 or n45764 n45765 ; po0731
g43331 and pi0575 n36139_not ; n45767
g43332 and pi0235 n36139 ; n45768
g43333 or n45767 n45768 ; po0732
g43334 and pi0576 n36139_not ; n45770
g43335 and pi0248 n36139 ; n45771
g43336 or n45770 n45771 ; po0733
g43337 and pi0577 n36111_not ; n45773
g43338 and pi0238 n36111 ; n45774
g43339 or n45773 n45774 ; po0734
g43340 and pi0578 n34783_not ; n45776
g43341 and pi0249 n34783 ; n45777
g43342 or n45776 n45777 ; po0735
g43343 and pi0579 n34775_not ; n45779
g43344 and pi0249 n34775 ; n45780
g43345 or n45779 n45780 ; po0736
g43346 and pi0580 n36111_not ; n45782
g43347 and pi0245 n36111 ; n45783
g43348 or n45782 n45783 ; po0737
g43349 and pi0581 n34783_not ; n45785
g43350 and pi0235 n34783 ; n45786
g43351 or n45785 n45786 ; po0738
g43352 and pi0582 n34783_not ; n45788
g43353 and pi0240 n34783 ; n45789
g43354 or n45788 n45789 ; po0739
g43355 and pi0584 n34783_not ; n45791
g43356 and pi0245 n34783 ; n45792
g43357 or n45791 n45792 ; po0741
g43358 and pi0585 n34783_not ; n45794
g43359 and pi0244 n34783 ; n45795
g43360 or n45794 n45795 ; po0742
g43361 and pi0586 n34783_not ; n45797
g43362 and pi0242 n34783 ; n45798
g43363 or n45797 n45798 ; po0743
g43364 and pi0230_not pi0587 ; n45800
g43365 and pi0230 n17168 ; n45801
g43366 and n20225_not n45801 ; n45802
g43367 and n35575_not n45802 ; n45803
g43368 and n20237 n45803 ; n45804
g43369 and n30797 n45804 ; n45805
g43370 or n45800 n45805 ; po0744
g43371 and pi0123_not n12373 ; n45807
g43372 nor pi0588 n45807 ; n45808
g43373 and pi0591_not n45807 ; n45809
g43374 and n44706 n45808_not ; n45810
g43375 and n45809_not n45810 ; po0745
g43376 and pi0204_not n45430 ; n45812
g43377 and pi0201_not n45454 ; n45813
g43378 and pi0233 n45812_not ; n45814
g43379 and n45813_not n45814 ; n45815
g43380 and pi0205_not n45430 ; n45816
g43381 and pi0202_not n45454 ; n45817
g43382 nor pi0233 n45816 ; n45818
g43383 and n45817_not n45818 ; n45819
g43384 nor n45815 n45819 ; n45820
g43385 and pi0237 n45820_not ; n45821
g43386 and pi0206_not n45430 ; n45822
g43387 and pi0220_not n45454 ; n45823
g43388 and pi0233 n45822_not ; n45824
g43389 and n45823_not n45824 ; n45825
g43390 and pi0218_not n45430 ; n45826
g43391 and pi0203_not n45454 ; n45827
g43392 nor pi0233 n45826 ; n45828
g43393 and n45827_not n45828 ; n45829
g43394 nor n45825 n45829 ; n45830
g43395 nor pi0237 n45830 ; n45831
g43396 nor n45821 n45831 ; po0746
g43397 and pi0588 n45807 ; n45833
g43398 and pi0590 n45807_not ; n45834
g43399 and n44706 n45833_not ; n45835
g43400 nand n45834_not n45835 ; po0747
g43401 nor pi0591 n45807 ; n45837
g43402 and pi0592_not n45807 ; n45838
g43403 and n44706 n45837_not ; n45839
g43404 and n45838_not n45839 ; po0748
g43405 nor pi0592 n45807 ; n45841
g43406 and pi0590_not n45807 ; n45842
g43407 and n44706 n45841_not ; n45843
g43408 and n45842_not n45843 ; po0749
g43409 and pi0234 n45454 ; n45845
g43410 and pi0518 n45845_not ; n45846
g43411 and pi0246 pi0520_not ; n45847
g43412 and pi0246_not pi0520 ; n45848
g43413 and pi0249 pi0578_not ; n45849
g43414 and pi0249_not pi0578 ; n45850
g43415 and pi0248 pi0521_not ; n45851
g43416 and pi0248_not pi0521 ; n45852
g43417 and pi0241 pi0574 ; n45853
g43418 nor pi0241 pi0574 ; n45854
g43419 nor n45853 n45854 ; n45855
g43420 nor pi0518 n45455 ; n45856
g43421 nor n45847 n45848 ; n45857
g43422 nor n45849 n45850 ; n45858
g43423 nor n45851 n45852 ; n45859
g43424 and n45858 n45859 ; n45860
g43425 and n45855_not n45857 ; n45861
g43426 and n45860 n45861 ; n45862
g43427 and n45846_not n45862 ; n45863
g43428 and n45856_not n45863 ; n45864
g43429 and pi0582 n45864 ; n45865
g43430 and pi0240 n45865_not ; n45866
g43431 and pi0582_not n45864 ; n45867
g43432 nor pi0240 n45867 ; n45868
g43433 nor n45866 n45868 ; n45869
g43434 and pi0239_not pi0519 ; n45870
g43435 and pi0239 pi0519_not ; n45871
g43436 nor n45870 n45871 ; n45872
g43437 and n45869 n45872_not ; n45873
g43438 and pi0242 pi0586 ; n45874
g43439 nor pi0242 pi0586 ; n45875
g43440 nor n45874 n45875 ; n45876
g43441 and n45873 n45876_not ; n45877
g43442 and pi0235 pi0581 ; n45878
g43443 nor pi0235 pi0581 ; n45879
g43444 nor n45878 n45879 ; n45880
g43445 and n45877 n45880_not ; n45881
g43446 and pi0585 n45881 ; n45882
g43447 and pi0244 n45882_not ; n45883
g43448 and pi0585_not n45881 ; n45884
g43449 nor pi0244 n45884 ; n45885
g43450 nor n45883 n45885 ; n45886
g43451 and pi0584 n45886 ; n45887
g43452 and pi0245 n45887_not ; n45888
g43453 and pi0584_not n45886 ; n45889
g43454 nor pi0245 n45889 ; n45890
g43455 nor n45888 n45890 ; n45891
g43456 nor pi0247 pi0561 ; n45892
g43457 and pi0247 pi0561 ; n45893
g43458 nor n45892 n45893 ; n45894
g43459 and n45891 n45894_not ; n45895
g43460 and pi0238 n45895 ; n45896
g43461 and pi0240 pi0542 ; n45897
g43462 nor pi0240 pi0542 ; n45898
g43463 nor n45897 n45898 ; n45899
g43464 nor pi0248 pi0501 ; n45900
g43465 and pi0248 pi0501 ; n45901
g43466 nor n45900 n45901 ; n45902
g43467 and pi0234 n45430 ; n45903
g43468 and pi0505 n45903_not ; n45904
g43469 nor pi0505 n45431 ; n45905
g43470 and pi0249 pi0496_not ; n45906
g43471 and pi0249_not pi0496 ; n45907
g43472 nor pi0246 pi0499 ; n45908
g43473 and pi0246 pi0499 ; n45909
g43474 nor n45908 n45909 ; n45910
g43475 nor n45906 n45907 ; n45911
g43476 and n45902_not n45911 ; n45912
g43477 and n45910_not n45912 ; n45913
g43478 and n45904_not n45913 ; n45914
g43479 and n45905_not n45914 ; n45915
g43480 nor pi0241 pi0500 ; n45916
g43481 and pi0241 pi0500 ; n45917
g43482 nor n45916 n45917 ; n45918
g43483 and n45915 n45918_not ; n45919
g43484 and n45899_not n45919 ; n45920
g43485 and pi0497 n45920 ; n45921
g43486 nor pi0239 n45921 ; n45922
g43487 and pi0497_not n45920 ; n45923
g43488 and pi0239 n45923_not ; n45924
g43489 nor n45922 n45924 ; n45925
g43490 and pi0539 n45925 ; n45926
g43491 and pi0242 n45926_not ; n45927
g43492 and pi0539_not n45925 ; n45928
g43493 nor pi0242 n45928 ; n45929
g43494 nor n45927 n45929 ; n45930
g43495 and pi0540 n45930 ; n45931
g43496 and pi0235 n45931_not ; n45932
g43497 and pi0540_not n45930 ; n45933
g43498 nor pi0235 n45933 ; n45934
g43499 nor n45932 n45934 ; n45935
g43500 and pi0244 pi0541 ; n45936
g43501 nor pi0244 pi0541 ; n45937
g43502 nor n45936 n45937 ; n45938
g43503 and n45935 n45938_not ; n45939
g43504 and pi0245 pi0503 ; n45940
g43505 nor pi0245 pi0503 ; n45941
g43506 nor n45940 n45941 ; n45942
g43507 and n45939 n45942_not ; n45943
g43508 and pi0502_not n45943 ; n45944
g43509 nor pi0247 n45944 ; n45945
g43510 and pi0502 n45943 ; n45946
g43511 and pi0247 n45946_not ; n45947
g43512 nor n45945 n45947 ; n45948
g43513 and pi0238_not n45948 ; n45949
g43514 and pi0522 n45896_not ; n45950
g43515 and n45949_not n45950 ; n45951
g43516 nor n45892 n45945 ; n45952
g43517 and pi0502 n45891_not ; n45953
g43518 and pi0500_not n45919 ; n45954
g43519 and n45915 n45917 ; n45955
g43520 nor n45864 n45955 ; n45956
g43521 and n45954_not n45956 ; n45957
g43522 nor pi0582 n45957 ; n45958
g43523 and pi0582 n45919 ; n45959
g43524 nor pi0240 n45959 ; n45960
g43525 and n45958_not n45960 ; n45961
g43526 nor n45866 n45961 ; n45962
g43527 nor pi0542 n45962 ; n45963
g43528 and pi0582 n45957_not ; n45964
g43529 and pi0582_not n45919 ; n45965
g43530 and pi0240 n45965_not ; n45966
g43531 and n45964_not n45966 ; n45967
g43532 nor n45868 n45967 ; n45968
g43533 and pi0542 n45968_not ; n45969
g43534 nor n45963 n45969 ; n45970
g43535 and pi0497_not n45970 ; n45971
g43536 and pi0497 n45869 ; n45972
g43537 and pi0239 n45972_not ; n45973
g43538 and n45971_not n45973 ; n45974
g43539 nor n45922 n45974 ; n45975
g43540 nor pi0519 n45975 ; n45976
g43541 and pi0497 n45970 ; n45977
g43542 and pi0497_not n45869 ; n45978
g43543 nor pi0239 n45978 ; n45979
g43544 and n45977_not n45979 ; n45980
g43545 nor n45924 n45980 ; n45981
g43546 and pi0519 n45981_not ; n45982
g43547 nor n45976 n45982 ; n45983
g43548 and pi0539_not n45983 ; n45984
g43549 and pi0539 n45873 ; n45985
g43550 nor pi0242 n45985 ; n45986
g43551 and n45984_not n45986 ; n45987
g43552 nor n45927 n45987 ; n45988
g43553 nor pi0586 n45988 ; n45989
g43554 and pi0539 n45983 ; n45990
g43555 and pi0539_not n45873 ; n45991
g43556 and pi0242 n45991_not ; n45992
g43557 and n45990_not n45992 ; n45993
g43558 nor n45929 n45993 ; n45994
g43559 and pi0586 n45994_not ; n45995
g43560 nor n45989 n45995 ; n45996
g43561 and pi0540_not n45996 ; n45997
g43562 and pi0540 n45877 ; n45998
g43563 nor pi0235 n45998 ; n45999
g43564 and n45997_not n45999 ; n46000
g43565 nor n45932 n46000 ; n46001
g43566 nor pi0581 n46001 ; n46002
g43567 and pi0540 n45996 ; n46003
g43568 and pi0540_not n45877 ; n46004
g43569 and pi0235 n46004_not ; n46005
g43570 and n46003_not n46005 ; n46006
g43571 nor n45934 n46006 ; n46007
g43572 and pi0581 n46007_not ; n46008
g43573 nor n46002 n46008 ; n46009
g43574 and pi0585_not n46009 ; n46010
g43575 and pi0585 n45935 ; n46011
g43576 nor pi0244 n46011 ; n46012
g43577 and n46010_not n46012 ; n46013
g43578 nor n45883 n46013 ; n46014
g43579 nor pi0541 n46014 ; n46015
g43580 and pi0585 n46009 ; n46016
g43581 and pi0585_not n45935 ; n46017
g43582 and pi0244 n46017_not ; n46018
g43583 and n46016_not n46018 ; n46019
g43584 nor n45885 n46019 ; n46020
g43585 and pi0541 n46020_not ; n46021
g43586 nor n46015 n46021 ; n46022
g43587 and pi0584_not n46022 ; n46023
g43588 and pi0584 n45939 ; n46024
g43589 nor pi0245 n46024 ; n46025
g43590 and n46023_not n46025 ; n46026
g43591 nor n45888 n46026 ; n46027
g43592 nor pi0503 n46027 ; n46028
g43593 and pi0584 n46022 ; n46029
g43594 and pi0584_not n45939 ; n46030
g43595 and pi0245 n46030_not ; n46031
g43596 and n46029_not n46031 ; n46032
g43597 nor n45890 n46032 ; n46033
g43598 and pi0503 n46033_not ; n46034
g43599 nor n46028 n46034 ; n46035
g43600 nor pi0502 n46035 ; n46036
g43601 nor pi0561 n45953 ; n46037
g43602 and n46036_not n46037 ; n46038
g43603 nor n45952 n46038 ; n46039
g43604 nor n45893 n45947 ; n46040
g43605 nor pi0502 n45891 ; n46041
g43606 and pi0502 n46035_not ; n46042
g43607 and pi0561 n46041_not ; n46043
g43608 and n46042_not n46043 ; n46044
g43609 nor n46040 n46044 ; n46045
g43610 nor n46039 n46045 ; n46046
g43611 and pi0238_not n46046 ; n46047
g43612 nor pi0522 n46047 ; n46048
g43613 nor pi0543 n45951 ; n46049
g43614 and n46048_not n46049 ; n46050
g43615 and pi0238_not n45895 ; n46051
g43616 and pi0238 n45948 ; n46052
g43617 nor pi0522 n46051 ; n46053
g43618 and n46052_not n46053 ; n46054
g43619 and pi0238 n46046 ; n46055
g43620 and pi0522 n46055_not ; n46056
g43621 and pi0543 n46054_not ; n46057
g43622 and n46056_not n46057 ; n46058
g43623 nor n46050 n46058 ; n46059
g43624 nor pi0233 n46059 ; n46060
g43625 and pi0246 pi0536 ; n46061
g43626 nor pi0246 pi0536 ; n46062
g43627 nor n46061 n46062 ; n46063
g43628 nor pi0557 n45431 ; n46064
g43629 and pi0557 n45903_not ; n46065
g43630 nor n46063 n46064 ; n46066
g43631 and n46065_not n46066 ; n46067
g43632 and pi0538_not n46067 ; n46068
g43633 nor pi0249 n46068 ; n46069
g43634 and pi0538 n46067 ; n46070
g43635 and pi0249 n46070_not ; n46071
g43636 nor n46069 n46071 ; n46072
g43637 and pi0537_not n46072 ; n46073
g43638 nor pi0248 n46073 ; n46074
g43639 and pi0537 n46072 ; n46075
g43640 and pi0248 n46075_not ; n46076
g43641 nor n46074 n46076 ; n46077
g43642 and pi0241 pi0506 ; n46078
g43643 nor pi0241 pi0506 ; n46079
g43644 nor n46078 n46079 ; n46080
g43645 and n46077 n46080_not ; n46081
g43646 and pi0240 pi0535 ; n46082
g43647 nor pi0240 pi0535 ; n46083
g43648 nor n46082 n46083 ; n46084
g43649 and n46081 n46084_not ; n46085
g43650 and pi0534 n46085 ; n46086
g43651 nor pi0239 n46086 ; n46087
g43652 and pi0534_not n46085 ; n46088
g43653 and pi0239 n46088_not ; n46089
g43654 nor n46087 n46089 ; n46090
g43655 and pi0504 n46090 ; n46091
g43656 and pi0242 n46091_not ; n46092
g43657 and pi0504_not n46090 ; n46093
g43658 nor pi0242 n46093 ; n46094
g43659 nor n46092 n46094 ; n46095
g43660 and pi0533 n46095 ; n46096
g43661 and pi0235 n46096_not ; n46097
g43662 and pi0533_not n46095 ; n46098
g43663 nor pi0235 n46098 ; n46099
g43664 nor n46097 n46099 ; n46100
g43665 and pi0558 n46100 ; n46101
g43666 and pi0244 n46101_not ; n46102
g43667 and pi0558_not n46100 ; n46103
g43668 nor pi0244 n46103 ; n46104
g43669 nor n46102 n46104 ; n46105
g43670 and pi0509 n46105 ; n46106
g43671 and pi0245 n46106_not ; n46107
g43672 and pi0509_not n46105 ; n46108
g43673 nor pi0245 n46108 ; n46109
g43674 nor n46107 n46109 ; n46110
g43675 and pi0508 n46110 ; n46111
g43676 and pi0247 n46111_not ; n46112
g43677 and pi0508_not n46110 ; n46113
g43678 nor pi0247 n46113 ; n46114
g43679 nor n46112 n46114 ; n46115
g43680 and pi0238_not n46115 ; n46116
g43681 and pi0248 pi0481 ; n46117
g43682 nor pi0248 pi0481 ; n46118
g43683 nor n46117 n46118 ; n46119
g43684 and pi0246 pi0487 ; n46120
g43685 nor pi0246 pi0487 ; n46121
g43686 nor n46120 n46121 ; n46122
g43687 nor pi0511 n45455 ; n46123
g43688 and pi0511 n45845_not ; n46124
g43689 nor n46122 n46123 ; n46125
g43690 and n46124_not n46125 ; n46126
g43691 nor pi0249 pi0579 ; n46127
g43692 and pi0249 pi0579 ; n46128
g43693 nor n46127 n46128 ; n46129
g43694 and n46126 n46129_not ; n46130
g43695 and n46119_not n46130 ; n46131
g43696 and pi0559 n46131 ; n46132
g43697 and pi0241 n46132_not ; n46133
g43698 and pi0559_not n46131 ; n46134
g43699 nor pi0241 n46134 ; n46135
g43700 nor n46133 n46135 ; n46136
g43701 and pi0515 n46136 ; n46137
g43702 and pi0240 n46137_not ; n46138
g43703 and pi0515_not n46136 ; n46139
g43704 nor pi0240 n46139 ; n46140
g43705 nor n46138 n46140 ; n46141
g43706 and pi0239_not pi0488 ; n46142
g43707 and pi0239 pi0488_not ; n46143
g43708 nor n46142 n46143 ; n46144
g43709 and n46141 n46144_not ; n46145
g43710 and pi0242 pi0510 ; n46146
g43711 nor pi0242 pi0510 ; n46147
g43712 nor n46146 n46147 ; n46148
g43713 and n46145 n46148_not ; n46149
g43714 and pi0235 pi0512 ; n46150
g43715 nor pi0235 pi0512 ; n46151
g43716 nor n46150 n46151 ; n46152
g43717 and n46149 n46152_not ; n46153
g43718 and pi0244 pi0513 ; n46154
g43719 nor pi0244 pi0513 ; n46155
g43720 nor n46154 n46155 ; n46156
g43721 and n46153 n46156_not ; n46157
g43722 and pi0245 pi0514 ; n46158
g43723 nor pi0245 pi0514 ; n46159
g43724 nor n46158 n46159 ; n46160
g43725 and n46157 n46160_not ; n46161
g43726 and pi0247 pi0516 ; n46162
g43727 nor pi0247 pi0516 ; n46163
g43728 nor n46162 n46163 ; n46164
g43729 and n46161 n46164_not ; n46165
g43730 and pi0238 n46165 ; n46166
g43731 and pi0517 n46166_not ; n46167
g43732 and n46116_not n46167 ; n46168
g43733 nor pi0579 n46130 ; n46169
g43734 and n46069_not n46126 ; n46170
g43735 and pi0579 n46170_not ; n46171
g43736 nor n46169 n46171 ; n46172
g43737 nor n46072 n46172 ; n46173
g43738 nor pi0537 n46173 ; n46174
g43739 and pi0537 n46130 ; n46175
g43740 nor pi0248 n46175 ; n46176
g43741 and n46174_not n46176 ; n46177
g43742 nor n46076 n46177 ; n46178
g43743 nor pi0481 n46178 ; n46179
g43744 and pi0537 n46173_not ; n46180
g43745 and pi0537_not n46130 ; n46181
g43746 and pi0248 n46181_not ; n46182
g43747 and n46180_not n46182 ; n46183
g43748 nor n46074 n46183 ; n46184
g43749 and pi0481 n46184_not ; n46185
g43750 nor n46179 n46185 ; n46186
g43751 and pi0559_not n46186 ; n46187
g43752 and pi0559 n46077 ; n46188
g43753 nor pi0241 n46188 ; n46189
g43754 and n46187_not n46189 ; n46190
g43755 nor n46133 n46190 ; n46191
g43756 nor pi0506 n46191 ; n46192
g43757 and pi0559 n46186 ; n46193
g43758 and pi0559_not n46077 ; n46194
g43759 and pi0241 n46194_not ; n46195
g43760 and n46193_not n46195 ; n46196
g43761 nor n46135 n46196 ; n46197
g43762 and pi0506 n46197_not ; n46198
g43763 nor n46192 n46198 ; n46199
g43764 and pi0515_not n46199 ; n46200
g43765 and pi0515 n46081 ; n46201
g43766 nor pi0240 n46201 ; n46202
g43767 and n46200_not n46202 ; n46203
g43768 nor n46138 n46203 ; n46204
g43769 nor pi0535 n46204 ; n46205
g43770 and pi0515 n46199 ; n46206
g43771 and pi0515_not n46081 ; n46207
g43772 and pi0240 n46207_not ; n46208
g43773 and n46206_not n46208 ; n46209
g43774 nor n46140 n46209 ; n46210
g43775 and pi0535 n46210_not ; n46211
g43776 nor n46205 n46211 ; n46212
g43777 and pi0534_not n46212 ; n46213
g43778 and pi0534 n46141 ; n46214
g43779 and pi0239 n46214_not ; n46215
g43780 and n46213_not n46215 ; n46216
g43781 nor n46087 n46216 ; n46217
g43782 nor pi0488 n46217 ; n46218
g43783 and pi0534 n46212 ; n46219
g43784 and pi0534_not n46141 ; n46220
g43785 nor pi0239 n46220 ; n46221
g43786 and n46219_not n46221 ; n46222
g43787 nor n46089 n46222 ; n46223
g43788 and pi0488 n46223_not ; n46224
g43789 nor n46218 n46224 ; n46225
g43790 and pi0504_not n46225 ; n46226
g43791 and pi0504 n46145 ; n46227
g43792 nor pi0242 n46227 ; n46228
g43793 and n46226_not n46228 ; n46229
g43794 nor n46092 n46229 ; n46230
g43795 nor pi0510 n46230 ; n46231
g43796 and pi0504 n46225 ; n46232
g43797 and pi0504_not n46145 ; n46233
g43798 and pi0242 n46233_not ; n46234
g43799 and n46232_not n46234 ; n46235
g43800 nor n46094 n46235 ; n46236
g43801 and pi0510 n46236_not ; n46237
g43802 nor n46231 n46237 ; n46238
g43803 and pi0533_not n46238 ; n46239
g43804 and pi0533 n46149 ; n46240
g43805 nor pi0235 n46240 ; n46241
g43806 and n46239_not n46241 ; n46242
g43807 nor n46097 n46242 ; n46243
g43808 nor pi0512 n46243 ; n46244
g43809 and pi0533 n46238 ; n46245
g43810 and pi0533_not n46149 ; n46246
g43811 and pi0235 n46246_not ; n46247
g43812 and n46245_not n46247 ; n46248
g43813 nor n46099 n46248 ; n46249
g43814 and pi0512 n46249_not ; n46250
g43815 nor n46244 n46250 ; n46251
g43816 and pi0558_not n46251 ; n46252
g43817 and pi0558 n46153 ; n46253
g43818 nor pi0244 n46253 ; n46254
g43819 and n46252_not n46254 ; n46255
g43820 nor n46102 n46255 ; n46256
g43821 nor pi0513 n46256 ; n46257
g43822 and pi0558 n46251 ; n46258
g43823 and pi0558_not n46153 ; n46259
g43824 and pi0244 n46259_not ; n46260
g43825 and n46258_not n46260 ; n46261
g43826 nor n46104 n46261 ; n46262
g43827 and pi0513 n46262_not ; n46263
g43828 nor n46257 n46263 ; n46264
g43829 and pi0509_not n46264 ; n46265
g43830 and pi0509 n46157 ; n46266
g43831 nor pi0245 n46266 ; n46267
g43832 and n46265_not n46267 ; n46268
g43833 nor n46107 n46268 ; n46269
g43834 nor pi0514 n46269 ; n46270
g43835 and pi0509 n46264 ; n46271
g43836 and pi0509_not n46157 ; n46272
g43837 and pi0245 n46272_not ; n46273
g43838 and n46271_not n46273 ; n46274
g43839 nor n46109 n46274 ; n46275
g43840 and pi0514 n46275_not ; n46276
g43841 nor n46270 n46276 ; n46277
g43842 and pi0508_not n46277 ; n46278
g43843 and pi0508 n46161 ; n46279
g43844 nor pi0247 n46279 ; n46280
g43845 and n46278_not n46280 ; n46281
g43846 nor n46112 n46281 ; n46282
g43847 nor pi0516 n46282 ; n46283
g43848 and pi0508 n46277 ; n46284
g43849 and pi0508_not n46161 ; n46285
g43850 and pi0247 n46285_not ; n46286
g43851 and n46284_not n46286 ; n46287
g43852 nor n46114 n46287 ; n46288
g43853 and pi0516 n46288_not ; n46289
g43854 nor n46283 n46289 ; n46290
g43855 and pi0238_not n46290 ; n46291
g43856 nor pi0517 n46291 ; n46292
g43857 nor pi0507 n46168 ; n46293
g43858 and n46292_not n46293 ; n46294
g43859 and pi0238 n46115 ; n46295
g43860 and pi0238_not n46165 ; n46296
g43861 nor pi0517 n46296 ; n46297
g43862 and n46295_not n46297 ; n46298
g43863 and pi0238 n46290 ; n46299
g43864 and pi0517 n46299_not ; n46300
g43865 and pi0507 n46298_not ; n46301
g43866 and n46300_not n46301 ; n46302
g43867 nor n46294 n46302 ; n46303
g43868 and pi0233 n46303_not ; n46304
g43869 and pi0237 n46060_not ; n46305
g43870 and n46304_not n46305 ; n46306
g43871 nor pi0240 pi0492 ; n46307
g43872 and pi0240 pi0492 ; n46308
g43873 nor n46307 n46308 ; n46309
g43874 and pi0241 pi0490 ; n46310
g43875 nor pi0241 pi0490 ; n46311
g43876 nor n46310 n46311 ; n46312
g43877 and pi0248 pi0548 ; n46313
g43878 nor pi0248 pi0548 ; n46314
g43879 nor n46313 n46314 ; n46315
g43880 and pi0249 pi0484 ; n46316
g43881 nor pi0249 pi0484 ; n46317
g43882 nor n46316 n46317 ; n46318
g43883 and pi0246 pi0546 ; n46319
g43884 nor pi0246 pi0546 ; n46320
g43885 nor n46319 n46320 ; n46321
g43886 nor pi0544 n45431 ; n46322
g43887 and pi0544 n45903_not ; n46323
g43888 nor n46315 n46318 ; n46324
g43889 and n46321_not n46324 ; n46325
g43890 and n46322_not n46325 ; n46326
g43891 and n46323_not n46326 ; n46327
g43892 and n46312_not n46327 ; n46328
g43893 and n46309_not n46328 ; n46329
g43894 and pi0494 n46329 ; n46330
g43895 nor pi0239 n46330 ; n46331
g43896 and pi0494_not n46329 ; n46332
g43897 and pi0239 n46332_not ; n46333
g43898 nor n46331 n46333 ; n46334
g43899 and pi0483 n46334 ; n46335
g43900 and pi0242 n46335_not ; n46336
g43901 and pi0483_not n46334 ; n46337
g43902 nor pi0242 n46337 ; n46338
g43903 nor n46336 n46338 ; n46339
g43904 and pi0495 n46339 ; n46340
g43905 and pi0235 n46340_not ; n46341
g43906 and pi0495_not n46339 ; n46342
g43907 nor pi0235 n46342 ; n46343
g43908 nor n46341 n46343 ; n46344
g43909 and pi0244 pi0493 ; n46345
g43910 nor pi0244 pi0493 ; n46346
g43911 nor n46345 n46346 ; n46347
g43912 and n46344 n46347_not ; n46348
g43913 and pi0545 n46348 ; n46349
g43914 and pi0245 n46349_not ; n46350
g43915 and pi0545_not n46348 ; n46351
g43916 nor pi0245 n46351 ; n46352
g43917 nor n46350 n46352 ; n46353
g43918 and pi0547 n46353 ; n46354
g43919 and pi0247 n46354_not ; n46355
g43920 and pi0547_not n46353 ; n46356
g43921 nor pi0247 n46356 ; n46357
g43922 nor n46355 n46357 ; n46358
g43923 and pi0238_not n46358 ; n46359
g43924 and pi0523 n45845_not ; n46360
g43925 and pi0248 pi0576 ; n46361
g43926 nor pi0248 pi0576 ; n46362
g43927 nor n46361 n46362 ; n46363
g43928 and pi0249 pi0528 ; n46364
g43929 nor pi0249 pi0528 ; n46365
g43930 nor n46364 n46365 ; n46366
g43931 and pi0246 pi0526 ; n46367
g43932 nor pi0246 pi0526 ; n46368
g43933 nor n46367 n46368 ; n46369
g43934 nor pi0523 n45455 ; n46370
g43935 nor n46363 n46366 ; n46371
g43936 and n46369_not n46371 ; n46372
g43937 and n46360_not n46372 ; n46373
g43938 and n46370_not n46373 ; n46374
g43939 and pi0571 n46374 ; n46375
g43940 and pi0241 n46375_not ; n46376
g43941 and pi0571_not n46374 ; n46377
g43942 nor pi0241 n46377 ; n46378
g43943 nor n46376 n46378 ; n46379
g43944 and pi0530_not n46379 ; n46380
g43945 nor pi0240 n46380 ; n46381
g43946 and pi0530 n46379 ; n46382
g43947 and pi0240 n46382_not ; n46383
g43948 nor n46381 n46383 ; n46384
g43949 and pi0239_not pi0524 ; n46385
g43950 and pi0239 pi0524_not ; n46386
g43951 nor n46385 n46386 ; n46387
g43952 and n46384 n46387_not ; n46388
g43953 and pi0242 pi0573 ; n46389
g43954 nor pi0242 pi0573 ; n46390
g43955 nor n46389 n46390 ; n46391
g43956 and n46388 n46391_not ; n46392
g43957 and pi0235 pi0575 ; n46393
g43958 nor pi0235 pi0575 ; n46394
g43959 nor n46393 n46394 ; n46395
g43960 and n46392 n46395_not ; n46396
g43961 and pi0572 n46396 ; n46397
g43962 and pi0244 n46397_not ; n46398
g43963 and pi0572_not n46396 ; n46399
g43964 nor pi0244 n46399 ; n46400
g43965 nor n46398 n46400 ; n46401
g43966 and pi0245 pi0525 ; n46402
g43967 nor pi0245 pi0525 ; n46403
g43968 nor n46402 n46403 ; n46404
g43969 and n46401 n46404_not ; n46405
g43970 and pi0247 pi0527 ; n46406
g43971 nor pi0247 pi0527 ; n46407
g43972 nor n46406 n46407 ; n46408
g43973 and n46405 n46408_not ; n46409
g43974 and pi0238 n46409 ; n46410
g43975 and pi0529 n46410_not ; n46411
g43976 and n46359_not n46411 ; n46412
g43977 nor n46307 n46381 ; n46413
g43978 and pi0530 n46328_not ; n46414
g43979 nor pi0241 n46327 ; n46415
g43980 and n46377_not n46415 ; n46416
g43981 nor n46376 n46416 ; n46417
g43982 nor pi0490 n46417 ; n46418
g43983 and pi0241 n46327_not ; n46419
g43984 and n46375_not n46419 ; n46420
g43985 nor n46378 n46420 ; n46421
g43986 and pi0490 n46421_not ; n46422
g43987 nor n46418 n46422 ; n46423
g43988 nor pi0530 n46423 ; n46424
g43989 nor pi0492 n46414 ; n46425
g43990 and n46424_not n46425 ; n46426
g43991 nor n46413 n46426 ; n46427
g43992 nor n46308 n46383 ; n46428
g43993 nor pi0530 n46328 ; n46429
g43994 and pi0530 n46423_not ; n46430
g43995 and pi0492 n46429_not ; n46431
g43996 and n46430_not n46431 ; n46432
g43997 nor n46428 n46432 ; n46433
g43998 nor n46427 n46433 ; n46434
g43999 and pi0494_not n46434 ; n46435
g44000 and pi0494 n46384 ; n46436
g44001 and pi0239 n46436_not ; n46437
g44002 and n46435_not n46437 ; n46438
g44003 nor n46331 n46438 ; n46439
g44004 nor pi0524 n46439 ; n46440
g44005 and pi0494 n46434 ; n46441
g44006 and pi0494_not n46384 ; n46442
g44007 nor pi0239 n46442 ; n46443
g44008 and n46441_not n46443 ; n46444
g44009 nor n46333 n46444 ; n46445
g44010 and pi0524 n46445_not ; n46446
g44011 nor n46440 n46446 ; n46447
g44012 and pi0483_not n46447 ; n46448
g44013 and pi0483 n46388 ; n46449
g44014 nor pi0242 n46449 ; n46450
g44015 and n46448_not n46450 ; n46451
g44016 nor n46336 n46451 ; n46452
g44017 nor pi0573 n46452 ; n46453
g44018 and pi0483 n46447 ; n46454
g44019 and pi0483_not n46388 ; n46455
g44020 and pi0242 n46455_not ; n46456
g44021 and n46454_not n46456 ; n46457
g44022 nor n46338 n46457 ; n46458
g44023 and pi0573 n46458_not ; n46459
g44024 nor n46453 n46459 ; n46460
g44025 and pi0495_not n46460 ; n46461
g44026 and pi0495 n46392 ; n46462
g44027 nor pi0235 n46462 ; n46463
g44028 and n46461_not n46463 ; n46464
g44029 nor n46341 n46464 ; n46465
g44030 nor pi0575 n46465 ; n46466
g44031 and pi0495 n46460 ; n46467
g44032 and pi0495_not n46392 ; n46468
g44033 and pi0235 n46468_not ; n46469
g44034 and n46467_not n46469 ; n46470
g44035 nor n46343 n46470 ; n46471
g44036 and pi0575 n46471_not ; n46472
g44037 nor n46466 n46472 ; n46473
g44038 and pi0572_not n46473 ; n46474
g44039 and pi0572 n46344 ; n46475
g44040 nor pi0244 n46475 ; n46476
g44041 and n46474_not n46476 ; n46477
g44042 nor n46398 n46477 ; n46478
g44043 nor pi0493 n46478 ; n46479
g44044 and pi0572 n46473 ; n46480
g44045 and pi0572_not n46344 ; n46481
g44046 and pi0244 n46481_not ; n46482
g44047 and n46480_not n46482 ; n46483
g44048 nor n46400 n46483 ; n46484
g44049 and pi0493 n46484_not ; n46485
g44050 nor n46479 n46485 ; n46486
g44051 and pi0545_not n46486 ; n46487
g44052 and pi0545 n46401 ; n46488
g44053 nor pi0245 n46488 ; n46489
g44054 and n46487_not n46489 ; n46490
g44055 nor n46350 n46490 ; n46491
g44056 nor pi0525 n46491 ; n46492
g44057 and pi0545 n46486 ; n46493
g44058 and pi0545_not n46401 ; n46494
g44059 and pi0245 n46494_not ; n46495
g44060 and n46493_not n46495 ; n46496
g44061 nor n46352 n46496 ; n46497
g44062 and pi0525 n46497_not ; n46498
g44063 nor n46492 n46498 ; n46499
g44064 and pi0547_not n46499 ; n46500
g44065 and pi0547 n46405 ; n46501
g44066 nor pi0247 n46501 ; n46502
g44067 and n46500_not n46502 ; n46503
g44068 nor n46355 n46503 ; n46504
g44069 nor pi0527 n46504 ; n46505
g44070 and pi0547 n46499 ; n46506
g44071 and pi0547_not n46405 ; n46507
g44072 and pi0247 n46507_not ; n46508
g44073 and n46506_not n46508 ; n46509
g44074 nor n46357 n46509 ; n46510
g44075 and pi0527 n46510_not ; n46511
g44076 nor n46505 n46511 ; n46512
g44077 and pi0238_not n46512 ; n46513
g44078 nor pi0529 n46513 ; n46514
g44079 nor pi0491 n46412 ; n46515
g44080 and n46514_not n46515 ; n46516
g44081 and pi0238 n46358 ; n46517
g44082 and pi0238_not n46409 ; n46518
g44083 nor pi0529 n46518 ; n46519
g44084 and n46517_not n46519 ; n46520
g44085 and pi0238 n46512 ; n46521
g44086 and pi0529 n46521_not ; n46522
g44087 and pi0491 n46520_not ; n46523
g44088 and n46522_not n46523 ; n46524
g44089 nor n46516 n46524 ; n46525
g44090 and pi0233 n46525_not ; n46526
g44091 and pi0485 n45903_not ; n46527
g44092 and pi0240 pi0551 ; n46528
g44093 nor pi0240 pi0551 ; n46529
g44094 nor n46528 n46529 ; n46530
g44095 and pi0249 pi0555_not ; n46531
g44096 and pi0249_not pi0555 ; n46532
g44097 and pi0241 pi0553_not ; n46533
g44098 and pi0241_not pi0553 ; n46534
g44099 and pi0248 pi0554_not ; n46535
g44100 and pi0248_not pi0554 ; n46536
g44101 and pi0246_not pi0563 ; n46537
g44102 and pi0246 pi0563_not ; n46538
g44103 nor pi0485 n45431 ; n46539
g44104 nor n46531 n46532 ; n46540
g44105 nor n46533 n46534 ; n46541
g44106 nor n46535 n46536 ; n46542
g44107 nor n46537 n46538 ; n46543
g44108 and n46542 n46543 ; n46544
g44109 and n46540 n46541 ; n46545
g44110 and n46530_not n46545 ; n46546
g44111 and n46544 n46546 ; n46547
g44112 and n46527_not n46547 ; n46548
g44113 and n46539_not n46548 ; n46549
g44114 and pi0550 n46549 ; n46550
g44115 nor pi0239 n46550 ; n46551
g44116 and pi0550_not n46549 ; n46552
g44117 and pi0239 n46552_not ; n46553
g44118 nor n46551 n46553 ; n46554
g44119 and pi0489_not n46554 ; n46555
g44120 nor pi0242 n46555 ; n46556
g44121 and pi0489 n46554 ; n46557
g44122 and pi0242 n46557_not ; n46558
g44123 nor n46556 n46558 ; n46559
g44124 and pi0549 n46559 ; n46560
g44125 and pi0235 n46560_not ; n46561
g44126 and pi0549_not n46559 ; n46562
g44127 nor pi0235 n46562 ; n46563
g44128 nor n46561 n46563 ; n46564
g44129 and pi0486 n46564 ; n46565
g44130 and pi0244 n46565_not ; n46566
g44131 and pi0486_not n46564 ; n46567
g44132 nor pi0244 n46567 ; n46568
g44133 nor n46566 n46568 ; n46569
g44134 and pi0245 pi0580 ; n46570
g44135 nor pi0245 pi0580 ; n46571
g44136 nor n46570 n46571 ; n46572
g44137 and n46569 n46572_not ; n46573
g44138 and pi0552 n46573 ; n46574
g44139 and pi0247 n46574_not ; n46575
g44140 and pi0552_not n46573 ; n46576
g44141 nor pi0247 n46576 ; n46577
g44142 nor n46575 n46577 ; n46578
g44143 and pi0238 n46578 ; n46579
g44144 nor pi0242 pi0556 ; n46580
g44145 and pi0242 pi0556 ; n46581
g44146 nor n46580 n46581 ; n46582
g44147 and pi0246 pi0564_not ; n46583
g44148 and pi0570 n45845_not ; n46584
g44149 and pi0246_not pi0564 ; n46585
g44150 and pi0249 pi0482_not ; n46586
g44151 and pi0249_not pi0482 ; n46587
g44152 and pi0241 pi0562 ; n46588
g44153 nor pi0241 pi0562 ; n46589
g44154 nor n46588 n46589 ; n46590
g44155 nor pi0570 n45455 ; n46591
g44156 nor n46585 n46586 ; n46592
g44157 and n46587_not n46592 ; n46593
g44158 and n46590_not n46593 ; n46594
g44159 and n46584_not n46594 ; n46595
g44160 and n46591_not n46595 ; n46596
g44161 and pi0248 pi0565_not ; n46597
g44162 and pi0248_not pi0565 ; n46598
g44163 nor n46597 n46598 ; n46599
g44164 and pi0240 pi0560 ; n46600
g44165 nor pi0240 pi0560 ; n46601
g44166 nor n46600 n46601 ; n46602
g44167 and n46583_not n46599 ; n46603
g44168 and n46602_not n46603 ; n46604
g44169 and n46596 n46604 ; n46605
g44170 nor pi0240 n46605 ; n46606
g44171 and pi0560 n46583_not ; n46607
g44172 and n46599 n46607 ; n46608
g44173 and n46596 n46608 ; n46609
g44174 and pi0240 n46609_not ; n46610
g44175 nor n46606 n46610 ; n46611
g44176 and pi0239_not pi0569 ; n46612
g44177 and pi0239 pi0569_not ; n46613
g44178 nor n46612 n46613 ; n46614
g44179 and n46611 n46614_not ; n46615
g44180 and n46582_not n46615 ; n46616
g44181 and pi0235 pi0531 ; n46617
g44182 nor pi0235 pi0531 ; n46618
g44183 nor n46617 n46618 ; n46619
g44184 and n46616 n46619_not ; n46620
g44185 and pi0244 pi0566 ; n46621
g44186 nor pi0244 pi0566 ; n46622
g44187 nor n46621 n46622 ; n46623
g44188 and n46620 n46623_not ; n46624
g44189 and pi0568 n46624 ; n46625
g44190 and pi0245 n46625_not ; n46626
g44191 and pi0568_not n46624 ; n46627
g44192 nor pi0245 n46627 ; n46628
g44193 nor n46626 n46628 ; n46629
g44194 and pi0247 pi0532 ; n46630
g44195 nor pi0247 pi0532 ; n46631
g44196 nor n46630 n46631 ; n46632
g44197 and n46629 n46632_not ; n46633
g44198 and pi0238_not n46633 ; n46634
g44199 and pi0577 n46634_not ; n46635
g44200 and n46579_not n46635 ; n46636
g44201 nor n46556 n46580 ; n46637
g44202 and pi0489 n46615_not ; n46638
g44203 and n46605 n46613 ; n46639
g44204 and pi0569 n46553_not ; n46640
g44205 and n46611 n46640 ; n46641
g44206 nor n46554 n46639 ; n46642
g44207 and n46641_not n46642 ; n46643
g44208 and pi0489_not n46643 ; n46644
g44209 nor pi0556 n46638 ; n46645
g44210 and n46644_not n46645 ; n46646
g44211 nor n46637 n46646 ; n46647
g44212 nor n46558 n46581 ; n46648
g44213 nor pi0489 n46615 ; n46649
g44214 and pi0489 n46643 ; n46650
g44215 and pi0556 n46649_not ; n46651
g44216 and n46650_not n46651 ; n46652
g44217 nor n46648 n46652 ; n46653
g44218 nor n46647 n46653 ; n46654
g44219 and pi0549_not n46654 ; n46655
g44220 and pi0549 n46616 ; n46656
g44221 nor pi0235 n46656 ; n46657
g44222 and n46655_not n46657 ; n46658
g44223 nor n46561 n46658 ; n46659
g44224 nor pi0531 n46659 ; n46660
g44225 and pi0549 n46654 ; n46661
g44226 and pi0549_not n46616 ; n46662
g44227 and pi0235 n46662_not ; n46663
g44228 and n46661_not n46663 ; n46664
g44229 nor n46563 n46664 ; n46665
g44230 and pi0531 n46665_not ; n46666
g44231 nor n46660 n46666 ; n46667
g44232 and pi0486_not n46667 ; n46668
g44233 and pi0486 n46620 ; n46669
g44234 nor pi0244 n46669 ; n46670
g44235 and n46668_not n46670 ; n46671
g44236 nor n46566 n46671 ; n46672
g44237 nor pi0566 n46672 ; n46673
g44238 and pi0486 n46667 ; n46674
g44239 and pi0486_not n46620 ; n46675
g44240 and pi0244 n46675_not ; n46676
g44241 and n46674_not n46676 ; n46677
g44242 nor n46568 n46677 ; n46678
g44243 and pi0566 n46678_not ; n46679
g44244 nor n46673 n46679 ; n46680
g44245 and pi0568_not n46680 ; n46681
g44246 and pi0568 n46569 ; n46682
g44247 nor pi0245 n46682 ; n46683
g44248 and n46681_not n46683 ; n46684
g44249 nor n46626 n46684 ; n46685
g44250 nor pi0580 n46685 ; n46686
g44251 and pi0568 n46680 ; n46687
g44252 and pi0568_not n46569 ; n46688
g44253 and pi0245 n46688_not ; n46689
g44254 and n46687_not n46689 ; n46690
g44255 nor n46628 n46690 ; n46691
g44256 and pi0580 n46691_not ; n46692
g44257 nor n46686 n46692 ; n46693
g44258 and pi0552_not n46693 ; n46694
g44259 and pi0552 n46629 ; n46695
g44260 nor pi0247 n46695 ; n46696
g44261 and n46694_not n46696 ; n46697
g44262 nor n46575 n46697 ; n46698
g44263 nor pi0532 n46698 ; n46699
g44264 and pi0552 n46693 ; n46700
g44265 and pi0552_not n46629 ; n46701
g44266 and pi0247 n46701_not ; n46702
g44267 and n46700_not n46702 ; n46703
g44268 nor n46577 n46703 ; n46704
g44269 and pi0532 n46704_not ; n46705
g44270 nor n46699 n46705 ; n46706
g44271 and pi0238_not n46706 ; n46707
g44272 nor pi0577 n46707 ; n46708
g44273 nor pi0498 n46636 ; n46709
g44274 and n46708_not n46709 ; n46710
g44275 and pi0238_not n46578 ; n46711
g44276 and pi0238 n46633 ; n46712
g44277 nor pi0577 n46712 ; n46713
g44278 and n46711_not n46713 ; n46714
g44279 and pi0238 n46706 ; n46715
g44280 and pi0577 n46715_not ; n46716
g44281 and pi0498 n46714_not ; n46717
g44282 and n46716_not n46717 ; n46718
g44283 nor n46710 n46718 ; n46719
g44284 nor pi0233 n46719 ; n46720
g44285 nor pi0237 n46720 ; n46721
g44286 and n46526_not n46721 ; n46722
g44287 nor n46306 n46722 ; po0750
g44288 and pi0806_not n45126 ; n46724
g44289 nor pi0332 pi0806 ; n46725
g44290 and pi0990 n46725 ; n46726
g44291 and pi0600 n46726 ; n46727
g44292 and pi0332_not pi0594 ; n46728
g44293 nor n46727 n46728 ; n46729
g44294 nor n46724 n46729 ; po0751
g44295 and pi0605 pi0806_not ; n46731
g44296 and n45109 n46731 ; n46732
g44297 nor pi0595 n46732 ; n46733
g44298 and pi0595 n46732 ; n46734
g44299 nor pi0332 n46733 ; n46735
g44300 and n46734_not n46735 ; po0752
g44301 and pi0332_not pi0596 ; n46737
g44302 and pi0595 n45108 ; n46738
g44303 and n46726 n46738 ; n46739
g44304 nor n46737 n46739 ; n46740
g44305 and pi0596 n46739 ; n46741
g44306 nor n46740 n46741 ; po0753
g44307 nor pi0597 n46724 ; n46743
g44308 and pi0597 n46724 ; n46744
g44309 nor pi0332 n46743 ; n46745
g44310 and n46744_not n46745 ; po0754
g44311 nor pi0882 po1038 ; n46747
g44312 and pi0947 n46747 ; n46748
g44313 and pi0598 n46748_not ; n46749
g44314 and pi0740 pi0780 ; n46750
g44315 and n6192 n46750 ; n46751
g44316 or n46749 n46751 ; po0755
g44317 and pi0332_not pi0599 ; n46753
g44318 nor n46741 n46753 ; n46754
g44319 and pi0599 n46741 ; n46755
g44320 nor n46754 n46755 ; po0756
g44321 and pi0332_not pi0600 ; n46757
g44322 nor n46726 n46757 ; n46758
g44323 nor n46727 n46758 ; po0757
g44324 nor pi0806 pi0989 ; n46760
g44325 and pi0601_not pi0806 ; n46761
g44326 nor pi0332 n46760 ; n46762
g44327 and n46761_not n46762 ; po0758
g44328 and pi0230_not pi0602 ; n46764
g44329 nor pi0715 pi1160 ; n46765
g44330 and pi0715 pi1160 ; n46766
g44331 and pi0790 n46765_not ; n46767
g44332 and n46766_not n46767 ; n46768
g44333 and pi0230 n16644 ; n46769
g44334 and n17856_not n46769 ; n46770
g44335 nor n19146 n19342 ; n46771
g44336 and n46768_not n46771 ; n46772
g44337 and n46770 n46772 ; n46773
g44338 and n19151 n46773 ; n46774
g44339 or n46764 n46774 ; po0759
g44340 and pi0871 pi0966 ; n46776
g44341 and pi0872 pi0966 ; n46777
g44342 and pi0832 pi1100_not ; n46778
g44343 and pi0980_not pi1038 ; n46779
g44344 and pi1060 n46779 ; n46780
g44345 and pi0952 pi1061_not ; n46781
g44346 and n46780 n46781 ; n46782
g44347 and n46778 n46782 ; n46783
g44348 and pi0832 n46782 ; po0897
g44349 nor pi0603 po0897 ; n46785
g44350 nor pi0966 n46783 ; n46786
g44351 and n46785_not n46786 ; n46787
g44352 nor n46776 n46777 ; n46788
g44353 nand n46787_not n46788 ; po0760
g44354 and pi0823 n16657 ; n46790
g44355 and pi0779_not n46790 ; n46791
g44356 and pi0299_not pi0983 ; n46792
g44357 and pi0907 n46792 ; n46793
g44358 and pi0604 n46793_not ; n46794
g44359 and n46790_not n46794 ; n46795
g44360 or n46791 n46795 ; po0761
g44361 nor pi0605 n46725 ; n46797
g44362 nor pi0332 n46731 ; n46798
g44363 and n46797_not n46798 ; po0762
g44364 nor pi0606 po0897 ; n46800
g44365 and pi1104_not po0897 ; n46801
g44366 nor n46800 n46801 ; n46802
g44367 nor pi0966 n46802 ; n46803
g44368 and pi0837_not pi0966 ; n46804
g44369 nor n46803 n46804 ; po0763
g44370 nor pi0607 po0897 ; n46806
g44371 and pi1107_not po0897 ; n46807
g44372 nor pi0966 n46806 ; n46808
g44373 and n46807_not n46808 ; po0764
g44374 nor pi0608 po0897 ; n46810
g44375 and pi1116_not po0897 ; n46811
g44376 nor pi0966 n46810 ; n46812
g44377 and n46811_not n46812 ; po0765
g44378 nor pi0609 po0897 ; n46814
g44379 and pi1118_not po0897 ; n46815
g44380 nor pi0966 n46814 ; n46816
g44381 and n46815_not n46816 ; po0766
g44382 nor pi0610 po0897 ; n46818
g44383 and pi1113_not po0897 ; n46819
g44384 nor pi0966 n46818 ; n46820
g44385 and n46819_not n46820 ; po0767
g44386 nor pi0611 po0897 ; n46822
g44387 and pi1114_not po0897 ; n46823
g44388 nor pi0966 n46822 ; n46824
g44389 and n46823_not n46824 ; po0768
g44390 nor pi0612 po0897 ; n46826
g44391 and pi1111_not po0897 ; n46827
g44392 nor pi0966 n46826 ; n46828
g44393 and n46827_not n46828 ; po0769
g44394 nor pi0613 po0897 ; n46830
g44395 and pi1115_not po0897 ; n46831
g44396 nor pi0966 n46830 ; n46832
g44397 and n46831_not n46832 ; po0770
g44398 nor pi0614 po0897 ; n46834
g44399 and pi1102_not po0897 ; n46835
g44400 nor pi0966 n46834 ; n46836
g44401 and n46835_not n46836 ; n46837
g44402 or n46776 n46837 ; po0771
g44403 and pi0907 n46747 ; n46839
g44404 nor pi0615 n46839 ; n46840
g44405 and pi0779 pi0797 ; n46841
g44406 and n6195 n46841 ; n46842
g44407 or n46840 n46842 ; po0772
g44408 nor pi0616 po0897 ; n46844
g44409 and pi1101_not po0897 ; n46845
g44410 nor pi0966 n46844 ; n46846
g44411 and n46845_not n46846 ; n46847
g44412 or n46777 n46847 ; po0773
g44413 nor pi0617 po0897 ; n46849
g44414 and pi1105_not po0897 ; n46850
g44415 nor n46849 n46850 ; n46851
g44416 nor pi0966 n46851 ; n46852
g44417 and pi0850_not pi0966 ; n46853
g44418 nor n46852 n46853 ; po0774
g44419 nor pi0618 po0897 ; n46855
g44420 and pi1117_not po0897 ; n46856
g44421 nor pi0966 n46855 ; n46857
g44422 and n46856_not n46857 ; po0775
g44423 nor pi0619 po0897 ; n46859
g44424 and pi1122_not po0897 ; n46860
g44425 nor pi0966 n46859 ; n46861
g44426 and n46860_not n46861 ; po0776
g44427 nor pi0620 po0897 ; n46863
g44428 and pi1112_not po0897 ; n46864
g44429 nor pi0966 n46863 ; n46865
g44430 and n46864_not n46865 ; po0777
g44431 nor pi0621 po0897 ; n46867
g44432 and pi1108_not po0897 ; n46868
g44433 nor pi0966 n46867 ; n46869
g44434 and n46868_not n46869 ; po0778
g44435 nor pi0622 po0897 ; n46871
g44436 and pi1109_not po0897 ; n46872
g44437 nor pi0966 n46871 ; n46873
g44438 and n46872_not n46873 ; po0779
g44439 nor pi0623 po0897 ; n46875
g44440 and pi1106_not po0897 ; n46876
g44441 nor pi0966 n46875 ; n46877
g44442 and n46876_not n46877 ; po0780
g44443 and pi0831 n17167 ; n46879
g44444 and pi0780_not n46879 ; n46880
g44445 and pi0947 n46792 ; n46881
g44446 and pi0624 n46881_not ; n46882
g44447 and n46879_not n46882 ; n46883
g44448 or n46880 n46883 ; po0781
g44449 and pi0832 pi0973_not ; n46885
g44450 and pi1054_not pi1066 ; n46886
g44451 and pi1088 n46886 ; n46887
g44452 and n46885 n46887 ; n46888
g44453 and pi0953_not n46888 ; po0954
g44454 nor pi0625 po0954 ; n46890
g44455 and pi1116_not po0954 ; n46891
g44456 nor pi0962 n46890 ; n46892
g44457 and n46891_not n46892 ; po0782
g44458 nor pi0626 po0897 ; n46894
g44459 and pi1121_not po0897 ; n46895
g44460 nor pi0966 n46894 ; n46896
g44461 and n46895_not n46896 ; po0783
g44462 nor pi0627 po0954 ; n46898
g44463 and pi1117_not po0954 ; n46899
g44464 nor pi0962 n46898 ; n46900
g44465 and n46899_not n46900 ; po0784
g44466 nor pi0628 po0954 ; n46902
g44467 and pi1119_not po0954 ; n46903
g44468 nor pi0962 n46902 ; n46904
g44469 and n46903_not n46904 ; po0785
g44470 nor pi0629 po0897 ; n46906
g44471 and pi1119_not po0897 ; n46907
g44472 nor pi0966 n46906 ; n46908
g44473 and n46907_not n46908 ; po0786
g44474 nor pi0630 po0897 ; n46910
g44475 and pi1120_not po0897 ; n46911
g44476 nor pi0966 n46910 ; n46912
g44477 and n46911_not n46912 ; po0787
g44478 and pi1113_not po0954 ; n46914
g44479 and pi0631 po0954_not ; n46915
g44480 nor pi0962 n46914 ; n46916
g44481 and n46915_not n46916 ; po0788
g44482 and pi1115_not po0954 ; n46918
g44483 and pi0632 po0954_not ; n46919
g44484 nor pi0962 n46918 ; n46920
g44485 and n46919_not n46920 ; po0789
g44486 nor pi0633 po0897 ; n46922
g44487 and pi1110_not po0897 ; n46923
g44488 nor pi0966 n46922 ; n46924
g44489 and n46923_not n46924 ; po0790
g44490 nor pi0634 po0954 ; n46926
g44491 and pi1110_not po0954 ; n46927
g44492 nor pi0962 n46926 ; n46928
g44493 and n46927_not n46928 ; po0791
g44494 and pi1112_not po0954 ; n46930
g44495 and pi0635 po0954_not ; n46931
g44496 nor pi0962 n46930 ; n46932
g44497 and n46931_not n46932 ; po0792
g44498 nor pi0636 po0897 ; n46934
g44499 and pi1127_not po0897 ; n46935
g44500 nor pi0966 n46934 ; n46936
g44501 and n46935_not n46936 ; po0793
g44502 nor pi0637 po0954 ; n46938
g44503 and pi1105_not po0954 ; n46939
g44504 nor pi0962 n46938 ; n46940
g44505 and n46939_not n46940 ; po0794
g44506 nor pi0638 po0954 ; n46942
g44507 and pi1107_not po0954 ; n46943
g44508 nor pi0962 n46942 ; n46944
g44509 and n46943_not n46944 ; po0795
g44510 nor pi0639 po0954 ; n46946
g44511 and pi1109_not po0954 ; n46947
g44512 nor pi0962 n46946 ; n46948
g44513 and n46947_not n46948 ; po0796
g44514 nor pi0640 po0897 ; n46950
g44515 and pi1128_not po0897 ; n46951
g44516 nor pi0966 n46950 ; n46952
g44517 and n46951_not n46952 ; po0797
g44518 nor pi0641 po0954 ; n46954
g44519 and pi1121_not po0954 ; n46955
g44520 nor pi0962 n46954 ; n46956
g44521 and n46955_not n46956 ; po0798
g44522 nor pi0642 po0897 ; n46958
g44523 and pi1103_not po0897 ; n46959
g44524 nor pi0966 n46958 ; n46960
g44525 and n46959_not n46960 ; po0799
g44526 nor pi0643 po0954 ; n46962
g44527 and pi1104_not po0954 ; n46963
g44528 nor pi0962 n46962 ; n46964
g44529 and n46963_not n46964 ; po0800
g44530 nor pi0644 po0897 ; n46966
g44531 and pi1123_not po0897 ; n46967
g44532 nor pi0966 n46966 ; n46968
g44533 and n46967_not n46968 ; po0801
g44534 nor pi0645 po0897 ; n46970
g44535 and pi1125_not po0897 ; n46971
g44536 nor pi0966 n46970 ; n46972
g44537 and n46971_not n46972 ; po0802
g44538 and pi1114_not po0954 ; n46974
g44539 and pi0646 po0954_not ; n46975
g44540 nor pi0962 n46974 ; n46976
g44541 and n46975_not n46976 ; po0803
g44542 nor pi0647 po0954 ; n46978
g44543 and pi1120_not po0954 ; n46979
g44544 nor pi0962 n46978 ; n46980
g44545 and n46979_not n46980 ; po0804
g44546 nor pi0648 po0954 ; n46982
g44547 and pi1122_not po0954 ; n46983
g44548 nor pi0962 n46982 ; n46984
g44549 and n46983_not n46984 ; po0805
g44550 and pi1126_not po0954 ; n46986
g44551 and pi0649 po0954_not ; n46987
g44552 nor pi0962 n46986 ; n46988
g44553 and n46987_not n46988 ; po0806
g44554 and pi1127_not po0954 ; n46990
g44555 and pi0650 po0954_not ; n46991
g44556 nor pi0962 n46990 ; n46992
g44557 and n46991_not n46992 ; po0807
g44558 nor pi0651 po0897 ; n46994
g44559 and pi1130_not po0897 ; n46995
g44560 nor pi0966 n46994 ; n46996
g44561 and n46995_not n46996 ; po0808
g44562 nor pi0652 po0897 ; n46998
g44563 and pi1131_not po0897 ; n46999
g44564 nor pi0966 n46998 ; n47000
g44565 and n46999_not n47000 ; po0809
g44566 nor pi0653 po0897 ; n47002
g44567 and pi1129_not po0897 ; n47003
g44568 nor pi0966 n47002 ; n47004
g44569 and n47003_not n47004 ; po0810
g44570 and pi1130_not po0954 ; n47006
g44571 and pi0654 po0954_not ; n47007
g44572 nor pi0962 n47006 ; n47008
g44573 and n47007_not n47008 ; po0811
g44574 and pi1124_not po0954 ; n47010
g44575 and pi0655 po0954_not ; n47011
g44576 nor pi0962 n47010 ; n47012
g44577 and n47011_not n47012 ; po0812
g44578 nor pi0656 po0897 ; n47014
g44579 and pi1126_not po0897 ; n47015
g44580 nor pi0966 n47014 ; n47016
g44581 and n47015_not n47016 ; po0813
g44582 and pi1131_not po0954 ; n47018
g44583 and pi0657 po0954_not ; n47019
g44584 nor pi0962 n47018 ; n47020
g44585 and n47019_not n47020 ; po0814
g44586 nor pi0658 po0897 ; n47022
g44587 and pi1124_not po0897 ; n47023
g44588 nor pi0966 n47022 ; n47024
g44589 and n47023_not n47024 ; po0815
g44590 and pi0266 pi0992 ; n47026
g44591 and pi0280_not n47026 ; n47027
g44592 and pi0269_not n47027 ; n47028
g44593 and pi0281_not n47028 ; n47029
g44594 nor pi0270 pi0277 ; n47030
g44595 and pi0282_not n47030 ; n47031
g44596 and n47029 n47031 ; n47032
g44597 and pi0264_not n47032 ; n47033
g44598 and pi0265_not n47033 ; n47034
g44599 and pi0274_not n47034 ; po0959
g44600 and pi0274 n47034_not ; n47036
g44601 nor po0959 n47036 ; po0816
g44602 nor pi0660 po0954 ; n47038
g44603 and pi1118_not po0954 ; n47039
g44604 nor pi0962 n47038 ; n47040
g44605 and n47039_not n47040 ; po0817
g44606 nor pi0661 po0954 ; n47042
g44607 and pi1101_not po0954 ; n47043
g44608 nor pi0962 n47042 ; n47044
g44609 and n47043_not n47044 ; po0818
g44610 nor pi0662 po0954 ; n47046
g44611 and pi1102_not po0954 ; n47047
g44612 nor pi0962 n47046 ; n47048
g44613 and n47047_not n47048 ; po0819
g44614 nor pi0223 pi0224 ; n47050
g44615 nor pi0199 pi0257 ; n47051
g44616 and pi0199 pi1065_not ; n47052
g44617 nor n47050 n47051 ; n47053
g44618 and n47052_not n47053 ; n47054
g44619 and pi0592_not n8041 ; n47055
g44620 and pi0464 n47055 ; n47056
g44621 and pi0588 n47056_not ; n47057
g44622 and pi0591_not pi0592 ; n47058
g44623 and pi0365 n47058 ; n47059
g44624 and pi0334 pi0591 ; n47060
g44625 and pi0592_not n47060 ; n47061
g44626 nor n47059 n47061 ; n47062
g44627 nor pi0590 n47062 ; n47063
g44628 and pi0590 pi0591_not ; n47064
g44629 and pi0592_not n47064 ; n47065
g44630 and pi0323 n47065 ; n47066
g44631 nor pi0588 n47066 ; n47067
g44632 and n47063_not n47067 ; n47068
g44633 and n47050 n47057_not ; n47069
g44634 and n47068_not n47069 ; n47070
g44635 nor n47054 n47070 ; n47071
g44636 and n7643 n47071_not ; n47072
g44637 nor pi1137 pi1138 ; n47073
g44638 and pi1134_not n47073 ; n47074
g44639 nor pi0784 pi1136 ; n47075
g44640 and pi0634_not pi1136 ; n47076
g44641 and pi1135 n47075_not ; n47077
g44642 and n47076_not n47077 ; n47078
g44643 nor pi0815 pi1136 ; n47079
g44644 and pi0633_not pi1136 ; n47080
g44645 nor pi1135 n47079 ; n47081
g44646 and n47080_not n47081 ; n47082
g44647 nor n47078 n47082 ; n47083
g44648 and n47074 n47083_not ; n47084
g44649 and pi1135 n47073 ; n47085
g44650 and pi1136 n47085_not ; n47086
g44651 and pi0766_not n47086 ; n47087
g44652 nor pi0855 pi1136 ; n47088
g44653 and pi0700_not pi1135 ; n47089
g44654 and pi1135 pi1136_not ; n47090
g44655 and pi1134 n47073 ; n47091
g44656 and n47090_not n47091 ; n47092
g44657 nor n47088 n47089 ; n47093
g44658 and n47092 n47093 ; n47094
g44659 and n47087_not n47094 ; n47095
g44660 nor n47084 n47095 ; n47096
g44661 nor n7643 n47096 ; n47097
g44662 or n47072 n47097 ; po0820
g44663 and pi0429 n47055 ; n47099
g44664 and pi0588 n47099_not ; n47100
g44665 and pi0590_not pi0591 ; n47101
g44666 and pi0404 n47101 ; n47102
g44667 and pi0590_not pi0592 ; n47103
g44668 nor pi0588 n47103 ; n47104
g44669 and n47102_not n47104 ; n47105
g44670 and pi0380 pi0591_not ; n47106
g44671 and pi0592 n47106_not ; n47107
g44672 nor n47105 n47107 ; n47108
g44673 and pi0355 n47065 ; n47109
g44674 nor n47108 n47109 ; n47110
g44675 and n47050 n47100_not ; n47111
g44676 and n47110_not n47111 ; n47112
g44677 nor pi0199 pi0292 ; n47113
g44678 and pi0199 pi1084_not ; n47114
g44679 nor n47050 n47113 ; n47115
g44680 and n47114_not n47115 ; n47116
g44681 nor n47112 n47116 ; n47117
g44682 and n7643 n47117_not ; n47118
g44683 nor pi1135 pi1136 ; n47119
g44684 and pi0872 n47119 ; n47120
g44685 nor pi0772 pi1135 ; n47121
g44686 and pi0727_not pi1135 ; n47122
g44687 and pi1136 n47121_not ; n47123
g44688 and n47122_not n47123 ; n47124
g44689 and pi1134 n47120_not ; n47125
g44690 and n47124_not n47125 ; n47126
g44691 and n7643_not n47073 ; n47127
g44692 and pi0614 pi1135_not ; n47128
g44693 and pi0662 pi1135 ; n47129
g44694 and pi1136 n47128_not ; n47130
g44695 and n47129_not n47130 ; n47131
g44696 and pi0811 pi1135_not ; n47132
g44697 and pi0785 pi1135 ; n47133
g44698 nor pi1136 n47132 ; n47134
g44699 and n47133_not n47134 ; n47135
g44700 nor n47131 n47135 ; n47136
g44701 nor pi1134 n47136 ; n47137
g44702 and n47126_not n47127 ; n47138
g44703 and n47137_not n47138 ; n47139
g44704 or n47118 n47139 ; po0821
g44705 nor pi0665 po0954 ; n47141
g44706 and pi1108_not po0954 ; n47142
g44707 nor pi0962 n47141 ; n47143
g44708 and n47142_not n47143 ; po0822
g44709 nor pi0607 pi1135 ; n47145
g44710 and pi0638_not pi1135 ; n47146
g44711 and pi1136 n47145_not ; n47147
g44712 and n47146_not n47147 ; n47148
g44713 and pi0790_not pi1135 ; n47149
g44714 and pi0799 pi1135_not ; n47150
g44715 nor pi1136 n47149 ; n47151
g44716 and n47150_not n47151 ; n47152
g44717 nor n47148 n47152 ; n47153
g44718 and n47074 n47153_not ; n47154
g44719 and pi0764_not n47086 ; n47155
g44720 and pi0691_not pi1135 ; n47156
g44721 nor pi0873 pi1136 ; n47157
g44722 nor n47156 n47157 ; n47158
g44723 and n47092 n47158 ; n47159
g44724 and n47155_not n47159 ; n47160
g44725 nor n47154 n47160 ; n47161
g44726 nor n7643 n47161 ; n47162
g44727 nor pi0199 pi0297 ; n47163
g44728 and pi0199 pi1044_not ; n47164
g44729 nor n47050 n47163 ; n47165
g44730 and n47164_not n47165 ; n47166
g44731 and pi0443 n47055 ; n47167
g44732 and pi0588 n47167_not ; n47168
g44733 and pi0456 n47101 ; n47169
g44734 and n47104 n47169_not ; n47170
g44735 and pi0337 pi0591_not ; n47171
g44736 and pi0592 n47171_not ; n47172
g44737 nor n47170 n47172 ; n47173
g44738 and pi0441 n47065 ; n47174
g44739 nor n47173 n47174 ; n47175
g44740 and n47050 n47168_not ; n47176
g44741 and n47175_not n47176 ; n47177
g44742 nor n47166 n47177 ; n47178
g44743 and n7643 n47178_not ; n47179
g44744 or n47162 n47179 ; po0823
g44745 and pi0444 n47055 ; n47181
g44746 and pi0588 n47181_not ; n47182
g44747 and pi0319 n47101 ; n47183
g44748 and n47104 n47183_not ; n47184
g44749 and pi0338 pi0591_not ; n47185
g44750 and pi0592 n47185_not ; n47186
g44751 nor n47184 n47186 ; n47187
g44752 and pi0458 n47065 ; n47188
g44753 nor n47187 n47188 ; n47189
g44754 and n47050 n47182_not ; n47190
g44755 and n47189_not n47190 ; n47191
g44756 nor pi0199 pi0294 ; n47192
g44757 and pi0199 pi1072_not ; n47193
g44758 nor n47050 n47192 ; n47194
g44759 and n47193_not n47194 ; n47195
g44760 nor n47191 n47195 ; n47196
g44761 and n7643 n47196_not ; n47197
g44762 and pi0871 n47119 ; n47198
g44763 nor pi0763 pi1135 ; n47199
g44764 and pi0699_not pi1135 ; n47200
g44765 and pi1136 n47199_not ; n47201
g44766 and n47200_not n47201 ; n47202
g44767 and pi1134 n47198_not ; n47203
g44768 and n47202_not n47203 ; n47204
g44769 and pi0792 pi1136_not ; n47205
g44770 and pi0681 pi1136 ; n47206
g44771 and pi1135 n47205_not ; n47207
g44772 and n47206_not n47207 ; n47208
g44773 nor pi0809 pi1136 ; n47209
g44774 and pi0642 pi1136 ; n47210
g44775 nor pi1135 n47209 ; n47211
g44776 and n47210_not n47211 ; n47212
g44777 nor n47208 n47212 ; n47213
g44778 nor pi1134 n47213 ; n47214
g44779 and n47127 n47204_not ; n47215
g44780 and n47214_not n47215 ; n47216
g44781 or n47197 n47216 ; po0824
g44782 nor pi0603 pi1135 ; n47218
g44783 and pi0680_not pi1135 ; n47219
g44784 and pi1136 n47218_not ; n47220
g44785 and n47219_not n47220 ; n47221
g44786 nor pi0981 pi1135 ; n47222
g44787 and pi0778_not pi1135 ; n47223
g44788 nor pi1136 n47222 ; n47224
g44789 and n47223_not n47224 ; n47225
g44790 nor n47221 n47225 ; n47226
g44791 and n47074 n47226_not ; n47227
g44792 and pi0759_not n47086 ; n47228
g44793 and pi0696_not pi1135 ; n47229
g44794 nor pi0837 pi1136 ; n47230
g44795 nor n47229 n47230 ; n47231
g44796 and n47092 n47231 ; n47232
g44797 and n47228_not n47232 ; n47233
g44798 nor n47227 n47233 ; n47234
g44799 nor n7643 n47234 ; n47235
g44800 nor pi0199 pi0291 ; n47236
g44801 and pi0199 pi1049_not ; n47237
g44802 nor n47050 n47236 ; n47238
g44803 and n47237_not n47238 ; n47239
g44804 and pi0414 n47055 ; n47240
g44805 and pi0588 n47240_not ; n47241
g44806 and pi0390 n47101 ; n47242
g44807 and n47104 n47242_not ; n47243
g44808 and pi0363 pi0591_not ; n47244
g44809 and pi0592 n47244_not ; n47245
g44810 nor n47243 n47245 ; n47246
g44811 and pi0342 n47065 ; n47247
g44812 nor n47246 n47247 ; n47248
g44813 and n47050 n47241_not ; n47249
g44814 and n47248_not n47249 ; n47250
g44815 nor n47239 n47250 ; n47251
g44816 and n7643 n47251_not ; n47252
g44817 or n47235 n47252 ; po0825
g44818 and pi1125_not po0954 ; n47254
g44819 and pi0669 po0954_not ; n47255
g44820 nor pi0962 n47254 ; n47256
g44821 and n47255_not n47256 ; po0826
g44822 nor pi0199 pi0258 ; n47258
g44823 and pi0199 pi1062_not ; n47259
g44824 nor n47050 n47258 ; n47260
g44825 and n47259_not n47260 ; n47261
g44826 and pi0415 n47055 ; n47262
g44827 and pi0588 n47262_not ; n47263
g44828 and pi0364 n47058 ; n47264
g44829 and pi0391 pi0591 ; n47265
g44830 and pi0592_not n47265 ; n47266
g44831 nor n47264 n47266 ; n47267
g44832 nor pi0590 n47267 ; n47268
g44833 and pi0343 n47065 ; n47269
g44834 nor pi0588 n47269 ; n47270
g44835 and n47268_not n47270 ; n47271
g44836 and n47050 n47263_not ; n47272
g44837 and n47271_not n47272 ; n47273
g44838 nor n47261 n47273 ; n47274
g44839 and n7643 n47274_not ; n47275
g44840 and pi0723 pi1135 ; n47276
g44841 nor pi0852 pi1136 ; n47277
g44842 and pi0745 n47086 ; n47278
g44843 nor n47276 n47277 ; n47279
g44844 and n47092 n47279 ; n47280
g44845 and n47278_not n47280 ; n47281
g44846 and pi0695 pi1135 ; n47282
g44847 and pi1136 n47073 ; n47283
g44848 nor pi0612 pi1135 ; n47284
g44849 nor pi1134 n47282 ; n47285
g44850 and n47284_not n47285 ; n47286
g44851 and n47283 n47286 ; n47287
g44852 nor n47281 n47287 ; n47288
g44853 nor n7643 n47288 ; n47289
g44854 or n47275 n47289 ; po0827
g44855 nor pi0199 pi0261 ; n47291
g44856 and pi0199 pi1040_not ; n47292
g44857 nor n47050 n47291 ; n47293
g44858 and n47292_not n47293 ; n47294
g44859 and pi0453 n47055 ; n47295
g44860 and pi0588 n47295_not ; n47296
g44861 and pi0447 n47058 ; n47297
g44862 and pi0333 pi0591 ; n47298
g44863 and pi0592_not n47298 ; n47299
g44864 nor n47297 n47299 ; n47300
g44865 nor pi0590 n47300 ; n47301
g44866 and pi0327 n47065 ; n47302
g44867 nor pi0588 n47302 ; n47303
g44868 and n47301_not n47303 ; n47304
g44869 and n47050 n47296_not ; n47305
g44870 and n47304_not n47305 ; n47306
g44871 nor n47294 n47306 ; n47307
g44872 and n7643 n47307_not ; n47308
g44873 and pi0724 pi1135 ; n47309
g44874 nor pi0865 pi1136 ; n47310
g44875 and pi0741 n47086 ; n47311
g44876 nor n47309 n47310 ; n47312
g44877 and n47092 n47312 ; n47313
g44878 and n47311_not n47313 ; n47314
g44879 and pi0646 pi1135 ; n47315
g44880 nor pi0611 pi1135 ; n47316
g44881 nor pi1134 n47315 ; n47317
g44882 and n47316_not n47317 ; n47318
g44883 and n47283 n47318 ; n47319
g44884 nor n47314 n47319 ; n47320
g44885 nor n7643 n47320 ; n47321
g44886 or n47308 n47321 ; po0828
g44887 nor pi0616 pi1135 ; n47323
g44888 and pi0661_not pi1135 ; n47324
g44889 and pi1136 n47323_not ; n47325
g44890 and n47324_not n47325 ; n47326
g44891 nor pi0808 pi1135 ; n47327
g44892 and pi0781_not pi1135 ; n47328
g44893 nor pi1136 n47327 ; n47329
g44894 and n47328_not n47329 ; n47330
g44895 nor n47326 n47330 ; n47331
g44896 and n47074 n47331_not ; n47332
g44897 and pi0758_not n47086 ; n47333
g44898 and pi0736_not pi1135 ; n47334
g44899 nor pi0850 pi1136 ; n47335
g44900 nor n47334 n47335 ; n47336
g44901 and n47092 n47336 ; n47337
g44902 and n47333_not n47337 ; n47338
g44903 nor n47332 n47338 ; n47339
g44904 nor n7643 n47339 ; n47340
g44905 nor pi0199 pi0290 ; n47341
g44906 and pi0199 pi1048_not ; n47342
g44907 nor n47050 n47341 ; n47343
g44908 and n47342_not n47343 ; n47344
g44909 and pi0422 n47055 ; n47345
g44910 and pi0588 n47345_not ; n47346
g44911 and pi0397 n47101 ; n47347
g44912 and n47104 n47347_not ; n47348
g44913 and pi0372 pi0591_not ; n47349
g44914 and pi0592 n47349_not ; n47350
g44915 nor n47348 n47350 ; n47351
g44916 and pi0320 n47065 ; n47352
g44917 nor n47351 n47352 ; n47353
g44918 and n47050 n47346_not ; n47354
g44919 and n47353_not n47354 ; n47355
g44920 nor n47344 n47355 ; n47356
g44921 and n7643 n47356_not ; n47357
g44922 or n47340 n47357 ; po0829
g44923 nor pi0617 pi1135 ; n47359
g44924 and pi0637_not pi1135 ; n47360
g44925 and pi1136 n47359_not ; n47361
g44926 and n47360_not n47361 ; n47362
g44927 and pi0788_not pi1135 ; n47363
g44928 and pi0814 pi1135_not ; n47364
g44929 nor pi1136 n47363 ; n47365
g44930 and n47364_not n47365 ; n47366
g44931 nor n47362 n47366 ; n47367
g44932 and n47074 n47367_not ; n47368
g44933 and pi0749_not n47086 ; n47369
g44934 and pi0706_not pi1135 ; n47370
g44935 nor pi0866 pi1136 ; n47371
g44936 nor n47370 n47371 ; n47372
g44937 and n47092 n47372 ; n47373
g44938 and n47369_not n47373 ; n47374
g44939 nor n47368 n47374 ; n47375
g44940 nor n7643 n47375 ; n47376
g44941 nor pi0199 pi0295 ; n47377
g44942 and pi0199 pi1053_not ; n47378
g44943 nor n47050 n47377 ; n47379
g44944 and n47378_not n47379 ; n47380
g44945 and pi0435 n47055 ; n47381
g44946 and pi0588 n47381_not ; n47382
g44947 and pi0411 n47101 ; n47383
g44948 and n47104 n47383_not ; n47384
g44949 and pi0387 pi0591_not ; n47385
g44950 and pi0592 n47385_not ; n47386
g44951 nor n47384 n47386 ; n47387
g44952 and pi0452 n47065 ; n47388
g44953 nor n47387 n47388 ; n47389
g44954 and n47050 n47382_not ; n47390
g44955 and n47389_not n47390 ; n47391
g44956 nor n47380 n47391 ; n47392
g44957 and n7643 n47392_not ; n47393
g44958 or n47376 n47393 ; po0830
g44959 nor pi0199 pi0256 ; n47395
g44960 and pi0199 pi1070_not ; n47396
g44961 nor n47050 n47395 ; n47397
g44962 and n47396_not n47397 ; n47398
g44963 and pi0437 n47055 ; n47399
g44964 and pi0588 n47399_not ; n47400
g44965 and pi0336 n47058 ; n47401
g44966 and pi0463 pi0591 ; n47402
g44967 and pi0592_not n47402 ; n47403
g44968 nor n47401 n47403 ; n47404
g44969 nor pi0590 n47404 ; n47405
g44970 and pi0362 n47065 ; n47406
g44971 nor pi0588 n47406 ; n47407
g44972 and n47405_not n47407 ; n47408
g44973 and n47050 n47400_not ; n47409
g44974 and n47408_not n47409 ; n47410
g44975 nor n47398 n47410 ; n47411
g44976 and n7643 n47411_not ; n47412
g44977 and pi0859 n47119 ; n47413
g44978 nor pi0743 pi1135 ; n47414
g44979 and pi0735_not pi1135 ; n47415
g44980 and pi1136 n47414_not ; n47416
g44981 and n47415_not n47416 ; n47417
g44982 and pi1134 n47413_not ; n47418
g44983 and n47417_not n47418 ; n47419
g44984 and pi0622 pi1135_not ; n47420
g44985 and pi0639 pi1135 ; n47421
g44986 and pi1136 n47420_not ; n47422
g44987 and n47421_not n47422 ; n47423
g44988 and pi0804 pi1135_not ; n47424
g44989 and pi0783 pi1135 ; n47425
g44990 nor pi1136 n47424 ; n47426
g44991 and n47425_not n47426 ; n47427
g44992 nor n47423 n47427 ; n47428
g44993 nor pi1134 n47428 ; n47429
g44994 and n47127 n47419_not ; n47430
g44995 and n47429_not n47430 ; n47431
g44996 or n47412 n47431 ; po0831
g44997 and pi0876 n47119 ; n47433
g44998 nor pi0748 pi1135 ; n47434
g44999 and pi0730_not pi1135 ; n47435
g45000 and pi1136 n47434_not ; n47436
g45001 and n47435_not n47436 ; n47437
g45002 nor n47433 n47437 ; n47438
g45003 and n47091 n47438_not ; n47439
g45004 and pi0623_not n47086 ; n47440
g45005 and pi0789 n47090 ; n47441
g45006 and pi0710_not pi1135 ; n47442
g45007 and pi1136 n47442_not ; n47443
g45008 nor pi0803 pi1135 ; n47444
g45009 nor n47441 n47444 ; n47445
g45010 and n47443_not n47445 ; n47446
g45011 and n47074 n47440_not ; n47447
g45012 and n47446_not n47447 ; n47448
g45013 nor n47439 n47448 ; n47449
g45014 nor n7643 n47449 ; n47450
g45015 nor pi0199 pi0296 ; n47451
g45016 and pi0199 pi1037_not ; n47452
g45017 nor n47050 n47451 ; n47453
g45018 and n47452_not n47453 ; n47454
g45019 and pi0436 n47055 ; n47455
g45020 and pi0588 n47455_not ; n47456
g45021 and pi0412 n47101 ; n47457
g45022 and n47104 n47457_not ; n47458
g45023 and pi0388 pi0591_not ; n47459
g45024 and pi0592 n47459_not ; n47460
g45025 nor n47458 n47460 ; n47461
g45026 and pi0455 n47065 ; n47462
g45027 nor n47461 n47462 ; n47463
g45028 and n47050 n47456_not ; n47464
g45029 and n47463_not n47464 ; n47465
g45030 nor n47454 n47465 ; n47466
g45031 and n7643 n47466_not ; n47467
g45032 or n47450 n47467 ; po0832
g45033 nor pi0606 pi1135 ; n47469
g45034 and pi0643_not pi1135 ; n47470
g45035 and pi1136 n47469_not ; n47471
g45036 and n47470_not n47471 ; n47472
g45037 and pi0787_not pi1135 ; n47473
g45038 and pi0812 pi1135_not ; n47474
g45039 nor pi1136 n47473 ; n47475
g45040 and n47474_not n47475 ; n47476
g45041 nor n47472 n47476 ; n47477
g45042 and n47074 n47477_not ; n47478
g45043 and pi0746_not n47086 ; n47479
g45044 and pi0729_not pi1135 ; n47480
g45045 nor pi0881 pi1136 ; n47481
g45046 nor n47480 n47481 ; n47482
g45047 and n47092 n47482 ; n47483
g45048 and n47479_not n47483 ; n47484
g45049 nor n47478 n47484 ; n47485
g45050 nor n7643 n47485 ; n47486
g45051 nor pi0199 pi0293 ; n47487
g45052 and pi0199 pi1059_not ; n47488
g45053 nor n47050 n47487 ; n47489
g45054 and n47488_not n47489 ; n47490
g45055 and pi0434 n47055 ; n47491
g45056 and pi0588 n47491_not ; n47492
g45057 and pi0410 n47101 ; n47493
g45058 and n47104 n47493_not ; n47494
g45059 and pi0386 pi0591_not ; n47495
g45060 and pi0592 n47495_not ; n47496
g45061 nor n47494 n47496 ; n47497
g45062 and pi0361 n47065 ; n47498
g45063 nor n47497 n47498 ; n47499
g45064 and n47050 n47492_not ; n47500
g45065 and n47499_not n47500 ; n47501
g45066 nor n47490 n47501 ; n47502
g45067 and n7643 n47502_not ; n47503
g45068 or n47486 n47503 ; po0833
g45069 nor pi0199 pi0259 ; n47505
g45070 and pi0199 pi1069_not ; n47506
g45071 nor n47050 n47505 ; n47507
g45072 and n47506_not n47507 ; n47508
g45073 and pi0416 n47055 ; n47509
g45074 and pi0588 n47509_not ; n47510
g45075 and pi0366 n47058 ; n47511
g45076 and pi0335 pi0591 ; n47512
g45077 and pi0592_not n47512 ; n47513
g45078 nor n47511 n47513 ; n47514
g45079 nor pi0590 n47514 ; n47515
g45080 and pi0344 n47065 ; n47516
g45081 nor pi0588 n47516 ; n47517
g45082 and n47515_not n47517 ; n47518
g45083 and n47050 n47510_not ; n47519
g45084 and n47518_not n47519 ; n47520
g45085 nor n47508 n47520 ; n47521
g45086 and n7643 n47521_not ; n47522
g45087 and pi0704 pi1135 ; n47523
g45088 nor pi0870 pi1136 ; n47524
g45089 and pi0742 n47086 ; n47525
g45090 nor n47523 n47524 ; n47526
g45091 and n47092 n47526 ; n47527
g45092 and n47525_not n47527 ; n47528
g45093 and pi0635 pi1135 ; n47529
g45094 nor pi0620 pi1135 ; n47530
g45095 nor pi1134 n47529 ; n47531
g45096 and n47530_not n47531 ; n47532
g45097 and n47283 n47532 ; n47533
g45098 nor n47528 n47533 ; n47534
g45099 nor n7643 n47534 ; n47535
g45100 or n47522 n47535 ; po0834
g45101 nor pi0199 pi0260 ; n47537
g45102 and pi0199 pi1067_not ; n47538
g45103 nor n47050 n47537 ; n47539
g45104 and n47538_not n47539 ; n47540
g45105 and pi0418 n47055 ; n47541
g45106 and pi0588 n47541_not ; n47542
g45107 and pi0368 n47058 ; n47543
g45108 and pi0393 pi0591 ; n47544
g45109 and pi0592_not n47544 ; n47545
g45110 nor n47543 n47545 ; n47546
g45111 nor pi0590 n47546 ; n47547
g45112 and pi0346 n47065 ; n47548
g45113 nor pi0588 n47548 ; n47549
g45114 and n47547_not n47549 ; n47550
g45115 and n47050 n47542_not ; n47551
g45116 and n47550_not n47551 ; n47552
g45117 nor n47540 n47552 ; n47553
g45118 and n7643 n47553_not ; n47554
g45119 and pi0688 pi1135 ; n47555
g45120 nor pi0856 pi1136 ; n47556
g45121 and pi0760 n47086 ; n47557
g45122 nor n47555 n47556 ; n47558
g45123 and n47092 n47558 ; n47559
g45124 and n47557_not n47559 ; n47560
g45125 and pi0632 pi1135 ; n47561
g45126 nor pi0613 pi1135 ; n47562
g45127 nor pi1134 n47561 ; n47563
g45128 and n47562_not n47563 ; n47564
g45129 and n47283 n47564 ; n47565
g45130 nor n47560 n47565 ; n47566
g45131 nor n7643 n47566 ; n47567
g45132 or n47554 n47567 ; po0835
g45133 nor pi0199 pi0255 ; n47569
g45134 and pi0199 pi1036_not ; n47570
g45135 nor n47050 n47569 ; n47571
g45136 and n47570_not n47571 ; n47572
g45137 and pi0438 n47055 ; n47573
g45138 and pi0588 n47573_not ; n47574
g45139 and pi0389 n47058 ; n47575
g45140 and pi0413 pi0591 ; n47576
g45141 and pi0592_not n47576 ; n47577
g45142 nor n47575 n47577 ; n47578
g45143 nor pi0590 n47578 ; n47579
g45144 and pi0450 n47065 ; n47580
g45145 nor pi0588 n47580 ; n47581
g45146 and n47579_not n47581 ; n47582
g45147 and n47050 n47574_not ; n47583
g45148 and n47582_not n47583 ; n47584
g45149 nor n47572 n47584 ; n47585
g45150 and n7643 n47585_not ; n47586
g45151 nor pi0791 pi1136 ; n47587
g45152 and pi0665_not pi1136 ; n47588
g45153 and pi1135 n47587_not ; n47589
g45154 and n47588_not n47589 ; n47590
g45155 nor pi0810 pi1136 ; n47591
g45156 and pi0621_not pi1136 ; n47592
g45157 nor pi1135 n47591 ; n47593
g45158 and n47592_not n47593 ; n47594
g45159 nor n47590 n47594 ; n47595
g45160 and n47074 n47595_not ; n47596
g45161 and pi0739_not n47086 ; n47597
g45162 nor pi0874 pi1136 ; n47598
g45163 and pi0690_not pi1135 ; n47599
g45164 nor n47598 n47599 ; n47600
g45165 and n47092 n47600 ; n47601
g45166 and n47597_not n47601 ; n47602
g45167 nor n47596 n47602 ; n47603
g45168 nor n7643 n47603 ; n47604
g45169 or n47586 n47604 ; po0836
g45170 nor pi0680 po0954 ; n47606
g45171 and pi1100_not po0954 ; n47607
g45172 nor pi0962 n47606 ; n47608
g45173 and n47607_not n47608 ; po0837
g45174 nor pi0681 po0954 ; n47610
g45175 and pi1103_not po0954 ; n47611
g45176 nor pi0962 n47610 ; n47612
g45177 and n47611_not n47612 ; po0838
g45178 nor pi0199 pi0251 ; n47614
g45179 and pi0199 pi1039_not ; n47615
g45180 nor n47050 n47614 ; n47616
g45181 and n47615_not n47616 ; n47617
g45182 and pi0417 n47055 ; n47618
g45183 and pi0588 n47618_not ; n47619
g45184 and pi0367 n47058 ; n47620
g45185 and pi0392 pi0591 ; n47621
g45186 and pi0592_not n47621 ; n47622
g45187 nor n47620 n47622 ; n47623
g45188 nor pi0590 n47623 ; n47624
g45189 and pi0345 n47065 ; n47625
g45190 nor pi0588 n47625 ; n47626
g45191 and n47624_not n47626 ; n47627
g45192 and n47050 n47619_not ; n47628
g45193 and n47627_not n47628 ; n47629
g45194 nor n47617 n47629 ; n47630
g45195 and n7643 n47630_not ; n47631
g45196 and pi0686 pi1135 ; n47632
g45197 nor pi0848 pi1136 ; n47633
g45198 and pi0757 n47086 ; n47634
g45199 nor n47632 n47633 ; n47635
g45200 and n47092 n47635 ; n47636
g45201 and n47634_not n47636 ; n47637
g45202 and pi0631 pi1135 ; n47638
g45203 nor pi0610 pi1135 ; n47639
g45204 nor pi1134 n47638 ; n47640
g45205 and n47639_not n47640 ; n47641
g45206 and n47283 n47641 ; n47642
g45207 nor n47637 n47642 ; n47643
g45208 nor n7643 n47643 ; n47644
g45209 or n47631 n47644 ; po0839
g45210 and pi0953 n46888 ; po0980
g45211 and pi1130_not po0980 ; n47647
g45212 and pi0684 po0980_not ; n47648
g45213 nor pi0962 n47647 ; n47649
g45214 and n47648_not n47649 ; po0841
g45215 and pi0590 pi0592_not ; n47651
g45216 and pi0357 n47651 ; n47652
g45217 and pi0382 n47103 ; n47653
g45218 nor n47652 n47653 ; n47654
g45219 nor pi0591 n47654 ; n47655
g45220 and pi0406 pi0592_not ; n47656
g45221 and n47101 n47656 ; n47657
g45222 nor n47655 n47657 ; n47658
g45223 nor pi0588 n47658 ; n47659
g45224 nor pi0591 pi0592 ; n47660
g45225 and pi0588 pi0590_not ; n47661
g45226 and pi0430 n47660 ; n47662
g45227 and n47661 n47662 ; n47663
g45228 nor n47659 n47663 ; n47664
g45229 and n47050 n47664_not ; n47665
g45230 and pi0199 pi1076_not ; n47666
g45231 nor n47050 n47666 ; n47667
g45232 and n42880_not n47667 ; n47668
g45233 nor n47665 n47668 ; n47669
g45234 and n7643 n47669_not ; n47670
g45235 and pi0860 n47119 ; n47671
g45236 and pi0744 pi1135_not ; n47672
g45237 and pi0728 pi1135 ; n47673
g45238 and pi1136 n47672_not ; n47674
g45239 and n47673_not n47674 ; n47675
g45240 nor n47671 n47675 ; n47676
g45241 and n47091 n47676_not ; n47677
g45242 and pi1136 n47073_not ; n47678
g45243 nor pi1134 n47678 ; n47679
g45244 nor pi0652 pi1135 ; n47680
g45245 and pi0657 pi1135 ; n47681
g45246 and pi1136 n47680_not ; n47682
g45247 and n47681_not n47682 ; n47683
g45248 and pi0813 n47073 ; n47684
g45249 and n47119 n47684 ; n47685
g45250 nor n47683 n47685 ; n47686
g45251 and n47679 n47686_not ; n47687
g45252 nor n47677 n47687 ; n47688
g45253 nor n7643 n47688 ; n47689
g45254 or n47670 n47689 ; po0842
g45255 and pi1113_not po0980 ; n47691
g45256 and pi0686 po0980_not ; n47692
g45257 nor pi0962 n47691 ; n47693
g45258 and n47692_not n47693 ; po0843
g45259 nor pi0687 po0980 ; n47695
g45260 and pi1127_not po0980 ; n47696
g45261 nor pi0962 n47695 ; n47697
g45262 and n47696_not n47697 ; po0844
g45263 and pi1115_not po0980 ; n47699
g45264 and pi0688 po0980_not ; n47700
g45265 nor pi0962 n47699 ; n47701
g45266 and n47700_not n47701 ; po0845
g45267 and pi0351 n47651 ; n47703
g45268 and pi0376 n47103 ; n47704
g45269 nor n47703 n47704 ; n47705
g45270 nor pi0591 n47705 ; n47706
g45271 and pi0401 pi0592_not ; n47707
g45272 and n47101 n47707 ; n47708
g45273 nor n47706 n47708 ; n47709
g45274 nor pi0588 n47709 ; n47710
g45275 and pi0426 n47660 ; n47711
g45276 and n47661 n47711 ; n47712
g45277 nor n47710 n47712 ; n47713
g45278 and n47050 n47713_not ; n47714
g45279 and pi0199 pi1079_not ; n47715
g45280 and pi0199_not n42849 ; n47716
g45281 nor n47050 n47715 ; n47717
g45282 and n47716_not n47717 ; n47718
g45283 nor n47714 n47718 ; n47719
g45284 and n7643 n47719_not ; n47720
g45285 and pi0798 n47119 ; n47721
g45286 nor pi0658 pi1135 ; n47722
g45287 and pi0655 pi1135 ; n47723
g45288 and pi1136 n47722_not ; n47724
g45289 and n47723_not n47724 ; n47725
g45290 nor n47721 n47725 ; n47726
g45291 and n47074 n47726_not ; n47727
g45292 and pi0752 n47086 ; n47728
g45293 and pi0703_not pi1135 ; n47729
g45294 nor pi0843 pi1136 ; n47730
g45295 nor n47729 n47730 ; n47731
g45296 and n47092 n47731 ; n47732
g45297 and n47728_not n47732 ; n47733
g45298 nor n47727 n47733 ; n47734
g45299 nor n7643 n47734 ; n47735
g45300 or n47720 n47735 ; po0846
g45301 nor pi0690 po0980 ; n47737
g45302 and pi1108_not po0980 ; n47738
g45303 nor pi0962 n47737 ; n47739
g45304 and n47738_not n47739 ; po0847
g45305 nor pi0691 po0980 ; n47741
g45306 and pi1107_not po0980 ; n47742
g45307 nor pi0962 n47741 ; n47743
g45308 and n47742_not n47743 ; po0848
g45309 and pi0352 n47651 ; n47745
g45310 and pi0317 n47103 ; n47746
g45311 nor n47745 n47746 ; n47747
g45312 nor pi0591 n47747 ; n47748
g45313 and pi0402 pi0592_not ; n47749
g45314 and n47101 n47749 ; n47750
g45315 nor n47748 n47750 ; n47751
g45316 nor pi0588 n47751 ; n47752
g45317 and pi0427 n47660 ; n47753
g45318 and n47661 n47753 ; n47754
g45319 nor n47752 n47754 ; n47755
g45320 and n47050 n47755_not ; n47756
g45321 and pi0199 pi1078_not ; n47757
g45322 and pi0199_not n42861 ; n47758
g45323 nor n47050 n47757 ; n47759
g45324 and n47758_not n47759 ; n47760
g45325 nor n47756 n47760 ; n47761
g45326 and n7643 n47761_not ; n47762
g45327 and pi0844 n47119 ; n47763
g45328 and pi0726_not pi1135 ; n47764
g45329 and pi0770 pi1135_not ; n47765
g45330 and pi1136 n47764_not ; n47766
g45331 and n47765_not n47766 ; n47767
g45332 and pi1134 n47763_not ; n47768
g45333 and n47767_not n47768 ; n47769
g45334 and pi0801 n47119 ; n47770
g45335 nor pi0656 pi1135 ; n47771
g45336 and pi0649 pi1135 ; n47772
g45337 and pi1136 n47771_not ; n47773
g45338 and n47772_not n47773 ; n47774
g45339 nor pi1134 n47770 ; n47775
g45340 and n47774_not n47775 ; n47776
g45341 and n47127 n47769_not ; n47777
g45342 and n47776_not n47777 ; n47778
g45343 or n47762 n47778 ; po0849
g45344 and pi1129_not po0954 ; n47780
g45345 and pi0693 po0954_not ; n47781
g45346 nor pi0962 n47780 ; n47782
g45347 and n47781_not n47782 ; po0850
g45348 and pi1128_not po0980 ; n47784
g45349 and pi0694 po0980_not ; n47785
g45350 nor pi0962 n47784 ; n47786
g45351 and n47785_not n47786 ; po0851
g45352 and pi1111_not po0954 ; n47788
g45353 and pi0695 po0954_not ; n47789
g45354 nor pi0962 n47788 ; n47790
g45355 and n47789_not n47790 ; po0852
g45356 nor pi0696 po0980 ; n47792
g45357 and pi1100_not po0980 ; n47793
g45358 nor pi0962 n47792 ; n47794
g45359 and n47793_not n47794 ; po0853
g45360 and pi1129_not po0980 ; n47796
g45361 and pi0697 po0980_not ; n47797
g45362 nor pi0962 n47796 ; n47798
g45363 and n47797_not n47798 ; po0854
g45364 and pi1116_not po0980 ; n47800
g45365 and pi0698 po0980_not ; n47801
g45366 nor pi0962 n47800 ; n47802
g45367 and n47801_not n47802 ; po0855
g45368 nor pi0699 po0980 ; n47804
g45369 and pi1103_not po0980 ; n47805
g45370 nor pi0962 n47804 ; n47806
g45371 and n47805_not n47806 ; po0856
g45372 nor pi0700 po0980 ; n47808
g45373 and pi1110_not po0980 ; n47809
g45374 nor pi0962 n47808 ; n47810
g45375 and n47809_not n47810 ; po0857
g45376 and pi1123_not po0980 ; n47812
g45377 and pi0701 po0980_not ; n47813
g45378 nor pi0962 n47812 ; n47814
g45379 and n47813_not n47814 ; po0858
g45380 and pi1117_not po0980 ; n47816
g45381 and pi0702 po0980_not ; n47817
g45382 nor pi0962 n47816 ; n47818
g45383 and n47817_not n47818 ; po0859
g45384 nor pi0703 po0980 ; n47820
g45385 and pi1124_not po0980 ; n47821
g45386 nor pi0962 n47820 ; n47822
g45387 and n47821_not n47822 ; po0860
g45388 and pi1112_not po0980 ; n47824
g45389 and pi0704 po0980_not ; n47825
g45390 nor pi0962 n47824 ; n47826
g45391 and n47825_not n47826 ; po0861
g45392 nor pi0705 po0980 ; n47828
g45393 and pi1125_not po0980 ; n47829
g45394 nor pi0962 n47828 ; n47830
g45395 and n47829_not n47830 ; po0862
g45396 nor pi0706 po0980 ; n47832
g45397 and pi1105_not po0980 ; n47833
g45398 nor pi0962 n47832 ; n47834
g45399 and n47833_not n47834 ; po0863
g45400 and pi0370 n47058 ; n47836
g45401 and pi0395 pi0591 ; n47837
g45402 and pi0592_not n47837 ; n47838
g45403 nor n47836 n47838 ; n47839
g45404 nor pi0590 n47839 ; n47840
g45405 and pi0347 n47065 ; n47841
g45406 nor n47840 n47841 ; n47842
g45407 and pi0588_not n47050 ; n47843
g45408 and n47842_not n47843 ; n47844
g45409 and pi0199 pi1055_not ; n47845
g45410 nor pi0200 pi0304 ; n47846
g45411 and pi0200 pi1048_not ; n47847
g45412 nor n47846 n47847 ; n47848
g45413 nor pi0199 n47848 ; n47849
g45414 nor n47050 n47845 ; n47850
g45415 and n47849_not n47850 ; n47851
g45416 and n47050 n47055 ; n47852
g45417 and pi0420 pi0588 ; n47853
g45418 and n47852 n47853 ; n47854
g45419 nor n47851 n47854 ; n47855
g45420 and n47844_not n47855 ; n47856
g45421 and n7643 n47856_not ; n47857
g45422 and pi0627_not pi1135 ; n47858
g45423 nor pi0618 pi1135 ; n47859
g45424 nor pi1134 n47858 ; n47860
g45425 and n47859_not n47860 ; n47861
g45426 and n47283 n47861 ; n47862
g45427 and pi0702 pi1135 ; n47863
g45428 nor pi0847 pi1136 ; n47864
g45429 and pi0753 n47086 ; n47865
g45430 nor n47863 n47864 ; n47866
g45431 and n47092 n47866 ; n47867
g45432 and n47865_not n47867 ; n47868
g45433 nor n47862 n47868 ; n47869
g45434 nor n7643 n47869 ; n47870
g45435 or n47857 n47870 ; po0864
g45436 and n47050 n47660 ; n47872
g45437 and pi0459 n47661 ; n47873
g45438 and n47872 n47873 ; n47874
g45439 and n47050 n47058 ; n47875
g45440 and pi0442 n47875 ; n47876
g45441 and pi0592_not n47050 ; n47877
g45442 and pi0328 pi0591 ; n47878
g45443 and n47877 n47878 ; n47879
g45444 nor n47876 n47879 ; n47880
g45445 nor pi0590 n47880 ; n47881
g45446 and pi0321 n47050 ; n47882
g45447 and n47065 n47882 ; n47883
g45448 nor n47881 n47883 ; n47884
g45449 nor pi0588 n47884 ; n47885
g45450 and pi0199 pi1058_not ; n47886
g45451 nor pi0200 pi0305 ; n47887
g45452 and pi0200 pi1084_not ; n47888
g45453 nor n47887 n47888 ; n47889
g45454 nor pi0199 n47889 ; n47890
g45455 nor n47050 n47886 ; n47891
g45456 and n47890_not n47891 ; n47892
g45457 and n7643 n47874_not ; n47893
g45458 and n47892_not n47893 ; n47894
g45459 and n47885_not n47894 ; n47895
g45460 nor pi0609 pi1135 ; n47896
g45461 and pi0660_not pi1135 ; n47897
g45462 nor pi1134 n47896 ; n47898
g45463 and n47897_not n47898 ; n47899
g45464 and n47283 n47899 ; n47900
g45465 and n47073 n47090_not ; n47901
g45466 and pi0709 pi1135 ; n47902
g45467 nor pi0857 pi1136 ; n47903
g45468 and pi0754 n47086 ; n47904
g45469 and pi1134 n47902_not ; n47905
g45470 and n47903_not n47905 ; n47906
g45471 and n47901 n47906 ; n47907
g45472 and n47904_not n47907 ; n47908
g45473 nor n7643 n47900 ; n47909
g45474 and n47908_not n47909 ; n47910
g45475 nor n47895 n47910 ; po0865
g45476 and pi1118_not po0980 ; n47912
g45477 and pi0709 po0980_not ; n47913
g45478 nor pi0962 n47912 ; n47914
g45479 and n47913_not n47914 ; po0866
g45480 nor pi0710 po0954 ; n47916
g45481 and pi1106_not po0954 ; n47917
g45482 nor pi0962 n47916 ; n47918
g45483 and n47917_not n47918 ; po0867
g45484 and pi0373 n47058 ; n47920
g45485 and pi0398 pi0591 ; n47921
g45486 and pi0592_not n47921 ; n47922
g45487 nor n47920 n47922 ; n47923
g45488 nor pi0590 n47923 ; n47924
g45489 and pi0348 n47065 ; n47925
g45490 nor n47924 n47925 ; n47926
g45491 and n47843 n47926_not ; n47927
g45492 and pi0199 pi1087_not ; n47928
g45493 nor pi0200 pi0306 ; n47929
g45494 and pi0200 pi1059_not ; n47930
g45495 nor n47929 n47930 ; n47931
g45496 nor pi0199 n47931 ; n47932
g45497 nor n47050 n47928 ; n47933
g45498 and n47932_not n47933 ; n47934
g45499 and pi0423 pi0588 ; n47935
g45500 and n47852 n47935 ; n47936
g45501 nor n47934 n47936 ; n47937
g45502 and n47927_not n47937 ; n47938
g45503 and n7643 n47938_not ; n47939
g45504 and pi0647_not pi1135 ; n47940
g45505 nor pi0630 pi1135 ; n47941
g45506 nor pi1134 n47940 ; n47942
g45507 and n47941_not n47942 ; n47943
g45508 and n47283 n47943 ; n47944
g45509 and pi0725 pi1135 ; n47945
g45510 nor pi0858 pi1136 ; n47946
g45511 and pi0755 n47086 ; n47947
g45512 nor n47945 n47946 ; n47948
g45513 and n47092 n47948 ; n47949
g45514 and n47947_not n47949 ; n47950
g45515 nor n47944 n47950 ; n47951
g45516 nor n7643 n47951 ; n47952
g45517 or n47939 n47952 ; po0868
g45518 and pi0701 pi1135 ; n47954
g45519 nor pi0842 pi1136 ; n47955
g45520 and pi0751 n47086 ; n47956
g45521 and pi1134 n47954_not ; n47957
g45522 and n47955_not n47957 ; n47958
g45523 and n47901 n47958 ; n47959
g45524 and n47956_not n47959 ; n47960
g45525 and pi0715_not pi1135 ; n47961
g45526 nor pi0644 pi1135 ; n47962
g45527 nor pi1134 n47961 ; n47963
g45528 and n47962_not n47963 ; n47964
g45529 and n47283 n47964 ; n47965
g45530 nor n47960 n47965 ; n47966
g45531 nor n7643 n47966 ; n47967
g45532 and pi0199 pi1035 ; n47968
g45533 and pi0298 n10809 ; n47969
g45534 and pi1044 n11444 ; n47970
g45535 nor n47050 n47968 ; n47971
g45536 and n47969_not n47971 ; n47972
g45537 and n47970_not n47972 ; n47973
g45538 and pi0425 n47660 ; n47974
g45539 and n47661 n47974 ; n47975
g45540 and pi0374 n47058 ; n47976
g45541 and pi0400 pi0591 ; n47977
g45542 and pi0592_not n47977 ; n47978
g45543 nor n47976 n47978 ; n47979
g45544 nor pi0590 n47979 ; n47980
g45545 and pi0350 n47065 ; n47981
g45546 nor n47980 n47981 ; n47982
g45547 nor pi0588 n47982 ; n47983
g45548 and n47050 n47975_not ; n47984
g45549 and n47983_not n47984 ; n47985
g45550 and n7643 n47973_not ; n47986
g45551 and n47985_not n47986 ; n47987
g45552 or n47967 n47987 ; po0869
g45553 and pi0371 n47058 ; n47989
g45554 and pi0396 pi0591 ; n47990
g45555 and pi0592_not n47990 ; n47991
g45556 nor n47989 n47991 ; n47992
g45557 nor pi0590 n47992 ; n47993
g45558 and pi0322 n47065 ; n47994
g45559 nor n47993 n47994 ; n47995
g45560 and n47843 n47995_not ; n47996
g45561 and pi0199 pi1051_not ; n47997
g45562 nor pi0200 pi0309 ; n47998
g45563 and pi0200 pi1072_not ; n47999
g45564 nor n47998 n47999 ; n48000
g45565 nor pi0199 n48000 ; n48001
g45566 nor n47050 n47997 ; n48002
g45567 and n48001_not n48002 ; n48003
g45568 and pi0421 pi0588 ; n48004
g45569 and n47852 n48004 ; n48005
g45570 nor n48003 n48005 ; n48006
g45571 and n47996_not n48006 ; n48007
g45572 and n7643 n48007_not ; n48008
g45573 and pi0628_not pi1135 ; n48009
g45574 nor pi0629 pi1135 ; n48010
g45575 nor pi1134 n48009 ; n48011
g45576 and n48010_not n48011 ; n48012
g45577 and n47283 n48012 ; n48013
g45578 and pi0734 pi1135 ; n48014
g45579 nor pi0854 pi1136 ; n48015
g45580 and pi0756 n47086 ; n48016
g45581 nor n48014 n48015 ; n48017
g45582 and n47092 n48017 ; n48018
g45583 and n48016_not n48018 ; n48019
g45584 nor n48013 n48019 ; n48020
g45585 nor n7643 n48020 ; n48021
g45586 or n48008 n48021 ; po0870
g45587 and pi0461 n47651 ; n48023
g45588 and pi0439 n47103 ; n48024
g45589 nor n48023 n48024 ; n48025
g45590 nor pi0591 n48025 ; n48026
g45591 and pi0326 pi0592_not ; n48027
g45592 and n47101 n48027 ; n48028
g45593 nor n48026 n48028 ; n48029
g45594 nor pi0588 n48029 ; n48030
g45595 and pi0449 n47660 ; n48031
g45596 and n47661 n48031 ; n48032
g45597 nor n48030 n48032 ; n48033
g45598 and n47050 n48033_not ; n48034
g45599 and pi0199 pi1057_not ; n48035
g45600 nor n47050 n48035 ; n48036
g45601 and n42339_not n48036 ; n48037
g45602 nor n48034 n48037 ; n48038
g45603 and n7643 n48038_not ; n48039
g45604 and pi0867 n47119 ; n48040
g45605 and pi0762 pi1135_not ; n48041
g45606 and pi0697 pi1135 ; n48042
g45607 and pi1136 n48041_not ; n48043
g45608 and n48042_not n48043 ; n48044
g45609 nor n48040 n48044 ; n48045
g45610 and n47091 n48045_not ; n48046
g45611 nor pi0653 pi1135 ; n48047
g45612 and pi0693 pi1135 ; n48048
g45613 and pi1136 n48047_not ; n48049
g45614 and n48048_not n48049 ; n48050
g45615 and pi0816 n47073 ; n48051
g45616 and n47119 n48051 ; n48052
g45617 nor n48050 n48052 ; n48053
g45618 and n47679 n48053_not ; n48054
g45619 nor n48046 n48054 ; n48055
g45620 nor n7643 n48055 ; n48056
g45621 or n48039 n48056 ; po0871
g45622 nor pi0715 po0954 ; n48058
g45623 and pi1123_not po0954 ; n48059
g45624 nor pi0962 n48058 ; n48060
g45625 and n48059_not n48060 ; po0872
g45626 and pi0454 n47661 ; n48062
g45627 and n47872 n48062 ; n48063
g45628 and pi0440 n47875 ; n48064
g45629 and pi0329 pi0591 ; n48065
g45630 and n47877 n48065 ; n48066
g45631 nor n48064 n48066 ; n48067
g45632 nor pi0590 n48067 ; n48068
g45633 and pi0349 n47050 ; n48069
g45634 and n47065 n48069 ; n48070
g45635 nor n48068 n48070 ; n48071
g45636 nor pi0588 n48071 ; n48072
g45637 and pi0199 pi1043_not ; n48073
g45638 nor pi0200 pi0307 ; n48074
g45639 and pi0200 pi1053_not ; n48075
g45640 nor n48074 n48075 ; n48076
g45641 nor pi0199 n48076 ; n48077
g45642 nor n47050 n48073 ; n48078
g45643 and n48077_not n48078 ; n48079
g45644 and n7643 n48063_not ; n48080
g45645 and n48079_not n48080 ; n48081
g45646 and n48072_not n48081 ; n48082
g45647 nor pi0626 pi1135 ; n48083
g45648 and pi0641_not pi1135 ; n48084
g45649 nor pi1134 n48083 ; n48085
g45650 and n48084_not n48085 ; n48086
g45651 and n47283 n48086 ; n48087
g45652 and pi0738 pi1135 ; n48088
g45653 nor pi0845 pi1136 ; n48089
g45654 and pi0761 n47086 ; n48090
g45655 and pi1134 n48088_not ; n48091
g45656 and n48089_not n48091 ; n48092
g45657 and n47901 n48092 ; n48093
g45658 and n48090_not n48093 ; n48094
g45659 nor n7643 n48087 ; n48095
g45660 and n48094_not n48095 ; n48096
g45661 nor n48082 n48096 ; po0873
g45662 and pi0318 pi0591 ; n48098
g45663 and pi0592_not n48098 ; n48099
g45664 and pi0591_not n8468 ; n48100
g45665 nor n48099 n48100 ; n48101
g45666 nor pi0590 n48101 ; n48102
g45667 and pi0462 n47065 ; n48103
g45668 nor n48102 n48103 ; n48104
g45669 and n47843 n48104_not ; n48105
g45670 and pi0199 pi1074_not ; n48106
g45671 and pi0199_not n42855 ; n48107
g45672 nor n47050 n48106 ; n48108
g45673 and n48107_not n48108 ; n48109
g45674 and pi0448 pi0588 ; n48110
g45675 and n47852 n48110 ; n48111
g45676 nor n48109 n48111 ; n48112
g45677 and n48105_not n48112 ; n48113
g45678 and n7643 n48113_not ; n48114
g45679 and pi0705_not pi1135 ; n48115
g45680 and pi0768 n47086 ; n48116
g45681 nor pi0839 pi1136 ; n48117
g45682 and pi1134 n48115_not ; n48118
g45683 and n48117_not n48118 ; n48119
g45684 and n47901 n48119 ; n48120
g45685 and n48116_not n48120 ; n48121
g45686 and pi0800 n47119 ; n48122
g45687 nor pi0645 pi1135 ; n48123
g45688 and pi0669 pi1135 ; n48124
g45689 and pi1136 n48123_not ; n48125
g45690 and n48124_not n48125 ; n48126
g45691 nor n48122 n48126 ; n48127
g45692 and n47074 n48127_not ; n48128
g45693 nor n48121 n48128 ; n48129
g45694 nor n7643 n48129 ; n48130
g45695 or n48114 n48130 ; po0874
g45696 and pi0419 n47661 ; n48132
g45697 and n47872 n48132 ; n48133
g45698 and pi0369 n47875 ; n48134
g45699 and pi0394 pi0591 ; n48135
g45700 and n47877 n48135 ; n48136
g45701 nor n48134 n48136 ; n48137
g45702 nor pi0590 n48137 ; n48138
g45703 and pi0315 n47050 ; n48139
g45704 and n47065 n48139 ; n48140
g45705 nor n48138 n48140 ; n48141
g45706 nor pi0588 n48141 ; n48142
g45707 and pi0199 pi1080_not ; n48143
g45708 nor pi0200 pi0303 ; n48144
g45709 and pi0200 pi1049_not ; n48145
g45710 nor n48144 n48145 ; n48146
g45711 nor pi0199 n48146 ; n48147
g45712 nor n47050 n48143 ; n48148
g45713 and n48147_not n48148 ; n48149
g45714 and n7643 n48133_not ; n48150
g45715 and n48149_not n48150 ; n48151
g45716 and n48142_not n48151 ; n48152
g45717 nor pi0608 pi1135 ; n48153
g45718 and pi0625_not pi1135 ; n48154
g45719 nor pi1134 n48153 ; n48155
g45720 and n48154_not n48155 ; n48156
g45721 and n47283 n48156 ; n48157
g45722 and pi0698 pi1135 ; n48158
g45723 nor pi0853 pi1136 ; n48159
g45724 and pi0767 n47086 ; n48160
g45725 and pi1134 n48158_not ; n48161
g45726 and n48159_not n48161 ; n48162
g45727 and n47901 n48162 ; n48163
g45728 and n48160_not n48163 ; n48164
g45729 nor n7643 n48157 ; n48165
g45730 and n48164_not n48165 ; n48166
g45731 nor n48152 n48166 ; po0875
g45732 and pi0378 n47058 ; n48168
g45733 and pi0325 pi0591 ; n48169
g45734 and pi0592_not n48169 ; n48170
g45735 nor n48168 n48170 ; n48171
g45736 nor pi0590 n48171 ; n48172
g45737 and pi0353 n47065 ; n48173
g45738 nor n48172 n48173 ; n48174
g45739 and n47843 n48174_not ; n48175
g45740 and pi0199 pi1063_not ; n48176
g45741 and pi0199_not n42867 ; n48177
g45742 nor n47050 n48176 ; n48178
g45743 and n48177_not n48178 ; n48179
g45744 and pi0451 pi0588 ; n48180
g45745 and n47852 n48180 ; n48181
g45746 nor n48179 n48181 ; n48182
g45747 and n48175_not n48182 ; n48183
g45748 and n7643 n48183_not ; n48184
g45749 and pi0687_not pi1135 ; n48185
g45750 and pi0774 n47086 ; n48186
g45751 nor pi0868 pi1136 ; n48187
g45752 and pi1134 n48185_not ; n48188
g45753 and n48187_not n48188 ; n48189
g45754 and n47901 n48189 ; n48190
g45755 and n48186_not n48190 ; n48191
g45756 and pi0807 n47119 ; n48192
g45757 nor pi0636 pi1135 ; n48193
g45758 and pi0650 pi1135 ; n48194
g45759 and pi1136 n48193_not ; n48195
g45760 and n48194_not n48195 ; n48196
g45761 nor n48192 n48196 ; n48197
g45762 and n47074 n48197_not ; n48198
g45763 nor n48191 n48198 ; n48199
g45764 nor n7643 n48199 ; n48200
g45765 or n48184 n48200 ; po0876
g45766 and pi0356 n47651 ; n48202
g45767 and pi0381 n47103 ; n48203
g45768 nor n48202 n48203 ; n48204
g45769 nor pi0591 n48204 ; n48205
g45770 and pi0405 pi0592_not ; n48206
g45771 and n47101 n48206 ; n48207
g45772 nor n48205 n48207 ; n48208
g45773 nor pi0588 n48208 ; n48209
g45774 and pi0445 n47660 ; n48210
g45775 and n47661 n48210 ; n48211
g45776 nor n48209 n48211 ; n48212
g45777 and n47050 n48212_not ; n48213
g45778 and pi0199 pi1081_not ; n48214
g45779 nor n47050 n48214 ; n48215
g45780 and n42887_not n48215 ; n48216
g45781 nor n48213 n48216 ; n48217
g45782 and n7643 n48217_not ; n48218
g45783 and pi0880 n47119 ; n48219
g45784 and pi0750 pi1135_not ; n48220
g45785 and pi0684 pi1135 ; n48221
g45786 and pi1136 n48220_not ; n48222
g45787 and n48221_not n48222 ; n48223
g45788 nor n48219 n48223 ; n48224
g45789 and n47091 n48224_not ; n48225
g45790 nor pi0651 pi1135 ; n48226
g45791 and pi0654 pi1135 ; n48227
g45792 and pi1136 n48226_not ; n48228
g45793 and n48227_not n48228 ; n48229
g45794 and pi0794 n47073 ; n48230
g45795 and n47119 n48230 ; n48231
g45796 nor n48229 n48231 ; n48232
g45797 and n47679 n48232_not ; n48233
g45798 nor n48225 n48233 ; n48234
g45799 nor n7643 n48234 ; n48235
g45800 or n48218 n48235 ; po0877
g45801 and pi0721 pi0775_not ; n48237
g45802 and pi0721 pi0813 ; n48238
g45803 nor pi0773 pi0801 ; n48239
g45804 and pi0773 pi0801 ; n48240
g45805 nor n48239 n48240 ; n48241
g45806 nor pi0771 pi0800 ; n48242
g45807 and pi0771 pi0800 ; n48243
g45808 nor n48242 n48243 ; n48244
g45809 nor pi0769 pi0794 ; n48245
g45810 and pi0769 pi0794 ; n48246
g45811 nor n48245 n48246 ; n48247
g45812 nor pi0765 pi0798 ; n48248
g45813 and pi0765 pi0798 ; n48249
g45814 nor n48248 n48249 ; n48250
g45815 and pi0807 n48250_not ; n48251
g45816 and pi0747 n48251 ; n48252
g45817 nor pi0747 pi0807 ; n48253
g45818 and n48250_not n48253 ; n48254
g45819 nor n48252 n48254 ; n48255
g45820 nor n48247 n48255 ; n48256
g45821 and n48244_not n48256 ; n48257
g45822 and n48241_not n48257 ; n48258
g45823 and n48238 n48258 ; n48259
g45824 nor pi0775 pi0816 ; n48260
g45825 and pi0775 pi0816 ; n48261
g45826 nor n48260 n48261 ; n48262
g45827 and n48259 n48262_not ; n48263
g45828 and n48237 n48263_not ; n48264
g45829 and pi0747 pi0773 ; n48265
g45830 and pi0769 n48265 ; n48266
g45831 and pi0721 n48266 ; n48267
g45832 nor pi0721 n48266 ; n48268
g45833 and pi0775 n48267_not ; n48269
g45834 and n48268_not n48269 ; n48270
g45835 and n48244_not n48251 ; n48271
g45836 nor pi0721 pi0813 ; n48272
g45837 and pi0794 pi0801 ; n48273
g45838 and n48272 n48273 ; n48274
g45839 and n48271 n48274 ; n48275
g45840 nor n48259 n48275 ; n48276
g45841 and pi0816 n48276_not ; n48277
g45842 and n48270 n48277_not ; n48278
g45843 and pi0795 n48278_not ; n48279
g45844 and pi0945_not pi0988 ; n48280
g45845 and pi0731 n48280 ; n48281
g45846 nor n48237 n48270 ; n48282
g45847 and n48281 n48282_not ; n48283
g45848 and n48279_not n48283 ; n48284
g45849 nor pi0731 pi0795 ; n48285
g45850 and pi0731 pi0795 ; n48286
g45851 nor n48285 n48286 ; n48287
g45852 and n48263 n48287_not ; n48288
g45853 and pi0721 n48281_not ; n48289
g45854 and n48288_not n48289 ; n48290
g45855 nor n48264 n48290 ; n48291
g45856 nand n48284_not n48291 ; po0878
g45857 and pi0379 n47058 ; n48293
g45858 and pi0403 pi0591 ; n48294
g45859 and pi0592_not n48294 ; n48295
g45860 nor n48293 n48295 ; n48296
g45861 nor pi0590 n48296 ; n48297
g45862 and pi0354 n47065 ; n48298
g45863 nor n48297 n48298 ; n48299
g45864 and n47843 n48299_not ; n48300
g45865 and pi0199 pi1045_not ; n48301
g45866 and pi0199_not n42873 ; n48302
g45867 nor n47050 n48301 ; n48303
g45868 and n48302_not n48303 ; n48304
g45869 and pi0428 pi0588 ; n48305
g45870 and n47852 n48305 ; n48306
g45871 nor n48304 n48306 ; n48307
g45872 and n48300_not n48307 ; n48308
g45873 and n7643 n48308_not ; n48309
g45874 nor pi0795 pi1134 ; n48310
g45875 and pi0851_not pi1134 ; n48311
g45876 nor pi1136 n48310 ; n48312
g45877 and n48311_not n48312 ; n48313
g45878 nor pi0640 pi1134 ; n48314
g45879 and pi0776 pi1134 ; n48315
g45880 and pi1136 n48314_not ; n48316
g45881 and n48315_not n48316 ; n48317
g45882 nor n48313 n48317 ; n48318
g45883 nor pi1135 n48318 ; n48319
g45884 and pi0694 pi1134 ; n48320
g45885 and pi0732 pi1134_not ; n48321
g45886 and pi1135 pi1136 ; n48322
g45887 and n48320_not n48322 ; n48323
g45888 and n48321_not n48323 ; n48324
g45889 nor n48319 n48324 ; n48325
g45890 and n47127 n48325_not ; n48326
g45891 or n48309 n48326 ; po0879
g45892 and pi1111_not po0980 ; n48328
g45893 and pi0723 po0980_not ; n48329
g45894 nor pi0962 n48328 ; n48330
g45895 and n48329_not n48330 ; po0880
g45896 and pi1114_not po0980 ; n48332
g45897 and pi0724 po0980_not ; n48333
g45898 nor pi0962 n48332 ; n48334
g45899 and n48333_not n48334 ; po0881
g45900 and pi1120_not po0980 ; n48336
g45901 and pi0725 po0980_not ; n48337
g45902 nor pi0962 n48336 ; n48338
g45903 and n48337_not n48338 ; po0882
g45904 nor pi0726 po0980 ; n48340
g45905 and pi1126_not po0980 ; n48341
g45906 nor pi0962 n48340 ; n48342
g45907 and n48341_not n48342 ; po0883
g45908 nor pi0727 po0980 ; n48344
g45909 and pi1102_not po0980 ; n48345
g45910 nor pi0962 n48344 ; n48346
g45911 and n48345_not n48346 ; po0884
g45912 and pi1131_not po0980 ; n48348
g45913 and pi0728 po0980_not ; n48349
g45914 nor pi0962 n48348 ; n48350
g45915 and n48349_not n48350 ; po0885
g45916 nor pi0729 po0980 ; n48352
g45917 and pi1104_not po0980 ; n48353
g45918 nor pi0962 n48352 ; n48354
g45919 and n48353_not n48354 ; po0886
g45920 nor pi0730 po0980 ; n48356
g45921 and pi1106_not po0980 ; n48357
g45922 nor pi0962 n48356 ; n48358
g45923 and n48357_not n48358 ; po0887
g45924 nor n48238 n48272 ; n48360
g45925 and n48258 n48360_not ; n48361
g45926 and pi0795 n48262_not ; n48362
g45927 and n48361 n48362 ; n48363
g45928 nor n48265 n48363 ; n48364
g45929 and n48281 n48364_not ; n48365
g45930 and pi0731 n48363_not ; n48366
g45931 nor n48262 n48360 ; n48367
g45932 and pi0795_not pi0801 ; n48368
g45933 and n48247_not n48368 ; n48369
g45934 and n48367 n48369 ; n48370
g45935 and n48271 n48370 ; n48371
g45936 and n48265 n48371_not ; n48372
g45937 nor pi0731 n48372 ; n48373
g45938 and n48280 n48373_not ; n48374
g45939 nor n48366 n48374 ; n48375
g45940 nor n48365 n48375 ; po0888
g45941 and pi1128_not po0954 ; n48377
g45942 and pi0732 po0954_not ; n48378
g45943 nor pi0962 n48377 ; n48379
g45944 and n48378_not n48379 ; po0889
g45945 and pi0424 n47661 ; n48381
g45946 and n47872 n48381 ; n48382
g45947 and pi0375 n47875 ; n48383
g45948 and pi0399 pi0591 ; n48384
g45949 and n47877 n48384 ; n48385
g45950 nor n48383 n48385 ; n48386
g45951 nor pi0590 n48386 ; n48387
g45952 and pi0316 n47050 ; n48388
g45953 and n47065 n48388 ; n48389
g45954 nor n48387 n48389 ; n48390
g45955 nor pi0588 n48390 ; n48391
g45956 and pi0199 pi1047_not ; n48392
g45957 nor pi0200 pi0308 ; n48393
g45958 and pi0200 pi1037_not ; n48394
g45959 nor n48393 n48394 ; n48395
g45960 nor pi0199 n48395 ; n48396
g45961 nor n47050 n48392 ; n48397
g45962 and n48396_not n48397 ; n48398
g45963 and n7643 n48382_not ; n48399
g45964 and n48398_not n48399 ; n48400
g45965 and n48391_not n48400 ; n48401
g45966 nor pi0619 pi1135 ; n48402
g45967 and pi0648_not pi1135 ; n48403
g45968 nor pi1134 n48402 ; n48404
g45969 and n48403_not n48404 ; n48405
g45970 and n47283 n48405 ; n48406
g45971 and pi0737 pi1135 ; n48407
g45972 nor pi0838 pi1136 ; n48408
g45973 and pi0777 n47086 ; n48409
g45974 and pi1134 n48407_not ; n48410
g45975 and n48408_not n48410 ; n48411
g45976 and n47901 n48411 ; n48412
g45977 and n48409_not n48412 ; n48413
g45978 nor n7643 n48406 ; n48414
g45979 and n48413_not n48414 ; n48415
g45980 nor n48401 n48415 ; po0890
g45981 and pi1119_not po0980 ; n48417
g45982 and pi0734 po0980_not ; n48418
g45983 nor pi0962 n48417 ; n48419
g45984 and n48418_not n48419 ; po0891
g45985 nor pi0735 po0980 ; n48421
g45986 and pi1109_not po0980 ; n48422
g45987 nor pi0962 n48421 ; n48423
g45988 and n48422_not n48423 ; po0892
g45989 nor pi0736 po0980 ; n48425
g45990 and pi1101_not po0980 ; n48426
g45991 nor pi0962 n48425 ; n48427
g45992 and n48426_not n48427 ; po0893
g45993 and pi1122_not po0980 ; n48429
g45994 and pi0737 po0980_not ; n48430
g45995 nor pi0962 n48429 ; n48431
g45996 and n48430_not n48431 ; po0894
g45997 and pi1121_not po0980 ; n48433
g45998 and pi0738 po0980_not ; n48434
g45999 nor pi0962 n48433 ; n48435
g46000 and n48434_not n48435 ; po0895
g46001 nor pi0952 pi1061 ; n48437
g46002 and n46780 n48437 ; n48438
g46003 and pi0832 n48438 ; po0988
g46004 and pi1108 po0988 ; n48440
g46005 and pi0739 po0988_not ; n48441
g46006 nor pi0966 n48440 ; n48442
g46007 nand n48441_not n48442 ; po0896
g46008 nor pi0741 po0988 ; n48444
g46009 and pi1114 po0988 ; n48445
g46010 nor pi0966 n48444 ; n48446
g46011 nand n48445_not n48446 ; po0898
g46012 nor pi0742 po0988 ; n48448
g46013 and pi1112 po0988 ; n48449
g46014 nor pi0966 n48448 ; n48450
g46015 nand n48449_not n48450 ; po0899
g46016 and pi1109 po0988 ; n48452
g46017 and pi0743 po0988_not ; n48453
g46018 nor pi0966 n48452 ; n48454
g46019 nand n48453_not n48454 ; po0900
g46020 nor pi0744 po0988 ; n48456
g46021 and pi1131 po0988 ; n48457
g46022 nor pi0966 n48456 ; n48458
g46023 nand n48457_not n48458 ; po0901
g46024 nor pi0745 po0988 ; n48460
g46025 and pi1111 po0988 ; n48461
g46026 nor pi0966 n48460 ; n48462
g46027 nand n48461_not n48462 ; po0902
g46028 and pi1104 po0988 ; n48464
g46029 and pi0746 po0988_not ; n48465
g46030 nor pi0966 n48464 ; n48466
g46031 nand n48465_not n48466 ; po0903
g46032 and pi0773 n48280 ; n48468
g46033 nor pi0747 n48468 ; n48469
g46034 and n48265 n48280 ; n48470
g46035 and n48287_not n48367 ; n48471
g46036 and pi0801 n48254 ; n48472
g46037 nor n48241 n48468 ; n48473
g46038 and n48251 n48473 ; n48474
g46039 nor n48472 n48474 ; n48475
g46040 nor n48244 n48247 ; n48476
g46041 and n48471 n48476 ; n48477
g46042 and n48475_not n48477 ; n48478
g46043 nor n48469 n48470 ; n48479
g46044 and n48478_not n48479 ; po0904
g46045 and pi1106 po0988 ; n48481
g46046 and pi0748 po0988_not ; n48482
g46047 nor pi0966 n48481 ; n48483
g46048 nand n48482_not n48483 ; po0905
g46049 and pi1105 po0988 ; n48485
g46050 and pi0749 po0988_not ; n48486
g46051 nor pi0966 n48485 ; n48487
g46052 nand n48486_not n48487 ; po0906
g46053 nor pi0750 po0988 ; n48489
g46054 and pi1130 po0988 ; n48490
g46055 nor pi0966 n48489 ; n48491
g46056 nand n48490_not n48491 ; po0907
g46057 nor pi0751 po0988 ; n48493
g46058 and pi1123 po0988 ; n48494
g46059 nor pi0966 n48493 ; n48495
g46060 nand n48494_not n48495 ; po0908
g46061 nor pi0752 po0988 ; n48497
g46062 and pi1124 po0988 ; n48498
g46063 nor pi0966 n48497 ; n48499
g46064 nand n48498_not n48499 ; po0909
g46065 nor pi0753 po0988 ; n48501
g46066 and pi1117 po0988 ; n48502
g46067 nor pi0966 n48501 ; n48503
g46068 nand n48502_not n48503 ; po0910
g46069 nor pi0754 po0988 ; n48505
g46070 and pi1118 po0988 ; n48506
g46071 nor pi0966 n48505 ; n48507
g46072 nand n48506_not n48507 ; po0911
g46073 nor pi0755 po0988 ; n48509
g46074 and pi1120 po0988 ; n48510
g46075 nor pi0966 n48509 ; n48511
g46076 nand n48510_not n48511 ; po0912
g46077 nor pi0756 po0988 ; n48513
g46078 and pi1119 po0988 ; n48514
g46079 nor pi0966 n48513 ; n48515
g46080 nand n48514_not n48515 ; po0913
g46081 nor pi0757 po0988 ; n48517
g46082 and pi1113 po0988 ; n48518
g46083 nor pi0966 n48517 ; n48519
g46084 nand n48518_not n48519 ; po0914
g46085 and pi1101 po0988 ; n48521
g46086 and pi0758 po0988_not ; n48522
g46087 nor pi0966 n48521 ; n48523
g46088 nand n48522_not n48523 ; po0915
g46089 nor pi0759 po0988 ; n48525
g46090 and n46778 n48438 ; n48526
g46091 nor n48525 n48526 ; n48527
g46092 or pi0966 n48527 ; po0916
g46093 nor pi0760 po0988 ; n48529
g46094 and pi1115 po0988 ; n48530
g46095 nor pi0966 n48529 ; n48531
g46096 nand n48530_not n48531 ; po0917
g46097 nor pi0761 po0988 ; n48533
g46098 and pi1121 po0988 ; n48534
g46099 nor pi0966 n48533 ; n48535
g46100 nand n48534_not n48535 ; po0918
g46101 nor pi0762 po0988 ; n48537
g46102 and pi1129 po0988 ; n48538
g46103 nor pi0966 n48537 ; n48539
g46104 nand n48538_not n48539 ; po0919
g46105 and pi1103 po0988 ; n48541
g46106 and pi0763 po0988_not ; n48542
g46107 nor pi0966 n48541 ; n48543
g46108 nand n48542_not n48543 ; po0920
g46109 and pi1107 po0988 ; n48545
g46110 and pi0764 po0988_not ; n48546
g46111 nor pi0966 n48545 ; n48547
g46112 nand n48546_not n48547 ; po0921
g46113 and n48258 n48471 ; po0978
g46114 and pi0765 po0978_not ; n48550
g46115 and pi0945 n48550_not ; n48551
g46116 nor n48259 n48272 ; n48552
g46117 nor pi0765 n48243 ; n48553
g46118 and n48246_not n48553 ; n48554
g46119 and n48252_not n48554 ; n48555
g46120 and n48239 n48555_not ; n48556
g46121 nor n48240 n48556 ; n48557
g46122 and n48257 n48557_not ; n48558
g46123 nor pi0721 n48558 ; n48559
g46124 and n48260 n48559_not ; n48560
g46125 and n48552_not n48560 ; n48561
g46126 and n48261 n48361 ; n48562
g46127 nor pi0765 n48562 ; n48563
g46128 and n48561_not n48563 ; n48564
g46129 nor pi0795 n48564 ; n48565
g46130 nor pi0731 n48565 ; n48566
g46131 and pi0795_not n48566 ; n48567
g46132 and pi0765 n48567_not ; n48568
g46133 nor n48366 n48566 ; n48569
g46134 nor n48568 n48569 ; n48570
g46135 nor pi0945 n48570 ; n48571
g46136 nor n48551 n48571 ; po0922
g46137 and pi1110 po0988 ; n48573
g46138 and pi0766 po0988_not ; n48574
g46139 nor pi0966 n48573 ; n48575
g46140 nand n48574_not n48575 ; po0923
g46141 nor pi0767 po0988 ; n48577
g46142 and pi1116 po0988 ; n48578
g46143 nor pi0966 n48577 ; n48579
g46144 nand n48578_not n48579 ; po0924
g46145 nor pi0768 po0988 ; n48581
g46146 and pi1125 po0988 ; n48582
g46147 nor pi0966 n48581 ; n48583
g46148 nand n48582_not n48583 ; po0925
g46149 and pi0794 n48241_not ; n48585
g46150 and n48244_not n48585 ; n48586
g46151 and n48367 n48586 ; n48587
g46152 and n48255_not n48587 ; n48588
g46153 and pi0775_not n48588 ; n48589
g46154 nor n48562 n48589 ; n48590
g46155 and pi0795 n48590_not ; n48591
g46156 and pi0775 n48265 ; n48592
g46157 and pi0769 n48592_not ; n48593
g46158 and pi0769_not n48592 ; n48594
g46159 nor n48593 n48594 ; n48595
g46160 and n48281 n48595_not ; n48596
g46161 and n48591_not n48596 ; n48597
g46162 and n48287_not n48588 ; n48598
g46163 and pi0769 n48281_not ; n48599
g46164 and n48598_not n48599 ; n48600
g46165 or n48597 n48600 ; po0926
g46166 nor pi0770 po0988 ; n48602
g46167 and pi1126 po0988 ; n48603
g46168 nor pi0966 n48602 ; n48604
g46169 nand n48603_not n48604 ; po0927
g46170 nor n48261 n48560 ; n48606
g46171 and n48285 n48606_not ; n48607
g46172 and n48262_not n48286 ; n48608
g46173 nor n48607 n48608 ; n48609
g46174 and n48361 n48609_not ; po0963
g46175 and pi0945_not pi0987 ; n48611
g46176 and po0963_not n48611 ; n48612
g46177 and pi0771 pi0945 ; n48613
g46178 and po0978_not n48613 ; n48614
g46179 or n48612 n48614 ; po0928
g46180 and pi1102 po0988 ; n48616
g46181 and pi0772 po0988_not ; n48617
g46182 nor pi0966 n48616 ; n48618
g46183 nand n48617_not n48618 ; po0929
g46184 and pi0801_not n48257 ; n48620
g46185 and po0963 n48620 ; n48621
g46186 and n48280 n48621_not ; n48622
g46187 and pi0801 n48471_not ; n48623
g46188 and n48258 n48623_not ; n48624
g46189 and pi0773 n48624_not ; n48625
g46190 nor n48622 n48625 ; n48626
g46191 nor n48468 n48626 ; po0930
g46192 nor pi0774 po0988 ; n48628
g46193 and pi1127 po0988 ; n48629
g46194 nor pi0966 n48628 ; n48630
g46195 nand n48629_not n48630 ; po0931
g46196 and pi0775 po0978_not ; n48632
g46197 and pi0731 pi0945_not ; n48633
g46198 and pi0765 pi0771 ; n48634
g46199 and n48265 n48634 ; n48635
g46200 and pi0795 pi0800 ; n48636
g46201 and pi0801 pi0816_not ; n48637
g46202 and n48636 n48637 ; n48638
g46203 and n48360_not n48638 ; n48639
g46204 and n48256 n48639 ; n48640
g46205 and n48635 n48640_not ; n48641
g46206 nor pi0775 n48641 ; n48642
g46207 and n48633 n48642_not ; n48643
g46208 nor n48632 n48643 ; n48644
g46209 nor n48363 n48635 ; n48645
g46210 and pi0775 n48633 ; n48646
g46211 and n48645_not n48646 ; n48647
g46212 nor n48644 n48647 ; po0932
g46213 nor pi0776 po0988 ; n48649
g46214 and pi1128 po0988 ; n48650
g46215 nor pi0966 n48649 ; n48651
g46216 nand n48650_not n48651 ; po0933
g46217 nor pi0777 po0988 ; n48653
g46218 and pi1122 po0988 ; n48654
g46219 nor pi0966 n48653 ; n48655
g46220 nand n48654_not n48655 ; po0934
g46221 and pi0832 pi0956 ; n48657
g46222 nor pi1046 pi1083 ; n48658
g46223 and pi1085 n48658 ; n48659
g46224 and n48657 n48659 ; n48660
g46225 and pi0968_not n48660 ; n48661
g46226 and pi0778 n48661_not ; n48662
g46227 and pi1100 n48661 ; n48663
g46228 or n48662 n48663 ; po0935
g46229 nand pi0779 n46839_not ; po0936
g46230 nand pi0780 n46748_not ; po0937
g46231 and pi0781 n48661_not ; n48667
g46232 and pi1101 n48661 ; n48668
g46233 or n48667 n48668 ; po0938
g46234 nor n42345 n46792 ; n48670
g46235 nand n46747_not n48670 ; po0939
g46236 and pi0783 n48661_not ; n48672
g46237 and pi1109 n48661 ; n48673
g46238 or n48672 n48673 ; po0940
g46239 and pi0784 n48661_not ; n48675
g46240 and pi1110 n48661 ; n48676
g46241 or n48675 n48676 ; po0941
g46242 and pi0785 n48661_not ; n48678
g46243 and pi1102 n48661 ; n48679
g46244 or n48678 n48679 ; po0942
g46245 and pi0024 pi0954_not ; n48681
g46246 and pi0786 pi0954 ; n48682
g46247 nor n48681 n48682 ; po0943
g46248 and pi0787 n48661_not ; n48684
g46249 and pi1104 n48661 ; n48685
g46250 or n48684 n48685 ; po0944
g46251 and pi0788 n48661_not ; n48687
g46252 and pi1105 n48661 ; n48688
g46253 or n48687 n48688 ; po0945
g46254 and pi0789 n48661_not ; n48690
g46255 and pi1106 n48661 ; n48691
g46256 or n48690 n48691 ; po0946
g46257 and pi0790 n48661_not ; n48693
g46258 and pi1107 n48661 ; n48694
g46259 or n48693 n48694 ; po0947
g46260 and pi0791 n48661_not ; n48696
g46261 and pi1108 n48661 ; n48697
g46262 or n48696 n48697 ; po0948
g46263 and pi0792 n48661_not ; n48699
g46264 and pi1103 n48661 ; n48700
g46265 or n48699 n48700 ; po0949
g46266 and pi0968 n48660 ; n48702
g46267 and pi0794 n48702_not ; n48703
g46268 and pi1130 n48702 ; n48704
g46269 or n48703 n48704 ; po0951
g46270 and pi0795 n48702_not ; n48706
g46271 and pi1128 n48702 ; n48707
g46272 or n48706 n48707 ; po0952
g46273 and pi0266 pi0269_not ; n48709
g46274 and pi0278 pi0279 ; n48710
g46275 and pi0280_not n48710 ; n48711
g46276 and n48709 n48711 ; n48712
g46277 and pi0281_not n48712 ; n48713
g46278 and n47031 n48713 ; n48714
g46279 and pi0264 n48714_not ; n48715
g46280 and pi0264_not n48714 ; n48716
g46281 nor n48715 n48716 ; po0953
g46282 and pi0798 n48702_not ; n48718
g46283 and pi1124 n48702 ; n48719
g46284 or n48718 n48719 ; po0955
g46285 and pi0799 n48702_not ; n48721
g46286 and pi1107_not n48702 ; n48722
g46287 nor n48721 n48722 ; po0956
g46288 and pi0800 n48702_not ; n48724
g46289 and pi1125 n48702 ; n48725
g46290 or n48724 n48725 ; po0957
g46291 and pi0801 n48702_not ; n48727
g46292 and pi1126 n48702 ; n48728
g46293 or n48727 n48728 ; po0958
g46294 and pi0803 n48702_not ; n48730
g46295 and pi1106_not n48702 ; n48731
g46296 nor n48730 n48731 ; po0960
g46297 and pi0804 n48702_not ; n48733
g46298 and pi1109 n48702 ; n48734
g46299 or n48733 n48734 ; po0961
g46300 and pi0282_not n47029 ; n48736
g46301 and pi0270_not n48736 ; n48737
g46302 and pi0270 n48736_not ; n48738
g46303 nor n48737 n48738 ; po0962
g46304 and pi0807 n48702_not ; n48740
g46305 and pi1127 n48702 ; n48741
g46306 or n48740 n48741 ; po0964
g46307 and pi0808 n48702_not ; n48743
g46308 and pi1101 n48702 ; n48744
g46309 or n48743 n48744 ; po0965
g46310 and pi0809 n48702_not ; n48746
g46311 and pi1103_not n48702 ; n48747
g46312 nor n48746 n48747 ; po0966
g46313 and pi0810 n48702_not ; n48749
g46314 and pi1108 n48702 ; n48750
g46315 or n48749 n48750 ; po0967
g46316 and pi0811 n48702_not ; n48752
g46317 and pi1102 n48702 ; n48753
g46318 or n48752 n48753 ; po0968
g46319 and pi0812 n48702_not ; n48755
g46320 and pi1104_not n48702 ; n48756
g46321 nor n48755 n48756 ; po0969
g46322 and pi0813 n48702_not ; n48758
g46323 and pi1131 n48702 ; n48759
g46324 or n48758 n48759 ; po0970
g46325 and pi0814 n48702_not ; n48761
g46326 and pi1105_not n48702 ; n48762
g46327 nor n48761 n48762 ; po0971
g46328 and pi0815 n48702_not ; n48764
g46329 and pi1110 n48702 ; n48765
g46330 or n48764 n48765 ; po0972
g46331 and pi0816 n48702_not ; n48767
g46332 and pi1129 n48702 ; n48768
g46333 or n48767 n48768 ; po0973
g46334 and pi0269 n47027_not ; n48770
g46335 nor n47028 n48770 ; po0974
g46336 and n7643 n14172 ; n48772
g46337 or n14025 n48772 ; po0975
g46338 and pi0265 n47033_not ; n48774
g46339 nor n47034 n48774 ; po0976
g46340 and pi0277 n48737_not ; n48776
g46341 nor n47032 n48776 ; po0977
g46342 nor pi0811 pi0893 ; po0979
g46343 nor pi0982 n10074 ; n48779
g46344 and n7626 n7643 ; n48780
g46345 nor n48779 n48780 ; n48781
g46346 and n2932 n48781_not ; po0981
g46347 and pi0123 n2604 ; n48783
g46348 and pi1131 n48783_not ; n48784
g46349 and pi1127 n48783_not ; n48785
g46350 nor n48784 n48785 ; n48786
g46351 and pi0825_not n48783 ; n48787
g46352 and n48786 n48787_not ; n48788
g46353 and pi1131 n48785 ; n48789
g46354 nor n48788 n48789 ; n48790
g46355 and pi1124 pi1130_not ; n48791
g46356 and pi1124_not pi1130 ; n48792
g46357 nor n48791 n48792 ; n48793
g46358 nor pi1128 pi1129 ; n48794
g46359 and pi1128 pi1129 ; n48795
g46360 nor n48794 n48795 ; n48796
g46361 nor pi1125 pi1126 ; n48797
g46362 and pi1125 pi1126 ; n48798
g46363 nor n48797 n48798 ; n48799
g46364 and n48796 n48799_not ; n48800
g46365 and n48796_not n48799 ; n48801
g46366 nor n48800 n48801 ; n48802
g46367 and n48793 n48802 ; n48803
g46368 nor n48793 n48802 ; n48804
g46369 nor n48803 n48804 ; n48805
g46370 nor n48790 n48805 ; n48806
g46371 and pi0825 n48783 ; n48807
g46372 and n48786 n48807_not ; n48808
g46373 and n48789_not n48805 ; n48809
g46374 and n48808_not n48809 ; n48810
g46375 nor n48806 n48810 ; po0982
g46376 and pi1123 n48783_not ; n48812
g46377 and pi1122 n48783_not ; n48813
g46378 nor n48812 n48813 ; n48814
g46379 and pi0826_not n48783 ; n48815
g46380 and n48814 n48815_not ; n48816
g46381 and pi1123 n48813 ; n48817
g46382 nor n48816 n48817 ; n48818
g46383 and pi1118 pi1119_not ; n48819
g46384 and pi1118_not pi1119 ; n48820
g46385 nor n48819 n48820 ; n48821
g46386 nor pi1120 pi1121 ; n48822
g46387 and pi1120 pi1121 ; n48823
g46388 nor n48822 n48823 ; n48824
g46389 nor pi1116 pi1117 ; n48825
g46390 and pi1116 pi1117 ; n48826
g46391 nor n48825 n48826 ; n48827
g46392 and n48824 n48827_not ; n48828
g46393 and n48824_not n48827 ; n48829
g46394 nor n48828 n48829 ; n48830
g46395 and n48821 n48830 ; n48831
g46396 nor n48821 n48830 ; n48832
g46397 nor n48831 n48832 ; n48833
g46398 nor n48818 n48833 ; n48834
g46399 and pi0826 n48783 ; n48835
g46400 and n48814 n48835_not ; n48836
g46401 and n48817_not n48833 ; n48837
g46402 and n48836_not n48837 ; n48838
g46403 nor n48834 n48838 ; po0983
g46404 and pi1100 n48783_not ; n48840
g46405 and pi1107 n48783_not ; n48841
g46406 nor n48840 n48841 ; n48842
g46407 and pi0827_not n48783 ; n48843
g46408 and n48842 n48843_not ; n48844
g46409 and pi1100 n48841 ; n48845
g46410 nor n48844 n48845 ; n48846
g46411 and pi1103 pi1105_not ; n48847
g46412 and pi1103_not pi1105 ; n48848
g46413 nor n48847 n48848 ; n48849
g46414 nor pi1101 pi1102 ; n48850
g46415 and pi1101 pi1102 ; n48851
g46416 nor n48850 n48851 ; n48852
g46417 nor pi1104 pi1106 ; n48853
g46418 and pi1104 pi1106 ; n48854
g46419 nor n48853 n48854 ; n48855
g46420 and n48852 n48855_not ; n48856
g46421 and n48852_not n48855 ; n48857
g46422 nor n48856 n48857 ; n48858
g46423 and n48849 n48858 ; n48859
g46424 nor n48849 n48858 ; n48860
g46425 nor n48859 n48860 ; n48861
g46426 nor n48846 n48861 ; n48862
g46427 and pi0827 n48783 ; n48863
g46428 and n48842 n48863_not ; n48864
g46429 and n48845_not n48861 ; n48865
g46430 and n48864_not n48865 ; n48866
g46431 nor n48862 n48866 ; po0984
g46432 and pi1115 n48783_not ; n48868
g46433 and pi1114 n48783_not ; n48869
g46434 nor n48868 n48869 ; n48870
g46435 and pi0828_not n48783 ; n48871
g46436 and n48870 n48871_not ; n48872
g46437 and pi1115 n48869 ; n48873
g46438 nor n48872 n48873 ; n48874
g46439 and pi1110 pi1111_not ; n48875
g46440 and pi1110_not pi1111 ; n48876
g46441 nor n48875 n48876 ; n48877
g46442 nor pi1112 pi1113 ; n48878
g46443 and pi1112 pi1113 ; n48879
g46444 nor n48878 n48879 ; n48880
g46445 nor pi1108 pi1109 ; n48881
g46446 and pi1108 pi1109 ; n48882
g46447 nor n48881 n48882 ; n48883
g46448 and n48880 n48883_not ; n48884
g46449 and n48880_not n48883 ; n48885
g46450 nor n48884 n48885 ; n48886
g46451 and n48877 n48886 ; n48887
g46452 nor n48877 n48886 ; n48888
g46453 nor n48887 n48888 ; n48889
g46454 nor n48874 n48889 ; n48890
g46455 and pi0828 n48783 ; n48891
g46456 and n48870 n48891_not ; n48892
g46457 and n48873_not n48889 ; n48893
g46458 and n48892_not n48893 ; n48894
g46459 nor n48890 n48894 ; po0985
g46460 and n2930 n7643 ; n48896
g46461 and pi0951 n48896_not ; n48897
g46462 and pi1092 n48897_not ; po0986
g46463 and pi0281 n48712_not ; n48899
g46464 nor n48713 n48899 ; po0987
g46465 and pi0832_not pi1091 ; n48901
g46466 and pi1162 n48901 ; n48902
g46467 and n8874 n48902 ; po0989
g46468 and pi0833 n2926_not ; n48904
g46469 or n16887 n48904 ; po0990
g46470 and pi0946 n2926 ; po0991
g46471 and pi0282 n47029_not ; n48907
g46472 nor n48736 n48907 ; po0992
g46473 and pi0955_not pi1049 ; n48909
g46474 and pi0837 pi0955 ; n48910
g46475 or n48909 n48910 ; po0993
g46476 and pi0955_not pi1047 ; n48912
g46477 and pi0838 pi0955 ; n48913
g46478 or n48912 n48913 ; po0994
g46479 and pi0955_not pi1074 ; n48915
g46480 and pi0839 pi0955 ; n48916
g46481 or n48915 n48916 ; po0995
g46482 and pi0840 n2926_not ; n48918
g46483 and pi1196 n2926 ; n48919
g46484 or n48918 n48919 ; po0996
g46485 and pi0033_not n8979 ; po0997
g46486 and pi0955_not pi1035 ; n48922
g46487 and pi0842 pi0955 ; n48923
g46488 or n48922 n48923 ; po0998
g46489 and pi0955_not pi1079 ; n48925
g46490 and pi0843 pi0955 ; n48926
g46491 or n48925 n48926 ; po0999
g46492 and pi0955_not pi1078 ; n48928
g46493 and pi0844 pi0955 ; n48929
g46494 or n48928 n48929 ; po1000
g46495 and pi0955_not pi1043 ; n48931
g46496 and pi0845 pi0955 ; n48932
g46497 or n48931 n48932 ; po1001
g46498 and pi0846 n42902_not ; n48934
g46499 and pi1134 n42902 ; n48935
g46500 or n48934 n48935 ; po1002
g46501 and pi0955_not pi1055 ; n48937
g46502 and pi0847 pi0955 ; n48938
g46503 or n48937 n48938 ; po1003
g46504 and pi0955_not pi1039 ; n48940
g46505 and pi0848 pi0955 ; n48941
g46506 or n48940 n48941 ; po1004
g46507 and pi0849 n2926_not ; n48943
g46508 and pi1198 n2926 ; n48944
g46509 or n48943 n48944 ; po1005
g46510 and pi0955_not pi1048 ; n48946
g46511 and pi0850 pi0955 ; n48947
g46512 or n48946 n48947 ; po1006
g46513 and pi0955_not pi1045 ; n48949
g46514 and pi0851 pi0955 ; n48950
g46515 or n48949 n48950 ; po1007
g46516 and pi0955_not pi1062 ; n48952
g46517 and pi0852 pi0955 ; n48953
g46518 or n48952 n48953 ; po1008
g46519 and pi0955_not pi1080 ; n48955
g46520 and pi0853 pi0955 ; n48956
g46521 or n48955 n48956 ; po1009
g46522 and pi0955_not pi1051 ; n48958
g46523 and pi0854 pi0955 ; n48959
g46524 or n48958 n48959 ; po1010
g46525 and pi0955_not pi1065 ; n48961
g46526 and pi0855 pi0955 ; n48962
g46527 or n48961 n48962 ; po1011
g46528 and pi0955_not pi1067 ; n48964
g46529 and pi0856 pi0955 ; n48965
g46530 or n48964 n48965 ; po1012
g46531 and pi0955_not pi1058 ; n48967
g46532 and pi0857 pi0955 ; n48968
g46533 or n48967 n48968 ; po1013
g46534 and pi0955_not pi1087 ; n48970
g46535 and pi0858 pi0955 ; n48971
g46536 or n48970 n48971 ; po1014
g46537 and pi0955_not pi1070 ; n48973
g46538 and pi0859 pi0955 ; n48974
g46539 or n48973 n48974 ; po1015
g46540 and pi0955_not pi1076 ; n48976
g46541 and pi0860 pi0955 ; n48977
g46542 or n48976 n48977 ; po1016
g46543 and pi1093 pi1141 ; n48979
g46544 and pi0861 pi1093_not ; n48980
g46545 nor n48979 n48980 ; n48981
g46546 nor pi0228 n48981 ; n48982
g46547 nor pi0123 pi1141 ; n48983
g46548 and pi0123 pi0861_not ; n48984
g46549 and pi0228 n48983_not ; n48985
g46550 and n48984_not n48985 ; n48986
g46551 or n48982 n48986 ; po1017
g46552 and pi0862 n42902_not ; n48988
g46553 and pi1139 n42902 ; n48989
g46554 or n48988 n48989 ; po1018
g46555 and pi0863 n2926_not ; n48991
g46556 and pi1199 n2926 ; n48992
g46557 or n48991 n48992 ; po1019
g46558 and pi0864 n2926_not ; n48994
g46559 and pi1197 n2926 ; n48995
g46560 or n48994 n48995 ; po1020
g46561 and pi0955_not pi1040 ; n48997
g46562 and pi0865 pi0955 ; n48998
g46563 or n48997 n48998 ; po1021
g46564 and pi0955_not pi1053 ; n49000
g46565 and pi0866 pi0955 ; n49001
g46566 or n49000 n49001 ; po1022
g46567 and pi0955_not pi1057 ; n49003
g46568 and pi0867 pi0955 ; n49004
g46569 or n49003 n49004 ; po1023
g46570 and pi0955_not pi1063 ; n49006
g46571 and pi0868 pi0955 ; n49007
g46572 or n49006 n49007 ; po1024
g46573 and pi1093 pi1140 ; n49009
g46574 and pi0869 pi1093_not ; n49010
g46575 nor n49009 n49010 ; n49011
g46576 nor pi0228 n49011 ; n49012
g46577 nor pi0123 pi1140 ; n49013
g46578 and pi0123 pi0869_not ; n49014
g46579 and pi0228 n49013_not ; n49015
g46580 and n49014_not n49015 ; n49016
g46581 or n49012 n49016 ; po1025
g46582 and pi0955_not pi1069 ; n49018
g46583 and pi0870 pi0955 ; n49019
g46584 or n49018 n49019 ; po1026
g46585 and pi0955_not pi1072 ; n49021
g46586 and pi0871 pi0955 ; n49022
g46587 or n49021 n49022 ; po1027
g46588 and pi0955_not pi1084 ; n49024
g46589 and pi0872 pi0955 ; n49025
g46590 or n49024 n49025 ; po1028
g46591 and pi0955_not pi1044 ; n49027
g46592 and pi0873 pi0955 ; n49028
g46593 or n49027 n49028 ; po1029
g46594 and pi0955_not pi1036 ; n49030
g46595 and pi0874 pi0955 ; n49031
g46596 or n49030 n49031 ; po1030
g46597 and pi1093 pi1136_not ; n49033
g46598 nor pi0875 pi1093 ; n49034
g46599 nor n49033 n49034 ; n49035
g46600 nor pi0228 n49035 ; n49036
g46601 and pi0123_not pi1136 ; n49037
g46602 and pi0123 pi0875 ; n49038
g46603 and pi0228 n49037_not ; n49039
g46604 and n49038_not n49039 ; n49040
g46605 nor n49036 n49040 ; po1031
g46606 and pi0955_not pi1037 ; n49042
g46607 and pi0876 pi0955 ; n49043
g46608 or n49042 n49043 ; po1032
g46609 and pi1093 pi1138 ; n49045
g46610 and pi0877 pi1093_not ; n49046
g46611 nor n49045 n49046 ; n49047
g46612 nor pi0228 n49047 ; n49048
g46613 nor pi0123 pi1138 ; n49049
g46614 and pi0123 pi0877_not ; n49050
g46615 and pi0228 n49049_not ; n49051
g46616 and n49050_not n49051 ; n49052
g46617 or n49048 n49052 ; po1033
g46618 and pi1093 pi1137 ; n49054
g46619 and pi0878 pi1093_not ; n49055
g46620 nor n49054 n49055 ; n49056
g46621 nor pi0228 n49056 ; n49057
g46622 nor pi0123 pi1137 ; n49058
g46623 and pi0123 pi0878_not ; n49059
g46624 and pi0228 n49058_not ; n49060
g46625 and n49059_not n49060 ; n49061
g46626 or n49057 n49061 ; po1034
g46627 and pi1093 pi1135 ; n49063
g46628 and pi0879 pi1093_not ; n49064
g46629 nor n49063 n49064 ; n49065
g46630 nor pi0228 n49065 ; n49066
g46631 nor pi0123 pi1135 ; n49067
g46632 and pi0123 pi0879_not ; n49068
g46633 and pi0228 n49067_not ; n49069
g46634 and n49068_not n49069 ; n49070
g46635 or n49066 n49070 ; po1035
g46636 and pi0955_not pi1081 ; n49072
g46637 and pi0880 pi0955 ; n49073
g46638 or n49072 n49073 ; po1036
g46639 and pi0955_not pi1059 ; n49075
g46640 and pi0881 pi0955 ; n49076
g46641 or n49075 n49076 ; po1037
g46642 and pi0883_not n48783 ; n49078
g46643 or n48841 n49078 ; po1039
g46644 and pi1124 n48783_not ; n49080
g46645 and pi0884_not n48783 ; n49081
g46646 or n49080 n49081 ; po1040
g46647 and pi1125 n48783_not ; n49083
g46648 and pi0885_not n48783 ; n49084
g46649 or n49083 n49084 ; po1041
g46650 and pi1109 n48783_not ; n49086
g46651 and pi0886_not n48783 ; n49087
g46652 or n49086 n49087 ; po1042
g46653 and pi0887_not n48783 ; n49089
g46654 or n48840 n49089 ; po1043
g46655 and pi1120 n48783_not ; n49091
g46656 and pi0888_not n48783 ; n49092
g46657 or n49091 n49092 ; po1044
g46658 and pi1103 n48783_not ; n49094
g46659 and pi0889_not n48783 ; n49095
g46660 or n49094 n49095 ; po1045
g46661 and pi1126 n48783_not ; n49097
g46662 and pi0890_not n48783 ; n49098
g46663 or n49097 n49098 ; po1046
g46664 and pi1116 n48783_not ; n49100
g46665 and pi0891_not n48783 ; n49101
g46666 or n49100 n49101 ; po1047
g46667 and pi1101 n48783_not ; n49103
g46668 and pi0892_not n48783 ; n49104
g46669 or n49103 n49104 ; po1048
g46670 and pi1119 n48783_not ; n49106
g46671 and pi0894_not n48783 ; n49107
g46672 or n49106 n49107 ; po1050
g46673 and pi1113 n48783_not ; n49109
g46674 and pi0895_not n48783 ; n49110
g46675 or n49109 n49110 ; po1051
g46676 and pi1118 n48783_not ; n49112
g46677 and pi0896_not n48783 ; n49113
g46678 or n49112 n49113 ; po1052
g46679 and pi1129 n48783_not ; n49115
g46680 and pi0898_not n48783 ; n49116
g46681 or n49115 n49116 ; po1054
g46682 and pi0899_not n48783 ; n49118
g46683 or n48868 n49118 ; po1055
g46684 and pi1110 n48783_not ; n49120
g46685 and pi0900_not n48783 ; n49121
g46686 or n49120 n49121 ; po1056
g46687 and pi1111 n48783_not ; n49123
g46688 and pi0902_not n48783 ; n49124
g46689 or n49123 n49124 ; po1058
g46690 and pi1121 n48783_not ; n49126
g46691 and pi0903_not n48783 ; n49127
g46692 or n49126 n49127 ; po1059
g46693 and pi0904_not n48783 ; n49129
g46694 or n48785 n49129 ; po1060
g46695 and pi0905_not n48783 ; n49131
g46696 or n48784 n49131 ; po1061
g46697 and pi1128 n48783_not ; n49133
g46698 and pi0906_not n48783 ; n49134
g46699 or n49133 n49134 ; po1062
g46700 nor pi0782 pi0907 ; n49136
g46701 nor pi0624 pi0979 ; n49137
g46702 and pi0598_not pi0979 ; n49138
g46703 and pi0782 n49137_not ; n49139
g46704 and n49138_not n49139 ; n49140
g46705 nor pi0604 pi0979 ; n49141
g46706 and pi0615 pi0979 ; n49142
g46707 nor n49141 n49142 ; n49143
g46708 and pi0782 n49143_not ; n49144
g46709 nor n49136 n49140 ; n49145
g46710 and n49144_not n49145 ; po1063
g46711 and pi0908_not n48783 ; n49147
g46712 or n48813 n49147 ; po1064
g46713 and pi1105 n48783_not ; n49149
g46714 and pi0909_not n48783 ; n49150
g46715 or n49149 n49150 ; po1065
g46716 and pi1117 n48783_not ; n49152
g46717 and pi0910_not n48783 ; n49153
g46718 or n49152 n49153 ; po1066
g46719 and pi1130 n48783_not ; n49155
g46720 and pi0911_not n48783 ; n49156
g46721 or n49155 n49156 ; po1067
g46722 and pi0912_not n48783 ; n49158
g46723 or n48869 n49158 ; po1068
g46724 and pi1106 n48783_not ; n49160
g46725 and pi0913_not n48783 ; n49161
g46726 or n49160 n49161 ; po1069
g46727 and pi0280 n47026_not ; n49163
g46728 nor n47027 n49163 ; po1070
g46729 and pi1108 n48783_not ; n49165
g46730 and pi0915_not n48783 ; n49166
g46731 or n49165 n49166 ; po1071
g46732 and pi0916_not n48783 ; n49168
g46733 or n48812 n49168 ; po1072
g46734 and pi1112 n48783_not ; n49170
g46735 and pi0917_not n48783 ; n49171
g46736 or n49170 n49171 ; po1073
g46737 and pi1104 n48783_not ; n49173
g46738 and pi0918_not n48783 ; n49174
g46739 or n49173 n49174 ; po1074
g46740 and pi1102 n48783_not ; n49176
g46741 and pi0919_not n48783 ; n49177
g46742 or n49176 n49177 ; po1075
g46743 and pi1093 pi1139 ; n49179
g46744 and pi0920 pi1093_not ; n49180
g46745 or n49179 n49180 ; po1076
g46746 and pi0921 pi1093_not ; n49182
g46747 or n49009 n49182 ; po1077
g46748 nor pi0922 pi1093 ; n49184
g46749 and pi1093 pi1152_not ; n49185
g46750 nor n49184 n49185 ; po1078
g46751 nor pi0923 pi1093 ; n49187
g46752 and pi1093 pi1154_not ; n49188
g46753 nor n49187 n49188 ; po1079
g46754 and pi0300_not pi0301 ; n49190
g46755 and pi0311 pi0312_not ; n49191
g46756 and n49190 n49191 ; po1080
g46757 nor pi0925 pi1093 ; n49193
g46758 and pi1093 pi1155_not ; n49194
g46759 nor n49193 n49194 ; po1081
g46760 nor pi0926 pi1093 ; n49196
g46761 and pi1093 pi1157_not ; n49197
g46762 nor n49196 n49197 ; po1082
g46763 nor pi0927 pi1093 ; n49199
g46764 and pi1093 pi1145_not ; n49200
g46765 nor n49199 n49200 ; po1083
g46766 nor pi0928 pi1093 ; n49202
g46767 nor n49033 n49202 ; po1084
g46768 nor pi0929 pi1093 ; n49204
g46769 and pi1093 pi1144_not ; n49205
g46770 nor n49204 n49205 ; po1085
g46771 nor pi0930 pi1093 ; n49207
g46772 and pi1093 pi1134_not ; n49208
g46773 nor n49207 n49208 ; po1086
g46774 nor pi0931 pi1093 ; n49210
g46775 and pi1093 pi1150_not ; n49211
g46776 nor n49210 n49211 ; po1087
g46777 and pi0932 pi1093_not ; n49213
g46778 or n42891 n49213 ; po1088
g46779 and pi0933 pi1093_not ; n49215
g46780 or n49054 n49215 ; po1089
g46781 nor pi0934 pi1093 ; n49217
g46782 and pi1093 pi1147_not ; n49218
g46783 nor n49217 n49218 ; po1090
g46784 and pi0935 pi1093_not ; n49220
g46785 or n48979 n49220 ; po1091
g46786 nor pi0936 pi1093 ; n49222
g46787 and pi1093 pi1149_not ; n49223
g46788 nor n49222 n49223 ; po1092
g46789 nor pi0937 pi1093 ; n49225
g46790 and pi1093 pi1148_not ; n49226
g46791 nor n49225 n49226 ; po1093
g46792 and pi0938 pi1093_not ; n49228
g46793 or n49063 n49228 ; po1094
g46794 nor pi0939 pi1093 ; n49230
g46795 and pi1093 pi1146_not ; n49231
g46796 nor n49230 n49231 ; po1095
g46797 and pi0940 pi1093_not ; n49233
g46798 or n49045 n49233 ; po1096
g46799 nor pi0941 pi1093 ; n49235
g46800 and pi1093 pi1153_not ; n49236
g46801 nor n49235 n49236 ; po1097
g46802 nor pi0942 pi1093 ; n49238
g46803 and pi1093 pi1156_not ; n49239
g46804 nor n49238 n49239 ; po1098
g46805 nor pi0943 pi1093 ; n49241
g46806 and pi1093 pi1151_not ; n49242
g46807 nor n49241 n49242 ; po1099
g46808 and pi1093 pi1143 ; n49244
g46809 and pi0944 pi1093_not ; n49245
g46810 or n49244 n49245 ; po1100
g46811 and pi0230 n2926 ; po1102
g46812 and pi0782_not pi0947 ; n49248
g46813 or n49140 n49248 ; po1103
g46814 nor pi0266 pi0992 ; n49250
g46815 nor n47026 n49250 ; po1104
g46816 nor pi0313 pi0954 ; n49252
g46817 and pi0949 pi0954 ; n49253
g46818 or n49252 n49253 ; po1105
g46819 and n7626_not n14271 ; po1107
g46820 and pi0957 pi1092 ; n49256
g46821 or pi0031 n49256 ; po1112
g46822 and pi0782_not pi0960 ; po1115
g46823 and pi0230_not pi0961 ; po1116
g46824 and pi0782_not pi0963 ; po1118
g46825 and pi0230_not pi0967 ; po1122
g46826 and pi0230_not pi0969 ; po1124
g46827 and pi0782_not pi0970 ; po1125
g46828 and pi0230_not pi0971 ; po1126
g46829 and pi0782_not pi0972 ; po1127
g46830 and pi0230_not pi0974 ; po1128
g46831 and pi0782_not pi0975 ; po1129
g46832 and pi0230_not pi0977 ; po1131
g46833 and pi0782_not pi0978 ; po1132
g46834 nand pi0598_not pi0615 ; po1133
g46835 and pi0824 pi1092 ; po1135
g46836 or pi0604 pi0624 ; po1137
g46974 not n3001 ; n3001_not
g46975 not n4000 ; n4000_not
g46976 not n3110 ; n3110_not
g46977 not n4010 ; n4010_not
g46978 not n5100 ; n5100_not
g46979 not n4110 ; n4110_not
g46980 not n3021 ; n3021_not
g46981 not n4101 ; n4101_not
g46982 not n3300 ; n3300_not
g46983 not n6000 ; n6000_not
g46984 not n3012 ; n3012_not
g46985 not n3120 ; n3120_not
g46986 not n3111 ; n3111_not
g46987 not n5010 ; n5010_not
g46988 not n4200 ; n4200_not
g46989 not n3103 ; n3103_not
g46990 not n6010 ; n6010_not
g46991 not n4012 ; n4012_not
g46992 not n3004 ; n3004_not
g46993 not n6100 ; n6100_not
g46994 not n4102 ; n4102_not
g46995 not n3220 ; n3220_not
g46996 not n3130 ; n3130_not
g46997 not n3202 ; n3202_not
g46998 not n3040 ; n3040_not
g46999 not n3022 ; n3022_not
g47000 not n5011 ; n5011_not
g47001 not n5201 ; n5201_not
g47002 not n4031 ; n4031_not
g47003 not n4301 ; n4301_not
g47004 not n4130 ; n4130_not
g47005 not n5102 ; n5102_not
g47006 not n7001 ; n7001_not
g47007 not n3122 ; n3122_not
g47008 not n4202 ; n4202_not
g47009 not n3302 ; n3302_not
g47010 not n5003 ; n5003_not
g47011 not n3041 ; n3041_not
g47012 not n3023 ; n3023_not
g47013 not n4112 ; n4112_not
g47014 not n5012 ; n5012_not
g47015 not n5210 ; n5210_not
g47016 not n4040 ; n4040_not
g47017 not n4310 ; n4310_not
g47018 not n3014 ; n3014_not
g47019 not n3104 ; n3104_not
g47020 not n3410 ; n3410_not
g47021 not n5021 ; n5021_not
g47022 not n6110 ; n6110_not
g47023 not n4022 ; n4022_not
g47024 not n7020 ; n7020_not
g47025 not n4140 ; n4140_not
g47026 not n7011 ; n7011_not
g47027 not n5211 ; n5211_not
g47028 not n3411 ; n3411_not
g47029 not n3213 ; n3213_not
g47030 not n5103 ; n5103_not
g47031 not n3222 ; n3222_not
g47032 not n3501 ; n3501_not
g47033 not n2610 ; n2610_not
g47034 not n2502 ; n2502_not
g47035 not n6012 ; n6012_not
g47036 not n6030 ; n6030_not
g47037 not n7101 ; n7101_not
g47038 not n3312 ; n3312_not
g47039 not n9000 ; n9000_not
g47040 not n8001 ; n8001_not
g47041 not n3600 ; n3600_not
g47042 not n4311 ; n4311_not
g47043 not n4203 ; n4203_not
g47044 not n2511 ; n2511_not
g47045 not n5031 ; n5031_not
g47046 not n4050 ; n4050_not
g47047 not n5022 ; n5022_not
g47048 not n3006 ; n3006_not
g47049 not n4041 ; n4041_not
g47050 not n3114 ; n3114_not
g47051 not n6102 ; n6102_not
g47052 not n3123 ; n3123_not
g47053 not n3402 ; n3402_not
g47054 not n4500 ; n4500_not
g47055 not n4032 ; n4032_not
g47056 not n3033 ; n3033_not
g47057 not n3141 ; n3141_not
g47058 not n3042 ; n3042_not
g47059 not n3150 ; n3150_not
g47060 not n4113 ; n4113_not
g47061 not n3051 ; n3051_not
g47062 not n2530 ; n2530_not
g47063 not n3052 ; n3052_not
g47064 not n4321 ; n4321_not
g47065 not n5410 ; n5410_not
g47066 not n2521 ; n2521_not
g47067 not n3403 ; n3403_not
g47068 not n3331 ; n3331_not
g47069 not n4312 ; n4312_not
g47070 not n2710 ; n2710_not
g47071 not n5230 ; n5230_not
g47072 not n3421 ; n3421_not
g47073 not n2800 ; n2800_not
g47074 not n3061 ; n3061_not
g47075 not n3043 ; n3043_not
g47076 not n3511 ; n3511_not
g47077 not n5221 ; n5221_not
g47078 not n4600 ; n4600_not
g47079 not n9010 ; n9010_not
g47080 not n3232 ; n3232_not
g47081 not n3241 ; n3241_not
g47082 not n3250 ; n3250_not
g47083 not n3142 ; n3142_not
g47084 not n3133 ; n3133_not
g47085 not n4501 ; n4501_not
g47086 not n3124 ; n3124_not
g47087 not n8011 ; n8011_not
g47088 not n3313 ; n3313_not
g47089 not n3340 ; n3340_not
g47090 not n2611 ; n2611_not
g47091 not n4330 ; n4330_not
g47092 not n2503 ; n2503_not
g47093 not n3016 ; n3016_not
g47094 not n2620 ; n2620_not
g47095 not n5104 ; n5104_not
g47096 not n6040 ; n6040_not
g47097 not n5032 ; n5032_not
g47098 not n5131 ; n5131_not
g47099 not n4114 ; n4114_not
g47100 not n4123 ; n4123_not
g47101 not n5014 ; n5014_not
g47102 not n5050 ; n5050_not
g47103 not n7003 ; n7003_not
g47104 not n4006 ; n4006_not
g47105 not n4231 ; n4231_not
g47106 not n3412 ; n3412_not
g47107 not n3502 ; n3502_not
g47108 not n6220 ; n6220_not
g47109 not n5212 ; n5212_not
g47110 not n4042 ; n4042_not
g47111 not n6022 ; n6022_not
g47112 not n3610 ; n3610_not
g47113 not n6112 ; n6112_not
g47114 not n7201 ; n7201_not
g47115 not n4204 ; n4204_not
g47116 not n6400 ; n6400_not
g47117 not n7120 ; n7120_not
g47118 not n4520 ; n4520_not
g47119 not n6230 ; n6230_not
g47120 not n3053 ; n3053_not
g47121 not n3062 ; n3062_not
g47122 not n3080 ; n3080_not
g47123 not n6320 ; n6320_not
g47124 not n6104 ; n6104_not
g47125 not n3305 ; n3305_not
g47126 not n7103 ; n7103_not
g47127 not n8012 ; n8012_not
g47128 not n8003 ; n8003_not
g47129 not n3341 ; n3341_not
g47130 not n7130 ; n7130_not
g47131 not n4331 ; n4331_not
g47132 not n4313 ; n4313_not
g47133 not n4322 ; n4322_not
g47134 not n4214 ; n4214_not
g47135 not n7301 ; n7301_not
g47136 not n7310 ; n7310_not
g47137 not n4232 ; n4232_not
g47138 not n3521 ; n3521_not
g47139 not n4250 ; n4250_not
g47140 not n3512 ; n3512_not
g47141 not n2441 ; n2441_not
g47142 not n3440 ; n3440_not
g47143 not n4223 ; n4223_not
g47144 not n3143 ; n3143_not
g47145 not n4124 ; n4124_not
g47146 not n4133 ; n4133_not
g47147 not n3161 ; n3161_not
g47148 not n3170 ; n3170_not
g47149 not n4412 ; n4412_not
g47150 not n4430 ; n4430_not
g47151 not n4142 ; n4142_not
g47152 not n3701 ; n3701_not
g47153 not n3224 ; n3224_not
g47154 not n6050 ; n6050_not
g47155 not n7013 ; n7013_not
g47156 not n8201 ; n8201_not
g47157 not n7022 ; n7022_not
g47158 not n3260 ; n3260_not
g47159 not n8120 ; n8120_not
g47160 not n4403 ; n4403_not
g47161 not n8111 ; n8111_not
g47162 not n4304 ; n4304_not
g47163 not n6032 ; n6032_not
g47164 not n3602 ; n3602_not
g47165 not n5213 ; n5213_not
g47166 not n5033 ; n5033_not
g47167 not n2900 ; n2900_not
g47168 not n5222 ; n5222_not
g47169 not n3017 ; n3017_not
g47170 not n2603 ; n2603_not
g47171 not n2801 ; n2801_not
g47172 not n5312 ; n5312_not
g47173 not n5060 ; n5060_not
g47174 not n2630 ; n2630_not
g47175 not n5123 ; n5123_not
g47176 not n5420 ; n5420_not
g47177 not n5402 ; n5402_not
g47178 not n9002 ; n9002_not
g47179 not n9011 ; n9011_not
g47180 not n5114 ; n5114_not
g47181 not n5150 ; n5150_not
g47182 not n9101 ; n9101_not
g47183 not n2711 ; n2711_not
g47184 not n5132 ; n5132_not
g47185 not n5231 ; n5231_not
g47186 not n5204 ; n5204_not
g47187 not n4700 ; n4700_not
g47188 not n2810 ; n2810_not
g47189 not n2513 ; n2513_not
g47190 not n2504 ; n2504_not
g47191 not n3026 ; n3026_not
g47192 not n9200 ; n9200_not
g47193 not n3035 ; n3035_not
g47194 not n5330 ; n5330_not
g47195 not n9210 ; n9210_not
g47196 not n5160 ; n5160_not
g47197 not n7320 ; n7320_not
g47198 not n2532 ; n2532_not
g47199 not n3531 ; n3531_not
g47200 not n3306 ; n3306_not
g47201 not n4233 ; n4233_not
g47202 not n7221 ; n7221_not
g47203 not n7212 ; n7212_not
g47204 not n5142 ; n5142_not
g47205 not n7203 ; n7203_not
g47206 not n2640 ; n2640_not
g47207 not n6006 ; n6006_not
g47208 not n5133 ; n5133_not
g47209 not n7113 ; n7113_not
g47210 not n3432 ; n3432_not
g47211 not n3342 ; n3342_not
g47212 not n4314 ; n4314_not
g47213 not n3450 ; n3450_not
g47214 not n2802 ; n2802_not
g47215 not n5214 ; n5214_not
g47216 not n7500 ; n7500_not
g47217 not n4260 ; n4260_not
g47218 not n2442 ; n2442_not
g47219 not n3504 ; n3504_not
g47220 not n4242 ; n4242_not
g47221 not n9300 ; n9300_not
g47222 not n6411 ; n6411_not
g47223 not n3801 ; n3801_not
g47224 not n6600 ; n6600_not
g47225 not n5043 ; n5043_not
g47226 not n4071 ; n4071_not
g47227 not n4053 ; n4053_not
g47228 not n4062 ; n4062_not
g47229 not n2523 ; n2523_not
g47230 not n6060 ; n6060_not
g47231 not n4044 ; n4044_not
g47232 not n6114 ; n6114_not
g47233 not n6123 ; n6123_not
g47234 not n6402 ; n6402_not
g47235 not n5007 ; n5007_not
g47236 not n3900 ; n3900_not
g47237 not n4008 ; n4008_not
g47238 not n6330 ; n6330_not
g47239 not n6141 ; n6141_not
g47240 not n6150 ; n6150_not
g47241 not n6213 ; n6213_not
g47242 not n2721 ; n2721_not
g47243 not n6024 ; n6024_not
g47244 not n3621 ; n3621_not
g47245 not n7041 ; n7041_not
g47246 not n4161 ; n4161_not
g47247 not n6042 ; n6042_not
g47248 not n7032 ; n7032_not
g47249 not n4116 ; n4116_not
g47250 not n9030 ; n9030_not
g47251 not n7005 ; n7005_not
g47252 not n2631 ; n2631_not
g47253 not n4134 ; n4134_not
g47254 not n6510 ; n6510_not
g47255 not n5052 ; n5052_not
g47256 not n8202 ; n8202_not
g47257 not n5610 ; n5610_not
g47258 not n3126 ; n3126_not
g47259 not n3054 ; n3054_not
g47260 not n3117 ; n3117_not
g47261 not n3081 ; n3081_not
g47262 not n3234 ; n3234_not
g47263 not n3261 ; n3261_not
g47264 not n4422 ; n4422_not
g47265 not n3216 ; n3216_not
g47266 not n5340 ; n5340_not
g47267 not n8400 ; n8400_not
g47268 not n8040 ; n8040_not
g47269 not n3243 ; n3243_not
g47270 not n5430 ; n5430_not
g47271 not n3252 ; n3252_not
g47272 not n3045 ; n3045_not
g47273 not n4620 ; n4620_not
g47274 not n8211 ; n8211_not
g47275 not n3063 ; n3063_not
g47276 not n4413 ; n4413_not
g47277 not n5403 ; n5403_not
g47278 not n8301 ; n8301_not
g47279 not n2703 ; n2703_not
g47280 not n4512 ; n4512_not
g47281 not n4404 ; n4404_not
g47282 not n5520 ; n5520_not
g47283 not n2505 ; n2505_not
g47284 not n3072 ; n3072_not
g47285 not n4440 ; n4440_not
g47286 not n3144 ; n3144_not
g47287 not n3270 ; n3270_not
g47288 not n4431 ; n4431_not
g47289 not n4602 ; n4602_not
g47290 not n8311 ; n8311_not
g47291 not n6205 ; n6205_not
g47292 not n5107 ; n5107_not
g47293 not n4153 ; n4153_not
g47294 not n9031 ; n9031_not
g47295 not n2533 ; n2533_not
g47296 not n7141 ; n7141_not
g47297 not n9022 ; n9022_not
g47298 not n5008 ; n5008_not
g47299 not n7024 ; n7024_not
g47300 not n6052 ; n6052_not
g47301 not n7420 ; n7420_not
g47302 not n3154 ; n3154_not
g47303 not n4180 ; n4180_not
g47304 not n7105 ; n7105_not
g47305 not n3640 ; n3640_not
g47306 not n3613 ; n3613_not
g47307 not n3172 ; n3172_not
g47308 not n3163 ; n3163_not
g47309 not n3028 ; n3028_not
g47310 not n5116 ; n5116_not
g47311 not n2722 ; n2722_not
g47312 not n7051 ; n7051_not
g47313 not n9121 ; n9121_not
g47314 not n7033 ; n7033_not
g47315 not n6061 ; n6061_not
g47316 not n6700 ; n6700_not
g47317 not n3118 ; n3118_not
g47318 not n6502 ; n6502_not
g47319 not n6511 ; n6511_not
g47320 not n5512 ; n5512_not
g47321 not n4081 ; n4081_not
g47322 not n2524 ; n2524_not
g47323 not n5044 ; n5044_not
g47324 not n3019 ; n3019_not
g47325 not n8401 ; n8401_not
g47326 not n3811 ; n3811_not
g47327 not n5035 ; n5035_not
g47328 not n6322 ; n6322_not
g47329 not n2803 ; n2803_not
g47330 not n2551 ; n2551_not
g47331 not n6106 ; n6106_not
g47332 not n4063 ; n4063_not
g47333 not n3820 ; n3820_not
g47334 not n3145 ; n3145_not
g47335 not n4810 ; n4810_not
g47336 not n3136 ; n3136_not
g47337 not n3703 ; n3703_not
g47338 not n5350 ; n5350_not
g47339 not n2641 ; n2641_not
g47340 not n4135 ; n4135_not
g47341 not n3127 ; n3127_not
g47342 not n2632 ; n2632_not
g47343 not n2560 ; n2560_not
g47344 not n8041 ; n8041_not
g47345 not n5080 ; n5080_not
g47346 not n4522 ; n4522_not
g47347 not n2605 ; n2605_not
g47348 not n5062 ; n5062_not
g47349 not n5026 ; n5026_not
g47350 not n9310 ; n9310_not
g47351 not n9130 ; n9130_not
g47352 not n2506 ; n2506_not
g47353 not n3361 ; n3361_not
g47354 not n3910 ; n3910_not
g47355 not n3406 ; n3406_not
g47356 not n5233 ; n5233_not
g47357 not n4711 ; n4711_not
g47358 not n3424 ; n3424_not
g47359 not n6304 ; n6304_not
g47360 not n4306 ; n4306_not
g47361 not n2740 ; n2740_not
g47362 not n2911 ; n2911_not
g47363 not n2902 ; n2902_not
g47364 not n3442 ; n3442_not
g47365 not n6232 ; n6232_not
g47366 not n3451 ; n3451_not
g47367 not n7510 ; n7510_not
g47368 not n8320 ; n8320_not
g47369 not n8032 ; n8032_not
g47370 not n4900 ; n4900_not
g47371 not n6214 ; n6214_not
g47372 not n8005 ; n8005_not
g47373 not n6250 ; n6250_not
g47374 not n3343 ; n3343_not
g47375 not n9301 ; n9301_not
g47376 not n5251 ; n5251_not
g47377 not n8122 ; n8122_not
g47378 not n2452 ; n2452_not
g47379 not n4351 ; n4351_not
g47380 not n5701 ; n5701_not
g47381 not n3325 ; n3325_not
g47382 not n3055 ; n3055_not
g47383 not n4333 ; n4333_not
g47384 not n8131 ; n8131_not
g47385 not n4702 ; n4702_not
g47386 not n3208 ; n3208_not
g47387 not n5314 ; n5314_not
g47388 not n8221 ; n8221_not
g47389 not n5530 ; n5530_not
g47390 not n7321 ; n7321_not
g47391 not n3550 ; n3550_not
g47392 not n4630 ; n4630_not
g47393 not n4216 ; n4216_not
g47394 not n2515 ; n2515_not
g47395 not n7231 ; n7231_not
g47396 not n4207 ; n4207_not
g47397 not n5071 ; n5071_not
g47398 not n6403 ; n6403_not
g47399 not n8302 ; n8302_not
g47400 not n3181 ; n3181_not
g47401 not n5611 ; n5611_not
g47402 not n3460 ; n3460_not
g47403 not n4540 ; n4540_not
g47404 not n4270 ; n4270_not
g47405 not n4261 ; n4261_not
g47406 not n7411 ; n7411_not
g47407 not n5206 ; n5206_not
g47408 not n3280 ; n3280_not
g47409 not n7402 ; n7402_not
g47410 not n4009 ; n4009_not
g47411 not n4423 ; n4423_not
g47412 not n3217 ; n3217_not
g47413 not n3505 ; n3505_not
g47414 not n5170 ; n5170_not
g47415 not n3514 ; n3514_not
g47416 not n4171 ; n4171_not
g47417 not n5161 ; n5161_not
g47418 not n2920 ; n2920_not
g47419 not n9103 ; n9103_not
g47420 not n3416 ; n3416_not
g47421 not n6224 ; n6224_not
g47422 not n4910 ; n4910_not
g47423 not n6152 ; n6152_not
g47424 not n4541 ; n4541_not
g47425 not n6125 ; n6125_not
g47426 not n4037 ; n4037_not
g47427 not n5441 ; n5441_not
g47428 not n4019 ; n4019_not
g47429 not n6116 ; n6116_not
g47430 not n5450 ; n5450_not
g47431 not n5162 ; n5162_not
g47432 not n4604 ; n4604_not
g47433 not n5135 ; n5135_not
g47434 not n4262 ; n4262_not
g47435 not n5072 ; n5072_not
g47436 not n6242 ; n6242_not
g47437 not n5351 ; n5351_not
g47438 not n4415 ; n4415_not
g47439 not n4235 ; n4235_not
g47440 not n4622 ; n4622_not
g47441 not n4172 ; n4172_not
g47442 not n4712 ; n4712_not
g47443 not n5234 ; n5234_not
g47444 not n4703 ; n4703_not
g47445 not n4334 ; n4334_not
g47446 not n4406 ; n4406_not
g47447 not n5261 ; n5261_not
g47448 not n4361 ; n4361_not
g47449 not n5720 ; n5720_not
g47450 not n5711 ; n5711_not
g47451 not n5702 ; n5702_not
g47452 not n5216 ; n5216_not
g47453 not n5306 ; n5306_not
g47454 not n4316 ; n4316_not
g47455 not n5333 ; n5333_not
g47456 not n4514 ; n4514_not
g47457 not n4073 ; n4073_not
g47458 not n6080 ; n6080_not
g47459 not n5522 ; n5522_not
g47460 not n6053 ; n6053_not
g47461 not n6062 ; n6062_not
g47462 not n4505 ; n4505_not
g47463 not n5054 ; n5054_not
g47464 not n5432 ; n5432_not
g47465 not n5081 ; n5081_not
g47466 not n5090 ; n5090_not
g47467 not n5405 ; n5405_not
g47468 not n4802 ; n4802_not
g47469 not n5108 ; n5108_not
g47470 not n6044 ; n6044_not
g47471 not n4163 ; n4163_not
g47472 not n5117 ; n5117_not
g47473 not n4181 ; n4181_not
g47474 not n5360 ; n5360_not
g47475 not n6017 ; n6017_not
g47476 not n4190 ; n4190_not
g47477 not n4208 ; n4208_not
g47478 not n4217 ; n4217_not
g47479 not n6008 ; n6008_not
g47480 not n3119 ; n3119_not
g47481 not n6170 ; n6170_not
g47482 not n9401 ; n9401_not
g47483 not n2732 ; n2732_not
g47484 not n7007 ; n7007_not
g47485 not n3407 ; n3407_not
g47486 not n6215 ; n6215_not
g47487 not n9311 ; n9311_not
g47488 not n8501 ; n8501_not
g47489 not n7034 ; n7034_not
g47490 not n3434 ; n3434_not
g47491 not n7052 ; n7052_not
g47492 not n7061 ; n7061_not
g47493 not n9212 ; n9212_not
g47494 not n2930 ; n2930_not
g47495 not n3146 ; n3146_not
g47496 not n6260 ; n6260_not
g47497 not n3137 ; n3137_not
g47498 not n2813 ; n2813_not
g47499 not n7601 ; n7601_not
g47500 not n3128 ; n3128_not
g47501 not n9122 ; n9122_not
g47502 not n7250 ; n7250_not
g47503 not n7304 ; n7304_not
g47504 not n7430 ; n7430_not
g47505 not n3533 ; n3533_not
g47506 not n9032 ; n9032_not
g47507 not n7340 ; n7340_not
g47508 not n9023 ; n9023_not
g47509 not n9014 ; n9014_not
g47510 not n2741 ; n2741_not
g47511 not n9230 ; n9230_not
g47512 not n3650 ; n3650_not
g47513 not n8510 ; n8510_not
g47514 not n3074 ; n3074_not
g47515 not n3632 ; n3632_not
g47516 not n3623 ; n3623_not
g47517 not n7511 ; n7511_not
g47518 not n7115 ; n7115_not
g47519 not n9203 ; n9203_not
g47520 not n3047 ; n3047_not
g47521 not n7205 ; n7205_not
g47522 not n7214 ; n7214_not
g47523 not n9104 ; n9104_not
g47524 not n3038 ; n3038_not
g47525 not n6440 ; n6440_not
g47526 not n8321 ; n8321_not
g47527 not n3353 ; n3353_not
g47528 not n6431 ; n6431_not
g47529 not n3173 ; n3173_not
g47530 not n6404 ; n6404_not
g47531 not n6413 ; n6413_not
g47532 not n2525 ; n2525_not
g47533 not n2444 ; n2444_not
g47534 not n3191 ; n3191_not
g47535 not n3218 ; n3218_not
g47536 not n8015 ; n8015_not
g47537 not n2543 ; n2543_not
g47538 not n2903 ; n2903_not
g47539 not n3209 ; n3209_not
g47540 not n6341 ; n6341_not
g47541 not n3155 ; n3155_not
g47542 not n6305 ; n6305_not
g47543 not n6512 ; n6512_not
g47544 not n8042 ; n8042_not
g47545 not n5460 ; n5460_not
g47546 not n3039 ; n3039_not
g47547 not n3273 ; n3273_not
g47548 not n2625 ; n2625_not
g47549 not n7620 ; n7620_not
g47550 not n3264 ; n3264_not
g47551 not n8223 ; n8223_not
g47552 not n4407 ; n4407_not
g47553 not n4533 ; n4533_not
g47554 not n8151 ; n8151_not
g47555 not n5451 ; n5451_not
g47556 not n8205 ; n8205_not
g47557 not n8160 ; n8160_not
g47558 not n5550 ; n5550_not
g47559 not n2571 ; n2571_not
g47560 not n5532 ; n5532_not
g47561 not n3138 ; n3138_not
g47562 not n8331 ; n8331_not
g47563 not n5442 ; n5442_not
g47564 not n8313 ; n8313_not
g47565 not n4506 ; n4506_not
g47566 not n4452 ; n4452_not
g47567 not n8403 ; n8403_not
g47568 not n3165 ; n3165_not
g47569 not n5514 ; n5514_not
g47570 not n3093 ; n3093_not
g47571 not n4425 ; n4425_not
g47572 not n3174 ; n3174_not
g47573 not n3183 ; n3183_not
g47574 not n4524 ; n4524_not
g47575 not n5505 ; n5505_not
g47576 not n3192 ; n3192_not
g47577 not n8241 ; n8241_not
g47578 not n3048 ; n3048_not
g47579 not n4812 ; n4812_not
g47580 not n2652 ; n2652_not
g47581 not n4731 ; n4731_not
g47582 not n4803 ; n4803_not
g47583 not n5154 ; n5154_not
g47584 not n2526 ; n2526_not
g47585 not n5145 ; n5145_not
g47586 not n2490 ; n2490_not
g47587 not n6207 ; n6207_not
g47588 not n4740 ; n4740_not
g47589 not n2445 ; n2445_not
g47590 not n2454 ; n2454_not
g47591 not n9150 ; n9150_not
g47592 not n5028 ; n5028_not
g47593 not n2562 ; n2562_not
g47594 not n5046 ; n5046_not
g47595 not n7602 ; n7602_not
g47596 not n2616 ; n2616_not
g47597 not n6405 ; n6405_not
g47598 not n4830 ; n4830_not
g47599 not n4821 ; n4821_not
g47600 not n5316 ; n5316_not
g47601 not n4650 ; n4650_not
g47602 not n5325 ; n5325_not
g47603 not n6135 ; n6135_not
g47604 not n5334 ; n5334_not
g47605 not n9132 ; n9132_not
g47606 not n5343 ; n5343_not
g47607 not n9123 ; n9123_not
g47608 not n2904 ; n2904_not
g47609 not n9105 ; n9105_not
g47610 not n4560 ; n4560_not
g47611 not n5361 ; n5361_not
g47612 not n5370 ; n5370_not
g47613 not n9024 ; n9024_not
g47614 not n5406 ; n5406_not
g47615 not n5352 ; n5352_not
g47616 not n5424 ; n5424_not
g47617 not n5217 ; n5217_not
g47618 not n5226 ; n5226_not
g47619 not n9510 ; n9510_not
g47620 not n2823 ; n2823_not
g47621 not n9411 ; n9411_not
g47622 not n5235 ; n5235_not
g47623 not n2841 ; n2841_not
g47624 not n9330 ; n9330_not
g47625 not n9321 ; n9321_not
g47626 not n9303 ; n9303_not
g47627 not n5244 ; n5244_not
g47628 not n9312 ; n9312_not
g47629 not n9051 ; n9051_not
g47630 not n5262 ; n5262_not
g47631 not n9231 ; n9231_not
g47632 not n9222 ; n9222_not
g47633 not n9204 ; n9204_not
g47634 not n5307 ; n5307_not
g47635 not n6432 ; n6432_not
g47636 not n7332 ; n7332_not
g47637 not n6441 ; n6441_not
g47638 not n6450 ; n6450_not
g47639 not n7323 ; n7323_not
g47640 not n7314 ; n7314_not
g47641 not n6504 ; n6504_not
g47642 not n7224 ; n7224_not
g47643 not n6009 ; n6009_not
g47644 not n4056 ; n4056_not
g47645 not n7125 ; n7125_not
g47646 not n6108 ; n6108_not
g47647 not n6018 ; n6018_not
g47648 not n3840 ; n3840_not
g47649 not n6513 ; n6513_not
g47650 not n3543 ; n3543_not
g47651 not n3462 ; n3462_not
g47652 not n7503 ; n7503_not
g47653 not n5811 ; n5811_not
g47654 not n5901 ; n5901_not
g47655 not n4029 ; n4029_not
g47656 not n7413 ; n7413_not
g47657 not n6054 ; n6054_not
g47658 not n4245 ; n4245_not
g47659 not n4254 ; n4254_not
g47660 not n6423 ; n6423_not
g47661 not n3507 ; n3507_not
g47662 not n7350 ; n7350_not
g47663 not n3525 ; n3525_not
g47664 not n3480 ; n3480_not
g47665 not n4146 ; n4146_not
g47666 not n3705 ; n3705_not
g47667 not n4137 ; n4137_not
g47668 not n3723 ; n3723_not
g47669 not n4128 ; n4128_not
g47670 not n6621 ; n6621_not
g47671 not n6612 ; n6612_not
g47672 not n6522 ; n6522_not
g47673 not n6702 ; n6702_not
g47674 not n6801 ; n6801_not
g47675 not n7116 ; n7116_not
g47676 not n3633 ; n3633_not
g47677 not n7107 ; n7107_not
g47678 not n7071 ; n7071_not
g47679 not n6027 ; n6027_not
g47680 not n4065 ; n4065_not
g47681 not n6531 ; n6531_not
g47682 not n3831 ; n3831_not
g47683 not n6036 ; n6036_not
g47684 not n3570 ; n3570_not
g47685 not n6333 ; n6333_not
g47686 not n7017 ; n7017_not
g47687 not n3804 ; n3804_not
g47688 not n4155 ; n4155_not
g47689 not n3714 ; n3714_not
g47690 not n4083 ; n4083_not
g47691 not n3327 ; n3327_not
g47692 not n3354 ; n3354_not
g47693 not n7800 ; n7800_not
g47694 not n6162 ; n6162_not
g47695 not n5802 ; n5802_not
g47696 not n4344 ; n4344_not
g47697 not n3318 ; n3318_not
g47698 not n6306 ; n6306_not
g47699 not n4335 ; n4335_not
g47700 not n3372 ; n3372_not
g47701 not n4326 ; n4326_not
g47702 not n3282 ; n3282_not
g47703 not n6225 ; n6225_not
g47704 not n8115 ; n8115_not
g47705 not n2607 ; n2607_not
g47706 not n8070 ; n8070_not
g47707 not n3291 ; n3291_not
g47708 not n8016 ; n8016_not
g47709 not n5703 ; n5703_not
g47710 not n8025 ; n8025_not
g47711 not n6252 ; n6252_not
g47712 not n5730 ; n5730_not
g47713 not n4362 ; n4362_not
g47714 not n6234 ; n6234_not
g47715 not n3453 ; n3453_not
g47716 not n6126 ; n6126_not
g47717 not n3903 ; n3903_not
g47718 not n3444 ; n3444_not
g47719 not n7530 ; n7530_not
g47720 not n3426 ; n3426_not
g47721 not n3912 ; n3912_not
g47722 not n6315 ; n6315_not
g47723 not n4317 ; n4317_not
g47724 not n6144 ; n6144_not
g47725 not n6226 ; n6226_not
g47726 not n6280 ; n6280_not
g47727 not n2608 ; n2608_not
g47728 not n9133 ; n9133_not
g47729 not n5164 ; n5164_not
g47730 not n4912 ; n4912_not
g47731 not n6406 ; n6406_not
g47732 not n2572 ; n2572_not
g47733 not n5074 ; n5074_not
g47734 not n9700 ; n9700_not
g47735 not n6244 ; n6244_not
g47736 not n6361 ; n6361_not
g47737 not n2914 ; n2914_not
g47738 not n5182 ; n5182_not
g47739 not n6370 ; n6370_not
g47740 not n5173 ; n5173_not
g47741 not n5191 ; n5191_not
g47742 not n5056 ; n5056_not
g47743 not n6712 ; n6712_not
g47744 not n6460 ; n6460_not
g47745 not n2923 ; n2923_not
g47746 not n6442 ; n6442_not
g47747 not n6145 ; n6145_not
g47748 not n2932 ; n2932_not
g47749 not n5092 ; n5092_not
g47750 not n6163 ; n6163_not
g47751 not n2743 ; n2743_not
g47752 not n6172 ; n6172_not
g47753 not n6343 ; n6343_not
g47754 not n6541 ; n6541_not
g47755 not n6181 ; n6181_not
g47756 not n9052 ; n9052_not
g47757 not n6424 ; n6424_not
g47758 not n5038 ; n5038_not
g47759 not n5083 ; n5083_not
g47760 not n6091 ; n6091_not
g47761 not n8404 ; n8404_not
g47762 not n7540 ; n7540_not
g47763 not n5506 ; n5506_not
g47764 not n8431 ; n8431_not
g47765 not n6136 ; n6136_not
g47766 not n5821 ; n5821_not
g47767 not n3508 ; n3508_not
g47768 not n7513 ; n7513_not
g47769 not n5470 ; n5470_not
g47770 not n3328 ; n3328_not
g47771 not n5902 ; n5902_not
g47772 not n8512 ; n8512_not
g47773 not n8602 ; n8602_not
g47774 not n5452 ; n5452_not
g47775 not n8611 ; n8611_not
g47776 not n5434 ; n5434_not
g47777 not n8116 ; n8116_not
g47778 not n8143 ; n8143_not
g47779 not n5632 ; n5632_not
g47780 not n8215 ; n8215_not
g47781 not n5623 ; n5623_not
g47782 not n8233 ; n8233_not
g47783 not n8260 ; n8260_not
g47784 not n5641 ; n5641_not
g47785 not n8305 ; n8305_not
g47786 not n5740 ; n5740_not
g47787 not n5605 ; n5605_not
g47788 not n8314 ; n8314_not
g47789 not n5560 ; n5560_not
g47790 not n5803 ; n5803_not
g47791 not n8341 ; n8341_not
g47792 not n5542 ; n5542_not
g47793 not n8350 ; n8350_not
g47794 not n7630 ; n7630_not
g47795 not n5524 ; n5524_not
g47796 not n9223 ; n9223_not
g47797 not n7063 ; n7063_not
g47798 not n5254 ; n5254_not
g47799 not n7045 ; n7045_not
g47800 not n5245 ; n5245_not
g47801 not n6046 ; n6046_not
g47802 not n9322 ; n9322_not
g47803 not n7009 ; n7009_not
g47804 not n9340 ; n9340_not
g47805 not n2716 ; n2716_not
g47806 not n6901 ; n6901_not
g47807 not n9430 ; n9430_not
g47808 not n9502 ; n9502_not
g47809 not n9601 ; n9601_not
g47810 not n9610 ; n9610_not
g47811 not n9250 ; n9250_not
g47812 not n9511 ; n9511_not
g47813 not n5218 ; n5218_not
g47814 not n6811 ; n6811_not
g47815 not n7360 ; n7360_not
g47816 not n9007 ; n9007_not
g47817 not n7351 ; n7351_not
g47818 not n9016 ; n9016_not
g47819 not n5362 ; n5362_not
g47820 not n9034 ; n9034_not
g47821 not n7333 ; n7333_not
g47822 not n7432 ; n7432_not
g47823 not n9106 ; n9106_not
g47824 not n9115 ; n9115_not
g47825 not n7243 ; n7243_not
g47826 not n5344 ; n5344_not
g47827 not n7225 ; n7225_not
g47828 not n7216 ; n7216_not
g47829 not n9151 ; n9151_not
g47830 not n9160 ; n9160_not
g47831 not n7153 ; n7153_not
g47832 not n5326 ; n5326_not
g47833 not n7135 ; n7135_not
g47834 not n7072 ; n7072_not
g47835 not n5281 ; n5281_not
g47836 not n9241 ; n9241_not
g47837 not n3184 ; n3184_not
g47838 not n2563 ; n2563_not
g47839 not n4606 ; n4606_not
g47840 not n4840 ; n4840_not
g47841 not n3247 ; n3247_not
g47842 not n4417 ; n4417_not
g47843 not n3931 ; n3931_not
g47844 not n3256 ; n3256_not
g47845 not n4732 ; n4732_not
g47846 not n4354 ; n4354_not
g47847 not n4516 ; n4516_not
g47848 not n4723 ; n4723_not
g47849 not n3832 ; n3832_not
g47850 not n3616 ; n3616_not
g47851 not n2545 ; n2545_not
g47852 not n4048 ; n4048_not
g47853 not n4714 ; n4714_not
g47854 not n3625 ; n3625_not
g47855 not n4165 ; n4165_not
g47856 not n4282 ; n4282_not
g47857 not n4705 ; n4705_not
g47858 not n2860 ; n2860_not
g47859 not n4345 ; n4345_not
g47860 not n3751 ; n3751_not
g47861 not n3571 ; n3571_not
g47862 not n3544 ; n3544_not
g47863 not n3733 ; n3733_not
g47864 not n3463 ; n3463_not
g47865 not n4264 ; n4264_not
g47866 not n4660 ; n4660_not
g47867 not n4381 ; n4381_not
g47868 not n3535 ; n3535_not
g47869 not n4192 ; n4192_not
g47870 not n4183 ; n4183_not
g47871 not n3580 ; n3580_not
g47872 not n2851 ; n2851_not
g47873 not n3238 ; n3238_not
g47874 not n4318 ; n4318_not
g47875 not n4534 ; n4534_not
g47876 not n4174 ; n4174_not
g47877 not n4750 ; n4750_not
g47878 not n3409 ; n3409_not
g47879 not n3652 ; n3652_not
g47880 not n3319 ; n3319_not
g47881 not n2905 ; n2905_not
g47882 not n3346 ; n3346_not
g47883 not n4093 ; n4093_not
g47884 not n4291 ; n4291_not
g47885 not n3391 ; n3391_not
g47886 not n2815 ; n2815_not
g47887 not n2761 ; n2761_not
g47888 not n3139 ; n3139_not
g47889 not n3364 ; n3364_not
g47890 not n2842 ; n2842_not
g47891 not n3373 ; n3373_not
g47892 not n3904 ; n3904_not
g47893 not n3337 ; n3337_not
g47894 not n3661 ; n3661_not
g47895 not n4426 ; n4426_not
g47896 not n2437 ; n2437_not
g47897 not n3085 ; n3085_not
g47898 not n3715 ; n3715_not
g47899 not n4480 ; n4480_not
g47900 not n2509 ; n2509_not
g47901 not n2473 ; n2473_not
g47902 not n4642 ; n4642_not
g47903 not n3436 ; n3436_not
g47904 not n3292 ; n3292_not
g47905 not n4273 ; n4273_not
g47906 not n4147 ; n4147_not
g47907 not n4075 ; n4075_not
g47908 not n3850 ; n3850_not
g47909 not n8522 ; n8522_not
g47910 not n2852 ; n2852_not
g47911 not n3680 ; n3680_not
g47912 not n6740 ; n6740_not
g47913 not n2537 ; n2537_not
g47914 not n6074 ; n6074_not
g47915 not n2924 ; n2924_not
g47916 not n2843 ; n2843_not
g47917 not n6713 ; n6713_not
g47918 not n4661 ; n4661_not
g47919 not n8504 ; n8504_not
g47920 not n2690 ; n2690_not
g47921 not n6056 ; n6056_not
g47922 not n2636 ; n2636_not
g47923 not n6911 ; n6911_not
g47924 not n9332 ; n9332_not
g47925 not n9323 ; n9323_not
g47926 not n3725 ; n3725_not
g47927 not n8315 ; n8315_not
g47928 not n5714 ; n5714_not
g47929 not n6830 ; n6830_not
g47930 not n4652 ; n4652_not
g47931 not n6821 ; n6821_not
g47932 not n6227 ; n6227_not
g47933 not n4373 ; n4373_not
g47934 not n6236 ; n6236_not
g47935 not n3734 ; n3734_not
g47936 not n9341 ; n9341_not
g47937 not n9305 ; n9305_not
g47938 not n8531 ; n8531_not
g47939 not n5741 ; n5741_not
g47940 not n4337 ; n4337_not
g47941 not n3095 ; n3095_not
g47942 not n3743 ; n3743_not
g47943 not n4058 ; n4058_not
g47944 not n2762 ; n2762_not
g47945 not n6434 ; n6434_not
g47946 not n6326 ; n6326_not
g47947 not n5561 ; n5561_not
g47948 not n5543 ; n5543_not
g47949 not n6263 ; n6263_not
g47950 not n5651 ; n5651_not
g47951 not n7451 ; n7451_not
g47952 not n6506 ; n6506_not
g47953 not n3842 ; n3842_not
g47954 not n4508 ; n4508_not
g47955 not n5516 ; n5516_not
g47956 not n6533 ; n6533_not
g47957 not n2870 ; n2870_not
g47958 not n4427 ; n4427_not
g47959 not n3923 ; n3923_not
g47960 not n4454 ; n4454_not
g47961 not n6344 ; n6344_not
g47962 not n5606 ; n5606_not
g47963 not n3905 ; n3905_not
g47964 not n6308 ; n6308_not
g47965 not n6317 ; n6317_not
g47966 not n6191 ; n6191_not
g47967 not n3383 ; n3383_not
g47968 not n9161 ; n9161_not
g47969 not n4418 ; n4418_not
g47970 not n9215 ; n9215_not
g47971 not n5633 ; n5633_not
g47972 not n6407 ; n6407_not
g47973 not n6425 ; n6425_not
g47974 not n6290 ; n6290_not
g47975 not n9116 ; n9116_not
g47976 not n3860 ; n3860_not
g47977 not n4553 ; n4553_not
g47978 not n5318 ; n5318_not
g47979 not n6605 ; n6605_not
g47980 not n6209 ; n6209_not
g47981 not n2483 ; n2483_not
g47982 not n5426 ; n5426_not
g47983 not n8720 ; n8720_not
g47984 not n6704 ; n6704_not
g47985 not n5417 ; n5417_not
g47986 not n6164 ; n6164_not
g47987 not n3761 ; n3761_not
g47988 not n3752 ; n3752_not
g47989 not n8711 ; n8711_not
g47990 not n6722 ; n6722_not
g47991 not n6524 ; n6524_not
g47992 not n6254 ; n6254_not
g47993 not n6560 ; n6560_not
g47994 not n3815 ; n3815_not
g47995 not n2960 ; n2960_not
g47996 not n5480 ; n5480_not
g47997 not n5471 ; n5471_not
g47998 not n4535 ; n4535_not
g47999 not n6173 ; n6173_not
g48000 not n2915 ; n2915_not
g48001 not n4544 ; n4544_not
g48002 not n9242 ; n9242_not
g48003 not n8810 ; n8810_not
g48004 not n5075 ; n5075_not
g48005 not n7415 ; n7415_not
g48006 not n5921 ; n5921_not
g48007 not n2564 ; n2564_not
g48008 not n8153 ; n8153_not
g48009 not n5930 ; n5930_not
g48010 not n3266 ; n3266_not
g48011 not n6272 ; n6272_not
g48012 not n5039 ; n5039_not
g48013 not n3473 ; n3473_not
g48014 not n3455 ; n3455_not
g48015 not n8090 ; n8090_not
g48016 not n4706 ; n4706_not
g48017 not n2438 ; n2438_not
g48018 not n7334 ; n7334_not
g48019 not n3527 ; n3527_not
g48020 not n4805 ; n4805_not
g48021 not n9314 ; n9314_not
g48022 not n3518 ; n3518_not
g48023 not n3239 ; n3239_not
g48024 not n7370 ; n7370_not
g48025 not n9440 ; n9440_not
g48026 not n5084 ; n5084_not
g48027 not n3248 ; n3248_not
g48028 not n4832 ; n4832_not
g48029 not n7406 ; n7406_not
g48030 not n3482 ; n3482_not
g48031 not n8009 ; n8009_not
g48032 not n3338 ; n3338_not
g48033 not n9602 ; n9602_not
g48034 not n9260 ; n9260_not
g48035 not n7622 ; n7622_not
g48036 not n7802 ; n7802_not
g48037 not n3356 ; n3356_not
g48038 not n3374 ; n3374_not
g48039 not n2456 ; n2456_not
g48040 not n4922 ; n4922_not
g48041 not n3365 ; n3365_not
g48042 not n4931 ; n4931_not
g48043 not n7721 ; n7721_not
g48044 not n7712 ; n7712_not
g48045 not n3464 ; n3464_not
g48046 not n7505 ; n7505_not
g48047 not n4283 ; n4283_not
g48048 not n7433 ; n7433_not
g48049 not n8054 ; n8054_not
g48050 not n8063 ; n8063_not
g48051 not n5903 ; n5903_not
g48052 not n3428 ; n3428_not
g48053 not n7541 ; n7541_not
g48054 not n2933 ; n2933_not
g48055 not n8036 ; n8036_not
g48056 not n7901 ; n7901_not
g48057 not n9611 ; n9611_not
g48058 not n6038 ; n6038_not
g48059 not n4355 ; n4355_not
g48060 not n7145 ; n7145_not
g48061 not n8306 ; n8306_not
g48062 not n7154 ; n7154_not
g48063 not n3185 ; n3185_not
g48064 not n4742 ; n4742_not
g48065 not n7172 ; n7172_not
g48066 not n4175 ; n4175_not
g48067 not n6029 ; n6029_not
g48068 not n2591 ; n2591_not
g48069 not n3194 ; n3194_not
g48070 not n3581 ; n3581_not
g48071 not n4184 ; n4184_not
g48072 not n2573 ; n2573_not
g48073 not n5183 ; n5183_not
g48074 not n9800 ; n9800_not
g48075 not n5705 ; n5705_not
g48076 not n4094 ; n4094_not
g48077 not n5237 ; n5237_not
g48078 not n6065 ; n6065_not
g48079 not n5273 ; n5273_not
g48080 not n7019 ; n7019_not
g48081 not n4670 ; n4670_not
g48082 not n5255 ; n5255_not
g48083 not n7082 ; n7082_not
g48084 not n2645 ; n2645_not
g48085 not n3644 ; n3644_not
g48086 not n2528 ; n2528_not
g48087 not n7109 ; n7109_not
g48088 not n7118 ; n7118_not
g48089 not n4157 ; n4157_not
g48090 not n8324 ; n8324_not
g48091 not n2834 ; n2834_not
g48092 not n6416 ; n6416_not
g48093 not n2807 ; n2807_not
g48094 not n3167 ; n3167_not
g48095 not n5129 ; n5129_not
g48096 not n9044 ; n9044_not
g48097 not n7262 ; n7262_not
g48098 not n8108 ; n8108_not
g48099 not n4229 ; n4229_not
g48100 not n7253 ; n7253_not
g48101 not n8180 ; n8180_not
g48102 not n3563 ; n3563_not
g48103 not n7235 ; n7235_not
g48104 not n7226 ; n7226_not
g48105 not n4760 ; n4760_not
g48106 not n3572 ; n3572_not
g48107 not n9612 ; n9612_not
g48108 not n4293 ; n4293_not
g48109 not n9342 ; n9342_not
g48110 not n6048 ; n6048_not
g48111 not n9630 ; n9630_not
g48112 not n6228 ; n6228_not
g48113 not n4275 ; n4275_not
g48114 not n6057 ; n6057_not
g48115 not n6066 ; n6066_not
g48116 not n2529 ; n2529_not
g48117 not n9252 ; n9252_not
g48118 not n4257 ; n4257_not
g48119 not n6093 ; n6093_not
g48120 not n3393 ; n3393_not
g48121 not n6219 ; n6219_not
g48122 not n5940 ; n5940_not
g48123 not n2835 ; n2835_not
g48124 not n9036 ; n9036_not
g48125 not n6156 ; n6156_not
g48126 not n6246 ; n6246_not
g48127 not n4167 ; n4167_not
g48128 not n9504 ; n9504_not
g48129 not n6129 ; n6129_not
g48130 not n4194 ; n4194_not
g48131 not n4086 ; n4086_not
g48132 not n3933 ; n3933_not
g48133 not n4176 ; n4176_not
g48134 not n5814 ; n5814_not
g48135 not n9441 ; n9441_not
g48136 not n9216 ; n9216_not
g48137 not n2871 ; n2871_not
g48138 not n9351 ; n9351_not
g48139 not n6165 ; n6165_not
g48140 not n6147 ; n6147_not
g48141 not n4149 ; n4149_not
g48142 not n3951 ; n3951_not
g48143 not n4077 ; n4077_not
g48144 not n7254 ; n7254_not
g48145 not n7245 ; n7245_not
g48146 not n7209 ; n7209_not
g48147 not n3195 ; n3195_not
g48148 not n8271 ; n8271_not
g48149 not n3591 ; n3591_not
g48150 not n7191 ; n7191_not
g48151 not n7137 ; n7137_not
g48152 not n7182 ; n7182_not
g48153 not n7164 ; n7164_not
g48154 not n7155 ; n7155_not
g48155 not n8172 ; n8172_not
g48156 not n8316 ; n8316_not
g48157 not n7128 ; n7128_not
g48158 not n3159 ; n3159_not
g48159 not n7029 ; n7029_not
g48160 not n8343 ; n8343_not
g48161 not n3654 ; n3654_not
g48162 not n3555 ; n3555_not
g48163 not n3663 ; n3663_not
g48164 not n8352 ; n8352_not
g48165 not n8370 ; n8370_not
g48166 not n3690 ; n3690_not
g48167 not n7722 ; n7722_not
g48168 not n7731 ; n7731_not
g48169 not n7542 ; n7542_not
g48170 not n7605 ; n7605_not
g48171 not n7821 ; n7821_not
g48172 not n7425 ; n7425_not
g48173 not n7920 ; n7920_not
g48174 not n7911 ; n7911_not
g48175 not n7551 ; n7551_not
g48176 not n7461 ; n7461_not
g48177 not n7533 ; n7533_not
g48178 not n8064 ; n8064_not
g48179 not n3438 ; n3438_not
g48180 not n8073 ; n8073_not
g48181 not n8082 ; n8082_not
g48182 not n8118 ; n8118_not
g48183 not n7263 ; n7263_not
g48184 not n7281 ; n7281_not
g48185 not n7308 ; n7308_not
g48186 not n7317 ; n7317_not
g48187 not n3456 ; n3456_not
g48188 not n3537 ; n3537_not
g48189 not n7326 ; n7326_not
g48190 not n8217 ; n8217_not
g48191 not n3492 ; n3492_not
g48192 not n8190 ; n8190_not
g48193 not n7371 ; n7371_not
g48194 not n7614 ; n7614_not
g48195 not n7434 ; n7434_not
g48196 not n7443 ; n7443_not
g48197 not n3258 ; n3258_not
g48198 not n8145 ; n8145_not
g48199 not n8811 ; n8811_not
g48200 not n6633 ; n6633_not
g48201 not n8820 ; n8820_not
g48202 not n6624 ; n6624_not
g48203 not n8613 ; n8613_not
g48204 not n7641 ; n7641_not
g48205 not n3807 ; n3807_not
g48206 not n6282 ; n6282_not
g48207 not n9009 ; n9009_not
g48208 not n6552 ; n6552_not
g48209 not n3825 ; n3825_not
g48210 not n3834 ; n3834_not
g48211 not n2943 ; n2943_not
g48212 not n9063 ; n9063_not
g48213 not n2745 ; n2745_not
g48214 not n9072 ; n9072_not
g48215 not n9090 ; n9090_not
g48216 not n6453 ; n6453_not
g48217 not n3861 ; n3861_not
g48218 not n9108 ; n9108_not
g48219 not n6426 ; n6426_not
g48220 not n3870 ; n3870_not
g48221 not n9135 ; n9135_not
g48222 not n9153 ; n9153_not
g48223 not n6354 ; n6354_not
g48224 not n6363 ; n6363_not
g48225 not n9171 ; n9171_not
g48226 not n6318 ; n6318_not
g48227 not n3096 ; n3096_not
g48228 not n8406 ; n8406_not
g48229 not n8433 ; n8433_not
g48230 not n8442 ; n8442_not
g48231 not n6921 ; n6921_not
g48232 not n3087 ; n3087_not
g48233 not n3069 ; n3069_not
g48234 not n6903 ; n6903_not
g48235 not n8541 ; n8541_not
g48236 not n8550 ; n8550_not
g48237 not n3717 ; n3717_not
g48238 not n6840 ; n6840_not
g48239 not n8802 ; n8802_not
g48240 not n6651 ; n6651_not
g48241 not n6660 ; n6660_not
g48242 not n8730 ; n8730_not
g48243 not n8712 ; n8712_not
g48244 not n3762 ; n3762_not
g48245 not n6714 ; n6714_not
g48246 not n6732 ; n6732_not
g48247 not n8640 ; n8640_not
g48248 not n3744 ; n3744_not
g48249 not n6417 ; n6417_not
g48250 not n6813 ; n6813_not
g48251 not n4518 ; n4518_not
g48252 not n6273 ; n6273_not
g48253 not n9711 ; n9711_not
g48254 not n5508 ; n5508_not
g48255 not n4671 ; n4671_not
g48256 not n5751 ; n5751_not
g48257 not n2547 ; n2547_not
g48258 not n5454 ; n5454_not
g48259 not n4851 ; n4851_not
g48260 not n4446 ; n4446_not
g48261 not n4842 ; n4842_not
g48262 not n5256 ; n5256_not
g48263 not n2646 ; n2646_not
g48264 not n5733 ; n5733_not
g48265 not n5526 ; n5526_not
g48266 not n5058 ; n5058_not
g48267 not n4644 ; n4644_not
g48268 not n4554 ; n4554_not
g48269 not n6192 ; n6192_not
g48270 not n2673 ; n2673_not
g48271 not n4653 ; n4653_not
g48272 not n9144 ; n9144_not
g48273 not n4536 ; n4536_not
g48274 not n4545 ; n4545_not
g48275 not n9801 ; n9801_not
g48276 not n5472 ; n5472_not
g48277 not n4662 ; n4662_not
g48278 not n9810 ; n9810_not
g48279 not n3447 ; n3447_not
g48280 not n5283 ; n5283_not
g48281 not n4356 ; n4356_not
g48282 not n4860 ; n4860_not
g48283 not n4473 ; n4473_not
g48284 not n5193 ; n5193_not
g48285 not n4752 ; n4752_not
g48286 not n2484 ; n2484_not
g48287 not n4455 ; n4455_not
g48288 not n5661 ; n5661_not
g48289 not n2772 ; n2772_not
g48290 not n5157 ; n5157_not
g48291 not n7452 ; n7452_not
g48292 not n5535 ; n5535_not
g48293 not n5175 ; n5175_not
g48294 not n5625 ; n5625_not
g48295 not n4437 ; n4437_not
g48296 not n5076 ; n5076_not
g48297 not n4491 ; n4491_not
g48298 not n4707 ; n4707_not
g48299 not n7506 ; n7506_not
g48300 not n4824 ; n4824_not
g48301 not n4725 ; n4725_not
g48302 not n4383 ; n4383_not
g48303 not n5094 ; n5094_not
g48304 not n4815 ; n4815_not
g48305 not n4734 ; n4734_not
g48306 not n2727 ; n2727_not
g48307 not n9414 ; n9414_not
g48308 not n2709 ; n2709_not
g48309 not n4617 ; n4617_not
g48310 not n2439 ; n2439_not
g48311 not n5553 ; n5553_not
g48312 not n4608 ; n4608_not
g48313 not n2628 ; n2628_not
g48314 not n5346 ; n5346_not
g48315 not n2592 ; n2592_not
g48316 not n4572 ; n4572_not
g48317 not n5391 ; n5391_not
g48318 not n5373 ; n5373_not
g48319 not n9702 ; n9702_not
g48320 not n5364 ; n5364_not
g48321 not n4941 ; n4941_not
g48322 not n4950 ; n4950_not
g48323 not n4527 ; n4527_not
g48324 not n5850 ; n5850_not
g48325 not n4590 ; n4590_not
g48326 not n5832 ; n5832_not
g48327 not n5418 ; n5418_not
g48328 not n2619 ; n2619_not
g48329 not n4581 ; n4581_not
g48330 not n5436 ; n5436_not
g48331 not n2475 ; n2475_not
g48332 not n5823 ; n5823_not
g48333 not n5328 ; n5328_not
g48334 not n7570 ; n7570_not
g48335 not n3871 ; n3871_not
g48336 not n3448 ; n3448_not
g48337 not n3862 ; n3862_not
g48338 not n4744 ; n4744_not
g48339 not n4726 ; n4726_not
g48340 not n6445 ; n6445_not
g48341 not n6841 ; n6841_not
g48342 not n3385 ; n3385_not
g48343 not n8317 ; n8317_not
g48344 not n7471 ; n7471_not
g48345 not n6436 ; n6436_not
g48346 not n8308 ; n8308_not
g48347 not n2692 ; n2692_not
g48348 not n6193 ; n6193_not
g48349 not n4483 ; n4483_not
g48350 not n7129 ; n7129_not
g48351 not n3727 ; n3727_not
g48352 not n6427 ; n6427_not
g48353 not n7147 ; n7147_not
g48354 not n2908 ; n2908_not
g48355 not n2755 ; n2755_not
g48356 not n2926 ; n2926_not
g48357 not n6724 ; n6724_not
g48358 not n4456 ; n4456_not
g48359 not n3907 ; n3907_not
g48360 not n9181 ; n9181_not
g48361 not n3916 ; n3916_not
g48362 not n6337 ; n6337_not
g48363 not n8632 ; n8632_not
g48364 not n9190 ; n9190_not
g48365 not n2683 ; n2683_not
g48366 not n6328 ; n6328_not
g48367 not n7228 ; n7228_not
g48368 not n3394 ; n3394_not
g48369 not n4762 ; n4762_not
g48370 not n8623 ; n8623_not
g48371 not n6139 ; n6139_not
g48372 not n7174 ; n7174_not
g48373 not n6742 ; n6742_not
g48374 not n9127 ; n9127_not
g48375 not n8263 ; n8263_not
g48376 not n2593 ; n2593_not
g48377 not n6265 ; n6265_not
g48378 not n8281 ; n8281_not
g48379 not n6373 ; n6373_not
g48380 not n6832 ; n6832_not
g48381 not n8614 ; n8614_not
g48382 not n4465 ; n4465_not
g48383 not n2773 ; n2773_not
g48384 not n6184 ; n6184_not
g48385 not n5185 ; n5185_not
g48386 not n6805 ; n6805_not
g48387 not n8407 ; n8407_not
g48388 not n5491 ; n5491_not
g48389 not n3808 ; n3808_not
g48390 not n5428 ; n5428_not
g48391 not n3691 ; n3691_not
g48392 not n2674 ; n2674_not
g48393 not n6562 ; n6562_not
g48394 not n6652 ; n6652_not
g48395 not n3817 ; n3817_not
g48396 not n5275 ; n5275_not
g48397 not n4618 ; n4618_not
g48398 not n7039 ; n7039_not
g48399 not n3718 ; n3718_not
g48400 not n8524 ; n8524_not
g48401 not n8506 ; n8506_not
g48402 not n2971 ; n2971_not
g48403 not n6643 ; n6643_not
g48404 not n5329 ; n5329_not
g48405 not n6625 ; n6625_not
g48406 not n6913 ; n6913_not
g48407 not n5455 ; n5455_not
g48408 not n8461 ; n8461_not
g48409 not n8452 ; n8452_not
g48410 not n8425 ; n8425_not
g48411 not n4537 ; n4537_not
g48412 not n8416 ; n8416_not
g48413 not n2647 ; n2647_not
g48414 not n3628 ; n3628_not
g48415 not n2719 ; n2719_not
g48416 not n6472 ; n6472_not
g48417 not n2728 ; n2728_not
g48418 not n9091 ; n9091_not
g48419 not n7417 ; n7417_not
g48420 not n3637 ; n3637_not
g48421 not n6463 ; n6463_not
g48422 not n8326 ; n8326_not
g48423 not n6454 ; n6454_not
g48424 not n3619 ; n3619_not
g48425 not n3169 ; n3169_not
g48426 not n5266 ; n5266_not
g48427 not n8731 ; n8731_not
g48428 not n5518 ; n5518_not
g48429 not n2953 ; n2953_not
g48430 not n6517 ; n6517_not
g48431 not n7057 ; n7057_not
g48432 not n3781 ; n3781_not
g48433 not n8344 ; n8344_not
g48434 not n3844 ; n3844_not
g48435 not n9037 ; n9037_not
g48436 not n6580 ; n6580_not
g48437 not n8551 ; n8551_not
g48438 not n8722 ; n8722_not
g48439 not n9055 ; n9055_not
g48440 not n3646 ; n3646_not
g48441 not n7093 ; n7093_not
g48442 not n8335 ; n8335_not
g48443 not n3268 ; n3268_not
g48444 not n5770 ; n5770_not
g48445 not n4159 ; n4159_not
g48446 not n4096 ; n4096_not
g48447 not n9109 ; n9109_not
g48448 not n9820 ; n9820_not
g48449 not n9802 ; n9802_not
g48450 not n4861 ; n4861_not
g48451 not n3286 ; n3286_not
g48452 not n4195 ; n4195_not
g48453 not n9361 ; n9361_not
g48454 not n2539 ; n2539_not
g48455 not n9370 ; n9370_not
g48456 not n7507 ; n7507_not
g48457 not n9424 ; n9424_not
g48458 not n8065 ; n8065_not
g48459 not n9433 ; n9433_not
g48460 not n5725 ; n5725_not
g48461 not n3475 ; n3475_not
g48462 not n4069 ; n4069_not
g48463 not n4366 ; n4366_not
g48464 not n4771 ; n4771_not
g48465 not n6094 ; n6094_not
g48466 not n8155 ; n8155_not
g48467 not n6157 ; n6157_not
g48468 not n5743 ; n5743_not
g48469 not n6085 ; n6085_not
g48470 not n4852 ; n4852_not
g48471 not n4087 ; n4087_not
g48472 not n6076 ; n6076_not
g48473 not n7444 ; n7444_not
g48474 not n8146 ; n8146_not
g48475 not n9901 ; n9901_not
g48476 not n9703 ; n9703_not
g48477 not n6058 ; n6058_not
g48478 not n5761 ; n5761_not
g48479 not n7462 ; n7462_not
g48480 not n9541 ; n9541_not
g48481 not n4285 ; n4285_not
g48482 not n9730 ; n9730_not
g48483 not n3358 ; n3358_not
g48484 not n4906 ; n4906_not
g48485 not n9118 ; n9118_not
g48486 not n7660 ; n7660_not
g48487 not n9613 ; n9613_not
g48488 not n9721 ; n9721_not
g48489 not n7723 ; n7723_not
g48490 not n9631 ; n9631_not
g48491 not n5815 ; n5815_not
g48492 not n3376 ; n3376_not
g48493 not n8119 ; n8119_not
g48494 not n5950 ; n5950_not
g48495 not n9460 ; n9460_not
g48496 not n9451 ; n9451_not
g48497 not n7561 ; n7561_not
g48498 not n5824 ; n5824_not
g48499 not n2827 ; n2827_not
g48500 not n5833 ; n5833_not
g48501 not n7840 ; n7840_not
g48502 not n4960 ; n4960_not
g48503 not n7804 ; n7804_not
g48504 not n7246 ; n7246_not
g48505 not n2485 ; n2485_not
g48506 not n9226 ; n9226_not
g48507 not n8209 ; n8209_not
g48508 not n5095 ; n5095_not
g48509 not n7345 ; n7345_not
g48510 not n9235 ; n9235_not
g48511 not n7336 ; n7336_not
g48512 not n7273 ; n7273_not
g48513 not n3529 ; n3529_not
g48514 not n7291 ; n7291_not
g48515 not n9280 ; n9280_not
g48516 not n5563 ; n5563_not
g48517 not n4636 ; n4636_not
g48518 not n2575 ; n2575_not
g48519 not n8236 ; n8236_not
g48520 not n9244 ; n9244_not
g48521 not n8227 ; n8227_not
g48522 not n6490 ; n6490_not
g48523 not n8128 ; n8128_not
g48524 not n9262 ; n9262_not
g48525 not n3547 ; n3547_not
g48526 not n9334 ; n9334_not
g48527 not n4834 ; n4834_not
g48528 not n3925 ; n3925_not
g48529 not n2881 ; n2881_not
g48530 not n4375 ; n4375_not
g48531 not n9325 ; n9325_not
g48532 not n7237 ; n7237_not
g48533 not n8254 ; n8254_not
g48534 not n7571 ; n7571_not
g48535 not n4772 ; n4772_not
g48536 not n8255 ; n8255_not
g48537 not n7193 ; n7193_not
g48538 not n8543 ; n8543_not
g48539 not n9209 ; n9209_not
g48540 not n5177 ; n5177_not
g48541 not n7706 ; n7706_not
g48542 not n9722 ; n9722_not
g48543 not n8291 ; n8291_not
g48544 not n6905 ; n6905_not
g48545 not n2927 ; n2927_not
g48546 not n3557 ; n3557_not
g48547 not n4781 ; n4781_not
g48548 not n8093 ; n8093_not
g48549 not n3728 ; n3728_not
g48550 not n7229 ; n7229_not
g48551 not n4871 ; n4871_not
g48552 not n6419 ; n6419_not
g48553 not n4628 ; n4628_not
g48554 not n7238 ; n7238_not
g48555 not n7850 ; n7850_not
g48556 not n5168 ; n5168_not
g48557 not n8516 ; n8516_not
g48558 not n3575 ; n3575_not
g48559 not n7724 ; n7724_not
g48560 not n2738 ; n2738_not
g48561 not n4592 ; n4592_not
g48562 not n8246 ; n8246_not
g48563 not n2585 ; n2585_not
g48564 not n3737 ; n3737_not
g48565 not n3719 ; n3719_not
g48566 not n7634 ; n7634_not
g48567 not n6761 ; n6761_not
g48568 not n6860 ; n6860_not
g48569 not n8561 ; n8561_not
g48570 not n4754 ; n4754_not
g48571 not n3197 ; n3197_not
g48572 not n4952 ; n4952_not
g48573 not n6815 ; n6815_not
g48574 not n7418 ; n7418_not
g48575 not n7283 ; n7283_not
g48576 not n8237 ; n8237_not
g48577 not n3584 ; n3584_not
g48578 not n4934 ; n4934_not
g48579 not n5195 ; n5195_not
g48580 not n7760 ; n7760_not
g48581 not n4970 ; n4970_not
g48582 not n6842 ; n6842_not
g48583 not n4691 ; n4691_not
g48584 not n6356 ; n6356_not
g48585 not n7058 ; n7058_not
g48586 not n8192 ; n8192_not
g48587 not n4673 ; n4673_not
g48588 not n7454 ; n7454_not
g48589 not n7049 ; n7049_not
g48590 not n7373 ; n7373_not
g48591 not n7463 ; n7463_not
g48592 not n5267 ; n5267_not
g48593 not n8354 ; n8354_not
g48594 not n8174 ; n8174_not
g48595 not n2639 ; n2639_not
g48596 not n3674 ; n3674_not
g48597 not n4817 ; n4817_not
g48598 not n8903 ; n8903_not
g48599 not n7346 ; n7346_not
g48600 not n6194 ; n6194_not
g48601 not n3638 ; n3638_not
g48602 not n3485 ; n3485_not
g48603 not n5249 ; n5249_not
g48604 not n7076 ; n7076_not
g48605 not n8183 ; n8183_not
g48606 not n4826 ; n4826_not
g48607 not n4844 ; n4844_not
g48608 not n4709 ; n4709_not
g48609 not n4853 ; n4853_not
g48610 not n5258 ; n5258_not
g48611 not n7391 ; n7391_not
g48612 not n3656 ; n3656_not
g48613 not n3089 ; n3089_not
g48614 not n4790 ; n4790_not
g48615 not n4880 ; n4880_not
g48616 not n3665 ; n3665_not
g48617 not n7508 ; n7508_not
g48618 not n6923 ; n6923_not
g48619 not n7157 ; n7157_not
g48620 not n6392 ; n6392_not
g48621 not n2747 ; n2747_not
g48622 not n7436 ; n7436_not
g48623 not n4646 ; n4646_not
g48624 not n3296 ; n3296_not
g48625 not n6491 ; n6491_not
g48626 not n3539 ; n3539_not
g48627 not n3683 ; n3683_not
g48628 not n8372 ; n8372_not
g48629 not n7337 ; n7337_not
g48630 not n5285 ; n5285_not
g48631 not n3467 ; n3467_not
g48632 not n7481 ; n7481_not
g48633 not n2648 ; n2648_not
g48634 not n7148 ; n7148_not
g48635 not n8408 ; n8408_not
g48636 not n8417 ; n8417_not
g48637 not n7490 ; n7490_not
g48638 not n4736 ; n4736_not
g48639 not n2666 ; n2666_not
g48640 not n2576 ; n2576_not
g48641 not n6077 ; n6077_not
g48642 not n9911 ; n9911_not
g48643 not n6509 ; n6509_not
g48644 not n5852 ; n5852_not
g48645 not n9038 ; n9038_not
g48646 not n9047 ; n9047_not
g48647 not n6086 ; n6086_not
g48648 not n4277 ; n4277_not
g48649 not n4079 ; n4079_not
g48650 not n9065 ; n9065_not
g48651 not n4367 ; n4367_not
g48652 not n9920 ; n9920_not
g48653 not n5726 ; n5726_not
g48654 not n4493 ; n4493_not
g48655 not n9335 ; n9335_not
g48656 not n6464 ; n6464_not
g48657 not n5717 ; n5717_not
g48658 not n3944 ; n3944_not
g48659 not n3746 ; n3746_not
g48660 not n4484 ; n4484_not
g48661 not n3809 ; n3809_not
g48662 not n3791 ; n3791_not
g48663 not n5780 ; n5780_not
g48664 not n5483 ; n5483_not
g48665 not n2837 ; n2837_not
g48666 not n5492 ; n5492_not
g48667 not n5942 ; n5942_not
g48668 not n9803 ; n9803_not
g48669 not n4529 ; n4529_not
g48670 not n4349 ; n4349_not
g48671 not n6554 ; n6554_not
g48672 not n9830 ; n9830_not
g48673 not n4358 ; n4358_not
g48674 not n6329 ; n6329_not
g48675 not n3386 ; n3386_not
g48676 not n2954 ; n2954_not
g48677 not n6518 ; n6518_not
g48678 not n6536 ; n6536_not
g48679 not n3827 ; n3827_not
g48680 not n3962 ; n3962_not
g48681 not n5474 ; n5474_not
g48682 not n4097 ; n4097_not
g48683 not n5753 ; n5753_not
g48684 not n3971 ; n3971_not
g48685 not n9164 ; n9164_not
g48686 not n9173 ; n9173_not
g48687 not n2891 ; n2891_not
g48688 not n6365 ; n6365_not
g48689 not n5681 ; n5681_not
g48690 not n6284 ; n6284_not
g48691 not n3917 ; n3917_not
g48692 not n2882 ; n2882_not
g48693 not n4439 ; n4439_not
g48694 not n5618 ; n5618_not
g48695 not n5627 ; n5627_not
g48696 not n2774 ; n2774_not
g48697 not n9902 ; n9902_not
g48698 not n6293 ; n6293_not
g48699 not n5636 ; n5636_not
g48700 not n2792 ; n2792_not
g48701 not n7472 ; n7472_not
g48702 not n3935 ; n3935_not
g48703 not n9236 ; n9236_not
g48704 not n6248 ; n6248_not
g48705 not n5663 ; n5663_not
g48706 not n6455 ; n6455_not
g48707 not n2909 ; n2909_not
g48708 not n3755 ; n3755_not
g48709 not n2486 ; n2486_not
g48710 not n6446 ; n6446_not
g48711 not n2729 ; n2729_not
g48712 not n5564 ; n5564_not
g48713 not n3863 ; n3863_not
g48714 not n5573 ; n5573_not
g48715 not n7643 ; n7643_not
g48716 not n4385 ; n4385_not
g48717 not n3980 ; n3980_not
g48718 not n2756 ; n2756_not
g48719 not n9128 ; n9128_not
g48720 not n3881 ; n3881_not
g48721 not n5672 ; n5672_not
g48722 not n5690 ; n5690_not
g48723 not n9290 ; n9290_not
g48724 not n4394 ; n4394_not
g48725 not n9272 ; n9272_not
g48726 not n6374 ; n6374_not
g48727 not n5393 ; n5393_not
g48728 not n8714 ; n8714_not
g48729 not n2819 ; n2819_not
g48730 not n4574 ; n4574_not
g48731 not n9740 ; n9740_not
g48732 not n2981 ; n2981_not
g48733 not n8741 ; n8741_not
g48734 not n5915 ; n5915_not
g48735 not n6527 ; n6527_not
g48736 not n5933 ; n5933_not
g48737 not n5438 ; n5438_not
g48738 not n6635 ; n6635_not
g48739 not n9461 ; n9461_not
g48740 not n4556 ; n4556_not
g48741 not n5825 ; n5825_not
g48742 not n4295 ; n4295_not
g48743 not n9704 ; n9704_not
g48744 not n8633 ; n8633_not
g48745 not n9605 ; n9605_not
g48746 not n9281 ; n9281_not
g48747 not n5870 ; n5870_not
g48748 not n9641 ; n9641_not
g48749 not n9614 ; n9614_not
g48750 not n2684 ; n2684_not
g48751 not n5384 ; n5384_not
g48752 not n5843 ; n5843_not
g48753 not n5294 ; n5294_not
g48754 not n6743 ; n6743_not
g48755 not n6734 ; n6734_not
g48756 not n9560 ; n9560_not
g48757 not n9542 ; n9542_not
g48758 not n5906 ; n5906_not
g48759 not n9443 ; n9443_not
g48760 not n9425 ; n9425_not
g48761 not n4268 ; n4268_not
g48762 not n5456 ; n5456_not
g48763 not n6572 ; n6572_not
g48764 not n6383 ; n6383_not
g48765 not n2828 ; n2828_not
g48766 not n2928 ; n2928_not
g48767 not n5682 ; n5682_not
g48768 not n9129 ; n9129_not
g48769 not n9723 ; n9723_not
g48770 not n9750 ; n9750_not
g48771 not n2487 ; n2487_not
g48772 not n5835 ; n5835_not
g48773 not n9426 ; n9426_not
g48774 not n3279 ; n3279_not
g48775 not n6771 ; n6771_not
g48776 not n9273 ; n9273_not
g48777 not n5790 ; n5790_not
g48778 not n9039 ; n9039_not
g48779 not n7428 ; n7428_not
g48780 not n9408 ; n9408_not
g48781 not n2865 ; n2865_not
g48782 not n6195 ; n6195_not
g48783 not n5691 ; n5691_not
g48784 not n7482 ; n7482_not
g48785 not n3486 ; n3486_not
g48786 not n7635 ; n7635_not
g48787 not n4881 ; n4881_not
g48788 not n9390 ; n9390_not
g48789 not n6249 ; n6249_not
g48790 not n3189 ; n3189_not
g48791 not n5808 ; n5808_not
g48792 not n9246 ; n9246_not
g48793 not n7626 ; n7626_not
g48794 not n7293 ; n7293_not
g48795 not n3954 ; n3954_not
g48796 not n7356 ; n7356_not
g48797 not n5862 ; n5862_not
g48798 not n9633 ; n9633_not
g48799 not n5880 ; n5880_not
g48800 not n3549 ; n3549_not
g48801 not n9624 ; n9624_not
g48802 not n7473 ; n7473_not
g48803 not n3369 ; n3369_not
g48804 not n4872 ; n4872_not
g48805 not n3288 ; n3288_not
g48806 not n2793 ; n2793_not
g48807 not n9264 ; n9264_not
g48808 not n7860 ; n7860_not
g48809 not n4908 ; n4908_not
g48810 not n5718 ; n5718_not
g48811 not n9507 ; n9507_not
g48812 not n4836 ; n4836_not
g48813 not n7941 ; n7941_not
g48814 not n2847 ; n2847_not
g48815 not n7581 ; n7581_not
g48816 not n9435 ; n9435_not
g48817 not n7932 ; n7932_not
g48818 not n7644 ; n7644_not
g48819 not n5961 ; n5961_not
g48820 not n6096 ; n6096_not
g48821 not n4089 ; n4089_not
g48822 not n7572 ; n7572_not
g48823 not n5934 ; n5934_not
g48824 not n5943 ; n5943_not
g48825 not n4098 ; n4098_not
g48826 not n3459 ; n3459_not
g48827 not n7455 ; n7455_not
g48828 not n9453 ; n9453_not
g48829 not n5952 ; n5952_not
g48830 not n6078 ; n6078_not
g48831 not n5907 ; n5907_not
g48832 not n9732 ; n9732_not
g48833 not n6159 ; n6159_not
g48834 not n4818 ; n4818_not
g48835 not n9741 ; n9741_not
g48836 not n9255 ; n9255_not
g48837 not n3387 ; n3387_not
g48838 not n4377 ; n4377_not
g48839 not n9534 ; n9534_not
g48840 not n7617 ; n7617_not
g48841 not n3990 ; n3990_not
g48842 not n9354 ; n9354_not
g48843 not n7383 ; n7383_not
g48844 not n7464 ; n7464_not
g48845 not n9444 ; n9444_not
g48846 not n9606 ; n9606_not
g48847 not n5673 ; n5673_not
g48848 not n7806 ; n7806_not
g48849 not n4962 ; n4962_not
g48850 not n9516 ; n9516_not
g48851 not n4278 ; n4278_not
g48852 not n8535 ; n8535_not
g48853 not n5277 ; n5277_not
g48854 not n6546 ; n6546_not
g48855 not n4458 ; n4458_not
g48856 not n3666 ; n3666_not
g48857 not n6519 ; n6519_not
g48858 not n8751 ; n8751_not
g48859 not n7059 ; n7059_not
g48860 not n2946 ; n2946_not
g48861 not n3846 ; n3846_not
g48862 not n7068 ; n7068_not
g48863 not n3648 ; n3648_not
g48864 not n8337 ; n8337_not
g48865 not n6681 ; n6681_not
g48866 not n9048 ; n9048_not
g48867 not n7086 ; n7086_not
g48868 not n6492 ; n6492_not
g48869 not n7095 ; n7095_not
g48870 not n8553 ; n8553_not
g48871 not n8706 ; n8706_not
g48872 not n6456 ; n6456_not
g48873 not n6465 ; n6465_not
g48874 not n7815 ; n7815_not
g48875 not n7554 ; n7554_not
g48876 not n7509 ; n7509_not
g48877 not n2667 ; n2667_not
g48878 not n8490 ; n8490_not
g48879 not n6582 ; n6582_not
g48880 not n8823 ; n8823_not
g48881 not n6924 ; n6924_not
g48882 not n6618 ; n6618_not
g48883 not n4557 ; n4557_not
g48884 not n8850 ; n8850_not
g48885 not n8463 ; n8463_not
g48886 not n9705 ; n9705_not
g48887 not n8841 ; n8841_not
g48888 not n4647 ; n4647_not
g48889 not n6915 ; n6915_not
g48890 not n8436 ; n8436_not
g48891 not n8805 ; n8805_not
g48892 not n8427 ; n8427_not
g48893 not n6663 ; n6663_not
g48894 not n8418 ; n8418_not
g48895 not n4395 ; n4395_not
g48896 not n8409 ; n8409_not
g48897 not n6573 ; n6573_not
g48898 not n3099 ; n3099_not
g48899 not n5484 ; n5484_not
g48900 not n5493 ; n5493_not
g48901 not n6933 ; n6933_not
g48902 not n6564 ; n6564_not
g48903 not n8391 ; n8391_not
g48904 not n8382 ; n8382_not
g48905 not n4665 ; n4665_not
g48906 not n7185 ; n7185_not
g48907 not n9138 ; n9138_not
g48908 not n8661 ; n8661_not
g48909 not n2892 ; n2892_not
g48910 not n4584 ; n4584_not
g48911 not n9156 ; n9156_not
g48912 not n9165 ; n9165_not
g48913 not n3558 ; n3558_not
g48914 not n8652 ; n8652_not
g48915 not n5358 ; n5358_not
g48916 not n3576 ; n3576_not
g48917 not n3891 ; n3891_not
g48918 not n6483 ; n6483_not
g48919 not n5178 ; n5178_not
g48920 not n3567 ; n3567_not
g48921 not n5637 ; n5637_not
g48922 not n6807 ; n6807_not
g48923 not n7248 ; n7248_not
g48924 not n3927 ; n3927_not
g48925 not n2577 ; n2577_not
g48926 not n5655 ; n5655_not
g48927 not n2874 ; n2874_not
g48928 not n6258 ; n6258_not
g48929 not n3747 ; n3747_not
g48930 not n9282 ; n9282_not
g48931 not n5376 ; n5376_not
g48932 not n4773 ; n4773_not
g48933 not n8175 ; n8175_not
g48934 not n3855 ; n3855_not
g48935 not n4719 ; n4719_not
g48936 not n4539 ; n4539_not
g48937 not n6447 ; n6447_not
g48938 not n4485 ; n4485_not
g48939 not n8571 ; n8571_not
g48940 not n5565 ; n5565_not
g48941 not n5574 ; n5574_not
g48942 not n6825 ; n6825_not
g48943 not n6735 ; n6735_not
g48944 not n2766 ; n2766_not
g48945 not n4728 ; n4728_not
g48946 not n4737 ; n4737_not
g48947 not n3882 ; n3882_not
g48948 not n7167 ; n7167_not
g48949 not n8590 ; n8590_not
g48950 not n6169 ; n6169_not
g48951 not n8806 ; n8806_not
g48952 not n9535 ; n9535_not
g48953 not n8473 ; n8473_not
g48954 not n8554 ; n8554_not
g48955 not n8815 ; n8815_not
g48956 not n9616 ; n9616_not
g48957 not n8572 ; n8572_not
g48958 not n8635 ; n8635_not
g48959 not n9490 ; n9490_not
g48960 not n7429 ; n7429_not
g48961 not n9526 ; n9526_not
g48962 not n2695 ; n2695_not
g48963 not n2983 ; n2983_not
g48964 not n8626 ; n8626_not
g48965 not n8752 ; n8752_not
g48966 not n8761 ; n8761_not
g48967 not n9715 ; n9715_not
g48968 not n9508 ; n9508_not
g48969 not n8545 ; n8545_not
g48970 not n7753 ; n7753_not
g48971 not n7645 ; n7645_not
g48972 not n8608 ; n8608_not
g48973 not n8518 ; n8518_not
g48974 not n7825 ; n7825_not
g48975 not n8770 ; n8770_not
g48976 not n7834 ; n7834_not
g48977 not n9652 ; n9652_not
g48978 not n2677 ; n2677_not
g48979 not n8671 ; n8671_not
g48980 not n8617 ; n8617_not
g48981 not n7780 ; n7780_not
g48982 not n2893 ; n2893_not
g48983 not n2758 ; n2758_not
g48984 not n2749 ; n2749_not
g48985 not n2857 ; n2857_not
g48986 not n9391 ; n9391_not
g48987 not n8266 ; n8266_not
g48988 not n9319 ; n9319_not
g48989 not n8194 ; n8194_not
g48990 not n8185 ; n8185_not
g48991 not n9931 ; n9931_not
g48992 not n9445 ; n9445_not
g48993 not n7636 ; n7636_not
g48994 not n8167 ; n8167_not
g48995 not n9328 ; n9328_not
g48996 not n6277 ; n6277_not
g48997 not n8158 ; n8158_not
g48998 not n8239 ; n8239_not
g48999 not n2767 ; n2767_not
g49000 not n2488 ; n2488_not
g49001 not n2875 ; n2875_not
g49002 not n8257 ; n8257_not
g49003 not n2587 ; n2587_not
g49004 not n3199 ; n3199_not
g49005 not n9265 ; n9265_not
g49006 not n9274 ; n9274_not
g49007 not n8275 ; n8275_not
g49008 not n9283 ; n9283_not
g49009 not n9148 ; n9148_not
g49010 not n2866 ; n2866_not
g49011 not n7474 ; n7474_not
g49012 not n9346 ; n9346_not
g49013 not n8419 ; n8419_not
g49014 not n8932 ; n8932_not
g49015 not n8428 ; n8428_not
g49016 not n8446 ; n8446_not
g49017 not n8860 ; n8860_not
g49018 not n8455 ; n8455_not
g49019 not n9436 ; n9436_not
g49020 not n3298 ; n3298_not
g49021 not n7465 ; n7465_not
g49022 not n7726 ; n7726_not
g49023 not n8833 ; n8833_not
g49024 not n8482 ; n8482_not
g49025 not n9067 ; n9067_not
g49026 not n9049 ; n9049_not
g49027 not n9913 ; n9913_not
g49028 not n9904 ; n9904_not
g49029 not n8149 ; n8149_not
g49030 not n8347 ; n8347_not
g49031 not n8356 ; n8356_not
g49032 not n2839 ; n2839_not
g49033 not n9733 ; n9733_not
g49034 not n9832 ; n9832_not
g49035 not n2965 ; n2965_not
g49036 not n9805 ; n9805_not
g49037 not n7357 ; n7357_not
g49038 not n4639 ; n4639_not
g49039 not n6790 ; n6790_not
g49040 not n5953 ; n5953_not
g49041 not n3739 ; n3739_not
g49042 not n6709 ; n6709_not
g49043 not n7555 ; n7555_not
g49044 not n5296 ; n5296_not
g49045 not n6817 ; n6817_not
g49046 not n6853 ; n6853_not
g49047 not n7528 ; n7528_not
g49048 not n5926 ; n5926_not
g49049 not n5377 ; n5377_not
g49050 not n3487 ; n3487_not
g49051 not n5917 ; n5917_not
g49052 not n6871 ; n6871_not
g49053 not n5782 ; n5782_not
g49054 not n6880 ; n6880_not
g49055 not n4585 ; n4585_not
g49056 not n3793 ; n3793_not
g49057 not n5089 ; n5089_not
g49058 not n6691 ; n6691_not
g49059 not n6088 ; n6088_not
g49060 not n4189 ; n4189_not
g49061 not n4756 ; n4756_not
g49062 not n3748 ; n3748_not
g49063 not n5197 ; n5197_not
g49064 not n6754 ; n6754_not
g49065 not n4693 ; n4693_not
g49066 not n4657 ; n4657_not
g49067 not n5269 ; n5269_not
g49068 not n6718 ; n6718_not
g49069 not n4666 ; n4666_not
g49070 not n5971 ; n5971_not
g49071 not n6772 ; n6772_not
g49072 not n7573 ; n7573_not
g49073 not n5593 ; n5593_not
g49074 not n7384 ; n7384_not
g49075 not n7375 ; n7375_not
g49076 not n7366 ; n7366_not
g49077 not n5629 ; n5629_not
g49078 not n5665 ; n5665_not
g49079 not n7285 ; n7285_not
g49080 not n7078 ; n7078_not
g49081 not n7267 ; n7267_not
g49082 not n5755 ; n5755_not
g49083 not n4369 ; n4369_not
g49084 not n5683 ; n5683_not
g49085 not n3559 ; n3559_not
g49086 not n3568 ; n3568_not
g49087 not n3595 ; n3595_not
g49088 not n7159 ; n7159_not
g49089 not n7168 ; n7168_not
g49090 not n5728 ; n5728_not
g49091 not n7195 ; n7195_not
g49092 not n4567 ; n4567_not
g49093 not n4558 ; n4558_not
g49094 not n4549 ; n4549_not
g49095 not n6907 ; n6907_not
g49096 not n7492 ; n7492_not
g49097 not n5890 ; n5890_not
g49098 not n5827 ; n5827_not
g49099 not n4468 ; n4468_not
g49100 not n6484 ; n6484_not
g49101 not n7447 ; n7447_not
g49102 not n6943 ; n6943_not
g49103 not n5872 ; n5872_not
g49104 not n4477 ; n4477_not
g49105 not n3478 ; n3478_not
g49106 not n5548 ; n5548_not
g49107 not n4297 ; n4297_not
g49108 not n6961 ; n6961_not
g49109 not n7393 ; n7393_not
g49110 not n5809 ; n5809_not
g49111 not n7654 ; n7654_not
g49112 not n4765 ; n4765_not
g49113 not n4972 ; n4972_not
g49114 not n3919 ; n3919_not
g49115 not n3775 ; n3775_not
g49116 not n6259 ; n6259_not
g49117 not n7609 ; n7609_not
g49118 not n7663 ; n7663_not
g49119 not n4954 ; n4954_not
g49120 not n6574 ; n6574_not
g49121 not n4909 ; n4909_not
g49122 not n3865 ; n3865_not
g49123 not n3379 ; n3379_not
g49124 not n4891 ; n4891_not
g49125 not n4990 ; n4990_not
g49126 not n6646 ; n6646_not
g49127 not n6466 ; n6466_not
g49128 not n6619 ; n6619_not
g49129 not n6628 ; n6628_not
g49130 not n6538 ; n6538_not
g49131 not n3838 ; n3838_not
g49132 not n6376 ; n6376_not
g49133 not n6394 ; n6394_not
g49134 not n6556 ; n6556_not
g49135 not n3883 ; n3883_not
g49136 not n6349 ; n6349_not
g49137 not n3892 ; n3892_not
g49138 not n7627 ; n7627_not
g49139 not n4792 ; n4792_not
g49140 not n4945 ; n4945_not
g49141 not n4981 ; n4981_not
g49142 not n6493 ; n6493_not
g49143 not n6367 ; n6367_not
g49144 not n4927 ; n4927_not
g49145 not n9608 ; n9608_not
g49146 not n6197 ; n6197_not
g49147 not n6926 ; n6926_not
g49148 not n6593 ; n6593_not
g49149 not n6764 ; n6764_not
g49150 not n6980 ; n6980_not
g49151 not n6962 ; n6962_not
g49152 not n9581 ; n9581_not
g49153 not n8951 ; n8951_not
g49154 not n3659 ; n3659_not
g49155 not n5882 ; n5882_not
g49156 not n6395 ; n6395_not
g49157 not n5855 ; n5855_not
g49158 not n9671 ; n9671_not
g49159 not n6953 ; n6953_not
g49160 not n9653 ; n9653_not
g49161 not n3866 ; n3866_not
g49162 not n2894 ; n2894_not
g49163 not n8933 ; n8933_not
g49164 not n8465 ; n8465_not
g49165 not n9644 ; n9644_not
g49166 not n8906 ; n8906_not
g49167 not n8474 ; n8474_not
g49168 not n3668 ; n3668_not
g49169 not n9851 ; n9851_not
g49170 not n8348 ; n8348_not
g49171 not n3848 ; n3848_not
g49172 not n7097 ; n7097_not
g49173 not n5747 ; n5747_not
g49174 not n3596 ; n3596_not
g49175 not n5585 ; n5585_not
g49176 not n9914 ; n9914_not
g49177 not n6494 ; n6494_not
g49178 not n2939 ; n2939_not
g49179 not n2966 ; n2966_not
g49180 not n7178 ; n7178_not
g49181 not n6566 ; n6566_not
g49182 not n5369 ; n5369_not
g49183 not n9932 ; n9932_not
g49184 not n8285 ; n8285_not
g49185 not n6458 ; n6458_not
g49186 not n6467 ; n6467_not
g49187 not n3488 ; n3488_not
g49188 not n9761 ; n9761_not
g49189 not n7628 ; n7628_not
g49190 not n9770 ; n9770_not
g49191 not n3695 ; n3695_not
g49192 not n5792 ; n5792_not
g49193 not n9815 ; n9815_not
g49194 not n9824 ; n9824_not
g49195 not n5774 ; n5774_not
g49196 not n8366 ; n8366_not
g49197 not n3677 ; n3677_not
g49198 not n7862 ; n7862_not
g49199 not n6476 ; n6476_not
g49200 not n9842 ; n9842_not
g49201 not n6665 ; n6665_not
g49202 not n3497 ; n3497_not
g49203 not n9284 ; n9284_not
g49204 not n8672 ; n8672_not
g49205 not n5981 ; n5981_not
g49206 not n5990 ; n5990_not
g49207 not n9419 ; n9419_not
g49208 not n9428 ; n9428_not
g49209 not n8780 ; n8780_not
g49210 not n8654 ; n8654_not
g49211 not n7475 ; n7475_not
g49212 not n9437 ; n9437_not
g49213 not n2867 ; n2867_not
g49214 not n8645 ; n8645_not
g49215 not n7961 ; n7961_not
g49216 not n3965 ; n3965_not
g49217 not n8636 ; n8636_not
g49218 not n8753 ; n8753_not
g49219 not n3992 ; n3992_not
g49220 not n6683 ; n6683_not
g49221 not n3983 ; n3983_not
g49222 not n9248 ; n9248_not
g49223 not n2849 ; n2849_not
g49224 not n8708 ; n8708_not
g49225 not n9257 ; n9257_not
g49226 not n8717 ; n8717_not
g49227 not n9356 ; n9356_not
g49228 not n4199 ; n4199_not
g49229 not n6728 ; n6728_not
g49230 not n9365 ; n9365_not
g49231 not n8690 ; n8690_not
g49232 not n6746 ; n6746_not
g49233 not n9527 ; n9527_not
g49234 not n5918 ; n5918_not
g49235 not n6359 ; n6359_not
g49236 not n9185 ; n9185_not
g49237 not n2885 ; n2885_not
g49238 not n7592 ; n7592_not
g49239 not n9158 ; n9158_not
g49240 not n8393 ; n8393_not
g49241 not n4289 ; n4289_not
g49242 not n9545 ; n9545_not
g49243 not n9554 ; n9554_not
g49244 not n9563 ; n9563_not
g49245 not n6890 ; n6890_not
g49246 not n8528 ; n8528_not
g49247 not n8870 ; n8870_not
g49248 not n6917 ; n6917_not
g49249 not n6647 ; n6647_not
g49250 not n3956 ; n3956_not
g49251 not n3938 ; n3938_not
g49252 not n9446 ; n9446_not
g49253 not n5963 ; n5963_not
g49254 not n5954 ; n5954_not
g49255 not n6809 ; n6809_not
g49256 not n3929 ; n3929_not
g49257 not n8609 ; n8609_not
g49258 not n5945 ; n5945_not
g49259 not n2777 ; n2777_not
g49260 not n5936 ; n5936_not
g49261 not n6827 ; n6827_not
g49262 not n8573 ; n8573_not
g49263 not n5927 ; n5927_not
g49264 not n7547 ; n7547_not
g49265 not n2678 ; n2678_not
g49266 not n7565 ; n7565_not
g49267 not n4649 ; n4649_not
g49268 not n4658 ; n4658_not
g49269 not n5279 ; n5279_not
g49270 not n4676 ; n4676_not
g49271 not n7970 ; n7970_not
g49272 not n7493 ; n7493_not
g49273 not n2759 ; n2759_not
g49274 not n7457 ; n7457_not
g49275 not n4487 ; n4487_not
g49276 not n4496 ; n4496_not
g49277 not n5495 ; n5495_not
g49278 not n5486 ; n5486_not
g49279 not n5468 ; n5468_not
g49280 not n5459 ; n5459_not
g49281 not n6485 ; n6485_not
g49282 not n4568 ; n4568_not
g49283 not n4577 ; n4577_not
g49284 not n2687 ; n2687_not
g49285 not n3389 ; n3389_not
g49286 not n8249 ; n8249_not
g49287 not n4991 ; n4991_not
g49288 not n7637 ; n7637_not
g49289 not n7772 ; n7772_not
g49290 not n7763 ; n7763_not
g49291 not n4955 ; n4955_not
g49292 not n4919 ; n4919_not
g49293 not n4937 ; n4937_not
g49294 not n4694 ; n4694_not
g49295 not n4685 ; n4685_not
g49296 not n4748 ; n4748_not
g49297 not n5189 ; n5189_not
g49298 not n7583 ; n7583_not
g49299 not n4766 ; n4766_not
g49300 not n7619 ; n7619_not
g49301 not n5099 ; n5099_not
g49302 not n9338 ; n9338_not
g49303 not n4838 ; n4838_not
g49304 not n7871 ; n7871_not
g49305 not n3398 ; n3398_not
g49306 not n7673 ; n7673_not
g49307 not n5648 ; n5648_not
g49308 not n2489 ; n2489_not
g49309 not n9950 ; n9950_not
g49310 not n7358 ; n7358_not
g49311 not n8177 ; n8177_not
g49312 not n7259 ; n7259_not
g49313 not n7277 ; n7277_not
g49314 not n9626 ; n9626_not
g49315 not n5576 ; n5576_not
g49316 not n8186 ; n8186_not
g49317 not n4397 ; n4397_not
g49318 not n4379 ; n4379_not
g49319 not n9941 ; n9941_not
g49320 not n8168 ; n8168_not
g49321 not n5657 ; n5657_not
g49322 not n7295 ; n7295_not
g49323 not n8267 ; n8267_not
g49324 not n8736 ; n8736_not
g49325 not n6198 ; n6198_not
g49326 not n9249 ; n9249_not
g49327 not n9339 ; n9339_not
g49328 not n3948 ; n3948_not
g49329 not n2976 ; n2976_not
g49330 not n3678 ; n3678_not
g49331 not n3975 ; n3975_not
g49332 not n6675 ; n6675_not
g49333 not n3993 ; n3993_not
g49334 not n7269 ; n7269_not
g49335 not n7926 ; n7926_not
g49336 not n6756 ; n6756_not
g49337 not n8754 ; n8754_not
g49338 not n7089 ; n7089_not
g49339 not n3984 ; n3984_not
g49340 not n9294 ; n9294_not
g49341 not n8772 ; n8772_not
g49342 not n4758 ; n4758_not
g49343 not n4767 ; n4767_not
g49344 not n5667 ; n5667_not
g49345 not n7944 ; n7944_not
g49346 not n7953 ; n7953_not
g49347 not n9393 ; n9393_not
g49348 not n9366 ; n9366_not
g49349 not n9375 ; n9375_not
g49350 not n3759 ; n3759_not
g49351 not n8682 ; n8682_not
g49352 not n5199 ; n5199_not
g49353 not n8718 ; n8718_not
g49354 not n7287 ; n7287_not
g49355 not n4776 ; n4776_not
g49356 not n8727 ; n8727_not
g49357 not n4785 ; n4785_not
g49358 not n6747 ; n6747_not
g49359 not n8169 ; n8169_not
g49360 not n9168 ; n9168_not
g49361 not n4983 ; n4983_not
g49362 not n6387 ; n6387_not
g49363 not n8907 ; n8907_not
g49364 not n2895 ; n2895_not
g49365 not n8934 ; n8934_not
g49366 not n9645 ; n9645_not
g49367 not n3867 ; n3867_not
g49368 not n4974 ; n4974_not
g49369 not n6459 ; n6459_not
g49370 not n7746 ; n7746_not
g49371 not n8268 ; n8268_not
g49372 not n6576 ; n6576_not
g49373 not n4398 ; n4398_not
g49374 not n4947 ; n4947_not
g49375 not n9924 ; n9924_not
g49376 not n6495 ; n6495_not
g49377 not n4938 ; n4938_not
g49378 not n9942 ; n9942_not
g49379 not n2949 ; n2949_not
g49380 not n7692 ; n7692_not
g49381 not n7197 ; n7197_not
g49382 not n6558 ; n6558_not
g49383 not n4848 ; n4848_not
g49384 not n9285 ; n9285_not
g49385 not n5685 ; n5685_not
g49386 not n4857 ; n4857_not
g49387 not n8790 ; n8790_not
g49388 not n3957 ; n3957_not
g49389 not n6657 ; n6657_not
g49390 not n5757 ; n5757_not
g49391 not n4884 ; n4884_not
g49392 not n6639 ; n6639_not
g49393 not n3777 ; n3777_not
g49394 not n7791 ; n7791_not
g49395 not n8817 ; n8817_not
g49396 not n2868 ; n2868_not
g49397 not n4893 ; n4893_not
g49398 not n6297 ; n6297_not
g49399 not n8835 ; n8835_not
g49400 not n3885 ; n3885_not
g49401 not n4866 ; n4866_not
g49402 not n3489 ; n3489_not
g49403 not n3768 ; n3768_not
g49404 not n2886 ; n2886_not
g49405 not n8547 ; n8547_not
g49406 not n6369 ; n6369_not
g49407 not n9573 ; n9573_not
g49408 not n4578 ; n4578_not
g49409 not n8178 ; n8178_not
g49410 not n8088 ; n8088_not
g49411 not n8079 ; n8079_not
g49412 not n5397 ; n5397_not
g49413 not n6990 ; n6990_not
g49414 not n6945 ; n6945_not
g49415 not n5919 ; n5919_not
g49416 not n8556 ; n8556_not
g49417 not n2679 ; n2679_not
g49418 not n8565 ; n8565_not
g49419 not n9762 ; n9762_not
g49420 not n8196 ; n8196_not
g49421 not n7548 ; n7548_not
g49422 not n4596 ; n4596_not
g49423 not n6828 ; n6828_not
g49424 not n6819 ; n6819_not
g49425 not n7494 ; n7494_not
g49426 not n5865 ; n5865_not
g49427 not n9717 ; n9717_not
g49428 not n8448 ; n8448_not
g49429 not n5586 ; n5586_not
g49430 not n5568 ; n5568_not
g49431 not n9726 ; n9726_not
g49432 not n6963 ; n6963_not
g49433 not n9636 ; n9636_not
g49434 not n8475 ; n8475_not
g49435 not n5595 ; n5595_not
g49436 not n4299 ; n4299_not
g49437 not n9627 ; n9627_not
g49438 not n9618 ; n9618_not
g49439 not n5784 ; n5784_not
g49440 not n7395 ; n7395_not
g49441 not n6936 ; n6936_not
g49442 not n7476 ; n7476_not
g49443 not n6837 ; n6837_not
g49444 not n6909 ; n6909_not
g49445 not n6972 ; n6972_not
g49446 not n5955 ; n5955_not
g49447 not n8628 ; n8628_not
g49448 not n5793 ; n5793_not
g49449 not n2859 ; n2859_not
g49450 not n7575 ; n7575_not
g49451 not n5973 ; n5973_not
g49452 not n4677 ; n4677_not
g49453 not n8619 ; n8619_not
g49454 not n5775 ; n5775_not
g49455 not n8376 ; n8376_not
g49456 not n5649 ; n5649_not
g49457 not n9474 ; n9474_not
g49458 not n8655 ; n8655_not
g49459 not n9834 ; n9834_not
g49460 not n9492 ; n9492_not
g49461 not n8592 ; n8592_not
g49462 not n9357 ; n9357_not
g49463 not n2778 ; n2778_not
g49464 not n4695 ; n4695_not
g49465 not n3859 ; n3859_not
g49466 not n5569 ; n5569_not
g49467 not n3769 ; n3769_not
g49468 not n9835 ; n9835_not
g49469 not n9916 ; n9916_not
g49470 not n9376 ; n9376_not
g49471 not n6478 ; n6478_not
g49472 not n9709 ; n9709_not
g49473 not n5965 ; n5965_not
g49474 not n5857 ; n5857_not
g49475 not n5839 ; n5839_not
g49476 not n9574 ; n9574_not
g49477 not n6496 ; n6496_not
g49478 not n4849 ; n4849_not
g49479 not n9367 ; n9367_not
g49480 not n5983 ; n5983_not
g49481 not n5587 ; n5587_not
g49482 not n5659 ; n5659_not
g49483 not n9727 ; n9727_not
g49484 not n9466 ; n9466_not
g49485 not n4939 ; n4939_not
g49486 not n9637 ; n9637_not
g49487 not n9385 ; n9385_not
g49488 not n8962 ; n8962_not
g49489 not n9295 ; n9295_not
g49490 not n4966 ; n4966_not
g49491 not n9439 ; n9439_not
g49492 not n5884 ; n5884_not
g49493 not n4498 ; n4498_not
g49494 not n9349 ; n9349_not
g49495 not n5686 ; n5686_not
g49496 not n9259 ; n9259_not
g49497 not n2896 ; n2896_not
g49498 not n4885 ; n4885_not
g49499 not n5389 ; n5389_not
g49500 not n4876 ; n4876_not
g49501 not n4768 ; n4768_not
g49502 not n5794 ; n5794_not
g49503 not n4867 ; n4867_not
g49504 not n4858 ; n4858_not
g49505 not n5299 ; n5299_not
g49506 not n4795 ; n4795_not
g49507 not n9286 ; n9286_not
g49508 not n4993 ; n4993_not
g49509 not n3976 ; n3976_not
g49510 not n9475 ; n9475_not
g49511 not n4786 ; n4786_not
g49512 not n9871 ; n9871_not
g49513 not n9862 ; n9862_not
g49514 not n6379 ; n6379_not
g49515 not n5938 ; n5938_not
g49516 not n9178 ; n9178_not
g49517 not n9844 ; n9844_not
g49518 not n5767 ; n5767_not
g49519 not n3499 ; n3499_not
g49520 not n9565 ; n9565_not
g49521 not n9547 ; n9547_not
g49522 not n4399 ; n4399_not
g49523 not n4579 ; n4579_not
g49524 not n2878 ; n2878_not
g49525 not n5947 ; n5947_not
g49526 not n6298 ; n6298_not
g49527 not n9907 ; n9907_not
g49528 not n4894 ; n4894_not
g49529 not n5749 ; n5749_not
g49530 not n9754 ; n9754_not
g49531 not n5785 ; n5785_not
g49532 not n7369 ; n7369_not
g49533 not n4777 ; n4777_not
g49534 not n5596 ; n5596_not
g49535 not n7099 ; n7099_not
g49536 not n8773 ; n8773_not
g49537 not n3598 ; n3598_not
g49538 not n6658 ; n6658_not
g49539 not n8287 ; n8287_not
g49540 not n7189 ; n7189_not
g49541 not n7297 ; n7297_not
g49542 not n8827 ; n8827_not
g49543 not n3778 ; n3778_not
g49544 not n8845 ; n8845_not
g49545 not n7468 ; n7468_not
g49546 not n7486 ; n7486_not
g49547 not n8089 ; n8089_not
g49548 not n7549 ; n7549_not
g49549 not n7567 ; n7567_not
g49550 not n7963 ; n7963_not
g49551 not n7954 ; n7954_not
g49552 not n6586 ; n6586_not
g49553 not n7585 ; n7585_not
g49554 not n7873 ; n7873_not
g49555 not n6928 ; n6928_not
g49556 not n8494 ; n8494_not
g49557 not n8539 ; n8539_not
g49558 not n6865 ; n6865_not
g49559 not n8566 ; n8566_not
g49560 not n6847 ; n6847_not
g49561 not n8575 ; n8575_not
g49562 not n8548 ; n8548_not
g49563 not n6937 ; n6937_not
g49564 not n6766 ; n6766_not
g49565 not n8629 ; n8629_not
g49566 not n8647 ; n8647_not
g49567 not n6955 ; n6955_not
g49568 not n8665 ; n8665_not
g49569 not n8395 ; n8395_not
g49570 not n6982 ; n6982_not
g49571 not n3697 ; n3697_not
g49572 not n3688 ; n3688_not
g49573 not n6685 ; n6685_not
g49574 not n3589 ; n3589_not
g49575 not n7846 ; n7846_not
g49576 not n7495 ; n7495_not
g49577 not n7639 ; n7639_not
g49578 not n7819 ; n7819_not
g49579 not n7693 ; n7693_not
g49580 not n6568 ; n6568_not
g49581 not n7648 ; n7648_not
g49582 not n7855 ; n7855_not
g49583 not n7199 ; n7199_not
g49584 not n3968 ; n3968_not
g49585 not n9458 ; n9458_not
g49586 not n6398 ; n6398_not
g49587 not n8783 ; n8783_not
g49588 not n5849 ; n5849_not
g49589 not n4994 ; n4994_not
g49590 not n5993 ; n5993_not
g49591 not n3599 ; n3599_not
g49592 not n2969 ; n2969_not
g49593 not n9908 ; n9908_not
g49594 not n9296 ; n9296_not
g49595 not n8819 ; n8819_not
g49596 not n7757 ; n7757_not
g49597 not n5669 ; n5669_not
g49598 not n7289 ; n7289_not
g49599 not n8468 ; n8468_not
g49600 not n4976 ; n4976_not
g49601 not n7775 ; n7775_not
g49602 not n8981 ; n8981_not
g49603 not n9971 ; n9971_not
g49604 not n5975 ; n5975_not
g49605 not n5687 ; n5687_not
g49606 not n6884 ; n6884_not
g49607 not n9953 ; n9953_not
g49608 not n8648 ; n8648_not
g49609 not n8657 ; n8657_not
g49610 not n9719 ; n9719_not
g49611 not n8792 ; n8792_not
g49612 not n9368 ; n9368_not
g49613 not n2987 ; n2987_not
g49614 not n9764 ; n9764_not
g49615 not n6695 ; n6695_not
g49616 not n9638 ; n9638_not
g49617 not n9359 ; n9359_not
g49618 not n9773 ; n9773_not
g49619 not n5795 ; n5795_not
g49620 not n8693 ; n8693_not
g49621 not n9746 ; n9746_not
g49622 not n6488 ; n6488_not
g49623 not n9386 ; n9386_not
g49624 not n9818 ; n9818_not
g49625 not n9539 ; n9539_not
g49626 not n6677 ; n6677_not
g49627 not n8378 ; n8378_not
g49628 not n7928 ; n7928_not
g49629 not n5876 ; n5876_not
g49630 not n8747 ; n8747_not
g49631 not n6497 ; n6497_not
g49632 not n6749 ; n6749_not
g49633 not n8756 ; n8756_not
g49634 not n9845 ; n9845_not
g49635 not n5759 ; n5759_not
g49636 not n9872 ; n9872_not
g49637 not n9863 ; n9863_not
g49638 not n9485 ; n9485_not
g49639 not n6965 ; n6965_not
g49640 not n6956 ; n6956_not
g49641 not n5957 ; n5957_not
g49642 not n5399 ; n5399_not
g49643 not n4589 ; n4589_not
g49644 not n9593 ; n9593_not
g49645 not n7766 ; n7766_not
g49646 not n4598 ; n4598_not
g49647 not n4877 ; n4877_not
g49648 not n6794 ; n6794_not
g49649 not n9683 ; n9683_not
g49650 not n7577 ; n7577_not
g49651 not n5867 ; n5867_not
g49652 not n6389 ; n6389_not
g49653 not n4697 ; n4697_not
g49654 not n7496 ; n7496_not
g49655 not n4769 ; n4769_not
g49656 not n6938 ; n6938_not
g49657 not n8954 ; n8954_not
g49658 not n9575 ; n9575_not
g49659 not n5894 ; n5894_not
g49660 not n6857 ; n6857_not
g49661 not n4796 ; n4796_not
g49662 not n6866 ; n6866_not
g49663 not n7865 ; n7865_not
g49664 not n7874 ; n7874_not
g49665 not n6587 ; n6587_not
g49666 not n8459 ; n8459_not
g49667 not n9584 ; n9584_not
g49668 not n6785 ; n6785_not
g49669 not n3779 ; n3779_not
g49670 not n8198 ; n8198_not
g49671 not n8189 ; n8189_not
g49672 not n5597 ; n5597_not
g49673 not n7676 ; n7676_not
g49674 not n2699 ; n2699_not
g49675 not n7397 ; n7397_not
g49676 not n9197 ; n9197_not
g49677 not n5579 ; n5579_not
g49678 not n9188 ; n9188_not
g49679 not n7487 ; n7487_not
g49680 not n5498 ; n5498_not
g49681 not n8972 ; n8972_not
g49682 not n6578 ; n6578_not
g49683 not n3788 ; n3788_not
g49684 not n3699 ; n3699_not
g49685 not n4959 ; n4959_not
g49686 not n6975 ; n6975_not
g49687 not n6489 ; n6489_not
g49688 not n6867 ; n6867_not
g49689 not n2997 ; n2997_not
g49690 not n5985 ; n5985_not
g49691 not n8658 ; n8658_not
g49692 not n8991 ; n8991_not
g49693 not n5859 ; n5859_not
g49694 not n8982 ; n8982_not
g49695 not n6876 ; n6876_not
g49696 not n9657 ; n9657_not
g49697 not n8694 ; n8694_not
g49698 not n6777 ; n6777_not
g49699 not n8469 ; n8469_not
g49700 not n2988 ; n2988_not
g49701 not n4968 ; n4968_not
g49702 not n8667 ; n8667_not
g49703 not n9729 ; n9729_not
g49704 not n5967 ; n5967_not
g49705 not n5868 ; n5868_not
g49706 not n9486 ; n9486_not
g49707 not n9738 ; n9738_not
g49708 not n8586 ; n8586_not
g49709 not n5994 ; n5994_not
g49710 not n9189 ; n9189_not
g49711 not n9495 ; n9495_not
g49712 not n8577 ; n8577_not
g49713 not n9639 ; n9639_not
g49714 not n9972 ; n9972_not
g49715 not n6849 ; n6849_not
g49716 not n5886 ; n5886_not
g49717 not n9990 ; n9990_not
g49718 not n9747 ; n9747_not
g49719 not n8829 ; n8829_not
g49720 not n7389 ; n7389_not
g49721 not n9594 ; n9594_not
g49722 not n8964 ; n8964_not
g49723 not n8892 ; n8892_not
g49724 not n3879 ; n3879_not
g49725 not n7569 ; n7569_not
g49726 not n7974 ; n7974_not
g49727 not n7956 ; n7956_not
g49728 not n7938 ; n7938_not
g49729 not n7596 ; n7596_not
g49730 not n9099 ; n9099_not
g49731 not n8937 ; n8937_not
g49732 not n4869 ; n4869_not
g49733 not n8946 ; n8946_not
g49734 not n6597 ; n6597_not
g49735 not n4788 ; n4788_not
g49736 not n9576 ; n9576_not
g49737 not n6993 ; n6993_not
g49738 not n9774 ; n9774_not
g49739 not n9783 ; n9783_not
g49740 not n6894 ; n6894_not
g49741 not n6687 ; n6687_not
g49742 not n8388 ; n8388_not
g49743 not n3978 ; n3978_not
g49744 not n9828 ; n9828_not
g49745 not n5778 ; n5778_not
g49746 not n9567 ; n9567_not
g49747 not n8757 ; n8757_not
g49748 not n9882 ; n9882_not
g49749 not n2799 ; n2799_not
g49750 not n7785 ; n7785_not
g49751 not n9936 ; n9936_not
g49752 not n9945 ; n9945_not
g49753 not n7695 ; n7695_not
g49754 not n4995 ; n4995_not
g49755 not n9927 ; n9927_not
g49756 not n8298 ; n8298_not
g49757 not n9918 ; n9918_not
g49758 not n8775 ; n8775_not
g49759 not n6669 ; n6669_not
g49760 not n8478 ; n8478_not
g49761 not n9649 ; n9649_not
g49762 not n7696 ; n7696_not
g49763 not n5797 ; n5797_not
g49764 not n5878 ; n5878_not
g49765 not n8488 ; n8488_not
g49766 not n5896 ; n5896_not
g49767 not n6949 ; n6949_not
g49768 not n9694 ; n9694_not
g49769 not n4987 ; n4987_not
g49770 not n9937 ; n9937_not
g49771 not n9946 ; n9946_not
g49772 not n9964 ; n9964_not
g49773 not n9982 ; n9982_not
g49774 not n9991 ; n9991_not
g49775 not n5599 ; n5599_not
g49776 not n7399 ; n7399_not
g49777 not n7498 ; n7498_not
g49778 not n9739 ; n9739_not
g49779 not n7588 ; n7588_not
g49780 not n4789 ; n4789_not
g49781 not n4798 ; n4798_not
g49782 not n7894 ; n7894_not
g49783 not n7867 ; n7867_not
g49784 not n5869 ; n5869_not
g49785 not n9658 ; n9658_not
g49786 not n7669 ; n7669_not
g49787 not n9667 ; n9667_not
g49788 not n9289 ; n9289_not
g49789 not n9676 ; n9676_not
g49790 not n5779 ; n5779_not
g49791 not n6967 ; n6967_not
g49792 not n6976 ; n6976_not
g49793 not n4879 ; n4879_not
g49794 not n9775 ; n9775_not
g49795 not n4978 ; n4978_not
g49796 not n8389 ; n8389_not
g49797 not n5788 ; n5788_not
g49798 not n9856 ; n9856_not
g49799 not n5986 ; n5986_not
g49800 not n6589 ; n6589_not
g49801 not n8659 ; n8659_not
g49802 not n6859 ; n6859_not
g49803 not n3979 ; n3979_not
g49804 not n8749 ; n8749_not
g49805 not n6679 ; n6679_not
g49806 not n9397 ; n9397_not
g49807 not n8596 ; n8596_not
g49808 not n6697 ; n6697_not
g49809 not n6886 ; n6886_not
g49810 not n8677 ; n8677_not
g49811 not n8686 ; n8686_not
g49812 not n2899 ; n2899_not
g49813 not n2989 ; n2989_not
g49814 not n8695 ; n8695_not
g49815 not n8767 ; n8767_not
g49816 not n8497 ; n8497_not
g49817 not n9298 ; n9298_not
g49818 not n8866 ; n8866_not
g49819 not n8857 ; n8857_not
g49820 not n8839 ; n8839_not
g49821 not n8992 ; n8992_not
g49822 not n5969 ; n5969_not
g49823 not n8768 ; n8768_not
g49824 not n4988 ; n4988_not
g49825 not n8777 ; n8777_not
g49826 not n6779 ; n6779_not
g49827 not n9875 ; n9875_not
g49828 not n9848 ; n9848_not
g49829 not n9398 ; n9398_not
g49830 not n6689 ; n6689_not
g49831 not n8687 ; n8687_not
g49832 not n9749 ; n9749_not
g49833 not n6986 ; n6986_not
g49834 not n9758 ; n9758_not
g49835 not n9785 ; n9785_not
g49836 not n5798 ; n5798_not
g49837 not n8399 ; n8399_not
g49838 not n5897 ; n5897_not
g49839 not n8858 ; n8858_not
g49840 not n5888 ; n5888_not
g49841 not n7499 ; n7499_not
g49842 not n6599 ; n6599_not
g49843 not n7958 ; n7958_not
g49844 not n7688 ; n7688_not
g49845 not n7589 ; n7589_not
g49846 not n8957 ; n8957_not
g49847 not n6869 ; n6869_not
g49848 not n9992 ; n9992_not
g49849 not n7877 ; n7877_not
g49850 not n9659 ; n9659_not
g49851 not n9578 ; n9578_not
g49852 not n8786 ; n8786_not
g49853 not n8579 ; n8579_not
g49854 not n7598 ; n7598_not
g49855 not n8984 ; n8984_not
g49856 not n5699 ; n5699_not
g49857 not n9686 ; n9686_not
g49858 not n6788 ; n6788_not
g49859 not n9677 ; n9677_not
g49860 not n7986 ; n7986_not
g49861 not n9795 ; n9795_not
g49862 not n4998 ; n4998_not
g49863 not n8985 ; n8985_not
g49864 not n8868 ; n8868_not
g49865 not n7788 ; n7788_not
g49866 not n3999 ; n3999_not
g49867 not n6699 ; n6699_not
g49868 not n9777 ; n9777_not
g49869 not n5988 ; n5988_not
g49870 not n7977 ; n7977_not
g49871 not n5799 ; n5799_not
g49872 not n7968 ; n7968_not
g49873 not n8796 ; n8796_not
g49874 not n7779 ; n7779_not
g49875 not n7995 ; n7995_not
g49876 not n7878 ; n7878_not
g49877 not n7887 ; n7887_not
g49878 not n9957 ; n9957_not
g49879 not n9876 ; n9876_not
g49880 not n9984 ; n9984_not
g49881 not n4989 ; n4989_not
g49882 not n9948 ; n9948_not
g49883 not n8679 ; n8679_not
g49884 not n5898 ; n5898_not
g49885 not n9669 ; n9669_not
g49886 not n9687 ; n9687_not
g49887 not n8697 ; n8697_not
g49888 not n8598 ; n8598_not
g49889 not n6798 ; n6798_not
g49890 not n9696 ; n9696_not
g49891 not n6897 ; n6897_not
g49892 not n9498 ; n9498_not
g49893 not n9588 ; n9588_not
g49894 not n9597 ; n9597_not
g49895 not n9768 ; n9768_not
g49896 not n6879 ; n6879_not
g49897 not n8994 ; n8994_not
g49898 not n4999 ; n4999_not
g49899 not n5998 ; n5998_not
g49900 not n5989 ; n5989_not
g49901 not n8698 ; n8698_not
g49902 not n9949 ; n9949_not
g49903 not n9679 ; n9679_not
g49904 not n7897 ; n7897_not
g49905 not n8959 ; n8959_not
g49906 not n9598 ; n9598_not
g49907 not n9994 ; n9994_not
g49908 not n6997 ; n6997_not
g49909 not n5899 ; n5899_not
g49910 not n9958 ; n9958_not
g49911 not n9976 ; n9976_not
g49912 not n8995 ; n8995_not
g49913 not n9697 ; n9697_not
g49914 not n7996 ; n7996_not
g49915 not n7969 ; n7969_not
g49916 not n9967 ; n9967_not
g49917 not n9986 ; n9986_not
g49918 not n9896 ; n9896_not
g49919 not n8888 ; n8888_not
g49920 not n9878 ; n9878_not
g49921 not n9698 ; n9698_not
g49922 not n8996 ; n8996_not
g49923 not n9779 ; n9779_not
g49924 not n9968 ; n9968_not
g49925 not n9977 ; n9977_not
g49926 not n7898 ; n7898_not
g49927 not n5999 ; n5999_not
g49928 not n8889 ; n8889_not
g49929 not n9978 ; n9978_not
g49930 not n7989 ; n7989_not
g49931 not n6999 ; n6999_not
g49932 not n9996 ; n9996_not
g49933 not n9988 ; n9988_not
g49934 not n8989 ; n8989_not
g49935 not n9889 ; n9889_not
g49936 not n8899 ; n8899_not
g49937 not n9799 ; n9799_not
g49938 not n7999 ; n7999_not
g49939 not n8999 ; n8999_not
g49940 not n10000 ; n10000_not
g49941 not n10002 ; n10002_not
g49942 not n11100 ; n11100_not
g49943 not n20001 ; n20001_not
g49944 not n30000 ; n30000_not
g49945 not n20010 ; n20010_not
g49946 not n21010 ; n21010_not
g49947 not n10210 ; n10210_not
g49948 not n40000 ; n40000_not
g49949 not n21001 ; n21001_not
g49950 not n10111 ; n10111_not
g49951 not n20002 ; n20002_not
g49952 not n20020 ; n20020_not
g49953 not n21100 ; n21100_not
g49954 not n10003 ; n10003_not
g49955 not n10021 ; n10021_not
g49956 not n20101 ; n20101_not
g49957 not n10012 ; n10012_not
g49958 not n11011 ; n11011_not
g49959 not n30100 ; n30100_not
g49960 not n10004 ; n10004_not
g49961 not n20120 ; n20120_not
g49962 not n11120 ; n11120_not
g49963 not n10040 ; n10040_not
g49964 not n20030 ; n20030_not
g49965 not n21110 ; n21110_not
g49966 not n20012 ; n20012_not
g49967 not n32000 ; n32000_not
g49968 not n22001 ; n22001_not
g49969 not n10103 ; n10103_not
g49970 not n11201 ; n11201_not
g49971 not n40010 ; n40010_not
g49972 not n10121 ; n10121_not
g49973 not n12011 ; n12011_not
g49974 not n12101 ; n12101_not
g49975 not n30002 ; n30002_not
g49976 not n40100 ; n40100_not
g49977 not n30020 ; n30020_not
g49978 not n10202 ; n10202_not
g49979 not n10220 ; n10220_not
g49980 not n10310 ; n10310_not
g49981 not n20201 ; n20201_not
g49982 not n11210 ; n11210_not
g49983 not n20111 ; n20111_not
g49984 not n13001 ; n13001_not
g49985 not n30110 ; n30110_not
g49986 not n10400 ; n10400_not
g49987 not n23000 ; n23000_not
g49988 not n12021 ; n12021_not
g49989 not n42000 ; n42000_not
g49990 not n12111 ; n12111_not
g49991 not n20013 ; n20013_not
g49992 not n12102 ; n12102_not
g49993 not n22011 ; n22011_not
g49994 not n11211 ; n11211_not
g49995 not n11004 ; n11004_not
g49996 not n21021 ; n21021_not
g49997 not n10221 ; n10221_not
g49998 not n10410 ; n10410_not
g49999 not n20040 ; n20040_not
g50000 not n12201 ; n12201_not
g50001 not n40200 ; n40200_not
g50002 not n20130 ; n20130_not
g50003 not n21030 ; n21030_not
g50004 not n10203 ; n10203_not
g50005 not n15000 ; n15000_not
g50006 not n13011 ; n13011_not
g50007 not n20220 ; n20220_not
g50008 not n10131 ; n10131_not
g50009 not n20211 ; n20211_not
g50010 not n40020 ; n40020_not
g50011 not n10140 ; n10140_not
g50012 not n30012 ; n30012_not
g50013 not n20400 ; n20400_not
g50014 not n10005 ; n10005_not
g50015 not n21201 ; n21201_not
g50016 not n31200 ; n31200_not
g50017 not n10023 ; n10023_not
g50018 not n20310 ; n20310_not
g50019 not n11130 ; n11130_not
g50020 not n10320 ; n10320_not
g50021 not n20121 ; n20121_not
g50022 not n10032 ; n10032_not
g50023 not n10302 ; n10302_not
g50024 not n10401 ; n10401_not
g50025 not n24000 ; n24000_not
g50026 not n10041 ; n10041_not
g50027 not n20301 ; n20301_not
g50028 not n22110 ; n22110_not
g50029 not n21112 ; n21112_not
g50030 not n23020 ; n23020_not
g50031 not n10312 ; n10312_not
g50032 not n30022 ; n30022_not
g50033 not n31003 ; n31003_not
g50034 not n12103 ; n12103_not
g50035 not n13111 ; n13111_not
g50036 not n21103 ; n21103_not
g50037 not n22210 ; n22210_not
g50038 not n42100 ; n42100_not
g50039 not n40111 ; n40111_not
g50040 not n11500 ; n11500_not
g50041 not n10321 ; n10321_not
g50042 not n23200 ; n23200_not
g50043 not n12040 ; n12040_not
g50044 not n11230 ; n11230_not
g50045 not n41110 ; n41110_not
g50046 not n41002 ; n41002_not
g50047 not n23002 ; n23002_not
g50048 not n12022 ; n12022_not
g50049 not n10330 ; n10330_not
g50050 not n10204 ; n10204_not
g50051 not n41011 ; n41011_not
g50052 not n21004 ; n21004_not
g50053 not n10510 ; n10510_not
g50054 not n14101 ; n14101_not
g50055 not n12310 ; n12310_not
g50056 not n12211 ; n12211_not
g50057 not n14020 ; n14020_not
g50058 not n22102 ; n22102_not
g50059 not n14002 ; n14002_not
g50060 not n11113 ; n11113_not
g50061 not n31102 ; n31102_not
g50062 not n11140 ; n11140_not
g50063 not n12220 ; n12220_not
g50064 not n11131 ; n11131_not
g50065 not n11122 ; n11122_not
g50066 not n12301 ; n12301_not
g50067 not n11032 ; n11032_not
g50068 not n11320 ; n11320_not
g50069 not n25000 ; n25000_not
g50070 not n21400 ; n21400_not
g50071 not n31210 ; n31210_not
g50072 not n16000 ; n16000_not
g50073 not n15010 ; n15010_not
g50074 not n31021 ; n31021_not
g50075 not n10411 ; n10411_not
g50076 not n23011 ; n23011_not
g50077 not n13021 ; n13021_not
g50078 not n32101 ; n32101_not
g50079 not n12112 ; n12112_not
g50080 not n13012 ; n13012_not
g50081 not n31030 ; n31030_not
g50082 not n34000 ; n34000_not
g50083 not n13300 ; n13300_not
g50084 not n13003 ; n13003_not
g50085 not n12121 ; n12121_not
g50086 not n11401 ; n11401_not
g50087 not n31120 ; n31120_not
g50088 not n21040 ; n21040_not
g50089 not n21121 ; n21121_not
g50090 not n10123 ; n10123_not
g50091 not n10105 ; n10105_not
g50092 not n10006 ; n10006_not
g50093 not n40012 ; n40012_not
g50094 not n40021 ; n40021_not
g50095 not n30103 ; n30103_not
g50096 not n21202 ; n21202_not
g50097 not n20320 ; n20320_not
g50098 not n40300 ; n40300_not
g50099 not n30202 ; n30202_not
g50100 not n10042 ; n10042_not
g50101 not n20230 ; n20230_not
g50102 not n10213 ; n10213_not
g50103 not n21301 ; n21301_not
g50104 not n20140 ; n20140_not
g50105 not n40120 ; n40120_not
g50106 not n10051 ; n10051_not
g50107 not n20005 ; n20005_not
g50108 not n21014 ; n21014_not
g50109 not n15020 ; n15020_not
g50110 not n15002 ; n15002_not
g50111 not n11114 ; n11114_not
g50112 not n31013 ; n31013_not
g50113 not n22031 ; n22031_not
g50114 not n15011 ; n15011_not
g50115 not n10106 ; n10106_not
g50116 not n12050 ; n12050_not
g50117 not n20024 ; n20024_not
g50118 not n43100 ; n43100_not
g50119 not n41012 ; n41012_not
g50120 not n34100 ; n34100_not
g50121 not n11204 ; n11204_not
g50122 not n20501 ; n20501_not
g50123 not n31031 ; n31031_not
g50124 not n22022 ; n22022_not
g50125 not n22004 ; n22004_not
g50126 not n42011 ; n42011_not
g50127 not n20510 ; n20510_not
g50128 not n32030 ; n32030_not
g50129 not n10520 ; n10520_not
g50130 not n23030 ; n23030_not
g50131 not n30122 ; n30122_not
g50132 not n40130 ; n40130_not
g50133 not n40121 ; n40121_not
g50134 not n31220 ; n31220_not
g50135 not n40112 ; n40112_not
g50136 not n23021 ; n23021_not
g50137 not n11240 ; n11240_not
g50138 not n10160 ; n10160_not
g50139 not n16100 ; n16100_not
g50140 not n22400 ; n22400_not
g50141 not n42200 ; n42200_not
g50142 not n12005 ; n12005_not
g50143 not n30005 ; n30005_not
g50144 not n40013 ; n40013_not
g50145 not n32201 ; n32201_not
g50146 not n30104 ; n30104_not
g50147 not n10115 ; n10115_not
g50148 not n13202 ; n13202_not
g50149 not n30140 ; n30140_not
g50150 not n21050 ; n21050_not
g50151 not n20114 ; n20114_not
g50152 not n33110 ; n33110_not
g50153 not n10601 ; n10601_not
g50154 not n22211 ; n22211_not
g50155 not n12311 ; n12311_not
g50156 not n30230 ; n30230_not
g50157 not n30221 ; n30221_not
g50158 not n12320 ; n12320_not
g50159 not n12410 ; n12410_not
g50160 not n20231 ; n20231_not
g50161 not n24110 ; n24110_not
g50162 not n11024 ; n11024_not
g50163 not n12302 ; n12302_not
g50164 not n30050 ; n30050_not
g50165 not n11033 ; n11033_not
g50166 not n24101 ; n24101_not
g50167 not n11042 ; n11042_not
g50168 not n12500 ; n12500_not
g50169 not n22301 ; n22301_not
g50170 not n22040 ; n22040_not
g50171 not n14111 ; n14111_not
g50172 not n14102 ; n14102_not
g50173 not n20033 ; n20033_not
g50174 not n10061 ; n10061_not
g50175 not n21104 ; n21104_not
g50176 not n21311 ; n21311_not
g50177 not n10052 ; n10052_not
g50178 not n12113 ; n12113_not
g50179 not n14012 ; n14012_not
g50180 not n12122 ; n12122_not
g50181 not n20060 ; n20060_not
g50182 not n30212 ; n30212_not
g50183 not n30203 ; n30203_not
g50184 not n31112 ; n31112_not
g50185 not n12140 ; n12140_not
g50186 not n21041 ; n21041_not
g50187 not n31211 ; n31211_not
g50188 not n11141 ; n11141_not
g50189 not n21401 ; n21401_not
g50190 not n33011 ; n33011_not
g50191 not n33101 ; n33101_not
g50192 not n24011 ; n24011_not
g50193 not n13310 ; n13310_not
g50194 not n12230 ; n12230_not
g50195 not n10403 ; n10403_not
g50196 not n13220 ; n13220_not
g50197 not n32012 ; n32012_not
g50198 not n30401 ; n30401_not
g50199 not n11600 ; n11600_not
g50200 not n40211 ; n40211_not
g50201 not n23102 ; n23102_not
g50202 not n11312 ; n11312_not
g50203 not n41111 ; n41111_not
g50204 not n20303 ; n20303_not
g50205 not n17000 ; n17000_not
g50206 not n10340 ; n10340_not
g50207 not n10223 ; n10223_not
g50208 not n21230 ; n21230_not
g50209 not n20222 ; n20222_not
g50210 not n10421 ; n10421_not
g50211 not n31301 ; n31301_not
g50212 not n20213 ; n20213_not
g50213 not n30032 ; n30032_not
g50214 not n30410 ; n30410_not
g50215 not n41300 ; n41300_not
g50216 not n31400 ; n31400_not
g50217 not n30320 ; n30320_not
g50218 not n30311 ; n30311_not
g50219 not n11501 ; n11501_not
g50220 not n30113 ; n30113_not
g50221 not n26000 ; n26000_not
g50222 not n33020 ; n33020_not
g50223 not n10017 ; n10017_not
g50224 not n22131 ; n22131_not
g50225 not n21114 ; n21114_not
g50226 not n10026 ; n10026_not
g50227 not n25101 ; n25101_not
g50228 not n10233 ; n10233_not
g50229 not n41202 ; n41202_not
g50230 not n32211 ; n32211_not
g50231 not n20052 ; n20052_not
g50232 not n30330 ; n30330_not
g50233 not n34011 ; n34011_not
g50234 not n20106 ; n20106_not
g50235 not n12402 ; n12402_not
g50236 not n30132 ; n30132_not
g50237 not n24300 ; n24300_not
g50238 not n30222 ; n30222_not
g50239 not n10350 ; n10350_not
g50240 not n41130 ; n41130_not
g50241 not n40401 ; n40401_not
g50242 not n30114 ; n30114_not
g50243 not n31113 ; n31113_not
g50244 not n12213 ; n12213_not
g50245 not n13500 ; n13500_not
g50246 not n22320 ; n22320_not
g50247 not n10224 ; n10224_not
g50248 not n23400 ; n23400_not
g50249 not n14121 ; n14121_not
g50250 not n44100 ; n44100_not
g50251 not n20232 ; n20232_not
g50252 not n32301 ; n32301_not
g50253 not n10062 ; n10062_not
g50254 not n18000 ; n18000_not
g50255 not n20304 ; n20304_not
g50256 not n22050 ; n22050_not
g50257 not n12105 ; n12105_not
g50258 not n20133 ; n20133_not
g50259 not n20412 ; n20412_not
g50260 not n14040 ; n14040_not
g50261 not n20223 ; n20223_not
g50262 not n12042 ; n12042_not
g50263 not n41220 ; n41220_not
g50264 not n20043 ; n20043_not
g50265 not n32121 ; n32121_not
g50266 not n12123 ; n12123_not
g50267 not n21024 ; n21024_not
g50268 not n40131 ; n40131_not
g50269 not n21222 ; n21222_not
g50270 not n20124 ; n20124_not
g50271 not n25200 ; n25200_not
g50272 not n24030 ; n24030_not
g50273 not n23004 ; n23004_not
g50274 not n41031 ; n41031_not
g50275 not n20403 ; n20403_not
g50276 not n10332 ; n10332_not
g50277 not n21420 ; n21420_not
g50278 not n40302 ; n40302_not
g50279 not n21402 ; n21402_not
g50280 not n41022 ; n41022_not
g50281 not n33120 ; n33120_not
g50282 not n21213 ; n21213_not
g50283 not n13014 ; n13014_not
g50284 not n11115 ; n11115_not
g50285 not n11511 ; n11511_not
g50286 not n26010 ; n26010_not
g50287 not n40320 ; n40320_not
g50288 not n25020 ; n25020_not
g50289 not n34020 ; n34020_not
g50290 not n32130 ; n32130_not
g50291 not n20340 ; n20340_not
g50292 not n12312 ; n12312_not
g50293 not n10314 ; n10314_not
g50294 not n12321 ; n12321_not
g50295 not n21312 ; n21312_not
g50296 not n20322 ; n20322_not
g50297 not n22203 ; n22203_not
g50298 not n13410 ; n13410_not
g50299 not n33003 ; n33003_not
g50300 not n21150 ; n21150_not
g50301 not n11025 ; n11025_not
g50302 not n24021 ; n24021_not
g50303 not n13311 ; n13311_not
g50304 not n13320 ; n13320_not
g50305 not n10341 ; n10341_not
g50306 not n34002 ; n34002_not
g50307 not n10305 ; n10305_not
g50308 not n11601 ; n11601_not
g50309 not n21033 ; n21033_not
g50310 not n33012 ; n33012_not
g50311 not n13212 ; n13212_not
g50312 not n24012 ; n24012_not
g50313 not n12303 ; n12303_not
g50314 not n13230 ; n13230_not
g50315 not n30402 ; n30402_not
g50316 not n40140 ; n40140_not
g50317 not n17010 ; n17010_not
g50318 not n21303 ; n21303_not
g50319 not n16011 ; n16011_not
g50320 not n10215 ; n10215_not
g50321 not n31131 ; n31131_not
g50322 not n11241 ; n11241_not
g50323 not n16002 ; n16002_not
g50324 not n40041 ; n40041_not
g50325 not n30015 ; n30015_not
g50326 not n40032 ; n40032_not
g50327 not n12006 ; n12006_not
g50328 not n42300 ; n42300_not
g50329 not n10620 ; n10620_not
g50330 not n31023 ; n31023_not
g50331 not n15021 ; n15021_not
g50332 not n10116 ; n10116_not
g50333 not n15102 ; n15102_not
g50334 not n12024 ; n12024_not
g50335 not n15111 ; n15111_not
g50336 not n20313 ; n20313_not
g50337 not n15210 ; n15210_not
g50338 not n11232 ; n11232_not
g50339 not n44001 ; n44001_not
g50340 not n15300 ; n15300_not
g50341 not n34110 ; n34110_not
g50342 not n10521 ; n10521_not
g50343 not n10440 ; n10440_not
g50344 not n22500 ; n22500_not
g50345 not n20601 ; n20601_not
g50346 not n42012 ; n42012_not
g50347 not n10206 ; n10206_not
g50348 not n23040 ; n23040_not
g50349 not n32031 ; n32031_not
g50350 not n10512 ; n10512_not
g50351 not n22401 ; n22401_not
g50352 not n42021 ; n42021_not
g50353 not n30033 ; n30033_not
g50354 not n42030 ; n42030_not
g50355 not n21141 ; n21141_not
g50356 not n23022 ; n23022_not
g50357 not n32112 ; n32112_not
g50358 not n16101 ; n16101_not
g50359 not n11304 ; n11304_not
g50360 not n16110 ; n16110_not
g50361 not n15003 ; n15003_not
g50362 not n31500 ; n31500_not
g50363 not n16200 ; n16200_not
g50364 not n24003 ; n24003_not
g50365 not n21132 ; n21132_not
g50366 not n31005 ; n31005_not
g50367 not n42111 ; n42111_not
g50368 not n42120 ; n42120_not
g50369 not n42102 ; n42102_not
g50370 not n30123 ; n30123_not
g50371 not n10530 ; n10530_not
g50372 not n17001 ; n17001_not
g50373 not n12051 ; n12051_not
g50374 not n10710 ; n10710_not
g50375 not n20610 ; n20610_not
g50376 not n23202 ; n23202_not
g50377 not n43110 ; n43110_not
g50378 not n40005 ; n40005_not
g50379 not n11223 ; n11223_not
g50380 not n20502 ; n20502_not
g50381 not n20205 ; n20205_not
g50382 not n11205 ; n11205_not
g50383 not n43011 ; n43011_not
g50384 not n11331 ; n11331_not
g50385 not n26001 ; n26001_not
g50386 not n10071 ; n10071_not
g50387 not n22005 ; n22005_not
g50388 not n43101 ; n43101_not
g50389 not n30510 ; n30510_not
g50390 not n20016 ; n20016_not
g50391 not n10431 ; n10431_not
g50392 not n12033 ; n12033_not
g50393 not n23112 ; n23112_not
g50394 not n21123 ; n21123_not
g50395 not n14211 ; n14211_not
g50396 not n11322 ; n11322_not
g50397 not n12060 ; n12060_not
g50398 not n10107 ; n10107_not
g50399 not n14202 ; n14202_not
g50400 not n23130 ; n23130_not
g50401 not n43210 ; n43210_not
g50402 not n20233 ; n20233_not
g50403 not n20314 ; n20314_not
g50404 not n22330 ; n22330_not
g50405 not n21304 ; n21304_not
g50406 not n12313 ; n12313_not
g50407 not n31411 ; n31411_not
g50408 not n22411 ; n22411_not
g50409 not n31222 ; n31222_not
g50410 not n10810 ; n10810_not
g50411 not n12043 ; n12043_not
g50412 not n20152 ; n20152_not
g50413 not n11710 ; n11710_not
g50414 not n20305 ; n20305_not
g50415 not n31231 ; n31231_not
g50416 not n12403 ; n12403_not
g50417 not n31402 ; n31402_not
g50418 not n32221 ; n32221_not
g50419 not n32014 ; n32014_not
g50420 not n12070 ; n12070_not
g50421 not n11431 ; n11431_not
g50422 not n20143 ; n20143_not
g50423 not n32410 ; n32410_not
g50424 not n34021 ; n34021_not
g50425 not n31420 ; n31420_not
g50426 not n12133 ; n12133_not
g50427 not n20323 ; n20323_not
g50428 not n24130 ; n24130_not
g50429 not n12232 ; n12232_not
g50430 not n11620 ; n11620_not
g50431 not n10108 ; n10108_not
g50432 not n11800 ; n11800_not
g50433 not n12223 ; n12223_not
g50434 not n22510 ; n22510_not
g50435 not n31213 ; n31213_not
g50436 not n30205 ; n30205_not
g50437 not n12025 ; n12025_not
g50438 not n33130 ; n33130_not
g50439 not n12205 ; n12205_not
g50440 not n32311 ; n32311_not
g50441 not n12304 ; n12304_not
g50442 not n32320 ; n32320_not
g50443 not n31312 ; n31312_not
g50444 not n12007 ; n12007_not
g50445 not n44020 ; n44020_not
g50446 not n30061 ; n30061_not
g50447 not n22402 ; n22402_not
g50448 not n20134 ; n20134_not
g50449 not n12115 ; n12115_not
g50450 not n33040 ; n33040_not
g50451 not n11521 ; n11521_not
g50452 not n12250 ; n12250_not
g50453 not n33310 ; n33310_not
g50454 not n12124 ; n12124_not
g50455 not n12241 ; n12241_not
g50456 not n20125 ; n20125_not
g50457 not n12034 ; n12034_not
g50458 not n32302 ; n32302_not
g50459 not n42112 ; n42112_not
g50460 not n40114 ; n40114_not
g50461 not n30025 ; n30025_not
g50462 not n42103 ; n42103_not
g50463 not n21142 ; n21142_not
g50464 not n40132 ; n40132_not
g50465 not n23041 ; n23041_not
g50466 not n40150 ; n40150_not
g50467 not n42004 ; n42004_not
g50468 not n21700 ; n21700_not
g50469 not n21601 ; n21601_not
g50470 not n21610 ; n21610_not
g50471 not n21520 ; n21520_not
g50472 not n40303 ; n40303_not
g50473 not n40060 ; n40060_not
g50474 not n17011 ; n17011_not
g50475 not n21511 ; n21511_not
g50476 not n36001 ; n36001_not
g50477 not n43003 ; n43003_not
g50478 not n40006 ; n40006_not
g50479 not n15013 ; n15013_not
g50480 not n15040 ; n15040_not
g50481 not n15112 ; n15112_not
g50482 not n15121 ; n15121_not
g50483 not n15220 ; n15220_not
g50484 not n10603 ; n10603_not
g50485 not n15400 ; n15400_not
g50486 not n40024 ; n40024_not
g50487 not n20530 ; n20530_not
g50488 not n42310 ; n42310_not
g50489 not n34201 ; n34201_not
g50490 not n40033 ; n40033_not
g50491 not n40105 ; n40105_not
g50492 not n16003 ; n16003_not
g50493 not n16012 ; n16012_not
g50494 not n16111 ; n16111_not
g50495 not n16120 ; n16120_not
g50496 not n16300 ; n16300_not
g50497 not n42130 ; n42130_not
g50498 not n40411 ; n40411_not
g50499 not n40231 ; n40231_not
g50500 not n41140 ; n41140_not
g50501 not n41113 ; n41113_not
g50502 not n30043 ; n30043_not
g50503 not n41014 ; n41014_not
g50504 not n41032 ; n41032_not
g50505 not n41023 ; n41023_not
g50506 not n40321 ; n40321_not
g50507 not n40330 ; n40330_not
g50508 not n21421 ; n21421_not
g50509 not n30340 ; n30340_not
g50510 not n30331 ; n30331_not
g50511 not n19000 ; n19000_not
g50512 not n40420 ; n40420_not
g50513 not n17101 ; n17101_not
g50514 not n40222 ; n40222_not
g50515 not n41311 ; n41311_not
g50516 not n30601 ; n30601_not
g50517 not n30502 ; n30502_not
g50518 not n30304 ; n30304_not
g50519 not n23212 ; n23212_not
g50520 not n23401 ; n23401_not
g50521 not n30430 ; n30430_not
g50522 not n27100 ; n27100_not
g50523 not n41410 ; n41410_not
g50524 not n18001 ; n18001_not
g50525 not n18010 ; n18010_not
g50526 not n23410 ; n23410_not
g50527 not n32131 ; n32131_not
g50528 not n41212 ; n41212_not
g50529 not n20350 ; n20350_not
g50530 not n13105 ; n13105_not
g50531 not n21025 ; n21025_not
g50532 not n13141 ; n13141_not
g50533 not n11422 ; n11422_not
g50534 not n13213 ; n13213_not
g50535 not n22204 ; n22204_not
g50536 not n20422 ; n20422_not
g50537 not n13303 ; n13303_not
g50538 not n13330 ; n13330_not
g50539 not n13312 ; n13312_not
g50540 not n21403 ; n21403_not
g50541 not n21070 ; n21070_not
g50542 not n13501 ; n13501_not
g50543 not n10504 ; n10504_not
g50544 not n21160 ; n21160_not
g50545 not n32005 ; n32005_not
g50546 not n13600 ; n13600_not
g50547 not n12421 ; n12421_not
g50548 not n21052 ; n21052_not
g50549 not n32230 ; n32230_not
g50550 not n24040 ; n24040_not
g50551 not n35110 ; n35110_not
g50552 not n31204 ; n31204_not
g50553 not n35020 ; n35020_not
g50554 not n24031 ; n24031_not
g50555 not n31132 ; n31132_not
g50556 not n21340 ; n21340_not
g50557 not n26200 ; n26200_not
g50558 not n25003 ; n25003_not
g50559 not n35002 ; n35002_not
g50560 not n25012 ; n25012_not
g50561 not n22240 ; n22240_not
g50562 not n22231 ; n22231_not
g50563 not n22222 ; n22222_not
g50564 not n32212 ; n32212_not
g50565 not n20332 ; n20332_not
g50566 not n13024 ; n13024_not
g50567 not n14050 ; n14050_not
g50568 not n20008 ; n20008_not
g50569 not n22060 ; n22060_not
g50570 not n22051 ; n22051_not
g50571 not n22042 ; n22042_not
g50572 not n20710 ; n20710_not
g50573 not n22033 ; n22033_not
g50574 not n14131 ; n14131_not
g50575 not n14140 ; n14140_not
g50576 not n20026 ; n20026_not
g50577 not n14212 ; n14212_not
g50578 not n14221 ; n14221_not
g50579 not n14041 ; n14041_not
g50580 not n20620 ; n20620_not
g50581 not n31060 ; n31060_not
g50582 not n14320 ; n14320_not
g50583 not n26011 ; n26011_not
g50584 not n31051 ; n31051_not
g50585 not n14410 ; n14410_not
g50586 not n43021 ; n43021_not
g50587 not n36010 ; n36010_not
g50588 not n34030 ; n34030_not
g50589 not n22141 ; n22141_not
g50590 not n21412 ; n21412_not
g50591 not n22132 ; n22132_not
g50592 not n20800 ; n20800_not
g50593 not n20062 ; n20062_not
g50594 not n34012 ; n34012_not
g50595 not n25102 ; n25102_not
g50596 not n20053 ; n20053_not
g50597 not n22123 ; n22123_not
g50598 not n22114 ; n22114_not
g50599 not n22105 ; n22105_not
g50600 not n14005 ; n14005_not
g50601 not n14014 ; n14014_not
g50602 not n20044 ; n20044_not
g50603 not n25201 ; n25201_not
g50604 not n26020 ; n26020_not
g50605 not n14032 ; n14032_not
g50606 not n10801 ; n10801_not
g50607 not n44200 ; n44200_not
g50608 not n10711 ; n10711_not
g50609 not n11080 ; n11080_not
g50610 not n10450 ; n10450_not
g50611 not n11134 ; n11134_not
g50612 not n11071 ; n11071_not
g50613 not n10117 ; n10117_not
g50614 not n10018 ; n10018_not
g50615 not n11233 ; n11233_not
g50616 not n10612 ; n10612_not
g50617 not n11341 ; n11341_not
g50618 not n10720 ; n10720_not
g50619 not n10126 ; n10126_not
g50620 not n10135 ; n10135_not
g50621 not n10306 ; n10306_not
g50622 not n10540 ; n10540_not
g50623 not n10261 ; n10261_not
g50624 not n10090 ; n10090_not
g50625 not n10009 ; n10009_not
g50626 not n11350 ; n11350_not
g50627 not n11206 ; n11206_not
g50628 not n10063 ; n10063_not
g50629 not n10360 ; n10360_not
g50630 not n10144 ; n10144_not
g50631 not n10072 ; n10072_not
g50632 not n10045 ; n10045_not
g50633 not n10441 ; n10441_not
g50634 not n11170 ; n11170_not
g50635 not n10270 ; n10270_not
g50636 not n30413 ; n30413_not
g50637 not n26102 ; n26102_not
g50638 not n22421 ; n22421_not
g50639 not n22430 ; n22430_not
g50640 not n20171 ; n20171_not
g50641 not n20162 ; n20162_not
g50642 not n30350 ; n30350_not
g50643 not n30341 ; n30341_not
g50644 not n30503 ; n30503_not
g50645 not n20207 ; n20207_not
g50646 not n20261 ; n20261_not
g50647 not n34103 ; n34103_not
g50648 not n12611 ; n12611_not
g50649 not n20243 ; n20243_not
g50650 not n21071 ; n21071_not
g50651 not n30440 ; n30440_not
g50652 not n22403 ; n22403_not
g50653 not n20225 ; n20225_not
g50654 not n30422 ; n30422_not
g50655 not n20216 ; n20216_not
g50656 not n26111 ; n26111_not
g50657 not n34022 ; n34022_not
g50658 not n26003 ; n26003_not
g50659 not n30161 ; n30161_not
g50660 not n30242 ; n30242_not
g50661 not n20018 ; n20018_not
g50662 not n13214 ; n13214_not
g50663 not n30251 ; n30251_not
g50664 not n22511 ; n22511_not
g50665 not n30260 ; n30260_not
g50666 not n22502 ; n22502_not
g50667 not n10028 ; n10028_not
g50668 not n13160 ; n13160_not
g50669 not n20072 ; n20072_not
g50670 not n13142 ; n13142_not
g50671 not n13124 ; n13124_not
g50672 not n10451 ; n10451_not
g50673 not n20081 ; n20081_not
g50674 not n13106 ; n13106_not
g50675 not n34004 ; n34004_not
g50676 not n17021 ; n17021_not
g50677 not n42500 ; n42500_not
g50678 not n13070 ; n13070_not
g50679 not n17003 ; n17003_not
g50680 not n13016 ; n13016_not
g50681 not n30215 ; n30215_not
g50682 not n34031 ; n34031_not
g50683 not n20144 ; n20144_not
g50684 not n13007 ; n13007_not
g50685 not n30314 ; n30314_not
g50686 not n30323 ; n30323_not
g50687 not n20153 ; n20153_not
g50688 not n12224 ; n12224_not
g50689 not n11135 ; n11135_not
g50690 not n11126 ; n11126_not
g50691 not n22016 ; n22016_not
g50692 not n12305 ; n12305_not
g50693 not n20702 ; n20702_not
g50694 not n22043 ; n22043_not
g50695 not n12332 ; n12332_not
g50696 not n12350 ; n12350_not
g50697 not n22070 ; n22070_not
g50698 not n42311 ; n42311_not
g50699 not n20513 ; n20513_not
g50700 not n11072 ; n11072_not
g50701 not n20630 ; n20630_not
g50702 not n31601 ; n31601_not
g50703 not n20621 ; n20621_not
g50704 not n12440 ; n12440_not
g50705 not n22106 ; n22106_not
g50706 not n42221 ; n42221_not
g50707 not n12071 ; n12071_not
g50708 not n31034 ; n31034_not
g50709 not n35030 ; n35030_not
g50710 not n31025 ; n31025_not
g50711 not n12080 ; n12080_not
g50712 not n31016 ; n31016_not
g50713 not n20900 ; n20900_not
g50714 not n46010 ; n46010_not
g50715 not n16400 ; n16400_not
g50716 not n12116 ; n12116_not
g50717 not n11153 ; n11153_not
g50718 not n12152 ; n12152_not
g50719 not n12161 ; n12161_not
g50720 not n35111 ; n35111_not
g50721 not n31502 ; n31502_not
g50722 not n31511 ; n31511_not
g50723 not n20801 ; n20801_not
g50724 not n30620 ; n30620_not
g50725 not n30611 ; n30611_not
g50726 not n12701 ; n12701_not
g50727 not n30602 ; n30602_not
g50728 not n22322 ; n22322_not
g50729 not n40160 ; n40160_not
g50730 not n20360 ; n20360_not
g50731 not n20333 ; n20333_not
g50732 not n20342 ; n20342_not
g50733 not n10910 ; n10910_not
g50734 not n20324 ; n20324_not
g50735 not n22340 ; n22340_not
g50736 not n34130 ; n34130_not
g50737 not n30512 ; n30512_not
g50738 not n34121 ; n34121_not
g50739 not n20603 ; n20603_not
g50740 not n22115 ; n22115_not
g50741 not n42032 ; n42032_not
g50742 not n10622 ; n10622_not
g50743 not n22124 ; n22124_not
g50744 not n12521 ; n12521_not
g50745 not n40124 ; n40124_not
g50746 not n20531 ; n20531_not
g50747 not n20522 ; n20522_not
g50748 not n30701 ; n30701_not
g50749 not n22250 ; n22250_not
g50750 not n20450 ; n20450_not
g50751 not n42410 ; n42410_not
g50752 not n20432 ; n20432_not
g50753 not n12602 ; n12602_not
g50754 not n22232 ; n22232_not
g50755 not n20414 ; n20414_not
g50756 not n40610 ; n40610_not
g50757 not n19001 ; n19001_not
g50758 not n33401 ; n33401_not
g50759 not n15023 ; n15023_not
g50760 not n41411 ; n41411_not
g50761 not n15113 ; n15113_not
g50762 not n32501 ; n32501_not
g50763 not n14213 ; n14213_not
g50764 not n41402 ; n41402_not
g50765 not n37100 ; n37100_not
g50766 not n14231 ; n14231_not
g50767 not n14240 ; n14240_not
g50768 not n40601 ; n40601_not
g50769 not n40151 ; n40151_not
g50770 not n25013 ; n25013_not
g50771 not n14303 ; n14303_not
g50772 not n10721 ; n10721_not
g50773 not n23420 ; n23420_not
g50774 not n25211 ; n25211_not
g50775 not n17300 ; n17300_not
g50776 not n10163 ; n10163_not
g50777 not n10820 ; n10820_not
g50778 not n40403 ; n40403_not
g50779 not n15212 ; n15212_not
g50780 not n41510 ; n41510_not
g50781 not n14033 ; n14033_not
g50782 not n14042 ; n14042_not
g50783 not n14051 ; n14051_not
g50784 not n40412 ; n40412_not
g50785 not n23600 ; n23600_not
g50786 not n41420 ; n41420_not
g50787 not n19010 ; n19010_not
g50788 not n15131 ; n15131_not
g50789 not n14123 ; n14123_not
g50790 not n33221 ; n33221_not
g50791 not n14600 ; n14600_not
g50792 not n10370 ; n10370_not
g50793 not n24401 ; n24401_not
g50794 not n41042 ; n41042_not
g50795 not n41051 ; n41051_not
g50796 not n33203 ; n33203_not
g50797 not n29000 ; n29000_not
g50798 not n10703 ; n10703_not
g50799 not n43040 ; n43040_not
g50800 not n33041 ; n33041_not
g50801 not n41141 ; n41141_not
g50802 not n43013 ; n43013_not
g50803 not n33104 ; n33104_not
g50804 not n33032 ; n33032_not
g50805 not n33122 ; n33122_not
g50806 not n33113 ; n33113_not
g50807 not n14330 ; n14330_not
g50808 not n25004 ; n25004_not
g50809 not n37001 ; n37001_not
g50810 not n41312 ; n41312_not
g50811 not n41303 ; n41303_not
g50812 not n10712 ; n10712_not
g50813 not n24104 ; n24104_not
g50814 not n43121 ; n43121_not
g50815 not n43112 ; n43112_not
g50816 not n24113 ; n24113_not
g50817 not n24122 ; n24122_not
g50818 not n13061 ; n13061_not
g50819 not n33302 ; n33302_not
g50820 not n14501 ; n14501_not
g50821 not n41114 ; n41114_not
g50822 not n24302 ; n24302_not
g50823 not n24311 ; n24311_not
g50824 not n23006 ; n23006_not
g50825 not n41105 ; n41105_not
g50826 not n17201 ; n17201_not
g50827 not n23033 ; n23033_not
g50828 not n23042 ; n23042_not
g50829 not n10460 ; n10460_not
g50830 not n28010 ; n28010_not
g50831 not n30053 ; n30053_not
g50832 not n10532 ; n10532_not
g50833 not n30044 ; n30044_not
g50834 not n23105 ; n23105_not
g50835 not n10505 ; n10505_not
g50836 not n30035 ; n30035_not
g50837 not n13520 ; n13520_not
g50838 not n10127 ; n10127_not
g50839 not n30008 ; n30008_not
g50840 not n23123 ; n23123_not
g50841 not n15221 ; n15221_not
g50842 not n17102 ; n17102_not
g50843 not n20009 ; n20009_not
g50844 not n17120 ; n17120_not
g50845 not n13304 ; n13304_not
g50846 not n30170 ; n30170_not
g50847 not n13313 ; n13313_not
g50848 not n30134 ; n30134_not
g50849 not n30125 ; n30125_not
g50850 not n22700 ; n22700_not
g50851 not n30116 ; n30116_not
g50852 not n30107 ; n30107_not
g50853 not n10433 ; n10433_not
g50854 not n32150 ; n32150_not
g50855 not n23240 ; n23240_not
g50856 not n40205 ; n40205_not
g50857 not n40232 ; n40232_not
g50858 not n32204 ; n32204_not
g50859 not n32213 ; n32213_not
g50860 not n40241 ; n40241_not
g50861 not n40250 ; n40250_not
g50862 not n23312 ; n23312_not
g50863 not n36101 ; n36101_not
g50864 not n32240 ; n32240_not
g50865 not n41600 ; n41600_not
g50866 not n43301 ; n43301_not
g50867 not n40313 ; n40313_not
g50868 not n32321 ; n32321_not
g50869 not n33500 ; n33500_not
g50870 not n23321 ; n23321_not
g50871 not n40331 ; n40331_not
g50872 not n40034 ; n40034_not
g50873 not n40043 ; n40043_not
g50874 not n40070 ; n40070_not
g50875 not n32024 ; n32024_not
g50876 not n43400 ; n43400_not
g50877 not n40106 ; n40106_not
g50878 not n32105 ; n32105_not
g50879 not n23213 ; n23213_not
g50880 not n13700 ; n13700_not
g50881 not n23222 ; n23222_not
g50882 not n32132 ; n32132_not
g50883 not n32141 ; n32141_not
g50884 not n16031 ; n16031_not
g50885 not n21062 ; n21062_not
g50886 not n21701 ; n21701_not
g50887 not n11243 ; n11243_not
g50888 not n21206 ; n21206_not
g50889 not n31151 ; n31151_not
g50890 not n21242 ; n21242_not
g50891 not n21503 ; n21503_not
g50892 not n27110 ; n27110_not
g50893 not n21161 ; n21161_not
g50894 not n21215 ; n21215_not
g50895 not n11225 ; n11225_not
g50896 not n44111 ; n44111_not
g50897 not n21530 ; n21530_not
g50898 not n11405 ; n11405_not
g50899 not n11900 ; n11900_not
g50900 not n21143 ; n21143_not
g50901 not n11234 ; n11234_not
g50902 not n21350 ; n21350_not
g50903 not n16103 ; n16103_not
g50904 not n11504 ; n11504_not
g50905 not n11441 ; n11441_not
g50906 not n42140 ; n42140_not
g50907 not n21125 ; n21125_not
g50908 not n44012 ; n44012_not
g50909 not n31070 ; n31070_not
g50910 not n31340 ; n31340_not
g50911 not n44102 ; n44102_not
g50912 not n44030 ; n44030_not
g50913 not n10217 ; n10217_not
g50914 not n44003 ; n44003_not
g50915 not n11720 ; n11720_not
g50916 not n21233 ; n21233_not
g50917 not n11702 ; n11702_not
g50918 not n11513 ; n11513_not
g50919 not n21710 ; n21710_not
g50920 not n11810 ; n11810_not
g50921 not n21521 ; n21521_not
g50922 not n27002 ; n27002_not
g50923 not n11801 ; n11801_not
g50924 not n31430 ; n31430_not
g50925 not n11621 ; n11621_not
g50926 not n27020 ; n27020_not
g50927 not n31331 ; n31331_not
g50928 not n11252 ; n11252_not
g50929 not n21080 ; n21080_not
g50930 not n10523 ; n10523_not
g50931 not n11315 ; n11315_not
g50932 not n11216 ; n11216_not
g50933 not n31250 ; n31250_not
g50934 not n31124 ; n31124_not
g50935 not n31241 ; n31241_not
g50936 not n11414 ; n11414_not
g50937 not n21800 ; n21800_not
g50938 not n42203 ; n42203_not
g50939 not n12008 ; n12008_not
g50940 not n42122 ; n42122_not
g50941 not n35003 ; n35003_not
g50942 not n16211 ; n16211_not
g50943 not n13017 ; n13017_not
g50944 not n21162 ; n21162_not
g50945 not n40431 ; n40431_not
g50946 not n40440 ; n40440_not
g50947 not n13008 ; n13008_not
g50948 not n21153 ; n21153_not
g50949 not n23610 ; n23610_not
g50950 not n20235 ; n20235_not
g50951 not n41421 ; n41421_not
g50952 not n30324 ; n30324_not
g50953 not n15150 ; n15150_not
g50954 not n36111 ; n36111_not
g50955 not n15141 ; n15141_not
g50956 not n10452 ; n10452_not
g50957 not n10038 ; n10038_not
g50958 not n10029 ; n10029_not
g50959 not n16302 ; n16302_not
g50960 not n13161 ; n13161_not
g50961 not n11811 ; n11811_not
g50962 not n13152 ; n13152_not
g50963 not n25140 ; n25140_not
g50964 not n13143 ; n13143_not
g50965 not n17031 ; n17031_not
g50966 not n16311 ; n16311_not
g50967 not n40143 ; n40143_not
g50968 not n25131 ; n25131_not
g50969 not n13134 ; n13134_not
g50970 not n16320 ; n16320_not
g50971 not n32430 ; n32430_not
g50972 not n30270 ; n30270_not
g50973 not n14115 ; n14115_not
g50974 not n30306 ; n30306_not
g50975 not n17112 ; n17112_not
g50976 not n13026 ; n13026_not
g50977 not n25113 ; n25113_not
g50978 not n13044 ; n13044_not
g50979 not n13053 ; n13053_not
g50980 not n21171 ; n21171_not
g50981 not n34014 ; n34014_not
g50982 not n10074 ; n10074_not
g50983 not n41403 ; n41403_not
g50984 not n19101 ; n19101_not
g50985 not n40413 ; n40413_not
g50986 not n31134 ; n31134_not
g50987 not n10911 ; n10911_not
g50988 not n37200 ; n37200_not
g50989 not n13116 ; n13116_not
g50990 not n34140 ; n34140_not
g50991 not n35301 ; n35301_not
g50992 not n30522 ; n30522_not
g50993 not n21333 ; n21333_not
g50994 not n14250 ; n14250_not
g50995 not n12801 ; n12801_not
g50996 not n34113 ; n34113_not
g50997 not n32511 ; n32511_not
g50998 not n44040 ; n44040_not
g50999 not n25041 ; n25041_not
g51000 not n20271 ; n20271_not
g51001 not n10461 ; n10461_not
g51002 not n25050 ; n25050_not
g51003 not n34104 ; n34104_not
g51004 not n14223 ; n14223_not
g51005 not n20361 ; n20361_not
g51006 not n43140 ; n43140_not
g51007 not n20352 ; n20352_not
g51008 not n26211 ; n26211_not
g51009 not n10371 ; n10371_not
g51010 not n15051 ; n15051_not
g51011 not n41340 ; n41340_not
g51012 not n21108 ; n21108_not
g51013 not n25023 ; n25023_not
g51014 not n22332 ; n22332_not
g51015 not n31143 ; n31143_not
g51016 not n20316 ; n20316_not
g51017 not n30531 ; n30531_not
g51018 not n40620 ; n40620_not
g51019 not n25032 ; n25032_not
g51020 not n20307 ; n20307_not
g51021 not n31431 ; n31431_not
g51022 not n26103 ; n26103_not
g51023 not n22413 ; n22413_not
g51024 not n14160 ; n14160_not
g51025 not n41412 ; n41412_not
g51026 not n20181 ; n20181_not
g51027 not n27111 ; n27111_not
g51028 not n34050 ; n34050_not
g51029 not n20172 ; n20172_not
g51030 not n30360 ; n30360_not
g51031 not n30351 ; n30351_not
g51032 not n14133 ; n14133_not
g51033 not n20163 ; n20163_not
g51034 not n10740 ; n10740_not
g51035 not n15105 ; n15105_not
g51036 not n20244 ; n20244_not
g51037 not n31305 ; n31305_not
g51038 not n45300 ; n45300_not
g51039 not n31152 ; n31152_not
g51040 not n10290 ; n10290_not
g51041 not n30432 ; n30432_not
g51042 not n30423 ; n30423_not
g51043 not n31161 ; n31161_not
g51044 not n33411 ; n33411_not
g51045 not n35310 ; n35310_not
g51046 not n40521 ; n40521_not
g51047 not n21135 ; n21135_not
g51048 not n40512 ; n40512_not
g51049 not n23700 ; n23700_not
g51050 not n32205 ; n32205_not
g51051 not n17301 ; n17301_not
g51052 not n21225 ; n21225_not
g51053 not n23052 ; n23052_not
g51054 not n31251 ; n31251_not
g51055 not n40242 ; n40242_not
g51056 not n13503 ; n13503_not
g51057 not n44400 ; n44400_not
g51058 not n23115 ; n23115_not
g51059 not n40233 ; n40233_not
g51060 not n10524 ; n10524_not
g51061 not n28101 ; n28101_not
g51062 not n16104 ; n16104_not
g51063 not n11712 ; n11712_not
g51064 not n23250 ; n23250_not
g51065 not n32061 ; n32061_not
g51066 not n40215 ; n40215_not
g51067 not n10209 ; n10209_not
g51068 not n11640 ; n11640_not
g51069 not n13422 ; n13422_not
g51070 not n32232 ; n32232_not
g51071 not n23331 ; n23331_not
g51072 not n23322 ; n23322_not
g51073 not n32223 ; n32223_not
g51074 not n30072 ; n30072_not
g51075 not n23232 ; n23232_not
g51076 not n28002 ; n28002_not
g51077 not n41610 ; n41610_not
g51078 not n25302 ; n25302_not
g51079 not n23061 ; n23061_not
g51080 not n30063 ; n30063_not
g51081 not n23070 ; n23070_not
g51082 not n31242 ; n31242_not
g51083 not n43320 ; n43320_not
g51084 not n23304 ; n23304_not
g51085 not n40071 ; n40071_not
g51086 not n25401 ; n25401_not
g51087 not n44112 ; n44112_not
g51088 not n15411 ; n15411_not
g51089 not n32142 ; n32142_not
g51090 not n43401 ; n43401_not
g51091 not n25500 ; n25500_not
g51092 not n36012 ; n36012_not
g51093 not n13710 ; n13710_not
g51094 not n32034 ; n32034_not
g51095 not n40161 ; n40161_not
g51096 not n23160 ; n23160_not
g51097 not n36021 ; n36021_not
g51098 not n32115 ; n32115_not
g51099 not n44211 ; n44211_not
g51100 not n23205 ; n23205_not
g51101 not n32106 ; n32106_not
g51102 not n25410 ; n25410_not
g51103 not n32070 ; n32070_not
g51104 not n40017 ; n40017_not
g51105 not n30018 ; n30018_not
g51106 not n13512 ; n13512_not
g51107 not n27003 ; n27003_not
g51108 not n30009 ; n30009_not
g51109 not n10425 ; n10425_not
g51110 not n23133 ; n23133_not
g51111 not n40044 ; n40044_not
g51112 not n41700 ; n41700_not
g51113 not n28200 ; n28200_not
g51114 not n40053 ; n40053_not
g51115 not n23142 ; n23142_not
g51116 not n23151 ; n23151_not
g51117 not n23223 ; n23223_not
g51118 not n15420 ; n15420_not
g51119 not n10605 ; n10605_not
g51120 not n43203 ; n43203_not
g51121 not n15222 ; n15222_not
g51122 not n23502 ; n23502_not
g51123 not n13251 ; n13251_not
g51124 not n42150 ; n42150_not
g51125 not n20019 ; n20019_not
g51126 not n41520 ; n41520_not
g51127 not n15231 ; n15231_not
g51128 not n25203 ; n25203_not
g51129 not n30234 ; n30234_not
g51130 not n19200 ; n19200_not
g51131 not n43221 ; n43221_not
g51132 not n30225 ; n30225_not
g51133 not n15240 ; n15240_not
g51134 not n30153 ; n30153_not
g51135 not n23430 ; n23430_not
g51136 not n13170 ; n13170_not
g51137 not n26022 ; n26022_not
g51138 not n41502 ; n41502_not
g51139 not n20046 ; n20046_not
g51140 not n27201 ; n27201_not
g51141 not n15204 ; n15204_not
g51142 not n10803 ; n10803_not
g51143 not n23520 ; n23520_not
g51144 not n11802 ; n11802_not
g51145 not n14016 ; n14016_not
g51146 not n20037 ; n20037_not
g51147 not n10272 ; n10272_not
g51148 not n11613 ; n11613_not
g51149 not n13224 ; n13224_not
g51150 not n16140 ; n16140_not
g51151 not n44220 ; n44220_not
g51152 not n13233 ; n13233_not
g51153 not n22521 ; n22521_not
g51154 not n32403 ; n32403_not
g51155 not n31107 ; n31107_not
g51156 not n15510 ; n15510_not
g51157 not n40305 ; n40305_not
g51158 not n13341 ; n13341_not
g51159 not n28011 ; n28011_not
g51160 not n30135 ; n30135_not
g51161 not n21612 ; n21612_not
g51162 not n33510 ; n33510_not
g51163 not n25230 ; n25230_not
g51164 not n44121 ; n44121_not
g51165 not n15501 ; n15501_not
g51166 not n11604 ; n11604_not
g51167 not n10830 ; n10830_not
g51168 not n23340 ; n23340_not
g51169 not n10821 ; n10821_not
g51170 not n40350 ; n40350_not
g51171 not n11622 ; n11622_not
g51172 not n31611 ; n31611_not
g51173 not n32340 ; n32340_not
g51174 not n21018 ; n21018_not
g51175 not n10902 ; n10902_not
g51176 not n11361 ; n11361_not
g51177 not n30162 ; n30162_not
g51178 not n40332 ; n40332_not
g51179 not n13323 ; n13323_not
g51180 not n25221 ; n25221_not
g51181 not n15042 ; n15042_not
g51182 not n40206 ; n40206_not
g51183 not n13332 ; n13332_not
g51184 not n43230 ; n43230_not
g51185 not n32304 ; n32304_not
g51186 not n30144 ; n30144_not
g51187 not n34302 ; n34302_not
g51188 not n12306 ; n12306_not
g51189 not n41232 ; n41232_not
g51190 not n24321 ; n24321_not
g51191 not n33231 ; n33231_not
g51192 not n12324 ; n12324_not
g51193 not n33222 ; n33222_not
g51194 not n34311 ; n34311_not
g51195 not n21045 ; n21045_not
g51196 not n29100 ; n29100_not
g51197 not n33240 ; n33240_not
g51198 not n12351 ; n12351_not
g51199 not n10614 ; n10614_not
g51200 not n22071 ; n22071_not
g51201 not n42312 ; n42312_not
g51202 not n42141 ; n42141_not
g51203 not n12252 ; n12252_not
g51204 not n10533 ; n10533_not
g51205 not n10335 ; n10335_not
g51206 not n38001 ; n38001_not
g51207 not n34320 ; n34320_not
g51208 not n22008 ; n22008_not
g51209 not n18111 ; n18111_not
g51210 not n20730 ; n20730_not
g51211 not n21423 ; n21423_not
g51212 not n41007 ; n41007_not
g51213 not n33213 ; n33213_not
g51214 not n22017 ; n22017_not
g51215 not n21414 ; n21414_not
g51216 not n14502 ; n14502_not
g51217 not n22107 ; n22107_not
g51218 not n31620 ; n31620_not
g51219 not n43104 ; n43104_not
g51220 not n21054 ; n21054_not
g51221 not n31332 ; n31332_not
g51222 not n32700 ; n32700_not
g51223 not n42114 ; n42114_not
g51224 not n11190 ; n11190_not
g51225 not n24141 ; n24141_not
g51226 not n24132 ; n24132_not
g51227 not n10623 ; n10623_not
g51228 not n24006 ; n24006_not
g51229 not n35211 ; n35211_not
g51230 not n24123 ; n24123_not
g51231 not n22152 ; n22152_not
g51232 not n21009 ; n21009_not
g51233 not n24114 ; n24114_not
g51234 not n24231 ; n24231_not
g51235 not n14520 ; n14520_not
g51236 not n14511 ; n14511_not
g51237 not n30810 ; n30810_not
g51238 not n11082 ; n11082_not
g51239 not n46101 ; n46101_not
g51240 not n18003 ; n18003_not
g51241 not n12405 ; n12405_not
g51242 not n30801 ; n30801_not
g51243 not n31080 ; n31080_not
g51244 not n44013 ; n44013_not
g51245 not n35022 ; n35022_not
g51246 not n31602 ; n31602_not
g51247 not n33303 ; n33303_not
g51248 not n42321 ; n42321_not
g51249 not n16401 ; n16401_not
g51250 not n41142 ; n41142_not
g51251 not n42240 ; n42240_not
g51252 not n31008 ; n31008_not
g51253 not n12036 ; n12036_not
g51254 not n12117 ; n12117_not
g51255 not n46020 ; n46020_not
g51256 not n11172 ; n11172_not
g51257 not n11163 ; n11163_not
g51258 not n24510 ; n24510_not
g51259 not n42105 ; n42105_not
g51260 not n31350 ; n31350_not
g51261 not n18201 ; n18201_not
g51262 not n33114 ; n33114_not
g51263 not n41151 ; n41151_not
g51264 not n33105 ; n33105_not
g51265 not n43014 ; n43014_not
g51266 not n12045 ; n12045_not
g51267 not n21801 ; n21801_not
g51268 not n18300 ; n18300_not
g51269 not n31017 ; n31017_not
g51270 not n12072 ; n12072_not
g51271 not n21810 ; n21810_not
g51272 not n35040 ; n35040_not
g51273 not n12090 ; n12090_not
g51274 not n16410 ; n16410_not
g51275 not n20910 ; n20910_not
g51276 not n33141 ; n33141_not
g51277 not n41016 ; n41016_not
g51278 not n41070 ; n41070_not
g51279 not n11154 ; n11154_not
g51280 not n12207 ; n12207_not
g51281 not n43050 ; n43050_not
g51282 not n41061 ; n41061_not
g51283 not n27030 ; n27030_not
g51284 not n41052 ; n41052_not
g51285 not n11118 ; n11118_not
g51286 not n16005 ; n16005_not
g51287 not n12234 ; n12234_not
g51288 not n35130 ; n35130_not
g51289 not n20721 ; n20721_not
g51290 not n11127 ; n11127_not
g51291 not n12135 ; n12135_not
g51292 not n41115 ; n41115_not
g51293 not n33033 ; n33033_not
g51294 not n12153 ; n12153_not
g51295 not n12162 ; n12162_not
g51296 not n11235 ; n11235_not
g51297 not n10317 ; n10317_not
g51298 not n35121 ; n35121_not
g51299 not n16500 ; n16500_not
g51300 not n12018 ; n12018_not
g51301 not n10362 ; n10362_not
g51302 not n33330 ; n33330_not
g51303 not n30621 ; n30621_not
g51304 not n22224 ; n22224_not
g51305 not n41304 ; n41304_not
g51306 not n12180 ; n12180_not
g51307 not n30405 ; n30405_not
g51308 not n24051 ; n24051_not
g51309 not n10650 ; n10650_not
g51310 not n24060 ; n24060_not
g51311 not n46200 ; n46200_not
g51312 not n42006 ; n42006_not
g51313 not n20514 ; n20514_not
g51314 not n10470 ; n10470_not
g51315 not n14403 ; n14403_not
g51316 not n34230 ; n34230_not
g51317 not n31125 ; n31125_not
g51318 not n12540 ; n12540_not
g51319 not n30612 ; n30612_not
g51320 not n12702 ; n12702_not
g51321 not n15033 ; n15033_not
g51322 not n22305 ; n22305_not
g51323 not n11523 ; n11523_not
g51324 not n43131 ; n43131_not
g51325 not n15015 ; n15015_not
g51326 not n42420 ; n42420_not
g51327 not n41322 ; n41322_not
g51328 not n11019 ; n11019_not
g51329 not n26301 ; n26301_not
g51330 not n20451 ; n20451_not
g51331 not n40125 ; n40125_not
g51332 not n15006 ; n15006_not
g51333 not n10704 ; n10704_not
g51334 not n11028 ; n11028_not
g51335 not n31116 ; n31116_not
g51336 not n22260 ; n22260_not
g51337 not n20460 ; n20460_not
g51338 not n41313 ; n41313_not
g51339 not n22242 ; n22242_not
g51340 not n40701 ; n40701_not
g51341 not n47100 ; n47100_not
g51342 not n30630 ; n30630_not
g51343 not n24015 ; n24015_not
g51344 not n27102 ; n27102_not
g51345 not n11262 ; n11262_not
g51346 not n20406 ; n20406_not
g51347 not n14304 ; n14304_not
g51348 not n35004 ; n35004_not
g51349 not n26400 ; n26400_not
g51350 not n12720 ; n12720_not
g51351 not n11514 ; n11514_not
g51352 not n12711 ; n12711_not
g51353 not n12513 ; n12513_not
g51354 not n20550 ; n20550_not
g51355 not n37020 ; n37020_not
g51356 not n14421 ; n14421_not
g51357 not n10506 ; n10506_not
g51358 not n30711 ; n30711_not
g51359 not n11037 ; n11037_not
g51360 not n23305 ; n23305_not
g51361 not n41080 ; n41080_not
g51362 not n23206 ; n23206_not
g51363 not n31405 ; n31405_not
g51364 not n17050 ; n17050_not
g51365 not n37003 ; n37003_not
g51366 not n40234 ; n40234_not
g51367 not n14233 ; n14233_not
g51368 not n43060 ; n43060_not
g51369 not n13801 ; n13801_not
g51370 not n43051 ; n43051_not
g51371 not n36031 ; n36031_not
g51372 not n32224 ; n32224_not
g51373 not n14332 ; n14332_not
g51374 not n41008 ; n41008_not
g51375 not n25042 ; n25042_not
g51376 not n43321 ; n43321_not
g51377 not n27121 ; n27121_not
g51378 not n32125 ; n32125_not
g51379 not n32512 ; n32512_not
g51380 not n11434 ; n11434_not
g51381 not n33133 ; n33133_not
g51382 not n24502 ; n24502_not
g51383 not n21433 ; n21433_not
g51384 not n10318 ; n10318_not
g51385 not n33601 ; n33601_not
g51386 not n21262 ; n21262_not
g51387 not n33403 ; n33403_not
g51388 not n23350 ; n23350_not
g51389 not n32260 ; n32260_not
g51390 not n32251 ; n32251_not
g51391 not n23161 ; n23161_not
g51392 not n13720 ; n13720_not
g51393 not n18400 ; n18400_not
g51394 not n10606 ; n10606_not
g51395 not n15232 ; n15232_not
g51396 not n42511 ; n42511_not
g51397 not n23341 ; n23341_not
g51398 not n36103 ; n36103_not
g51399 not n32242 ; n32242_not
g51400 not n41602 ; n41602_not
g51401 not n21451 ; n21451_not
g51402 not n37012 ; n37012_not
g51403 not n10732 ; n10732_not
g51404 not n10651 ; n10651_not
g51405 not n40531 ; n40531_not
g51406 not n40144 ; n40144_not
g51407 not n43303 ; n43303_not
g51408 not n16231 ; n16231_not
g51409 not n32107 ; n32107_not
g51410 not n23314 ; n23314_not
g51411 not n13810 ; n13810_not
g51412 not n31360 ; n31360_not
g51413 not n41332 ; n41332_not
g51414 not n21370 ; n21370_not
g51415 not n10237 ; n10237_not
g51416 not n42700 ; n42700_not
g51417 not n13702 ; n13702_not
g51418 not n15052 ; n15052_not
g51419 not n18130 ; n18130_not
g51420 not n14323 ; n14323_not
g51421 not n18310 ; n18310_not
g51422 not n16123 ; n16123_not
g51423 not n32170 ; n32170_not
g51424 not n10309 ; n10309_not
g51425 not n41116 ; n41116_not
g51426 not n25015 ; n25015_not
g51427 not n25312 ; n25312_not
g51428 not n23242 ; n23242_not
g51429 not n32161 ; n32161_not
g51430 not n40612 ; n40612_not
g51431 not n33052 ; n33052_not
g51432 not n21271 ; n21271_not
g51433 not n15061 ; n15061_not
g51434 not n14710 ; n14710_not
g51435 not n32152 ; n32152_not
g51436 not n21442 ; n21442_not
g51437 not n15322 ; n15322_not
g51438 not n41044 ; n41044_not
g51439 not n15043 ; n15043_not
g51440 not n23233 ; n23233_not
g51441 not n10417 ; n10417_not
g51442 not n17122 ; n17122_not
g51443 not n40405 ; n40405_not
g51444 not n47011 ; n47011_not
g51445 not n18220 ; n18220_not
g51446 not n31261 ; n31261_not
g51447 not n14242 ; n14242_not
g51448 not n33007 ; n33007_not
g51449 not n40243 ; n40243_not
g51450 not n41143 ; n41143_not
g51451 not n32215 ; n32215_not
g51452 not n25033 ; n25033_not
g51453 not n16132 ; n16132_not
g51454 not n11632 ; n11632_not
g51455 not n25402 ; n25402_not
g51456 not n47110 ; n47110_not
g51457 not n16213 ; n16213_not
g51458 not n21361 ; n21361_not
g51459 not n14260 ; n14260_not
g51460 not n24610 ; n24610_not
g51461 not n21280 ; n21280_not
g51462 not n18301 ; n18301_not
g51463 not n41350 ; n41350_not
g51464 not n18211 ; n18211_not
g51465 not n10219 ; n10219_not
g51466 not n24511 ; n24511_not
g51467 not n40225 ; n40225_not
g51468 not n25006 ; n25006_not
g51469 not n41620 ; n41620_not
g51470 not n21460 ; n21460_not
g51471 not n27022 ; n27022_not
g51472 not n17032 ; n17032_not
g51473 not n19120 ; n19120_not
g51474 not n14503 ; n14503_not
g51475 not n25150 ; n25150_not
g51476 not n32422 ; n32422_not
g51477 not n19003 ; n19003_not
g51478 not n41251 ; n41251_not
g51479 not n41026 ; n41026_not
g51480 not n21505 ; n21505_not
g51481 not n14035 ; n14035_not
g51482 not n31414 ; n31414_not
g51483 not n40450 ; n40450_not
g51484 not n41422 ; n41422_not
g51485 not n33331 ; n33331_not
g51486 not n32314 ; n32314_not
g51487 not n10822 ; n10822_not
g51488 not n24205 ; n24205_not
g51489 not n20902 ; n20902_not
g51490 not n16222 ; n16222_not
g51491 not n24232 ; n24232_not
g51492 not n32413 ; n32413_not
g51493 not n10714 ; n10714_not
g51494 not n25123 ; n25123_not
g51495 not n24223 ; n24223_not
g51496 not n41224 ; n41224_not
g51497 not n41512 ; n41512_not
g51498 not n10381 ; n10381_not
g51499 not n18013 ; n18013_not
g51500 not n10750 ; n10750_not
g51501 not n31270 ; n31270_not
g51502 not n14404 ; n14404_not
g51503 not n24070 ; n24070_not
g51504 not n21316 ; n21316_not
g51505 not n40810 ; n40810_not
g51506 not n14107 ; n14107_not
g51507 not n21541 ; n21541_not
g51508 not n40432 ; n40432_not
g51509 not n40333 ; n40333_not
g51510 not n33421 ; n33421_not
g51511 not n33322 ; n33322_not
g51512 not n23602 ; n23602_not
g51513 not n15160 ; n15160_not
g51514 not n14116 ; n14116_not
g51515 not n43114 ; n43114_not
g51516 not n36211 ; n36211_not
g51517 not n36202 ; n36202_not
g51518 not n25105 ; n25105_not
g51519 not n24151 ; n24151_not
g51520 not n14134 ; n14134_not
g51521 not n33304 ; n33304_not
g51522 not n19111 ; n19111_not
g51523 not n44410 ; n44410_not
g51524 not n10570 ; n10570_not
g51525 not n43123 ; n43123_not
g51526 not n42430 ; n42430_not
g51527 not n14071 ; n14071_not
g51528 not n14062 ; n14062_not
g51529 not n40414 ; n40414_not
g51530 not n48001 ; n48001_not
g51531 not n14080 ; n14080_not
g51532 not n32440 ; n32440_not
g51533 not n40342 ; n40342_not
g51534 not n40423 ; n40423_not
g51535 not n32611 ; n32611_not
g51536 not n14206 ; n14206_not
g51537 not n15007 ; n15007_not
g51538 not n40324 ; n40324_not
g51539 not n18112 ; n18112_not
g51540 not n11470 ; n11470_not
g51541 not n11623 ; n11623_not
g51542 not n41035 ; n41035_not
g51543 not n16204 ; n16204_not
g51544 not n25222 ; n25222_not
g51545 not n31306 ; n31306_not
g51546 not n32332 ; n32332_not
g51547 not n23404 ; n23404_not
g51548 not n21550 ; n21550_not
g51549 not n48010 ; n48010_not
g51550 not n11524 ; n11524_not
g51551 not n33205 ; n33205_not
g51552 not n40306 ; n40306_not
g51553 not n21343 ; n21343_not
g51554 not n40702 ; n40702_not
g51555 not n33520 ; n33520_not
g51556 not n24430 ; n24430_not
g51557 not n21352 ; n21352_not
g51558 not n29020 ; n29020_not
g51559 not n14215 ; n14215_not
g51560 not n19300 ; n19300_not
g51561 not n10741 ; n10741_not
g51562 not n25231 ; n25231_not
g51563 not n41314 ; n41314_not
g51564 not n24322 ; n24322_not
g51565 not n41233 ; n41233_not
g51566 not n24034 ; n24034_not
g51567 not n10390 ; n10390_not
g51568 not n41260 ; n41260_not
g51569 not n21334 ; n21334_not
g51570 not n33232 ; n33232_not
g51571 not n36301 ; n36301_not
g51572 not n15214 ; n15214_not
g51573 not n40207 ; n40207_not
g51574 not n33241 ; n33241_not
g51575 not n41242 ; n41242_not
g51576 not n23503 ; n23503_not
g51577 not n23512 ; n23512_not
g51578 not n24241 ; n24241_not
g51579 not n10273 ; n10273_not
g51580 not n18022 ; n18022_not
g51581 not n36121 ; n36121_not
g51582 not n15250 ; n15250_not
g51583 not n14611 ; n14611_not
g51584 not n40522 ; n40522_not
g51585 not n32620 ; n32620_not
g51586 not n40540 ; n40540_not
g51587 not n23413 ; n23413_not
g51588 not n15115 ; n15115_not
g51589 not n32350 ; n32350_not
g51590 not n33214 ; n33214_not
g51591 not n43240 ; n43240_not
g51592 not n24007 ; n24007_not
g51593 not n24340 ; n24340_not
g51594 not n25204 ; n25204_not
g51595 not n43231 ; n43231_not
g51596 not n33223 ; n33223_not
g51597 not n34501 ; n34501_not
g51598 not n40360 ; n40360_not
g51599 not n10633 ; n10633_not
g51600 not n20380 ; n20380_not
g51601 not n20371 ; n20371_not
g51602 not n20362 ; n20362_not
g51603 not n11911 ; n11911_not
g51604 not n20344 ; n20344_not
g51605 not n42124 ; n42124_not
g51606 not n22333 ; n22333_not
g51607 not n20254 ; n20254_not
g51608 not n26122 ; n26122_not
g51609 not n26203 ; n26203_not
g51610 not n11290 ; n11290_not
g51611 not n20326 ; n20326_not
g51612 not n22324 ; n22324_not
g51613 not n30451 ; n30451_not
g51614 not n22342 ; n22342_not
g51615 not n46210 ; n46210_not
g51616 not n22351 ; n22351_not
g51617 not n21091 ; n21091_not
g51618 not n12811 ; n12811_not
g51619 not n31144 ; n31144_not
g51620 not n20281 ; n20281_not
g51621 not n34114 ; n34114_not
g51622 not n40315 ; n40315_not
g51623 not n30712 ; n30712_not
g51624 not n20506 ; n20506_not
g51625 not n34213 ; n34213_not
g51626 not n41800 ; n41800_not
g51627 not n22234 ; n22234_not
g51628 not n20416 ; n20416_not
g51629 not n22261 ; n22261_not
g51630 not n12316 ; n12316_not
g51631 not n16015 ; n16015_not
g51632 not n11263 ; n11263_not
g51633 not n26311 ; n26311_not
g51634 not n10615 ; n10615_not
g51635 not n34204 ; n34204_not
g51636 not n22270 ; n22270_not
g51637 not n12631 ; n12631_not
g51638 not n12604 ; n12604_not
g51639 not n21073 ; n21073_not
g51640 not n31108 ; n31108_not
g51641 not n20425 ; n20425_not
g51642 not n22252 ; n22252_not
g51643 not n20407 ; n20407_not
g51644 not n12181 ; n12181_not
g51645 not n12703 ; n12703_not
g51646 not n34042 ; n34042_not
g51647 not n20146 ; n20146_not
g51648 not n21136 ; n21136_not
g51649 not n11308 ; n11308_not
g51650 not n42142 ; n42142_not
g51651 not n31423 ; n31423_not
g51652 not n15601 ; n15601_not
g51653 not n44230 ; n44230_not
g51654 not n42502 ; n42502_not
g51655 not n21163 ; n21163_not
g51656 not n30208 ; n30208_not
g51657 not n16051 ; n16051_not
g51658 not n13054 ; n13054_not
g51659 not n45211 ; n45211_not
g51660 not n10453 ; n10453_not
g51661 not n30280 ; n30280_not
g51662 not n20092 ; n20092_not
g51663 not n11821 ; n11821_not
g51664 not n30190 ; n30190_not
g51665 not n11812 ; n11812_not
g51666 not n27211 ; n27211_not
g51667 not n16024 ; n16024_not
g51668 not n31702 ; n31702_not
g51669 not n35302 ; n35302_not
g51670 not n20263 ; n20263_not
g51671 not n42133 ; n42133_not
g51672 not n34105 ; n34105_not
g51673 not n30460 ; n30460_not
g51674 not n20245 ; n20245_not
g51675 not n30406 ; n30406_not
g51676 not n31153 ; n31153_not
g51677 not n30433 ; n30433_not
g51678 not n16042 ; n16042_not
g51679 not n12901 ; n12901_not
g51680 not n44050 ; n44050_not
g51681 not n12910 ; n12910_not
g51682 not n31711 ; n31711_not
g51683 not n10642 ; n10642_not
g51684 not n34060 ; n34060_not
g51685 not n39010 ; n39010_not
g51686 not n22423 ; n22423_not
g51687 not n31171 ; n31171_not
g51688 not n30361 ; n30361_not
g51689 not n22432 ; n22432_not
g51690 not n21145 ; n21145_not
g51691 not n31432 ; n31432_not
g51692 not n16501 ; n16501_not
g51693 not n12190 ; n12190_not
g51694 not n20821 ; n20821_not
g51695 not n20812 ; n20812_not
g51696 not n20803 ; n20803_not
g51697 not n12217 ; n12217_not
g51698 not n20713 ; n20713_not
g51699 not n11146 ; n11146_not
g51700 not n11137 ; n11137_not
g51701 not n31063 ; n31063_not
g51702 not n12226 ; n12226_not
g51703 not n16510 ; n16510_not
g51704 not n12244 ; n12244_not
g51705 not n26320 ; n26320_not
g51706 not n34321 ; n34321_not
g51707 not n22009 ; n22009_not
g51708 not n12271 ; n12271_not
g51709 not n41404 ; n41404_not
g51710 not n12280 ; n12280_not
g51711 not n11119 ; n11119_not
g51712 not n20722 ; n20722_not
g51713 not n22018 ; n22018_not
g51714 not n42205 ; n42205_not
g51715 not n35023 ; n35023_not
g51716 not n46003 ; n46003_not
g51717 not n38110 ; n38110_not
g51718 not n42223 ; n42223_not
g51719 not n12073 ; n12073_not
g51720 not n35032 ; n35032_not
g51721 not n12082 ; n12082_not
g51722 not n31018 ; n31018_not
g51723 not n31009 ; n31009_not
g51724 not n12109 ; n12109_not
g51725 not n42241 ; n42241_not
g51726 not n38101 ; n38101_not
g51727 not n46030 ; n46030_not
g51728 not n42106 ; n42106_not
g51729 not n12136 ; n12136_not
g51730 not n17041 ; n17041_not
g51731 not n35104 ; n35104_not
g51732 not n10534 ; n10534_not
g51733 not n21910 ; n21910_not
g51734 not n12172 ; n12172_not
g51735 not n20830 ; n20830_not
g51736 not n10525 ; n10525_not
g51737 not n20623 ; n20623_not
g51738 not n20434 ; n20434_not
g51739 not n12424 ; n12424_not
g51740 not n20614 ; n20614_not
g51741 not n12442 ; n12442_not
g51742 not n46111 ; n46111_not
g51743 not n20605 ; n20605_not
g51744 not n31621 ; n31621_not
g51745 not n31081 ; n31081_not
g51746 not n22144 ; n22144_not
g51747 not n31630 ; n31630_not
g51748 not n30730 ; n30730_not
g51749 not n20560 ; n20560_not
g51750 not n42016 ; n42016_not
g51751 not n22171 ; n22171_not
g51752 not n44302 ; n44302_not
g51753 not n11038 ; n11038_not
g51754 not n35212 ; n35212_not
g51755 not n12523 ; n12523_not
g51756 not n11047 ; n11047_not
g51757 not n21712 ; n21712_not
g51758 not n12550 ; n12550_not
g51759 not n31090 ; n31090_not
g51760 not n30901 ; n30901_not
g51761 not n31540 ; n31540_not
g51762 not n34312 ; n34312_not
g51763 not n12307 ; n12307_not
g51764 not n22027 ; n22027_not
g51765 not n22036 ; n22036_not
g51766 not n11245 ; n11245_not
g51767 not n16006 ; n16006_not
g51768 not n12334 ; n12334_not
g51769 not n21028 ; n21028_not
g51770 not n22054 ; n22054_not
g51771 not n27400 ; n27400_not
g51772 not n22063 ; n22063_not
g51773 not n42304 ; n42304_not
g51774 not n31072 ; n31072_not
g51775 not n21721 ; n21721_not
g51776 not n12361 ; n12361_not
g51777 not n20443 ; n20443_not
g51778 not n12370 ; n12370_not
g51779 not n16402 ; n16402_not
g51780 not n30820 ; n30820_not
g51781 not n35203 ; n35203_not
g51782 not n22090 ; n22090_not
g51783 not n20641 ; n20641_not
g51784 not n42232 ; n42232_not
g51785 not n20632 ; n20632_not
g51786 not n13360 ; n13360_not
g51787 not n16060 ; n16060_not
g51788 not n21217 ; n21217_not
g51789 not n22711 ; n22711_not
g51790 not n22702 ; n22702_not
g51791 not n22720 ; n22720_not
g51792 not n43501 ; n43501_not
g51793 not n28021 ; n28021_not
g51794 not n30091 ; n30091_not
g51795 not n22801 ; n22801_not
g51796 not n22810 ; n22810_not
g51797 not n30082 ; n30082_not
g51798 not n10426 ; n10426_not
g51799 not n13414 ; n13414_not
g51800 not n34402 ; n34402_not
g51801 not n23008 ; n23008_not
g51802 not n31234 ; n31234_not
g51803 not n13450 ; n13450_not
g51804 not n23044 ; n23044_not
g51805 not n30073 ; n30073_not
g51806 not n22540 ; n22540_not
g51807 not n31216 ; n31216_not
g51808 not n10903 ; n10903_not
g51809 not n33700 ; n33700_not
g51810 not n13315 ; n13315_not
g51811 not n15520 ; n15520_not
g51812 not n28003 ; n28003_not
g51813 not n22612 ; n22612_not
g51814 not n31225 ; n31225_not
g51815 not n42160 ; n42160_not
g51816 not n22630 ; n22630_not
g51817 not n22621 ; n22621_not
g51818 not n13342 ; n13342_not
g51819 not n13351 ; n13351_not
g51820 not n15511 ; n15511_not
g51821 not n40045 ; n40045_not
g51822 not n15421 ; n15421_not
g51823 not n23152 ; n23152_not
g51824 not n11704 ; n11704_not
g51825 not n32017 ; n32017_not
g51826 not n43402 ; n43402_not
g51827 not n15403 ; n15403_not
g51828 not n32026 ; n32026_not
g51829 not n40090 ; n40090_not
g51830 not n13612 ; n13612_not
g51831 not n45121 ; n45121_not
g51832 not n16105 ; n16105_not
g51833 not n13621 ; n13621_not
g51834 not n44104 ; n44104_not
g51835 not n32035 ; n32035_not
g51836 not n32044 ; n32044_not
g51837 not n13630 ; n13630_not
g51838 not n42520 ; n42520_not
g51839 not n10183 ; n10183_not
g51840 not n32062 ; n32062_not
g51841 not n42601 ; n42601_not
g51842 not n45112 ; n45112_not
g51843 not n10192 ; n10192_not
g51844 not n40126 ; n40126_not
g51845 not n23053 ; n23053_not
g51846 not n23062 ; n23062_not
g51847 not n37300 ; n37300_not
g51848 not n47200 ; n47200_not
g51849 not n30046 ; n30046_not
g51850 not n30028 ; n30028_not
g51851 not n28102 ; n28102_not
g51852 not n17113 ; n17113_not
g51853 not n13504 ; n13504_not
g51854 not n40009 ; n40009_not
g51855 not n11713 ; n11713_not
g51856 not n41710 ; n41710_not
g51857 not n13513 ; n13513_not
g51858 not n40018 ; n40018_not
g51859 not n23116 ; n23116_not
g51860 not n30019 ; n30019_not
g51861 not n28120 ; n28120_not
g51862 not n40036 ; n40036_not
g51863 not n31900 ; n31900_not
g51864 not n13261 ; n13261_not
g51865 not n21622 ; n21622_not
g51866 not n13243 ; n13243_not
g51867 not n22504 ; n22504_not
g51868 not n30235 ; n30235_not
g51869 not n21631 ; n21631_not
g51870 not n22522 ; n22522_not
g51871 not n21181 ; n21181_not
g51872 not n10912 ; n10912_not
g51873 not n31207 ; n31207_not
g51874 not n43510 ; n43510_not
g51875 not n10039 ; n10039_not
g51876 not n17230 ; n17230_not
g51877 not n11803 ; n11803_not
g51878 not n46300 ; n46300_not
g51879 not n26014 ; n26014_not
g51880 not n10921 ; n10921_not
g51881 not n10327 ; n10327_not
g51882 not n13225 ; n13225_not
g51883 not n10057 ; n10057_not
g51884 not n22513 ; n22513_not
g51885 not n13234 ; n13234_not
g51886 not n20065 ; n20065_not
g51887 not n30226 ; n30226_not
g51888 not n20056 ; n20056_not
g51889 not n16303 ; n16303_not
g51890 not n13270 ; n13270_not
g51891 not n13216 ; n13216_not
g51892 not n22531 ; n22531_not
g51893 not n42215 ; n42215_not
g51894 not n42080 ; n42080_not
g51895 not n41441 ; n41441_not
g51896 not n41216 ; n41216_not
g51897 not n17060 ; n17060_not
g51898 not n33206 ; n33206_not
g51899 not n25322 ; n25322_not
g51900 not n15332 ; n15332_not
g51901 not n10373 ; n10373_not
g51902 not n25610 ; n25610_not
g51903 not n40145 ; n40145_not
g51904 not n14612 ; n14612_not
g51905 not n34412 ; n34412_not
g51906 not n23081 ; n23081_not
g51907 not n10427 ; n10427_not
g51908 not n17033 ; n17033_not
g51909 not n47210 ; n47210_not
g51910 not n16106 ; n16106_not
g51911 not n34520 ; n34520_not
g51912 not n25115 ; n25115_not
g51913 not n34340 ; n34340_not
g51914 not n33125 ; n33125_not
g51915 not n33800 ; n33800_not
g51916 not n18131 ; n18131_not
g51917 not n27140 ; n27140_not
g51918 not n27131 ; n27131_not
g51919 not n33251 ; n33251_not
g51920 not n34034 ; n34034_not
g51921 not n41243 ; n41243_not
g51922 not n28103 ; n28103_not
g51923 not n18032 ; n18032_not
g51924 not n27410 ; n27410_not
g51925 not n42305 ; n42305_not
g51926 not n26510 ; n26510_not
g51927 not n18041 ; n18041_not
g51928 not n34511 ; n34511_not
g51929 not n27122 ; n27122_not
g51930 not n10391 ; n10391_not
g51931 not n24602 ; n24602_not
g51932 not n33512 ; n33512_not
g51933 not n35150 ; n35150_not
g51934 not n41153 ; n41153_not
g51935 not n17330 ; n17330_not
g51936 not n10607 ; n10607_not
g51937 not n15341 ; n15341_not
g51938 not n34304 ; n34304_not
g51939 not n40514 ; n40514_not
g51940 not n41630 ; n41630_not
g51941 not n36311 ; n36311_not
g51942 not n40235 ; n40235_not
g51943 not n21641 ; n21641_not
g51944 not n10544 ; n10544_not
g51945 not n14810 ; n14810_not
g51946 not n16340 ; n16340_not
g51947 not n10526 ; n10526_not
g51948 not n26024 ; n26024_not
g51949 not n42107 ; n42107_not
g51950 not n18212 ; n18212_not
g51951 not n10571 ; n10571_not
g51952 not n42251 ; n42251_not
g51953 not n36500 ; n36500_not
g51954 not n10562 ; n10562_not
g51955 not n18221 ; n18221_not
g51956 not n34403 ; n34403_not
g51957 not n44501 ; n44501_not
g51958 not n20570 ; n20570_not
g51959 not n16241 ; n16241_not
g51960 not n16412 ; n16412_not
g51961 not n33143 ; n33143_not
g51962 not n18230 ; n18230_not
g51963 not n18104 ; n18104_not
g51964 not n36023 ; n36023_not
g51965 not n17420 ; n17420_not
g51966 not n34421 ; n34421_not
g51967 not n28400 ; n28400_not
g51968 not n16232 ; n16232_not
g51969 not n24620 ; n24620_not
g51970 not n41162 ; n41162_not
g51971 not n16421 ; n16421_not
g51972 not n41207 ; n41207_not
g51973 not n17402 ; n17402_not
g51974 not n28031 ; n28031_not
g51975 not n28130 ; n28130_not
g51976 not n35024 ; n35024_not
g51977 not n15170 ; n15170_not
g51978 not n26051 ; n26051_not
g51979 not n41450 ; n41450_not
g51980 not n16331 ; n16331_not
g51981 not n27005 ; n27005_not
g51982 not n10445 ; n10445_not
g51983 not n17015 ; n17015_not
g51984 not n42206 ; n42206_not
g51985 not n24413 ; n24413_not
g51986 not n42611 ; n42611_not
g51987 not n33161 ; n33161_not
g51988 not n35123 ; n35123_not
g51989 not n41306 ; n41306_not
g51990 not n40181 ; n40181_not
g51991 not n36014 ; n36014_not
g51992 not n24710 ; n24710_not
g51993 not n35114 ; n35114_not
g51994 not n33170 ; n33170_not
g51995 not n14513 ; n14513_not
g51996 not n33620 ; n33620_not
g51997 not n26600 ; n26600_not
g51998 not n26240 ; n26240_not
g51999 not n41333 ; n41333_not
g52000 not n40208 ; n40208_not
g52001 not n28310 ; n28310_not
g52002 not n41405 ; n41405_not
g52003 not n26231 ; n26231_not
g52004 not n42710 ; n42710_not
g52005 not n25061 ; n25061_not
g52006 not n41324 ; n41324_not
g52007 not n27104 ; n27104_not
g52008 not n16016 ; n16016_not
g52009 not n42431 ; n42431_not
g52010 not n10661 ; n10661_not
g52011 not n42530 ; n42530_not
g52012 not n34070 ; n34070_not
g52013 not n10652 ; n10652_not
g52014 not n15017 ; n15017_not
g52015 not n47102 ; n47102_not
g52016 not n33341 ; n33341_not
g52017 not n47120 ; n47120_not
g52018 not n26303 ; n26303_not
g52019 not n40172 ; n40172_not
g52020 not n15503 ; n15503_not
g52021 not n27221 ; n27221_not
g52022 not n42422 ; n42422_not
g52023 not n41513 ; n41513_not
g52024 not n28301 ; n28301_not
g52025 not n15071 ; n15071_not
g52026 not n25214 ; n25214_not
g52027 not n17105 ; n17105_not
g52028 not n33503 ; n33503_not
g52029 not n10463 ; n10463_not
g52030 not n15080 ; n15080_not
g52031 not n42440 ; n42440_not
g52032 not n34124 ; n34124_not
g52033 not n16214 ; n16214_not
g52034 not n34025 ; n34025_not
g52035 not n15242 ; n15242_not
g52036 not n26141 ; n26141_not
g52037 not n41603 ; n41603_not
g52038 not n26150 ; n26150_not
g52039 not n26123 ; n26123_not
g52040 not n10436 ; n10436_not
g52041 not n26213 ; n26213_not
g52042 not n17123 ; n17123_not
g52043 not n15107 ; n15107_not
g52044 not n15053 ; n15053_not
g52045 not n15521 ; n15521_not
g52046 not n27014 ; n27014_not
g52047 not n25016 ; n25016_not
g52048 not n40073 ; n40073_not
g52049 not n34133 ; n34133_not
g52050 not n26132 ; n26132_not
g52051 not n26114 ; n26114_not
g52052 not n42152 ; n42152_not
g52053 not n16133 ; n16133_not
g52054 not n15134 ; n15134_not
g52055 not n33305 ; n33305_not
g52056 not n41252 ; n41252_not
g52057 not n41801 ; n41801_not
g52058 not n16403 ; n16403_not
g52059 not n41810 ; n41810_not
g52060 not n16205 ; n16205_not
g52061 not n41261 ; n41261_not
g52062 not n27320 ; n27320_not
g52063 not n26420 ; n26420_not
g52064 not n17600 ; n17600_not
g52065 not n42350 ; n42350_not
g52066 not n41270 ; n41270_not
g52067 not n33314 ; n33314_not
g52068 not n42062 ; n42062_not
g52069 not n33260 ; n33260_not
g52070 not n18023 ; n18023_not
g52071 not n41360 ; n41360_not
g52072 not n25304 ; n25304_not
g52073 not n16043 ; n16043_not
g52074 not n42053 ; n42053_not
g52075 not n15143 ; n15143_not
g52076 not n15152 ; n15152_not
g52077 not n41720 ; n41720_not
g52078 not n16250 ; n16250_not
g52079 not n41702 ; n41702_not
g52080 not n41423 ; n41423_not
g52081 not n17231 ; n17231_not
g52082 not n26042 ; n26042_not
g52083 not n35222 ; n35222_not
g52084 not n10643 ; n10643_not
g52085 not n35231 ; n35231_not
g52086 not n34223 ; n34223_not
g52087 not n35240 ; n35240_not
g52088 not n33413 ; n33413_not
g52089 not n34061 ; n34061_not
g52090 not n17150 ; n17150_not
g52091 not n25250 ; n25250_not
g52092 not n34214 ; n34214_not
g52093 not n40127 ; n40127_not
g52094 not n42404 ; n42404_not
g52095 not n26006 ; n26006_not
g52096 not n35321 ; n35321_not
g52097 not n42143 ; n42143_not
g52098 not n17213 ; n17213_not
g52099 not n36221 ; n36221_not
g52100 not n42026 ; n42026_not
g52101 not n17204 ; n17204_not
g52102 not n35510 ; n35510_not
g52103 not n35501 ; n35501_not
g52104 not n16160 ; n16160_not
g52105 not n26411 ; n26411_not
g52106 not n33323 ; n33323_not
g52107 not n10490 ; n10490_not
g52108 not n16052 ; n16052_not
g52109 not n42017 ; n42017_not
g52110 not n17312 ; n17312_not
g52111 not n10508 ; n10508_not
g52112 not n34043 ; n34043_not
g52113 not n27041 ; n27041_not
g52114 not n10922 ; n10922_not
g52115 not n30254 ; n30254_not
g52116 not n43502 ; n43502_not
g52117 not n30182 ; n30182_not
g52118 not n13181 ; n13181_not
g52119 not n45203 ; n45203_not
g52120 not n13172 ; n13172_not
g52121 not n30263 ; n30263_not
g52122 not n20075 ; n20075_not
g52123 not n13118 ; n13118_not
g52124 not n10940 ; n10940_not
g52125 not n30272 ; n30272_not
g52126 not n20084 ; n20084_not
g52127 not n22460 ; n22460_not
g52128 not n13055 ; n13055_not
g52129 not n13037 ; n13037_not
g52130 not n22451 ; n22451_not
g52131 not n13352 ; n13352_not
g52132 not n22631 ; n22631_not
g52133 not n30146 ; n30146_not
g52134 not n13325 ; n13325_not
g52135 not n22604 ; n22604_not
g52136 not n10328 ; n10328_not
g52137 not n30191 ; n30191_not
g52138 not n39110 ; n39110_not
g52139 not n30218 ; n30218_not
g52140 not n13262 ; n13262_not
g52141 not n10076 ; n10076_not
g52142 not n13253 ; n13253_not
g52143 not n13244 ; n13244_not
g52144 not n30245 ; n30245_not
g52145 not n13217 ; n13217_not
g52146 not n13235 ; n13235_not
g52147 not n22514 ; n22514_not
g52148 not n31712 ; n31712_not
g52149 not n30452 ; n30452_not
g52150 not n22370 ; n22370_not
g52151 not n30470 ; n30470_not
g52152 not n30425 ; n30425_not
g52153 not n31703 ; n31703_not
g52154 not n12830 ; n12830_not
g52155 not n30506 ; n30506_not
g52156 not n31514 ; n31514_not
g52157 not n30515 ; n30515_not
g52158 not n22352 ; n22352_not
g52159 not n43520 ; n43520_not
g52160 not n30542 ; n30542_not
g52161 not n20336 ; n20336_not
g52162 not n30551 ; n30551_not
g52163 not n20354 ; n20354_not
g52164 not n45221 ; n45221_not
g52165 not n13019 ; n13019_not
g52166 not n30317 ; n30317_not
g52167 not n30335 ; n30335_not
g52168 not n22433 ; n22433_not
g52169 not n30353 ; n30353_not
g52170 not n20165 ; n20165_not
g52171 not n31730 ; n31730_not
g52172 not n31523 ; n31523_not
g52173 not n20174 ; n20174_not
g52174 not n20183 ; n20183_not
g52175 not n31721 ; n31721_not
g52176 not n22415 ; n22415_not
g52177 not n12920 ; n12920_not
g52178 not n22406 ; n22406_not
g52179 not n30416 ; n30416_not
g52180 not n12902 ; n12902_not
g52181 not n32180 ; n32180_not
g52182 not n23243 ; n23243_not
g52183 not n40190 ; n40190_not
g52184 not n32144 ; n32144_not
g52185 not n13721 ; n13721_not
g52186 not n13703 ; n13703_not
g52187 not n32126 ; n32126_not
g52188 not n40154 ; n40154_not
g52189 not n13640 ; n13640_not
g52190 not n23171 ; n23171_not
g52191 not n45113 ; n45113_not
g52192 not n40118 ; n40118_not
g52193 not n13622 ; n13622_not
g52194 not n10823 ; n10823_not
g52195 not n40307 ; n40307_not
g52196 not n32261 ; n32261_not
g52197 not n23351 ; n23351_not
g52198 not n23342 ; n23342_not
g52199 not n23315 ; n23315_not
g52200 not n10238 ; n10238_not
g52201 not n13820 ; n13820_not
g52202 not n40280 ; n40280_not
g52203 not n13811 ; n13811_not
g52204 not n10850 ; n10850_not
g52205 not n43322 ; n43322_not
g52206 not n40262 ; n40262_not
g52207 not n43340 ; n43340_not
g52208 not n32207 ; n32207_not
g52209 not n10229 ; n10229_not
g52210 not n40226 ; n40226_not
g52211 not n43430 ; n43430_not
g52212 not n13460 ; n13460_not
g52213 not n43421 ; n43421_not
g52214 not n13433 ; n13433_not
g52215 not n30065 ; n30065_not
g52216 not n23027 ; n23027_not
g52217 not n23018 ; n23018_not
g52218 not n37400 ; n37400_not
g52219 not n22730 ; n22730_not
g52220 not n22703 ; n22703_not
g52221 not n22712 ; n22712_not
g52222 not n30119 ; n30119_not
g52223 not n22622 ; n22622_not
g52224 not n32036 ; n32036_not
g52225 not n23162 ; n23162_not
g52226 not n40082 ; n40082_not
g52227 not n10535 ; n10535_not
g52228 not n31901 ; n31901_not
g52229 not n40046 ; n40046_not
g52230 not n23126 ; n23126_not
g52231 not n43412 ; n43412_not
g52232 not n13541 ; n13541_not
g52233 not n13532 ; n13532_not
g52234 not n30029 ; n30029_not
g52235 not n13523 ; n13523_not
g52236 not n13514 ; n13514_not
g52237 not n13505 ; n13505_not
g52238 not n30038 ; n30038_not
g52239 not n23108 ; n23108_not
g52240 not n30047 ; n30047_not
g52241 not n31424 ; n31424_not
g52242 not n21092 ; n21092_not
g52243 not n11903 ; n11903_not
g52244 not n44213 ; n44213_not
g52245 not n21119 ; n21119_not
g52246 not n21038 ; n21038_not
g52247 not n21137 ; n21137_not
g52248 not n38201 ; n38201_not
g52249 not n31172 ; n31172_not
g52250 not n31190 ; n31190_not
g52251 not n11309 ; n11309_not
g52252 not n44060 ; n44060_not
g52253 not n21173 ; n21173_not
g52254 not n11813 ; n11813_not
g52255 not n11183 ; n11183_not
g52256 not n11192 ; n11192_not
g52257 not n12092 ; n12092_not
g52258 not n21830 ; n21830_not
g52259 not n20921 ; n20921_not
g52260 not n21821 ; n21821_not
g52261 not n12038 ; n12038_not
g52262 not n12056 ; n12056_not
g52263 not n38102 ; n38102_not
g52264 not n11147 ; n11147_not
g52265 not n11219 ; n11219_not
g52266 not n46004 ; n46004_not
g52267 not n12029 ; n12029_not
g52268 not n21731 ; n21731_not
g52269 not n31442 ; n31442_not
g52270 not n31451 ; n31451_not
g52271 not n31082 ; n31082_not
g52272 not n21542 ; n21542_not
g52273 not n21560 ; n21560_not
g52274 not n11633 ; n11633_not
g52275 not n11624 ; n11624_not
g52276 not n44123 ; n44123_not
g52277 not n21308 ; n21308_not
g52278 not n44204 ; n44204_not
g52279 not n21074 ; n21074_not
g52280 not n31307 ; n31307_not
g52281 not n21515 ; n21515_not
g52282 not n21362 ; n21362_not
g52283 not n11507 ; n11507_not
g52284 not n21506 ; n21506_not
g52285 not n31370 ; n31370_not
g52286 not n21425 ; n21425_not
g52287 not n21452 ; n21452_not
g52288 not n21155 ; n21155_not
g52289 not n21623 ; n21623_not
g52290 not n31037 ; n31037_not
g52291 not n21209 ; n21209_not
g52292 not n31226 ; n31226_not
g52293 not n21614 ; n21614_not
g52294 not n31235 ; n31235_not
g52295 not n11750 ; n11750_not
g52296 not n21605 ; n21605_not
g52297 not n31244 ; n31244_not
g52298 not n31415 ; n31415_not
g52299 not n31046 ; n31046_not
g52300 not n31253 ; n31253_not
g52301 not n44114 ; n44114_not
g52302 not n21254 ; n21254_not
g52303 not n11363 ; n11363_not
g52304 not n30713 ; n30713_not
g52305 not n11039 ; n11039_not
g52306 not n20534 ; n20534_not
g52307 not n30722 ; n30722_not
g52308 not n22181 ; n22181_not
g52309 not n22172 ; n22172_not
g52310 not n22163 ; n22163_not
g52311 not n22145 ; n22145_not
g52312 not n22136 ; n22136_not
g52313 not n12470 ; n12470_not
g52314 not n12452 ; n12452_not
g52315 not n22118 ; n22118_not
g52316 not n12434 ; n12434_not
g52317 not n30803 ; n30803_not
g52318 not n20651 ; n20651_not
g52319 not n30830 ; n30830_not
g52320 not n22325 ; n22325_not
g52321 not n30614 ; n30614_not
g52322 not n20390 ; n20390_not
g52323 not n30623 ; n30623_not
g52324 not n30632 ; n30632_not
g52325 not n12650 ; n12650_not
g52326 not n20435 ; n20435_not
g52327 not n12623 ; n12623_not
g52328 not n12605 ; n12605_not
g52329 not n30650 ; n30650_not
g52330 not n22262 ; n22262_not
g52331 not n12614 ; n12614_not
g52332 not n22244 ; n22244_not
g52333 not n30704 ; n30704_not
g52334 not n20507 ; n20507_not
g52335 not n12560 ; n12560_not
g52336 not n11156 ; n11156_not
g52337 not n20741 ; n20741_not
g52338 not n12182 ; n12182_not
g52339 not n12173 ; n12173_not
g52340 not n12164 ; n12164_not
g52341 not n11912 ; n11912_not
g52342 not n21902 ; n21902_not
g52343 not n12155 ; n12155_not
g52344 not n20831 ; n20831_not
g52345 not n11417 ; n11417_not
g52346 not n12146 ; n12146_not
g52347 not n11165 ; n11165_not
g52348 not n12137 ; n12137_not
g52349 not n12065 ; n12065_not
g52350 not n12128 ; n12128_not
g52351 not n12119 ; n12119_not
g52352 not n20660 ; n20660_not
g52353 not n20525 ; n20525_not
g52354 not n22073 ; n22073_not
g52355 not n12344 ; n12344_not
g52356 not n22046 ; n22046_not
g52357 not n12326 ; n12326_not
g52358 not n20714 ; n20714_not
g52359 not n22028 ; n22028_not
g52360 not n30902 ; n30902_not
g52361 not n12263 ; n12263_not
g52362 not n20750 ; n20750_not
g52363 not n38003 ; n38003_not
g52364 not n38021 ; n38021_not
g52365 not n12236 ; n12236_not
g52366 not n12191 ; n12191_not
g52367 not n20822 ; n20822_not
g52368 not n24350 ; n24350_not
g52369 not n24251 ; n24251_not
g52370 not n14144 ; n14144_not
g52371 not n40451 ; n40451_not
g52372 not n40460 ; n40460_not
g52373 not n37112 ; n37112_not
g52374 not n37121 ; n37121_not
g52375 not n10319 ; n10319_not
g52376 not n18500 ; n18500_not
g52377 not n43151 ; n43151_not
g52378 not n40532 ; n40532_not
g52379 not n14180 ; n14180_not
g52380 not n24323 ; n24323_not
g52381 not n23711 ; n23711_not
g52382 not n24314 ; n24314_not
g52383 not n32810 ; n32810_not
g52384 not n10733 ; n10733_not
g52385 not n32801 ; n32801_not
g52386 not n24305 ; n24305_not
g52387 not n23810 ; n23810_not
g52388 not n40604 ; n40604_not
g52389 not n14054 ; n14054_not
g52390 not n32900 ; n32900_not
g52391 not n14081 ; n14081_not
g52392 not n10337 ; n10337_not
g52393 not n40343 ; n40343_not
g52394 not n14045 ; n14045_not
g52395 not n14090 ; n14090_not
g52396 not n29012 ; n29012_not
g52397 not n47003 ; n47003_not
g52398 not n23603 ; n23603_not
g52399 not n14117 ; n14117_not
g52400 not n10751 ; n10751_not
g52401 not n29030 ; n29030_not
g52402 not n41027 ; n41027_not
g52403 not n40442 ; n40442_not
g52404 not n19031 ; n19031_not
g52405 not n23630 ; n23630_not
g52406 not n14603 ; n14603_not
g52407 not n14504 ; n14504_not
g52408 not n19013 ; n19013_not
g52409 not n14135 ; n14135_not
g52410 not n23900 ; n23900_not
g52411 not n14333 ; n14333_not
g52412 not n24143 ; n24143_not
g52413 not n32711 ; n32711_not
g52414 not n40703 ; n40703_not
g52415 not n32702 ; n32702_not
g52416 not n14351 ; n14351_not
g52417 not n14360 ; n14360_not
g52418 not n40820 ; n40820_not
g52419 not n37004 ; n37004_not
g52420 not n40721 ; n40721_not
g52421 not n40730 ; n40730_not
g52422 not n14441 ; n14441_not
g52423 not n14450 ; n14450_not
g52424 not n32630 ; n32630_not
g52425 not n24062 ; n24062_not
g52426 not n40802 ; n40802_not
g52427 not n24116 ; n24116_not
g52428 not n43124 ; n43124_not
g52429 not n24107 ; n24107_not
g52430 not n43016 ; n43016_not
g52431 not n43142 ; n43142_not
g52432 not n14261 ; n14261_not
g52433 not n40622 ; n40622_not
g52434 not n29111 ; n29111_not
g52435 not n14252 ; n14252_not
g52436 not n14270 ; n14270_not
g52437 not n14531 ; n14531_not
g52438 not n11444 ; n11444_not
g52439 not n24215 ; n24215_not
g52440 not n24206 ; n24206_not
g52441 not n37040 ; n37040_not
g52442 not n32504 ; n32504_not
g52443 not n17051 ; n17051_not
g52444 not n37031 ; n37031_not
g52445 not n14306 ; n14306_not
g52446 not n10724 ; n10724_not
g52447 not n24161 ; n24161_not
g52448 not n14324 ; n14324_not
g52449 not n10292 ; n10292_not
g52450 not n33071 ; n33071_not
g52451 not n33062 ; n33062_not
g52452 not n18320 ; n18320_not
g52453 not n41072 ; n41072_not
g52454 not n43025 ; n43025_not
g52455 not n23441 ; n23441_not
g52456 not n41135 ; n41135_not
g52457 not n43214 ; n43214_not
g52458 not n40370 ; n40370_not
g52459 not n14720 ; n14720_not
g52460 not n33053 ; n33053_not
g52461 not n37211 ; n37211_not
g52462 not n24521 ; n24521_not
g52463 not n43205 ; n43205_not
g52464 not n14702 ; n14702_not
g52465 not n32405 ; n32405_not
g52466 not n43043 ; n43043_not
g52467 not n24512 ; n24512_not
g52468 not n10814 ; n10814_not
g52469 not n33116 ; n33116_not
g52470 not n43007 ; n43007_not
g52471 not n40316 ; n40316_not
g52472 not n33107 ; n33107_not
g52473 not n24404 ; n24404_not
g52474 not n43223 ; n43223_not
g52475 not n33080 ; n33080_not
g52476 not n41009 ; n41009_not
g52477 not n13901 ; n13901_not
g52478 not n40334 ; n40334_not
g52479 not n32324 ; n32324_not
g52480 not n32333 ; n32333_not
g52481 not n23333 ; n23333_not
g52482 not n40352 ; n40352_not
g52483 not n44420 ; n44420_not
g52484 not n43250 ; n43250_not
g52485 not n33008 ; n33008_not
g52486 not n19121 ; n19121_not
g52487 not n10346 ; n10346_not
g52488 not n10805 ; n10805_not
g52489 not n24503 ; n24503_not
g52490 not n32423 ; n32423_not
g52491 not n37202 ; n37202_not
g52492 not n14018 ; n14018_not
g52493 not n41235 ; n41235_not
g52494 not n36420 ; n36420_not
g52495 not n21309 ; n21309_not
g52496 not n21147 ; n21147_not
g52497 not n40830 ; n40830_not
g52498 not n41055 ; n41055_not
g52499 not n24153 ; n24153_not
g52500 not n21372 ; n21372_not
g52501 not n24018 ; n24018_not
g52502 not n26502 ; n26502_not
g52503 not n41163 ; n41163_not
g52504 not n11373 ; n11373_not
g52505 not n22065 ; n22065_not
g52506 not n20661 ; n20661_not
g52507 not n26511 ; n26511_not
g52508 not n21525 ; n21525_not
g52509 not n38013 ; n38013_not
g52510 not n16512 ; n16512_not
g52511 not n21543 ; n21543_not
g52512 not n16224 ; n16224_not
g52513 not n21156 ; n21156_not
g52514 not n17052 ; n17052_not
g52515 not n17025 ; n17025_not
g52516 not n36240 ; n36240_not
g52517 not n18141 ; n18141_not
g52518 not n46041 ; n46041_not
g52519 not n36402 ; n36402_not
g52520 not n20742 ; n20742_not
g52521 not n24612 ; n24612_not
g52522 not n16530 ; n16530_not
g52523 not n36411 ; n36411_not
g52524 not n10527 ; n10527_not
g52525 not n35142 ; n35142_not
g52526 not n18006 ; n18006_not
g52527 not n21183 ; n21183_not
g52528 not n24162 ; n24162_not
g52529 not n16602 ; n16602_not
g52530 not n18411 ; n18411_not
g52531 not n21426 ; n21426_not
g52532 not n21471 ; n21471_not
g52533 not n22128 ; n22128_not
g52534 not n36204 ; n36204_not
g52535 not n26430 ; n26430_not
g52536 not n16611 ; n16611_not
g52537 not n41082 ; n41082_not
g52538 not n26421 ; n26421_not
g52539 not n21174 ; n21174_not
g52540 not n22146 ; n22146_not
g52541 not n42171 ; n42171_not
g52542 not n20571 ; n20571_not
g52543 not n16323 ; n16323_not
g52544 not n22155 ; n22155_not
g52545 not n21444 ; n21444_not
g52546 not n36213 ; n36213_not
g52547 not n22164 ; n22164_not
g52548 not n42072 ; n42072_not
g52549 not n22074 ; n22074_not
g52550 not n41244 ; n41244_not
g52551 not n35160 ; n35160_not
g52552 not n21642 ; n21642_not
g52553 not n16305 ; n16305_not
g52554 not n22083 ; n22083_not
g52555 not n21633 ; n21633_not
g52556 not n21165 ; n21165_not
g52557 not n20652 ; n20652_not
g52558 not n21381 ; n21381_not
g52559 not n42054 ; n42054_not
g52560 not n22092 ; n22092_not
g52561 not n24135 ; n24135_not
g52562 not n41145 ; n41145_not
g52563 not n40812 ; n40812_not
g52564 not n42045 ; n42045_not
g52565 not n16206 ; n16206_not
g52566 not n42036 ; n42036_not
g52567 not n24126 ; n24126_not
g52568 not n24342 ; n24342_not
g52569 not n21606 ; n21606_not
g52570 not n20904 ; n20904_not
g52571 not n21705 ; n21705_not
g52572 not n35016 ; n35016_not
g52573 not n20940 ; n20940_not
g52574 not n21822 ; n21822_not
g52575 not n34431 ; n34431_not
g52576 not n24315 ; n24315_not
g52577 not n16431 ; n16431_not
g52578 not n38211 ; n38211_not
g52579 not n18510 ; n18510_not
g52580 not n24360 ; n24360_not
g52581 not n36303 ; n36303_not
g52582 not n38103 ; n38103_not
g52583 not n47301 ; n47301_not
g52584 not n41091 ; n41091_not
g52585 not n41217 ; n41217_not
g52586 not n42162 ; n42162_not
g52587 not n21714 ; n21714_not
g52588 not n34701 ; n34701_not
g52589 not n15333 ; n15333_not
g52590 not n21219 ; n21219_not
g52591 not n41019 ; n41019_not
g52592 not n16233 ; n16233_not
g52593 not n34602 ; n34602_not
g52594 not n41226 ; n41226_not
g52595 not n21057 ; n21057_not
g52596 not n10554 ; n10554_not
g52597 not n36330 ; n36330_not
g52598 not n24333 ; n24333_not
g52599 not n16251 ; n16251_not
g52600 not n16413 ; n16413_not
g52601 not n21066 ; n21066_not
g52602 not n11445 ; n11445_not
g52603 not n41073 ; n41073_not
g52604 not n24261 ; n24261_not
g52605 not n20841 ; n20841_not
g52606 not n21570 ; n21570_not
g52607 not n18123 ; n18123_not
g52608 not n20832 ; n20832_not
g52609 not n34521 ; n34521_not
g52610 not n21921 ; n21921_not
g52611 not n41208 ; n41208_not
g52612 not n41190 ; n41190_not
g52613 not n21291 ; n21291_not
g52614 not n42126 ; n42126_not
g52615 not n40902 ; n40902_not
g52616 not n20733 ; n20733_not
g52617 not n21552 ; n21552_not
g52618 not n18024 ; n18024_not
g52619 not n18240 ; n18240_not
g52620 not n35133 ; n35133_not
g52621 not n21840 ; n21840_not
g52622 not n41181 ; n41181_not
g52623 not n21228 ; n21228_not
g52624 not n21237 ; n21237_not
g52625 not n24306 ; n24306_not
g52626 not n46023 ; n46023_not
g52627 not n18033 ; n18033_not
g52628 not n35007 ; n35007_not
g52629 not n38301 ; n38301_not
g52630 not n35061 ; n35061_not
g52631 not n16242 ; n16242_not
g52632 not n38400 ; n38400_not
g52633 not n24900 ; n24900_not
g52634 not n18051 ; n18051_not
g52635 not n24702 ; n24702_not
g52636 not n36600 ; n36600_not
g52637 not n34710 ; n34710_not
g52638 not n24270 ; n24270_not
g52639 not n24405 ; n24405_not
g52640 not n17133 ; n17133_not
g52641 not n17430 ; n17430_not
g52642 not n36150 ; n36150_not
g52643 not n35601 ; n35601_not
g52644 not n37320 ; n37320_not
g52645 not n19104 ; n19104_not
g52646 not n17313 ; n17313_not
g52647 not n19122 ; n19122_not
g52648 not n10095 ; n10095_not
g52649 not n23118 ; n23118_not
g52650 not n23532 ; n23532_not
g52651 not n37203 ; n37203_not
g52652 not n41712 ; n41712_not
g52653 not n25602 ; n25602_not
g52654 not n36132 ; n36132_not
g52655 not n23514 ; n23514_not
g52656 not n25170 ; n25170_not
g52657 not n19131 ; n19131_not
g52658 not n40038 ; n40038_not
g52659 not n40146 ; n40146_not
g52660 not n23136 ; n23136_not
g52661 not n40056 ; n40056_not
g52662 not n25413 ; n25413_not
g52663 not n23145 ; n23145_not
g52664 not n25521 ; n25521_not
g52665 not n23073 ; n23073_not
g52666 not n25512 ; n25512_not
g52667 not n19014 ; n19014_not
g52668 not n39120 ; n39120_not
g52669 not n41424 ; n41424_not
g52670 not n39210 ; n39210_not
g52671 not n17124 ; n17124_not
g52672 not n23640 ; n23640_not
g52673 not n23622 ; n23622_not
g52674 not n35403 ; n35403_not
g52675 not n47121 ; n47121_not
g52676 not n35412 ; n35412_not
g52677 not n39300 ; n39300_not
g52678 not n23604 ; n23604_not
g52679 not n17151 ; n17151_not
g52680 not n22740 ; n22740_not
g52681 not n40119 ; n40119_not
g52682 not n22902 ; n22902_not
g52683 not n40083 ; n40083_not
g52684 not n46410 ; n46410_not
g52685 not n40434 ; n40434_not
g52686 not n41442 ; n41442_not
g52687 not n35520 ; n35520_not
g52688 not n17214 ; n17214_not
g52689 not n17223 ; n17223_not
g52690 not n23235 ; n23235_not
g52691 not n37230 ; n37230_not
g52692 not n44511 ; n44511_not
g52693 not n17520 ; n17520_not
g52694 not n23424 ; n23424_not
g52695 not n25332 ; n25332_not
g52696 not n25314 ; n25314_not
g52697 not n25134 ; n25134_not
g52698 not n25215 ; n25215_not
g52699 not n40218 ; n40218_not
g52700 not n41622 ; n41622_not
g52701 not n40263 ; n40263_not
g52702 not n25260 ; n25260_not
g52703 not n25224 ; n25224_not
g52704 not n41604 ; n41604_not
g52705 not n10266 ; n10266_not
g52706 not n10239 ; n10239_not
g52707 not n23334 ; n23334_not
g52708 not n40317 ; n40317_not
g52709 not n23352 ; n23352_not
g52710 not n25233 ; n25233_not
g52711 not n19320 ; n19320_not
g52712 not n23307 ; n23307_not
g52713 not n25242 ; n25242_not
g52714 not n17610 ; n17610_not
g52715 not n25161 ; n25161_not
g52716 not n19302 ; n19302_not
g52717 not n19401 ; n19401_not
g52718 not n25503 ; n25503_not
g52719 not n23154 ; n23154_not
g52720 not n36123 ; n36123_not
g52721 not n19140 ; n19140_not
g52722 not n37302 ; n37302_not
g52723 not n41514 ; n41514_not
g52724 not n45114 ; n45114_not
g52725 not n23505 ; n23505_not
g52726 not n10419 ; n10419_not
g52727 not n40128 ; n40128_not
g52728 not n23271 ; n23271_not
g52729 not n25422 ; n25422_not
g52730 not n37221 ; n37221_not
g52731 not n40371 ; n40371_not
g52732 not n41523 ; n41523_not
g52733 not n46500 ; n46500_not
g52734 not n36024 ; n36024_not
g52735 not n23217 ; n23217_not
g52736 not n40362 ; n40362_not
g52737 not n40155 ; n40155_not
g52738 not n19212 ; n19212_not
g52739 not n17502 ; n17502_not
g52740 not n40173 ; n40173_not
g52741 not n25350 ; n25350_not
g52742 not n23433 ; n23433_not
g52743 not n20391 ; n20391_not
g52744 not n22308 ; n22308_not
g52745 not n26250 ; n26250_not
g52746 not n40704 ; n40704_not
g52747 not n37014 ; n37014_not
g52748 not n23910 ; n23910_not
g52749 not n22326 ; n22326_not
g52750 not n20346 ; n20346_not
g52751 not n26205 ; n26205_not
g52752 not n25008 ; n25008_not
g52753 not n22335 ; n22335_not
g52754 not n22344 ; n22344_not
g52755 not n22362 ; n22362_not
g52756 not n35304 ; n35304_not
g52757 not n41910 ; n41910_not
g52758 not n26106 ; n26106_not
g52759 not n20292 ; n20292_not
g52760 not n20283 ; n20283_not
g52761 not n20274 ; n20274_not
g52762 not n20265 ; n20265_not
g52763 not n20256 ; n20256_not
g52764 not n40641 ; n40641_not
g52765 not n26142 ; n26142_not
g52766 not n20463 ; n20463_not
g52767 not n10509 ; n10509_not
g52768 not n20472 ; n20472_not
g52769 not n24108 ; n24108_not
g52770 not n35223 ; n35223_not
g52771 not n24054 ; n24054_not
g52772 not n20526 ; n20526_not
g52773 not n24072 ; n24072_not
g52774 not n22209 ; n22209_not
g52775 not n24045 ; n24045_not
g52776 not n22218 ; n22218_not
g52777 not n22227 ; n22227_not
g52778 not n22236 ; n22236_not
g52779 not n10491 ; n10491_not
g52780 not n26322 ; n26322_not
g52781 not n26313 ; n26313_not
g52782 not n40731 ; n40731_not
g52783 not n35241 ; n35241_not
g52784 not n41316 ; n41316_not
g52785 not n26304 ; n26304_not
g52786 not n20427 ; n20427_not
g52787 not n22272 ; n22272_not
g52788 not n40713 ; n40713_not
g52789 not n10473 ; n10473_not
g52790 not n22470 ; n22470_not
g52791 not n20094 ; n20094_not
g52792 not n22443 ; n22443_not
g52793 not n22461 ; n22461_not
g52794 not n20085 ; n20085_not
g52795 not n40560 ; n40560_not
g52796 not n20076 ; n20076_not
g52797 not n40542 ; n40542_not
g52798 not n17061 ; n17061_not
g52799 not n20049 ; n20049_not
g52800 not n23703 ; n23703_not
g52801 not n22506 ; n22506_not
g52802 not n26016 ; n26016_not
g52803 not n41406 ; n41406_not
g52804 not n40506 ; n40506_not
g52805 not n37131 ; n37131_not
g52806 not n40533 ; n40533_not
g52807 not n41415 ; n41415_not
g52808 not n37140 ; n37140_not
g52809 not n25071 ; n25071_not
g52810 not n22533 ; n22533_not
g52811 not n47202 ; n47202_not
g52812 not n35313 ; n35313_not
g52813 not n40182 ; n40182_not
g52814 not n22380 ; n22380_not
g52815 not n37050 ; n37050_not
g52816 not n26115 ; n26115_not
g52817 not n22407 ; n22407_not
g52818 not n40632 ; n40632_not
g52819 not n20193 ; n20193_not
g52820 not n41343 ; n41343_not
g52821 not n20184 ; n20184_not
g52822 not n22425 ; n22425_not
g52823 not n35331 ; n35331_not
g52824 not n25026 ; n25026_not
g52825 not n41820 ; n41820_not
g52826 not n39021 ; n39021_not
g52827 not n26061 ; n26061_not
g52828 not n25035 ; n25035_not
g52829 not n45240 ; n45240_not
g52830 not n41370 ; n41370_not
g52831 not n23802 ; n23802_not
g52832 not n45231 ; n45231_not
g52833 not n25044 ; n25044_not
g52834 not n25053 ; n25053_not
g52835 not n29400 ; n29400_not
g52836 not n14172 ; n14172_not
g52837 not n12813 ; n12813_not
g52838 not n30372 ; n30372_not
g52839 not n10635 ; n10635_not
g52840 not n15720 ; n15720_not
g52841 not n34143 ; n34143_not
g52842 not n30525 ; n30525_not
g52843 not n10617 ; n10617_not
g52844 not n32505 ; n32505_not
g52845 not n30345 ; n30345_not
g52846 not n30534 ; n30534_not
g52847 not n43701 ; n43701_not
g52848 not n14208 ; n14208_not
g52849 not n44340 ; n44340_not
g52850 not n12750 ; n12750_not
g52851 not n30561 ; n30561_not
g52852 not n44322 ; n44322_not
g52853 not n30570 ; n30570_not
g52854 not n12723 ; n12723_not
g52855 not n14235 ; n14235_not
g52856 not n12714 ; n12714_not
g52857 not n12705 ; n12705_not
g52858 not n14244 ; n14244_not
g52859 not n14253 ; n14253_not
g52860 not n12408 ; n12408_not
g52861 not n30633 ; n30633_not
g52862 not n30327 ; n30327_not
g52863 not n10752 ; n10752_not
g52864 not n43161 ; n43161_not
g52865 not n34071 ; n34071_not
g52866 not n14091 ; n14091_not
g52867 not n30390 ; n30390_not
g52868 not n28311 ; n28311_not
g52869 not n12903 ; n12903_not
g52870 not n30426 ; n30426_not
g52871 not n30444 ; n30444_not
g52872 not n34107 ; n34107_not
g52873 not n43620 ; n43620_not
g52874 not n28320 ; n28320_not
g52875 not n34116 ; n34116_not
g52876 not n14163 ; n14163_not
g52877 not n34125 ; n34125_not
g52878 not n30462 ; n30462_not
g52879 not n30480 ; n30480_not
g52880 not n12840 ; n12840_not
g52881 not n34134 ; n34134_not
g52882 not n33432 ; n33432_not
g52883 not n12462 ; n12462_not
g52884 not n29310 ; n29310_not
g52885 not n12444 ; n12444_not
g52886 not n31605 ; n31605_not
g52887 not n15180 ; n15180_not
g52888 not n14361 ; n14361_not
g52889 not n30804 ; n30804_not
g52890 not n32604 ; n32604_not
g52891 not n30813 ; n30813_not
g52892 not n47400 ; n47400_not
g52893 not n29301 ; n29301_not
g52894 not n12390 ; n12390_not
g52895 not n10716 ; n10716_not
g52896 not n12381 ; n12381_not
g52897 not n32613 ; n32613_not
g52898 not n28401 ; n28401_not
g52899 not n29211 ; n29211_not
g52900 not n12363 ; n12363_not
g52901 not n32622 ; n32622_not
g52902 not n15162 ; n15162_not
g52903 not n14028 ; n14028_not
g52904 not n12345 ; n12345_not
g52905 not n43116 ; n43116_not
g52906 not n14433 ; n14433_not
g52907 not n29220 ; n29220_not
g52908 not n27420 ; n27420_not
g52909 not n42315 ; n42315_not
g52910 not n30840 ; n30840_not
g52911 not n27600 ; n27600_not
g52912 not n34152 ; n34152_not
g52913 not n30642 ; n30642_not
g52914 not n43152 ; n43152_not
g52915 not n32550 ; n32550_not
g52916 not n44313 ; n44313_not
g52917 not n12570 ; n12570_not
g52918 not n42414 ; n42414_not
g52919 not n27501 ; n27501_not
g52920 not n14280 ; n14280_not
g52921 not n31641 ; n31641_not
g52922 not n12273 ; n12273_not
g52923 not n12561 ; n12561_not
g52924 not n12552 ; n12552_not
g52925 not n14046 ; n14046_not
g52926 not n12534 ; n12534_not
g52927 not n12525 ; n12525_not
g52928 not n15144 ; n15144_not
g52929 not n10725 ; n10725_not
g52930 not n34224 ; n34224_not
g52931 not n30732 ; n30732_not
g52932 not n34233 ; n34233_not
g52933 not n30741 ; n30741_not
g52934 not n30750 ; n30750_not
g52935 not n14334 ; n14334_not
g52936 not n14343 ; n14343_not
g52937 not n43314 ; n43314_not
g52938 not n15405 ; n15405_not
g52939 not n31830 ; n31830_not
g52940 not n10536 ; n10536_not
g52941 not n28140 ; n28140_not
g52942 not n13524 ; n13524_not
g52943 not n31911 ; n31911_not
g52944 not n31902 ; n31902_not
g52945 not n32244 ; n32244_not
g52946 not n13551 ; n13551_not
g52947 not n43305 ; n43305_not
g52948 not n42603 ; n42603_not
g52949 not n33612 ; n33612_not
g52950 not n43422 ; n43422_not
g52951 not n13515 ; n13515_not
g52952 not n10833 ; n10833_not
g52953 not n48300 ; n48300_not
g52954 not n31821 ; n31821_not
g52955 not n33603 ; n33603_not
g52956 not n10644 ; n10644_not
g52957 not n28050 ; n28050_not
g52958 not n30066 ; n30066_not
g52959 not n32271 ; n32271_not
g52960 not n13425 ; n13425_not
g52961 not n28041 ; n28041_not
g52962 not n32325 ; n32325_not
g52963 not n30075 ; n30075_not
g52964 not n43260 ; n43260_not
g52965 not n13407 ; n13407_not
g52966 not n13740 ; n13740_not
g52967 not n32154 ; n32154_not
g52968 not n28113 ; n28113_not
g52969 not n15432 ; n15432_not
g52970 not n28122 ; n28122_not
g52971 not n13731 ; n13731_not
g52972 not n32145 ; n32145_not
g52973 not n15423 ; n15423_not
g52974 not n13722 ; n13722_not
g52975 not n32136 ; n32136_not
g52976 not n10860 ; n10860_not
g52977 not n15441 ; n15441_not
g52978 not n32118 ; n32118_not
g52979 not n32073 ; n32073_not
g52980 not n33621 ; n33621_not
g52981 not n32082 ; n32082_not
g52982 not n13641 ; n13641_not
g52983 not n15414 ; n15414_not
g52984 not n32217 ; n32217_not
g52985 not n15450 ; n15450_not
g52986 not n13605 ; n13605_not
g52987 not n13803 ; n13803_not
g52988 not n10851 ; n10851_not
g52989 not n43413 ; n43413_not
g52990 not n15135 ; n15135_not
g52991 not n13218 ; n13218_not
g52992 not n15306 ; n15306_not
g52993 not n10329 ; n10329_not
g52994 not n10923 ; n10923_not
g52995 not n30255 ; n30255_not
g52996 not n43503 ; n43503_not
g52997 not n11427 ; n11427_not
g52998 not n43512 ; n43512_not
g52999 not n30264 ; n30264_not
g53000 not n14109 ; n14109_not
g53001 not n34017 ; n34017_not
g53002 not n31740 ; n31740_not
g53003 not n10932 ; n10932_not
g53004 not n43521 ; n43521_not
g53005 not n13137 ; n13137_not
g53006 not n13092 ; n13092_not
g53007 not n14127 ; n14127_not
g53008 not n13074 ; n13074_not
g53009 not n42513 ; n42513_not
g53010 not n30291 ; n30291_not
g53011 not n12183 ; n12183_not
g53012 not n28221 ; n28221_not
g53013 not n33513 ; n33513_not
g53014 not n10950 ; n10950_not
g53015 not n30318 ; n30318_not
g53016 not n34053 ; n34053_not
g53017 not n32343 ; n32343_not
g53018 not n43242 ; n43242_not
g53019 not n15351 ; n15351_not
g53020 not n43251 ; n43251_not
g53021 not n13371 ; n13371_not
g53022 not n30129 ; n30129_not
g53023 not n15531 ; n15531_not
g53024 not n32307 ; n32307_not
g53025 not n30138 ; n30138_not
g53026 not n10815 ; n10815_not
g53027 not n10653 ; n10653_not
g53028 not n44403 ; n44403_not
g53029 not n14037 ; n14037_not
g53030 not n13308 ; n13308_not
g53031 not n30183 ; n30183_not
g53032 not n13290 ; n13290_not
g53033 not n33810 ; n33810_not
g53034 not n10572 ; n10572_not
g53035 not n30228 ; n30228_not
g53036 not n30237 ; n30237_not
g53037 not n32451 ; n32451_not
g53038 not n15324 ; n15324_not
g53039 not n13254 ; n13254_not
g53040 not n32460 ; n32460_not
g53041 not n10770 ; n10770_not
g53042 not n16008 ; n16008_not
g53043 not n11922 ; n11922_not
g53044 not n15900 ; n15900_not
g53045 not n31128 ; n31128_not
g53046 not n43062 ; n43062_not
g53047 not n11904 ; n11904_not
g53048 not n16026 ; n16026_not
g53049 not n15027 ; n15027_not
g53050 not n31434 ; n31434_not
g53051 not n44034 ; n44034_not
g53052 not n42207 ; n42207_not
g53053 not n43044 ; n43044_not
g53054 not n31164 ; n31164_not
g53055 not n11823 ; n11823_not
g53056 not n11832 ; n11832_not
g53057 not n11841 ; n11841_not
g53058 not n31182 ; n31182_not
g53059 not n31191 ; n31191_not
g53060 not n16035 ; n16035_not
g53061 not n16044 ; n16044_not
g53062 not n33333 ; n33333_not
g53063 not n44052 ; n44052_not
g53064 not n27303 ; n27303_not
g53065 not n31038 ; n31038_not
g53066 not n44241 ; n44241_not
g53067 not n10608 ; n10608_not
g53068 not n43071 ; n43071_not
g53069 not n14505 ; n14505_not
g53070 not n12039 ; n12039_not
g53071 not n14604 ; n14604_not
g53072 not n15063 ; n15063_not
g53073 not n11238 ; n11238_not
g53074 not n29022 ; n29022_not
g53075 not n44016 ; n44016_not
g53076 not n34422 ; n34422_not
g53077 not n11940 ; n11940_not
g53078 not n14631 ; n14631_not
g53079 not n29013 ; n29013_not
g53080 not n11247 ; n11247_not
g53081 not n42225 ; n42225_not
g53082 not n33351 ; n33351_not
g53083 not n42216 ; n42216_not
g53084 not n44430 ; n44430_not
g53085 not n31353 ; n31353_not
g53086 not n14811 ; n14811_not
g53087 not n31290 ; n31290_not
g53088 not n33270 ; n33270_not
g53089 not n11580 ; n11580_not
g53090 not n27060 ; n27060_not
g53091 not n33252 ; n33252_not
g53092 not n33180 ; n33180_not
g53093 not n44133 ; n44133_not
g53094 not n16170 ; n16170_not
g53095 not n44142 ; n44142_not
g53096 not n16143 ; n16143_not
g53097 not n11490 ; n11490_not
g53098 not n16152 ; n16152_not
g53099 not n11481 ; n11481_not
g53100 not n31344 ; n31344_not
g53101 not n16161 ; n16161_not
g53102 not n31317 ; n31317_not
g53103 not n44412 ; n44412_not
g53104 not n31371 ; n31371_not
g53105 not n34512 ; n34512_not
g53106 not n42180 ; n42180_not
g53107 not n43035 ; n43035_not
g53108 not n42711 ; n42711_not
g53109 not n33045 ; n33045_not
g53110 not n11814 ; n11814_not
g53111 not n31425 ; n31425_not
g53112 not n33072 ; n33072_not
g53113 not n11760 ; n11760_not
g53114 not n33315 ; n33315_not
g53115 not n16062 ; n16062_not
g53116 not n27204 ; n27204_not
g53117 not n31119 ; n31119_not
g53118 not n11733 ; n11733_not
g53119 not n41118 ; n41118_not
g53120 not n44106 ; n44106_not
g53121 not n43008 ; n43008_not
g53122 not n11346 ; n11346_not
g53123 not n39111 ; n39111_not
g53124 not n11670 ; n11670_not
g53125 not n11661 ; n11661_not
g53126 not n14442 ; n14442_not
g53127 not n14514 ; n14514_not
g53128 not n33135 ; n33135_not
g53129 not n31263 ; n31263_not
g53130 not n14802 ; n14802_not
g53131 not n32730 ; n32730_not
g53132 not n12084 ; n12084_not
g53133 not n12219 ; n12219_not
g53134 not n41046 ; n41046_not
g53135 not n10707 ; n10707_not
g53136 not n11193 ; n11193_not
g53137 not n15117 ; n15117_not
g53138 not n31515 ; n31515_not
g53139 not n27321 ; n27321_not
g53140 not n14532 ; n14532_not
g53141 not n15126 ; n15126_not
g53142 not n11166 ; n11166_not
g53143 not n11175 ; n11175_not
g53144 not n30912 ; n30912_not
g53145 not n34305 ; n34305_not
g53146 not n29103 ; n29103_not
g53147 not n14523 ; n14523_not
g53148 not n12156 ; n12156_not
g53149 not n12066 ; n12066_not
g53150 not n12291 ; n12291_not
g53151 not n34332 ; n34332_not
g53152 not n12147 ; n12147_not
g53153 not n43080 ; n43080_not
g53154 not n12138 ; n12138_not
g53155 not n42261 ; n42261_not
g53156 not n12174 ; n12174_not
g53157 not n42243 ; n42243_not
g53158 not n15081 ; n15081_not
g53159 not n42306 ; n42306_not
g53160 not n12228 ; n12228_not
g53161 not n12246 ; n12246_not
g53162 not n27411 ; n27411_not
g53163 not n28212 ; n28212_not
g53164 not n32272 ; n32272_not
g53165 not n18205 ; n18205_not
g53166 not n14812 ; n14812_not
g53167 not n19312 ; n19312_not
g53168 not n32281 ; n32281_not
g53169 not n23362 ; n23362_not
g53170 not n47023 ; n47023_not
g53171 not n10834 ; n10834_not
g53172 not n19321 ; n19321_not
g53173 not n41182 ; n41182_not
g53174 not n41191 ; n41191_not
g53175 not n24145 ; n24145_not
g53176 not n40831 ; n40831_not
g53177 not n40381 ; n40381_not
g53178 not n32704 ; n32704_not
g53179 not n32263 ; n32263_not
g53180 not n33136 ; n33136_not
g53181 not n43216 ; n43216_not
g53182 not n32371 ; n32371_not
g53183 not n23452 ; n23452_not
g53184 not n32362 ; n32362_not
g53185 not n16630 ; n16630_not
g53186 not n24613 ; n24613_not
g53187 not n23443 ; n23443_not
g53188 not n32353 ; n32353_not
g53189 not n23416 ; n23416_not
g53190 not n23227 ; n23227_not
g53191 not n24181 ; n24181_not
g53192 not n23407 ; n23407_not
g53193 not n23254 ; n23254_not
g53194 not n13921 ; n13921_not
g53195 not n32335 ; n32335_not
g53196 not n33154 ; n33154_not
g53197 not n40840 ; n40840_not
g53198 not n24631 ; n24631_not
g53199 not n13903 ; n13903_not
g53200 not n40327 ; n40327_not
g53201 not n19204 ; n19204_not
g53202 not n14803 ; n14803_not
g53203 not n32317 ; n32317_not
g53204 not n32290 ; n32290_not
g53205 not n18214 ; n18214_not
g53206 not n40066 ; n40066_not
g53207 not n42460 ; n42460_not
g53208 not n46510 ; n46510_not
g53209 not n41209 ; n41209_not
g53210 not n13741 ; n13741_not
g53211 not n23281 ; n23281_not
g53212 not n24082 ; n24082_not
g53213 not n24811 ; n24811_not
g53214 not n19411 ; n19411_not
g53215 not n23272 ; n23272_not
g53216 not n17233 ; n17233_not
g53217 not n36340 ; n36340_not
g53218 not n32209 ; n32209_not
g53219 not n40237 ; n40237_not
g53220 not n24064 ; n24064_not
g53221 not n39112 ; n39112_not
g53222 not n29212 ; n29212_not
g53223 not n32182 ; n32182_not
g53224 not n33217 ; n33217_not
g53225 not n36304 ; n36304_not
g53226 not n36331 ; n36331_not
g53227 not n32173 ; n32173_not
g53228 not n32533 ; n32533_not
g53229 not n43108 ; n43108_not
g53230 not n17404 ; n17404_not
g53231 not n18070 ; n18070_not
g53232 not n33226 ; n33226_not
g53233 not n42604 ; n42604_not
g53234 not n40813 ; n40813_not
g53235 not n14452 ; n14452_not
g53236 not n32245 ; n32245_not
g53237 not n24019 ; n24019_not
g53238 not n23344 ; n23344_not
g53239 not n36430 ; n36430_not
g53240 not n19330 ; n19330_not
g53241 not n33181 ; n33181_not
g53242 not n24730 ; n24730_not
g53243 not n23326 ; n23326_not
g53244 not n29203 ; n29203_not
g53245 not n24703 ; n24703_not
g53246 not n40741 ; n40741_not
g53247 not n18700 ; n18700_not
g53248 not n13822 ; n13822_not
g53249 not n43333 ; n43333_not
g53250 not n40255 ; n40255_not
g53251 not n18124 ; n18124_not
g53252 not n40246 ; n40246_not
g53253 not n14407 ; n14407_not
g53254 not n24802 ; n24802_not
g53255 not n40273 ; n40273_not
g53256 not n10366 ; n10366_not
g53257 not n40750 ; n40750_not
g53258 not n33208 ; n33208_not
g53259 not n10843 ; n10843_not
g53260 not n18142 ; n18142_not
g53261 not n23308 ; n23308_not
g53262 not n32560 ; n32560_not
g53263 not n32227 ; n32227_not
g53264 not n40282 ; n40282_not
g53265 not n33190 ; n33190_not
g53266 not n23821 ; n23821_not
g53267 not n18520 ; n18520_not
g53268 not n14623 ; n14623_not
g53269 not n37123 ; n37123_not
g53270 not n41056 ; n41056_not
g53271 not n10753 ; n10753_not
g53272 not n14650 ; n14650_not
g53273 not n18403 ; n18403_not
g53274 not n32551 ; n32551_not
g53275 not n14029 ; n14029_not
g53276 not n40462 ; n40462_not
g53277 not n36610 ; n36610_not
g53278 not n24316 ; n24316_not
g53279 not n24226 ; n24226_not
g53280 not n14551 ; n14551_not
g53281 not n40633 ; n40633_not
g53282 not n40453 ; n40453_not
g53283 not n14155 ; n14155_not
g53284 not n36700 ; n36700_not
g53285 not n29401 ; n29401_not
g53286 not n23830 ; n23830_not
g53287 not n37060 ; n37060_not
g53288 not n44611 ; n44611_not
g53289 not n19006 ; n19006_not
g53290 not n40642 ; n40642_not
g53291 not n32911 ; n32911_not
g53292 not n10348 ; n10348_not
g53293 not n19024 ; n19024_not
g53294 not n24271 ; n24271_not
g53295 not n32506 ; n32506_not
g53296 not n23803 ; n23803_not
g53297 not n23722 ; n23722_not
g53298 not n20923 ; n20923_not
g53299 not n44413 ; n44413_not
g53300 not n14218 ; n14218_not
g53301 not n40570 ; n40570_not
g53302 not n29050 ; n29050_not
g53303 not n10744 ; n10744_not
g53304 not n24244 ; n24244_not
g53305 not n37105 ; n37105_not
g53306 not n29005 ; n29005_not
g53307 not n32542 ; n32542_not
g53308 not n32830 ; n32830_not
g53309 not n41029 ; n41029_not
g53310 not n14605 ; n14605_not
g53311 not n29023 ; n29023_not
g53312 not n18502 ; n18502_not
g53313 not n40543 ; n40543_not
g53314 not n23812 ; n23812_not
g53315 not n24325 ; n24325_not
g53316 not n14506 ; n14506_not
g53317 not n40615 ; n40615_not
g53318 not n41047 ; n41047_not
g53319 not n14164 ; n14164_not
g53320 not n40165 ; n40165_not
g53321 not n32821 ; n32821_not
g53322 not n14641 ; n14641_not
g53323 not n18304 ; n18304_not
g53324 not n32605 ; n32605_not
g53325 not n14083 ; n14083_not
g53326 not n40417 ; n40417_not
g53327 not n33055 ; n33055_not
g53328 not n14362 ; n14362_not
g53329 not n19105 ; n19105_not
g53330 not n14056 ; n14056_not
g53331 not n43018 ; n43018_not
g53332 not n32434 ; n32434_not
g53333 not n19114 ; n19114_not
g53334 not n40408 ; n40408_not
g53335 not n18106 ; n18106_not
g53336 not n10771 ; n10771_not
g53337 not n41083 ; n41083_not
g53338 not n13453 ; n13453_not
g53339 not n23524 ; n23524_not
g53340 not n32416 ; n32416_not
g53341 not n32731 ; n32731_not
g53342 not n10816 ; n10816_not
g53343 not n23515 ; n23515_not
g53344 not n36520 ; n36520_not
g53345 not n36403 ; n36403_not
g53346 not n41155 ; n41155_not
g53347 not n18250 ; n18250_not
g53348 not n10825 ; n10825_not
g53349 not n40390 ; n40390_not
g53350 not n40651 ; n40651_not
g53351 not n24442 ; n24442_not
g53352 not n41128 ; n41128_not
g53353 not n43045 ; n43045_not
g53354 not n37015 ; n37015_not
g53355 not n14128 ; n14128_not
g53356 not n40444 ; n40444_not
g53357 not n23623 ; n23623_not
g53358 not n29113 ; n29113_not
g53359 not n14119 ; n14119_not
g53360 not n33037 ; n33037_not
g53361 not n23614 ; n23614_not
g53362 not n10645 ; n10645_not
g53363 not n37150 ; n37150_not
g53364 not n14713 ; n14713_not
g53365 not n24523 ; n24523_not
g53366 not n24262 ; n24262_not
g53367 not n29320 ; n29320_not
g53368 not n33046 ; n33046_not
g53369 not n24532 ; n24532_not
g53370 not n33019 ; n33019_not
g53371 not n24541 ; n24541_not
g53372 not n29122 ; n29122_not
g53373 not n24550 ; n24550_not
g53374 not n10618 ; n10618_not
g53375 not n14731 ; n14731_not
g53376 not n18313 ; n18313_not
g53377 not n24235 ; n24235_not
g53378 not n21850 ; n21850_not
g53379 not n31480 ; n31480_not
g53380 not n44242 ; n44242_not
g53381 not n11176 ; n11176_not
g53382 not n20860 ; n20860_not
g53383 not n21094 ; n21094_not
g53384 not n31507 ; n31507_not
g53385 not n38410 ; n38410_not
g53386 not n20824 ; n20824_not
g53387 not n20815 ; n20815_not
g53388 not n46033 ; n46033_not
g53389 not n12193 ; n12193_not
g53390 not n20806 ; n20806_not
g53391 not n30940 ; n30940_not
g53392 not n11149 ; n11149_not
g53393 not n38041 ; n38041_not
g53394 not n30931 ; n30931_not
g53395 not n38032 ; n38032_not
g53396 not n44260 ; n44260_not
g53397 not n21922 ; n21922_not
g53398 not n12256 ; n12256_not
g53399 not n34900 ; n34900_not
g53400 not n21724 ; n21724_not
g53401 not n44008 ; n44008_not
g53402 not n38311 ; n38311_not
g53403 not n21751 ; n21751_not
g53404 not n38320 ; n38320_not
g53405 not n20905 ; n20905_not
g53406 not n12049 ; n12049_not
g53407 not n12067 ; n12067_not
g53408 not n20950 ; n20950_not
g53409 not n20941 ; n20941_not
g53410 not n31462 ; n31462_not
g53411 not n20932 ; n20932_not
g53412 not n20914 ; n20914_not
g53413 not n12094 ; n12094_not
g53414 not n11194 ; n11194_not
g53415 not n12184 ; n12184_not
g53416 not n11077 ; n11077_not
g53417 not n30832 ; n30832_not
g53418 not n31570 ; n31570_not
g53419 not n20644 ; n20644_not
g53420 not n20635 ; n20635_not
g53421 not n20626 ; n20626_not
g53422 not n30805 ; n30805_not
g53423 not n12427 ; n12427_not
g53424 not n20617 ; n20617_not
g53425 not n31624 ; n31624_not
g53426 not n20590 ; n20590_not
g53427 not n46132 ; n46132_not
g53428 not n20581 ; n20581_not
g53429 not n22138 ; n22138_not
g53430 not n31552 ; n31552_not
g53431 not n12481 ; n12481_not
g53432 not n20563 ; n20563_not
g53433 not n22156 ; n22156_not
g53434 not n12508 ; n12508_not
g53435 not n12517 ; n12517_not
g53436 not n30724 ; n30724_not
g53437 not n30922 ; n30922_not
g53438 not n46042 ; n46042_not
g53439 not n20734 ; n20734_not
g53440 not n12283 ; n12283_not
g53441 not n30904 ; n30904_not
g53442 not n12292 ; n12292_not
g53443 not n11095 ; n11095_not
g53444 not n22039 ; n22039_not
g53445 not n12319 ; n12319_not
g53446 not n12328 ; n12328_not
g53447 not n20680 ; n20680_not
g53448 not n12346 ; n12346_not
g53449 not n30850 ; n30850_not
g53450 not n22066 ; n22066_not
g53451 not n20671 ; n20671_not
g53452 not n12355 ; n12355_not
g53453 not n30841 ; n30841_not
g53454 not n11572 ; n11572_not
g53455 not n11563 ; n11563_not
g53456 not n31408 ; n31408_not
g53457 not n31291 ; n31291_not
g53458 not n11590 ; n11590_not
g53459 not n31273 ; n31273_not
g53460 not n21328 ; n21328_not
g53461 not n21535 ; n21535_not
g53462 not n21319 ; n21319_not
g53463 not n11608 ; n11608_not
g53464 not n11617 ; n11617_not
g53465 not n21544 ; n21544_not
g53466 not n11365 ; n11365_not
g53467 not n21292 ; n21292_not
g53468 not n21562 ; n21562_not
g53469 not n21283 ; n21283_not
g53470 not n11653 ; n11653_not
g53471 not n21274 ; n21274_not
g53472 not n21580 ; n21580_not
g53473 not n21256 ; n21256_not
g53474 not n11680 ; n11680_not
g53475 not n31255 ; n31255_not
g53476 not n31309 ; n31309_not
g53477 not n31381 ; n31381_not
g53478 not n21463 ; n21463_not
g53479 not n21436 ; n21436_not
g53480 not n31363 ; n31363_not
g53481 not n11464 ; n11464_not
g53482 not n21427 ; n21427_not
g53483 not n21490 ; n21490_not
g53484 not n21409 ; n21409_not
g53485 not n11482 ; n11482_not
g53486 not n31336 ; n31336_not
g53487 not n31327 ; n31327_not
g53488 not n21391 ; n21391_not
g53489 not n11518 ; n11518_not
g53490 not n21382 ; n21382_not
g53491 not n11527 ; n11527_not
g53492 not n21517 ; n21517_not
g53493 not n31318 ; n31318_not
g53494 not n21364 ; n21364_not
g53495 not n11824 ; n11824_not
g53496 not n38203 ; n38203_not
g53497 not n45601 ; n45601_not
g53498 not n21166 ; n21166_not
g53499 not n21157 ; n21157_not
g53500 not n11842 ; n11842_not
g53501 not n31174 ; n31174_not
g53502 not n21139 ; n21139_not
g53503 not n44053 ; n44053_not
g53504 not n31075 ; n31075_not
g53505 not n31147 ; n31147_not
g53506 not n11905 ; n11905_not
g53507 not n21670 ; n21670_not
g53508 not n11914 ; n11914_not
g53509 not n21085 ; n21085_not
g53510 not n21706 ; n21706_not
g53511 not n31093 ; n31093_not
g53512 not n11257 ; n11257_not
g53513 not n11950 ; n11950_not
g53514 not n11707 ; n11707_not
g53515 not n21247 ; n21247_not
g53516 not n10069 ; n10069_not
g53517 not n21238 ; n21238_not
g53518 not n21229 ; n21229_not
g53519 not n11734 ; n11734_not
g53520 not n44215 ; n44215_not
g53521 not n11752 ; n11752_not
g53522 not n31228 ; n31228_not
g53523 not n31219 ; n31219_not
g53524 not n31417 ; n31417_not
g53525 not n21616 ; n21616_not
g53526 not n21193 ; n21193_not
g53527 not n44224 ; n44224_not
g53528 not n44071 ; n44071_not
g53529 not n44062 ; n44062_not
g53530 not n11806 ; n11806_not
g53531 not n44044 ; n44044_not
g53532 not n21175 ; n21175_not
g53533 not n11815 ; n11815_not
g53534 not n22921 ; n22921_not
g53535 not n22930 ; n22930_not
g53536 not n37411 ; n37411_not
g53537 not n43450 ; n43450_not
g53538 not n13417 ; n13417_not
g53539 not n30076 ; n30076_not
g53540 not n13426 ; n13426_not
g53541 not n23029 ; n23029_not
g53542 not n37321 ; n37321_not
g53543 not n43441 ; n43441_not
g53544 not n30067 ; n30067_not
g53545 not n17422 ; n17422_not
g53546 not n13471 ; n13471_not
g53547 not n30058 ; n30058_not
g53548 not n43423 ; n43423_not
g53549 not n37312 ; n37312_not
g53550 not n23074 ; n23074_not
g53551 not n23092 ; n23092_not
g53552 not n13516 ; n13516_not
g53553 not n13345 ; n13345_not
g53554 not n22642 ; n22642_not
g53555 not n13354 ; n13354_not
g53556 not n22606 ; n22606_not
g53557 not n30139 ; n30139_not
g53558 not n22651 ; n22651_not
g53559 not n39310 ; n39310_not
g53560 not n31804 ; n31804_not
g53561 not n13372 ; n13372_not
g53562 not n37600 ; n37600_not
g53563 not n22723 ; n22723_not
g53564 not n30094 ; n30094_not
g53565 not n39400 ; n39400_not
g53566 not n22732 ; n22732_not
g53567 not n39202 ; n39202_not
g53568 not n30085 ; n30085_not
g53569 not n31813 ; n31813_not
g53570 not n37501 ; n37501_not
g53571 not n22813 ; n22813_not
g53572 not n22804 ; n22804_not
g53573 not n22912 ; n22912_not
g53574 not n13462 ; n13462_not
g53575 not n23083 ; n23083_not
g53576 not n13624 ; n13624_not
g53577 not n13633 ; n13633_not
g53578 not n32047 ; n32047_not
g53579 not n32056 ; n32056_not
g53580 not n10195 ; n10195_not
g53581 not n13651 ; n13651_not
g53582 not n32074 ; n32074_not
g53583 not n40138 ; n40138_not
g53584 not n23173 ; n23173_not
g53585 not n40147 ; n40147_not
g53586 not n48220 ; n48220_not
g53587 not n32029 ; n32029_not
g53588 not n23209 ; n23209_not
g53589 not n32128 ; n32128_not
g53590 not n19501 ; n19501_not
g53591 not n40174 ; n40174_not
g53592 not n10609 ; n10609_not
g53593 not n40183 ; n40183_not
g53594 not n32164 ; n32164_not
g53595 not n13525 ; n13525_not
g53596 not n10537 ; n10537_not
g53597 not n10870 ; n10870_not
g53598 not n13534 ; n13534_not
g53599 not n23119 ; n23119_not
g53600 not n31840 ; n31840_not
g53601 not n44404 ; n44404_not
g53602 not n23047 ; n23047_not
g53603 not n40039 ; n40039_not
g53604 not n45124 ; n45124_not
g53605 not n23137 ; n23137_not
g53606 not n40048 ; n40048_not
g53607 not n13570 ; n13570_not
g53608 not n23065 ; n23065_not
g53609 not n43414 ; n43414_not
g53610 not n23146 ; n23146_not
g53611 not n37303 ; n37303_not
g53612 not n40075 ; n40075_not
g53613 not n13606 ; n13606_not
g53614 not n13615 ; n13615_not
g53615 not n12724 ; n12724_not
g53616 not n22327 ; n22327_not
g53617 not n20356 ; n20356_not
g53618 not n30571 ; n30571_not
g53619 not n44332 ; n44332_not
g53620 not n30544 ; n30544_not
g53621 not n20329 ; n20329_not
g53622 not n45340 ; n45340_not
g53623 not n30535 ; n30535_not
g53624 not n30526 ; n30526_not
g53625 not n12805 ; n12805_not
g53626 not n46213 ; n46213_not
g53627 not n12823 ; n12823_not
g53628 not n12832 ; n12832_not
g53629 not n30490 ; n30490_not
g53630 not n43630 ; n43630_not
g53631 not n30463 ; n30463_not
g53632 not n31705 ; n31705_not
g53633 not n20239 ; n20239_not
g53634 not n30445 ; n30445_not
g53635 not n30436 ; n30436_not
g53636 not n12922 ; n12922_not
g53637 not n22192 ; n22192_not
g53638 not n12544 ; n12544_not
g53639 not n30715 ; n30715_not
g53640 not n20518 ; n20518_not
g53641 not n12571 ; n12571_not
g53642 not n22228 ; n22228_not
g53643 not n31651 ; n31651_not
g53644 not n22246 ; n22246_not
g53645 not n20473 ; n20473_not
g53646 not n22255 ; n22255_not
g53647 not n20455 ; n20455_not
g53648 not n12616 ; n12616_not
g53649 not n22264 ; n22264_not
g53650 not n12634 ; n12634_not
g53651 not n20428 ; n20428_not
g53652 not n20419 ; n20419_not
g53653 not n22282 ; n22282_not
g53654 not n22291 ; n22291_not
g53655 not n20392 ; n20392_not
g53656 not n22309 ; n22309_not
g53657 not n22318 ; n22318_not
g53658 not n30580 ; n30580_not
g53659 not n10915 ; n10915_not
g53660 not n13237 ; n13237_not
g53661 not n13246 ; n13246_not
g53662 not n46303 ; n46303_not
g53663 not n10078 ; n10078_not
g53664 not n30238 ; n30238_not
g53665 not n39103 ; n39103_not
g53666 not n10096 ; n10096_not
g53667 not n13273 ; n13273_not
g53668 not n46060 ; n46060_not
g53669 not n22543 ; n22543_not
g53670 not n22552 ; n22552_not
g53671 not n22561 ; n22561_not
g53672 not n31750 ; n31750_not
g53673 not n46321 ; n46321_not
g53674 not n30157 ; n30157_not
g53675 not n39220 ; n39220_not
g53676 not n46312 ; n46312_not
g53677 not n13336 ; n13336_not
g53678 not n39004 ; n39004_not
g53679 not n12931 ; n12931_not
g53680 not n22417 ; n22417_not
g53681 not n30382 ; n30382_not
g53682 not n30364 ; n30364_not
g53683 not n30355 ; n30355_not
g53684 not n31732 ; n31732_not
g53685 not n30337 ; n30337_not
g53686 not n20149 ; n20149_not
g53687 not n39022 ; n39022_not
g53688 not n10960 ; n10960_not
g53689 not n12841 ; n12841_not
g53690 not n30283 ; n30283_not
g53691 not n20095 ; n20095_not
g53692 not n13093 ; n13093_not
g53693 not n10942 ; n10942_not
g53694 not n20068 ; n20068_not
g53695 not n13147 ; n13147_not
g53696 not n13165 ; n13165_not
g53697 not n10933 ; n10933_not
g53698 not n20059 ; n20059_not
g53699 not n11419 ; n11419_not
g53700 not n13228 ; n13228_not
g53701 not n36124 ; n36124_not
g53702 not n16711 ; n16711_not
g53703 not n33451 ; n33451_not
g53704 not n42622 ; n42622_not
g53705 not n26332 ; n26332_not
g53706 not n41506 ; n41506_not
g53707 not n25162 ; n25162_not
g53708 not n10492 ; n10492_not
g53709 not n35242 ; n35242_not
g53710 not n11446 ; n11446_not
g53711 not n42370 ; n42370_not
g53712 not n35224 ; n35224_not
g53713 not n15190 ; n15190_not
g53714 not n33442 ; n33442_not
g53715 not n35215 ; n35215_not
g53716 not n34243 ; n34243_not
g53717 not n41470 ; n41470_not
g53718 not n34261 ; n34261_not
g53719 not n42019 ; n42019_not
g53720 not n26404 ; n26404_not
g53721 not n41461 ; n41461_not
g53722 not n34270 ; n34270_not
g53723 not n10519 ; n10519_not
g53724 not n41452 ; n41452_not
g53725 not n10465 ; n10465_not
g53726 not n26224 ; n26224_not
g53727 not n36115 ; n36115_not
g53728 not n25153 ; n25153_not
g53729 not n41830 ; n41830_not
g53730 not n33505 ; n33505_not
g53731 not n34153 ; n34153_not
g53732 not n26251 ; n26251_not
g53733 not n41551 ; n41551_not
g53734 not n15244 ; n15244_not
g53735 not n26260 ; n26260_not
g53736 not n10528 ; n10528_not
g53737 not n41533 ; n41533_not
g53738 not n35260 ; n35260_not
g53739 not n10474 ; n10474_not
g53740 not n15226 ; n15226_not
g53741 not n15217 ; n15217_not
g53742 not n14443 ; n14443_not
g53743 not n17701 ; n17701_not
g53744 not n40525 ; n40525_not
g53745 not n34207 ; n34207_not
g53746 not n44422 ; n44422_not
g53747 not n26530 ; n26530_not
g53748 not n28420 ; n28420_not
g53749 not n15910 ; n15910_not
g53750 not n35143 ; n35143_not
g53751 not n25063 ; n25063_not
g53752 not n34324 ; n34324_not
g53753 not n41407 ; n41407_not
g53754 not n15127 ; n15127_not
g53755 not n42082 ; n42082_not
g53756 not n35134 ; n35134_not
g53757 not n34333 ; n34333_not
g53758 not n42280 ; n42280_not
g53759 not n33406 ; n33406_not
g53760 not n42271 ; n42271_not
g53761 not n17143 ; n17143_not
g53762 not n35107 ; n35107_not
g53763 not n27313 ; n27313_not
g53764 not n41371 ; n41371_not
g53765 not n33370 ; n33370_not
g53766 not n33361 ; n33361_not
g53767 not n16450 ; n16450_not
g53768 not n41317 ; n41317_not
g53769 not n42253 ; n42253_not
g53770 not n26602 ; n26602_not
g53771 not n41353 ; n41353_not
g53772 not n16441 ; n16441_not
g53773 not n15172 ; n15172_not
g53774 not n15820 ; n15820_not
g53775 not n42352 ; n42352_not
g53776 not n10627 ; n10627_not
g53777 not n14515 ; n14515_not
g53778 not n41335 ; n41335_not
g53779 not n27250 ; n27250_not
g53780 not n16603 ; n16603_not
g53781 not n15154 ; n15154_not
g53782 not n36151 ; n36151_not
g53783 not n25108 ; n25108_not
g53784 not n27241 ; n27241_not
g53785 not n35170 ; n35170_not
g53786 not n47122 ; n47122_not
g53787 not n35152 ; n35152_not
g53788 not n42073 ; n42073_not
g53789 not n28411 ; n28411_not
g53790 not n17800 ; n17800_not
g53791 not n36160 ; n36160_not
g53792 not n16531 ; n16531_not
g53793 not n26503 ; n26503_not
g53794 not n15145 ; n15145_not
g53795 not n16540 ; n16540_not
g53796 not n26521 ; n26521_not
g53797 not n35440 ; n35440_not
g53798 not n25540 ; n25540_not
g53799 not n28042 ; n28042_not
g53800 not n35431 ; n35431_not
g53801 not n25531 ; n25531_not
g53802 not n15505 ; n15505_not
g53803 not n35422 ; n35422_not
g53804 not n28015 ; n28015_not
g53805 not n25513 ; n25513_not
g53806 not n42541 ; n42541_not
g53807 not n17431 ; n17431_not
g53808 not n25504 ; n25504_not
g53809 not n15514 ; n15514_not
g53810 not n17116 ; n17116_not
g53811 not n35206 ; n35206_not
g53812 not n33712 ; n33712_not
g53813 not n33730 ; n33730_not
g53814 not n36016 ; n36016_not
g53815 not n25441 ; n25441_not
g53816 not n33622 ; n33622_not
g53817 not n15550 ; n15550_not
g53818 not n26017 ; n26017_not
g53819 not n17305 ; n17305_not
g53820 not n35701 ; n35701_not
g53821 not n41731 ; n41731_not
g53822 not n15460 ; n15460_not
g53823 not n28105 ; n28105_not
g53824 not n25720 ; n25720_not
g53825 not n25711 ; n25711_not
g53826 not n17242 ; n17242_not
g53827 not n41722 ; n41722_not
g53828 not n25810 ; n25810_not
g53829 not n35620 ; n35620_not
g53830 not n25630 ; n25630_not
g53831 not n42550 ; n42550_not
g53832 not n28060 ; n28060_not
g53833 not n35530 ; n35530_not
g53834 not n35521 ; n35521_not
g53835 not n28024 ; n28024_not
g53836 not n35503 ; n35503_not
g53837 not n41713 ; n41713_not
g53838 not n41704 ; n41704_not
g53839 not n41740 ; n41740_not
g53840 not n15442 ; n15442_not
g53841 not n25900 ; n25900_not
g53842 not n41632 ; n41632_not
g53843 not n26080 ; n26080_not
g53844 not n35332 ; n35332_not
g53845 not n28222 ; n28222_not
g53846 not n15343 ; n15343_not
g53847 not n15640 ; n15640_not
g53848 not n34063 ; n34063_not
g53849 not n26107 ; n26107_not
g53850 not n41623 ; n41623_not
g53851 not n34081 ; n34081_not
g53852 not n27700 ; n27700_not
g53853 not n41614 ; n41614_not
g53854 not n15325 ; n15325_not
g53855 not n26125 ; n26125_not
g53856 not n25252 ; n25252_not
g53857 not n40714 ; n40714_not
g53858 not n15316 ; n15316_not
g53859 not n26161 ; n26161_not
g53860 not n12373 ; n12373_not
g53861 not n17620 ; n17620_not
g53862 not n34144 ; n34144_not
g53863 not n41920 ; n41920_not
g53864 not n26206 ; n26206_not
g53865 not n15280 ; n15280_not
g53866 not n25414 ; n25414_not
g53867 not n33604 ; n33604_not
g53868 not n15370 ; n15370_not
g53869 not n42532 ; n42532_not
g53870 not n36034 ; n36034_not
g53871 not n17008 ; n17008_not
g53872 not n25360 ; n25360_not
g53873 not n36052 ; n36052_not
g53874 not n17062 ; n17062_not
g53875 not n33820 ; n33820_not
g53876 not n33541 ; n33541_not
g53877 not n17044 ; n17044_not
g53878 not n26035 ; n26035_not
g53879 not n25351 ; n25351_not
g53880 not n36007 ; n36007_not
g53881 not n33703 ; n33703_not
g53882 not n28204 ; n28204_not
g53883 not n36061 ; n36061_not
g53884 not n42505 ; n42505_not
g53885 not n41641 ; n41641_not
g53886 not n16702 ; n16702_not
g53887 not n26062 ; n26062_not
g53888 not n15334 ; n15334_not
g53889 not n41803 ; n41803_not
g53890 not n26071 ; n26071_not
g53891 not n15613 ; n15613_not
g53892 not n41380 ; n41380_not
g53893 not n33271 ; n33271_not
g53894 not n33334 ; n33334_not
g53895 not n44440 ; n44440_not
g53896 not n16351 ; n16351_not
g53897 not n16036 ; n16036_not
g53898 not n27007 ; n27007_not
g53899 not n15019 ; n15019_not
g53900 not n16234 ; n16234_not
g53901 not n26701 ; n26701_not
g53902 not n27223 ; n27223_not
g53903 not n16135 ; n16135_not
g53904 not n27115 ; n27115_not
g53905 not n15028 ; n15028_not
g53906 not n16225 ; n16225_not
g53907 not n16126 ; n16126_not
g53908 not n41326 ; n41326_not
g53909 not n16162 ; n16162_not
g53910 not n24910 ; n24910_not
g53911 not n16018 ; n16018_not
g53912 not n24901 ; n24901_not
g53913 not n15901 ; n15901_not
g53914 not n16405 ; n16405_not
g53915 not n18052 ; n18052_not
g53916 not n34531 ; n34531_not
g53917 not n27232 ; n27232_not
g53918 not n33235 ; n33235_not
g53919 not n16153 ; n16153_not
g53920 not n34351 ; n34351_not
g53921 not n34315 ; n34315_not
g53922 not n36214 ; n36214_not
g53923 not n34720 ; n34720_not
g53924 not n10681 ; n10681_not
g53925 not n34450 ; n34450_not
g53926 not n41263 ; n41263_not
g53927 not n16072 ; n16072_not
g53928 not n27205 ; n27205_not
g53929 not n16063 ; n16063_not
g53930 not n10384 ; n10384_not
g53931 not n47311 ; n47311_not
g53932 not n27160 ; n27160_not
g53933 not n16261 ; n16261_not
g53934 not n16315 ; n16315_not
g53935 not n27214 ; n27214_not
g53936 not n41308 ; n41308_not
g53937 not n10591 ; n10591_not
g53938 not n10555 ; n10555_not
g53939 not n42721 ; n42721_not
g53940 not n40309 ; n40309_not
g53941 not n16054 ; n16054_not
g53942 not n36223 ; n36223_not
g53943 not n34540 ; n34540_not
g53944 not n41290 ; n41290_not
g53945 not n18016 ; n18016_not
g53946 not n16333 ; n16333_not
g53947 not n36205 ; n36205_not
g53948 not n42730 ; n42730_not
g53949 not n34612 ; n34612_not
g53950 not n34504 ; n34504_not
g53951 not n36313 ; n36313_not
g53952 not n34522 ; n34522_not
g53953 not n18061 ; n18061_not
g53954 not n27034 ; n27034_not
g53955 not n27061 ; n27061_not
g53956 not n25027 ; n25027_not
g53957 not n36322 ; n36322_not
g53958 not n15073 ; n15073_not
g53959 not n42109 ; n42109_not
g53960 not n41344 ; n41344_not
g53961 not n35044 ; n35044_not
g53962 not n41236 ; n41236_not
g53963 not n20069 ; n20069_not
g53964 not n11366 ; n11366_not
g53965 not n34604 ; n34604_not
g53966 not n27161 ; n27161_not
g53967 not n30266 ; n30266_not
g53968 not n13175 ; n13175_not
g53969 not n31850 ; n31850_not
g53970 not n27152 ; n27152_not
g53971 not n43730 ; n43730_not
g53972 not n11384 ; n11384_not
g53973 not n16253 ; n16253_not
g53974 not n27800 ; n27800_not
g53975 not n15470 ; n15470_not
g53976 not n42506 ; n42506_not
g53977 not n13148 ; n13148_not
g53978 not n34028 ; n34028_not
g53979 not n11627 ; n11627_not
g53980 not n19142 ; n19142_not
g53981 not n20078 ; n20078_not
g53982 not n43523 ; n43523_not
g53983 not n15614 ; n15614_not
g53984 not n22490 ; n22490_not
g53985 not n10943 ; n10943_not
g53986 not n22445 ; n22445_not
g53987 not n30275 ; n30275_not
g53988 not n31265 ; n31265_not
g53989 not n21554 ; n21554_not
g53990 not n41813 ; n41813_not
g53991 not n20096 ; n20096_not
g53992 not n21455 ; n21455_not
g53993 not n13274 ; n13274_not
g53994 not n47204 ; n47204_not
g53995 not n15461 ; n15461_not
g53996 not n10592 ; n10592_not
g53997 not n17054 ; n17054_not
g53998 not n31373 ; n31373_not
g53999 not n33902 ; n33902_not
g54000 not n48302 ; n48302_not
g54001 not n17117 ; n17117_not
g54002 not n10088 ; n10088_not
g54003 not n35351 ; n35351_not
g54004 not n13256 ; n13256_not
g54005 not n13544 ; n13544_not
g54006 not n27134 ; n27134_not
g54007 not n17612 ; n17612_not
g54008 not n10907 ; n10907_not
g54009 not n38231 ; n38231_not
g54010 not n27143 ; n27143_not
g54011 not n22364 ; n22364_not
g54012 not n13238 ; n13238_not
g54013 not n26045 ; n26045_not
g54014 not n35630 ; n35630_not
g54015 not n31274 ; n31274_not
g54016 not n38510 ; n38510_not
g54017 not n17243 ; n17243_not
g54018 not n17027 ; n17027_not
g54019 not n30248 ; n30248_not
g54020 not n26054 ; n26054_not
g54021 not n47510 ; n47510_not
g54022 not n30257 ; n30257_not
g54023 not n20168 ; n20168_not
g54024 not n34514 ; n34514_not
g54025 not n42443 ; n42443_not
g54026 not n13571 ; n13571_not
g54027 not n12950 ; n12950_not
g54028 not n16631 ; n16631_not
g54029 not n31715 ; n31715_not
g54030 not n16721 ; n16721_not
g54031 not n40049 ; n40049_not
g54032 not n20177 ; n20177_not
g54033 not n30383 ; n30383_not
g54034 not n12941 ; n12941_not
g54035 not n21257 ; n21257_not
g54036 not n31724 ; n31724_not
g54037 not n33641 ; n33641_not
g54038 not n27710 ; n27710_not
g54039 not n49013 ; n49013_not
g54040 not n34703 ; n34703_not
g54041 not n38222 ; n38222_not
g54042 not n26135 ; n26135_not
g54043 not n12923 ; n12923_not
g54044 not n34091 ; n34091_not
g54045 not n20195 ; n20195_not
g54046 not n12680 ; n12680_not
g54047 not n45260 ; n45260_not
g54048 not n44207 ; n44207_not
g54049 not n16910 ; n16910_not
g54050 not n46232 ; n46232_not
g54051 not n22409 ; n22409_not
g54052 not n15623 ; n15623_not
g54053 not n45206 ; n45206_not
g54054 not n22481 ; n22481_not
g54055 not n16280 ; n16280_not
g54056 not n26072 ; n26072_not
g54057 not n17270 ; n17270_not
g54058 not n11357 ; n11357_not
g54059 not n41822 ; n41822_not
g54060 not n39041 ; n39041_not
g54061 not n15632 ; n15632_not
g54062 not n13058 ; n13058_not
g54063 not n30293 ; n30293_not
g54064 not n43541 ; n43541_not
g54065 not n35342 ; n35342_not
g54066 not n26081 ; n26081_not
g54067 not n34613 ; n34613_not
g54068 not n10961 ; n10961_not
g54069 not n12905 ; n12905_not
g54070 not n31913 ; n31913_not
g54071 not n45251 ; n45251_not
g54072 not n21446 ; n21446_not
g54073 not n41831 ; n41831_not
g54074 not n21284 ; n21284_not
g54075 not n20159 ; n20159_not
g54076 not n31382 ; n31382_not
g54077 not n11654 ; n11654_not
g54078 not n23129 ; n23129_not
g54079 not n16082 ; n16082_not
g54080 not n15650 ; n15650_not
g54081 not n22814 ; n22814_not
g54082 not n37511 ; n37511_not
g54083 not n27026 ; n27026_not
g54084 not n35423 ; n35423_not
g54085 not n37520 ; n37520_not
g54086 not n22760 ; n22760_not
g54087 not n22724 ; n22724_not
g54088 not n22742 ; n22742_not
g54089 not n31328 ; n31328_not
g54090 not n30095 ; n30095_not
g54091 not n39410 ; n39410_not
g54092 not n44144 ; n44144_not
g54093 not n16172 ; n16172_not
g54094 not n35513 ; n35513_not
g54095 not n43433 ; n43433_not
g54096 not n15830 ; n15830_not
g54097 not n39401 ; n39401_not
g54098 not n23066 ; n23066_not
g54099 not n11519 ; n11519_not
g54100 not n16136 ; n16136_not
g54101 not n42533 ; n42533_not
g54102 not n37313 ; n37313_not
g54103 not n13391 ; n13391_not
g54104 not n21473 ; n21473_not
g54105 not n48320 ; n48320_not
g54106 not n28007 ; n28007_not
g54107 not n39320 ; n39320_not
g54108 not n31805 ; n31805_not
g54109 not n17207 ; n17207_not
g54110 not n34505 ; n34505_not
g54111 not n46430 ; n46430_not
g54112 not n25901 ; n25901_not
g54113 not n41057 ; n41057_not
g54114 not n27035 ; n27035_not
g54115 not n25910 ; n25910_not
g54116 not n21482 ; n21482_not
g54117 not n35414 ; n35414_not
g54118 not n13436 ; n13436_not
g54119 not n46421 ; n46421_not
g54120 not n37331 ; n37331_not
g54121 not n37340 ; n37340_not
g54122 not n17144 ; n17144_not
g54123 not n35450 ; n35450_not
g54124 not n37403 ; n37403_not
g54125 not n42551 ; n42551_not
g54126 not n28034 ; n28034_not
g54127 not n37430 ; n37430_not
g54128 not n42524 ; n42524_not
g54129 not n35432 ; n35432_not
g54130 not n37421 ; n37421_not
g54131 not n38240 ; n38240_not
g54132 not n40931 ; n40931_not
g54133 not n27107 ; n27107_not
g54134 not n28052 ; n28052_not
g54135 not n22922 ; n22922_not
g54136 not n17162 ; n17162_not
g54137 not n43442 ; n43442_not
g54138 not n22940 ; n22940_not
g54139 not n39302 ; n39302_not
g54140 not n35504 ; n35504_not
g54141 not n21419 ; n21419_not
g54142 not n46322 ; n46322_not
g54143 not n26018 ; n26018_not
g54144 not n13490 ; n13490_not
g54145 not n31751 ; n31751_not
g54146 not n21356 ; n21356_not
g54147 not n10880 ; n10880_not
g54148 not n13508 ; n13508_not
g54149 not n45170 ; n45170_not
g54150 not n11573 ; n11573_not
g54151 not n27125 ; n27125_not
g54152 not n22553 ; n22553_not
g54153 not n39140 ; n39140_not
g54154 not n33650 ; n33650_not
g54155 not n31490 ; n31490_not
g54156 not n16118 ; n16118_not
g54157 not n17135 ; n17135_not
g54158 not n21527 ; n21527_not
g54159 not n39131 ; n39131_not
g54160 not n15560 ; n15560_not
g54161 not n46304 ; n46304_not
g54162 not n31742 ; n31742_not
g54163 not n28070 ; n28070_not
g54164 not n13526 ; n13526_not
g54165 not n21347 ; n21347_not
g54166 not n17072 ; n17072_not
g54167 not n17126 ; n17126_not
g54168 not n15812 ; n15812_not
g54169 not n42182 ; n42182_not
g54170 not n44360 ; n44360_not
g54171 not n21338 ; n21338_not
g54172 not n33704 ; n33704_not
g54173 not n27017 ; n27017_not
g54174 not n46340 ; n46340_not
g54175 not n11537 ; n11537_not
g54176 not n13364 ; n13364_not
g54177 not n21518 ; n21518_not
g54178 not n22643 ; n22643_not
g54179 not n22661 ; n22661_not
g54180 not n13481 ; n13481_not
g54181 not n15542 ; n15542_not
g54182 not n40652 ; n40652_not
g54183 not n23084 ; n23084_not
g54184 not n10439 ; n10439_not
g54185 not n11456 ; n11456_not
g54186 not n37304 ; n37304_not
g54187 not n13337 ; n13337_not
g54188 not n13319 ; n13319_not
g54189 not n35126 ; n35126_not
g54190 not n48311 ; n48311_not
g54191 not n15551 ; n15551_not
g54192 not n16127 ; n16127_not
g54193 not n22607 ; n22607_not
g54194 not n26009 ; n26009_not
g54195 not n39212 ; n39212_not
g54196 not n30158 ; n30158_not
g54197 not n13328 ; n13328_not
g54198 not n31409 ; n31409_not
g54199 not n43451 ; n43451_not
g54200 not n22616 ; n22616_not
g54201 not n39230 ; n39230_not
g54202 not n17090 ; n17090_not
g54203 not n30149 ; n30149_not
g54204 not n30923 ; n30923_not
g54205 not n31436 ; n31436_not
g54206 not n21095 ; n21095_not
g54207 not n12266 ; n12266_not
g54208 not n26360 ; n26360_not
g54209 not n38501 ; n38501_not
g54210 not n42119 ; n42119_not
g54211 not n46052 ; n46052_not
g54212 not n16019 ; n16019_not
g54213 not n30905 ; n30905_not
g54214 not n27413 ; n27413_not
g54215 not n26441 ; n26441_not
g54216 not n31535 ; n31535_not
g54217 not n30824 ; n30824_not
g54218 not n42056 ; n42056_not
g54219 not n31553 ; n31553_not
g54220 not n20807 ; n20807_not
g54221 not n21716 ; n21716_not
g54222 not n11951 ; n11951_not
g54223 not n42290 ; n42290_not
g54224 not n38420 ; n38420_not
g54225 not n21950 ; n21950_not
g54226 not n26522 ; n26522_not
g54227 not n15902 ; n15902_not
g54228 not n11942 ; n11942_not
g54229 not n41840 ; n41840_not
g54230 not n16550 ; n16550_not
g54231 not n21077 ; n21077_not
g54232 not n26513 ; n26513_not
g54233 not n27404 ; n27404_not
g54234 not n20762 ; n20762_not
g54235 not n38024 ; n38024_not
g54236 not n30932 ; n30932_not
g54237 not n27332 ; n27332_not
g54238 not n16622 ; n16622_not
g54239 not n20654 ; n20654_not
g54240 not n21662 ; n21662_not
g54241 not n26414 ; n26414_not
g54242 not n20645 ; n20645_not
g54243 not n11294 ; n11294_not
g54244 not n22094 ; n22094_not
g54245 not n20636 ; n20636_not
g54246 not n26612 ; n26612_not
g54247 not n11870 ; n11870_not
g54248 not n11681 ; n11681_not
g54249 not n46106 ; n46106_not
g54250 not n26711 ; n26711_not
g54251 not n42128 ; n42128_not
g54252 not n26720 ; n26720_not
g54253 not n27422 ; n27422_not
g54254 not n27431 ; n27431_not
g54255 not n42038 ; n42038_not
g54256 not n46070 ; n46070_not
g54257 not n15740 ; n15740_not
g54258 not n17234 ; n17234_not
g54259 not n20690 ; n20690_not
g54260 not n12338 ; n12338_not
g54261 not n35207 ; n35207_not
g54262 not n16604 ; n16604_not
g54263 not n16028 ; n16028_not
g54264 not n30851 ; n30851_not
g54265 not n42029 ; n42029_not
g54266 not n16613 ; n16613_not
g54267 not n34280 ; n34280_not
g54268 not n20663 ; n20663_not
g54269 not n31562 ; n31562_not
g54270 not n16316 ; n16316_not
g54271 not n42263 ; n42263_not
g54272 not n12068 ; n12068_not
g54273 not n10538 ; n10538_not
g54274 not n21725 ; n21725_not
g54275 not n31463 ; n31463_not
g54276 not n20924 ; n20924_not
g54277 not n27314 ; n27314_not
g54278 not n35063 ; n35063_not
g54279 not n42092 ; n42092_not
g54280 not n17018 ; n17018_not
g54281 not n21824 ; n21824_not
g54282 not n12077 ; n12077_not
g54283 not n12086 ; n12086_not
g54284 not n12095 ; n12095_not
g54285 not n42137 ; n42137_not
g54286 not n42272 ; n42272_not
g54287 not n38321 ; n38321_not
g54288 not n38132 ; n38132_not
g54289 not n10817 ; n10817_not
g54290 not n31058 ; n31058_not
g54291 not n38141 ; n38141_not
g54292 not n42236 ; n42236_not
g54293 not n16406 ; n16406_not
g54294 not n26630 ; n26630_not
g54295 not n38330 ; n38330_not
g54296 not n38114 ; n38114_not
g54297 not n16451 ; n16451_not
g54298 not n42254 ; n42254_not
g54299 not n21815 ; n21815_not
g54300 not n35072 ; n35072_not
g54301 not n20843 ; n20843_not
g54302 not n16514 ; n16514_not
g54303 not n44018 ; n44018_not
g54304 not n20753 ; n20753_not
g54305 not n42209 ; n42209_not
g54306 not n42218 ; n42218_not
g54307 not n16523 ; n16523_not
g54308 not n12185 ; n12185_not
g54309 not n31508 ; n31508_not
g54310 not n11159 ; n11159_not
g54311 not n44027 ; n44027_not
g54312 not n31085 ; n31085_not
g54313 not n21059 ; n21059_not
g54314 not n20816 ; n20816_not
g54315 not n15911 ; n15911_not
g54316 not n21932 ; n21932_not
g54317 not n21833 ; n21833_not
g54318 not n31472 ; n31472_not
g54319 not n31076 ; n31076_not
g54320 not n20906 ; n20906_not
g54321 not n46007 ; n46007_not
g54322 not n35117 ; n35117_not
g54323 not n21851 ; n21851_not
g54324 not n34352 ; n34352_not
g54325 not n11177 ; n11177_not
g54326 not n46016 ; n46016_not
g54327 not n10295 ; n10295_not
g54328 not n27242 ; n27242_not
g54329 not n16505 ; n16505_not
g54330 not n26540 ; n26540_not
g54331 not n12149 ; n12149_not
g54332 not n20375 ; n20375_not
g54333 not n27602 ; n27602_not
g54334 not n30563 ; n30563_not
g54335 not n42434 ; n42434_not
g54336 not n27611 ; n27611_not
g54337 not n20249 ; n20249_not
g54338 not n12734 ; n12734_not
g54339 not n11762 ; n11762_not
g54340 not n26243 ; n26243_not
g54341 not n42902 ; n42902_not
g54342 not n44090 ; n44090_not
g54343 not n34730 ; n34730_not
g54344 not n20348 ; n20348_not
g54345 not n31238 ; n31238_not
g54346 not n26234 ; n26234_not
g54347 not n11744 ; n11744_not
g54348 not n34163 ; n34163_not
g54349 not n12662 ; n12662_not
g54350 not n20384 ; n20384_not
g54351 not n30626 ; n30626_not
g54352 not n26261 ; n26261_not
g54353 not n21194 ; n21194_not
g54354 not n30617 ; n30617_not
g54355 not n12707 ; n12707_not
g54356 not n30608 ; n30608_not
g54357 not n31661 ; n31661_not
g54358 not n44072 ; n44072_not
g54359 not n10367 ; n10367_not
g54360 not n34127 ; n34127_not
g54361 not n20267 ; n20267_not
g54362 not n31247 ; n31247_not
g54363 not n34037 ; n34037_not
g54364 not n26180 ; n26180_not
g54365 not n35306 ; n35306_not
g54366 not n26171 ; n26171_not
g54367 not n47420 ; n47420_not
g54368 not n41903 ; n41903_not
g54369 not n30455 ; n30455_not
g54370 not n38213 ; n38213_not
g54371 not n46223 ; n46223_not
g54372 not n21248 ; n21248_not
g54373 not n26153 ; n26153_not
g54374 not n42461 ; n42461_not
g54375 not n12752 ; n12752_not
g54376 not n43703 ; n43703_not
g54377 not n16307 ; n16307_not
g54378 not n30545 ; n30545_not
g54379 not n12770 ; n12770_not
g54380 not n16820 ; n16820_not
g54381 not n41930 ; n41930_not
g54382 not n27620 ; n27620_not
g54383 not n30518 ; n30518_not
g54384 not n43505 ; n43505_not
g54385 not n46214 ; n46214_not
g54386 not n26207 ; n26207_not
g54387 not n30509 ; n30509_not
g54388 not n20285 ; n20285_not
g54389 not n20276 ; n20276_not
g54390 not n43640 ; n43640_not
g54391 not n31184 ; n31184_not
g54392 not n12491 ; n12491_not
g54393 not n44306 ; n44306_not
g54394 not n47411 ; n47411_not
g54395 not n43820 ; n43820_not
g54396 not n20474 ; n20474_not
g54397 not n20546 ; n20546_not
g54398 not n22184 ; n22184_not
g54399 not n17504 ; n17504_not
g54400 not n35243 ; n35243_not
g54401 not n26333 ; n26333_not
g54402 not n11834 ; n11834_not
g54403 not n46160 ; n46160_not
g54404 not n20519 ; n20519_not
g54405 not n11825 ; n11825_not
g54406 not n21167 ; n21167_not
g54407 not n34802 ; n34802_not
g54408 not n12563 ; n12563_not
g54409 not n26405 ; n26405_not
g54410 not n12428 ; n12428_not
g54411 not n20609 ; n20609_not
g54412 not n11852 ; n11852_not
g54413 not n12446 ; n12446_not
g54414 not n46124 ; n46124_not
g54415 not n12464 ; n12464_not
g54416 not n15803 ; n15803_not
g54417 not n20591 ; n20591_not
g54418 not n42362 ; n42362_not
g54419 not n30770 ; n30770_not
g54420 not n30743 ; n30743_not
g54421 not n30752 ; n30752_not
g54422 not n34244 ; n34244_not
g54423 not n16352 ; n16352_not
g54424 not n34226 ; n34226_not
g54425 not n22256 ; n22256_not
g54426 not n35252 ; n35252_not
g54427 not n16730 ; n16730_not
g54428 not n22265 ; n22265_not
g54429 not n42146 ; n42146_not
g54430 not n12626 ; n12626_not
g54431 not n27512 ; n27512_not
g54432 not n30644 ; n30644_not
g54433 not n12644 ; n12644_not
g54434 not n44315 ; n44315_not
g54435 not n26810 ; n26810_not
g54436 not n47033 ; n47033_not
g54437 not n34442 ; n34442_not
g54438 not n22283 ; n22283_not
g54439 not n22274 ; n22274_not
g54440 not n47240 ; n47240_not
g54441 not n30707 ; n30707_not
g54442 not n16712 ; n16712_not
g54443 not n43811 ; n43811_not
g54444 not n12581 ; n12581_not
g54445 not n27215 ; n27215_not
g54446 not n22229 ; n22229_not
g54447 not n12590 ; n12590_not
g54448 not n10628 ; n10628_not
g54449 not n22238 ; n22238_not
g54450 not n42407 ; n42407_not
g54451 not n30680 ; n30680_not
g54452 not n34172 ; n34172_not
g54453 not n16334 ; n16334_not
g54454 not n30662 ; n30662_not
g54455 not n32444 ; n32444_not
g54456 not n14930 ; n14930_not
g54457 not n15119 ; n15119_not
g54458 not n40418 ; n40418_not
g54459 not n24506 ; n24506_not
g54460 not n41444 ; n41444_not
g54461 not n14075 ; n14075_not
g54462 not n14066 ; n14066_not
g54463 not n25271 ; n25271_not
g54464 not n10781 ; n10781_not
g54465 not n10673 ; n10673_not
g54466 not n41129 ; n41129_not
g54467 not n10718 ; n10718_not
g54468 not n14705 ; n14705_not
g54469 not n32426 ; n32426_not
g54470 not n18134 ; n18134_not
g54471 not n10682 ; n10682_not
g54472 not n32417 ; n32417_not
g54473 not n14714 ; n14714_not
g54474 not n43172 ; n43172_not
g54475 not n18332 ; n18332_not
g54476 not n14435 ; n14435_not
g54477 not n25307 ; n25307_not
g54478 not n36044 ; n36044_not
g54479 not n10277 ; n10277_not
g54480 not n24533 ; n24533_not
g54481 not n42731 ; n42731_not
g54482 not n19034 ; n19034_not
g54483 not n23642 ; n23642_not
g54484 not n40436 ; n40436_not
g54485 not n41390 ; n41390_not
g54486 not n17630 ; n17630_not
g54487 not n32903 ; n32903_not
g54488 not n41093 ; n41093_not
g54489 not n33524 ; n33524_not
g54490 not n43055 ; n43055_not
g54491 not n29420 ; n29420_not
g54492 not n40706 ; n40706_not
g54493 not n25127 ; n25127_not
g54494 not n33542 ; n33542_not
g54495 not n33344 ; n33344_not
g54496 not n23606 ; n23606_not
g54497 not n25253 ; n25253_not
g54498 not n17603 ; n17603_not
g54499 not n43163 ; n43163_not
g54500 not n15308 ; n15308_not
g54501 not n10772 ; n10772_not
g54502 not n42632 ; n42632_not
g54503 not n10664 ; n10664_not
g54504 not n43046 ; n43046_not
g54505 not n33029 ; n33029_not
g54506 not n41606 ; n41606_not
g54507 not n46700 ; n46700_not
g54508 not n17108 ; n17108_not
g54509 not n19160 ; n19160_not
g54510 not n36062 ; n36062_not
g54511 not n43217 ; n43217_not
g54512 not n25325 ; n25325_not
g54513 not n28430 ; n28430_not
g54514 not n23453 ; n23453_not
g54515 not n10844 ; n10844_not
g54516 not n32363 ; n32363_not
g54517 not n41273 ; n41273_not
g54518 not n43226 ; n43226_not
g54519 not n19214 ; n19214_not
g54520 not n17540 ; n17540_not
g54521 not n32354 ; n32354_not
g54522 not n23426 ; n23426_not
g54523 not n29123 ; n29123_not
g54524 not n10394 ; n10394_not
g54525 not n43235 ; n43235_not
g54526 not n24254 ; n24254_not
g54527 not n14750 ; n14750_not
g54528 not n19232 ; n19232_not
g54529 not n40742 ; n40742_not
g54530 not n33092 ; n33092_not
g54531 not n33317 ; n33317_not
g54532 not n13940 ; n13940_not
g54533 not n41147 ; n41147_not
g54534 not n24038 ; n24038_not
g54535 not n19241 ; n19241_not
g54536 not n23417 ; n23417_not
g54537 not n43181 ; n43181_not
g54538 not n15335 ; n15335_not
g54539 not n36206 ; n36206_not
g54540 not n36071 ; n36071_not
g54541 not n41138 ; n41138_not
g54542 not n14723 ; n14723_not
g54543 not n17324 ; n17324_not
g54544 not n32390 ; n32390_not
g54545 not n25316 ; n25316_not
g54546 not n23903 ; n23903_not
g54547 not n18323 ; n18323_not
g54548 not n40724 ; n40724_not
g54549 not n25118 ; n25118_not
g54550 not n41282 ; n41282_not
g54551 not n18314 ; n18314_not
g54552 not n10826 ; n10826_not
g54553 not n33065 ; n33065_not
g54554 not n23480 ; n23480_not
g54555 not n32624 ; n32624_not
g54556 not n36143 ; n36143_not
g54557 not n23471 ; n23471_not
g54558 not n32615 ; n32615_not
g54559 not n40373 ; n40373_not
g54560 not n18305 ; n18305_not
g54561 not n23462 ; n23462_not
g54562 not n37223 ; n37223_not
g54563 not n40481 ; n40481_not
g54564 not n14237 ; n14237_not
g54565 not n36116 ; n36116_not
g54566 not n17081 ; n17081_not
g54567 not n37025 ; n37025_not
g54568 not n43136 ; n43136_not
g54569 not n15218 ; n15218_not
g54570 not n18602 ; n18602_not
g54571 not n33380 ; n33380_not
g54572 not n44414 ; n44414_not
g54573 not n29330 ; n29330_not
g54574 not n43154 ; n43154_not
g54575 not n14219 ; n14219_not
g54576 not n44603 ; n44603_not
g54577 not n14561 ; n14561_not
g54578 not n15191 ; n15191_not
g54579 not n40562 ; n40562_not
g54580 not n23750 ; n23750_not
g54581 not n24371 ; n24371_not
g54582 not n37016 ; n37016_not
g54583 not n41525 ; n41525_not
g54584 not n40553 ; n40553_not
g54585 not n14507 ; n14507_not
g54586 not n33353 ; n33353_not
g54587 not n28331 ; n28331_not
g54588 not n15038 ; n15038_not
g54589 not n29033 ; n29033_not
g54590 not n33371 ; n33371_not
g54591 not n43073 ; n43073_not
g54592 not n18503 ; n18503_not
g54593 not n43145 ; n43145_not
g54594 not n14291 ; n14291_not
g54595 not n33362 ; n33362_not
g54596 not n25154 ; n25154_not
g54597 not n23840 ; n23840_not
g54598 not n41354 ; n41354_not
g54599 not n32813 ; n32813_not
g54600 not n40634 ; n40634_not
g54601 not n40274 ; n40274_not
g54602 not n29042 ; n29042_not
g54603 not n10529 ; n10529_not
g54604 not n18422 ; n18422_not
g54605 not n33452 ; n33452_not
g54606 not n36620 ; n36620_not
g54607 not n32570 ; n32570_not
g54608 not n15209 ; n15209_not
g54609 not n28502 ; n28502_not
g54610 not n40616 ; n40616_not
g54611 not n14516 ; n14516_not
g54612 not n28250 ; n28250_not
g54613 not n24353 ; n24353_not
g54614 not n17711 ; n17711_not
g54615 not n23741 ; n23741_not
g54616 not n32534 ; n32534_not
g54617 not n25172 ; n25172_not
g54618 not n14633 ; n14633_not
g54619 not n36701 ; n36701_not
g54620 not n24452 ; n24452_not
g54621 not n23651 ; n23651_not
g54622 not n15254 ; n15254_not
g54623 not n28304 ; n28304_not
g54624 not n24218 ; n24218_not
g54625 not n15047 ; n15047_not
g54626 not n29006 ; n29006_not
g54627 not n28520 ; n28520_not
g54628 not n15272 ; n15272_not
g54629 not n41471 ; n41471_not
g54630 not n15281 ; n15281_not
g54631 not n19016 ; n19016_not
g54632 not n44612 ; n44612_not
g54633 not n14138 ; n14138_not
g54634 not n14651 ; n14651_not
g54635 not n10754 ; n10754_not
g54636 not n37007 ; n37007_not
g54637 not n32480 ; n32480_not
g54638 not n24461 ; n24461_not
g54639 not n40382 ; n40382_not
g54640 not n23921 ; n23921_not
g54641 not n19025 ; n19025_not
g54642 not n14660 ; n14660_not
g54643 not n37142 ; n37142_not
g54644 not n24290 ; n24290_not
g54645 not n28223 ; n28223_not
g54646 not n24281 ; n24281_not
g54647 not n29240 ; n29240_not
g54648 not n48104 ; n48104_not
g54649 not n24308 ; n24308_not
g54650 not n14084 ; n14084_not
g54651 not n37106 ; n37106_not
g54652 not n14192 ; n14192_not
g54653 not n14624 ; n14624_not
g54654 not n47114 ; n47114_not
g54655 not n23912 ; n23912_not
g54656 not n40517 ; n40517_not
g54657 not n17900 ; n17900_not
g54658 not n14174 ; n14174_not
g54659 not n25208 ; n25208_not
g54660 not n41480 ; n41480_not
g54661 not n14336 ; n14336_not
g54662 not n40508 ; n40508_not
g54663 not n24425 ; n24425_not
g54664 not n40490 ; n40490_not
g54665 not n41561 ; n41561_not
g54666 not n18431 ; n18431_not
g54667 not n15065 ; n15065_not
g54668 not n14444 ; n14444_not
g54669 not n24443 ; n24443_not
g54670 not n40472 ; n40472_not
g54671 not n29402 ; n29402_not
g54672 not n37133 ; n37133_not
g54673 not n14921 ; n14921_not
g54674 not n13751 ; n13751_not
g54675 not n23264 ; n23264_not
g54676 not n32192 ; n32192_not
g54677 not n13760 ; n13760_not
g54678 not n41723 ; n41723_not
g54679 not n18026 ; n18026_not
g54680 not n36242 ; n36242_not
g54681 not n18035 ; n18035_not
g54682 not n44720 ; n44720_not
g54683 not n18620 ; n18620_not
g54684 not n14912 ; n14912_not
g54685 not n48221 ; n48221_not
g54686 not n19430 ; n19430_not
g54687 not n23246 ; n23246_not
g54688 not n24740 ; n24740_not
g54689 not n32174 ; n32174_not
g54690 not n17045 ; n17045_not
g54691 not n47150 ; n47150_not
g54692 not n42335 ; n42335_not
g54693 not n25343 ; n25343_not
g54694 not n32165 ; n32165_not
g54695 not n17351 ; n17351_not
g54696 not n32660 ; n32660_not
g54697 not n15425 ; n15425_not
g54698 not n24155 ; n24155_not
g54699 not n33164 ; n33164_not
g54700 not n32219 ; n32219_not
g54701 not n47015 ; n47015_not
g54702 not n42812 ; n42812_not
g54703 not n43325 ; n43325_not
g54704 not n41417 ; n41417_not
g54705 not n17450 ; n17450_not
g54706 not n32651 ; n32651_not
g54707 not n43406 ; n43406_not
g54708 not n36233 ; n36233_not
g54709 not n17441 ; n17441_not
g54710 not n33173 ; n33173_not
g54711 not n25334 ; n25334_not
g54712 not n25730 ; n25730_not
g54713 not n40238 ; n40238_not
g54714 not n40805 ; n40805_not
g54715 not n24119 ; n24119_not
g54716 not n28133 ; n28133_not
g54717 not n16811 ; n16811_not
g54718 not n10691 ; n10691_not
g54719 not n15416 ; n15416_not
g54720 not n10853 ; n10853_not
g54721 not n43343 ; n43343_not
g54722 not n25604 ; n25604_not
g54723 not n32714 ; n32714_not
g54724 not n10862 ; n10862_not
g54725 not n48212 ; n48212_not
g54726 not n28700 ; n28700_not
g54727 not n25082 ; n25082_not
g54728 not n42803 ; n42803_not
g54729 not n13670 ; n13670_not
g54730 not n14462 ; n14462_not
g54731 not n13661 ; n13661_not
g54732 not n18116 ; n18116_not
g54733 not n40148 ; n40148_not
g54734 not n14840 ; n14840_not
g54735 not n10196 ; n10196_not
g54736 not n25640 ; n25640_not
g54737 not n14741 ; n14741_not
g54738 not n32066 ; n32066_not
g54739 not n35810 ; n35810_not
g54740 not n35801 ; n35801_not
g54741 not n23165 ; n23165_not
g54742 not n33191 ; n33191_not
g54743 not n23237 ; n23237_not
g54744 not n24164 ; n24164_not
g54745 not n29141 ; n29141_not
g54746 not n32039 ; n32039_not
g54747 not n43352 ; n43352_not
g54748 not n29150 ; n29150_not
g54749 not n13733 ; n13733_not
g54750 not n40247 ; n40247_not
g54751 not n25550 ; n25550_not
g54752 not n18143 ; n18143_not
g54753 not n25703 ; n25703_not
g54754 not n24821 ; n24821_not
g54755 not n33245 ; n33245_not
g54756 not n19502 ; n19502_not
g54757 not n13724 ; n13724_not
g54758 not n10709 ; n10709_not
g54759 not n32138 ; n32138_not
g54760 not n23219 ; n23219_not
g54761 not n43370 ; n43370_not
g54762 not n36350 ; n36350_not
g54763 not n33128 ; n33128_not
g54764 not n41237 ; n41237_not
g54765 not n17306 ; n17306_not
g54766 not n41156 ; n41156_not
g54767 not n32255 ; n32255_not
g54768 not n36170 ; n36170_not
g54769 not n23372 ; n23372_not
g54770 not n18701 ; n18701_not
g54771 not n32282 ; n32282_not
g54772 not n15353 ; n15353_not
g54773 not n25406 ; n25406_not
g54774 not n33137 ; n33137_not
g54775 not n24605 ; n24605_not
g54776 not n17405 ; n17405_not
g54777 not n19322 ; n19322_not
g54778 not n28403 ; n28403_not
g54779 not n14372 ; n14372_not
g54780 not n24614 ; n24614_not
g54781 not n41255 ; n41255_not
g54782 not n41048 ; n41048_not
g54783 not n43127 ; n43127_not
g54784 not n36026 ; n36026_not
g54785 not n46520 ; n46520_not
g54786 not n19250 ; n19250_not
g54787 not n23408 ; n23408_not
g54788 not n41264 ; n41264_not
g54789 not n48041 ; n48041_not
g54790 not n32336 ; n32336_not
g54791 not n37232 ; n37232_not
g54792 not n32633 ; n32633_not
g54793 not n14390 ; n14390_not
g54794 not n17522 ; n17522_not
g54795 not n33119 ; n33119_not
g54796 not n24146 ; n24146_not
g54797 not n23381 ; n23381_not
g54798 not n32327 ; n32327_not
g54799 not n18260 ; n18260_not
g54800 not n41651 ; n41651_not
g54801 not n10646 ; n10646_not
g54802 not n29600 ; n29600_not
g54803 not n17513 ; n17513_not
g54804 not n37241 ; n37241_not
g54805 not n32642 ; n32642_not
g54806 not n43271 ; n43271_not
g54807 not n48113 ; n48113_not
g54808 not n42515 ; n42515_not
g54809 not n33281 ; n33281_not
g54810 not n14417 ; n14417_not
g54811 not n13823 ; n13823_not
g54812 not n28601 ; n28601_not
g54813 not n28610 ; n28610_not
g54814 not n32228 ; n32228_not
g54815 not n41228 ; n41228_not
g54816 not n24092 ; n24092_not
g54817 not n18224 ; n18224_not
g54818 not n13814 ; n13814_not
g54819 not n29132 ; n29132_not
g54820 not n18062 ; n18062_not
g54821 not n41174 ; n41174_not
g54822 not n25064 ; n25064_not
g54823 not n28412 ; n28412_not
g54824 not n13805 ; n13805_not
g54825 not n32723 ; n32723_not
g54826 not n40067 ; n40067_not
g54827 not n15380 ; n15380_not
g54828 not n42830 ; n42830_not
g54829 not n13562 ; n13562_not
g54830 not n10259 ; n10259_not
g54831 not n42821 ; n42821_not
g54832 not n44711 ; n44711_not
g54833 not n33227 ; n33227_not
g54834 not n31940 ; n31940_not
g54835 not n23345 ; n23345_not
g54836 not n28151 ; n28151_not
g54837 not n24065 ; n24065_not
g54838 not n24227 ; n24227_not
g54839 not n25109 ; n25109_not
g54840 not n19331 ; n19331_not
g54841 not n19601 ; n19601_not
g54842 not n40913 ; n40913_not
g54843 not n23318 ; n23318_not
g54844 not n18233 ; n18233_not
g54845 not n41408 ; n41408_not
g54846 not n23327 ; n23327_not
g54847 not n13715 ; n13715_not
g54848 not n13832 ; n13832_not
g54849 not n10376 ; n10376_not
g54850 not n40292 ; n40292_not
g54851 not n43307 ; n43307_not
g54852 not n21942 ; n21942_not
g54853 not n29160 ; n29160_not
g54854 not n25038 ; n25038_not
g54855 not n17046 ; n17046_not
g54856 not n36162 ; n36162_not
g54857 not n29052 ; n29052_not
g54858 not n27333 ; n27333_not
g54859 not n32733 ; n32733_not
g54860 not n24264 ; n24264_not
g54861 not n38070 ; n38070_not
g54862 not n38106 ; n38106_not
g54863 not n24219 ; n24219_not
g54864 not n35127 ; n35127_not
g54865 not n46017 ; n46017_not
g54866 not n36720 ; n36720_not
g54867 not n21861 ; n21861_not
g54868 not n34344 ; n34344_not
g54869 not n29115 ; n29115_not
g54870 not n31482 ; n31482_not
g54871 not n25065 ; n25065_not
g54872 not n21870 ; n21870_not
g54873 not n25056 ; n25056_not
g54874 not n36711 ; n36711_not
g54875 not n35082 ; n35082_not
g54876 not n35091 ; n35091_not
g54877 not n32814 ; n32814_not
g54878 not n25047 ; n25047_not
g54879 not n29070 ; n29070_not
g54880 not n21924 ; n21924_not
g54881 not n30951 ; n30951_not
g54882 not n33390 ; n33390_not
g54883 not n26316 ; n26316_not
g54884 not n21807 ; n21807_not
g54885 not n24174 ; n24174_not
g54886 not n36810 ; n36810_not
g54887 not n24291 ; n24291_not
g54888 not n30870 ; n30870_not
g54889 not n21915 ; n21915_not
g54890 not n24273 ; n24273_not
g54891 not n32742 ; n32742_not
g54892 not n21906 ; n21906_not
g54893 not n36171 ; n36171_not
g54894 not n27153 ; n27153_not
g54895 not n21573 ; n21573_not
g54896 not n16533 ; n16533_not
g54897 not n28800 ; n28800_not
g54898 not n24606 ; n24606_not
g54899 not n47304 ; n47304_not
g54900 not n21564 ; n21564_not
g54901 not n31257 ; n31257_not
g54902 not n24624 ; n24624_not
g54903 not n47331 ; n47331_not
g54904 not n33129 ; n33129_not
g54905 not n36504 ; n36504_not
g54906 not n49014 ; n49014_not
g54907 not n34605 ; n34605_not
g54908 not n33156 ; n33156_not
g54909 not n33147 ; n33147_not
g54910 not n33084 ; n33084_not
g54911 not n34812 ; n34812_not
g54912 not n48042 ; n48042_not
g54913 not n24552 ; n24552_not
g54914 not n26802 ; n26802_not
g54915 not n36225 ; n36225_not
g54916 not n33309 ; n33309_not
g54917 not n34452 ; n34452_not
g54918 not n36540 ; n36540_not
g54919 not n34461 ; n34461_not
g54920 not n48033 ; n48033_not
g54921 not n34713 ; n34713_not
g54922 not n26901 ; n26901_not
g54923 not n27171 ; n27171_not
g54924 not n27180 ; n27180_not
g54925 not n26910 ; n26910_not
g54926 not n21582 ; n21582_not
g54927 not n36405 ; n36405_not
g54928 not n24903 ; n24903_not
g54929 not n28710 ; n28710_not
g54930 not n27108 ; n27108_not
g54931 not n33237 ; n33237_not
g54932 not n17037 ; n17037_not
g54933 not n21492 ; n21492_not
g54934 not n34407 ; n34407_not
g54935 not n36342 ; n36342_not
g54936 not n31392 ; n31392_not
g54937 not n21483 ; n21483_not
g54938 not n24831 ; n24831_not
g54939 not n27036 ; n27036_not
g54940 not n21465 ; n21465_not
g54941 not n33219 ; n33219_not
g54942 not n36324 ; n36324_not
g54943 not n33228 ; n33228_not
g54944 not n28611 ; n28611_not
g54945 not n24642 ; n24642_not
g54946 not n27144 ; n27144_not
g54947 not n24651 ; n24651_not
g54948 not n33273 ; n33273_not
g54949 not n33174 ; n33174_not
g54950 not n24660 ; n24660_not
g54951 not n31293 ; n31293_not
g54952 not n47034 ; n47034_not
g54953 not n47043 ; n47043_not
g54954 not n17154 ; n17154_not
g54955 not n36423 ; n36423_not
g54956 not n47052 ; n47052_not
g54957 not n24750 ; n24750_not
g54958 not n49050 ; n49050_not
g54959 not n24912 ; n24912_not
g54960 not n34533 ; n34533_not
g54961 not n16641 ; n16641_not
g54962 not n26631 ; n26631_not
g54963 not n24381 ; n24381_not
g54964 not n24390 ; n24390_not
g54965 not n36441 ; n36441_not
g54966 not n38151 ; n38151_not
g54967 not n35055 ; n35055_not
g54968 not n29016 ; n29016_not
g54969 not n36180 ; n36180_not
g54970 not n34425 ; n34425_not
g54971 not n33354 ; n33354_not
g54972 not n28512 ; n28512_not
g54973 not n27234 ; n27234_not
g54974 not n28521 ; n28521_not
g54975 not n38052 ; n38052_not
g54976 not n24327 ; n24327_not
g54977 not n34371 ; n34371_not
g54978 not n35064 ; n35064_not
g54979 not n32823 ; n32823_not
g54980 not n29043 ; n29043_not
g54981 not n26622 ; n26622_not
g54982 not n21780 ; n21780_not
g54983 not n24354 ; n24354_not
g54984 not n21771 ; n21771_not
g54985 not n25029 ; n25029_not
g54986 not n29034 ; n29034_not
g54987 not n24363 ; n24363_not
g54988 not n21753 ; n21753_not
g54989 not n17433 ; n17433_not
g54990 not n21744 ; n21744_not
g54991 not n21735 ; n21735_not
g54992 not n34920 ; n34920_not
g54993 not n34434 ; n34434_not
g54994 not n31194 ; n31194_not
g54995 not n31176 ; n31176_not
g54996 not n47241 ; n47241_not
g54997 not n31167 ; n31167_not
g54998 not n33327 ; n33327_not
g54999 not n31428 ; n31428_not
g55000 not n38205 ; n38205_not
g55001 not n34821 ; n34821_not
g55002 not n21618 ; n21618_not
g55003 not n26820 ; n26820_not
g55004 not n36216 ; n36216_not
g55005 not n33318 ; n33318_not
g55006 not n33075 ; n33075_not
g55007 not n32850 ; n32850_not
g55008 not n24471 ; n24471_not
g55009 not n47007 ; n47007_not
g55010 not n21681 ; n21681_not
g55011 not n21672 ; n21672_not
g55012 not n36612 ; n36612_not
g55013 not n21654 ; n21654_not
g55014 not n32913 ; n32913_not
g55015 not n21645 ; n21645_not
g55016 not n31077 ; n31077_not
g55017 not n26703 ; n26703_not
g55018 not n32922 ; n32922_not
g55019 not n31158 ; n31158_not
g55020 not n47106 ; n47106_not
g55021 not n31347 ; n31347_not
g55022 not n24444 ; n24444_not
g55023 not n17631 ; n17631_not
g55024 not n26721 ; n26721_not
g55025 not n22527 ; n22527_not
g55026 not n36036 ; n36036_not
g55027 not n29610 ; n29610_not
g55028 not n16650 ; n16650_not
g55029 not n33813 ; n33813_not
g55030 not n36054 ; n36054_not
g55031 not n33912 ; n33912_not
g55032 not n29601 ; n29601_not
g55033 not n26037 ; n26037_not
g55034 not n23391 ; n23391_not
g55035 not n33921 ; n33921_not
g55036 not n33930 ; n33930_not
g55037 not n26028 ; n26028_not
g55038 not n30249 ; n30249_not
g55039 not n46521 ; n46521_not
g55040 not n29430 ; n29430_not
g55041 not n47214 ; n47214_not
g55042 not n22482 ; n22482_not
g55043 not n26055 ; n26055_not
g55044 not n37620 ; n37620_not
g55045 not n33741 ; n33741_not
g55046 not n33750 ; n33750_not
g55047 not n22626 ; n22626_not
g55048 not n31770 ; n31770_not
g55049 not n48123 ; n48123_not
g55050 not n25452 ; n25452_not
g55051 not n23337 ; n23337_not
g55052 not n46323 ; n46323_not
g55053 not n28143 ; n28143_not
g55054 not n22590 ; n22590_not
g55055 not n22563 ; n22563_not
g55056 not n37251 ; n37251_not
g55057 not n28161 ; n28161_not
g55058 not n32247 ; n32247_not
g55059 not n30195 ; n30195_not
g55060 not n22545 ; n22545_not
g55061 not n22554 ; n22554_not
g55062 not n25407 ; n25407_not
g55063 not n36072 ; n36072_not
g55064 not n26082 ; n26082_not
g55065 not n48510 ; n48510_not
g55066 not n23508 ; n23508_not
g55067 not n34065 ; n34065_not
g55068 not n33552 ; n33552_not
g55069 not n18072 ; n18072_not
g55070 not n29511 ; n29511_not
g55071 not n34074 ; n34074_not
g55072 not n25308 ; n25308_not
g55073 not n29502 ; n29502_not
g55074 not n34056 ; n34056_not
g55075 not n23526 ; n23526_not
g55076 not n22419 ; n22419_not
g55077 not n36081 ; n36081_not
g55078 not n25290 ; n25290_not
g55079 not n47421 ; n47421_not
g55080 not n23544 ; n23544_not
g55081 not n25281 ; n25281_not
g55082 not n25335 ; n25335_not
g55083 not n32346 ; n32346_not
g55084 not n47502 ; n47502_not
g55085 not n23427 ; n23427_not
g55086 not n34038 ; n34038_not
g55087 not n31734 ; n31734_not
g55088 not n34047 ; n34047_not
g55089 not n23445 ; n23445_not
g55090 not n30285 ; n30285_not
g55091 not n33417 ; n33417_not
g55092 not n32382 ; n32382_not
g55093 not n48105 ; n48105_not
g55094 not n37215 ; n37215_not
g55095 not n22455 ; n22455_not
g55096 not n31608 ; n31608_not
g55097 not n23490 ; n23490_not
g55098 not n22446 ; n22446_not
g55099 not n23283 ; n23283_not
g55100 not n37206 ; n37206_not
g55101 not n32067 ; n32067_not
g55102 not n25632 ; n25632_not
g55103 not n10197 ; n10197_not
g55104 not n35541 ; n35541_not
g55105 not n23175 ; n23175_not
g55106 not n25614 ; n25614_not
g55107 not n28053 ; n28053_not
g55108 not n35514 ; n35514_not
g55109 not n35901 ; n35901_not
g55110 not n23193 ; n23193_not
g55111 not n28044 ; n28044_not
g55112 not n35910 ; n35910_not
g55113 not n25560 ; n25560_not
g55114 not n16803 ; n16803_not
g55115 not n32148 ; n32148_not
g55116 not n37341 ; n37341_not
g55117 not n37332 ; n37332_not
g55118 not n37350 ; n37350_not
g55119 not n35703 ; n35703_not
g55120 not n23139 ; n23139_not
g55121 not n23148 ; n23148_not
g55122 not n28080 ; n28080_not
g55123 not n25740 ; n25740_not
g55124 not n35721 ; n35721_not
g55125 not n25731 ; n25731_not
g55126 not n35640 ; n35640_not
g55127 not n31824 ; n31824_not
g55128 not n31905 ; n31905_not
g55129 not n33633 ; n33633_not
g55130 not n35631 ; n35631_not
g55131 not n23157 ; n23157_not
g55132 not n25803 ; n25803_not
g55133 not n35613 ; n35613_not
g55134 not n25704 ; n25704_not
g55135 not n35604 ; n35604_not
g55136 not n28107 ; n28107_not
g55137 not n28071 ; n28071_not
g55138 not n35820 ; n35820_not
g55139 not n35550 ; n35550_not
g55140 not n25506 ; n25506_not
g55141 not n28134 ; n28134_not
g55142 not n22725 ; n22725_not
g55143 not n33624 ; n33624_not
g55144 not n23292 ; n23292_not
g55145 not n48321 ; n48321_not
g55146 not n47142 ; n47142_not
g55147 not n22707 ; n22707_not
g55148 not n35370 ; n35370_not
g55149 not n47133 ; n47133_not
g55150 not n36009 ; n36009_not
g55151 not n22671 ; n22671_not
g55152 not n46332 ; n46332_not
g55153 not n22653 ; n22653_not
g55154 not n47205 ; n47205_not
g55155 not n22644 ; n22644_not
g55156 not n25461 ; n25461_not
g55157 not n22842 ; n22842_not
g55158 not n37161 ; n37161_not
g55159 not n25425 ; n25425_not
g55160 not n22941 ; n22941_not
g55161 not n25551 ; n25551_not
g55162 not n22932 ; n22932_not
g55163 not n22923 ; n22923_not
g55164 not n22905 ; n22905_not
g55165 not n37413 ; n37413_not
g55166 not n25524 ; n25524_not
g55167 not n22815 ; n22815_not
g55168 not n22860 ; n22860_not
g55169 not n22851 ; n22851_not
g55170 not n46404 ; n46404_not
g55171 not n37521 ; n37521_not
g55172 not n23265 ; n23265_not
g55173 not n25515 ; n25515_not
g55174 not n22734 ; n22734_not
g55175 not n32085 ; n32085_not
g55176 not n34236 ; n34236_not
g55177 not n33435 ; n33435_not
g55178 not n30771 ; n30771_not
g55179 not n30654 ; n30654_not
g55180 not n29313 ; n29313_not
g55181 not n34254 ; n34254_not
g55182 not n27270 ; n27270_not
g55183 not n26325 ; n26325_not
g55184 not n26406 ; n26406_not
g55185 not n29232 ; n29232_not
g55186 not n37611 ; n37611_not
g55187 not n25128 ; n25128_not
g55188 not n29304 ; n29304_not
g55189 not n25119 ; n25119_not
g55190 not n30807 ; n30807_not
g55191 not n31590 ; n31590_not
g55192 not n32607 ; n32607_not
g55193 not n46530 ; n46530_not
g55194 not n23841 ; n23841_not
g55195 not n36126 ; n36126_not
g55196 not n33453 ; n33453_not
g55197 not n37035 ; n37035_not
g55198 not n22185 ; n22185_not
g55199 not n33444 ; n33444_not
g55200 not n46602 ; n46602_not
g55201 not n34218 ; n34218_not
g55202 not n22176 ; n22176_not
g55203 not n26343 ; n26343_not
g55204 not n26361 ; n26361_not
g55205 not n30735 ; n30735_not
g55206 not n46152 ; n46152_not
g55207 not n29322 ; n29322_not
g55208 not n22149 ; n22149_not
g55209 not n47223 ; n47223_not
g55210 not n35181 ; n35181_not
g55211 not n31554 ; n31554_not
g55212 not n23904 ; n23904_not
g55213 not n35172 ; n35172_not
g55214 not n36801 ; n36801_not
g55215 not n30915 ; n30915_not
g55216 not n35163 ; n35163_not
g55217 not n32652 ; n32652_not
g55218 not n32661 ; n32661_not
g55219 not n26505 ; n26505_not
g55220 not n38016 ; n38016_not
g55221 not n38025 ; n38025_not
g55222 not n32670 ; n32670_not
g55223 not n25092 ; n25092_not
g55224 not n34308 ; n34308_not
g55225 not n24129 ; n24129_not
g55226 not n21960 ; n21960_not
g55227 not n21951 ; n21951_not
g55228 not n38034 ; n38034_not
g55229 not n21933 ; n21933_not
g55230 not n24138 ; n24138_not
g55231 not n46035 ; n46035_not
g55232 not n24147 ; n24147_not
g55233 not n30816 ; n30816_not
g55234 not n22086 ; n22086_not
g55235 not n46701 ; n46701_not
g55236 not n35208 ; n35208_not
g55237 not n24039 ; n24039_not
g55238 not n27450 ; n27450_not
g55239 not n26424 ; n26424_not
g55240 not n27441 ; n27441_not
g55241 not n24048 ; n24048_not
g55242 not n34290 ; n34290_not
g55243 not n22059 ; n22059_not
g55244 not n46080 ; n46080_not
g55245 not n26433 ; n26433_not
g55246 not n24066 ; n24066_not
g55247 not n26442 ; n26442_not
g55248 not n24075 ; n24075_not
g55249 not n24084 ; n24084_not
g55250 not n26451 ; n26451_not
g55251 not n29241 ; n29241_not
g55252 not n22365 ; n22365_not
g55253 not n23634 ; n23634_not
g55254 not n30519 ; n30519_not
g55255 not n25236 ; n25236_not
g55256 not n33507 ; n33507_not
g55257 not n30528 ; n30528_not
g55258 not n35280 ; n35280_not
g55259 not n34146 ; n34146_not
g55260 not n22338 ; n22338_not
g55261 not n37143 ; n37143_not
g55262 not n30546 ; n30546_not
g55263 not n26226 ; n26226_not
g55264 not n29412 ; n29412_not
g55265 not n26217 ; n26217_not
g55266 not n31644 ; n31644_not
g55267 not n46206 ; n46206_not
g55268 not n25227 ; n25227_not
g55269 not n30564 ; n30564_not
g55270 not n31653 ; n31653_not
g55271 not n37008 ; n37008_not
g55272 not n25182 ; n25182_not
g55273 not n23562 ; n23562_not
g55274 not n23571 ; n23571_not
g55275 not n32436 ; n32436_not
g55276 not n28251 ; n28251_not
g55277 not n26145 ; n26145_not
g55278 not n37170 ; n37170_not
g55279 not n46233 ; n46233_not
g55280 not n23580 ; n23580_not
g55281 not n26154 ; n26154_not
g55282 not n32454 ; n32454_not
g55283 not n35307 ; n35307_not
g55284 not n22374 ; n22374_not
g55285 not n30474 ; n30474_not
g55286 not n25254 ; n25254_not
g55287 not n25245 ; n25245_not
g55288 not n30483 ; n30483_not
g55289 not n34137 ; n34137_not
g55290 not n33534 ; n33534_not
g55291 not n26190 ; n26190_not
g55292 not n33525 ; n33525_not
g55293 not n27630 ; n27630_not
g55294 not n28341 ; n28341_not
g55295 not n23742 ; n23742_not
g55296 not n22275 ; n22275_not
g55297 not n30645 ; n30645_not
g55298 not n26280 ; n26280_not
g55299 not n22266 ; n22266_not
g55300 not n33471 ; n33471_not
g55301 not n23760 ; n23760_not
g55302 not n30672 ; n30672_not
g55303 not n37080 ; n37080_not
g55304 not n31635 ; n31635_not
g55305 not n37071 ; n37071_not
g55306 not n46170 ; n46170_not
g55307 not n27540 ; n27540_not
g55308 not n46116 ; n46116_not
g55309 not n28314 ; n28314_not
g55310 not n23670 ; n23670_not
g55311 not n26244 ; n26244_not
g55312 not n25218 ; n25218_not
g55313 not n37125 ; n37125_not
g55314 not n30573 ; n30573_not
g55315 not n31671 ; n31671_not
g55316 not n37116 ; n37116_not
g55317 not n27531 ; n27531_not
g55318 not n32490 ; n32490_not
g55319 not n35271 ; n35271_not
g55320 not n37800 ; n37800_not
g55321 not n28323 ; n28323_not
g55322 not n47124 ; n47124_not
g55323 not n23706 ; n23706_not
g55324 not n23715 ; n23715_not
g55325 not n30627 ; n30627_not
g55326 not n47700 ; n47700_not
g55327 not n28332 ; n28332_not
g55328 not n37107 ; n37107_not
g55329 not n35235 ; n35235_not
g55330 not n30636 ; n30636_not
g55331 not n15507 ; n15507_not
g55332 not n20259 ; n20259_not
g55333 not n15525 ; n15525_not
g55334 not n11187 ; n11187_not
g55335 not n40941 ; n40941_not
g55336 not n45306 ; n45306_not
g55337 not n40932 ; n40932_not
g55338 not n45162 ; n45162_not
g55339 not n13752 ; n13752_not
g55340 not n41904 ; n41904_not
g55341 not n41913 ; n41913_not
g55342 not n40905 ; n40905_not
g55343 not n20196 ; n20196_not
g55344 not n20187 ; n20187_not
g55345 not n12762 ; n12762_not
g55346 not n20178 ; n20178_not
g55347 not n10971 ; n10971_not
g55348 not n39015 ; n39015_not
g55349 not n43344 ; n43344_not
g55350 not n42732 ; n42732_not
g55351 not n42525 ; n42525_not
g55352 not n44244 ; n44244_not
g55353 not n18504 ; n18504_not
g55354 not n41832 ; n41832_not
g55355 not n20376 ; n20376_not
g55356 not n42516 ; n42516_not
g55357 not n20349 ; n20349_not
g55358 not n15480 ; n15480_not
g55359 not n11448 ; n11448_not
g55360 not n18513 ; n18513_not
g55361 not n18531 ; n18531_not
g55362 not n40914 ; n40914_not
g55363 not n45315 ; n45315_not
g55364 not n20295 ; n20295_not
g55365 not n42543 ; n42543_not
g55366 not n43560 ; n43560_not
g55367 not n15039 ; n15039_not
g55368 not n39060 ; n39060_not
g55369 not n39006 ; n39006_not
g55370 not n16713 ; n16713_not
g55371 not n39123 ; n39123_not
g55372 not n14355 ; n14355_not
g55373 not n12915 ; n12915_not
g55374 not n14364 ; n14364_not
g55375 not n44550 ; n44550_not
g55376 not n10494 ; n10494_not
g55377 not n42534 ; n42534_not
g55378 not n39150 ; n39150_not
g55379 not n15327 ; n15327_not
g55380 not n16623 ; n16623_not
g55381 not n12168 ; n12168_not
g55382 not n18720 ; n18720_not
g55383 not n42048 ; n42048_not
g55384 not n14337 ; n14337_not
g55385 not n14328 ; n14328_not
g55386 not n15561 ; n15561_not
g55387 not n16812 ; n16812_not
g55388 not n12096 ; n12096_not
g55389 not n12942 ; n12942_not
g55390 not n45207 ; n45207_not
g55391 not n12933 ; n12933_not
g55392 not n43128 ; n43128_not
g55393 not n15570 ; n15570_not
g55394 not n20088 ; n20088_not
g55395 not n18612 ; n18612_not
g55396 not n41940 ; n41940_not
g55397 not n11169 ; n11169_not
g55398 not n10467 ; n10467_not
g55399 not n40815 ; n40815_not
g55400 not n14382 ; n14382_not
g55401 not n43119 ; n43119_not
g55402 not n15273 ; n15273_not
g55403 not n18324 ; n18324_not
g55404 not n11295 ; n11295_not
g55405 not n38610 ; n38610_not
g55406 not n42642 ; n42642_not
g55407 not n15291 ; n15291_not
g55408 not n20592 ; n20592_not
g55409 not n13149 ; n13149_not
g55410 not n18333 ; n18333_not
g55411 not n44037 ; n44037_not
g55412 not n18342 ; n18342_not
g55413 not n15318 ; n15318_not
g55414 not n10647 ; n10647_not
g55415 not n18351 ; n18351_not
g55416 not n20574 ; n20574_not
g55417 not n11916 ; n11916_not
g55418 not n17163 ; n17163_not
g55419 not n10908 ; n10908_not
g55420 not n20709 ; n20709_not
g55421 not n13266 ; n13266_not
g55422 not n13626 ; n13626_not
g55423 not n10359 ; n10359_not
g55424 not n41166 ; n41166_not
g55425 not n18243 ; n18243_not
g55426 not n20691 ; n20691_not
g55427 not n18261 ; n18261_not
g55428 not n11691 ; n11691_not
g55429 not n10863 ; n10863_not
g55430 not n13644 ; n13644_not
g55431 not n20673 ; n20673_not
g55432 not n17190 ; n17190_not
g55433 not n13653 ; n13653_not
g55434 not n15255 ; n15255_not
g55435 not n43515 ; n43515_not
g55436 not n10854 ; n10854_not
g55437 not n11961 ; n11961_not
g55438 not n17073 ; n17073_not
g55439 not n15408 ; n15408_not
g55440 not n14463 ; n14463_not
g55441 not n10944 ; n10944_not
g55442 not n43362 ; n43362_not
g55443 not n10926 ; n10926_not
g55444 not n20448 ; n20448_not
g55445 not n43614 ; n43614_not
g55446 not n15435 ; n15435_not
g55447 not n10449 ; n10449_not
g55448 not n42570 ; n42570_not
g55449 not n17028 ; n17028_not
g55450 not n12744 ; n12744_not
g55451 not n18414 ; n18414_not
g55452 not n10458 ; n10458_not
g55453 not n15462 ; n15462_not
g55454 not n20394 ; n20394_not
g55455 not n15471 ; n15471_not
g55456 not n41751 ; n41751_not
g55457 not n38430 ; n38430_not
g55458 not n20547 ; n20547_not
g55459 not n43524 ; n43524_not
g55460 not n41067 ; n41067_not
g55461 not n20538 ; n20538_not
g55462 not n44226 ; n44226_not
g55463 not n41058 ; n41058_not
g55464 not n15363 ; n15363_not
g55465 not n43083 ; n43083_not
g55466 not n18423 ; n18423_not
g55467 not n15372 ; n15372_not
g55468 not n38700 ; n38700_not
g55469 not n11934 ; n11934_not
g55470 not n17109 ; n17109_not
g55471 not n43371 ; n43371_not
g55472 not n11943 ; n11943_not
g55473 not n20484 ; n20484_not
g55474 not n41760 ; n41760_not
g55475 not n18441 ; n18441_not
g55476 not n40095 ; n40095_not
g55477 not n43821 ; n43821_not
g55478 not n12519 ; n12519_not
g55479 not n19701 ; n19701_not
g55480 not n42237 ; n42237_not
g55481 not n10485 ; n10485_not
g55482 not n12546 ; n12546_not
g55483 not n42228 ; n42228_not
g55484 not n19206 ; n19206_not
g55485 not n15903 ; n15903_not
g55486 not n16263 ; n16263_not
g55487 not n12708 ; n12708_not
g55488 not n16245 ; n16245_not
g55489 not n12573 ; n12573_not
g55490 not n16029 ; n16029_not
g55491 not n19224 ; n19224_not
g55492 not n16254 ; n16254_not
g55493 not n12582 ; n12582_not
g55494 not n42183 ; n42183_not
g55495 not n19413 ; n19413_not
g55496 not n43254 ; n43254_not
g55497 not n12438 ; n12438_not
g55498 not n40437 ; n40437_not
g55499 not n13932 ; n13932_not
g55500 not n15921 ; n15921_not
g55501 not n12456 ; n12456_not
g55502 not n44442 ; n44442_not
g55503 not n12474 ; n12474_not
g55504 not n13941 ; n13941_not
g55505 not n19107 ; n19107_not
g55506 not n42264 ; n42264_not
g55507 not n19116 ; n19116_not
g55508 not n12483 ; n12483_not
g55509 not n19134 ; n19134_not
g55510 not n12717 ; n12717_not
g55511 not n16317 ; n16317_not
g55512 not n42255 ; n42255_not
g55513 not n40635 ; n40635_not
g55514 not n19161 ; n19161_not
g55515 not n16281 ; n16281_not
g55516 not n43173 ; n43173_not
g55517 not n16209 ; n16209_not
g55518 not n19512 ; n19512_not
g55519 not n40167 ; n40167_not
g55520 not n42174 ; n42174_not
g55521 not n19341 ; n19341_not
g55522 not n12672 ; n12672_not
g55523 not n40194 ; n40194_not
g55524 not n16191 ; n16191_not
g55525 not n42192 ; n42192_not
g55526 not n40086 ; n40086_not
g55527 not n12654 ; n12654_not
g55528 not n19422 ; n19422_not
g55529 not n16146 ; n16146_not
g55530 not n10818 ; n10818_not
g55531 not n16164 ; n16164_not
g55532 not n40257 ; n40257_not
g55533 not n19404 ; n19404_not
g55534 not n10827 ; n10827_not
g55535 not n15147 ; n15147_not
g55536 not n16065 ; n16065_not
g55537 not n19611 ; n19611_not
g55538 not n10791 ; n10791_not
g55539 not n40347 ; n40347_not
g55540 not n19602 ; n19602_not
g55541 not n19260 ; n19260_not
g55542 not n45117 ; n45117_not
g55543 not n12591 ; n12591_not
g55544 not n16056 ; n16056_not
g55545 not n16236 ; n16236_not
g55546 not n15282 ; n15282_not
g55547 not n16227 ; n16227_not
g55548 not n19305 ; n19305_not
g55549 not n19521 ; n19521_not
g55550 not n40158 ; n40158_not
g55551 not n16173 ; n16173_not
g55552 not n39312 ; n39312_not
g55553 not n16506 ; n16506_not
g55554 not n15705 ; n15705_not
g55555 not n14256 ; n14256_not
g55556 not n42084 ; n42084_not
g55557 not n15714 ; n15714_not
g55558 not n17226 ; n17226_not
g55559 not n12834 ; n12834_not
g55560 not n42435 ; n42435_not
g55561 not n15723 ; n15723_not
g55562 not n16443 ; n16443_not
g55563 not n16470 ; n16470_not
g55564 not n40077 ; n40077_not
g55565 not n13860 ; n13860_not
g55566 not n40590 ; n40590_not
g55567 not n43632 ; n43632_not
g55568 not n12807 ; n12807_not
g55569 not n40572 ; n40572_not
g55570 not n42417 ; n42417_not
g55571 not n39213 ; n39213_not
g55572 not n12870 ; n12870_not
g55573 not n40734 ; n40734_not
g55574 not n42480 ; n42480_not
g55575 not n15651 ; n15651_not
g55576 not n12195 ; n12195_not
g55577 not n39024 ; n39024_not
g55578 not n39240 ; n39240_not
g55579 not n13833 ; n13833_not
g55580 not n16560 ; n16560_not
g55581 not n18810 ; n18810_not
g55582 not n12267 ; n12267_not
g55583 not n42075 ; n42075_not
g55584 not n18801 ; n18801_not
g55585 not n13851 ; n13851_not
g55586 not n39303 ; n39303_not
g55587 not n42462 ; n42462_not
g55588 not n14265 ; n14265_not
g55589 not n14148 ; n14148_not
g55590 not n43272 ; n43272_not
g55591 not n15831 ; n15831_not
g55592 not n40446 ; n40446_not
g55593 not n40455 ; n40455_not
g55594 not n10287 ; n10287_not
g55595 not n16353 ; n16353_not
g55596 not n43263 ; n43263_not
g55597 not n13914 ; n13914_not
g55598 not n42318 ; n42318_not
g55599 not n39420 ; n39420_not
g55600 not n12492 ; n12492_not
g55601 not n12276 ; n12276_not
g55602 not n19044 ; n19044_not
g55603 not n19053 ; n19053_not
g55604 not n42291 ; n42291_not
g55605 not n39600 ; n39600_not
g55606 not n42381 ; n42381_not
g55607 not n16416 ; n16416_not
g55608 not n38601 ; n38601_not
g55609 not n14193 ; n14193_not
g55610 not n39501 ; n39501_not
g55611 not n14175 ; n14175_not
g55612 not n14166 ; n14166_not
g55613 not n12339 ; n12339_not
g55614 not n16407 ; n16407_not
g55615 not n12348 ; n12348_not
g55616 not n44343 ; n44343_not
g55617 not n14157 ; n14157_not
g55618 not n40509 ; n40509_not
g55619 not n10629 ; n10629_not
g55620 not n15813 ; n15813_not
g55621 not n40491 ; n40491_not
g55622 not n43281 ; n43281_not
g55623 not n16371 ; n16371_not
g55624 not n16362 ; n16362_not
g55625 not n38250 ; n38250_not
g55626 not n15093 ; n15093_not
g55627 not n41481 ; n41481_not
g55628 not n43902 ; n43902_not
g55629 not n21294 ; n21294_not
g55630 not n41409 ; n41409_not
g55631 not n15075 ; n15075_not
g55632 not n14751 ; n14751_not
g55633 not n17505 ; n17505_not
g55634 not n21087 ; n21087_not
g55635 not n11664 ; n11664_not
g55636 not n14508 ; n14508_not
g55637 not n17334 ; n17334_not
g55638 not n20871 ; n20871_not
g55639 not n11529 ; n11529_not
g55640 not n17352 ; n17352_not
g55641 not n10386 ; n10386_not
g55642 not n15057 ; n15057_not
g55643 not n13581 ; n13581_not
g55644 not n18081 ; n18081_not
g55645 not n41274 ; n41274_not
g55646 not n41463 ; n41463_not
g55647 not n21348 ; n21348_not
g55648 not n18162 ; n18162_not
g55649 not n11565 ; n11565_not
g55650 not n17721 ; n17721_not
g55651 not n18144 ; n18144_not
g55652 not n11781 ; n11781_not
g55653 not n45720 ; n45720_not
g55654 not n11637 ; n11637_not
g55655 not n41508 ; n41508_not
g55656 not n14904 ; n14904_not
g55657 not n38313 ; n38313_not
g55658 not n43056 ; n43056_not
g55659 not n20835 ; n20835_not
g55660 not n41283 ; n41283_not
g55661 not n14823 ; n14823_not
g55662 not n14733 ; n14733_not
g55663 not n44370 ; n44370_not
g55664 not n17541 ; n17541_not
g55665 not n17424 ; n17424_not
g55666 not n44136 ; n44136_not
g55667 not n38403 ; n38403_not
g55668 not n41490 ; n41490_not
g55669 not n11646 ; n11646_not
g55670 not n14814 ; n14814_not
g55671 not n13356 ; n13356_not
g55672 not n14517 ; n14517_not
g55673 not n20916 ; n20916_not
g55674 not n14661 ; n14661_not
g55675 not n11709 ; n11709_not
g55676 not n38340 ; n38340_not
g55677 not n13563 ; n13563_not
g55678 not n10683 ; n10683_not
g55679 not n11466 ; n11466_not
g55680 not n18045 ; n18045_not
g55681 not n43416 ; n43416_not
g55682 not n11736 ; n11736_not
g55683 not n44154 ; n44154_not
g55684 not n18009 ; n18009_not
g55685 not n16902 ; n16902_not
g55686 not n17811 ; n17811_not
g55687 not n10692 ; n10692_not
g55688 not n13518 ; n13518_not
g55689 not n13365 ; n13365_not
g55690 not n41427 ; n41427_not
g55691 not n14760 ; n14760_not
g55692 not n11754 ; n11754_not
g55693 not n41382 ; n41382_not
g55694 not n13392 ; n13392_not
g55695 not n41454 ; n41454_not
g55696 not n17415 ; n17415_not
g55697 not n17370 ; n17370_not
g55698 not n41238 ; n41238_not
g55699 not n41337 ; n41337_not
g55700 not n41670 ; n41670_not
g55701 not n21186 ; n21186_not
g55702 not n41436 ; n41436_not
g55703 not n14625 ; n14625_not
g55704 not n14805 ; n14805_not
g55705 not n42912 ; n42912_not
g55706 not n38322 ; n38322_not
g55707 not n42921 ; n42921_not
g55708 not n40860 ; n40860_not
g55709 not n38331 ; n38331_not
g55710 not n41256 ; n41256_not
g55711 not n14562 ; n14562_not
g55712 not n41418 ; n41418_not
g55713 not n14607 ; n14607_not
g55714 not n41580 ; n41580_not
g55715 not n14526 ; n14526_not
g55716 not n41733 ; n41733_not
g55717 not n14832 ; n14832_not
g55718 not n13284 ; n13284_not
g55719 not n11808 ; n11808_not
g55720 not n41175 ; n41175_not
g55721 not n41571 ; n41571_not
g55722 not n13590 ; n13590_not
g55723 not n11583 ; n11583_not
g55724 not n41562 ; n41562_not
g55725 not n13473 ; n13473_not
g55726 not n14931 ; n14931_not
g55727 not n41193 ; n41193_not
g55728 not n20772 ; n20772_not
g55729 not n41346 ; n41346_not
g55730 not n11835 ; n11835_not
g55731 not n14742 ; n14742_not
g55732 not n21393 ; n21393_not
g55733 not n13617 ; n13617_not
g55734 not n21429 ; n21429_not
g55735 not n44055 ; n44055_not
g55736 not n14850 ; n14850_not
g55737 not n21438 ; n21438_not
g55738 not n17910 ; n17910_not
g55739 not n13545 ; n13545_not
g55740 not n17613 ; n17613_not
g55741 not n13464 ; n13464_not
g55742 not n38304 ; n38304_not
g55743 not n41328 ; n41328_not
g55744 not n44190 ; n44190_not
g55745 not n20754 ; n20754_not
g55746 not n17451 ; n17451_not
g55747 not n17262 ; n17262_not
g55748 not n13455 ; n13455_not
g55749 not n38241 ; n38241_not
g55750 not n21375 ; n21375_not
g55751 not n43452 ; n43452_not
g55752 not n18171 ; n18171_not
g55753 not n13536 ; n13536_not
g55754 not n10881 ; n10881_not
g55755 not n10548 ; n10548_not
g55756 not n20790 ; n20790_not
g55757 not n14706 ; n14706_not
g55758 not n44172 ; n44172_not
g55759 not n17316 ; n17316_not
g55760 not n10746 ; n10746_not
g55761 not n15129 ; n15129_not
g55762 not n42804 ; n42804_not
g55763 not n18135 ; n18135_not
g55764 not n45432 ; n45432_not
g55765 not n41625 ; n41625_not
g55766 not n39700 ; n39700_not
g55767 not n23662 ; n23662_not
g55768 not n23536 ; n23536_not
g55769 not n23842 ; n23842_not
g55770 not n23770 ; n23770_not
g55771 not n26623 ; n26623_not
g55772 not n30565 ; n30565_not
g55773 not n25057 ; n25057_not
g55774 not n43264 ; n43264_not
g55775 not n23833 ; n23833_not
g55776 not n40474 ; n40474_not
g55777 not n16417 ; n16417_not
g55778 not n30556 ; n30556_not
g55779 not n37063 ; n37063_not
g55780 not n32329 ; n32329_not
g55781 not n43255 ; n43255_not
g55782 not n25075 ; n25075_not
g55783 not n25084 ; n25084_not
g55784 not n19027 ; n19027_not
g55785 not n35128 ; n35128_not
g55786 not n40555 ; n40555_not
g55787 not n35047 ; n35047_not
g55788 not n16426 ; n16426_not
g55789 not n41662 ; n41662_not
g55790 not n13906 ; n13906_not
g55791 not n19009 ; n19009_not
g55792 not n26641 ; n26641_not
g55793 not n41815 ; n41815_not
g55794 not n16435 ; n16435_not
g55795 not n44461 ; n44461_not
g55796 not n41680 ; n41680_not
g55797 not n38413 ; n38413_not
g55798 not n40645 ; n40645_not
g55799 not n23653 ; n23653_not
g55800 not n30538 ; n30538_not
g55801 not n36019 ; n36019_not
g55802 not n37135 ; n37135_not
g55803 not n17470 ; n17470_not
g55804 not n40609 ; n40609_not
g55805 not n16453 ; n16453_not
g55806 not n25426 ; n25426_not
g55807 not n25372 ; n25372_not
g55808 not n31681 ; n31681_not
g55809 not n31834 ; n31834_not
g55810 not n10288 ; n10288_not
g55811 not n43282 ; n43282_not
g55812 not n37090 ; n37090_not
g55813 not n23806 ; n23806_not
g55814 not n31690 ; n31690_not
g55815 not n13528 ; n13528_not
g55816 not n16462 ; n16462_not
g55817 not n42706 ; n42706_not
g55818 not n12826 ; n12826_not
g55819 not n23707 ; n23707_not
g55820 not n16408 ; n16408_not
g55821 not n40528 ; n40528_not
g55822 not n41383 ; n41383_not
g55823 not n23716 ; n23716_not
g55824 not n13384 ; n13384_not
g55825 not n12817 ; n12817_not
g55826 not n40564 ; n40564_not
g55827 not n25048 ; n25048_not
g55828 not n13537 ; n13537_not
g55829 not n42094 ; n42094_not
g55830 not n19342 ; n19342_not
g55831 not n41347 ; n41347_not
g55832 not n30493 ; n30493_not
g55833 not n48115 ; n48115_not
g55834 not n41419 ; n41419_not
g55835 not n16363 ; n16363_not
g55836 not n36145 ; n36145_not
g55837 not n26605 ; n26605_not
g55838 not n23824 ; n23824_not
g55839 not n36172 ; n36172_not
g55840 not n30367 ; n30367_not
g55841 not n30439 ; n30439_not
g55842 not n37117 ; n37117_not
g55843 not n40618 ; n40618_not
g55844 not n23815 ; n23815_not
g55845 not n29620 ; n29620_not
g55846 not n40276 ; n40276_not
g55847 not n29530 ; n29530_not
g55848 not n25192 ; n25192_not
g55849 not n34543 ; n34543_not
g55850 not n34354 ; n34354_not
g55851 not n23392 ; n23392_not
g55852 not n19270 ; n19270_not
g55853 not n16246 ; n16246_not
g55854 not n37018 ; n37018_not
g55855 not n16228 ; n16228_not
g55856 not n44326 ; n44326_not
g55857 not n25291 ; n25291_not
g55858 not n36091 ; n36091_not
g55859 not n27019 ; n27019_not
g55860 not n42166 ; n42166_not
g55861 not n15760 ; n15760_not
g55862 not n17524 ; n17524_not
g55863 not n23446 ; n23446_not
g55864 not n34615 ; n34615_not
g55865 not n25327 ; n25327_not
g55866 not n19216 ; n19216_not
g55867 not n23428 ; n23428_not
g55868 not n17236 ; n17236_not
g55869 not n17551 ; n17551_not
g55870 not n16723 ; n16723_not
g55871 not n31825 ; n31825_not
g55872 not n19234 ; n19234_not
g55873 not n40357 ; n40357_not
g55874 not n16255 ; n16255_not
g55875 not n13483 ; n13483_not
g55876 not n34570 ; n34570_not
g55877 not n41626 ; n41626_not
g55878 not n34561 ; n34561_not
g55879 not n30088 ; n30088_not
g55880 not n17704 ; n17704_not
g55881 not n25237 ; n25237_not
g55882 not n34525 ; n34525_not
g55883 not n44551 ; n44551_not
g55884 not n25246 ; n25246_not
g55885 not n19351 ; n19351_not
g55886 not n40285 ; n40285_not
g55887 not n27073 ; n27073_not
g55888 not n16174 ; n16174_not
g55889 not n37261 ; n37261_not
g55890 not n27046 ; n27046_not
g55891 not n10576 ; n10576_not
g55892 not n41608 ; n41608_not
g55893 not n30637 ; n30637_not
g55894 not n17623 ; n17623_not
g55895 not n43183 ; n43183_not
g55896 not n17128 ; n17128_not
g55897 not n13465 ; n13465_not
g55898 not n19315 ; n19315_not
g55899 not n30079 ; n30079_not
g55900 not n23365 ; n23365_not
g55901 not n42139 ; n42139_not
g55902 not n25264 ; n25264_not
g55903 not n19324 ; n19324_not
g55904 not n25273 ; n25273_not
g55905 not n41581 ; n41581_not
g55906 not n13429 ; n13429_not
g55907 not n23356 ; n23356_not
g55908 not n12673 ; n12673_not
g55909 not n17254 ; n17254_not
g55910 not n15823 ; n15823_not
g55911 not n32392 ; n32392_not
g55912 not n29521 ; n29521_not
g55913 not n17641 ; n17641_not
g55914 not n47251 ; n47251_not
g55915 not n43714 ; n43714_not
g55916 not n26803 ; n26803_not
g55917 not n40429 ; n40429_not
g55918 not n13933 ; n13933_not
g55919 not n32266 ; n32266_not
g55920 not n40393 ; n40393_not
g55921 not n30574 ; n30574_not
g55922 not n34822 ; n34822_not
g55923 not n17803 ; n17803_not
g55924 not n12727 ; n12727_not
g55925 not n32347 ; n32347_not
g55926 not n36046 ; n36046_not
g55927 not n43246 ; n43246_not
g55928 not n23554 ; n23554_not
g55929 not n10279 ; n10279_not
g55930 not n30097 ; n30097_not
g55931 not n13924 ; n13924_not
g55932 not n23617 ; n23617_not
g55933 not n16345 ; n16345_not
g55934 not n23626 ; n23626_not
g55935 not n36037 ; n36037_not
g55936 not n19054 ; n19054_not
g55937 not n16930 ; n16930_not
g55938 not n40780 ; n40780_not
g55939 not n19063 ; n19063_not
g55940 not n34840 ; n34840_not
g55941 not n43426 ; n43426_not
g55942 not n40438 ; n40438_not
g55943 not n47242 ; n47242_not
g55944 not n16327 ; n16327_not
g55945 not n34831 ; n34831_not
g55946 not n37162 ; n37162_not
g55947 not n12736 ; n12736_not
g55948 not n25129 ; n25129_not
g55949 not n37207 ; n37207_not
g55950 not n32365 ; n32365_not
g55951 not n40384 ; n40384_not
g55952 not n26911 ; n26911_not
g55953 not n17506 ; n17506_not
g55954 not n32293 ; n32293_not
g55955 not n32374 ; n32374_not
g55956 not n23455 ; n23455_not
g55957 not n31654 ; n31654_not
g55958 not n47323 ; n47323_not
g55959 not n34642 ; n34642_not
g55960 not n41644 ; n41644_not
g55961 not n43723 ; n43723_not
g55962 not n37225 ; n37225_not
g55963 not n19117 ; n19117_not
g55964 not n42148 ; n42148_not
g55965 not n46522 ; n46522_not
g55966 not n34804 ; n34804_not
g55967 not n19126 ; n19126_not
g55968 not n23527 ; n23527_not
g55969 not n23518 ; n23518_not
g55970 not n32356 ; n32356_not
g55971 not n34732 ; n34732_not
g55972 not n23509 ; n23509_not
g55973 not n43228 ; n43228_not
g55974 not n30583 ; n30583_not
g55975 not n34723 ; n34723_not
g55976 not n19162 ; n19162_not
g55977 not n30592 ; n30592_not
g55978 not n21637 ; n21637_not
g55979 not n17065 ; n17065_not
g55980 not n18127 ; n18127_not
g55981 not n24805 ; n24805_not
g55982 not n31753 ; n31753_not
g55983 not n35803 ; n35803_not
g55984 not n35821 ; n35821_not
g55985 not n31942 ; n31942_not
g55986 not n18109 ; n18109_not
g55987 not n24814 ; n24814_not
g55988 not n17038 ; n17038_not
g55989 not n10945 ; n10945_not
g55990 not n42733 ; n42733_not
g55991 not n35344 ; n35344_not
g55992 not n48502 ; n48502_not
g55993 not n24373 ; n24373_not
g55994 not n10954 ; n10954_not
g55995 not n25633 ; n25633_not
g55996 not n36451 ; n36451_not
g55997 not n48250 ; n48250_not
g55998 not n36406 ; n36406_not
g55999 not n25714 ; n25714_not
g56000 not n31933 ; n31933_not
g56001 not n35353 ; n35353_not
g56002 not n35119 ; n35119_not
g56003 not n24427 ; n24427_not
g56004 not n18406 ; n18406_not
g56005 not n25921 ; n25921_not
g56006 not n24418 ; n24418_not
g56007 not n36361 ; n36361_not
g56008 not n35731 ; n35731_not
g56009 not n47206 ; n47206_not
g56010 not n18451 ; n18451_not
g56011 not n30286 ; n30286_not
g56012 not n24724 ; n24724_not
g56013 not n29800 ; n29800_not
g56014 not n31915 ; n31915_not
g56015 not n18073 ; n18073_not
g56016 not n40159 ; n40159_not
g56017 not n35317 ; n35317_not
g56018 not n44353 ; n44353_not
g56019 not n13573 ; n13573_not
g56020 not n18541 ; n18541_not
g56021 not n35902 ; n35902_not
g56022 not n41707 ; n41707_not
g56023 not n26119 ; n26119_not
g56024 not n47080 ; n47080_not
g56025 not n10891 ; n10891_not
g56026 not n12970 ; n12970_not
g56027 not n32158 ; n32158_not
g56028 not n26092 ; n26092_not
g56029 not n25363 ; n25363_not
g56030 not n10855 ; n10855_not
g56031 not n24274 ; n24274_not
g56032 not n31744 ; n31744_not
g56033 not n13726 ; n13726_not
g56034 not n43543 ; n43543_not
g56035 not n10459 ; n10459_not
g56036 not n41806 ; n41806_not
g56037 not n10963 ; n10963_not
g56038 not n48160 ; n48160_not
g56039 not n35335 ; n35335_not
g56040 not n31735 ; n31735_not
g56041 not n24841 ; n24841_not
g56042 not n41824 ; n41824_not
g56043 not n36334 ; n36334_not
g56044 not n24850 ; n24850_not
g56045 not n24238 ; n24238_not
g56046 not n36622 ; n36622_not
g56047 not n47071 ; n47071_not
g56048 not n18514 ; n18514_not
g56049 not n24319 ; n24319_not
g56050 not n41185 ; n41185_not
g56051 not n48430 ; n48430_not
g56052 not n25804 ; n25804_not
g56053 not n18271 ; n18271_not
g56054 not n36532 ; n36532_not
g56055 not n36541 ; n36541_not
g56056 not n24580 ; n24580_not
g56057 not n35515 ; n35515_not
g56058 not n10927 ; n10927_not
g56059 not n41149 ; n41149_not
g56060 not n24571 ; n24571_not
g56061 not n13195 ; n13195_not
g56062 not n32086 ; n32086_not
g56063 not n13177 ; n13177_not
g56064 not n24562 ; n24562_not
g56065 not n36460 ; n36460_not
g56066 not n25822 ; n25822_not
g56067 not n13267 ; n13267_not
g56068 not n18217 ; n18217_not
g56069 not n18208 ; n18208_not
g56070 not n35614 ; n35614_not
g56071 not n25831 ; n25831_not
g56072 not n13258 ; n13258_not
g56073 not n13618 ; n13618_not
g56074 not n25651 ; n25651_not
g56075 not n24616 ; n24616_not
g56076 not n24490 ; n24490_not
g56077 not n13249 ; n13249_not
g56078 not n18253 ; n18253_not
g56079 not n25813 ; n25813_not
g56080 not n44506 ; n44506_not
g56081 not n13609 ; n13609_not
g56082 not n24517 ; n24517_not
g56083 not n18352 ; n18352_not
g56084 not n41725 ; n41725_not
g56085 not n18361 ; n18361_not
g56086 not n25723 ; n25723_not
g56087 not n10936 ; n10936_not
g56088 not n36604 ; n36604_not
g56089 not n24751 ; n24751_not
g56090 not n40096 ; n40096_not
g56091 not n36415 ; n36415_not
g56092 not n13096 ; n13096_not
g56093 not n41077 ; n41077_not
g56094 not n24472 ; n24472_not
g56095 not n30187 ; n30187_not
g56096 not n41770 ; n41770_not
g56097 not n41068 ; n41068_not
g56098 not n18415 ; n18415_not
g56099 not n17182 ; n17182_not
g56100 not n24391 ; n24391_not
g56101 not n13285 ; n13285_not
g56102 not n13672 ; n13672_not
g56103 not n18118 ; n18118_not
g56104 not n30169 ; n30169_not
g56105 not n13681 ; n13681_not
g56106 not n48232 ; n48232_not
g56107 not n25930 ; n25930_not
g56108 not n35452 ; n35452_not
g56109 not n13690 ; n13690_not
g56110 not n13582 ; n13582_not
g56111 not n25750 ; n25750_not
g56112 not n35713 ; n35713_not
g56113 not n18343 ; n18343_not
g56114 not n24526 ; n24526_not
g56115 not n35443 ; n35443_not
g56116 not n24733 ; n24733_not
g56117 not n43480 ; n43480_not
g56118 not n30196 ; n30196_not
g56119 not n17164 ; n17164_not
g56120 not n16624 ; n16624_not
g56121 not n36208 ; n36208_not
g56122 not n40744 ; n40744_not
g56123 not n43606 ; n43606_not
g56124 not n43309 ; n43309_not
g56125 not n12880 ; n12880_not
g56126 not n26434 ; n26434_not
g56127 not n42049 ; n42049_not
g56128 not n40735 ; n40735_not
g56129 not n17425 ; n17425_not
g56130 not n12871 ; n12871_not
g56131 not n43615 ; n43615_not
g56132 not n31708 ; n31708_not
g56133 not n42058 ; n42058_not
g56134 not n41329 ; n41329_not
g56135 not n26452 ; n26452_not
g56136 not n35191 ; n35191_not
g56137 not n26308 ; n26308_not
g56138 not n16714 ; n16714_not
g56139 not n36190 ; n36190_not
g56140 not n35245 ; n35245_not
g56141 not n26326 ; n26326_not
g56142 not n41275 ; n41275_not
g56143 not n48124 ; n48124_not
g56144 not n31852 ; n31852_not
g56145 not n35227 ; n35227_not
g56146 not n43417 ; n43417_not
g56147 not n13780 ; n13780_not
g56148 not n24076 ; n24076_not
g56149 not n40762 ; n40762_not
g56150 not n35218 ; n35218_not
g56151 not n16642 ; n16642_not
g56152 not n40753 ; n40753_not
g56153 not n43318 ; n43318_not
g56154 not n48241 ; n48241_not
g56155 not n40690 ; n40690_not
g56156 not n12853 ; n12853_not
g56157 not n44650 ; n44650_not
g56158 not n16561 ; n16561_not
g56159 not n23905 ; n23905_not
g56160 not n36181 ; n36181_not
g56161 not n40681 ; n40681_not
g56162 not n25480 ; n25480_not
g56163 not n26515 ; n26515_not
g56164 not n12745 ; n12745_not
g56165 not n25471 ; n25471_not
g56166 not n10837 ; n10837_not
g56167 not n40654 ; n40654_not
g56168 not n26542 ; n26542_not
g56169 not n25462 ; n25462_not
g56170 not n31843 ; n31843_not
g56171 not n40726 ; n40726_not
g56172 not n10819 ; n10819_not
g56173 not n12844 ; n12844_not
g56174 not n12862 ; n12862_not
g56175 not n35173 ; n35173_not
g56176 not n24931 ; n24931_not
g56177 not n43624 ; n43624_not
g56178 not n16570 ; n16570_not
g56179 not n23950 ; n23950_not
g56180 not n17137 ; n17137_not
g56181 not n30466 ; n30466_not
g56182 not n40717 ; n40717_not
g56183 not n40708 ; n40708_not
g56184 not n35155 ; n35155_not
g56185 not n35146 ; n35146_not
g56186 not n36730 ; n36730_not
g56187 not n36262 ; n36262_not
g56188 not n48403 ; n48403_not
g56189 not n41914 ; n41914_not
g56190 not n24913 ; n24913_not
g56191 not n35290 ; n35290_not
g56192 not n10972 ; n10972_not
g56193 not n31816 ; n31816_not
g56194 not n36523 ; n36523_not
g56195 not n24193 ; n24193_not
g56196 not n12907 ; n12907_not
g56197 not n32185 ; n32185_not
g56198 not n25552 ; n25552_not
g56199 not n35281 ; n35281_not
g56200 not n41923 ; n41923_not
g56201 not n26209 ; n26209_not
g56202 not n25543 ; n25543_not
g56203 not n36811 ; n36811_not
g56204 not n13339 ; n13339_not
g56205 not n40672 ; n40672_not
g56206 not n26146 ; n26146_not
g56207 not n13348 ; n13348_not
g56208 not n32167 ; n32167_not
g56209 not n40933 ; n40933_not
g56210 not n38701 ; n38701_not
g56211 not n40870 ; n40870_not
g56212 not n26164 ; n26164_not
g56213 not n40087 ; n40087_not
g56214 not n32176 ; n32176_not
g56215 not n43453 ; n43453_not
g56216 not n13357 ; n13357_not
g56217 not n40915 ; n40915_not
g56218 not n41905 ; n41905_not
g56219 not n17380 ; n17380_not
g56220 not n41239 ; n41239_not
g56221 not n30358 ; n30358_not
g56222 not n24940 ; n24940_not
g56223 not n40834 ; n40834_not
g56224 not n41248 ; n41248_not
g56225 not n38431 ; n38431_not
g56226 not n48142 ; n48142_not
g56227 not n31870 ; n31870_not
g56228 not n48133 ; n48133_not
g56229 not n26272 ; n26272_not
g56230 not n35263 ; n35263_not
g56231 not n40807 ; n40807_not
g56232 not n30394 ; n30394_not
g56233 not n36820 ; n36820_not
g56234 not n26281 ; n26281_not
g56235 not n41257 ; n41257_not
g56236 not n35254 ; n35254_not
g56237 not n13771 ; n13771_not
g56238 not n40771 ; n40771_not
g56239 not n46711 ; n46711_not
g56240 not n13762 ; n13762_not
g56241 not n16831 ; n16831_not
g56242 not n24922 ; n24922_not
g56243 not n25534 ; n25534_not
g56244 not n26128 ; n26128_not
g56245 not n24166 ; n24166_not
g56246 not n36253 ; n36253_not
g56247 not n41932 ; n41932_not
g56248 not n40852 ; n40852_not
g56249 not n36244 ; n36244_not
g56250 not n17407 ; n17407_not
g56251 not n24157 ; n24157_not
g56252 not n40843 ; n40843_not
g56253 not n18019 ; n18019_not
g56254 not n16804 ; n16804_not
g56255 not n24139 ; n24139_not
g56256 not n44614 ; n44614_not
g56257 not n35272 ; n35272_not
g56258 not n28063 ; n28063_not
g56259 not n20386 ; n20386_not
g56260 not n33634 ; n33634_not
g56261 not n22294 ; n22294_not
g56262 not n11188 ; n11188_not
g56263 not n47611 ; n47611_not
g56264 not n22285 ; n22285_not
g56265 not n42571 ; n42571_not
g56266 not n43516 ; n43516_not
g56267 not n28018 ; n28018_not
g56268 not n15445 ; n15445_not
g56269 not n22276 ; n22276_not
g56270 not n11980 ; n11980_not
g56271 not n11971 ; n11971_not
g56272 not n20458 ; n20458_not
g56273 not n15148 ; n15148_not
g56274 not n46180 ; n46180_not
g56275 not n22249 ; n22249_not
g56276 not n15409 ; n15409_not
g56277 not n45280 ; n45280_not
g56278 not n45154 ; n45154_not
g56279 not n14437 ; n14437_not
g56280 not n33733 ; n33733_not
g56281 not n15535 ; n15535_not
g56282 not n33724 ; n33724_not
g56283 not n11197 ; n11197_not
g56284 not n12079 ; n12079_not
g56285 not n29233 ; n29233_not
g56286 not n22384 ; n22384_not
g56287 not n15508 ; n15508_not
g56288 not n20296 ; n20296_not
g56289 not n33661 ; n33661_not
g56290 not n22348 ; n22348_not
g56291 not n15490 ; n15490_not
g56292 not n32545 ; n32545_not
g56293 not n46207 ; n46207_not
g56294 not n20377 ; n20377_not
g56295 not n20467 ; n20467_not
g56296 not n33562 ; n33562_not
g56297 not n15256 ; n15256_not
g56298 not n46144 ; n46144_not
g56299 not n33535 ; n33535_not
g56300 not n15292 ; n15292_not
g56301 not n38620 ; n38620_not
g56302 not n15283 ; n15283_not
g56303 not n42643 ; n42643_not
g56304 not n22096 ; n22096_not
g56305 not n20629 ; n20629_not
g56306 not n20638 ; n20638_not
g56307 not n15247 ; n15247_not
g56308 not n14914 ; n14914_not
g56309 not n22078 ; n22078_not
g56310 not n20665 ; n20665_not
g56311 not n38602 ; n38602_not
g56312 not n28324 ; n28324_not
g56313 not n15238 ; n15238_not
g56314 not n10648 ; n10648_not
g56315 not n28153 ; n28153_not
g56316 not n33616 ; n33616_not
g56317 not n15382 ; n15382_not
g56318 not n28171 ; n28171_not
g56319 not n11935 ; n11935_not
g56320 not n31438 ; n31438_not
g56321 not n11269 ; n11269_not
g56322 not n15364 ; n15364_not
g56323 not n22195 ; n22195_not
g56324 not n42616 ; n42616_not
g56325 not n32716 ; n32716_not
g56326 not n22186 ; n22186_not
g56327 not n42625 ; n42625_not
g56328 not n28207 ; n28207_not
g56329 not n22168 ; n22168_not
g56330 not n33571 ; n33571_not
g56331 not n11917 ; n11917_not
g56332 not n22159 ; n22159_not
g56333 not n30943 ; n30943_not
g56334 not n32590 ; n32590_not
g56335 not n43138 ; n43138_not
g56336 not n10486 ; n10486_not
g56337 not n12187 ; n12187_not
g56338 not n22591 ; n22591_not
g56339 not n15319 ; n15319_not
g56340 not n47440 ; n47440_not
g56341 not n42454 ; n42454_not
g56342 not n22582 ; n22582_not
g56343 not n15328 ; n15328_not
g56344 not n22573 ; n22573_not
g56345 not n39160 ; n39160_not
g56346 not n30961 ; n30961_not
g56347 not n29314 ; n29314_not
g56348 not n42508 ; n42508_not
g56349 not n15526 ; n15526_not
g56350 not n29305 ; n29305_not
g56351 not n22546 ; n22546_not
g56352 not n22555 ; n22555_not
g56353 not n39133 ; n39133_not
g56354 not n22672 ; n22672_not
g56355 not n34084 ; n34084_not
g56356 not n36028 ; n36028_not
g56357 not n29341 ; n29341_not
g56358 not n22663 ; n22663_not
g56359 not n27703 ; n27703_not
g56360 not n30925 ; n30925_not
g56361 not n30934 ; n30934_not
g56362 not n34075 ; n34075_not
g56363 not n42472 ; n42472_not
g56364 not n15661 ; n15661_not
g56365 not n22645 ; n22645_not
g56366 not n44254 ; n44254_not
g56367 not n30862 ; n30862_not
g56368 not n22636 ; n22636_not
g56369 not n19900 ; n19900_not
g56370 not n15643 ; n15643_not
g56371 not n39232 ; n39232_not
g56372 not n16840 ; n16840_not
g56373 not n22618 ; n22618_not
g56374 not n22483 ; n22483_not
g56375 not n20098 ; n20098_not
g56376 not n33814 ; n33814_not
g56377 not n42526 ; n42526_not
g56378 not n45217 ; n45217_not
g56379 not n27721 ; n27721_not
g56380 not n39034 ; n39034_not
g56381 not n22465 ; n22465_not
g56382 not n33805 ; n33805_not
g56383 not n46252 ; n46252_not
g56384 not n22429 ; n22429_not
g56385 not n39016 ; n39016_not
g56386 not n15553 ; n15553_not
g56387 not n42535 ; n42535_not
g56388 not n14419 ; n14419_not
g56389 not n20188 ; n20188_not
g56390 not n15544 ; n15544_not
g56391 not n33742 ; n33742_not
g56392 not n45271 ; n45271_not
g56393 not n33715 ; n33715_not
g56394 not n39124 ; n39124_not
g56395 not n22519 ; n22519_not
g56396 not n32608 ; n32608_not
g56397 not n39115 ; n39115_not
g56398 not n33940 ; n33940_not
g56399 not n14374 ; n14374_not
g56400 not n33922 ; n33922_not
g56401 not n33913 ; n33913_not
g56402 not n47521 ; n47521_not
g56403 not n31456 ; n31456_not
g56404 not n27712 ; n27712_not
g56405 not n32626 ; n32626_not
g56406 not n33841 ; n33841_not
g56407 not n33823 ; n33823_not
g56408 not n43129 ; n43129_not
g56409 not n22492 ; n22492_not
g56410 not n33832 ; n33832_not
g56411 not n47530 ; n47530_not
g56412 not n31465 ; n31465_not
g56413 not n14608 ; n14608_not
g56414 not n21088 ; n21088_not
g56415 not n38170 ; n38170_not
g56416 not n11593 ; n11593_not
g56417 not n21628 ; n21628_not
g56418 not n14617 ; n14617_not
g56419 not n21673 ; n21673_not
g56420 not n42904 ; n42904_not
g56421 not n44137 ; n44137_not
g56422 not n11539 ; n11539_not
g56423 not n21646 ; n21646_not
g56424 not n14815 ; n14815_not
g56425 not n21169 ; n21169_not
g56426 not n33058 ; n33058_not
g56427 not n21196 ; n21196_not
g56428 not n33139 ; n33139_not
g56429 not n11476 ; n11476_not
g56430 not n28801 ; n28801_not
g56431 not n48016 ; n48016_not
g56432 not n21592 ; n21592_not
g56433 not n21754 ; n21754_not
g56434 not n33265 ; n33265_not
g56435 not n11656 ; n11656_not
g56436 not n33256 ; n33256_not
g56437 not n33247 ; n33247_not
g56438 not n14905 ; n14905_not
g56439 not n21745 ; n21745_not
g56440 not n21736 ; n21736_not
g56441 not n11638 ; n11638_not
g56442 not n21727 ; n21727_not
g56443 not n45910 ; n45910_not
g56444 not n42760 ; n42760_not
g56445 not n10387 ; n10387_not
g56446 not n31276 ; n31276_not
g56447 not n31267 ; n31267_not
g56448 not n38305 ; n38305_not
g56449 not n42841 ; n42841_not
g56450 not n48007 ; n48007_not
g56451 not n14851 ; n14851_not
g56452 not n11386 ; n11386_not
g56453 not n32833 ; n32833_not
g56454 not n21367 ; n21367_not
g56455 not n33049 ; n33049_not
g56456 not n14716 ; n14716_not
g56457 not n21376 ; n21376_not
g56458 not n31366 ; n31366_not
g56459 not n32806 ; n32806_not
g56460 not n14671 ; n14671_not
g56461 not n21493 ; n21493_not
g56462 not n31375 ; n31375_not
g56463 not n14662 ; n14662_not
g56464 not n32950 ; n32950_not
g56465 not n44191 ; n44191_not
g56466 not n21475 ; n21475_not
g56467 not n32941 ; n32941_not
g56468 not n32932 ; n32932_not
g56469 not n43048 ; n43048_not
g56470 not n44416 ; n44416_not
g56471 not n31393 ; n31393_not
g56472 not n32923 ; n32923_not
g56473 not n21448 ; n21448_not
g56474 not n47026 ; n47026_not
g56475 not n38215 ; n38215_not
g56476 not n21583 ; n21583_not
g56477 not n31348 ; n31348_not
g56478 not n21574 ; n21574_not
g56479 not n21268 ; n21268_not
g56480 not n32842 ; n32842_not
g56481 not n14743 ; n14743_not
g56482 not n21277 ; n21277_not
g56483 not n11467 ; n11467_not
g56484 not n33085 ; n33085_not
g56485 not n21556 ; n21556_not
g56486 not n33076 ; n33076_not
g56487 not n21547 ; n21547_not
g56488 not n31357 ; n31357_not
g56489 not n45703 ; n45703_not
g56490 not n14653 ; n14653_not
g56491 not n21538 ; n21538_not
g56492 not n45712 ; n45712_not
g56493 not n45820 ; n45820_not
g56494 not n21529 ; n21529_not
g56495 not n21349 ; n21349_not
g56496 not n15175 ; n15175_not
g56497 not n15166 ; n15166_not
g56498 not n33427 ; n33427_not
g56499 not n28405 ; n28405_not
g56500 not n42409 ; n42409_not
g56501 not n38035 ; n38035_not
g56502 not n21952 ; n21952_not
g56503 not n40951 ; n40951_not
g56504 not n20782 ; n20782_not
g56505 not n28216 ; n28216_not
g56506 not n38053 ; n38053_not
g56507 not n29116 ; n29116_not
g56508 not n10639 ; n10639_not
g56509 not n42661 ; n42661_not
g56510 not n28432 ; n28432_not
g56511 not n21934 ; n21934_not
g56512 not n33409 ; n33409_not
g56513 not n46036 ; n46036_not
g56514 not n20809 ; n20809_not
g56515 not n11863 ; n11863_not
g56516 not n44056 ; n44056_not
g56517 not n11854 ; n11854_not
g56518 not n11764 ; n11764_not
g56519 not n28342 ; n28342_not
g56520 not n33490 ; n33490_not
g56521 not n31177 ; n31177_not
g56522 not n38530 ; n38530_not
g56523 not n14509 ; n14509_not
g56524 not n33472 ; n33472_not
g56525 not n15184 ; n15184_not
g56526 not n46054 ; n46054_not
g56527 not n42652 ; n42652_not
g56528 not n38512 ; n38512_not
g56529 not n38503 ; n38503_not
g56530 not n11827 ; n11827_not
g56531 not n29125 ; n29125_not
g56532 not n20746 ; n20746_not
g56533 not n14518 ; n14518_not
g56534 not n11818 ; n11818_not
g56535 not n33436 ; n33436_not
g56536 not n10675 ; n10675_not
g56537 not n42715 ; n42715_not
g56538 not n42742 ; n42742_not
g56539 not n42751 ; n42751_not
g56540 not n20944 ; n20944_not
g56541 not n38107 ; n38107_not
g56542 not n20953 ; n20953_not
g56543 not n11719 ; n11719_not
g56544 not n20908 ; n20908_not
g56545 not n20971 ; n20971_not
g56546 not n38116 ; n38116_not
g56547 not n33292 ; n33292_not
g56548 not n43075 ; n43075_not
g56549 not n32815 ; n32815_not
g56550 not n20980 ; n20980_not
g56551 not n21781 ; n21781_not
g56552 not n11665 ; n11665_not
g56553 not n29062 ; n29062_not
g56554 not n31258 ; n31258_not
g56555 not n38134 ; n38134_not
g56556 not n20818 ; n20818_not
g56557 not n10666 ; n10666_not
g56558 not n20827 ; n20827_not
g56559 not n21916 ; n21916_not
g56560 not n38404 ; n38404_not
g56561 not n21907 ; n21907_not
g56562 not n15094 ; n15094_not
g56563 not n20845 ; n20845_not
g56564 not n33382 ; n33382_not
g56565 not n21880 ; n21880_not
g56566 not n20872 ; n20872_not
g56567 not n15067 ; n15067_not
g56568 not n28513 ; n28513_not
g56569 not n20881 ; n20881_not
g56570 not n21862 ; n21862_not
g56571 not n28531 ; n28531_not
g56572 not n32761 ; n32761_not
g56573 not n38350 ; n38350_not
g56574 not n31339 ; n31339_not
g56575 not n44218 ; n44218_not
g56576 not n33337 ; n33337_not
g56577 not n21844 ; n21844_not
g56578 not n10765 ; n10765_not
g56579 not n15805 ; n15805_not
g56580 not n37414 ; n37414_not
g56581 not n42292 ; n42292_not
g56582 not n15904 ; n15904_not
g56583 not n22951 ; n22951_not
g56584 not n15049 ; n15049_not
g56585 not n31609 ; n31609_not
g56586 not n34318 ; n34318_not
g56587 not n43840 ; n43840_not
g56588 not n15913 ; n15913_not
g56589 not n22960 ; n22960_not
g56590 not n30781 ; n30781_not
g56591 not n12448 ; n12448_not
g56592 not n30772 ; n30772_not
g56593 not n37360 ; n37360_not
g56594 not n32464 ; n32464_not
g56595 not n34345 ; n34345_not
g56596 not n27352 ; n27352_not
g56597 not n12484 ; n12484_not
g56598 not n29440 ; n29440_not
g56599 not n15931 ; n15931_not
g56600 not n37333 ; n37333_not
g56601 not n30745 ; n30745_not
g56602 not n46423 ; n46423_not
g56603 not n30754 ; n30754_not
g56604 not n27325 ; n27325_not
g56605 not n42274 ; n42274_not
g56606 not n37531 ; n37531_not
g56607 not n27550 ; n27550_not
g56608 not n46360 ; n46360_not
g56609 not n22753 ; n22753_not
g56610 not n30871 ; n30871_not
g56611 not n27532 ; n27532_not
g56612 not n42373 ; n42373_not
g56613 not n34228 ; n34228_not
g56614 not n42364 ; n42364_not
g56615 not n34237 ; n34237_not
g56616 not n34246 ; n34246_not
g56617 not n22825 ; n22825_not
g56618 not n27505 ; n27505_not
g56619 not n10756 ; n10756_not
g56620 not n34291 ; n34291_not
g56621 not n42337 ; n42337_not
g56622 not n39520 ; n39520_not
g56623 not n27442 ; n27442_not
g56624 not n29413 ; n29413_not
g56625 not n19801 ; n19801_not
g56626 not n37432 ; n37432_not
g56627 not n27451 ; n27451_not
g56628 not n34273 ; n34273_not
g56629 not n34264 ; n34264_not
g56630 not n32482 ; n32482_not
g56631 not n14149 ; n14149_not
g56632 not n34255 ; n34255_not
g56633 not n22843 ; n22843_not
g56634 not n44290 ; n44290_not
g56635 not n36631 ; n36631_not
g56636 not n16075 ; n16075_not
g56637 not n34471 ; n34471_not
g56638 not n23167 ; n23167_not
g56639 not n27082 ; n27082_not
g56640 not n19531 ; n19531_not
g56641 not n42175 ; n42175_not
g56642 not n12592 ; n12592_not
g56643 not n30664 ; n30664_not
g56644 not n27163 ; n27163_not
g56645 not n32419 ; n32419_not
g56646 not n16084 ; n16084_not
g56647 not n34480 ; n34480_not
g56648 not n39412 ; n39412_not
g56649 not n19522 ; n19522_not
g56650 not n27154 ; n27154_not
g56651 not n19513 ; n19513_not
g56652 not n43741 ; n43741_not
g56653 not n17605 ; n17605_not
g56654 not n44407 ; n44407_not
g56655 not n40186 ; n40186_not
g56656 not n44722 ; n44722_not
g56657 not n12619 ; n12619_not
g56658 not n12637 ; n12637_not
g56659 not n16138 ; n16138_not
g56660 not n27118 ; n27118_not
g56661 not n19414 ; n19414_not
g56662 not n34327 ; n34327_not
g56663 not n23284 ; n23284_not
g56664 not n37270 ; n37270_not
g56665 not n46441 ; n46441_not
g56666 not n42265 ; n42265_not
g56667 not n10774 ; n10774_not
g56668 not n34381 ; n34381_not
g56669 not n43831 ; n43831_not
g56670 not n30736 ; n30736_not
g56671 not n34390 ; n34390_not
g56672 not n14086 ; n14086_not
g56673 not n37315 ; n37315_not
g56674 not n19720 ; n19720_not
g56675 not n27280 ; n27280_not
g56676 not n30727 ; n30727_not
g56677 not n27262 ; n27262_not
g56678 not n42247 ; n42247_not
g56679 not n14077 ; n14077_not
g56680 not n19621 ; n19621_not
g56681 not n19630 ; n19630_not
g56682 not n16057 ; n16057_not
g56683 not n27226 ; n27226_not
g56684 not n43813 ; n43813_not
g56685 not n12565 ; n12565_not
g56686 not n12556 ; n12556_not
g56687 not n27235 ; n27235_not
g56688 not n30709 ; n30709_not
g56689 not n32446 ; n32446_not
g56690 not n12538 ; n12538_not
g56691 not n30718 ; n30718_not
g56692 not n30880 ; n30880_not
g56693 not n31528 ; n31528_not
g56694 not n37540 ; n37540_not
g56695 not n47413 ; n47413_not
g56696 not n30916 ; n30916_not
g56697 not n31537 ; n31537_not
g56698 not n22717 ; n22717_not
g56699 not n32554 ; n32554_not
g56700 not n27631 ; n27631_not
g56701 not n15724 ; n15724_not
g56702 not n34165 ; n34165_not
g56703 not n39421 ; n39421_not
g56704 not n39340 ; n39340_not
g56705 not n22726 ; n22726_not
g56706 not n12286 ; n12286_not
g56707 not n30835 ; n30835_not
g56708 not n14239 ; n14239_not
g56709 not n32509 ; n32509_not
g56710 not n42436 ; n42436_not
g56711 not n34183 ; n34183_not
g56712 not n22744 ; n22744_not
g56713 not n44425 ; n44425_not
g56714 not n22681 ; n22681_not
g56715 not n42445 ; n42445_not
g56716 not n15715 ; n15715_not
g56717 not n14951 ; n14951_not
g56718 not n35912 ; n35912_not
g56719 not n25571 ; n25571_not
g56720 not n42248 ; n42248_not
g56721 not n13565 ; n13565_not
g56722 not n16490 ; n16490_not
g56723 not n29072 ; n29072_not
g56724 not n16265 ; n16265_not
g56725 not n35138 ; n35138_not
g56726 not n17381 ; n17381_not
g56727 not n25544 ; n25544_not
g56728 not n32807 ; n32807_not
g56729 not n26444 ; n26444_not
g56730 not n26921 ; n26921_not
g56731 not n17075 ; n17075_not
g56732 not n17336 ; n17336_not
g56733 not n28550 ; n28550_not
g56734 not n17048 ; n17048_not
g56735 not n47153 ; n47153_not
g56736 not n25562 ; n25562_not
g56737 not n14960 ; n14960_not
g56738 not n34706 ; n34706_not
g56739 not n42725 ; n42725_not
g56740 not n10982 ; n10982_not
g56741 not n34634 ; n34634_not
g56742 not n29540 ; n29540_not
g56743 not n27560 ; n27560_not
g56744 not n34616 ; n34616_not
g56745 not n34427 ; n34427_not
g56746 not n42428 ; n42428_not
g56747 not n17417 ; n17417_not
g56748 not n48107 ; n48107_not
g56749 not n28622 ; n28622_not
g56750 not n33257 ; n33257_not
g56751 not n32546 ; n32546_not
g56752 not n35192 ; n35192_not
g56753 not n33248 ; n33248_not
g56754 not n16049 ; n16049_not
g56755 not n47333 ; n47333_not
g56756 not n26462 ; n26462_not
g56757 not n34607 ; n34607_not
g56758 not n14654 ; n14654_not
g56759 not n10685 ; n10685_not
g56760 not n34418 ; n34418_not
g56761 not n31808 ; n31808_not
g56762 not n32528 ; n32528_not
g56763 not n16643 ; n16643_not
g56764 not n25535 ; n25535_not
g56765 not n47324 ; n47324_not
g56766 not n29333 ; n29333_not
g56767 not n26543 ; n26543_not
g56768 not n34058 ; n34058_not
g56769 not n10658 ; n10658_not
g56770 not n10775 ; n10775_not
g56771 not n33275 ; n33275_not
g56772 not n28604 ; n28604_not
g56773 not n17408 ; n17408_not
g56774 not n26804 ; n26804_not
g56775 not n25616 ; n25616_not
g56776 not n25715 ; n25715_not
g56777 not n13862 ; n13862_not
g56778 not n26417 ; n26417_not
g56779 not n17327 ; n17327_not
g56780 not n28451 ; n28451_not
g56781 not n35732 ; n35732_not
g56782 not n15950 ; n15950_not
g56783 not n26561 ; n26561_not
g56784 not n31952 ; n31952_not
g56785 not n29108 ; n29108_not
g56786 not n35741 ; n35741_not
g56787 not n34724 ; n34724_not
g56788 not n47090 ; n47090_not
g56789 not n16616 ; n16616_not
g56790 not n15464 ; n15464_not
g56791 not n25733 ; n25733_not
g56792 not n17309 ; n17309_not
g56793 not n17804 ; n17804_not
g56794 not n34760 ; n34760_not
g56795 not n34742 ; n34742_not
g56796 not n15941 ; n15941_not
g56797 not n32285 ; n32285_not
g56798 not n35714 ; n35714_not
g56799 not n14339 ; n14339_not
g56800 not n28433 ; n28433_not
g56801 not n35723 ; n35723_not
g56802 not n27317 ; n27317_not
g56803 not n29117 ; n29117_not
g56804 not n25724 ; n25724_not
g56805 not n14249 ; n14249_not
g56806 not n14924 ; n14924_not
g56807 not n17237 ; n17237_not
g56808 not n26435 ; n26435_not
g56809 not n16274 ; n16274_not
g56810 not n34715 ; n34715_not
g56811 not n33347 ; n33347_not
g56812 not n42482 ; n42482_not
g56813 not n47360 ; n47360_not
g56814 not n13556 ; n13556_not
g56815 not n25607 ; n25607_not
g56816 not n10667 ; n10667_not
g56817 not n28523 ; n28523_not
g56818 not n41852 ; n41852_not
g56819 not n32762 ; n32762_not
g56820 not n26912 ; n26912_not
g56821 not n28541 ; n28541_not
g56822 not n31907 ; n31907_not
g56823 not n47171 ; n47171_not
g56824 not n28460 ; n28460_not
g56825 not n21674 ; n21674_not
g56826 not n19433 ; n19433_not
g56827 not n33383 ; n33383_not
g56828 not n16607 ; n16607_not
g56829 not n15095 ; n15095_not
g56830 not n35831 ; n35831_not
g56831 not n14546 ; n14546_not
g56832 not n25652 ; n25652_not
g56833 not n35840 ; n35840_not
g56834 not n23078 ; n23078_not
g56835 not n15086 ; n15086_not
g56836 not n14528 ; n14528_not
g56837 not n41447 ; n41447_not
g56838 not n33365 ; n33365_not
g56839 not n15608 ; n15608_not
g56840 not n28505 ; n28505_not
g56841 not n25328 ; n25328_not
g56842 not n33068 ; n33068_not
g56843 not n48314 ; n48314_not
g56844 not n14285 ; n14285_not
g56845 not n10595 ; n10595_not
g56846 not n25319 ; n25319_not
g56847 not n17552 ; n17552_not
g56848 not n27047 ; n27047_not
g56849 not n10577 ; n10577_not
g56850 not n17561 ; n17561_not
g56851 not n27056 ; n27056_not
g56852 not n13844 ; n13844_not
g56853 not n34517 ; n34517_not
g56854 not n27065 ; n27065_not
g56855 not n14708 ; n14708_not
g56856 not n43175 ; n43175_not
g56857 not n15815 ; n15815_not
g56858 not n27038 ; n27038_not
g56859 not n25373 ; n25373_not
g56860 not n42194 ; n42194_not
g56861 not n41654 ; n41654_not
g56862 not n13493 ; n13493_not
g56863 not n13673 ; n13673_not
g56864 not n43058 ; n43058_not
g56865 not n16553 ; n16553_not
g56866 not n25355 ; n25355_not
g56867 not n35156 ; n35156_not
g56868 not n27137 ; n27137_not
g56869 not n14537 ; n14537_not
g56870 not n26372 ; n26372_not
g56871 not n14465 ; n14465_not
g56872 not n17525 ; n17525_not
g56873 not n29252 ; n29252_not
g56874 not n32780 ; n32780_not
g56875 not n28910 ; n28910_not
g56876 not n32960 ; n32960_not
g56877 not n16139 ; n16139_not
g56878 not n25175 ; n25175_not
g56879 not n34508 ; n34508_not
g56880 not n27092 ; n27092_not
g56881 not n16148 ; n16148_not
g56882 not n42185 ; n42185_not
g56883 not n32915 ; n32915_not
g56884 not n40628 ; n40628_not
g56885 not n14438 ; n14438_not
g56886 not n42077 ; n42077_not
g56887 not n15671 ; n15671_not
g56888 not n25256 ; n25256_not
g56889 not n42464 ; n42464_not
g56890 not n16184 ; n16184_not
g56891 not n17246 ; n17246_not
g56892 not n14681 ; n14681_not
g56893 not n36065 ; n36065_not
g56894 not n36056 ; n36056_not
g56895 not n27128 ; n27128_not
g56896 not n48053 ; n48053_not
g56897 not n41618 ; n41618_not
g56898 not n34094 ; n34094_not
g56899 not n32573 ; n32573_not
g56900 not n32852 ; n32852_not
g56901 not n26507 ; n26507_not
g56902 not n35543 ; n35543_not
g56903 not n32870 ; n32870_not
g56904 not n27191 ; n27191_not
g56905 not n32429 ; n32429_not
g56906 not n16544 ; n16544_not
g56907 not n16247 ; n16247_not
g56908 not n11477 ; n11477_not
g56909 not n35174 ; n35174_not
g56910 not n42905 ; n42905_not
g56911 not n14834 ; n14834_not
g56912 not n25445 ; n25445_not
g56913 not n16067 ; n16067_not
g56914 not n26525 ; n26525_not
g56915 not n26471 ; n26471_not
g56916 not n32834 ; n32834_not
g56917 not n14591 ; n14591_not
g56918 not n14825 ; n14825_not
g56919 not n17471 ; n17471_not
g56920 not n41690 ; n41690_not
g56921 not n27209 ; n27209_not
g56922 not n16526 ; n16526_not
g56923 not n42806 ; n42806_not
g56924 not n13448 ; n13448_not
g56925 not n42815 ; n42815_not
g56926 not n47342 ; n47342_not
g56927 not n34445 ; n34445_not
g56928 not n47126 ; n47126_not
g56929 not n48116 ; n48116_not
g56930 not n34454 ; n34454_not
g56931 not n15644 ; n15644_not
g56932 not n31844 ; n31844_not
g56933 not n14861 ; n14861_not
g56934 not n32384 ; n32384_not
g56935 not n34544 ; n34544_not
g56936 not n29036 ; n29036_not
g56937 not n29018 ; n29018_not
g56938 not n28811 ; n28811_not
g56939 not n42068 ; n42068_not
g56940 not n36038 ; n36038_not
g56941 not n14276 ; n14276_not
g56942 not n14771 ; n14771_not
g56943 not n32843 ; n32843_not
g56944 not n10793 ; n10793_not
g56945 not n29009 ; n29009_not
g56946 not n15653 ; n15653_not
g56947 not n44435 ; n44435_not
g56948 not n14294 ; n14294_not
g56949 not n27146 ; n27146_not
g56950 not n36047 ; n36047_not
g56951 not n33095 ; n33095_not
g56952 not n34490 ; n34490_not
g56953 not n10874 ; n10874_not
g56954 not n29027 ; n29027_not
g56955 not n33185 ; n33185_not
g56956 not n25418 ; n25418_not
g56957 not n34535 ; n34535_not
g56958 not n35147 ; n35147_not
g56959 not n13853 ; n13853_not
g56960 not n17480 ; n17480_not
g56961 not n16229 ; n16229_not
g56962 not n34481 ; n34481_not
g56963 not n33167 ; n33167_not
g56964 not n15662 ; n15662_not
g56965 not n26480 ; n26480_not
g56966 not n42932 ; n42932_not
g56967 not n41663 ; n41663_not
g56968 not n28802 ; n28802_not
g56969 not n27713 ; n27713_not
g56970 not n26084 ; n26084_not
g56971 not n27506 ; n27506_not
g56972 not n15806 ; n15806_not
g56973 not n29720 ; n29720_not
g56974 not n28073 ; n28073_not
g56975 not n42536 ; n42536_not
g56976 not n28082 ; n28082_not
g56977 not n29405 ; n29405_not
g56978 not n26066 ; n26066_not
g56979 not n27605 ; n27605_not
g56980 not n43355 ; n43355_not
g56981 not n28091 ; n28091_not
g56982 not n13736 ; n13736_not
g56983 not n32681 ; n32681_not
g56984 not n32483 ; n32483_not
g56985 not n42518 ; n42518_not
g56986 not n16931 ; n16931_not
g56987 not n28037 ; n28037_not
g56988 not n16382 ; n16382_not
g56989 not n41843 ; n41843_not
g56990 not n42554 ; n42554_not
g56991 not n40637 ; n40637_not
g56992 not n35318 ; n35318_not
g56993 not n28046 ; n28046_not
g56994 not n43067 ; n43067_not
g56995 not n26093 ; n26093_not
g56996 not n16814 ; n16814_not
g56997 not n15482 ; n15482_not
g56998 not n29207 ; n29207_not
g56999 not n35327 ; n35327_not
g57000 not n41834 ; n41834_not
g57001 not n28064 ; n28064_not
g57002 not n15572 ; n15572_not
g57003 not n13709 ; n13709_not
g57004 not n27461 ; n27461_not
g57005 not n15824 ; n15824_not
g57006 not n34283 ; n34283_not
g57007 not n28136 ; n28136_not
g57008 not n15833 ; n15833_not
g57009 not n35354 ; n35354_not
g57010 not n28127 ; n28127_not
g57011 not n15581 ; n15581_not
g57012 not n10757 ; n10757_not
g57013 not n28163 ; n28163_not
g57014 not n47630 ; n47630_not
g57015 not n47405 ; n47405_not
g57016 not n10829 ; n10829_not
g57017 not n27335 ; n27335_not
g57018 not n26048 ; n26048_not
g57019 not n13727 ; n13727_not
g57020 not n34274 ; n34274_not
g57021 not n44480 ; n44480_not
g57022 not n27470 ; n27470_not
g57023 not n15455 ; n15455_not
g57024 not n26714 ; n26714_not
g57025 not n44444 ; n44444_not
g57026 not n13772 ; n13772_not
g57027 not n17039 ; n17039_not
g57028 not n15446 ; n15446_not
g57029 not n40619 ; n40619_not
g57030 not n28109 ; n28109_not
g57031 not n15428 ; n15428_not
g57032 not n26732 ; n26732_not
g57033 not n14393 ; n14393_not
g57034 not n43346 ; n43346_not
g57035 not n33761 ; n33761_not
g57036 not n26633 ; n26633_not
g57037 not n16436 ; n16436_not
g57038 not n42455 ; n42455_not
g57039 not n26192 ; n26192_not
g57040 not n13754 ; n13754_not
g57041 not n32645 ; n32645_not
g57042 not n26183 ; n26183_not
g57043 not n15770 ; n15770_not
g57044 not n13880 ; n13880_not
g57045 not n26651 ; n26651_not
g57046 not n27902 ; n27902_not
g57047 not n35066 ; n35066_not
g57048 not n16805 ; n16805_not
g57049 not n26615 ; n26615_not
g57050 not n16463 ; n16463_not
g57051 not n16454 ; n16454_not
g57052 not n32636 ; n32636_not
g57053 not n32294 ; n32294_not
g57054 not n15761 ; n15761_not
g57055 not n47414 ; n47414_not
g57056 not n15554 ; n15554_not
g57057 not n15563 ; n15563_not
g57058 not n27803 ; n27803_not
g57059 not n33572 ; n33572_not
g57060 not n33770 ; n33770_not
g57061 not n33518 ; n33518_not
g57062 not n32195 ; n32195_not
g57063 not n16760 ; n16760_not
g57064 not n15527 ; n15527_not
g57065 not n41744 ; n41744_not
g57066 not n26138 ; n26138_not
g57067 not n33671 ; n33671_not
g57068 not n15518 ; n15518_not
g57069 not n41861 ; n41861_not
g57070 not n15734 ; n15734_not
g57071 not n28019 ; n28019_not
g57072 not n14384 ; n14384_not
g57073 not n28028 ; n28028_not
g57074 not n33833 ; n33833_not
g57075 not n32492 ; n32492_not
g57076 not n26660 ; n26660_not
g57077 not n26174 ; n26174_not
g57078 not n35039 ; n35039_not
g57079 not n26237 ; n26237_not
g57080 not n41906 ; n41906_not
g57081 not n35273 ; n35273_not
g57082 not n26255 ; n26255_not
g57083 not n34166 ; n34166_not
g57084 not n40952 ; n40952_not
g57085 not n33716 ; n33716_not
g57086 not n13745 ; n13745_not
g57087 not n26156 ; n26156_not
g57088 not n32654 ; n32654_not
g57089 not n16904 ; n16904_not
g57090 not n34337 ; n34337_not
g57091 not n25841 ; n25841_not
g57092 not n31970 ; n31970_not
g57093 not n28352 ; n28352_not
g57094 not n27362 ; n27362_not
g57095 not n16328 ; n16328_not
g57096 not n26381 ; n26381_not
g57097 not n42275 ; n42275_not
g57098 not n28361 ; n28361_not
g57099 not n33455 ; n33455_not
g57100 not n35219 ; n35219_not
g57101 not n28370 ; n28370_not
g57102 not n35615 ; n35615_not
g57103 not n15194 ; n15194_not
g57104 not n14492 ; n14492_not
g57105 not n27353 ; n27353_not
g57106 not n35237 ; n35237_not
g57107 not n29144 ; n29144_not
g57108 not n26570 ; n26570_not
g57109 not n15239 ; n15239_not
g57110 not n41735 ; n41735_not
g57111 not n28334 ; n28334_not
g57112 not n35552 ; n35552_not
g57113 not n13637 ; n13637_not
g57114 not n15923 ; n15923_not
g57115 not n25850 ; n25850_not
g57116 not n42086 ; n42086_not
g57117 not n29135 ; n29135_not
g57118 not n33482 ; n33482_not
g57119 not n17282 ; n17282_not
g57120 not n34364 ; n34364_not
g57121 not n41726 ; n41726_not
g57122 not n15158 ; n15158_not
g57123 not n43409 ; n43409_not
g57124 not n25760 ; n25760_not
g57125 not n25625 ; n25625_not
g57126 not n47801 ; n47801_not
g57127 not n25751 ; n25751_not
g57128 not n28415 ; n28415_not
g57129 not n15149 ; n15149_not
g57130 not n27326 ; n27326_not
g57131 not n16634 ; n16634_not
g57132 not n13817 ; n13817_not
g57133 not n28262 ; n28262_not
g57134 not n15932 ; n15932_not
g57135 not n27281 ; n27281_not
g57136 not n15185 ; n15185_not
g57137 not n29126 ; n29126_not
g57138 not n35624 ; n35624_not
g57139 not n10568 ; n10568_not
g57140 not n34814 ; n34814_not
g57141 not n17255 ; n17255_not
g57142 not n48224 ; n48224_not
g57143 not n41771 ; n41771_not
g57144 not n15509 ; n15509_not
g57145 not n16940 ; n16940_not
g57146 not n26327 ; n26327_not
g57147 not n27344 ; n27344_not
g57148 not n42662 ; n42662_not
g57149 not n27425 ; n27425_not
g57150 not n14366 ; n14366_not
g57151 not n16670 ; n16670_not
g57152 not n44426 ; n44426_not
g57153 not n15347 ; n15347_not
g57154 not n27416 ; n27416_not
g57155 not n35426 ; n35426_not
g57156 not n27614 ; n27614_not
g57157 not n13916 ; n13916_not
g57158 not n17156 ; n17156_not
g57159 not n32717 ; n32717_not
g57160 not n28226 ; n28226_not
g57161 not n15329 ; n15329_not
g57162 not n10766 ; n10766_not
g57163 not n27407 ; n27407_not
g57164 not n15374 ; n15374_not
g57165 not n35363 ; n35363_not
g57166 not n16724 ; n16724_not
g57167 not n28181 ; n28181_not
g57168 not n16355 ; n16355_not
g57169 not n35246 ; n35246_not
g57170 not n27434 ; n27434_not
g57171 not n35075 ; n35075_not
g57172 not n42329 ; n42329_not
g57173 not n40178 ; n40178_not
g57174 not n25913 ; n25913_not
g57175 not n43373 ; n43373_not
g57176 not n42617 ; n42617_not
g57177 not n27308 ; n27308_not
g57178 not n15356 ; n15356_not
g57179 not n35381 ; n35381_not
g57180 not n35390 ; n35390_not
g57181 not n15266 ; n15266_not
g57182 not n16706 ; n16706_not
g57183 not n13781 ; n13781_not
g57184 not n28307 ; n28307_not
g57185 not n27830 ; n27830_not
g57186 not n15248 ; n15248_not
g57187 not n35507 ; n35507_not
g57188 not n27623 ; n27623_not
g57189 not n27632 ; n27632_not
g57190 not n28325 ; n28325_not
g57191 not n42284 ; n42284_not
g57192 not n42761 ; n42761_not
g57193 not n32078 ; n32078_not
g57194 not n35525 ; n35525_not
g57195 not n34832 ; n34832_not
g57196 not n34328 ; n34328_not
g57197 not n29153 ; n29153_not
g57198 not n13691 ; n13691_not
g57199 not n42635 ; n42635_not
g57200 not n29810 ; n29810_not
g57201 not n34049 ; n34049_not
g57202 not n33428 ; n33428_not
g57203 not n28271 ; n28271_not
g57204 not n34850 ; n34850_not
g57205 not n15284 ; n15284_not
g57206 not n16337 ; n16337_not
g57207 not n14672 ; n14672_not
g57208 not n25922 ; n25922_not
g57209 not n35462 ; n35462_not
g57210 not n42293 ; n42293_not
g57211 not n35471 ; n35471_not
g57212 not n31736 ; n31736_not
g57213 not n20675 ; n20675_not
g57214 not n37901 ; n37901_not
g57215 not n23483 ; n23483_not
g57216 not n11864 ; n11864_not
g57217 not n22079 ; n22079_not
g57218 not n24329 ; n24329_not
g57219 not n20657 ; n20657_not
g57220 not n18434 ; n18434_not
g57221 not n18506 ; n18506_not
g57222 not n20648 ; n20648_not
g57223 not n46091 ; n46091_not
g57224 not n44048 ; n44048_not
g57225 not n31727 ; n31727_not
g57226 not n43841 ; n43841_not
g57227 not n22709 ; n22709_not
g57228 not n11882 ; n11882_not
g57229 not n39206 ; n39206_not
g57230 not n31547 ; n31547_not
g57231 not n23465 ; n23465_not
g57232 not n18452 ; n18452_not
g57233 not n17363 ; n17363_not
g57234 not n22736 ; n22736_not
g57235 not n24392 ; n24392_not
g57236 not n36650 ; n36650_not
g57237 not n24383 ; n24383_not
g57238 not n38414 ; n38414_not
g57239 not n30890 ; n30890_not
g57240 not n43715 ; n43715_not
g57241 not n24347 ; n24347_not
g57242 not n39404 ; n39404_not
g57243 not n31178 ; n31178_not
g57244 not n12296 ; n12296_not
g57245 not n24356 ; n24356_not
g57246 not n23474 ; n23474_not
g57247 not n44606 ; n44606_not
g57248 not n19154 ; n19154_not
g57249 not n18560 ; n18560_not
g57250 not n42527 ; n42527_not
g57251 not n24257 ; n24257_not
g57252 not n24248 ; n24248_not
g57253 not n19145 ; n19145_not
g57254 not n36713 ; n36713_not
g57255 not n24239 ; n24239_not
g57256 not n38612 ; n38612_not
g57257 not n23519 ; n23519_not
g57258 not n44039 ; n44039_not
g57259 not n40925 ; n40925_not
g57260 not n43580 ; n43580_not
g57261 not n12953 ; n12953_not
g57262 not n37604 ; n37604_not
g57263 not n40880 ; n40880_not
g57264 not n36740 ; n36740_not
g57265 not n30368 ; n30368_not
g57266 not n18524 ; n18524_not
g57267 not n48530 ; n48530_not
g57268 not n24293 ; n24293_not
g57269 not n24284 ; n24284_not
g57270 not n11891 ; n11891_not
g57271 not n30593 ; n30593_not
g57272 not n12971 ; n12971_not
g57273 not n46811 ; n46811_not
g57274 not n31664 ; n31664_not
g57275 not n20594 ; n20594_not
g57276 not n40943 ; n40943_not
g57277 not n24266 ; n24266_not
g57278 not n18551 ; n18551_not
g57279 not n24590 ; n24590_not
g57280 not n37532 ; n37532_not
g57281 not n21935 ; n21935_not
g57282 not n40349 ; n40349_not
g57283 not n19244 ; n19244_not
g57284 not n24581 ; n24581_not
g57285 not n43490 ; n43490_not
g57286 not n47027 ; n47027_not
g57287 not n40907 ; n40907_not
g57288 not n36380 ; n36380_not
g57289 not n36425 ; n36425_not
g57290 not n22763 ; n22763_not
g57291 not n21962 ; n21962_not
g57292 not n18281 ; n18281_not
g57293 not n10928 ; n10928_not
g57294 not n31655 ; n31655_not
g57295 not n38036 ; n38036_not
g57296 not n24554 ; n24554_not
g57297 not n21971 ; n21971_not
g57298 not n24635 ; n24635_not
g57299 not n18227 ; n18227_not
g57300 not n37235 ; n37235_not
g57301 not n36506 ; n36506_not
g57302 not n37523 ; n37523_not
g57303 not n23384 ; n23384_not
g57304 not n18236 ; n18236_not
g57305 not n38072 ; n38072_not
g57306 not n18263 ; n18263_not
g57307 not n24608 ; n24608_not
g57308 not n19262 ; n19262_not
g57309 not n18272 ; n18272_not
g57310 not n19181 ; n19181_not
g57311 not n20837 ; n20837_not
g57312 not n11783 ; n11783_not
g57313 not n19253 ; n19253_not
g57314 not n36524 ; n36524_not
g57315 not n11792 ; n11792_not
g57316 not n20747 ; n20747_not
g57317 not n31196 ; n31196_not
g57318 not n11828 ; n11828_not
g57319 not n20738 ; n20738_not
g57320 not n13097 ; n13097_not
g57321 not n37550 ; n37550_not
g57322 not n41078 ; n41078_not
g57323 not n38504 ; n38504_not
g57324 not n13088 ; n13088_not
g57325 not n36623 ; n36623_not
g57326 not n30278 ; n30278_not
g57327 not n40367 ; n40367_not
g57328 not n24437 ; n24437_not
g57329 not n38513 ; n38513_not
g57330 not n46055 ; n46055_not
g57331 not n36632 ; n36632_not
g57332 not n31187 ; n31187_not
g57333 not n30287 ; n30287_not
g57334 not n43517 ; n43517_not
g57335 not n36416 ; n36416_not
g57336 not n24545 ; n24545_not
g57337 not n18326 ; n18326_not
g57338 not n41087 ; n41087_not
g57339 not n24536 ; n24536_not
g57340 not n21926 ; n21926_not
g57341 not n37226 ; n37226_not
g57342 not n23438 ; n23438_not
g57343 not n30269 ; n30269_not
g57344 not n23447 ; n23447_not
g57345 not n19190 ; n19190_not
g57346 not n41096 ; n41096_not
g57347 not n24491 ; n24491_not
g57348 not n23456 ; n23456_not
g57349 not n23717 ; n23717_not
g57350 not n36902 ; n36902_not
g57351 not n40727 ; n40727_not
g57352 not n18902 ; n18902_not
g57353 not n11990 ; n11990_not
g57354 not n22376 ; n22376_not
g57355 not n10487 ; n10487_not
g57356 not n31493 ; n31493_not
g57357 not n22538 ; n22538_not
g57358 not n37703 ; n37703_not
g57359 not n22394 ; n22394_not
g57360 not n12629 ; n12629_not
g57361 not n39107 ; n39107_not
g57362 not n30476 ; n30476_not
g57363 not n46226 ; n46226_not
g57364 not n40556 ; n40556_not
g57365 not n40745 ; n40745_not
g57366 not n20369 ; n20369_not
g57367 not n22565 ; n22565_not
g57368 not n40736 ; n40736_not
g57369 not n18731 ; n18731_not
g57370 not n40484 ; n40484_not
g57371 not n45326 ; n45326_not
g57372 not n40493 ; n40493_not
g57373 not n37118 ; n37118_not
g57374 not n30449 ; n30449_not
g57375 not n36911 ; n36911_not
g57376 not n23690 ; n23690_not
g57377 not n22349 ; n22349_not
g57378 not n30548 ; n30548_not
g57379 not n40529 ; n40529_not
g57380 not n12773 ; n12773_not
g57381 not n39062 ; n39062_not
g57382 not n23834 ; n23834_not
g57383 not n37055 ; n37055_not
g57384 not n22457 ; n22457_not
g57385 not n12836 ; n12836_not
g57386 not n46271 ; n46271_not
g57387 not n45218 ; n45218_not
g57388 not n12098 ; n12098_not
g57389 not n23825 ; n23825_not
g57390 not n22475 ; n22475_not
g57391 not n30494 ; n30494_not
g57392 not n23780 ; n23780_not
g57393 not n40592 ; n40592_not
g57394 not n22484 ; n22484_not
g57395 not n11189 ; n11189_not
g57396 not n31475 ; n31475_not
g57397 not n40682 ; n40682_not
g57398 not n20198 ; n20198_not
g57399 not n20189 ; n20189_not
g57400 not n40664 ; n40664_not
g57401 not n17183 ; n17183_not
g57402 not n43652 ; n43652_not
g57403 not n40655 ; n40655_not
g57404 not n12089 ; n12089_not
g57405 not n45191 ; n45191_not
g57406 not n30458 ; n30458_not
g57407 not n12791 ; n12791_not
g57408 not n23852 ; n23852_not
g57409 not n39080 ; n39080_not
g57410 not n46262 ; n46262_not
g57411 not n23861 ; n23861_not
g57412 not n40646 ; n40646_not
g57413 not n22196 ; n22196_not
g57414 not n30854 ; n30854_not
g57415 not n31673 ; n31673_not
g57416 not n23933 ; n23933_not
g57417 not n22655 ; n22655_not
g57418 not n19082 ; n19082_not
g57419 not n37154 ; n37154_not
g57420 not n18641 ; n18641_not
g57421 not n10298 ; n10298_not
g57422 not n19073 ; n19073_not
g57423 not n39251 ; n39251_not
g57424 not n30395 ; n30395_not
g57425 not n12566 ; n12566_not
g57426 not n40790 ; n40790_not
g57427 not n38801 ; n38801_not
g57428 not n23609 ; n23609_not
g57429 not n22628 ; n22628_not
g57430 not n12719 ; n12719_not
g57431 not n24194 ; n24194_not
g57432 not n12269 ; n12269_not
g57433 not n36803 ; n36803_not
g57434 not n38702 ; n38702_not
g57435 not n24185 ; n24185_not
g57436 not n39314 ; n39314_not
g57437 not n12944 ; n12944_not
g57438 not n24176 ; n24176_not
g57439 not n40862 ; n40862_not
g57440 not n24158 ; n24158_not
g57441 not n23546 ; n23546_not
g57442 not n22178 ; n22178_not
g57443 not n24149 ; n24149_not
g57444 not n11288 ; n11288_not
g57445 not n40817 ; n40817_not
g57446 not n43733 ; n43733_not
g57447 not n19019 ; n19019_not
g57448 not n40457 ; n40457_not
g57449 not n37073 ; n37073_not
g57450 not n40763 ; n40763_not
g57451 not n43940 ; n43940_not
g57452 not n22295 ; n22295_not
g57453 not n37631 ; n37631_not
g57454 not n39413 ; n39413_not
g57455 not n30953 ; n30953_not
g57456 not n24059 ; n24059_not
g57457 not n40754 ; n40754_not
g57458 not n39170 ; n39170_not
g57459 not n18704 ; n18704_not
g57460 not n37127 ; n37127_not
g57461 not n20477 ; n20477_not
g57462 not n19910 ; n19910_not
g57463 not n31718 ; n31718_not
g57464 not n46181 ; n46181_not
g57465 not n23924 ; n23924_not
g57466 not n22619 ; n22619_not
g57467 not n39215 ; n39215_not
g57468 not n36830 ; n36830_not
g57469 not n24095 ; n24095_not
g57470 not n38810 ; n38810_not
g57471 not n23636 ; n23636_not
g57472 not n24086 ; n24086_not
g57473 not n40376 ; n40376_not
g57474 not n19028 ; n19028_not
g57475 not n23645 ; n23645_not
g57476 not n19640 ; n19640_not
g57477 not n43850 ; n43850_not
g57478 not n13376 ; n13376_not
g57479 not n44561 ; n44561_not
g57480 not n12584 ; n12584_not
g57481 not n41294 ; n41294_not
g57482 not n21197 ; n21197_not
g57483 not n22934 ; n22934_not
g57484 not n37415 ; n37415_not
g57485 not n40079 ; n40079_not
g57486 not n21188 ; n21188_not
g57487 not n41267 ; n41267_not
g57488 not n21629 ; n21629_not
g57489 not n45119 ; n45119_not
g57490 not n36227 ; n36227_not
g57491 not n17291 ; n17291_not
g57492 not n45164 ; n45164_not
g57493 not n41348 ; n41348_not
g57494 not n21593 ; n21593_not
g57495 not n17903 ; n17903_not
g57496 not n45155 ; n45155_not
g57497 not n22961 ; n22961_not
g57498 not n48341 ; n48341_not
g57499 not n39602 ; n39602_not
g57500 not n22952 ; n22952_not
g57501 not n37406 ; n37406_not
g57502 not n31628 ; n31628_not
g57503 not n38270 ; n38270_not
g57504 not n44309 ; n44309_not
g57505 not n18056 ; n18056_not
g57506 not n45560 ; n45560_not
g57507 not n30683 ; n30683_not
g57508 not n30674 ; n30674_not
g57509 not n11567 ; n11567_not
g57510 not n36290 ; n36290_not
g57511 not n21692 ; n21692_not
g57512 not n21089 ; n21089_not
g57513 not n38153 ; n38153_not
g57514 not n31286 ; n31286_not
g57515 not n12395 ; n12395_not
g57516 not n45902 ; n45902_not
g57517 not n30656 ; n30656_not
g57518 not n39710 ; n39710_not
g57519 not n36317 ; n36317_not
g57520 not n44381 ; n44381_not
g57521 not n24860 ; n24860_not
g57522 not n23168 ; n23168_not
g57523 not n36236 ; n36236_not
g57524 not n18029 ; n18029_not
g57525 not n21179 ; n21179_not
g57526 not n18038 ; n18038_not
g57527 not n44291 ; n44291_not
g57528 not n22925 ; n22925_not
g57529 not n19541 ; n19541_not
g57530 not n11387 ; n11387_not
g57531 not n30692 ; n30692_not
g57532 not n23186 ; n23186_not
g57533 not n11558 ; n11558_not
g57534 not n38180 ; n38180_not
g57535 not n21665 ; n21665_not
g57536 not n39530 ; n39530_not
g57537 not n17705 ; n17705_not
g57538 not n25193 ; n25193_not
g57539 not n17714 ; n17714_not
g57540 not n25139 ; n25139_not
g57541 not n39800 ; n39800_not
g57542 not n36128 ; n36128_not
g57543 not n45740 ; n45740_not
g57544 not n17084 ; n17084_not
g57545 not n21485 ; n21485_not
g57546 not n25166 ; n25166_not
g57547 not n17732 ; n17732_not
g57548 not n45731 ; n45731_not
g57549 not n30728 ; n30728_not
g57550 not n12485 ; n12485_not
g57551 not n17741 ; n17741_not
g57552 not n19712 ; n19712_not
g57553 not n30764 ; n30764_not
g57554 not n17606 ; n17606_not
g57555 not n17615 ; n17615_not
g57556 not n25247 ; n25247_not
g57557 not n41591 ; n41591_not
g57558 not n16751 ; n16751_not
g57559 not n21458 ; n21458_not
g57560 not n30746 ; n30746_not
g57561 not n17660 ; n17660_not
g57562 not n10883 ; n10883_not
g57563 not n12449 ; n12449_not
g57564 not n21467 ; n21467_not
g57565 not n39701 ; n39701_not
g57566 not n41555 ; n41555_not
g57567 not n44552 ; n44552_not
g57568 not n31817 ; n31817_not
g57569 not n46424 ; n46424_not
g57570 not n38234 ; n38234_not
g57571 not n41519 ; n41519_not
g57572 not n17813 ; n17813_not
g57573 not n23096 ; n23096_not
g57574 not n36164 ; n36164_not
g57575 not n25067 ; n25067_not
g57576 not n13385 ; n13385_not
g57577 not n25058 ; n25058_not
g57578 not n21287 ; n21287_not
g57579 not n38252 ; n38252_not
g57580 not n21566 ; n21566_not
g57581 not n41393 ; n41393_not
g57582 not n12557 ; n12557_not
g57583 not n21269 ; n21269_not
g57584 not n47117 ; n47117_not
g57585 not n41375 ; n41375_not
g57586 not n11468 ; n11468_not
g57587 not n41366 ; n41366_not
g57588 not n38261 ; n38261_not
g57589 not n13394 ; n13394_not
g57590 not n37352 ; n37352_not
g57591 not n45812 ; n45812_not
g57592 not n43454 ; n43454_not
g57593 not n36146 ; n36146_not
g57594 not n38243 ; n38243_not
g57595 not n31367 ; n31367_not
g57596 not n12458 ; n12458_not
g57597 not n41456 ; n41456_not
g57598 not n41438 ; n41438_not
g57599 not n41429 ; n41429_not
g57600 not n44165 ; n44165_not
g57601 not n45704 ; n45704_not
g57602 not n36155 ; n36155_not
g57603 not n21548 ; n21548_not
g57604 not n39611 ; n39611_not
g57605 not n38342 ; n38342_not
g57606 not n41195 ; n41195_not
g57607 not n40286 ; n40286_not
g57608 not n19361 ; n19361_not
g57609 not n20909 ; n20909_not
g57610 not n12359 ; n12359_not
g57611 not n21827 ; n21827_not
g57612 not n11738 ; n11738_not
g57613 not n24743 ; n24743_not
g57614 not n39503 ; n39503_not
g57615 not n24770 ; n24770_not
g57616 not n47063 ; n47063_not
g57617 not n43913 ; n43913_not
g57618 not n12656 ; n12656_not
g57619 not n21809 ; n21809_not
g57620 not n20963 ; n20963_not
g57621 not n30638 ; n30638_not
g57622 not n19370 ; n19370_not
g57623 not n40259 ; n40259_not
g57624 not n38117 ; n38117_not
g57625 not n21791 ; n21791_not
g57626 not n30179 ; n30179_not
g57627 not n36362 ; n36362_not
g57628 not n19406 ; n19406_not
g57629 not n18137 ; n18137_not
g57630 not n36353 ; n36353_not
g57631 not n24806 ; n24806_not
g57632 not n43904 ; n43904_not
g57633 not n22871 ; n22871_not
g57634 not n31259 ; n31259_not
g57635 not n18119 ; n18119_not
g57636 not n23249 ; n23249_not
g57637 not n21881 ; n21881_not
g57638 not n23375 ; n23375_not
g57639 not n38360 ; n38360_not
g57640 not n44318 ; n44318_not
g57641 not n46370 ; n46370_not
g57642 not n18191 ; n18191_not
g57643 not n36470 ; n36470_not
g57644 not n23348 ; n23348_not
g57645 not n21854 ; n21854_not
g57646 not n48422 ; n48422_not
g57647 not n19811 ; n19811_not
g57648 not n24680 ; n24680_not
g57649 not n48413 ; n48413_not
g57650 not n20891 ; n20891_not
g57651 not n30863 ; n30863_not
g57652 not n13286 ; n13286_not
g57653 not n21845 ; n21845_not
g57654 not n46514 ; n46514_not
g57655 not n36443 ; n36443_not
g57656 not n19352 ; n19352_not
g57657 not n43481 ; n43481_not
g57658 not n21836 ; n21836_not
g57659 not n37505 ; n37505_not
g57660 not n36434 ; n36434_not
g57661 not n24725 ; n24725_not
g57662 not n40187 ; n40187_not
g57663 not n44129 ; n44129_not
g57664 not n36344 ; n36344_not
g57665 not n38063 ; n38063_not
g57666 not n24851 ; n24851_not
g57667 not n38630 ; n38630_not
g57668 not n36335 ; n36335_not
g57669 not n18092 ; n18092_not
g57670 not n12386 ; n12386_not
g57671 not n24824 ; n24824_not
g57672 not n31763 ; n31763_not
g57673 not n22808 ; n22808_not
g57674 not n30647 ; n30647_not
g57675 not n23276 ; n23276_not
g57676 not n24815 ; n24815_not
g57677 not n18083 ; n18083_not
g57678 not n27345 ; n27345_not
g57679 not n39072 ; n39072_not
g57680 not n22854 ; n22854_not
g57681 not n22908 ; n22908_not
g57682 not n15582 ; n15582_not
g57683 not n27570 ; n27570_not
g57684 not n39126 ; n39126_not
g57685 not n37515 ; n37515_not
g57686 not n33960 ; n33960_not
g57687 not n17625 ; n17625_not
g57688 not n27435 ; n27435_not
g57689 not n27840 ; n27840_not
g57690 not n39432 ; n39432_not
g57691 not n39621 ; n39621_not
g57692 not n27354 ; n27354_not
g57693 not n43914 ; n43914_not
g57694 not n20559 ; n20559_not
g57695 not n27804 ; n27804_not
g57696 not n22548 ; n22548_not
g57697 not n27426 ; n27426_not
g57698 not n40863 ; n40863_not
g57699 not n16635 ; n16635_not
g57700 not n22818 ; n22818_not
g57701 not n34185 ; n34185_not
g57702 not n12396 ; n12396_not
g57703 not n12468 ; n12468_not
g57704 not n31494 ; n31494_not
g57705 not n30972 ; n30972_not
g57706 not n39333 ; n39333_not
g57707 not n10659 ; n10659_not
g57708 not n34194 ; n34194_not
g57709 not n31557 ; n31557_not
g57710 not n29307 ; n29307_not
g57711 not n27750 ; n27750_not
g57712 not n14358 ; n14358_not
g57713 not n39513 ; n39513_not
g57714 not n45903 ; n45903_not
g57715 not n39612 ; n39612_not
g57716 not n15852 ; n15852_not
g57717 not n33870 ; n33870_not
g57718 not n32619 ; n32619_not
g57719 not n31485 ; n31485_not
g57720 not n37218 ; n37218_not
g57721 not n22791 ; n22791_not
g57722 not n38514 ; n38514_not
g57723 not n29280 ; n29280_not
g57724 not n22773 ; n22773_not
g57725 not n14196 ; n14196_not
g57726 not n44283 ; n44283_not
g57727 not n33852 ; n33852_not
g57728 not n15771 ; n15771_not
g57729 not n27444 ; n27444_not
g57730 not n10983 ; n10983_not
g57731 not n31629 ; n31629_not
g57732 not n29361 ; n29361_not
g57733 not n37641 ; n37641_not
g57734 not n22494 ; n22494_not
g57735 not n19821 ; n19821_not
g57736 not n27453 ; n27453_not
g57737 not n39522 ; n39522_not
g57738 not n39324 ; n39324_not
g57739 not n33933 ; n33933_not
g57740 not n37407 ; n37407_not
g57741 not n44571 ; n44571_not
g57742 not n16653 ; n16653_not
g57743 not n27642 ; n27642_not
g57744 not n33924 ; n33924_not
g57745 not n19470 ; n19470_not
g57746 not n30756 ; n30756_not
g57747 not n33915 ; n33915_not
g57748 not n48090 ; n48090_not
g57749 not n10749 ; n10749_not
g57750 not n15933 ; n15933_not
g57751 not n48360 ; n48360_not
g57752 not n33906 ; n33906_not
g57753 not n32538 ; n32538_not
g57754 not n37533 ; n37533_not
g57755 not n27651 ; n27651_not
g57756 not n34365 ; n34365_not
g57757 not n15762 ; n15762_not
g57758 not n31593 ; n31593_not
g57759 not n44256 ; n44256_not
g57760 not n30873 ; n30873_not
g57761 not n16644 ; n16644_not
g57762 not n14268 ; n14268_not
g57763 not n22863 ; n22863_not
g57764 not n30828 ; n30828_not
g57765 not n42474 ; n42474_not
g57766 not n34257 ; n34257_not
g57767 not n44292 ; n44292_not
g57768 not n42357 ; n42357_not
g57769 not n19902 ; n19902_not
g57770 not n22746 ; n22746_not
g57771 not n39225 ; n39225_not
g57772 not n30792 ; n30792_not
g57773 not n15816 ; n15816_not
g57774 not n14295 ; n14295_not
g57775 not n37443 ; n37443_not
g57776 not n15672 ; n15672_not
g57777 not n16743 ; n16743_not
g57778 not n22872 ; n22872_not
g57779 not n29343 ; n29343_not
g57780 not n44274 ; n44274_not
g57781 not n37452 ; n37452_not
g57782 not n15681 ; n15681_not
g57783 not n34149 ; n34149_not
g57784 not n46335 ; n46335_not
g57785 not n22674 ; n22674_not
g57786 not n39270 ; n39270_not
g57787 not n15861 ; n15861_not
g57788 not n22665 ; n22665_not
g57789 not n27615 ; n27615_not
g57790 not n34086 ; n34086_not
g57791 not n43941 ; n43941_not
g57792 not n15726 ; n15726_not
g57793 not n27219 ; n27219_not
g57794 not n43860 ; n43860_not
g57795 not n27705 ; n27705_not
g57796 not n44238 ; n44238_not
g57797 not n44418 ; n44418_not
g57798 not n39450 ; n39450_not
g57799 not n42294 ; n42294_not
g57800 not n37173 ; n37173_not
g57801 not n30855 ; n30855_not
g57802 not n34167 ; n34167_not
g57803 not n22584 ; n22584_not
g57804 not n15708 ; n15708_not
g57805 not n30819 ; n30819_not
g57806 not n29433 ; n29433_not
g57807 not n14349 ; n14349_not
g57808 not n42366 ; n42366_not
g57809 not n43950 ; n43950_not
g57810 not n30783 ; n30783_not
g57811 not n27507 ; n27507_not
g57812 not n43815 ; n43815_not
g57813 not n14259 ; n14259_not
g57814 not n15627 ; n15627_not
g57815 not n29316 ; n29316_not
g57816 not n15591 ; n15591_not
g57817 not n30909 ; n30909_not
g57818 not n19803 ; n19803_not
g57819 not n15753 ; n15753_not
g57820 not n39162 ; n39162_not
g57821 not n47415 ; n47415_not
g57822 not n27372 ; n27372_not
g57823 not n42456 ; n42456_not
g57824 not n12369 ; n12369_not
g57825 not n12288 ; n12288_not
g57826 not n29325 ; n29325_not
g57827 not n15636 ; n15636_not
g57828 not n42447 ; n42447_not
g57829 not n27390 ; n27390_not
g57830 not n12189 ; n12189_not
g57831 not n43923 ; n43923_not
g57832 not n15690 ; n15690_not
g57833 not n15915 ; n15915_not
g57834 not n15735 ; n15735_not
g57835 not n27381 ; n27381_not
g57836 not n37425 ; n37425_not
g57837 not n47442 ; n47442_not
g57838 not n30954 ; n30954_not
g57839 not n15609 ; n15609_not
g57840 not n16941 ; n16941_not
g57841 not n15744 ; n15744_not
g57842 not n22593 ; n22593_not
g57843 not n22755 ; n22755_not
g57844 not n29370 ; n29370_not
g57845 not n27624 ; n27624_not
g57846 not n38127 ; n38127_not
g57847 not n38325 ; n38325_not
g57848 not n14556 ; n14556_not
g57849 not n20973 ; n20973_not
g57850 not n20928 ; n20928_not
g57851 not n42771 ; n42771_not
g57852 not n42762 ; n42762_not
g57853 not n14970 ; n14970_not
g57854 not n11739 ; n11739_not
g57855 not n20937 ; n20937_not
g57856 not n32727 ; n32727_not
g57857 not n48072 ; n48072_not
g57858 not n14961 ; n14961_not
g57859 not n42735 ; n42735_not
g57860 not n10677 ; n10677_not
g57861 not n32781 ; n32781_not
g57862 not n21837 ; n21837_not
g57863 not n20865 ; n20865_not
g57864 not n33339 ; n33339_not
g57865 not n28551 ; n28551_not
g57866 not n29082 ; n29082_not
g57867 not n42717 ; n42717_not
g57868 not n11649 ; n11649_not
g57869 not n42528 ; n42528_not
g57870 not n20991 ; n20991_not
g57871 not n38145 ; n38145_not
g57872 not n14916 ; n14916_not
g57873 not n38316 ; n38316_not
g57874 not n38082 ; n38082_not
g57875 not n43077 ; n43077_not
g57876 not n14565 ; n14565_not
g57877 not n16275 ; n16275_not
g57878 not n28632 ; n28632_not
g57879 not n29055 ; n29055_not
g57880 not n11667 ; n11667_not
g57881 not n21765 ; n21765_not
g57882 not n14925 ; n14925_not
g57883 not n21774 ; n21774_not
g57884 not n42780 ; n42780_not
g57885 not n33276 ; n33276_not
g57886 not n32817 ; n32817_not
g57887 not n28614 ; n28614_not
g57888 not n14934 ; n14934_not
g57889 not n28605 ; n28605_not
g57890 not n11685 ; n11685_not
g57891 not n43752 ; n43752_not
g57892 not n33375 ; n33375_not
g57893 not n11784 ; n11784_not
g57894 not n15096 ; n15096_not
g57895 not n28470 ; n28470_not
g57896 not n46029 ; n46029_not
g57897 not n14439 ; n14439_not
g57898 not n20838 ; n20838_not
g57899 not n28920 ; n28920_not
g57900 not n21936 ; n21936_not
g57901 not n38415 ; n38415_not
g57902 not n21945 ; n21945_not
g57903 not n21954 ; n21954_not
g57904 not n48702 ; n48702_not
g57905 not n21963 ; n21963_not
g57906 not n20775 ; n20775_not
g57907 not n28416 ; n28416_not
g57908 not n28542 ; n28542_not
g57909 not n33348 ; n33348_not
g57910 not n38352 ; n38352_not
g57911 not n44094 ; n44094_not
g57912 not n11757 ; n11757_not
g57913 not n28524 ; n28524_not
g57914 not n21864 ; n21864_not
g57915 not n20874 ; n20874_not
g57916 not n11766 ; n11766_not
g57917 not n28515 ; n28515_not
g57918 not n42690 ; n42690_not
g57919 not n38361 ; n38361_not
g57920 not n15069 ; n15069_not
g57921 not n28443 ; n28443_not
g57922 not n33357 ; n33357_not
g57923 not n38370 ; n38370_not
g57924 not n15078 ; n15078_not
g57925 not n44085 ; n44085_not
g57926 not n21891 ; n21891_not
g57927 not n21378 ; n21378_not
g57928 not n21369 ; n21369_not
g57929 not n45813 ; n45813_not
g57930 not n14718 ; n14718_not
g57931 not n14466 ; n14466_not
g57932 not n48045 ; n48045_not
g57933 not n21297 ; n21297_not
g57934 not n33078 ; n33078_not
g57935 not n21558 ; n21558_not
g57936 not n14754 ; n14754_not
g57937 not n33087 ; n33087_not
g57938 not n45822 ; n45822_not
g57939 not n10695 ; n10695_not
g57940 not n38217 ; n38217_not
g57941 not n11487 ; n11487_not
g57942 not n14763 ; n14763_not
g57943 not n28830 ; n28830_not
g57944 not n10686 ; n10686_not
g57945 not n42339 ; n42339_not
g57946 not n42951 ; n42951_not
g57947 not n14457 ; n14457_not
g57948 not n31386 ; n31386_not
g57949 not n21459 ; n21459_not
g57950 not n32925 ; n32925_not
g57951 not n45750 ; n45750_not
g57952 not n32916 ; n32916_not
g57953 not n38235 ; n38235_not
g57954 not n48063 ; n48063_not
g57955 not n14664 ; n14664_not
g57956 not n32754 ; n32754_not
g57957 not n32862 ; n32862_not
g57958 not n45732 ; n45732_not
g57959 not n19434 ; n19434_not
g57960 not n14691 ; n14691_not
g57961 not n21387 ; n21387_not
g57962 not n21657 ; n21657_not
g57963 not n21666 ; n21666_not
g57964 not n28740 ; n28740_not
g57965 not n14826 ; n14826_not
g57966 not n42906 ; n42906_not
g57967 not n28722 ; n28722_not
g57968 not n28713 ; n28713_not
g57969 not n38163 ; n38163_not
g57970 not n21693 ; n21693_not
g57971 not n42843 ; n42843_not
g57972 not n14862 ; n14862_not
g57973 not n31278 ; n31278_not
g57974 not n29046 ; n29046_not
g57975 not n31269 ; n31269_not
g57976 not n14583 ; n14583_not
g57977 not n21729 ; n21729_not
g57978 not n38307 ; n38307_not
g57979 not n42960 ; n42960_not
g57980 not n43068 ; n43068_not
g57981 not n14781 ; n14781_not
g57982 not n28812 ; n28812_not
g57983 not n42933 ; n42933_not
g57984 not n14637 ; n14637_not
g57985 not n19146 ; n19146_not
g57986 not n49143 ; n49143_not
g57987 not n14628 ; n14628_not
g57988 not n38280 ; n38280_not
g57989 not n21189 ; n21189_not
g57990 not n14808 ; n14808_not
g57991 not n42915 ; n42915_not
g57992 not n33168 ; n33168_not
g57993 not n44148 ; n44148_not
g57994 not n32745 ; n32745_not
g57995 not n33177 ; n33177_not
g57996 not n38190 ; n38190_not
g57997 not n39711 ; n39711_not
g57998 not n32673 ; n32673_not
g57999 not n29208 ; n29208_not
g58000 not n33465 ; n33465_not
g58001 not n47550 ; n47550_not
g58002 not n15465 ; n15465_not
g58003 not n37803 ; n37803_not
g58004 not n42564 ; n42564_not
g58005 not n20388 ; n20388_not
g58006 not n15474 ; n15474_not
g58007 not n15483 ; n15483_not
g58008 not n37740 ; n37740_not
g58009 not n15492 ; n15492_not
g58010 not n28038 ; n28038_not
g58011 not n47541 ; n47541_not
g58012 not n37731 ; n37731_not
g58013 not n42591 ; n42591_not
g58014 not n28146 ; n28146_not
g58015 not n46173 ; n46173_not
g58016 not n11928 ; n11928_not
g58017 not n29190 ; n29190_not
g58018 not n20469 ; n20469_not
g58019 not n14448 ; n14448_not
g58020 not n31449 ; n31449_not
g58021 not n32691 ; n32691_not
g58022 not n22269 ; n22269_not
g58023 not n15177 ; n15177_not
g58024 not n15438 ; n15438_not
g58025 not n15447 ; n15447_not
g58026 not n11973 ; n11973_not
g58027 not n22278 ; n22278_not
g58028 not n11982 ; n11982_not
g58029 not n33618 ; n33618_not
g58030 not n43806 ; n43806_not
g58031 not n22287 ; n22287_not
g58032 not n32475 ; n32475_not
g58033 not n20397 ; n20397_not
g58034 not n27741 ; n27741_not
g58035 not n32646 ; n32646_not
g58036 not n39018 ; n39018_not
g58037 not n46245 ; n46245_not
g58038 not n45246 ; n45246_not
g58039 not n29253 ; n29253_not
g58040 not n32466 ; n32466_not
g58041 not n33771 ; n33771_not
g58042 not n32637 ; n32637_not
g58043 not n45228 ; n45228_not
g58044 not n27930 ; n27930_not
g58045 not n27921 ; n27921_not
g58046 not n22458 ; n22458_not
g58047 not n22467 ; n22467_not
g58048 not n29262 ; n29262_not
g58049 not n27912 ; n27912_not
g58050 not n29271 ; n29271_not
g58051 not n39054 ; n39054_not
g58052 not n31476 ; n31476_not
g58053 not n46272 ; n46272_not
g58054 not n11199 ; n11199_not
g58055 not n33663 ; n33663_not
g58056 not n45318 ; n45318_not
g58057 not n32664 ; n32664_not
g58058 not n20298 ; n20298_not
g58059 not n20289 ; n20289_not
g58060 not n33654 ; n33654_not
g58061 not n22377 ; n22377_not
g58062 not n33708 ; n33708_not
g58063 not n15528 ; n15528_not
g58064 not n13665 ; n13665_not
g58065 not n22386 ; n22386_not
g58066 not n33564 ; n33564_not
g58067 not n15537 ; n15537_not
g58068 not n45291 ; n45291_not
g58069 not n46236 ; n46236_not
g58070 not n33753 ; n33753_not
g58071 not n44058 ; n44058_not
g58072 not n46065 ; n46065_not
g58073 not n11847 ; n11847_not
g58074 not n38550 ; n38550_not
g58075 not n33492 ; n33492_not
g58076 not n28236 ; n28236_not
g58077 not n42636 ; n42636_not
g58078 not n43581 ; n43581_not
g58079 not n37911 ; n37911_not
g58080 not n28335 ; n28335_not
g58081 not n29145 ; n29145_not
g58082 not n20667 ; n20667_not
g58083 not n38604 ; n38604_not
g58084 not n43563 ; n43563_not
g58085 not n11883 ; n11883_not
g58086 not n15276 ; n15276_not
g58087 not n28290 ; n28290_not
g58088 not n15294 ; n15294_not
g58089 not n46119 ; n46119_not
g58090 not n28407 ; n28407_not
g58091 not n39045 ; n39045_not
g58092 not n38442 ; n38442_not
g58093 not n20766 ; n20766_not
g58094 not n38028 ; n38028_not
g58095 not n21990 ; n21990_not
g58096 not n15186 ; n15186_not
g58097 not n38019 ; n38019_not
g58098 not n37722 ; n37722_not
g58099 not n33438 ; n33438_not
g58100 not n15195 ; n15195_not
g58101 not n28380 ; n28380_not
g58102 not n42654 ; n42654_not
g58103 not n31188 ; n31188_not
g58104 not n33447 ; n33447_not
g58105 not n11838 ; n11838_not
g58106 not n46056 ; n46056_not
g58107 not n28362 ; n28362_not
g58108 not n33474 ; n33474_not
g58109 not n38523 ; n38523_not
g58110 not n28353 ; n28353_not
g58111 not n11289 ; n11289_not
g58112 not n38703 ; n38703_not
g58113 not n29172 ; n29172_not
g58114 not n46164 ; n46164_not
g58115 not n15375 ; n15375_not
g58116 not n33609 ; n33609_not
g58117 not n38532 ; n38532_not
g58118 not n20496 ; n20496_not
g58119 not n42609 ; n42609_not
g58120 not n15384 ; n15384_not
g58121 not n20487 ; n20487_not
g58122 not n20478 ; n20478_not
g58123 not n42582 ; n42582_not
g58124 not n37623 ; n37623_not
g58125 not n38622 ; n38622_not
g58126 not n28263 ; n28263_not
g58127 not n29154 ; n29154_not
g58128 not n46137 ; n46137_not
g58129 not n17445 ; n17445_not
g58130 not n44229 ; n44229_not
g58131 not n28245 ; n28245_not
g58132 not n20577 ; n20577_not
g58133 not n38631 ; n38631_not
g58134 not n29163 ; n29163_not
g58135 not n47073 ; n47073_not
g58136 not n15348 ; n15348_not
g58137 not n28218 ; n28218_not
g58138 not n28209 ; n28209_not
g58139 not n37830 ; n37830_not
g58140 not n38640 ; n38640_not
g58141 not n11919 ; n11919_not
g58142 not n37821 ; n37821_not
g58143 not n48522 ; n48522_not
g58144 not n18525 ; n18525_not
g58145 not n10965 ; n10965_not
g58146 not n40890 ; n40890_not
g58147 not n10947 ; n10947_not
g58148 not n40665 ; n40665_not
g58149 not n41817 ; n41817_not
g58150 not n41808 ; n41808_not
g58151 not n35346 ; n35346_not
g58152 not n18480 ; n18480_not
g58153 not n26058 ; n26058_not
g58154 not n46911 ; n46911_not
g58155 not n26049 ; n26049_not
g58156 not n30297 ; n30297_not
g58157 not n24366 ; n24366_not
g58158 not n18471 ; n18471_not
g58159 not n10857 ; n10857_not
g58160 not n36660 ; n36660_not
g58161 not n18462 ; n18462_not
g58162 not n30279 ; n30279_not
g58163 not n36651 ; n36651_not
g58164 not n16851 ; n16851_not
g58165 not n36804 ; n36804_not
g58166 not n29730 ; n29730_not
g58167 not n16860 ; n16860_not
g58168 not n26184 ; n26184_not
g58169 not n40926 ; n40926_not
g58170 not n41907 ; n41907_not
g58171 not n18570 ; n18570_not
g58172 not n26175 ; n26175_not
g58173 not n36705 ; n36705_not
g58174 not n24258 ; n24258_not
g58175 not n26157 ; n26157_not
g58176 not n26148 ; n26148_not
g58177 not n16905 ; n16905_not
g58178 not n26076 ; n26076_not
g58179 not n18534 ; n18534_not
g58180 not n43347 ; n43347_not
g58181 not n12972 ; n12972_not
g58182 not n24285 ; n24285_not
g58183 not n40971 ; n40971_not
g58184 not n18345 ; n18345_not
g58185 not n18336 ; n18336_not
g58186 not n24537 ; n24537_not
g58187 not n41565 ; n41565_not
g58188 not n18291 ; n18291_not
g58189 not n24555 ; n24555_not
g58190 not n25914 ; n25914_not
g58191 not n35472 ; n35472_not
g58192 not n17175 ; n17175_not
g58193 not n32097 ; n32097_not
g58194 not n16716 ; n16716_not
g58195 not n17184 ; n17184_not
g58196 not n17193 ; n17193_not
g58197 not n35517 ; n35517_not
g58198 not n32079 ; n32079_not
g58199 not n43491 ; n43491_not
g58200 not n31728 ; n31728_not
g58201 not n36516 ; n36516_not
g58202 not n44364 ; n44364_not
g58203 not n35535 ; n35535_not
g58204 not n41790 ; n41790_not
g58205 not n43365 ; n43365_not
g58206 not n41781 ; n41781_not
g58207 not n36642 ; n36642_not
g58208 not n17094 ; n17094_not
g58209 not n18435 ; n18435_not
g58210 not n36633 ; n36633_not
g58211 not n35373 ; n35373_not
g58212 not n36615 ; n36615_not
g58213 not n41763 ; n41763_not
g58214 not n24483 ; n24483_not
g58215 not n36606 ; n36606_not
g58216 not n35418 ; n35418_not
g58217 not n18363 ; n18363_not
g58218 not n29811 ; n29811_not
g58219 not n18354 ; n18354_not
g58220 not n13692 ; n13692_not
g58221 not n18066 ; n18066_not
g58222 not n16608 ; n16608_not
g58223 not n16617 ; n16617_not
g58224 not n18147 ; n18147_not
g58225 not n46704 ; n46704_not
g58226 not n32088 ; n32088_not
g58227 not n10839 ; n10839_not
g58228 not n12882 ; n12882_not
g58229 not n40746 ; n40746_not
g58230 not n40755 ; n40755_not
g58231 not n44454 ; n44454_not
g58232 not n43608 ; n43608_not
g58233 not n16662 ; n16662_not
g58234 not n26373 ; n26373_not
g58235 not n35229 ; n35229_not
g58236 not n24078 ; n24078_not
g58237 not n44481 ; n44481_not
g58238 not n26355 ; n26355_not
g58239 not n26265 ; n26265_not
g58240 not n36921 ; n36921_not
g58241 not n43626 ; n43626_not
g58242 not n30459 ; n30459_not
g58243 not n26472 ; n26472_not
g58244 not n36930 ; n36930_not
g58245 not n26463 ; n26463_not
g58246 not n35193 ; n35193_not
g58247 not n12864 ; n12864_not
g58248 not n46632 ; n46632_not
g58249 not n16581 ; n16581_not
g58250 not n12873 ; n12873_not
g58251 not n46641 ; n46641_not
g58252 not n46650 ; n46650_not
g58253 not n26445 ; n26445_not
g58254 not n43572 ; n43572_not
g58255 not n16590 ; n16590_not
g58256 not n13827 ; n13827_not
g58257 not n18732 ; n18732_not
g58258 not n40818 ; n40818_not
g58259 not n40809 ; n40809_not
g58260 not n36813 ; n36813_not
g58261 not n41970 ; n41970_not
g58262 not n13764 ; n13764_not
g58263 not n26247 ; n26247_not
g58264 not n32196 ; n32196_not
g58265 not n26238 ; n26238_not
g58266 not n18615 ; n18615_not
g58267 not n18606 ; n18606_not
g58268 not n40845 ; n40845_not
g58269 not n40872 ; n40872_not
g58270 not n41925 ; n41925_not
g58271 not n26346 ; n26346_not
g58272 not n39414 ; n39414_not
g58273 not n43329 ; n43329_not
g58274 not n13782 ; n13782_not
g58275 not n10488 ; n10488_not
g58276 not n12918 ; n12918_not
g58277 not n48252 ; n48252_not
g58278 not n36822 ; n36822_not
g58279 not n16725 ; n16725_not
g58280 not n31719 ; n31719_not
g58281 not n29712 ; n29712_not
g58282 not n12909 ; n12909_not
g58283 not n10479 ; n10479_not
g58284 not n40791 ; n40791_not
g58285 not n12927 ; n12927_not
g58286 not n29721 ; n29721_not
g58287 not n35265 ; n35265_not
g58288 not n30387 ; n30387_not
g58289 not n47145 ; n47145_not
g58290 not n25482 ; n25482_not
g58291 not n13377 ; n13377_not
g58292 not n43419 ; n43419_not
g58293 not n17940 ; n17940_not
g58294 not n17931 ; n17931_not
g58295 not n13548 ; n13548_not
g58296 not n41682 ; n41682_not
g58297 not n17841 ; n17841_not
g58298 not n17913 ; n17913_not
g58299 not n44508 ; n44508_not
g58300 not n25455 ; n25455_not
g58301 not n36174 ; n36174_not
g58302 not n48333 ; n48333_not
g58303 not n25446 ; n25446_not
g58304 not n24960 ; n24960_not
g58305 not n25374 ; n25374_not
g58306 not n41394 ; n41394_not
g58307 not n25428 ; n25428_not
g58308 not n36273 ; n36273_not
g58309 not n25563 ; n25563_not
g58310 not n18048 ; n18048_not
g58311 not n36264 ; n36264_not
g58312 not n25554 ; n25554_not
g58313 not n17832 ; n17832_not
g58314 not n17373 ; n17373_not
g58315 not n31782 ; n31782_not
g58316 not n41691 ; n41691_not
g58317 not n13359 ; n13359_not
g58318 not n18039 ; n18039_not
g58319 not n36255 ; n36255_not
g58320 not n24924 ; n24924_not
g58321 not n25527 ; n25527_not
g58322 not n17166 ; n17166_not
g58323 not n36228 ; n36228_not
g58324 not n31863 ; n31863_not
g58325 not n25518 ; n25518_not
g58326 not n36219 ; n36219_not
g58327 not n25509 ; n25509_not
g58328 not n13368 ; n13368_not
g58329 not n31827 ; n31827_not
g58330 not n44544 ; n44544_not
g58331 not n41637 ; n41637_not
g58332 not n41493 ; n41493_not
g58333 not n25158 ; n25158_not
g58334 not n17544 ; n17544_not
g58335 not n10875 ; n10875_not
g58336 not n17742 ; n17742_not
g58337 not n13485 ; n13485_not
g58338 not n36075 ; n36075_not
g58339 not n25185 ; n25185_not
g58340 not n17715 ; n17715_not
g58341 not n13476 ; n13476_not
g58342 not n36084 ; n36084_not
g58343 not n41538 ; n41538_not
g58344 not n25284 ; n25284_not
g58345 not n36093 ; n36093_not
g58346 not n41556 ; n41556_not
g58347 not n41574 ; n41574_not
g58348 not n17319 ; n17319_not
g58349 not n25239 ; n25239_not
g58350 not n48315 ; n48315_not
g58351 not n25437 ; n25437_not
g58352 not n17472 ; n17472_not
g58353 not n25419 ; n25419_not
g58354 not n13386 ; n13386_not
g58355 not n41673 ; n41673_not
g58356 not n43455 ; n43455_not
g58357 not n41664 ; n41664_not
g58358 not n17823 ; n17823_not
g58359 not n17814 ; n17814_not
g58360 not n25095 ; n25095_not
g58361 not n36039 ; n36039_not
g58362 not n31809 ; n31809_not
g58363 not n13494 ; n13494_not
g58364 not n41466 ; n41466_not
g58365 not n41475 ; n41475_not
g58366 not n36147 ; n36147_not
g58367 not n17508 ; n17508_not
g58368 not n13395 ; n13395_not
g58369 not n25149 ; n25149_not
g58370 not n10866 ; n10866_not
g58371 not n35634 ; n35634_not
g58372 not n35580 ; n35580_not
g58373 not n18192 ; n18192_not
g58374 not n17265 ; n17265_not
g58375 not n43059 ; n43059_not
g58376 not n35652 ; n35652_not
g58377 not n13593 ; n13593_not
g58378 not n41187 ; n41187_not
g58379 not n36444 ; n36444_not
g58380 not n24447 ; n24447_not
g58381 not n31971 ; n31971_not
g58382 not n18183 ; n18183_not
g58383 not n25743 ; n25743_not
g58384 not n24744 ; n24744_not
g58385 not n13584 ; n13584_not
g58386 not n31746 ; n31746_not
g58387 not n24762 ; n24762_not
g58388 not n25860 ; n25860_not
g58389 not n35553 ; n35553_not
g58390 not n35562 ; n35562_not
g58391 not n18246 ; n18246_not
g58392 not n35544 ; n35544_not
g58393 not n24618 ; n24618_not
g58394 not n10497 ; n10497_not
g58395 not n13629 ; n13629_not
g58396 not n18237 ; n18237_not
g58397 not n35607 ; n35607_not
g58398 not n18228 ; n18228_not
g58399 not n48441 ; n48441_not
g58400 not n24645 ; n24645_not
g58401 not n41178 ; n41178_not
g58402 not n13278 ; n13278_not
g58403 not n17238 ; n17238_not
g58404 not n25806 ; n25806_not
g58405 not n47019 ; n47019_not
g58406 not n18174 ; n18174_not
g58407 not n36480 ; n36480_not
g58408 not n36462 ; n36462_not
g58409 not n35625 ; n35625_not
g58410 not n31926 ; n31926_not
g58411 not n36336 ; n36336_not
g58412 not n17355 ; n17355_not
g58413 not n25617 ; n25617_not
g58414 not n24843 ; n24843_not
g58415 not n17364 ; n17364_not
g58416 not n10893 ; n10893_not
g58417 not n25590 ; n25590_not
g58418 not n13557 ; n13557_not
g58419 not n25581 ; n25581_not
g58420 not n31908 ; n31908_not
g58421 not n44391 ; n44391_not
g58422 not n35931 ; n35931_not
g58423 not n24663 ; n24663_not
g58424 not n36390 ; n36390_not
g58425 not n29910 ; n29910_not
g58426 not n43464 ; n43464_not
g58427 not n16815 ; n16815_not
g58428 not n47181 ; n47181_not
g58429 not n43437 ; n43437_not
g58430 not n31962 ; n31962_not
g58431 not n35751 ; n35751_not
g58432 not n35760 ; n35760_not
g58433 not n31755 ; n31755_not
g58434 not n17337 ; n17337_not
g58435 not n31953 ; n31953_not
g58436 not n24672 ; n24672_not
g58437 not n24825 ; n24825_not
g58438 not n35841 ; n35841_not
g58439 not n25644 ; n25644_not
g58440 not n19209 ; n19209_not
g58441 not n40368 ; n40368_not
g58442 not n47316 ; n47316_not
g58443 not n34626 ; n34626_not
g58444 not n34653 ; n34653_not
g58445 not n26940 ; n26940_not
g58446 not n34662 ; n34662_not
g58447 not n47307 ; n47307_not
g58448 not n19182 ; n19182_not
g58449 not n16158 ; n16158_not
g58450 not n34707 ; n34707_not
g58451 not n26922 ; n26922_not
g58452 not n29550 ; n29550_not
g58453 not n23475 ; n23475_not
g58454 not n40377 ; n40377_not
g58455 not n47271 ; n47271_not
g58456 not n23484 ; n23484_not
g58457 not n37209 ; n37209_not
g58458 not n31665 ; n31665_not
g58459 not n19290 ; n19290_not
g58460 not n34527 ; n34527_not
g58461 not n23376 ; n23376_not
g58462 not n19281 ; n19281_not
g58463 not n23385 ; n23385_not
g58464 not n37236 ; n37236_not
g58465 not n16239 ; n16239_not
g58466 not n42159 ; n42159_not
g58467 not n23394 ; n23394_not
g58468 not n26742 ; n26742_not
g58469 not n43194 ; n43194_not
g58470 not n19254 ; n19254_not
g58471 not n34563 ; n34563_not
g58472 not n32385 ; n32385_not
g58473 not n19245 ; n19245_not
g58474 not n16257 ; n16257_not
g58475 not n19227 ; n19227_not
g58476 not n48603 ; n48603_not
g58477 not n37227 ; n37227_not
g58478 not n34635 ; n34635_not
g58479 not n37182 ; n37182_not
g58480 not n16329 ; n16329_not
g58481 not n19092 ; n19092_not
g58482 not n23583 ; n23583_not
g58483 not n12738 ; n12738_not
g58484 not n37155 ; n37155_not
g58485 not n47244 ; n47244_not
g58486 not n23619 ; n23619_not
g58487 not n13926 ; n13926_not
g58488 not n19047 ; n19047_not
g58489 not n23628 ; n23628_not
g58490 not n37146 ; n37146_not
g58491 not n23637 ; n23637_not
g58492 not n16347 ; n16347_not
g58493 not n23493 ; n23493_not
g58494 not n40386 ; n40386_not
g58495 not n34725 ; n34725_not
g58496 not n40395 ; n40395_not
g58497 not n47262 ; n47262_not
g58498 not n34743 ; n34743_not
g58499 not n19128 ; n19128_not
g58500 not n34752 ; n34752_not
g58501 not n34770 ; n34770_not
g58502 not n13953 ; n13953_not
g58503 not n26850 ; n26850_not
g58504 not n23529 ; n23529_not
g58505 not n34806 ; n34806_not
g58506 not n23538 ; n23538_not
g58507 not n37191 ; n37191_not
g58508 not n23556 ; n23556_not
g58509 not n26832 ; n26832_not
g58510 not n26823 ; n26823_not
g58511 not n23565 ; n23565_not
g58512 not n23574 ; n23574_not
g58513 not n14079 ; n14079_not
g58514 not n46461 ; n46461_not
g58515 not n14673 ; n14673_not
g58516 not n32439 ; n32439_not
g58517 not n45129 ; n45129_not
g58518 not n34437 ; n34437_not
g58519 not n44436 ; n44436_not
g58520 not n19425 ; n19425_not
g58521 not n16059 ; n16059_not
g58522 not n19614 ; n19614_not
g58523 not n31638 ; n31638_not
g58524 not n19605 ; n19605_not
g58525 not n27192 ; n27192_not
g58526 not n34464 ; n34464_not
g58527 not n23169 ; n23169_not
g58528 not n19551 ; n19551_not
g58529 not n16077 ; n16077_not
g58530 not n32457 ; n32457_not
g58531 not n27309 ; n27309_not
g58532 not n34374 ; n34374_not
g58533 not n29451 ; n29451_not
g58534 not n39801 ; n39801_not
g58535 not n12495 ; n12495_not
g58536 not n37317 ; n37317_not
g58537 not n39810 ; n39810_not
g58538 not n32448 ; n32448_not
g58539 not n19704 ; n19704_not
g58540 not n23079 ; n23079_not
g58541 not n23088 ; n23088_not
g58542 not n27255 ; n27255_not
g58543 not n39027 ; n39027_not
g58544 not n37308 ; n37308_not
g58545 not n23277 ; n23277_not
g58546 not n29505 ; n29505_not
g58547 not n19407 ; n19407_not
g58548 not n37272 ; n37272_not
g58549 not n43185 ; n43185_not
g58550 not n23295 ; n23295_not
g58551 not n29514 ; n29514_not
g58552 not n19371 ; n19371_not
g58553 not n19362 ; n19362_not
g58554 not n19344 ; n19344_not
g58555 not n16185 ; n16185_not
g58556 not n27057 ; n27057_not
g58557 not n42177 ; n42177_not
g58558 not n37254 ; n37254_not
g58559 not n12666 ; n12666_not
g58560 not n19335 ; n19335_not
g58561 not n42168 ; n42168_not
g58562 not n23358 ; n23358_not
g58563 not n27165 ; n27165_not
g58564 not n23196 ; n23196_not
g58565 not n37290 ; n37290_not
g58566 not n16086 ; n16086_not
g58567 not n46506 ; n46506_not
g58568 not n37281 ; n37281_not
g58569 not n19515 ; n19515_not
g58570 not n19506 ; n19506_not
g58571 not n40179 ; n40179_not
g58572 not n40188 ; n40188_not
g58573 not n27138 ; n27138_not
g58574 not n48621 ; n48621_not
g58575 not n27129 ; n27129_not
g58576 not n43176 ; n43176_not
g58577 not n12639 ; n12639_not
g58578 not n12648 ; n12648_not
g58579 not n42186 ; n42186_not
g58580 not n16419 ; n16419_not
g58581 not n16509 ; n16509_not
g58582 not n16437 ; n16437_not
g58583 not n37038 ; n37038_not
g58584 not n32259 ; n32259_not
g58585 not n34932 ; n34932_not
g58586 not n26625 ; n26625_not
g58587 not n40647 ; n40647_not
g58588 not n26526 ; n26526_not
g58589 not n46614 ; n46614_not
g58590 not n29622 ; n29622_not
g58591 not n16545 ; n16545_not
g58592 not n29442 ; n29442_not
g58593 not n40539 ; n40539_not
g58594 not n23781 ; n23781_not
g58595 not n16770 ; n16770_not
g58596 not n40494 ; n40494_not
g58597 not n26517 ; n26517_not
g58598 not n12846 ; n12846_not
g58599 not n32286 ; n32286_not
g58600 not n37074 ; n37074_not
g58601 not n48117 ; n48117_not
g58602 not n23844 ; n23844_not
g58603 not n42087 ; n42087_not
g58604 not n46560 ; n46560_not
g58605 not n26652 ; n26652_not
g58606 not n23763 ; n23763_not
g58607 not n18921 ; n18921_not
g58608 not n23754 ; n23754_not
g58609 not n18912 ; n18912_not
g58610 not n23835 ; n23835_not
g58611 not n40638 ; n40638_not
g58612 not n47226 ; n47226_not
g58613 not n26580 ; n26580_not
g58614 not n26661 ; n26661_not
g58615 not n16428 ; n16428_not
g58616 not n13863 ; n13863_not
g58617 not n26634 ; n26634_not
g58618 not n13872 ; n13872_not
g58619 not n12783 ; n12783_not
g58620 not n35094 ; n35094_not
g58621 not n37047 ; n37047_not
g58622 not n23727 ; n23727_not
g58623 not n16563 ; n16563_not
g58624 not n35139 ; n35139_not
g58625 not n26724 ; n26724_not
g58626 not n12819 ; n12819_not
g58627 not n29613 ; n29613_not
g58628 not n31584 ; n31584_not
g58629 not n17157 ; n17157_not
g58630 not n43275 ; n43275_not
g58631 not n40584 ; n40584_not
g58632 not n34923 ; n34923_not
g58633 not n23925 ; n23925_not
g58634 not n12747 ; n12747_not
g58635 not n26490 ; n26490_not
g58636 not n29604 ; n29604_not
g58637 not n30468 ; n30468_not
g58638 not n16365 ; n16365_not
g58639 not n18813 ; n18813_not
g58640 not n40485 ; n40485_not
g58641 not n42096 ; n42096_not
g58642 not n26715 ; n26715_not
g58643 not n35148 ; n35148_not
g58644 not n40692 ; n40692_not
g58645 not n12855 ; n12855_not
g58646 not n26553 ; n26553_not
g58647 not n46623 ; n46623_not
g58648 not n23691 ; n23691_not
g58649 not n16374 ; n16374_not
g58650 not n12919 ; n12919_not
g58651 not n44383 ; n44383_not
g58652 not n31288 ; n31288_not
g58653 not n29407 ; n29407_not
g58654 not n10849 ; n10849_not
g58655 not n43753 ; n43753_not
g58656 not n32683 ; n32683_not
g58657 not n31765 ; n31765_not
g58658 not n31567 ; n31567_not
g58659 not n11956 ; n11956_not
g58660 not n31855 ; n31855_not
g58661 not n17851 ; n17851_not
g58662 not n10876 ; n10876_not
g58663 not n29416 ; n29416_not
g58664 not n48262 ; n48262_not
g58665 not n44158 ; n44158_not
g58666 not n43861 ; n43861_not
g58667 not n43771 ; n43771_not
g58668 not n31693 ; n31693_not
g58669 not n48640 ; n48640_not
g58670 not n13558 ; n13558_not
g58671 not n31891 ; n31891_not
g58672 not n31882 ; n31882_not
g58673 not n11965 ; n11965_not
g58674 not n30496 ; n30496_not
g58675 not n11587 ; n11587_not
g58676 not n31909 ; n31909_not
g58677 not n31297 ; n31297_not
g58678 not n29704 ; n29704_not
g58679 not n31783 ; n31783_not
g58680 not n43762 ; n43762_not
g58681 not n29272 ; n29272_not
g58682 not n30829 ; n30829_not
g58683 not n11569 ; n11569_not
g58684 not n31873 ; n31873_not
g58685 not n48550 ; n48550_not
g58686 not n31774 ; n31774_not
g58687 not n43744 ; n43744_not
g58688 not n32467 ; n32467_not
g58689 not n49144 ; n49144_not
g58690 not n43960 ; n43960_not
g58691 not n29245 ; n29245_not
g58692 not n30775 ; n30775_not
g58693 not n18076 ; n18076_not
g58694 not n43429 ; n43429_not
g58695 not n30766 ; n30766_not
g58696 not n44176 ; n44176_not
g58697 not n44185 ; n44185_not
g58698 not n43825 ; n43825_not
g58699 not n31378 ; n31378_not
g58700 not n13486 ; n13486_not
g58701 not n32872 ; n32872_not
g58702 not n43834 ; n43834_not
g58703 not n30469 ; n30469_not
g58704 not n13693 ; n13693_not
g58705 not n44194 ; n44194_not
g58706 not n32908 ; n32908_not
g58707 not n14674 ; n14674_not
g58708 not n32449 ; n32449_not
g58709 not n32917 ; n32917_not
g58710 not n31396 ; n31396_not
g58711 not n10885 ; n10885_not
g58712 not n30739 ; n30739_not
g58713 not n43447 ; n43447_not
g58714 not n13828 ; n13828_not
g58715 not n14449 ; n14449_not
g58716 not n12487 ; n12487_not
g58717 not n29443 ; n29443_not
g58718 not n32836 ; n32836_not
g58719 not n14629 ; n14629_not
g58720 not n32557 ; n32557_not
g58721 not n31648 ; n31648_not
g58722 not n43591 ; n43591_not
g58723 not n14638 ; n14638_not
g58724 not n48244 ; n48244_not
g58725 not n30667 ; n30667_not
g58726 not n30676 ; n30676_not
g58727 not n31585 ; n31585_not
g58728 not n43870 ; n43870_not
g58729 not n10759 ; n10759_not
g58730 not n13855 ; n13855_not
g58731 not n29650 ; n29650_not
g58732 not n43168 ; n43168_not
g58733 not n12892 ; n12892_not
g58734 not n11479 ; n11479_not
g58735 not n30487 ; n30487_not
g58736 not n14647 ; n14647_not
g58737 not n43807 ; n43807_not
g58738 not n48325 ; n48325_not
g58739 not n12838 ; n12838_not
g58740 not n30694 ; n30694_not
g58741 not n31468 ; n31468_not
g58742 not n31459 ; n31459_not
g58743 not n14458 ; n14458_not
g58744 not n43609 ; n43609_not
g58745 not n31837 ; n31837_not
g58746 not n31684 ; n31684_not
g58747 not n10948 ; n10948_not
g58748 not n32746 ; n32746_not
g58749 not n32539 ; n32539_not
g58750 not n32359 ; n32359_not
g58751 not n14539 ; n14539_not
g58752 not n44356 ; n44356_not
g58753 not n43573 ; n43573_not
g58754 not n13954 ; n13954_not
g58755 not n43348 ; n43348_not
g58756 not n13189 ; n13189_not
g58757 not n32719 ; n32719_not
g58758 not n11794 ; n11794_not
g58759 not n29740 ; n29740_not
g58760 not n32098 ; n32098_not
g58761 not n12757 ; n12757_not
g58762 not n14476 ; n14476_not
g58763 not n43096 ; n43096_not
g58764 not n43663 ; n43663_not
g58765 not n13279 ; n13279_not
g58766 not n13882 ; n13882_not
g58767 not n44266 ; n44266_not
g58768 not n42583 ; n42583_not
g58769 not n12298 ; n12298_not
g58770 not n32368 ; n32368_not
g58771 not n29164 ; n29164_not
g58772 not n12289 ; n12289_not
g58773 not n30595 ; n30595_not
g58774 not n32179 ; n32179_not
g58775 not n13963 ; n13963_not
g58776 not n29560 ; n29560_not
g58777 not n13639 ; n13639_not
g58778 not n31495 ; n31495_not
g58779 not n47029 ; n47029_not
g58780 not n48712 ; n48712_not
g58781 not n24385 ; n24385_not
g58782 not n42538 ; n42538_not
g58783 not n31675 ; n31675_not
g58784 not n30559 ; n30559_not
g58785 not n11875 ; n11875_not
g58786 not n30289 ; n30289_not
g58787 not n32584 ; n32584_not
g58788 not n43087 ; n43087_not
g58789 not n13738 ; n13738_not
g58790 not n12991 ; n12991_not
g58791 not n13729 ; n13729_not
g58792 not n12199 ; n12199_not
g58793 not n30955 ; n30955_not
g58794 not n13918 ; n13918_not
g58795 not n44248 ; n44248_not
g58796 not n30946 ; n30946_not
g58797 not n10957 ; n10957_not
g58798 not n48217 ; n48217_not
g58799 not n43384 ; n43384_not
g58800 not n41098 ; n41098_not
g58801 not n11893 ; n11893_not
g58802 not n30919 ; n30919_not
g58803 not n17059 ; n17059_not
g58804 not n30577 ; n30577_not
g58805 not n43933 ; n43933_not
g58806 not n29335 ; n29335_not
g58807 not n48154 ; n48154_not
g58808 not n31198 ; n31198_not
g58809 not n30928 ; n30928_not
g58810 not n29812 ; n29812_not
g58811 not n29803 ; n29803_not
g58812 not n43276 ; n43276_not
g58813 not n48514 ; n48514_not
g58814 not n30937 ; n30937_not
g58815 not n31738 ; n31738_not
g58816 not n29182 ; n29182_not
g58817 not n13990 ; n13990_not
g58818 not n32593 ; n32593_not
g58819 not n31945 ; n31945_not
g58820 not n14197 ; n14197_not
g58821 not n14557 ; n14557_not
g58822 not n12694 ; n12694_not
g58823 not n43645 ; n43645_not
g58824 not n14377 ; n14377_not
g58825 not n12937 ; n12937_not
g58826 not n12793 ; n12793_not
g58827 not n29065 ; n29065_not
g58828 not n11686 ; n11686_not
g58829 not n31549 ; n31549_not
g58830 not n30991 ; n30991_not
g58831 not n11938 ; n11938_not
g58832 not n29911 ; n29911_not
g58833 not n48127 ; n48127_not
g58834 not n32827 ; n32827_not
g58835 not n11596 ; n11596_not
g58836 not n13567 ; n13567_not
g58837 not n14584 ; n14584_not
g58838 not n43924 ; n43924_not
g58839 not n31558 ; n31558_not
g58840 not n29641 ; n29641_not
g58841 not n14467 ; n14467_not
g58842 not n43195 ; n43195_not
g58843 not n43069 ; n43069_not
g58844 not n13774 ; n13774_not
g58845 not n31936 ; n31936_not
g58846 not n48226 ; n48226_not
g58847 not n30883 ; n30883_not
g58848 not n43285 ; n43285_not
g58849 not n32773 ; n32773_not
g58850 not n32377 ; n32377_not
g58851 not n32188 ; n32188_not
g58852 not n43078 ; n43078_not
g58853 not n29632 ; n29632_not
g58854 not n29533 ; n29533_not
g58855 not n38443 ; n38443_not
g58856 not n14368 ; n14368_not
g58857 not n14179 ; n14179_not
g58858 not n13972 ; n13972_not
g58859 not n38434 ; n38434_not
g58860 not n31486 ; n31486_not
g58861 not n29524 ; n29524_not
g58862 not n29173 ; n29173_not
g58863 not n31963 ; n31963_not
g58864 not n44329 ; n44329_not
g58865 not n30982 ; n30982_not
g58866 not n43465 ; n43465_not
g58867 not n31747 ; n31747_not
g58868 not n29380 ; n29380_not
g58869 not n13297 ; n13297_not
g58870 not n29083 ; n29083_not
g58871 not n31972 ; n31972_not
g58872 not n32386 ; n32386_not
g58873 not n30199 ; n30199_not
g58874 not n17275 ; n17275_not
g58875 not n18544 ; n18544_not
g58876 not n40936 ; n40936_not
g58877 not n18382 ; n18382_not
g58878 not n40918 ; n40918_not
g58879 not n36742 ; n36742_not
g58880 not n36751 ; n36751_not
g58881 not n36535 ; n36535_not
g58882 not n24178 ; n24178_not
g58883 not n46714 ; n46714_not
g58884 not n18670 ; n18670_not
g58885 not n40783 ; n40783_not
g58886 not n36823 ; n36823_not
g58887 not n36832 ; n36832_not
g58888 not n40774 ; n40774_not
g58889 not n24088 ; n24088_not
g58890 not n24079 ; n24079_not
g58891 not n40738 ; n40738_not
g58892 not n36850 ; n36850_not
g58893 not n23962 ; n23962_not
g58894 not n18724 ; n18724_not
g58895 not n16690 ; n16690_not
g58896 not n46615 ; n46615_not
g58897 not n36319 ; n36319_not
g58898 not n36913 ; n36913_not
g58899 not n23980 ; n23980_not
g58900 not n36283 ; n36283_not
g58901 not n36904 ; n36904_not
g58902 not n36940 ; n36940_not
g58903 not n18751 ; n18751_not
g58904 not n18760 ; n18760_not
g58905 not n44644 ; n44644_not
g58906 not n24529 ; n24529_not
g58907 not n18364 ; n18364_not
g58908 not n18373 ; n18373_not
g58909 not n24484 ; n24484_not
g58910 not n24475 ; n24475_not
g58911 not n18427 ; n18427_not
g58912 not n24439 ; n24439_not
g58913 not n36634 ; n36634_not
g58914 not n18454 ; n18454_not
g58915 not n36643 ; n36643_not
g58916 not n18391 ; n18391_not
g58917 not n36661 ; n36661_not
g58918 not n40981 ; n40981_not
g58919 not n24376 ; n24376_not
g58920 not n40954 ; n40954_not
g58921 not n36706 ; n36706_not
g58922 not n18535 ; n18535_not
g58923 not n46831 ; n46831_not
g58924 not n18526 ; n18526_not
g58925 not n46903 ; n46903_not
g58926 not n18445 ; n18445_not
g58927 not n18508 ; n18508_not
g58928 not n40990 ; n40990_not
g58929 not n44617 ; n44617_not
g58930 not n18481 ; n18481_not
g58931 not n36670 ; n36670_not
g58932 not n18472 ; n18472_not
g58933 not n24367 ; n24367_not
g58934 not n23683 ; n23683_not
g58935 not n39640 ; n39640_not
g58936 not n18841 ; n18841_not
g58937 not n23692 ; n23692_not
g58938 not n23674 ; n23674_not
g58939 not n37129 ; n37129_not
g58940 not n40477 ; n40477_not
g58941 not n19039 ; n19039_not
g58942 not n19057 ; n19057_not
g58943 not n19066 ; n19066_not
g58944 not n44653 ; n44653_not
g58945 not n23593 ; n23593_not
g58946 not n37174 ; n37174_not
g58947 not n37192 ; n37192_not
g58948 not n18742 ; n18742_not
g58949 not n19129 ; n19129_not
g58950 not n19138 ; n19138_not
g58951 not n23287 ; n23287_not
g58952 not n19165 ; n19165_not
g58953 not n23494 ; n23494_not
g58954 not n19174 ; n19174_not
g58955 not n36562 ; n36562_not
g58956 not n37219 ; n37219_not
g58957 not n19219 ; n19219_not
g58958 not n19228 ; n19228_not
g58959 not n19237 ; n19237_not
g58960 not n19273 ; n19273_not
g58961 not n37246 ; n37246_not
g58962 not n19309 ; n19309_not
g58963 not n23917 ; n23917_not
g58964 not n40675 ; n40675_not
g58965 not n23908 ; n23908_not
g58966 not n40684 ; n40684_not
g58967 not n18814 ; n18814_not
g58968 not n23890 ; n23890_not
g58969 not n37039 ; n37039_not
g58970 not n23872 ; n23872_not
g58971 not n38641 ; n38641_not
g58972 not n16924 ; n16924_not
g58973 not n46552 ; n46552_not
g58974 not n23827 ; n23827_not
g58975 not n23818 ; n23818_not
g58976 not n23809 ; n23809_not
g58977 not n40567 ; n40567_not
g58978 not n23719 ; n23719_not
g58979 not n18931 ; n18931_not
g58980 not n23728 ; n23728_not
g58981 not n23737 ; n23737_not
g58982 not n46525 ; n46525_not
g58983 not n40549 ; n40549_not
g58984 not n23746 ; n23746_not
g58985 not n37066 ; n37066_not
g58986 not n23773 ; n23773_not
g58987 not n18904 ; n18904_not
g58988 not n37093 ; n37093_not
g58989 not n37084 ; n37084_not
g58990 not n23791 ; n23791_not
g58991 not n37075 ; n37075_not
g58992 not n17464 ; n17464_not
g58993 not n25447 ; n25447_not
g58994 not n25438 ; n25438_not
g58995 not n17473 ; n17473_not
g58996 not n41656 ; n41656_not
g58997 not n47128 ; n47128_not
g58998 not n36049 ; n36049_not
g58999 not n17167 ; n17167_not
g59000 not n25348 ; n25348_not
g59001 not n36067 ; n36067_not
g59002 not n17554 ; n17554_not
g59003 not n17563 ; n17563_not
g59004 not n25294 ; n25294_not
g59005 not n25285 ; n25285_not
g59006 not n25258 ; n25258_not
g59007 not n17626 ; n17626_not
g59008 not n17644 ; n17644_not
g59009 not n17653 ; n17653_not
g59010 not n40729 ; n40729_not
g59011 not n17068 ; n17068_not
g59012 not n41566 ; n41566_not
g59013 not n41548 ; n41548_not
g59014 not n17680 ; n17680_not
g59015 not n25195 ; n25195_not
g59016 not n17716 ; n17716_not
g59017 not n17752 ; n17752_not
g59018 not n36139 ; n36139_not
g59019 not n41458 ; n41458_not
g59020 not n35815 ; n35815_not
g59021 not n47164 ; n47164_not
g59022 not n35833 ; n35833_not
g59023 not n25645 ; n25645_not
g59024 not n35851 ; n35851_not
g59025 not n41719 ; n41719_not
g59026 not n17356 ; n17356_not
g59027 not n25609 ; n25609_not
g59028 not n47155 ; n47155_not
g59029 not n17365 ; n17365_not
g59030 not n35914 ; n35914_not
g59031 not n35923 ; n35923_not
g59032 not n35941 ; n35941_not
g59033 not n17374 ; n17374_not
g59034 not n25465 ; n25465_not
g59035 not n17455 ; n17455_not
g59036 not n25474 ; n25474_not
g59037 not n17194 ; n17194_not
g59038 not n25483 ; n25483_not
g59039 not n47137 ; n47137_not
g59040 not n41683 ; n41683_not
g59041 not n25492 ; n25492_not
g59042 not n35950 ; n35950_not
g59043 not n17428 ; n17428_not
g59044 not n47146 ; n47146_not
g59045 not n41692 ; n41692_not
g59046 not n25519 ; n25519_not
g59047 not n25528 ; n25528_not
g59048 not n25537 ; n25537_not
g59049 not n25546 ; n25546_not
g59050 not n24790 ; n24790_not
g59051 not n24763 ; n24763_not
g59052 not n36418 ; n36418_not
g59053 not n47056 ; n47056_not
g59054 not n24646 ; n24646_not
g59055 not n18175 ; n18175_not
g59056 not n36427 ; n36427_not
g59057 not n47047 ; n47047_not
g59058 not n36454 ; n36454_not
g59059 not n24691 ; n24691_not
g59060 not n36463 ; n36463_not
g59061 not n24664 ; n24664_not
g59062 not n36490 ; n36490_not
g59063 not n41179 ; n41179_not
g59064 not n24628 ; n24628_not
g59065 not n18247 ; n18247_not
g59066 not n18256 ; n18256_not
g59067 not n36508 ; n36508_not
g59068 not n36517 ; n36517_not
g59069 not n24583 ; n24583_not
g59070 not n24466 ; n24466_not
g59071 not n24574 ; n24574_not
g59072 not n36544 ; n36544_not
g59073 not n18274 ; n18274_not
g59074 not n36553 ; n36553_not
g59075 not n24565 ; n24565_not
g59076 not n17347 ; n17347_not
g59077 not n36580 ; n36580_not
g59078 not n24493 ; n24493_not
g59079 not n25096 ; n25096_not
g59080 not n36157 ; n36157_not
g59081 not n25069 ; n25069_not
g59082 not n17842 ; n17842_not
g59083 not n17833 ; n17833_not
g59084 not n41359 ; n41359_not
g59085 not n17923 ; n17923_not
g59086 not n36184 ; n36184_not
g59087 not n41287 ; n41287_not
g59088 not n41278 ; n41278_not
g59089 not n24961 ; n24961_not
g59090 not n36238 ; n36238_not
g59091 not n36247 ; n36247_not
g59092 not n36265 ; n36265_not
g59093 not n24736 ; n24736_not
g59094 not n24808 ; n24808_not
g59095 not n24826 ; n24826_not
g59096 not n24844 ; n24844_not
g59097 not n24853 ; n24853_not
g59098 not n44572 ; n44572_not
g59099 not n18058 ; n18058_not
g59100 not n36292 ; n36292_not
g59101 not n47083 ; n47083_not
g59102 not n36274 ; n36274_not
g59103 not n24907 ; n24907_not
g59104 not n24916 ; n24916_not
g59105 not n38533 ; n38533_not
g59106 not n46156 ; n46156_not
g59107 not n22189 ; n22189_not
g59108 not n37822 ; n37822_not
g59109 not n20578 ; n20578_not
g59110 not n20587 ; n20587_not
g59111 not n46129 ; n46129_not
g59112 not n20596 ; n20596_not
g59113 not n22099 ; n22099_not
g59114 not n20668 ; n20668_not
g59115 not n37903 ; n37903_not
g59116 not n20677 ; n20677_not
g59117 not n46084 ; n46084_not
g59118 not n46075 ; n46075_not
g59119 not n38524 ; n38524_not
g59120 not n38452 ; n38452_not
g59121 not n37921 ; n37921_not
g59122 not n38515 ; n38515_not
g59123 not n37930 ; n37930_not
g59124 not n46048 ; n46048_not
g59125 not n20758 ; n20758_not
g59126 not n21982 ; n21982_not
g59127 not n21973 ; n21973_not
g59128 not n20794 ; n20794_not
g59129 not n21928 ; n21928_not
g59130 not n38065 ; n38065_not
g59131 not n20839 ; n20839_not
g59132 not n38074 ; n38074_not
g59133 not n45184 ; n45184_not
g59134 not n38731 ; n38731_not
g59135 not n19921 ; n19921_not
g59136 not n39055 ; n39055_not
g59137 not n39046 ; n39046_not
g59138 not n37660 ; n37660_not
g59139 not n45238 ; n45238_not
g59140 not n39019 ; n39019_not
g59141 not n46246 ; n46246_not
g59142 not n37705 ; n37705_not
g59143 not n37723 ; n37723_not
g59144 not n46219 ; n46219_not
g59145 not n38920 ; n38920_not
g59146 not n45337 ; n45337_not
g59147 not n46174 ; n46174_not
g59148 not n34915 ; n34915_not
g59149 not n38803 ; n38803_not
g59150 not n38812 ; n38812_not
g59151 not n38821 ; n38821_not
g59152 not n37804 ; n37804_not
g59153 not n38830 ; n38830_not
g59154 not n38173 ; n38173_not
g59155 not n21658 ; n21658_not
g59156 not n21649 ; n21649_not
g59157 not n38191 ; n38191_not
g59158 not n38281 ; n38281_not
g59159 not n45841 ; n45841_not
g59160 not n45643 ; n45643_not
g59161 not n45823 ; n45823_not
g59162 not n45652 ; n45652_not
g59163 not n45661 ; n45661_not
g59164 not n21298 ; n21298_not
g59165 not n45634 ; n45634_not
g59166 not n38245 ; n38245_not
g59167 not n45706 ; n45706_not
g59168 not n45724 ; n45724_not
g59169 not n45733 ; n45733_not
g59170 not n21388 ; n21388_not
g59171 not n21478 ; n21478_not
g59172 not n21469 ; n21469_not
g59173 not n38371 ; n38371_not
g59174 not n21874 ; n21874_not
g59175 not n21865 ; n21865_not
g59176 not n38353 ; n38353_not
g59177 not n20884 ; n20884_not
g59178 not n21856 ; n21856_not
g59179 not n38344 ; n38344_not
g59180 not n21847 ; n21847_not
g59181 not n20929 ; n20929_not
g59182 not n38335 ; n38335_not
g59183 not n20956 ; n20956_not
g59184 not n20965 ; n20965_not
g59185 not n38119 ; n38119_not
g59186 not n45931 ; n45931_not
g59187 not n21784 ; n21784_not
g59188 not n20983 ; n20983_not
g59189 not n21676 ; n21676_not
g59190 not n38155 ; n38155_not
g59191 not n21739 ; n21739_not
g59192 not n45904 ; n45904_not
g59193 not n20992 ; n20992_not
g59194 not n21766 ; n21766_not
g59195 not n38083 ; n38083_not
g59196 not n46471 ; n46471_not
g59197 not n23089 ; n23089_not
g59198 not n37309 ; n37309_not
g59199 not n39820 ; n39820_not
g59200 not n39811 ; n39811_not
g59201 not n39802 ; n39802_not
g59202 not n19732 ; n19732_not
g59203 not n39721 ; n39721_not
g59204 not n39712 ; n39712_not
g59205 not n46435 ; n46435_not
g59206 not n39703 ; n39703_not
g59207 not n37327 ; n37327_not
g59208 not n46327 ; n46327_not
g59209 not n39613 ; n39613_not
g59210 not n37354 ; n37354_not
g59211 not n37228 ; n37228_not
g59212 not n37372 ; n37372_not
g59213 not n22972 ; n22972_not
g59214 not n37381 ; n37381_not
g59215 not n37390 ; n37390_not
g59216 not n22963 ; n22963_not
g59217 not n22954 ; n22954_not
g59218 not n39604 ; n39604_not
g59219 not n37408 ; n37408_not
g59220 not n22945 ; n22945_not
g59221 not n39550 ; n39550_not
g59222 not n39541 ; n39541_not
g59223 not n22936 ; n22936_not
g59224 not n39190 ; n39190_not
g59225 not n19318 ; n19318_not
g59226 not n19327 ; n19327_not
g59227 not n19345 ; n19345_not
g59228 not n40297 ; n40297_not
g59229 not n17329 ; n17329_not
g59230 not n44716 ; n44716_not
g59231 not n40279 ; n40279_not
g59232 not n19372 ; n19372_not
g59233 not n37255 ; n37255_not
g59234 not n23269 ; n23269_not
g59235 not n19426 ; n19426_not
g59236 not n19444 ; n19444_not
g59237 not n19453 ; n19453_not
g59238 not n45166 ; n45166_not
g59239 not n39145 ; n39145_not
g59240 not n19633 ; n19633_not
g59241 not n19624 ; n19624_not
g59242 not n19615 ; n19615_not
g59243 not n19606 ; n19606_not
g59244 not n19561 ; n19561_not
g59245 not n19534 ; n19534_not
g59246 not n23188 ; n23188_not
g59247 not n23179 ; n23179_not
g59248 not n46480 ; n46480_not
g59249 not n19525 ; n19525_not
g59250 not n46507 ; n46507_not
g59251 not n19390 ; n19390_not
g59252 not n37282 ; n37282_not
g59253 not n19462 ; n19462_not
g59254 not n39361 ; n39361_not
g59255 not n39352 ; n39352_not
g59256 not n46354 ; n46354_not
g59257 not n22693 ; n22693_not
g59258 not n39217 ; n39217_not
g59259 not n22675 ; n22675_not
g59260 not n39280 ; n39280_not
g59261 not n39271 ; n39271_not
g59262 not n39244 ; n39244_not
g59263 not n37615 ; n37615_not
g59264 not n22657 ; n22657_not
g59265 not n22648 ; n22648_not
g59266 not n39262 ; n39262_not
g59267 not n46309 ; n46309_not
g59268 not n39253 ; n39253_not
g59269 not n22639 ; n22639_not
g59270 not n39226 ; n39226_not
g59271 not n39208 ; n39208_not
g59272 not n38650 ; n38650_not
g59273 not n22594 ; n22594_not
g59274 not n39181 ; n39181_not
g59275 not n22576 ; n22576_not
g59276 not n22567 ; n22567_not
g59277 not n39154 ; n39154_not
g59278 not n39118 ; n39118_not
g59279 not n39082 ; n39082_not
g59280 not n22927 ; n22927_not
g59281 not n39532 ; n39532_not
g59282 not n22918 ; n22918_not
g59283 not n39523 ; n39523_not
g59284 not n37417 ; n37417_not
g59285 not n22909 ; n22909_not
g59286 not n19723 ; n19723_not
g59287 not n39514 ; n39514_not
g59288 not n22891 ; n22891_not
g59289 not n37435 ; n37435_not
g59290 not n46408 ; n46408_not
g59291 not n19804 ; n19804_not
g59292 not n37462 ; n37462_not
g59293 not n22855 ; n22855_not
g59294 not n39505 ; n39505_not
g59295 not n38425 ; n38425_not
g59296 not n39415 ; n39415_not
g59297 not n22729 ; n22729_not
g59298 not n22738 ; n22738_not
g59299 not n39433 ; n39433_not
g59300 not n37534 ; n37534_not
g59301 not n39460 ; n39460_not
g59302 not n37525 ; n37525_not
g59303 not n22792 ; n22792_not
g59304 not n37516 ; n37516_not
g59305 not n22819 ; n22819_not
g59306 not n22828 ; n22828_not
g59307 not n22837 ; n22837_not
g59308 not n15718 ; n15718_not
g59309 not n34159 ; n34159_not
g59310 not n42394 ; n42394_not
g59311 not n34177 ; n34177_not
g59312 not n27571 ; n27571_not
g59313 not n34195 ; n34195_not
g59314 not n27517 ; n27517_not
g59315 not n27544 ; n27544_not
g59316 not n15781 ; n15781_not
g59317 not n34249 ; n34249_not
g59318 not n42358 ; n42358_not
g59319 not n27490 ; n27490_not
g59320 not n27274 ; n27274_not
g59321 not n34267 ; n34267_not
g59322 not n27463 ; n27463_not
g59323 not n34276 ; n34276_not
g59324 not n15835 ; n15835_not
g59325 not n34285 ; n34285_not
g59326 not n15862 ; n15862_not
g59327 not n15880 ; n15880_not
g59328 not n27382 ; n27382_not
g59329 not n15925 ; n15925_not
g59330 not n42268 ; n42268_not
g59331 not n34384 ; n34384_not
g59332 not n34393 ; n34393_not
g59333 not n33952 ; n33952_not
g59334 not n33961 ; n33961_not
g59335 not n27823 ; n27823_not
g59336 not n33727 ; n33727_not
g59337 not n47515 ; n47515_not
g59338 not n47506 ; n47506_not
g59339 not n47470 ; n47470_not
g59340 not n47452 ; n47452_not
g59341 not n47443 ; n47443_not
g59342 not n42457 ; n42457_not
g59343 not n47434 ; n47434_not
g59344 not n27751 ; n27751_not
g59345 not n15637 ; n15637_not
g59346 not n42484 ; n42484_not
g59347 not n27733 ; n27733_not
g59348 not n27706 ; n27706_not
g59349 not n15664 ; n15664_not
g59350 not n34087 ; n34087_not
g59351 not n47425 ; n47425_not
g59352 not n15673 ; n15673_not
g59353 not n15682 ; n15682_not
g59354 not n15691 ; n15691_not
g59355 not n27553 ; n27553_not
g59356 not n15709 ; n15709_not
g59357 not n27634 ; n27634_not
g59358 not n27625 ; n27625_not
g59359 not n34636 ; n34636_not
g59360 not n34645 ; n34645_not
g59361 not n34663 ; n34663_not
g59362 not n16267 ; n16267_not
g59363 not n34681 ; n34681_not
g59364 not n34708 ; n34708_not
g59365 not n26914 ; n26914_not
g59366 not n16285 ; n16285_not
g59367 not n47263 ; n47263_not
g59368 not n34735 ; n34735_not
g59369 not n34672 ; n34672_not
g59370 not n34744 ; n34744_not
g59371 not n26842 ; n26842_not
g59372 not n34609 ; n34609_not
g59373 not n26815 ; n26815_not
g59374 not n34843 ; n34843_not
g59375 not n34861 ; n34861_not
g59376 not n34870 ; n34870_not
g59377 not n26752 ; n26752_not
g59378 not n16348 ; n16348_not
g59379 not n26734 ; n26734_not
g59380 not n34933 ; n34933_not
g59381 not n15961 ; n15961_not
g59382 not n27265 ; n27265_not
g59383 not n15970 ; n15970_not
g59384 not n14962 ; n14962_not
g59385 not n44428 ; n44428_not
g59386 not n27229 ; n27229_not
g59387 not n24754 ; n24754_not
g59388 not n16069 ; n16069_not
g59389 not n34456 ; n34456_not
g59390 not n34474 ; n34474_not
g59391 not n27076 ; n27076_not
g59392 not n27157 ; n27157_not
g59393 not n34483 ; n34483_not
g59394 not n34492 ; n34492_not
g59395 not n10588 ; n10588_not
g59396 not n16096 ; n16096_not
g59397 not n47353 ; n47353_not
g59398 not n16159 ; n16159_not
g59399 not n16177 ; n16177_not
g59400 not n42178 ; n42178_not
g59401 not n34339 ; n34339_not
g59402 not n34528 ; n34528_not
g59403 not n34546 ; n34546_not
g59404 not n34537 ; n34537_not
g59405 not n16249 ; n16249_not
g59406 not n34573 ; n34573_not
g59407 not n16258 ; n16258_not
g59408 not n33259 ; n33259_not
g59409 not n42781 ; n42781_not
g59410 not n28624 ; n28624_not
g59411 not n33277 ; n33277_not
g59412 not n14935 ; n14935_not
g59413 not n14944 ; n14944_not
g59414 not n10687 ; n10687_not
g59415 not n42754 ; n42754_not
g59416 not n42745 ; n42745_not
g59417 not n42448 ; n42448_not
g59418 not n28570 ; n28570_not
g59419 not n42727 ; n42727_not
g59420 not n42718 ; n42718_not
g59421 not n10669 ; n10669_not
g59422 not n28534 ; n28534_not
g59423 not n33349 ; n33349_not
g59424 not n33376 ; n33376_not
g59425 not n47902 ; n47902_not
g59426 not n42691 ; n42691_not
g59427 not n47821 ; n47821_not
g59428 not n28435 ; n28435_not
g59429 not n42682 ; n42682_not
g59430 not n42673 ; n42673_not
g59431 not n28192 ; n28192_not
g59432 not n32926 ; n32926_not
g59433 not n32935 ; n32935_not
g59434 not n28930 ; n28930_not
g59435 not n32944 ; n32944_not
g59436 not n32953 ; n32953_not
g59437 not n28912 ; n28912_not
g59438 not n14665 ; n14665_not
g59439 not n14737 ; n14737_not
g59440 not n14485 ; n14485_not
g59441 not n33088 ; n33088_not
g59442 not n14755 ; n14755_not
g59443 not n14773 ; n14773_not
g59444 not n28804 ; n28804_not
g59445 not n42934 ; n42934_not
g59446 not n14791 ; n14791_not
g59447 not n42925 ; n42925_not
g59448 not n42916 ; n42916_not
g59449 not n14818 ; n14818_not
g59450 not n33187 ; n33187_not
g59451 not n33196 ; n33196_not
g59452 not n28732 ; n28732_not
g59453 not n14836 ; n14836_not
g59454 not n28705 ; n28705_not
g59455 not n42826 ; n42826_not
g59456 not n42817 ; n42817_not
g59457 not n42808 ; n42808_not
g59458 not n28642 ; n28642_not
g59459 not n33637 ; n33637_not
g59460 not n47542 ; n47542_not
g59461 not n28057 ; n28057_not
g59462 not n33655 ; n33655_not
g59463 not n42556 ; n42556_not
g59464 not n42547 ; n42547_not
g59465 not n15484 ; n15484_not
g59466 not n33709 ; n33709_not
g59467 not n33736 ; n33736_not
g59468 not n15538 ; n15538_not
g59469 not n33718 ; n33718_not
g59470 not n33745 ; n33745_not
g59471 not n27940 ; n27940_not
g59472 not n33763 ; n33763_not
g59473 not n27922 ; n27922_not
g59474 not n33808 ; n33808_not
g59475 not n15565 ; n15565_not
g59476 not n27913 ; n27913_not
g59477 not n33817 ; n33817_not
g59478 not n33835 ; n33835_not
g59479 not n33862 ; n33862_not
g59480 not n33691 ; n33691_not
g59481 not n33547 ; n33547_not
g59482 not n33943 ; n33943_not
g59483 not n15574 ; n15574_not
g59484 not n42655 ; n42655_not
g59485 not n15196 ; n15196_not
g59486 not n47722 ; n47722_not
g59487 not n47713 ; n47713_not
g59488 not n28183 ; n28183_not
g59489 not n28327 ; n28327_not
g59490 not n42646 ; n42646_not
g59491 not n15286 ; n15286_not
g59492 not n15295 ; n15295_not
g59493 not n42637 ; n42637_not
g59494 not n33529 ; n33529_not
g59495 not n33538 ; n33538_not
g59496 not n28255 ; n28255_not
g59497 not n28228 ; n28228_not
g59498 not n33565 ; n33565_not
g59499 not n33583 ; n33583_not
g59500 not n33592 ; n33592_not
g59501 not n15358 ; n15358_not
g59502 not n42880 ; n42880_not
g59503 not n28174 ; n28174_not
g59504 not n28165 ; n28165_not
g59505 not n28156 ; n28156_not
g59506 not n28147 ; n28147_not
g59507 not n15187 ; n15187_not
g59508 not n15457 ; n15457_not
g59509 not n44464 ; n44464_not
g59510 not n35284 ; n35284_not
g59511 not n47182 ; n47182_not
g59512 not n42088 ; n42088_not
g59513 not n41917 ; n41917_not
g59514 not n16807 ; n16807_not
g59515 not n26167 ; n26167_not
g59516 not n41746 ; n41746_not
g59517 not n16681 ; n16681_not
g59518 not n26338 ; n26338_not
g59519 not n42097 ; n42097_not
g59520 not n35563 ; n35563_not
g59521 not n35554 ; n35554_not
g59522 not n35095 ; n35095_not
g59523 not n41728 ; n41728_not
g59524 not n35473 ; n35473_not
g59525 not n16465 ; n16465_not
g59526 not n16906 ; n16906_not
g59527 not n17176 ; n17176_not
g59528 not n16447 ; n16447_not
g59529 not n16429 ; n16429_not
g59530 not n35059 ; n35059_not
g59531 not n25753 ; n25753_not
g59532 not n25825 ; n25825_not
g59533 not n16636 ; n16636_not
g59534 not n25816 ; n25816_not
g59535 not n35617 ; n35617_not
g59536 not n44473 ; n44473_not
g59537 not n25807 ; n25807_not
g59538 not n26437 ; n26437_not
g59539 not n16834 ; n16834_not
g59540 not n35176 ; n35176_not
g59541 not n10498 ; n10498_not
g59542 not n26365 ; n26365_not
g59543 not n17257 ; n17257_not
g59544 not n35446 ; n35446_not
g59545 not n41953 ; n41953_not
g59546 not n16555 ; n16555_not
g59547 not n26509 ; n26509_not
g59548 not n35635 ; n35635_not
g59549 not n25627 ; n25627_not
g59550 not n41908 ; n41908_not
g59551 not n16546 ; n16546_not
g59552 not n16528 ; n16528_not
g59553 not n16519 ; n16519_not
g59554 not n47218 ; n47218_not
g59555 not n25834 ; n25834_not
g59556 not n26545 ; n26545_not
g59557 not n17284 ; n17284_not
g59558 not n40198 ; n40198_not
g59559 not n41764 ; n41764_not
g59560 not n10399 ; n10399_not
g59561 not n41818 ; n41818_not
g59562 not n41773 ; n41773_not
g59563 not n25717 ; n25717_not
g59564 not n41782 ; n41782_not
g59565 not n25933 ; n25933_not
g59566 not n35257 ; n35257_not
g59567 not n26257 ; n26257_not
g59568 not n41791 ; n41791_not
g59569 not n26275 ; n26275_not
g59570 not n35266 ; n35266_not
g59571 not n44446 ; n44446_not
g59572 not n26068 ; n26068_not
g59573 not n35347 ; n35347_not
g59574 not n34951 ; n34951_not
g59575 not n25708 ; n25708_not
g59576 not n35743 ; n35743_not
g59577 not n35716 ; n35716_not
g59578 not n41737 ; n41737_not
g59579 not n35383 ; n35383_not
g59580 not n41962 ; n41962_not
g59581 not n26644 ; n26644_not
g59582 not n16726 ; n16726_not
g59583 not n26680 ; n26680_not
g59584 not n25870 ; n25870_not
g59585 not n37814 ; n37814_not
g59586 not n38912 ; n38912_not
g59587 not n35465 ; n35465_not
g59588 not n46184 ; n46184_not
g59589 not n41369 ; n41369_not
g59590 not n42647 ; n42647_not
g59591 not n48308 ; n48308_not
g59592 not n36059 ; n36059_not
g59593 not n38813 ; n38813_not
g59594 not n38741 ; n38741_not
g59595 not n36077 ; n36077_not
g59596 not n43754 ; n43754_not
g59597 not n34907 ; n34907_not
g59598 not n41387 ; n41387_not
g59599 not n33467 ; n33467_not
g59600 not n38804 ; n38804_not
g59601 not n46166 ; n46166_not
g59602 not n38903 ; n38903_not
g59603 not n33485 ; n33485_not
g59604 not n46193 ; n46193_not
g59605 not n38750 ; n38750_not
g59606 not n33494 ; n33494_not
g59607 not n38831 ; n38831_not
g59608 not n35456 ; n35456_not
g59609 not n43970 ; n43970_not
g59610 not n43097 ; n43097_not
g59611 not n41756 ; n41756_not
g59612 not n44573 ; n44573_not
g59613 not n33629 ; n33629_not
g59614 not n39128 ; n39128_not
g59615 not n39137 ; n39137_not
g59616 not n39146 ; n39146_not
g59617 not n43376 ; n43376_not
g59618 not n32684 ; n32684_not
g59619 not n33638 ; n33638_not
g59620 not n48623 ; n48623_not
g59621 not n37634 ; n37634_not
g59622 not n39173 ; n39173_not
g59623 not n35375 ; n35375_not
g59624 not n39191 ; n39191_not
g59625 not n40874 ; n40874_not
g59626 not n37625 ; n37625_not
g59627 not n39182 ; n39182_not
g59628 not n47570 ; n47570_not
g59629 not n39218 ; n39218_not
g59630 not n39236 ; n39236_not
g59631 not n33656 ; n33656_not
g59632 not n48164 ; n48164_not
g59633 not n41792 ; n41792_not
g59634 not n33692 ; n33692_not
g59635 not n39263 ; n39263_not
g59636 not n32657 ; n32657_not
g59637 not n34943 ; n34943_not
g59638 not n35339 ; n35339_not
g59639 not n45329 ; n45329_not
g59640 not n41585 ; n41585_not
g59641 not n38921 ; n38921_not
g59642 not n38930 ; n38930_not
g59643 not n35429 ; n35429_not
g59644 not n37715 ; n37715_not
g59645 not n43439 ; n43439_not
g59646 not n45266 ; n45266_not
g59647 not n42782 ; n42782_not
g59648 not n35447 ; n35447_not
g59649 not n32495 ; n32495_not
g59650 not n31469 ; n31469_not
g59651 not n46265 ; n46265_not
g59652 not n35294 ; n35294_not
g59653 not n32693 ; n32693_not
g59654 not n48650 ; n48650_not
g59655 not n35438 ; n35438_not
g59656 not n41747 ; n41747_not
g59657 not n39056 ; n39056_not
g59658 not n37652 ; n37652_not
g59659 not n47624 ; n47624_not
g59660 not n37643 ; n37643_not
g59661 not n39065 ; n39065_not
g59662 not n39029 ; n39029_not
g59663 not n46292 ; n46292_not
g59664 not n47615 ; n47615_not
g59665 not n39083 ; n39083_not
g59666 not n42962 ; n42962_not
g59667 not n45842 ; n45842_not
g59668 not n42944 ; n42944_not
g59669 not n35870 ; n35870_not
g59670 not n49037 ; n49037_not
g59671 not n42935 ; n42935_not
g59672 not n35906 ; n35906_not
g59673 not n40676 ; n40676_not
g59674 not n35915 ; n35915_not
g59675 not n38174 ; n38174_not
g59676 not n35933 ; n35933_not
g59677 not n38309 ; n38309_not
g59678 not n16493 ; n16493_not
g59679 not n33197 ; n33197_not
g59680 not n35942 ; n35942_not
g59681 not n38147 ; n38147_not
g59682 not n35690 ; n35690_not
g59683 not n42836 ; n42836_not
g59684 not n42827 ; n42827_not
g59685 not n45455 ; n45455_not
g59686 not n35681 ; n35681_not
g59687 not n45905 ; n45905_not
g59688 not n42818 ; n42818_not
g59689 not n31892 ; n31892_not
g59690 not n16853 ; n16853_not
g59691 not n35762 ; n35762_not
g59692 not n32945 ; n32945_not
g59693 not n38237 ; n38237_not
g59694 not n31946 ; n31946_not
g59695 not n32756 ; n32756_not
g59696 not n32954 ; n32954_not
g59697 not n44177 ; n44177_not
g59698 not n35726 ; n35726_not
g59699 not n32882 ; n32882_not
g59700 not n35843 ; n35843_not
g59701 not n32963 ; n32963_not
g59702 not n32972 ; n32972_not
g59703 not n45707 ; n45707_not
g59704 not n32990 ; n32990_not
g59705 not n32855 ; n32855_not
g59706 not n45680 ; n45680_not
g59707 not n38228 ; n38228_not
g59708 not n38255 ; n38255_not
g59709 not n31919 ; n31919_not
g59710 not n48047 ; n48047_not
g59711 not n47183 ; n47183_not
g59712 not n31928 ; n31928_not
g59713 not n35852 ; n35852_not
g59714 not n45833 ; n45833_not
g59715 not n38273 ; n38273_not
g59716 not n33098 ; n33098_not
g59717 not n32846 ; n32846_not
g59718 not n35717 ; n35717_not
g59719 not n38282 ; n38282_not
g59720 not n48038 ; n48038_not
g59721 not n42467 ; n42467_not
g59722 not n42692 ; n42692_not
g59723 not n41675 ; n41675_not
g59724 not n48281 ; n48281_not
g59725 not n37913 ; n37913_not
g59726 not n38552 ; n38552_not
g59727 not n38543 ; n38543_not
g59728 not n33395 ; n33395_not
g59729 not n47813 ; n47813_not
g59730 not n47129 ; n47129_not
g59731 not n38606 ; n38606_not
g59732 not n42674 ; n42674_not
g59733 not n38615 ; n38615_not
g59734 not n47723 ; n47723_not
g59735 not n43385 ; n43385_not
g59736 not n46148 ; n46148_not
g59737 not n37832 ; n37832_not
g59738 not n38633 ; n38633_not
g59739 not n38705 ; n38705_not
g59740 not n32738 ; n32738_not
g59741 not n38723 ; n38723_not
g59742 not n38732 ; n38732_not
g59743 not n48227 ; n48227_not
g59744 not n45923 ; n45923_not
g59745 not n41693 ; n41693_not
g59746 not n42791 ; n42791_not
g59747 not n35672 ; n35672_not
g59748 not n35663 ; n35663_not
g59749 not n35645 ; n35645_not
g59750 not n31856 ; n31856_not
g59751 not n35960 ; n35960_not
g59752 not n32819 ; n32819_not
g59753 not n33278 ; n33278_not
g59754 not n31847 ; n31847_not
g59755 not n38354 ; n38354_not
g59756 not n38084 ; n38084_not
g59757 not n38372 ; n38372_not
g59758 not n38075 ; n38075_not
g59759 not n38390 ; n38390_not
g59760 not n32792 ; n32792_not
g59761 not n35609 ; n35609_not
g59762 not n38444 ; n38444_not
g59763 not n32774 ; n32774_not
g59764 not n44069 ; n44069_not
g59765 not n48263 ; n48263_not
g59766 not n47903 ; n47903_not
g59767 not n38462 ; n38462_not
g59768 not n35591 ; n35591_not
g59769 not n38471 ; n38471_not
g59770 not n38480 ; n38480_not
g59771 not n35186 ; n35186_not
g59772 not n37166 ; n37166_not
g59773 not n35168 ; n35168_not
g59774 not n41918 ; n41918_not
g59775 not n40739 ; n40739_not
g59776 not n35159 ; n35159_not
g59777 not n36608 ; n36608_not
g59778 not n40469 ; n40469_not
g59779 not n37094 ; n37094_not
g59780 not n36617 ; n36617_not
g59781 not n42188 ; n42188_not
g59782 not n43709 ; n43709_not
g59783 not n44438 ; n44438_not
g59784 not n32396 ; n32396_not
g59785 not n43682 ; n43682_not
g59786 not n42179 ; n42179_not
g59787 not n48461 ; n48461_not
g59788 not n43673 ; n43673_not
g59789 not n43655 ; n43655_not
g59790 not n43187 ; n43187_not
g59791 not n40568 ; n40568_not
g59792 not n43646 ; n43646_not
g59793 not n34529 ; n34529_not
g59794 not n43619 ; n43619_not
g59795 not n36653 ; n36653_not
g59796 not n32378 ; n32378_not
g59797 not n43538 ; n43538_not
g59798 not n34556 ; n34556_not
g59799 not n40595 ; n40595_not
g59800 not n47345 ; n47345_not
g59801 not n36491 ; n36491_not
g59802 not n44483 ; n44483_not
g59803 not n37265 ; n37265_not
g59804 not n37256 ; n37256_not
g59805 not n44456 ; n44456_not
g59806 not n41954 ; n41954_not
g59807 not n36482 ; n36482_not
g59808 not n34286 ; n34286_not
g59809 not n47219 ; n47219_not
g59810 not n34295 ; n34295_not
g59811 not n47381 ; n47381_not
g59812 not n43736 ; n43736_not
g59813 not n42287 ; n42287_not
g59814 not n43484 ; n43484_not
g59815 not n46517 ; n46517_not
g59816 not n39074 ; n39074_not
g59817 not n37229 ; n37229_not
g59818 not n34349 ; n34349_not
g59819 not n36536 ; n36536_not
g59820 not n32459 ; n32459_not
g59821 not n42269 ; n42269_not
g59822 not n41882 ; n41882_not
g59823 not n44474 ; n44474_not
g59824 not n36554 ; n36554_not
g59825 not n31667 ; n31667_not
g59826 not n40397 ; n40397_not
g59827 not n41873 ; n41873_not
g59828 not n37193 ; n37193_not
g59829 not n46823 ; n46823_not
g59830 not n40757 ; n40757_not
g59831 not n36842 ; n36842_not
g59832 not n43583 ; n43583_not
g59833 not n43259 ; n43259_not
g59834 not n40766 ; n40766_not
g59835 not n47237 ; n47237_not
g59836 not n47228 ; n47228_not
g59837 not n40775 ; n40775_not
g59838 not n34835 ; n34835_not
g59839 not n36824 ; n36824_not
g59840 not n43556 ; n43556_not
g59841 not n48542 ; n48542_not
g59842 not n46715 ; n46715_not
g59843 not n36707 ; n36707_not
g59844 not n40793 ; n40793_not
g59845 not n36815 ; n36815_not
g59846 not n44627 ; n44627_not
g59847 not n46526 ; n46526_not
g59848 not n40856 ; n40856_not
g59849 not n36770 ; n36770_not
g59850 not n36761 ; n36761_not
g59851 not n40937 ; n40937_not
g59852 not n34961 ; n34961_not
g59853 not n36266 ; n36266_not
g59854 not n40892 ; n40892_not
g59855 not n36725 ; n36725_not
g59856 not n40199 ; n40199_not
g59857 not n37067 ; n37067_not
g59858 not n46931 ; n46931_not
g59859 not n35078 ; n35078_not
g59860 not n34664 ; n34664_not
g59861 not n42548 ; n42548_not
g59862 not n35069 ; n35069_not
g59863 not n40667 ; n40667_not
g59864 not n44618 ; n44618_not
g59865 not n32369 ; n32369_not
g59866 not n34709 ; n34709_not
g59867 not n34727 ; n34727_not
g59868 not n40982 ; n40982_not
g59869 not n48506 ; n48506_not
g59870 not n36950 ; n36950_not
g59871 not n46625 ; n46625_not
g59872 not n34772 ; n34772_not
g59873 not n36923 ; n36923_not
g59874 not n36914 ; n36914_not
g59875 not n46634 ; n46634_not
g59876 not n34817 ; n34817_not
g59877 not n40964 ; n40964_not
g59878 not n46553 ; n46553_not
g59879 not n47255 ; n47255_not
g59880 not n46661 ; n46661_not
g59881 not n40748 ; n40748_not
g59882 not n43907 ; n43907_not
g59883 not n37490 ; n37490_not
g59884 not n33890 ; n33890_not
g59885 not n41864 ; n41864_not
g59886 not n36257 ; n36257_not
g59887 not n33944 ; n33944_not
g59888 not n39506 ; n39506_not
g59889 not n37445 ; n37445_not
g59890 not n37436 ; n37436_not
g59891 not n31991 ; n31991_not
g59892 not n36275 ; n36275_not
g59893 not n33953 ; n33953_not
g59894 not n33971 ; n33971_not
g59895 not n41819 ; n41819_not
g59896 not n44276 ; n44276_not
g59897 not n47075 ; n47075_not
g59898 not n39560 ; n39560_not
g59899 not n43844 ; n43844_not
g59900 not n42485 ; n42485_not
g59901 not n47435 ; n47435_not
g59902 not n32594 ; n32594_not
g59903 not n39605 ; n39605_not
g59904 not n47057 ; n47057_not
g59905 not n37391 ; n37391_not
g59906 not n37382 ; n37382_not
g59907 not n48353 ; n48353_not
g59908 not n33746 ; n33746_not
g59909 not n32648 ; n32648_not
g59910 not n33755 ; n33755_not
g59911 not n39326 ; n39326_not
g59912 not n33764 ; n33764_not
g59913 not n32639 ; n32639_not
g59914 not n39371 ; n39371_not
g59915 not n39380 ; n39380_not
g59916 not n36185 ; n36185_not
g59917 not n37571 ; n37571_not
g59918 not n36194 ; n36194_not
g59919 not n41279 ; n41279_not
g59920 not n37553 ; n37553_not
g59921 not n37544 ; n37544_not
g59922 not n33809 ; n33809_not
g59923 not n31784 ; n31784_not
g59924 not n41855 ; n41855_not
g59925 not n33845 ; n33845_not
g59926 not n48371 ; n48371_not
g59927 not n46382 ; n46382_not
g59928 not n33863 ; n33863_not
g59929 not n47525 ; n47525_not
g59930 not n31559 ; n31559_not
g59931 not n33872 ; n33872_not
g59932 not n46391 ; n46391_not
g59933 not n33881 ; n33881_not
g59934 not n43763 ; n43763_not
g59935 not n41963 ; n41963_not
g59936 not n41198 ; n41198_not
g59937 not n39902 ; n39902_not
g59938 not n39911 ; n39911_not
g59939 not n39920 ; n39920_not
g59940 not n32198 ; n32198_not
g59941 not n38651 ; n38651_not
g59942 not n36437 ; n36437_not
g59943 not n46481 ; n46481_not
g59944 not n48407 ; n48407_not
g59945 not n34169 ; n34169_not
g59946 not n39713 ; n39713_not
g59947 not n34187 ; n34187_not
g59948 not n31649 ; n31649_not
g59949 not n36455 ; n36455_not
g59950 not n37292 ; n37292_not
g59951 not n44753 ; n44753_not
g59952 not n42395 ; n42395_not
g59953 not n44726 ; n44726_not
g59954 not n43808 ; n43808_not
g59955 not n37283 ; n37283_not
g59956 not n38570 ; n38570_not
g59957 not n47039 ; n47039_not
g59958 not n35258 ; n35258_not
g59959 not n42368 ; n42368_not
g59960 not n36464 ; n36464_not
g59961 not n35249 ; n35249_not
g59962 not n48434 ; n48434_not
g59963 not n37274 ; n37274_not
g59964 not n47408 ; n47408_not
g59965 not n34259 ; n34259_not
g59966 not n43835 ; n43835_not
g59967 not n35285 ; n35285_not
g59968 not n32189 ; n32189_not
g59969 not n34079 ; n34079_not
g59970 not n37346 ; n37346_not
g59971 not n39623 ; n39623_not
g59972 not n39632 ; n39632_not
g59973 not n46328 ; n46328_not
g59974 not n37337 ; n37337_not
g59975 not n36356 ; n36356_not
g59976 not n39641 ; n39641_not
g59977 not n38561 ; n38561_not
g59978 not n34097 ; n34097_not
g59979 not n46436 ; n46436_not
g59980 not n36365 ; n36365_not
g59981 not n32558 ; n32558_not
g59982 not n36383 ; n36383_not
g59983 not n41945 ; n41945_not
g59984 not n46445 ; n46445_not
g59985 not n46454 ; n46454_not
g59986 not n41189 ; n41189_not
g59987 not n43826 ; n43826_not
g59988 not n42449 ; n42449_not
g59989 not n39812 ; n39812_not
g59990 not n47417 ; n47417_not
g59991 not n43817 ; n43817_not
g59992 not n28823 ; n28823_not
g59993 not n28814 ; n28814_not
g59994 not n18185 ; n18185_not
g59995 not n18095 ; n18095_not
g59996 not n18167 ; n18167_not
g59997 not n18248 ; n18248_not
g59998 not n18257 ; n18257_not
g59999 not n18266 ; n18266_not
g60000 not n18275 ; n18275_not
g60001 not n18329 ; n18329_not
g60002 not n18392 ; n18392_not
g60003 not n18383 ; n18383_not
g60004 not n18419 ; n18419_not
g60005 not n18428 ; n18428_not
g60006 not n18455 ; n18455_not
g60007 not n28733 ; n28733_not
g60008 not n18554 ; n18554_not
g60009 not n18563 ; n18563_not
g60010 not n18581 ; n18581_not
g60011 not n28670 ; n28670_not
g60012 not n16970 ; n16970_not
g60013 not n28652 ; n28652_not
g60014 not n18617 ; n18617_not
g60015 not n18626 ; n18626_not
g60016 not n28634 ; n28634_not
g60017 not n18662 ; n18662_not
g60018 not n28607 ; n28607_not
g60019 not n17348 ; n17348_not
g60020 not n17366 ; n17366_not
g60021 not n17375 ; n17375_not
g60022 not n17456 ; n17456_not
g60023 not n17168 ; n17168_not
g60024 not n28904 ; n28904_not
g60025 not n17519 ; n17519_not
g60026 not n17528 ; n17528_not
g60027 not n17537 ; n17537_not
g60028 not n16727 ; n16727_not
g60029 not n17609 ; n17609_not
g60030 not n17645 ; n17645_not
g60031 not n17663 ; n17663_not
g60032 not n17672 ; n17672_not
g60033 not n17708 ; n17708_not
g60034 not n17726 ; n17726_not
g60035 not n17735 ; n17735_not
g60036 not n17762 ; n17762_not
g60037 not n17096 ; n17096_not
g60038 not n28751 ; n28751_not
g60039 not n17771 ; n17771_not
g60040 not n17825 ; n17825_not
g60041 not n28850 ; n28850_not
g60042 not n17924 ; n17924_not
g60043 not n28841 ; n28841_not
g60044 not n28832 ; n28832_not
g60045 not n17906 ; n17906_not
g60046 not n28418 ; n28418_not
g60047 not n19148 ; n19148_not
g60048 not n28274 ; n28274_not
g60049 not n19238 ; n19238_not
g60050 not n19247 ; n19247_not
g60051 not n19256 ; n19256_not
g60052 not n19265 ; n19265_not
g60053 not n19193 ; n19193_not
g60054 not n19283 ; n19283_not
g60055 not n28373 ; n28373_not
g60056 not n19346 ; n19346_not
g60057 not n28364 ; n28364_not
g60058 not n19373 ; n19373_not
g60059 not n28355 ; n28355_not
g60060 not n19391 ; n19391_not
g60061 not n28346 ; n28346_not
g60062 not n28337 ; n28337_not
g60063 not n19418 ; n19418_not
g60064 not n17546 ; n17546_not
g60065 not n19490 ; n19490_not
g60066 not n19481 ; n19481_not
g60067 not n19544 ; n19544_not
g60068 not n19562 ; n19562_not
g60069 not n19625 ; n19625_not
g60070 not n28256 ; n28256_not
g60071 not n19634 ; n19634_not
g60072 not n19643 ; n19643_not
g60073 not n19652 ; n19652_not
g60074 not n19670 ; n19670_not
g60075 not n18680 ; n18680_not
g60076 not n18752 ; n18752_not
g60077 not n28580 ; n28580_not
g60078 not n18806 ; n18806_not
g60079 not n28562 ; n28562_not
g60080 not n28481 ; n28481_not
g60081 not n18743 ; n18743_not
g60082 not n28553 ; n28553_not
g60083 not n28544 ; n28544_not
g60084 not n28535 ; n28535_not
g60085 not n28454 ; n28454_not
g60086 not n28517 ; n28517_not
g60087 not n28508 ; n28508_not
g60088 not n18905 ; n18905_not
g60089 not n28490 ; n28490_not
g60090 not n18833 ; n18833_not
g60091 not n19058 ; n19058_not
g60092 not n19067 ; n19067_not
g60093 not n19076 ; n19076_not
g60094 not n19085 ; n19085_not
g60095 not n19139 ; n19139_not
g60096 not n19175 ; n19175_not
g60097 not n28427 ; n28427_not
g60098 not n28409 ; n28409_not
g60099 not n15395 ; n15395_not
g60100 not n29435 ; n29435_not
g60101 not n15386 ; n15386_not
g60102 not n15476 ; n15476_not
g60103 not n15494 ; n15494_not
g60104 not n15377 ; n15377_not
g60105 not n29390 ; n29390_not
g60106 not n15584 ; n15584_not
g60107 not n15593 ; n15593_not
g60108 not n29381 ; n29381_not
g60109 not n13685 ; n13685_not
g60110 not n15629 ; n15629_not
g60111 not n15638 ; n15638_not
g60112 not n15647 ; n15647_not
g60113 not n15674 ; n15674_not
g60114 not n29354 ; n29354_not
g60115 not n15719 ; n15719_not
g60116 not n15728 ; n15728_not
g60117 not n15764 ; n15764_not
g60118 not n29336 ; n29336_not
g60119 not n14657 ; n14657_not
g60120 not n15773 ; n15773_not
g60121 not n14666 ; n14666_not
g60122 not n15809 ; n15809_not
g60123 not n15827 ; n15827_not
g60124 not n15836 ; n15836_not
g60125 not n15872 ; n15872_not
g60126 not n15908 ; n15908_not
g60127 not n29255 ; n29255_not
g60128 not n14486 ; n14486_not
g60129 not n11669 ; n11669_not
g60130 not n14639 ; n14639_not
g60131 not n14459 ; n14459_not
g60132 not n14693 ; n14693_not
g60133 not n14648 ; n14648_not
g60134 not n14765 ; n14765_not
g60135 not n14774 ; n14774_not
g60136 not n14792 ; n14792_not
g60137 not n14828 ; n14828_not
g60138 not n14738 ; n14738_not
g60139 not n10976 ; n10976_not
g60140 not n29543 ; n29543_not
g60141 not n14882 ; n14882_not
g60142 not n29534 ; n29534_not
g60143 not n29480 ; n29480_not
g60144 not n29525 ; n29525_not
g60145 not n14927 ; n14927_not
g60146 not n14963 ; n14963_not
g60147 not n14972 ; n14972_not
g60148 not n14990 ; n14990_not
g60149 not n14936 ; n14936_not
g60150 not n15188 ; n15188_not
g60151 not n15368 ; n15368_not
g60152 not n16466 ; n16466_not
g60153 not n29129 ; n29129_not
g60154 not n16583 ; n16583_not
g60155 not n29093 ; n29093_not
g60156 not n16619 ; n16619_not
g60157 not n16637 ; n16637_not
g60158 not n16646 ; n16646_not
g60159 not n16673 ; n16673_not
g60160 not n16691 ; n16691_not
g60161 not n29075 ; n29075_not
g60162 not n16718 ; n16718_not
g60163 not n16736 ; n16736_not
g60164 not n16781 ; n16781_not
g60165 not n29039 ; n29039_not
g60166 not n16835 ; n16835_not
g60167 not n16844 ; n16844_not
g60168 not n16862 ; n16862_not
g60169 not n16916 ; n16916_not
g60170 not n17069 ; n17069_not
g60171 not n17087 ; n17087_not
g60172 not n17159 ; n17159_not
g60173 not n17267 ; n17267_not
g60174 not n17294 ; n17294_not
g60175 not n15881 ; n15881_not
g60176 not n29219 ; n29219_not
g60177 not n15917 ; n15917_not
g60178 not n15935 ; n15935_not
g60179 not n29246 ; n29246_not
g60180 not n14585 ; n14585_not
g60181 not n29237 ; n29237_not
g60182 not n15944 ; n15944_not
g60183 not n15962 ; n15962_not
g60184 not n15971 ; n15971_not
g60185 not n15980 ; n15980_not
g60186 not n16079 ; n16079_not
g60187 not n16097 ; n16097_not
g60188 not n16169 ; n16169_not
g60189 not n16196 ; n16196_not
g60190 not n16277 ; n16277_not
g60191 not n16349 ; n16349_not
g60192 not n15845 ; n15845_not
g60193 not n16367 ; n16367_not
g60194 not n16385 ; n16385_not
g60195 not n15746 ; n15746_not
g60196 not n29147 ; n29147_not
g60197 not n16439 ; n16439_not
g60198 not n29138 ; n29138_not
g60199 not n16448 ; n16448_not
g60200 not n24566 ; n24566_not
g60201 not n24575 ; n24575_not
g60202 not n26960 ; n26960_not
g60203 not n24593 ; n24593_not
g60204 not n26951 ; n26951_not
g60205 not n24629 ; n24629_not
g60206 not n24656 ; n24656_not
g60207 not n26942 ; n26942_not
g60208 not n26933 ; n26933_not
g60209 not n24692 ; n24692_not
g60210 not n24719 ; n24719_not
g60211 not n24737 ; n24737_not
g60212 not n26924 ; n26924_not
g60213 not n24773 ; n24773_not
g60214 not n24782 ; n24782_not
g60215 not n24818 ; n24818_not
g60216 not n24674 ; n24674_not
g60217 not n24836 ; n24836_not
g60218 not n24845 ; n24845_not
g60219 not n24854 ; n24854_not
g60220 not n24863 ; n24863_not
g60221 not n24872 ; n24872_not
g60222 not n24881 ; n24881_not
g60223 not n24917 ; n24917_not
g60224 not n24935 ; n24935_not
g60225 not n26843 ; n26843_not
g60226 not n24980 ; n24980_not
g60227 not n26780 ; n26780_not
g60228 not n23792 ; n23792_not
g60229 not n23819 ; n23819_not
g60230 not n27185 ; n27185_not
g60231 not n23846 ; n23846_not
g60232 not n27194 ; n27194_not
g60233 not n23873 ; n23873_not
g60234 not n23882 ; n23882_not
g60235 not n23918 ; n23918_not
g60236 not n23945 ; n23945_not
g60237 not n27167 ; n27167_not
g60238 not n23963 ; n23963_not
g60239 not n27149 ; n27149_not
g60240 not n23972 ; n23972_not
g60241 not n27068 ; n27068_not
g60242 not n27095 ; n27095_not
g60243 not n27086 ; n27086_not
g60244 not n27077 ; n27077_not
g60245 not n24098 ; n24098_not
g60246 not n24179 ; n24179_not
g60247 not n24197 ; n24197_not
g60248 not n24278 ; n24278_not
g60249 not n24287 ; n24287_not
g60250 not n24296 ; n24296_not
g60251 not n26861 ; n26861_not
g60252 not n24359 ; n24359_not
g60253 not n24377 ; n24377_not
g60254 not n24467 ; n24467_not
g60255 not n24539 ; n24539_not
g60256 not n24548 ; n24548_not
g60257 not n26618 ; n26618_not
g60258 not n26609 ; n26609_not
g60259 not n25835 ; n25835_not
g60260 not n25844 ; n25844_not
g60261 not n25853 ; n25853_not
g60262 not n25655 ; n25655_not
g60263 not n25871 ; n25871_not
g60264 not n25880 ; n25880_not
g60265 not n25934 ; n25934_not
g60266 not n25943 ; n25943_not
g60267 not n25952 ; n25952_not
g60268 not n26537 ; n26537_not
g60269 not n25961 ; n25961_not
g60270 not n26519 ; n26519_not
g60271 not n26528 ; n26528_not
g60272 not n26384 ; n26384_not
g60273 not n26087 ; n26087_not
g60274 not n26168 ; n26168_not
g60275 not n26177 ; n26177_not
g60276 not n26186 ; n26186_not
g60277 not n26483 ; n26483_not
g60278 not n26195 ; n26195_not
g60279 not n26474 ; n26474_not
g60280 not n26267 ; n26267_not
g60281 not n26465 ; n26465_not
g60282 not n26285 ; n26285_not
g60283 not n26366 ; n26366_not
g60284 not n26456 ; n26456_not
g60285 not n26447 ; n26447_not
g60286 not n25169 ; n25169_not
g60287 not n26762 ; n26762_not
g60288 not n25358 ; n25358_not
g60289 not n25475 ; n25475_not
g60290 not n25493 ; n25493_not
g60291 not n26744 ; n26744_not
g60292 not n26708 ; n26708_not
g60293 not n25556 ; n25556_not
g60294 not n26717 ; n26717_not
g60295 not n25367 ; n25367_not
g60296 not n25583 ; n25583_not
g60297 not n26690 ; n26690_not
g60298 not n25637 ; n25637_not
g60299 not n25664 ; n25664_not
g60300 not n25673 ; n25673_not
g60301 not n25682 ; n25682_not
g60302 not n25691 ; n25691_not
g60303 not n25727 ; n25727_not
g60304 not n25736 ; n25736_not
g60305 not n25763 ; n25763_not
g60306 not n26672 ; n26672_not
g60307 not n26591 ; n26591_not
g60308 not n25781 ; n25781_not
g60309 not n26663 ; n26663_not
g60310 not n26654 ; n26654_not
g60311 not n25826 ; n25826_not
g60312 not n26645 ; n26645_not
g60313 not n26564 ; n26564_not
g60314 not n26627 ; n26627_not
g60315 not n20849 ; n20849_not
g60316 not n27860 ; n27860_not
g60317 not n20885 ; n20885_not
g60318 not n20894 ; n20894_not
g60319 not n20984 ; n20984_not
g60320 not n21398 ; n21398_not
g60321 not n27833 ; n27833_not
g60322 not n21479 ; n21479_not
g60323 not n21578 ; n21578_not
g60324 not n27824 ; n27824_not
g60325 not n27752 ; n27752_not
g60326 not n21587 ; n21587_not
g60327 not n21686 ; n21686_not
g60328 not n21695 ; n21695_not
g60329 not n21794 ; n21794_not
g60330 not n27815 ; n27815_not
g60331 not n21857 ; n21857_not
g60332 not n21884 ; n21884_not
g60333 not n21947 ; n21947_not
g60334 not n21965 ; n21965_not
g60335 not n21956 ; n21956_not
g60336 not n21992 ; n21992_not
g60337 not n22199 ; n22199_not
g60338 not n22289 ; n22289_not
g60339 not n22298 ; n22298_not
g60340 not n22388 ; n22388_not
g60341 not n28184 ; n28184_not
g60342 not n19724 ; n19724_not
g60343 not n28157 ; n28157_not
g60344 not n19742 ; n19742_not
g60345 not n28139 ; n28139_not
g60346 not n28094 ; n28094_not
g60347 not n19760 ; n19760_not
g60348 not n28085 ; n28085_not
g60349 not n19715 ; n19715_not
g60350 not n28076 ; n28076_not
g60351 not n28067 ; n28067_not
g60352 not n28049 ; n28049_not
g60353 not n19805 ; n19805_not
g60354 not n19814 ; n19814_not
g60355 not n19832 ; n19832_not
g60356 not n19850 ; n19850_not
g60357 not n19904 ; n19904_not
g60358 not n19913 ; n19913_not
g60359 not n19931 ; n19931_not
g60360 not n27806 ; n27806_not
g60361 not n27941 ; n27941_not
g60362 not n27932 ; n27932_not
g60363 not n27905 ; n27905_not
g60364 not n20669 ; n20669_not
g60365 not n20687 ; n20687_not
g60366 not n20696 ; n20696_not
g60367 not n20759 ; n20759_not
g60368 not n20786 ; n20786_not
g60369 not n20858 ; n20858_not
g60370 not n22775 ; n22775_not
g60371 not n27491 ; n27491_not
g60372 not n22982 ; n22982_not
g60373 not n27473 ; n27473_not
g60374 not n22784 ; n22784_not
g60375 not n22991 ; n22991_not
g60376 not n27455 ; n27455_not
g60377 not n27428 ; n27428_not
g60378 not n27419 ; n27419_not
g60379 not n27392 ; n27392_not
g60380 not n23288 ; n23288_not
g60381 not n27383 ; n27383_not
g60382 not n23369 ; n23369_not
g60383 not n23378 ; n23378_not
g60384 not n23459 ; n23459_not
g60385 not n27365 ; n27365_not
g60386 not n23477 ; n23477_not
g60387 not n23549 ; n23549_not
g60388 not n23558 ; n23558_not
g60389 not n27329 ; n27329_not
g60390 not n23576 ; n23576_not
g60391 not n23639 ; n23639_not
g60392 not n23657 ; n23657_not
g60393 not n27284 ; n27284_not
g60394 not n23675 ; n23675_not
g60395 not n23738 ; n23738_not
g60396 not n27257 ; n27257_not
g60397 not n23783 ; n23783_not
g60398 not n27239 ; n27239_not
g60399 not n22379 ; n22379_not
g60400 not n27680 ; n27680_not
g60401 not n22397 ; n22397_not
g60402 not n22469 ; n22469_not
g60403 not n22478 ; n22478_not
g60404 not n27662 ; n27662_not
g60405 not n22487 ; n22487_not
g60406 not n22496 ; n22496_not
g60407 not n22559 ; n22559_not
g60408 not n22586 ; n22586_not
g60409 not n27617 ; n27617_not
g60410 not n22649 ; n22649_not
g60411 not n27608 ; n27608_not
g60412 not n22667 ; n22667_not
g60413 not n22685 ; n22685_not
g60414 not n27509 ; n27509_not
g60415 not n22748 ; n22748_not
g60416 not n22757 ; n22757_not
g60417 not n27581 ; n27581_not
g60418 not n22766 ; n22766_not
g60419 not n27563 ; n27563_not
g60420 not n22847 ; n22847_not
g60421 not n27536 ; n27536_not
g60422 not n27527 ; n27527_not
g60423 not n27518 ; n27518_not
g60424 not n29804 ; n29804_not
g60425 not n13946 ; n13946_not
g60426 not n29930 ; n29930_not
g60427 not n29750 ; n29750_not
g60428 not n14297 ; n14297_not
g60429 not n14378 ; n14378_not
g60430 not n11678 ; n11678_not
g60431 not n13559 ; n13559_not
g60432 not n11795 ; n11795_not
g60433 not n14387 ; n14387_not
g60434 not n30938 ; n30938_not
g60435 not n30389 ; n30389_not
g60436 not n11975 ; n11975_not
g60437 not n11984 ; n11984_not
g60438 not n12848 ; n12848_not
g60439 not n14396 ; n14396_not
g60440 not n11687 ; n11687_not
g60441 not n30992 ; n30992_not
g60442 not n12389 ; n12389_not
g60443 not n12596 ; n12596_not
g60444 not n29903 ; n29903_not
g60445 not n14279 ; n14279_not
g60446 not n29831 ; n29831_not
g60447 not n14288 ; n14288_not
g60448 not n30686 ; n30686_not
g60449 not n11777 ; n11777_not
g60450 not n11885 ; n11885_not
g60451 not n29822 ; n29822_not
g60452 not n13937 ; n13937_not
g60453 not n30947 ; n30947_not
g60454 not n13388 ; n13388_not
g60455 not n13892 ; n13892_not
g60456 not n14099 ; n14099_not
g60457 not n11876 ; n11876_not
g60458 not n30695 ; n30695_not
g60459 not n10877 ; n10877_not
g60460 not n12776 ; n12776_not
g60461 not n11858 ; n11858_not
g60462 not n12974 ; n12974_not
g60463 not n13784 ; n13784_not
g60464 not n30893 ; n30893_not
g60465 not n30965 ; n30965_not
g60466 not n13694 ; n13694_not
g60467 not n10895 ; n10895_not
g60468 not n13964 ; n13964_not
g60469 not n31379 ; n31379_not
g60470 not n29660 ; n29660_not
g60471 not n13199 ; n13199_not
g60472 not n14549 ; n14549_not
g60473 not n30974 ; n30974_not
g60474 not n13982 ; n13982_not
g60475 not n10868 ; n10868_not
g60476 not n13577 ; n13577_not
g60477 not n13586 ; n13586_not
g60478 not n13955 ; n13955_not
g60479 not n11489 ; n11489_not
g60480 not n12938 ; n12938_not
g60481 not n13766 ; n13766_not
g60482 not n12758 ; n12758_not
g60483 not n10697 ; n10697_not
g60484 not n13838 ; n13838_not
g60485 not n30758 ; n30758_not
g60486 not n45159 ; n45159_not
g60487 not n21399 ; n21399_not
g60488 not n45258 ; n45258_not
g60489 not n43791 ; n43791_not
g60490 not n27825 ; n27825_not
g60491 not n21579 ; n21579_not
g60492 not n38247 ; n38247_not
g60493 not n33954 ; n33954_not
g60494 not n33963 ; n33963_not
g60495 not n21489 ; n21489_not
g60496 not n27870 ; n27870_not
g60497 not n31767 ; n31767_not
g60498 not n44664 ; n44664_not
g60499 not n33756 ; n33756_not
g60500 not n17862 ; n17862_not
g60501 not n38409 ; n38409_not
g60502 not n20787 ; n20787_not
g60503 not n38436 ; n38436_not
g60504 not n20778 ; n20778_not
g60505 not n38454 ; n38454_not
g60506 not n38553 ; n38553_not
g60507 not n38562 ; n38562_not
g60508 not n38580 ; n38580_not
g60509 not n20976 ; n20976_not
g60510 not n27843 ; n27843_not
g60511 not n33936 ; n33936_not
g60512 not n20949 ; n20949_not
g60513 not n20895 ; n20895_not
g60514 not n27852 ; n27852_not
g60515 not n38346 ; n38346_not
g60516 not n33927 ; n33927_not
g60517 not n27861 ; n27861_not
g60518 not n38355 ; n38355_not
g60519 not n33918 ; n33918_not
g60520 not n20877 ; n20877_not
g60521 not n38364 ; n38364_not
g60522 not n20868 ; n20868_not
g60523 not n33909 ; n33909_not
g60524 not n22488 ; n22488_not
g60525 not n27663 ; n27663_not
g60526 not n37635 ; n37635_not
g60527 not n27672 ; n27672_not
g60528 not n37680 ; n37680_not
g60529 not n45654 ; n45654_not
g60530 not n22389 ; n22389_not
g60531 not n37707 ; n37707_not
g60532 not n30399 ; n30399_not
g60533 not n37716 ; n37716_not
g60534 not n31596 ; n31596_not
g60535 not n45645 ; n45645_not
g60536 not n37743 ; n37743_not
g60537 not n27690 ; n27690_not
g60538 not n37752 ; n37752_not
g60539 not n34791 ; n34791_not
g60540 not n22299 ; n22299_not
g60541 not n37518 ; n37518_not
g60542 not n27573 ; n27573_not
g60543 not n22776 ; n22776_not
g60544 not n34188 ; n34188_not
g60545 not n37536 ; n37536_not
g60546 not n27582 ; n27582_not
g60547 not n37581 ; n37581_not
g60548 not n37590 ; n37590_not
g60549 not n17187 ; n17187_not
g60550 not n27609 ; n27609_not
g60551 not n22659 ; n22659_not
g60552 not n45735 ; n45735_not
g60553 not n22578 ; n22578_not
g60554 not n22569 ; n22569_not
g60555 not n27636 ; n27636_not
g60556 not n45690 ; n45690_not
g60557 not n21957 ; n21957_not
g60558 not n38058 ; n38058_not
g60559 not n21894 ; n21894_not
g60560 not n21795 ; n21795_not
g60561 not n21777 ; n21777_not
g60562 not n27816 ; n27816_not
g60563 not n21768 ; n21768_not
g60564 not n21759 ; n21759_not
g60565 not n38139 ; n38139_not
g60566 not n21696 ; n21696_not
g60567 not n38157 ; n38157_not
g60568 not n38184 ; n38184_not
g60569 not n21597 ; n21597_not
g60570 not n24549 ; n24549_not
g60571 not n36636 ; n36636_not
g60572 not n37833 ; n37833_not
g60573 not n27726 ; n27726_not
g60574 not n17457 ; n17457_not
g60575 not n37860 ; n37860_not
g60576 not n37923 ; n37923_not
g60577 not n37734 ; n37734_not
g60578 not n21975 ; n21975_not
g60579 not n27780 ; n27780_not
g60580 not n19572 ; n19572_not
g60581 not n19554 ; n19554_not
g60582 not n28275 ; n28275_not
g60583 not n31848 ; n31848_not
g60584 not n19518 ; n19518_not
g60585 not n16944 ; n16944_not
g60586 not n19509 ; n19509_not
g60587 not n16926 ; n16926_not
g60588 not n44646 ; n44646_not
g60589 not n19437 ; n19437_not
g60590 not n19419 ; n19419_not
g60591 not n15297 ; n15297_not
g60592 not n28329 ; n28329_not
g60593 not n44637 ; n44637_not
g60594 not n39714 ; n39714_not
g60595 not n28176 ; n28176_not
g60596 not n39804 ; n39804_not
g60597 not n19716 ; n19716_not
g60598 not n31794 ; n31794_not
g60599 not n39831 ; n39831_not
g60600 not n39903 ; n39903_not
g60601 not n39930 ; n39930_not
g60602 not n19662 ; n19662_not
g60603 not n19653 ; n19653_not
g60604 not n44754 ; n44754_not
g60605 not n19644 ; n19644_not
g60606 not n10797 ; n10797_not
g60607 not n19194 ; n19194_not
g60608 not n19149 ; n19149_not
g60609 not n44394 ; n44394_not
g60610 not n19158 ; n19158_not
g60611 not n10887 ; n10887_not
g60612 not n40389 ; n40389_not
g60613 not n19095 ; n19095_not
g60614 not n10878 ; n10878_not
g60615 not n19086 ; n19086_not
g60616 not n18726 ; n18726_not
g60617 not n33387 ; n33387_not
g60618 not n19077 ; n19077_not
g60619 not n44367 ; n44367_not
g60620 not n10968 ; n10968_not
g60621 not n18960 ; n18960_not
g60622 not n44619 ; n44619_not
g60623 not n19383 ; n19383_not
g60624 not n44466 ; n44466_not
g60625 not n44493 ; n44493_not
g60626 not n19356 ; n19356_not
g60627 not n31866 ; n31866_not
g60628 not n19338 ; n19338_not
g60629 not n33459 ; n33459_not
g60630 not n40299 ; n40299_not
g60631 not n44475 ; n44475_not
g60632 not n19293 ; n19293_not
g60633 not n19275 ; n19275_not
g60634 not n28383 ; n28383_not
g60635 not n10599 ; n10599_not
g60636 not n10689 ; n10689_not
g60637 not n19167 ; n19167_not
g60638 not n10788 ; n10788_not
g60639 not n28392 ; n28392_not
g60640 not n39048 ; n39048_not
g60641 not n39084 ; n39084_not
g60642 not n39165 ; n39165_not
g60643 not n39183 ; n39183_not
g60644 not n38661 ; n38661_not
g60645 not n19932 ; n19932_not
g60646 not n39246 ; n39246_not
g60647 not n38805 ; n38805_not
g60648 not n38535 ; n38535_not
g60649 not n39309 ; n39309_not
g60650 not n33855 ; n33855_not
g60651 not n20598 ; n20598_not
g60652 not n38625 ; n38625_not
g60653 not n38670 ; n38670_not
g60654 not n38715 ; n38715_not
g60655 not n27906 ; n27906_not
g60656 not n38742 ; n38742_not
g60657 not n38760 ; n38760_not
g60658 not n27915 ; n27915_not
g60659 not n27924 ; n27924_not
g60660 not n38850 ; n38850_not
g60661 not n38931 ; n38931_not
g60662 not n19950 ; n19950_not
g60663 not n28086 ; n28086_not
g60664 not n39606 ; n39606_not
g60665 not n39624 ; n39624_not
g60666 not n28095 ; n28095_not
g60667 not n19752 ; n19752_not
g60668 not n39651 ; n39651_not
g60669 not n19707 ; n19707_not
g60670 not n39327 ; n39327_not
g60671 not n39363 ; n39363_not
g60672 not n39372 ; n39372_not
g60673 not n19842 ; n19842_not
g60674 not n39408 ; n39408_not
g60675 not n39435 ; n39435_not
g60676 not n19815 ; n19815_not
g60677 not n39471 ; n39471_not
g60678 not n39525 ; n39525_not
g60679 not n33675 ; n33675_not
g60680 not n39543 ; n39543_not
g60681 not n33666 ; n33666_not
g60682 not n39552 ; n39552_not
g60683 not n26781 ; n26781_not
g60684 not n25089 ; n25089_not
g60685 not n25098 ; n25098_not
g60686 not n26790 ; n26790_not
g60687 not n16980 ; n16980_not
g60688 not n24990 ; n24990_not
g60689 not n24981 ; n24981_not
g60690 not n36177 ; n36177_not
g60691 not n35880 ; n35880_not
g60692 not n34809 ; n34809_not
g60693 not n30876 ; n30876_not
g60694 not n24936 ; n24936_not
g60695 not n24927 ; n24927_not
g60696 not n47742 ; n47742_not
g60697 not n36258 ; n36258_not
g60698 not n24918 ; n24918_not
g60699 not n47913 ; n47913_not
g60700 not n25485 ; n25485_not
g60701 not n34854 ; n34854_not
g60702 not n47904 ; n47904_not
g60703 not n25476 ; n25476_not
g60704 not n25458 ; n25458_not
g60705 not n25377 ; n25377_not
g60706 not n25278 ; n25278_not
g60707 not n34863 ; n34863_not
g60708 not n25287 ; n25287_not
g60709 not n36096 ; n36096_not
g60710 not n34845 ; n34845_not
g60711 not n47805 ; n47805_not
g60712 not n25197 ; n25197_not
g60713 not n25188 ; n25188_not
g60714 not n25179 ; n25179_not
g60715 not n24792 ; n24792_not
g60716 not n34728 ; n34728_not
g60717 not n47562 ; n47562_not
g60718 not n24783 ; n24783_not
g60719 not n36393 ; n36393_not
g60720 not n26907 ; n26907_not
g60721 not n24774 ; n24774_not
g60722 not n26916 ; n26916_not
g60723 not n47553 ; n47553_not
g60724 not n24756 ; n24756_not
g60725 not n24747 ; n24747_not
g60726 not n17169 ; n17169_not
g60727 not n36429 ; n36429_not
g60728 not n24729 ; n24729_not
g60729 not n24639 ; n24639_not
g60730 not n36456 ; n36456_not
g60731 not n47463 ; n47463_not
g60732 not n36267 ; n36267_not
g60733 not n24891 ; n24891_not
g60734 not n24882 ; n24882_not
g60735 not n16818 ; n16818_not
g60736 not n24873 ; n24873_not
g60737 not n34737 ; n34737_not
g60738 not n34746 ; n34746_not
g60739 not n30957 ; n30957_not
g60740 not n26862 ; n26862_not
g60741 not n47634 ; n47634_not
g60742 not n47607 ; n47607_not
g60743 not n36339 ; n36339_not
g60744 not n24828 ; n24828_not
g60745 not n36348 ; n36348_not
g60746 not n30948 ; n30948_not
g60747 not n48642 ; n48642_not
g60748 not n48624 ; n48624_not
g60749 not n25953 ; n25953_not
g60750 not n48471 ; n48471_not
g60751 not n35448 ; n35448_not
g60752 not n48606 ; n48606_not
g60753 not n25926 ; n25926_not
g60754 not n35493 ; n35493_not
g60755 not n48255 ; n48255_not
g60756 not n48561 ; n48561_not
g60757 not n25863 ; n25863_not
g60758 not n25854 ; n25854_not
g60759 not n35088 ; n35088_not
g60760 not n48552 ; n48552_not
g60761 not n48246 ; n48246_not
g60762 not n35574 ; n35574_not
g60763 not n35079 ; n35079_not
g60764 not n31389 ; n31389_not
g60765 not n26439 ; n26439_not
g60766 not n35196 ; n35196_not
g60767 not n26385 ; n26385_not
g60768 not n49137 ; n49137_not
g60769 not n49038 ; n49038_not
g60770 not n35178 ; n35178_not
g60771 not n48714 ; n48714_not
g60772 not n35268 ; n35268_not
g60773 not n35286 ; n35286_not
g60774 not n35169 ; n35169_not
g60775 not n35349 ; n35349_not
g60776 not n26493 ; n26493_not
g60777 not n35358 ; n35358_not
g60778 not n35295 ; n35295_not
g60779 not n34953 ; n34953_not
g60780 not n25980 ; n25980_not
g60781 not n35394 ; n35394_not
g60782 not n48183 ; n48183_not
g60783 not n35826 ; n35826_not
g60784 not n48174 ; n48174_not
g60785 not n48147 ; n48147_not
g60786 not n35871 ; n35871_not
g60787 not n35862 ; n35862_not
g60788 not n34962 ; n34962_not
g60789 not n25584 ; n25584_not
g60790 not n48084 ; n48084_not
g60791 not n25566 ; n25566_not
g60792 not n48048 ; n48048_not
g60793 not n26727 ; n26727_not
g60794 not n35943 ; n35943_not
g60795 not n25548 ; n25548_not
g60796 not n35952 ; n35952_not
g60797 not n35970 ; n35970_not
g60798 not n26592 ; n26592_not
g60799 not n48534 ; n48534_not
g60800 not n25845 ; n25845_not
g60801 not n48453 ; n48453_not
g60802 not n26619 ; n26619_not
g60803 not n48426 ; n48426_not
g60804 not n34935 ; n34935_not
g60805 not n48408 ; n48408_not
g60806 not n26583 ; n26583_not
g60807 not n48363 ; n48363_not
g60808 not n25764 ; n25764_not
g60809 not n35691 ; n35691_not
g60810 not n25746 ; n25746_not
g60811 not n48345 ; n48345_not
g60812 not n48282 ; n48282_not
g60813 not n26682 ; n26682_not
g60814 not n35772 ; n35772_not
g60815 not n25656 ; n25656_not
g60816 not n46590 ; n46590_not
g60817 not n23568 ; n23568_not
g60818 not n46572 ; n46572_not
g60819 not n27348 ; n27348_not
g60820 not n46527 ; n46527_not
g60821 not n37176 ; n37176_not
g60822 not n23496 ; n23496_not
g60823 not n30687 ; n30687_not
g60824 not n46455 ; n46455_not
g60825 not n23397 ; n23397_not
g60826 not n23388 ; n23388_not
g60827 not n37239 ; n37239_not
g60828 not n46347 ; n46347_not
g60829 not n37257 ; n37257_not
g60830 not n27393 ; n27393_not
g60831 not n23298 ; n23298_not
g60832 not n31659 ; n31659_not
g60833 not n46662 ; n46662_not
g60834 not n46644 ; n46644_not
g60835 not n27258 ; n27258_not
g60836 not n27267 ; n27267_not
g60837 not n27276 ; n27276_not
g60838 not n23694 ; n23694_not
g60839 not n23676 ; n23676_not
g60840 not n34395 ; n34395_not
g60841 not n23658 ; n23658_not
g60842 not n30696 ; n30696_not
g60843 not n23586 ; n23586_not
g60844 not n34377 ; n34377_not
g60845 not n37158 ; n37158_not
g60846 not n23595 ; n23595_not
g60847 not n37167 ; n37167_not
g60848 not n23577 ; n23577_not
g60849 not n37185 ; n37185_not
g60850 not n22929 ; n22929_not
g60851 not n37419 ; n37419_not
g60852 not n22875 ; n22875_not
g60853 not n37446 ; n37446_not
g60854 not n31677 ; n31677_not
g60855 not n37464 ; n37464_not
g60856 not n27528 ; n27528_not
g60857 not n45942 ; n45942_not
g60858 not n37473 ; n37473_not
g60859 not n37482 ; n37482_not
g60860 not n22848 ; n22848_not
g60861 not n45834 ; n45834_not
g60862 not n34197 ; n34197_not
g60863 not n45807 ; n45807_not
g60864 not n37509 ; n37509_not
g60865 not n27294 ; n27294_not
g60866 not n37284 ; n37284_not
g60867 not n23199 ; n23199_not
g60868 not n46284 ; n46284_not
g60869 not n37329 ; n37329_not
g60870 not n27438 ; n27438_not
g60871 not n22992 ; n22992_not
g60872 not n27447 ; n27447_not
g60873 not n22866 ; n22866_not
g60874 not n46275 ; n46275_not
g60875 not n31668 ; n31668_not
g60876 not n27465 ; n27465_not
g60877 not n22983 ; n22983_not
g60878 not n27474 ; n27474_not
g60879 not n37356 ; n37356_not
g60880 not n37149 ; n37149_not
g60881 not n46239 ; n46239_not
g60882 not n46194 ; n46194_not
g60883 not n36582 ; n36582_not
g60884 not n36591 ; n36591_not
g60885 not n47364 ; n47364_not
g60886 not n36645 ; n36645_not
g60887 not n16647 ; n16647_not
g60888 not n47346 ; n47346_not
g60889 not n34566 ; n34566_not
g60890 not n36663 ; n36663_not
g60891 not n36690 ; n36690_not
g60892 not n47328 ; n47328_not
g60893 not n47292 ; n47292_not
g60894 not n34548 ; n34548_not
g60895 not n47274 ; n47274_not
g60896 not n24189 ; n24189_not
g60897 not n36717 ; n36717_not
g60898 not n24684 ; n24684_not
g60899 not n36474 ; n36474_not
g60900 not n34647 ; n34647_not
g60901 not n34674 ; n34674_not
g60902 not n36438 ; n36438_not
g60903 not n36483 ; n36483_not
g60904 not n24657 ; n24657_not
g60905 not n30894 ; n30894_not
g60906 not n36528 ; n36528_not
g60907 not n34638 ; n34638_not
g60908 not n30867 ; n30867_not
g60909 not n34629 ; n34629_not
g60910 not n36555 ; n36555_not
g60911 not n47382 ; n47382_not
g60912 not n36573 ; n36573_not
g60913 not n26970 ; n26970_not
g60914 not n36924 ; n36924_not
g60915 not n47076 ; n47076_not
g60916 not n36933 ; n36933_not
g60917 not n36942 ; n36942_not
g60918 not n27159 ; n27159_not
g60919 not n46923 ; n46923_not
g60920 not n46860 ; n46860_not
g60921 not n34467 ; n34467_not
g60922 not n46815 ; n46815_not
g60923 not n23892 ; n23892_not
g60924 not n46761 ; n46761_not
g60925 not n46734 ; n46734_not
g60926 not n46716 ; n46716_not
g60927 not n23757 ; n23757_not
g60928 not n23838 ; n23838_not
g60929 not n37086 ; n37086_not
g60930 not n36726 ; n36726_not
g60931 not n34539 ; n34539_not
g60932 not n36735 ; n36735_not
g60933 not n36762 ; n36762_not
g60934 not n36771 ; n36771_not
g60935 not n24198 ; n24198_not
g60936 not n36807 ; n36807_not
g60937 not n47193 ; n47193_not
g60938 not n24099 ; n24099_not
g60939 not n27069 ; n27069_not
g60940 not n47175 ; n47175_not
g60941 not n17970 ; n17970_not
g60942 not n27096 ; n27096_not
g60943 not n47085 ; n47085_not
g60944 not n36861 ; n36861_not
g60945 not n36870 ; n36870_not
g60946 not n23964 ; n23964_not
g60947 not n43593 ; n43593_not
g60948 not n29058 ; n29058_not
g60949 not n16782 ; n16782_not
g60950 not n29049 ; n29049_not
g60951 not n12849 ; n12849_not
g60952 not n41937 ; n41937_not
g60953 not n43638 ; n43638_not
g60954 not n41919 ; n41919_not
g60955 not n12795 ; n12795_not
g60956 not n41892 ; n41892_not
g60957 not n16881 ; n16881_not
g60958 not n41883 ; n41883_not
g60959 not n28923 ; n28923_not
g60960 not n41865 ; n41865_not
g60961 not n12777 ; n12777_not
g60962 not n32865 ; n32865_not
g60963 not n41856 ; n41856_not
g60964 not n16935 ; n16935_not
g60965 not n16953 ; n16953_not
g60966 not n16962 ; n16962_not
g60967 not n41829 ; n41829_not
g60968 not n32883 ; n32883_not
g60969 not n41577 ; n41577_not
g60970 not n41793 ; n41793_not
g60971 not n41784 ; n41784_not
g60972 not n17097 ; n17097_not
g60973 not n41775 ; n41775_not
g60974 not n41766 ; n41766_not
g60975 not n43377 ; n43377_not
g60976 not n43467 ; n43467_not
g60977 not n29715 ; n29715_not
g60978 not n16359 ; n16359_not
g60979 not n43485 ; n43485_not
g60980 not n29175 ; n29175_not
g60981 not n16368 ; n16368_not
g60982 not n16386 ; n16386_not
g60983 not n29805 ; n29805_not
g60984 not n29166 ; n29166_not
g60985 not n29157 ; n29157_not
g60986 not n43548 ; n43548_not
g60987 not n29814 ; n29814_not
g60988 not n32739 ; n32739_not
g60989 not n13686 ; n13686_not
g60990 not n15738 ; n15738_not
g60991 not n41991 ; n41991_not
g60992 not n29733 ; n29733_not
g60993 not n32766 ; n32766_not
g60994 not n16575 ; n16575_not
g60995 not n16584 ; n16584_not
g60996 not n29094 ; n29094_not
g60997 not n16593 ; n16593_not
g60998 not n12894 ; n12894_not
g60999 not n41757 ; n41757_not
g61000 not n29085 ; n29085_not
g61001 not n16674 ; n16674_not
g61002 not n16692 ; n16692_not
g61003 not n17628 ; n17628_not
g61004 not n41559 ; n41559_not
g61005 not n43872 ; n43872_not
g61006 not n17664 ; n17664_not
g61007 not n41568 ; n41568_not
g61008 not n17673 ; n17673_not
g61009 not n17682 ; n17682_not
g61010 not n12399 ; n12399_not
g61011 not n17718 ; n17718_not
g61012 not n43881 ; n43881_not
g61013 not n43908 ; n43908_not
g61014 not n41478 ; n41478_not
g61015 not n41379 ; n41379_not
g61016 not n17808 ; n17808_not
g61017 not n17817 ; n17817_not
g61018 not n43935 ; n43935_not
g61019 not n28860 ; n28860_not
g61020 not n41388 ; n41388_not
g61021 not n31992 ; n31992_not
g61022 not n17880 ; n17880_not
g61023 not n33099 ; n33099_not
g61024 not n17907 ; n17907_not
g61025 not n43944 ; n43944_not
g61026 not n17934 ; n17934_not
g61027 not n17943 ; n17943_not
g61028 not n17952 ; n17952_not
g61029 not n28941 ; n28941_not
g61030 not n12678 ; n12678_not
g61031 not n17259 ; n17259_not
g61032 not n12669 ; n12669_not
g61033 not n28932 ; n28932_not
g61034 not n17349 ; n17349_not
g61035 not n43737 ; n43737_not
g61036 not n17376 ; n17376_not
g61037 not n43746 ; n43746_not
g61038 not n17439 ; n17439_not
g61039 not n17448 ; n17448_not
g61040 not n12579 ; n12579_not
g61041 not n32964 ; n32964_not
g61042 not n43782 ; n43782_not
g61043 not n32784 ; n32784_not
g61044 not n32973 ; n32973_not
g61045 not n43809 ; n43809_not
g61046 not n32982 ; n32982_not
g61047 not n41649 ; n41649_not
g61048 not n43827 ; n43827_not
g61049 not n12489 ; n12489_not
g61050 not n17493 ; n17493_not
g61051 not n17556 ; n17556_not
g61052 not n43854 ; n43854_not
g61053 not n14388 ; n14388_not
g61054 not n42837 ; n42837_not
g61055 not n42828 ; n42828_not
g61056 not n32379 ; n32379_not
g61057 not n29544 ; n29544_not
g61058 not n42747 ; n42747_not
g61059 not n14919 ; n14919_not
g61060 not n32388 ; n32388_not
g61061 not n14298 ; n14298_not
g61062 not n29517 ; n29517_not
g61063 not n14928 ; n14928_not
g61064 not n42774 ; n42774_not
g61065 not n29508 ; n29508_not
g61066 not n42738 ; n42738_not
g61067 not n15099 ; n15099_not
g61068 not n14937 ; n14937_not
g61069 not n14199 ; n14199_not
g61070 not n42675 ; n42675_not
g61071 not n29481 ; n29481_not
g61072 not n15288 ; n15288_not
g61073 not n13992 ; n13992_not
g61074 not n42594 ; n42594_not
g61075 not n43197 ; n43197_not
g61076 not n29436 ; n29436_not
g61077 not n13965 ; n13965_not
g61078 not n42576 ; n42576_not
g61079 not n15477 ; n15477_not
g61080 not n15486 ; n15486_not
g61081 not n15495 ; n15495_not
g61082 not n14559 ; n14559_not
g61083 not n14649 ; n14649_not
g61084 not n14676 ; n14676_not
g61085 not n14694 ; n14694_not
g61086 not n29454 ; n29454_not
g61087 not n40983 ; n40983_not
g61088 not n32298 ; n32298_not
g61089 not n43089 ; n43089_not
g61090 not n14496 ; n14496_not
g61091 not n14469 ; n14469_not
g61092 not n14748 ; n14748_not
g61093 not n14757 ; n14757_not
g61094 not n29625 ; n29625_not
g61095 not n14766 ; n14766_not
g61096 not n29616 ; n29616_not
g61097 not n42990 ; n42990_not
g61098 not n29607 ; n29607_not
g61099 not n42981 ; n42981_not
g61100 not n42972 ; n42972_not
g61101 not n38544 ; n38544_not
g61102 not n14775 ; n14775_not
g61103 not n14577 ; n14577_not
g61104 not n42927 ; n42927_not
g61105 not n42936 ; n42936_not
g61106 not n29571 ; n29571_not
g61107 not n40965 ; n40965_not
g61108 not n29553 ; n29553_not
g61109 not n14838 ; n14838_not
g61110 not n29292 ; n29292_not
g61111 not n15855 ; n15855_not
g61112 not n15864 ; n15864_not
g61113 not n15891 ; n15891_not
g61114 not n42297 ; n42297_not
g61115 not n29760 ; n29760_not
g61116 not n42288 ; n42288_not
g61117 not n13776 ; n13776_not
g61118 not n13758 ; n13758_not
g61119 not n29265 ; n29265_not
g61120 not n13749 ; n13749_not
g61121 not n43359 ; n43359_not
g61122 not n15927 ; n15927_not
g61123 not n13695 ; n13695_not
g61124 not n13677 ; n13677_not
g61125 not n15945 ; n15945_not
g61126 not n43386 ; n43386_not
g61127 not n13587 ; n13587_not
g61128 not n29229 ; n29229_not
g61129 not n15981 ; n15981_not
g61130 not n32667 ; n32667_not
g61131 not n15990 ; n15990_not
g61132 not n15279 ; n15279_not
g61133 not n42198 ; n42198_not
g61134 not n16089 ; n16089_not
g61135 not n32676 ; n32676_not
g61136 not n32685 ; n32685_not
g61137 not n13479 ; n13479_not
g61138 not n15756 ; n15756_not
g61139 not n29184 ; n29184_not
g61140 not n32487 ; n32487_not
g61141 not n29391 ; n29391_not
g61142 not n13947 ; n13947_not
g61143 not n15576 ; n15576_not
g61144 not n29724 ; n29724_not
g61145 not n42495 ; n42495_not
g61146 not n29373 ; n29373_not
g61147 not n13938 ; n13938_not
g61148 not n15639 ; n15639_not
g61149 not n42477 ; n42477_not
g61150 not n15648 ; n15648_not
g61151 not n29364 ; n29364_not
g61152 not n42459 ; n42459_not
g61153 not n13929 ; n13929_not
g61154 not n15684 ; n15684_not
g61155 not n15693 ; n15693_not
g61156 not n15729 ; n15729_not
g61157 not n29751 ; n29751_not
g61158 not n32577 ; n32577_not
g61159 not n29337 ; n29337_not
g61160 not n15774 ; n15774_not
g61161 not n13839 ; n13839_not
g61162 not n29328 ; n29328_not
g61163 not n15783 ; n15783_not
g61164 not n32595 ; n32595_not
g61165 not n29319 ; n29319_not
g61166 not n13794 ; n13794_not
g61167 not n15846 ; n15846_not
g61168 not n40938 ; n40938_not
g61169 not n11859 ; n11859_not
g61170 not n18564 ; n18564_not
g61171 not n18573 ; n18573_not
g61172 not n28680 ; n28680_not
g61173 not n40893 ; n40893_not
g61174 not n40884 ; n40884_not
g61175 not n28671 ; n28671_not
g61176 not n40875 ; n40875_not
g61177 not n40866 ; n40866_not
g61178 not n18591 ; n18591_not
g61179 not n29922 ; n29922_not
g61180 not n40848 ; n40848_not
g61181 not n18609 ; n18609_not
g61182 not n44079 ; n44079_not
g61183 not n16791 ; n16791_not
g61184 not n18645 ; n18645_not
g61185 not n18195 ; n18195_not
g61186 not n18177 ; n18177_not
g61187 not n11949 ; n11949_not
g61188 not n18294 ; n18294_not
g61189 not n11895 ; n11895_not
g61190 not n18339 ; n18339_not
g61191 not n18348 ; n18348_not
g61192 not n18375 ; n18375_not
g61193 not n28752 ; n28752_not
g61194 not n43845 ; n43845_not
g61195 not n18438 ; n18438_not
g61196 not n18447 ; n18447_not
g61197 not n18465 ; n18465_not
g61198 not n18474 ; n18474_not
g61199 not n18483 ; n18483_not
g61200 not n18492 ; n18492_not
g61201 not n43575 ; n43575_not
g61202 not n18528 ; n18528_not
g61203 not n11679 ; n11679_not
g61204 not n18834 ; n18834_not
g61205 not n11598 ; n11598_not
g61206 not n18870 ; n18870_not
g61207 not n44178 ; n44178_not
g61208 not n28473 ; n28473_not
g61209 not n44196 ; n44196_not
g61210 not n40596 ; n40596_not
g61211 not n40587 ; n40587_not
g61212 not n28509 ; n28509_not
g61213 not n10977 ; n10977_not
g61214 not n40569 ; n40569_not
g61215 not n18915 ; n18915_not
g61216 not n43719 ; n43719_not
g61217 not n28482 ; n28482_not
g61218 not n18942 ; n18942_not
g61219 not n18654 ; n18654_not
g61220 not n11769 ; n11769_not
g61221 not n18663 ; n18663_not
g61222 not n18672 ; n18672_not
g61223 not n28617 ; n28617_not
g61224 not n18627 ; n18627_not
g61225 not n33288 ; n33288_not
g61226 not n16539 ; n16539_not
g61227 not n18717 ; n18717_not
g61228 not n33297 ; n33297_not
g61229 not n18735 ; n18735_not
g61230 not n18762 ; n18762_not
g61231 not n18771 ; n18771_not
g61232 not n28572 ; n28572_not
g61233 not n39642 ; n39642_not
g61234 not n40659 ; n40659_not
g61235 not n40686 ; n40686_not
g61236 not n18816 ; n18816_not
g61237 not n40677 ; n40677_not
g61238 not n41298 ; n41298_not
g61239 not n17961 ; n17961_not
g61240 not n43962 ; n43962_not
g61241 not n43980 ; n43980_not
g61242 not n18069 ; n18069_not
g61243 not n18096 ; n18096_not
g61244 not n28806 ; n28806_not
g61245 not n18168 ; n18168_not
g61246 not n40795 ; n40795_not
g61247 not n24892 ; n24892_not
g61248 not n13948 ; n13948_not
g61249 not n36268 ; n36268_not
g61250 not n42496 ; n42496_not
g61251 not n18754 ; n18754_not
g61252 not n40993 ; n40993_not
g61253 not n16639 ; n16639_not
g61254 not n38707 ; n38707_not
g61255 not n17863 ; n17863_not
g61256 not n15568 ; n15568_not
g61257 not n15559 ; n15559_not
g61258 not n13957 ; n13957_not
g61259 not n19366 ; n19366_not
g61260 not n44638 ; n44638_not
g61261 not n17845 ; n17845_not
g61262 not n13849 ; n13849_not
g61263 not n14965 ; n14965_not
g61264 not n24973 ; n24973_not
g61265 not n13885 ; n13885_not
g61266 not n17980 ; n17980_not
g61267 not n19528 ; n19528_not
g61268 not n38365 ; n38365_not
g61269 not n42469 ; n42469_not
g61270 not n18691 ; n18691_not
g61271 not n15658 ; n15658_not
g61272 not n41596 ; n41596_not
g61273 not n47680 ; n47680_not
g61274 not n44647 ; n44647_not
g61275 not n47716 ; n47716_not
g61276 not n41389 ; n41389_not
g61277 not n17485 ; n17485_not
g61278 not n36295 ; n36295_not
g61279 not n36286 ; n36286_not
g61280 not n18727 ; n18727_not
g61281 not n43189 ; n43189_not
g61282 not n36097 ; n36097_not
g61283 not n35485 ; n35485_not
g61284 not n47833 ; n47833_not
g61285 not n36088 ; n36088_not
g61286 not n42595 ; n42595_not
g61287 not n36079 ; n36079_not
g61288 not n19348 ; n19348_not
g61289 not n25297 ; n25297_not
g61290 not n15298 ; n15298_not
g61291 not n34783 ; n34783_not
g61292 not n35980 ; n35980_not
g61293 not n47842 ; n47842_not
g61294 not n25369 ; n25369_not
g61295 not n35890 ; n35890_not
g61296 not n40885 ; n40885_not
g61297 not n25396 ; n25396_not
g61298 not n42649 ; n42649_not
g61299 not n18781 ; n18781_not
g61300 not n36196 ; n36196_not
g61301 not n19384 ; n19384_not
g61302 not n36187 ; n36187_not
g61303 not n42568 ; n42568_not
g61304 not n38680 ; n38680_not
g61305 not n15397 ; n15397_not
g61306 not n41299 ; n41299_not
g61307 not n20797 ; n20797_not
g61308 not n34765 ; n34765_not
g61309 not n47761 ; n47761_not
g61310 not n42586 ; n42586_not
g61311 not n25189 ; n25189_not
g61312 not n15388 ; n15388_not
g61313 not n40687 ; n40687_not
g61314 not n34891 ; n34891_not
g61315 not n15379 ; n15379_not
g61316 not n38545 ; n38545_not
g61317 not n17791 ; n17791_not
g61318 not n47392 ; n47392_not
g61319 not n24577 ; n24577_not
g61320 not n36259 ; n36259_not
g61321 not n24586 ; n24586_not
g61322 not n39463 ; n39463_not
g61323 not n47419 ; n47419_not
g61324 not n47446 ; n47446_not
g61325 not n36529 ; n36529_not
g61326 not n24478 ; n24478_not
g61327 not n47455 ; n47455_not
g61328 not n24649 ; n24649_not
g61329 not n36493 ; n36493_not
g61330 not n42298 ; n42298_not
g61331 not n17917 ; n17917_not
g61332 not n39841 ; n39841_not
g61333 not n38608 ; n38608_not
g61334 not n36637 ; n36637_not
g61335 not n36628 ; n36628_not
g61336 not n17548 ; n17548_not
g61337 not n47356 ; n47356_not
g61338 not n24487 ; n24487_not
g61339 not n13687 ; n13687_not
g61340 not n40786 ; n40786_not
g61341 not n39904 ; n39904_not
g61342 not n13696 ; n13696_not
g61343 not n47383 ; n47383_not
g61344 not n39913 ; n39913_not
g61345 not n24559 ; n24559_not
g61346 not n18628 ; n18628_not
g61347 not n20878 ; n20878_not
g61348 not n24568 ; n24568_not
g61349 not n15919 ; n15919_not
g61350 not n19582 ; n19582_not
g61351 not n44098 ; n44098_not
g61352 not n15766 ; n15766_not
g61353 not n19573 ; n19573_not
g61354 not n19564 ; n19564_not
g61355 not n15775 ; n15775_not
g61356 not n43297 ; n43297_not
g61357 not n38419 ; n38419_not
g61358 not n15757 ; n15757_not
g61359 not n36385 ; n36385_not
g61360 not n40759 ; n40759_not
g61361 not n19537 ; n19537_not
g61362 not n13876 ; n13876_not
g61363 not n19429 ; n19429_not
g61364 not n36484 ; n36484_not
g61365 not n15856 ; n15856_not
g61366 not n38356 ; n38356_not
g61367 not n16819 ; n16819_not
g61368 not n38761 ; n38761_not
g61369 not n15847 ; n15847_not
g61370 not n13786 ; n13786_not
g61371 not n17818 ; n17818_not
g61372 not n42379 ; n42379_not
g61373 not n36448 ; n36448_not
g61374 not n38752 ; n38752_not
g61375 not n47491 ; n47491_not
g61376 not n15784 ; n15784_not
g61377 not n36439 ; n36439_not
g61378 not n47509 ; n47509_not
g61379 not n19627 ; n19627_not
g61380 not n44089 ; n44089_not
g61381 not n47518 ; n47518_not
g61382 not n19168 ; n19168_not
g61383 not n35548 ; n35548_not
g61384 not n35539 ; n35539_not
g61385 not n39481 ; n39481_not
g61386 not n20599 ; n20599_not
g61387 not n35494 ; n35494_not
g61388 not n42964 ; n42964_not
g61389 not n35458 ; n35458_not
g61390 not n25918 ; n25918_not
g61391 not n14776 ; n14776_not
g61392 not n25927 ; n25927_not
g61393 not n42973 ; n42973_not
g61394 not n44296 ; n44296_not
g61395 not n40399 ; n40399_not
g61396 not n10888 ; n10888_not
g61397 not n25936 ; n25936_not
g61398 not n40579 ; n40579_not
g61399 not n25639 ; n25639_not
g61400 not n48409 ; n48409_not
g61401 not n48418 ; n48418_not
g61402 not n25828 ; n25828_not
g61403 not n10798 ; n10798_not
g61404 not n48445 ; n48445_not
g61405 not n14848 ; n14848_not
g61406 not n48490 ; n48490_not
g61407 not n19186 ; n19186_not
g61408 not n40588 ; n40588_not
g61409 not n42928 ; n42928_not
g61410 not n17971 ; n17971_not
g61411 not n20698 ; n20698_not
g61412 not n35557 ; n35557_not
g61413 not n44395 ; n44395_not
g61414 not n25594 ; n25594_not
g61415 not n17944 ; n17944_not
g61416 not n48661 ; n48661_not
g61417 not n17953 ; n17953_not
g61418 not n18925 ; n18925_not
g61419 not n21679 ; n21679_not
g61420 not n26269 ; n26269_not
g61421 not n26278 ; n26278_not
g61422 not n18709 ; n18709_not
g61423 not n18916 ; n18916_not
g61424 not n49138 ; n49138_not
g61425 not n26377 ; n26377_not
g61426 not n18952 ; n18952_not
g61427 not n14587 ; n14587_not
g61428 not n14578 ; n14578_not
g61429 not n14659 ; n14659_not
g61430 not n10978 ; n10978_not
g61431 not n19096 ; n19096_not
g61432 not n35377 ; n35377_not
g61433 not n43954 ; n43954_not
g61434 not n35368 ; n35368_not
g61435 not n43099 ; n43099_not
g61436 not n35359 ; n35359_not
g61437 not n20689 ; n20689_not
g61438 not n38581 ; n38581_not
g61439 not n34990 ; n34990_not
g61440 not n44467 ; n44467_not
g61441 not n25567 ; n25567_not
g61442 not n14956 ; n14956_not
g61443 not n14974 ; n14974_not
g61444 not n16657 ; n16657_not
g61445 not n35863 ; n35863_not
g61446 not n48094 ; n48094_not
g61447 not n17926 ; n17926_not
g61448 not n38617 ; n38617_not
g61449 not n38464 ; n38464_not
g61450 not n14299 ; n14299_not
g61451 not n15199 ; n15199_not
g61452 not n17890 ; n17890_not
g61453 not n14785 ; n14785_not
g61454 not n25486 ; n25486_not
g61455 not n44485 ; n44485_not
g61456 not n25387 ; n25387_not
g61457 not n40669 ; n40669_not
g61458 not n47932 ; n47932_not
g61459 not n35971 ; n35971_not
g61460 not n38662 ; n38662_not
g61461 not n38653 ; n38653_not
g61462 not n14983 ; n14983_not
g61463 not n47941 ; n47941_not
g61464 not n42739 ; n42739_not
g61465 not n25558 ; n25558_not
g61466 not n35674 ; n35674_not
g61467 not n44179 ; n44179_not
g61468 not n38518 ; n38518_not
g61469 not n48364 ; n48364_not
g61470 not n14884 ; n14884_not
g61471 not n25774 ; n25774_not
g61472 not n48247 ; n48247_not
g61473 not n35656 ; n35656_not
g61474 not n48373 ; n48373_not
g61475 not n35638 ; n35638_not
g61476 not n35629 ; n35629_not
g61477 not n48382 ; n48382_not
g61478 not n25792 ; n25792_not
g61479 not n48391 ; n48391_not
g61480 not n42775 ; n42775_not
g61481 not n25819 ; n25819_not
g61482 not n35845 ; n35845_not
g61483 not n25648 ; n25648_not
g61484 not n19276 ; n19276_not
g61485 not n48175 ; n48175_not
g61486 not n35809 ; n35809_not
g61487 not n42766 ; n42766_not
g61488 not n16945 ; n16945_not
g61489 not n48193 ; n48193_not
g61490 not n35764 ; n35764_not
g61491 not n10699 ; n10699_not
g61492 not n18862 ; n18862_not
g61493 not n35737 ; n35737_not
g61494 not n48337 ; n48337_not
g61495 not n16684 ; n16684_not
g61496 not n42793 ; n42793_not
g61497 not n14875 ; n14875_not
g61498 not n35683 ; n35683_not
g61499 not n25756 ; n25756_not
g61500 not n37465 ; n37465_not
g61501 not n16990 ; n16990_not
g61502 not n35575 ; n35575_not
g61503 not n39373 ; n39373_not
g61504 not n45808 ; n45808_not
g61505 not n22768 ; n22768_not
g61506 not n38437 ; n38437_not
g61507 not n11878 ; n11878_not
g61508 not n45286 ; n45286_not
g61509 not n38905 ; n38905_not
g61510 not n45817 ; n45817_not
g61511 not n38833 ; n38833_not
g61512 not n41848 ; n41848_not
g61513 not n16936 ; n16936_not
g61514 not n37492 ; n37492_not
g61515 not n41767 ; n41767_not
g61516 not n37636 ; n37636_not
g61517 not n41785 ; n41785_not
g61518 not n39382 ; n39382_not
g61519 not n16765 ; n16765_not
g61520 not n22687 ; n22687_not
g61521 not n37573 ; n37573_not
g61522 not n22966 ; n22966_not
g61523 not n41893 ; n41893_not
g61524 not n37384 ; n37384_not
g61525 not n17692 ; n17692_not
g61526 not n37375 ; n37375_not
g61527 not n36970 ; n36970_not
g61528 not n37366 ; n37366_not
g61529 not n16873 ; n16873_not
g61530 not n22975 ; n22975_not
g61531 not n37339 ; n37339_not
g61532 not n46249 ; n46249_not
g61533 not n46258 ; n46258_not
g61534 not n12787 ; n12787_not
g61535 not n39472 ; n39472_not
g61536 not n37348 ; n37348_not
g61537 not n39490 ; n39490_not
g61538 not n38725 ; n38725_not
g61539 not n37294 ; n37294_not
g61540 not n39418 ; n39418_not
g61541 not n45880 ; n45880_not
g61542 not n37474 ; n37474_not
g61543 not n41857 ; n41857_not
g61544 not n39409 ; n39409_not
g61545 not n19825 ; n19825_not
g61546 not n46096 ; n46096_not
g61547 not n43873 ; n43873_not
g61548 not n39445 ; n39445_not
g61549 not n22867 ; n22867_not
g61550 not n16909 ; n16909_not
g61551 not n37447 ; n37447_not
g61552 not n18466 ; n18466_not
g61553 not n46069 ; n46069_not
g61554 not n41875 ; n41875_not
g61555 not n22948 ; n22948_not
g61556 not n43855 ; n43855_not
g61557 not n22957 ; n22957_not
g61558 not n11977 ; n11977_not
g61559 not n21985 ; n21985_not
g61560 not n21994 ; n21994_not
g61561 not n17476 ; n17476_not
g61562 not n37951 ; n37951_not
g61563 not n37942 ; n37942_not
g61564 not n37933 ; n37933_not
g61565 not n11968 ; n11968_not
g61566 not n17467 ; n17467_not
g61567 not n37915 ; n37915_not
g61568 not n37906 ; n37906_not
g61569 not n17449 ; n17449_not
g61570 not n43864 ; n43864_not
g61571 not n37852 ; n37852_not
g61572 not n37825 ; n37825_not
g61573 not n18286 ; n18286_not
g61574 not n41587 ; n41587_not
g61575 not n39067 ; n39067_not
g61576 not n43990 ; n43990_not
g61577 not n43837 ; n43837_not
g61578 not n21877 ; n21877_not
g61579 not n21886 ; n21886_not
g61580 not n39094 ; n39094_not
g61581 not n38491 ; n38491_not
g61582 not n38059 ; n38059_not
g61583 not n19960 ; n19960_not
g61584 not n18178 ; n18178_not
g61585 not n19951 ; n19951_not
g61586 not n21958 ; n21958_not
g61587 not n41659 ; n41659_not
g61588 not n39184 ; n39184_not
g61589 not n17494 ; n17494_not
g61590 not n38194 ; n38194_not
g61591 not n37591 ; n37591_not
g61592 not n18367 ; n18367_not
g61593 not n45646 ; n45646_not
g61594 not n39319 ; n39319_not
g61595 not n11896 ; n11896_not
g61596 not n39328 ; n39328_not
g61597 not n37672 ; n37672_not
g61598 not n37663 ; n37663_not
g61599 not n45664 ; n45664_not
g61600 not n41758 ; n41758_not
g61601 not n45673 ; n45673_not
g61602 not n19861 ; n19861_not
g61603 not n45709 ; n45709_not
g61604 not n22498 ; n22498_not
g61605 not n45718 ; n45718_not
g61606 not n19852 ; n19852_not
g61607 not n17089 ; n17089_not
g61608 not n17395 ; n17395_not
g61609 not n37645 ; n37645_not
g61610 not n17386 ; n17386_not
g61611 not n38950 ; n38950_not
g61612 not n17377 ; n17377_not
g61613 not n37807 ; n37807_not
g61614 not n39229 ; n39229_not
g61615 not n45349 ; n45349_not
g61616 not n37762 ; n37762_not
g61617 not n37753 ; n37753_not
g61618 not n43729 ; n43729_not
g61619 not n18358 ; n18358_not
g61620 not n37735 ; n37735_not
g61621 not n39256 ; n39256_not
g61622 not n12688 ; n12688_not
g61623 not n39283 ; n39283_not
g61624 not n41668 ; n41668_not
g61625 not n45196 ; n45196_not
g61626 not n46951 ; n46951_not
g61627 not n47068 ; n47068_not
g61628 not n36925 ; n36925_not
g61629 not n39661 ; n39661_not
g61630 not n18088 ; n18088_not
g61631 not n40876 ; n40876_not
g61632 not n36907 ; n36907_not
g61633 not n39706 ; n39706_not
g61634 not n16279 ; n16279_not
g61635 not n16297 ; n16297_not
g61636 not n36853 ; n36853_not
g61637 not n18079 ; n18079_not
g61638 not n39724 ; n39724_not
g61639 not n47167 ; n47167_not
g61640 not n43459 ; n43459_not
g61641 not n39742 ; n39742_not
g61642 not n14596 ; n14596_not
g61643 not n23848 ; n23848_not
g61644 not n46744 ; n46744_not
g61645 not n41488 ; n41488_not
g61646 not n46807 ; n46807_not
g61647 not n23875 ; n23875_not
g61648 not n19753 ; n19753_not
g61649 not n20959 ; n20959_not
g61650 not n23866 ; n23866_not
g61651 not n11788 ; n11788_not
g61652 not n43495 ; n43495_not
g61653 not n23938 ; n23938_not
g61654 not n39670 ; n39670_not
g61655 not n23947 ; n23947_not
g61656 not n46915 ; n46915_not
g61657 not n16378 ; n16378_not
g61658 not n16369 ; n16369_not
g61659 not n17755 ; n17755_not
g61660 not n36709 ; n36709_not
g61661 not n17575 ; n17575_not
g61662 not n47248 ; n47248_not
g61663 not n11779 ; n11779_not
g61664 not n39823 ; n39823_not
g61665 not n47284 ; n47284_not
g61666 not n13579 ; n13579_not
g61667 not n15973 ; n15973_not
g61668 not n15937 ; n15937_not
g61669 not n36619 ; n36619_not
g61670 not n47347 ; n47347_not
g61671 not n17782 ; n17782_not
g61672 not n15946 ; n15946_not
g61673 not n36466 ; n36466_not
g61674 not n36655 ; n36655_not
g61675 not n24397 ; n24397_not
g61676 not n13399 ; n13399_not
g61677 not n47185 ; n47185_not
g61678 not n36826 ; n36826_not
g61679 not n36547 ; n36547_not
g61680 not n16189 ; n16189_not
g61681 not n36817 ; n36817_not
g61682 not n43909 ; n43909_not
g61683 not n39643 ; n39643_not
g61684 not n16099 ; n16099_not
g61685 not n36574 ; n36574_not
g61686 not n36736 ; n36736_not
g61687 not n43918 ; n43918_not
g61688 not n15991 ; n15991_not
g61689 not n12859 ; n12859_not
g61690 not n46375 ; n46375_not
g61691 not n46429 ; n46429_not
g61692 not n12868 ; n12868_not
g61693 not n12877 ; n12877_not
g61694 not n12886 ; n12886_not
g61695 not n38860 ; n38860_not
g61696 not n46474 ; n46474_not
g61697 not n39535 ; n39535_not
g61698 not n38275 ; n38275_not
g61699 not n18538 ; n18538_not
g61700 not n23569 ; n23569_not
g61701 not n16666 ; n16666_not
g61702 not n40957 ; n40957_not
g61703 not n39553 ; n39553_not
g61704 not n46285 ; n46285_not
g61705 not n41929 ; n41929_not
g61706 not n16792 ; n16792_not
g61707 not n41947 ; n41947_not
g61708 not n19807 ; n19807_not
g61709 not n19735 ; n19735_not
g61710 not n17557 ; n17557_not
g61711 not n37267 ; n37267_not
g61712 not n39517 ; n39517_not
g61713 not n41956 ; n41956_not
g61714 not n37276 ; n37276_not
g61715 not n16783 ; n16783_not
g61716 not n38266 ; n38266_not
g61717 not n37258 ; n37258_not
g61718 not n39526 ; n39526_not
g61719 not n16747 ; n16747_not
g61720 not n39616 ; n39616_not
g61721 not n23758 ; n23758_not
g61722 not n46582 ; n46582_not
g61723 not n20968 ; n20968_not
g61724 not n23767 ; n23767_not
g61725 not n23776 ; n23776_not
g61726 not n16486 ; n16486_not
g61727 not n23785 ; n23785_not
g61728 not n12976 ; n12976_not
g61729 not n46681 ; n46681_not
g61730 not n37078 ; n37078_not
g61731 not n46708 ; n46708_not
g61732 not n37069 ; n37069_not
g61733 not n23749 ; n23749_not
g61734 not n18583 ; n18583_not
g61735 not n12985 ; n12985_not
g61736 not n16396 ; n16396_not
g61737 not n18547 ; n18547_not
g61738 not n23578 ; n23578_not
g61739 not n39562 ; n39562_not
g61740 not n39571 ; n39571_not
g61741 not n11869 ; n11869_not
g61742 not n43576 ; n43576_not
g61743 not n39580 ; n39580_not
g61744 not n41497 ; n41497_not
g61745 not n41974 ; n41974_not
g61746 not n23659 ; n23659_not
g61747 not n46591 ; n46591_not
g61748 not n23668 ; n23668_not
g61749 not n46609 ; n46609_not
g61750 not n16558 ; n16558_not
g61751 not n23686 ; n23686_not
g61752 not n17746 ; n17746_not
g61753 not n16549 ; n16549_not
g61754 not n33289 ; n33289_not
g61755 not n28618 ; n28618_not
g61756 not n31795 ; n31795_not
g61757 not n28627 ; n28627_not
g61758 not n27079 ; n27079_not
g61759 not n29905 ; n29905_not
g61760 not n29455 ; n29455_not
g61761 not n28636 ; n28636_not
g61762 not n34495 ; n34495_not
g61763 not n28645 ; n28645_not
g61764 not n33829 ; n33829_not
g61765 not n32785 ; n32785_not
g61766 not n34486 ; n34486_not
g61767 not n29068 ; n29068_not
g61768 not n34477 ; n34477_not
g61769 not n27745 ; n27745_not
g61770 not n26737 ; n26737_not
g61771 not n34558 ; n34558_not
g61772 not n31894 ; n31894_not
g61773 not n34927 ; n34927_not
g61774 not n26728 ; n26728_not
g61775 not n26980 ; n26980_not
g61776 not n33757 ; n33757_not
g61777 not n29374 ; n29374_not
g61778 not n27934 ; n27934_not
g61779 not n28573 ; n28573_not
g61780 not n33784 ; n33784_not
g61781 not n30787 ; n30787_not
g61782 not n31786 ; n31786_not
g61783 not n33775 ; n33775_not
g61784 not n34981 ; n34981_not
g61785 not n28591 ; n28591_not
g61786 not n29707 ; n29707_not
g61787 not n33928 ; n33928_not
g61788 not n30499 ; n30499_not
g61789 not n27853 ; n27853_not
g61790 not n33937 ; n33937_not
g61791 not n31696 ; n31696_not
g61792 not n34396 ; n34396_not
g61793 not n29545 ; n29545_not
g61794 not n33946 ; n33946_not
g61795 not n27286 ; n27286_not
g61796 not n29428 ; n29428_not
g61797 not n29554 ; n29554_not
g61798 not n34378 ; n34378_not
g61799 not n26584 ; n26584_not
g61800 not n35098 ; n35098_not
g61801 not n29563 ; n29563_not
g61802 not n31498 ; n31498_not
g61803 not n33982 ; n33982_not
g61804 not n29572 ; n29572_not
g61805 not n32875 ; n32875_not
g61806 not n28654 ; n28654_not
g61807 not n26683 ; n26683_not
g61808 not n29491 ; n29491_not
g61809 not n27178 ; n27178_not
g61810 not n31597 ; n31597_not
g61811 not n33874 ; n33874_not
g61812 not n30985 ; n30985_not
g61813 not n29509 ; n29509_not
g61814 not n28744 ; n28744_not
g61815 not n29059 ; n29059_not
g61816 not n29419 ; n29419_not
g61817 not n29770 ; n29770_not
g61818 not n29518 ; n29518_not
g61819 not n31984 ; n31984_not
g61820 not n29527 ; n29527_not
g61821 not n32839 ; n32839_not
g61822 not n31687 ; n31687_not
g61823 not n26638 ; n26638_not
g61824 not n27871 ; n27871_not
g61825 not n28771 ; n28771_not
g61826 not n26746 ; n26746_not
g61827 not n30598 ; n30598_not
g61828 not n26809 ; n26809_not
g61829 not n29842 ; n29842_not
g61830 not n28168 ; n28168_not
g61831 not n30589 ; n30589_not
g61832 not n33478 ; n33478_not
g61833 not n33595 ; n33595_not
g61834 not n32578 ; n32578_not
g61835 not n33487 ; n33487_not
g61836 not n34684 ; n34684_not
g61837 not n33469 ; n33469_not
g61838 not n32668 ; n32668_not
g61839 not n34675 ; n34675_not
g61840 not n29329 ; n29329_not
g61841 not n34666 ; n34666_not
g61842 not n26764 ; n26764_not
g61843 not n34657 ; n34657_not
g61844 not n26854 ; n26854_not
g61845 not n33559 ; n33559_not
g61846 not n34756 ; n34756_not
g61847 not n29284 ; n29284_not
g61848 not n34747 ; n34747_not
g61849 not n29275 ; n29275_not
g61850 not n31876 ; n31876_not
g61851 not n28267 ; n28267_not
g61852 not n26881 ; n26881_not
g61853 not n29860 ; n29860_not
g61854 not n32587 ; n32587_not
g61855 not n28177 ; n28177_not
g61856 not n34819 ; n34819_not
g61857 not n28294 ; n28294_not
g61858 not n32695 ; n32695_not
g61859 not n33379 ; n33379_not
g61860 not n29185 ; n29185_not
g61861 not n26773 ; n26773_not
g61862 not n28474 ; n28474_not
g61863 not n29356 ; n29356_not
g61864 not n29347 ; n29347_not
g61865 not n34576 ; n34576_not
g61866 not n33739 ; n33739_not
g61867 not n28492 ; n28492_not
g61868 not n28528 ; n28528_not
g61869 not n34567 ; n34567_not
g61870 not n27961 ; n27961_not
g61871 not n33748 ; n33748_not
g61872 not n28384 ; n28384_not
g61873 not n32569 ; n32569_not
g61874 not n31768 ; n31768_not
g61875 not n28096 ; n28096_not
g61876 not n34837 ; n34837_not
g61877 not n28393 ; n28393_not
g61878 not n32677 ; n32677_not
g61879 not n26755 ; n26755_not
g61880 not n29194 ; n29194_not
g61881 not n28447 ; n28447_not
g61882 not n34594 ; n34594_not
g61883 not n33667 ; n33667_not
g61884 not n33388 ; n33388_not
g61885 not n33397 ; n33397_not
g61886 not n26971 ; n26971_not
g61887 not n34873 ; n34873_not
g61888 not n33676 ; n33676_not
g61889 not n31885 ; n31885_not
g61890 not n32929 ; n32929_not
g61891 not n27682 ; n27682_not
g61892 not n31957 ; n31957_not
g61893 not n29635 ; n29635_not
g61894 not n31579 ; n31579_not
g61895 not n27493 ; n27493_not
g61896 not n29950 ; n29950_not
g61897 not n29923 ; n29923_not
g61898 not n31399 ; n31399_not
g61899 not n27628 ; n27628_not
g61900 not n34279 ; n34279_not
g61901 not n28663 ; n28663_not
g61902 not n32893 ; n32893_not
g61903 not n30796 ; n30796_not
g61904 not n31975 ; n31975_not
g61905 not n27457 ; n27457_not
g61906 not n26296 ; n26296_not
g61907 not n29671 ; n29671_not
g61908 not n27736 ; n27736_not
g61909 not n29743 ; n29743_not
g61910 not n26557 ; n26557_not
g61911 not n28960 ; n28960_not
g61912 not n27547 ; n27547_not
g61913 not n27385 ; n27385_not
g61914 not n28924 ; n28924_not
g61915 not n32938 ; n32938_not
g61916 not n34189 ; n34189_not
g61917 not n31939 ; n31939_not
g61918 not n29716 ; n29716_not
g61919 not n28870 ; n28870_not
g61920 not n26287 ; n26287_not
g61921 not n30886 ; n30886_not
g61922 not n29644 ; n29644_not
g61923 not n32947 ; n32947_not
g61924 not n31858 ; n31858_not
g61925 not n26494 ; n26494_not
g61926 not n28861 ; n28861_not
g61927 not n34198 ; n34198_not
g61928 not n30859 ; n30859_not
g61929 not n27592 ; n27592_not
g61930 not n29590 ; n29590_not
g61931 not n34918 ; n34918_not
g61932 not n27692 ; n27692_not
g61933 not n33686 ; n33686_not
g61934 not n37754 ; n37754_not
g61935 not n36593 ; n36593_not
g61936 not n46583 ; n46583_not
g61937 not n48185 ; n48185_not
g61938 not n29258 ; n29258_not
g61939 not n29816 ; n29816_not
g61940 not n26837 ; n26837_not
g61941 not n36548 ; n36548_not
g61942 not n27980 ; n27980_not
g61943 not n12959 ; n12959_not
g61944 not n43577 ; n43577_not
g61945 not n27665 ; n27665_not
g61946 not n37673 ; n37673_not
g61947 not n37691 ; n37691_not
g61948 not n37682 ; n37682_not
g61949 not n36566 ; n36566_not
g61950 not n26963 ; n26963_not
g61951 not n37439 ; n37439_not
g61952 not n39455 ; n39455_not
g61953 not n12968 ; n12968_not
g61954 not n14498 ; n14498_not
g61955 not n48194 ; n48194_not
g61956 not n19781 ; n19781_not
g61957 not n27656 ; n27656_not
g61958 not n36584 ; n36584_not
g61959 not n37727 ; n37727_not
g61960 not n29663 ; n29663_not
g61961 not n19790 ; n19790_not
g61962 not n15695 ; n15695_not
g61963 not n30698 ; n30698_not
g61964 not n15668 ; n15668_not
g61965 not n37394 ; n37394_not
g61966 not n36656 ; n36656_not
g61967 not n36638 ; n36638_not
g61968 not n39356 ; n39356_not
g61969 not n39338 ; n39338_not
g61970 not n27962 ; n27962_not
g61971 not n15659 ; n15659_not
g61972 not n22967 ; n22967_not
g61973 not n36665 ; n36665_not
g61974 not n14669 ; n14669_not
g61975 not n19871 ; n19871_not
g61976 not n46655 ; n46655_not
g61977 not n39293 ; n39293_not
g61978 not n36674 ; n36674_not
g61979 not n39266 ; n39266_not
g61980 not n30896 ; n30896_not
g61981 not n37376 ; n37376_not
g61982 not n39239 ; n39239_not
g61983 not n37844 ; n37844_not
g61984 not n22976 ; n22976_not
g61985 not n27485 ; n27485_not
g61986 not n37367 ; n37367_not
g61987 not n27467 ; n27467_not
g61988 not n19907 ; n19907_not
g61989 not n14678 ; n14678_not
g61990 not n24299 ; n24299_not
g61991 not n47456 ; n47456_not
g61992 not n37466 ; n37466_not
g61993 not n24479 ; n24479_not
g61994 not n17882 ; n17882_not
g61995 not n48158 ; n48158_not
g61996 not n36728 ; n36728_not
g61997 not n46619 ; n46619_not
g61998 not n39437 ; n39437_not
g61999 not n40868 ; n40868_not
g62000 not n40994 ; n40994_not
g62001 not n19826 ; n19826_not
g62002 not n36629 ; n36629_not
g62003 not n48149 ; n48149_not
g62004 not n42569 ; n42569_not
g62005 not n39428 ; n39428_not
g62006 not n44657 ; n44657_not
g62007 not n37772 ; n37772_not
g62008 not n12995 ; n12995_not
g62009 not n47474 ; n47474_not
g62010 not n24398 ; n24398_not
g62011 not n29654 ; n29654_not
g62012 not n19835 ; n19835_not
g62013 not n39392 ; n39392_not
g62014 not n26882 ; n26882_not
g62015 not n22697 ; n22697_not
g62016 not n46493 ; n46493_not
g62017 not n39860 ; n39860_not
g62018 not n43667 ; n43667_not
g62019 not n48329 ; n48329_not
g62020 not n26891 ; n26891_not
g62021 not n27557 ; n27557_not
g62022 not n39662 ; n39662_not
g62023 not n15785 ; n15785_not
g62024 not n22688 ; n22688_not
g62025 not n33596 ; n33596_not
g62026 not n39806 ; n39806_not
g62027 not n43658 ; n43658_not
g62028 not n24776 ; n24776_not
g62029 not n24767 ; n24767_not
g62030 not n12797 ; n12797_not
g62031 not n27539 ; n27539_not
g62032 not n24758 ; n24758_not
g62033 not n26918 ; n26918_not
g62034 not n42389 ; n42389_not
g62035 not n24875 ; n24875_not
g62036 not n24686 ; n24686_not
g62037 not n19646 ; n19646_not
g62038 not n27575 ; n27575_not
g62039 not n29285 ; n29285_not
g62040 not n22769 ; n22769_not
g62041 not n37538 ; n37538_not
g62042 not n27566 ; n27566_not
g62043 not n46448 ; n46448_not
g62044 not n24866 ; n24866_not
g62045 not n39149 ; n39149_not
g62046 not n19655 ; n19655_not
g62047 not n24857 ; n24857_not
g62048 not n34748 ; n34748_not
g62049 not n31967 ; n31967_not
g62050 not n37493 ; n37493_not
g62051 not n24839 ; n24839_not
g62052 not n22796 ; n22796_not
g62053 not n27593 ; n27593_not
g62054 not n19664 ; n19664_not
g62055 not n26873 ; n26873_not
g62056 not n34739 ; n34739_not
g62057 not n43685 ; n43685_not
g62058 not n30689 ; n30689_not
g62059 not n39581 ; n39581_not
g62060 not n15839 ; n15839_not
g62061 not n46484 ; n46484_not
g62062 not n15749 ; n15749_not
g62063 not n39680 ; n39680_not
g62064 not n26945 ; n26945_not
g62065 not n37655 ; n37655_not
g62066 not n38825 ; n38825_not
g62067 not n39644 ; n39644_not
g62068 not n22859 ; n22859_not
g62069 not n34649 ; n34649_not
g62070 not n19763 ; n19763_not
g62071 not n39545 ; n39545_not
g62072 not n24596 ; n24596_not
g62073 not n46565 ; n46565_not
g62074 not n47429 ; n47429_not
g62075 not n47438 ; n47438_not
g62076 not n28088 ; n28088_not
g62077 not n19772 ; n19772_not
g62078 not n46574 ; n46574_not
g62079 not n28079 ; n28079_not
g62080 not n26954 ; n26954_not
g62081 not n45845 ; n45845_not
g62082 not n39743 ; n39743_not
g62083 not n29843 ; n29843_not
g62084 not n39761 ; n39761_not
g62085 not n27548 ; n27548_not
g62086 not n39752 ; n39752_not
g62087 not n48284 ; n48284_not
g62088 not n42398 ; n42398_not
g62089 not n37484 ; n37484_not
g62090 not n37628 ; n37628_not
g62091 not n24695 ; n24695_not
g62092 not n39734 ; n39734_not
g62093 not n34685 ; n34685_not
g62094 not n19736 ; n19736_not
g62095 not n37619 ; n37619_not
g62096 not n12869 ; n12869_not
g62097 not n39716 ; n39716_not
g62098 not n24677 ; n24677_not
g62099 not n32579 ; n32579_not
g62100 not n29339 ; n29339_not
g62101 not n15758 ; n15758_not
g62102 not n26936 ; n26936_not
g62103 not n37475 ; n37475_not
g62104 not n27638 ; n27638_not
g62105 not n31859 ; n31859_not
g62106 not n46943 ; n46943_not
g62107 not n13769 ; n13769_not
g62108 not n33866 ; n33866_not
g62109 not n38456 ; n38456_not
g62110 not n13778 ; n13778_not
g62111 not n38447 ; n38447_not
g62112 not n37277 ; n37277_not
g62113 not n42776 ; n42776_not
g62114 not n13787 ; n13787_not
g62115 not n33893 ; n33893_not
g62116 not n20789 ; n20789_not
g62117 not n37079 ; n37079_not
g62118 not n38429 ; n38429_not
g62119 not n14768 ; n14768_not
g62120 not n29537 ; n29537_not
g62121 not n38483 ; n38483_not
g62122 not n47618 ; n47618_not
g62123 not n29762 ; n29762_not
g62124 not n23777 ; n23777_not
g62125 not n38069 ; n38069_not
g62126 not n27395 ; n27395_not
g62127 not n13796 ; n13796_not
g62128 not n36971 ; n36971_not
g62129 not n37970 ; n37970_not
g62130 not n38528 ; n38528_not
g62131 not n27881 ; n27881_not
g62132 not n20699 ; n20699_not
g62133 not n40985 ; n40985_not
g62134 not n34469 ; n34469_not
g62135 not n40859 ; n40859_not
g62136 not n27089 ; n27089_not
g62137 not n14966 ; n14966_not
g62138 not n47582 ; n47582_not
g62139 not n27755 ; n27755_not
g62140 not n19475 ; n19475_not
g62141 not n21986 ; n21986_not
g62142 not n42587 ; n42587_not
g62143 not n27188 ; n27188_not
g62144 not n23885 ; n23885_not
g62145 not n27197 ; n27197_not
g62146 not n47825 ; n47825_not
g62147 not n31778 ; n31778_not
g62148 not n21788 ; n21788_not
g62149 not n38258 ; n38258_not
g62150 not n13895 ; n13895_not
g62151 not n29753 ; n29753_not
g62152 not n38249 ; n38249_not
g62153 not n27836 ; n27836_not
g62154 not n14759 ; n14759_not
g62155 not n33965 ; n33965_not
g62156 not n37187 ; n37187_not
g62157 not n47681 ; n47681_not
g62158 not n21599 ; n21599_not
g62159 not n14795 ; n14795_not
g62160 not n33983 ; n33983_not
g62161 not n47726 ; n47726_not
g62162 not n27368 ; n27368_not
g62163 not n14786 ; n14786_not
g62164 not n42947 ; n42947_not
g62165 not n38177 ; n38177_not
g62166 not n44729 ; n44729_not
g62167 not n30959 ; n30959_not
g62168 not n13859 ; n13859_not
g62169 not n27359 ; n27359_not
g62170 not n38168 ; n38168_not
g62171 not n38159 ; n38159_not
g62172 not n33992 ; n33992_not
g62173 not n31589 ; n31589_not
g62174 not n47087 ; n47087_not
g62175 not n47627 ; n47627_not
g62176 not n27863 ; n27863_not
g62177 not n14894 ; n14894_not
g62178 not n38357 ; n38357_not
g62179 not n38348 ; n38348_not
g62180 not n38078 ; n38078_not
g62181 not n27854 ; n27854_not
g62182 not n42974 ; n42974_not
g62183 not n20969 ; n20969_not
g62184 not n21878 ; n21878_not
g62185 not n21869 ; n21869_not
g62186 not n47771 ; n47771_not
g62187 not n42965 ; n42965_not
g62188 not n16856 ; n16856_not
g62189 not n29591 ; n29591_not
g62190 not n14777 ; n14777_not
g62191 not n14876 ; n14876_not
g62192 not n42839 ; n42839_not
g62193 not n13868 ; n13868_not
g62194 not n47672 ; n47672_not
g62195 not n38591 ; n38591_not
g62196 not n23597 ; n23597_not
g62197 not n43298 ; n43298_not
g62198 not n14858 ; n14858_not
g62199 not n38276 ; n38276_not
g62200 not n15569 ; n15569_not
g62201 not n19916 ; n19916_not
g62202 not n36773 ; n36773_not
g62203 not n30788 ; n30788_not
g62204 not n15488 ; n15488_not
g62205 not n13985 ; n13985_not
g62206 not n36782 ; n36782_not
g62207 not n27476 ; n27476_not
g62208 not n14687 ; n14687_not
g62209 not n22985 ; n22985_not
g62210 not n27728 ; n27728_not
g62211 not n38960 ; n38960_not
g62212 not n43379 ; n43379_not
g62213 not n29780 ; n29780_not
g62214 not n29870 ; n29870_not
g62215 not n38942 ; n38942_not
g62216 not n38933 ; n38933_not
g62217 not n33794 ; n33794_not
g62218 not n38924 ; n38924_not
g62219 not n46790 ; n46790_not
g62220 not n38744 ; n38744_not
g62221 not n22994 ; n22994_not
g62222 not n13598 ; n13598_not
g62223 not n27458 ; n27458_not
g62224 not n38843 ; n38843_not
g62225 not n27926 ; n27926_not
g62226 not n27944 ; n27944_not
g62227 not n26990 ; n26990_not
g62228 not n48077 ; n48077_not
g62229 not n37862 ; n37862_not
g62230 not n33767 ; n33767_not
g62231 not n19943 ; n19943_not
g62232 not n43478 ; n43478_not
g62233 not n38645 ; n38645_not
g62234 not n48059 ; n48059_not
g62235 not n43469 ; n43469_not
g62236 not n39194 ; n39194_not
g62237 not n42488 ; n42488_not
g62238 not n26864 ; n26864_not
g62239 not n39176 ; n39176_not
g62240 not n15596 ; n15596_not
g62241 not n36746 ; n36746_not
g62242 not n46691 ; n46691_not
g62243 not n36719 ; n36719_not
g62244 not n33776 ; n33776_not
g62245 not n47492 ; n47492_not
g62246 not n36755 ; n36755_not
g62247 not n15587 ; n15587_not
g62248 not n36368 ; n36368_not
g62249 not n36764 ; n36764_not
g62250 not n15578 ; n15578_not
g62251 not n38762 ; n38762_not
g62252 not n37934 ; n37934_not
g62253 not n30986 ; n30986_not
g62254 not n36917 ; n36917_not
g62255 not n37556 ; n37556_not
g62256 not n37943 ; n37943_not
g62257 not n27890 ; n27890_not
g62258 not n14597 ; n14597_not
g62259 not n37961 ; n37961_not
g62260 not n36935 ; n36935_not
g62261 not n38636 ; n38636_not
g62262 not n38609 ; n38609_not
g62263 not n38627 ; n38627_not
g62264 not n33848 ; n33848_not
g62265 not n47573 ; n47573_not
g62266 not n42686 ; n42686_not
g62267 not n23957 ; n23957_not
g62268 not n46907 ; n46907_not
g62269 not n47168 ; n47168_not
g62270 not n29708 ; n29708_not
g62271 not n29933 ; n29933_not
g62272 not n29447 ; n29447_not
g62273 not n38834 ; n38834_not
g62274 not n36845 ; n36845_not
g62275 not n37907 ; n37907_not
g62276 not n13976 ; n13976_not
g62277 not n36854 ; n36854_not
g62278 not n30995 ; n30995_not
g62279 not n34289 ; n34289_not
g62280 not n46835 ; n46835_not
g62281 not n38807 ; n38807_not
g62282 not n36863 ; n36863_not
g62283 not n34496 ; n34496_not
g62284 not n43397 ; n43397_not
g62285 not n37763 ; n37763_not
g62286 not n36881 ; n36881_not
g62287 not n38573 ; n38573_not
g62288 not n27791 ; n27791_not
g62289 not n28853 ; n28853_not
g62290 not n18719 ; n18719_not
g62291 not n41399 ; n41399_not
g62292 not n33299 ; n33299_not
g62293 not n43892 ; n43892_not
g62294 not n17855 ; n17855_not
g62295 not n45971 ; n45971_not
g62296 not n17189 ; n17189_not
g62297 not n18773 ; n18773_not
g62298 not n40697 ; n40697_not
g62299 not n17837 ; n17837_not
g62300 not n25892 ; n25892_not
g62301 not n25973 ; n25973_not
g62302 not n44378 ; n44378_not
g62303 not n35882 ; n35882_not
g62304 not n40679 ; n40679_not
g62305 not n40688 ; n40688_not
g62306 not n18809 ; n18809_not
g62307 not n41795 ; n41795_not
g62308 not n28574 ; n28574_not
g62309 not n18818 ; n18818_not
g62310 not n16667 ; n16667_not
g62311 not n25946 ; n25946_not
g62312 not n28628 ; n28628_not
g62313 not n32777 ; n32777_not
g62314 not n26558 ; n26558_not
g62315 not n18665 ; n18665_not
g62316 not n40787 ; n40787_not
g62317 not n18656 ; n18656_not
g62318 not n11978 ; n11978_not
g62319 not n34991 ; n34991_not
g62320 not n25658 ; n25658_not
g62321 not n26549 ; n26549_not
g62322 not n43937 ; n43937_not
g62323 not n35828 ; n35828_not
g62324 not n40778 ; n40778_not
g62325 not n43919 ; n43919_not
g62326 not n16595 ; n16595_not
g62327 not n18683 ; n18683_not
g62328 not n18674 ; n18674_not
g62329 not n49067 ; n49067_not
g62330 not n10898 ; n10898_not
g62331 not n32894 ; n32894_not
g62332 not n29078 ; n29078_not
g62333 not n28547 ; n28547_not
g62334 not n26738 ; n26738_not
g62335 not n28961 ; n28961_not
g62336 not n17765 ; n17765_not
g62337 not n16973 ; n16973_not
g62338 not n28880 ; n28880_not
g62339 not n25991 ; n25991_not
g62340 not n16496 ; n16496_not
g62341 not n18890 ; n18890_not
g62342 not n40598 ; n40598_not
g62343 not n28538 ; n28538_not
g62344 not n18881 ; n18881_not
g62345 not n35963 ; n35963_not
g62346 not n40589 ; n40589_not
g62347 not n17756 ; n17756_not
g62348 not n43586 ; n43586_not
g62349 not n41768 ; n41768_not
g62350 not n35981 ; n35981_not
g62351 not n34775 ; n34775_not
g62352 not n16469 ; n16469_not
g62353 not n18917 ; n18917_not
g62354 not n35396 ; n35396_not
g62355 not n32759 ; n32759_not
g62356 not n28565 ; n28565_not
g62357 not n16955 ; n16955_not
g62358 not n17828 ; n17828_not
g62359 not n35891 ; n35891_not
g62360 not n16919 ; n16919_not
g62361 not n17819 ; n17819_not
g62362 not n18845 ; n18845_not
g62363 not n25586 ; n25586_not
g62364 not n16937 ; n16937_not
g62365 not n26387 ; n26387_not
g62366 not n43865 ; n43865_not
g62367 not n25982 ; n25982_not
g62368 not n35918 ; n35918_not
g62369 not n35387 ; n35387_not
g62370 not n35909 ; n35909_not
g62371 not n28556 ; n28556_not
g62372 not n29096 ; n29096_not
g62373 not n43496 ; n43496_not
g62374 not n16946 ; n16946_not
g62375 not n16568 ; n16568_not
g62376 not n17774 ; n17774_not
g62377 not n35945 ; n35945_not
g62378 not n28763 ; n28763_not
g62379 not n26666 ; n26666_not
g62380 not n41948 ; n41948_not
g62381 not n35558 ; n35558_not
g62382 not n32849 ; n32849_not
g62383 not n35648 ; n35648_not
g62384 not n45728 ; n45728_not
g62385 not n45827 ; n45827_not
g62386 not n25775 ; n25775_not
g62387 not n45737 ; n45737_not
g62388 not n25856 ; n25856_not
g62389 not n28745 ; n28745_not
g62390 not n35675 ; n35675_not
g62391 not n25766 ; n25766_not
g62392 not n35684 ; n35684_not
g62393 not n18089 ; n18089_not
g62394 not n41966 ; n41966_not
g62395 not n28808 ; n28808_not
g62396 not n26675 ; n26675_not
g62397 not n35693 ; n35693_not
g62398 not n28736 ; n28736_not
g62399 not n31688 ; n31688_not
g62400 not n28772 ; n28772_not
g62401 not n25838 ; n25838_not
g62402 not n45809 ; n45809_not
g62403 not n18278 ; n18278_not
g62404 not n35594 ; n35594_not
g62405 not n31697 ; n31697_not
g62406 not n28781 ; n28781_not
g62407 not n26648 ; n26648_not
g62408 not n16892 ; n16892_not
g62409 not n18197 ; n18197_not
g62410 not n41885 ; n41885_not
g62411 not n18368 ; n18368_not
g62412 not n26657 ; n26657_not
g62413 not n16838 ; n16838_not
g62414 not n18188 ; n18188_not
g62415 not n16829 ; n16829_not
g62416 not n16757 ; n16757_not
g62417 not n35567 ; n35567_not
g62418 not n25847 ; n25847_not
g62419 not n31985 ; n31985_not
g62420 not n18179 ; n18179_not
g62421 not n25784 ; n25784_not
g62422 not n45638 ; n45638_not
g62423 not n28844 ; n28844_not
g62424 not n17927 ; n17927_not
g62425 not n17873 ; n17873_not
g62426 not n16694 ; n16694_not
g62427 not n45926 ; n45926_not
g62428 not n32885 ; n32885_not
g62429 not n18593 ; n18593_not
g62430 not n35774 ; n35774_not
g62431 not n28727 ; n28727_not
g62432 not n28655 ; n28655_not
g62433 not n49049 ; n49049_not
g62434 not n35783 ; n35783_not
g62435 not n45278 ; n45278_not
g62436 not n18629 ; n18629_not
g62437 not n49058 ; n49058_not
g62438 not n32858 ; n32858_not
g62439 not n25865 ; n25865_not
g62440 not n41975 ; n41975_not
g62441 not n41849 ; n41849_not
g62442 not n25739 ; n25739_not
g62443 not n48824 ; n48824_not
g62444 not n43991 ; n43991_not
g62445 not n45683 ; n45683_not
g62446 not n26684 ; n26684_not
g62447 not n28826 ; n28826_not
g62448 not n28835 ; n28835_not
g62449 not n40958 ; n40958_not
g62450 not n48815 ; n48815_not
g62451 not n45872 ; n45872_not
g62452 not n29069 ; n29069_not
g62453 not n45656 ; n45656_not
g62454 not n18548 ; n18548_not
g62455 not n18557 ; n18557_not
g62456 not n41984 ; n41984_not
g62457 not n18566 ; n18566_not
g62458 not n35756 ; n35756_not
g62459 not n19376 ; n19376_not
g62460 not n28349 ; n28349_not
g62461 not n11789 ; n11789_not
g62462 not n11798 ; n11798_not
g62463 not n33497 ; n33497_not
g62464 not n14984 ; n14984_not
g62465 not n46259 ; n46259_not
g62466 not n17549 ; n17549_not
g62467 not n24983 ; n24983_not
g62468 not n14993 ; n14993_not
g62469 not n31949 ; n31949_not
g62470 not n15929 ; n15929_not
g62471 not n26468 ; n26468_not
g62472 not n34829 ; n34829_not
g62473 not n36188 ; n36188_not
g62474 not n32984 ; n32984_not
g62475 not n32975 ; n32975_not
g62476 not n24947 ; n24947_not
g62477 not n36197 ; n36197_not
g62478 not n26288 ; n26288_not
g62479 not n19484 ; n19484_not
g62480 not n19187 ; n19187_not
g62481 not n19259 ; n19259_not
g62482 not n19268 ; n19268_not
g62483 not n41588 ; n41588_not
g62484 not n19277 ; n19277_not
g62485 not n26189 ; n26189_not
g62486 not n46187 ; n46187_not
g62487 not n28376 ; n28376_not
g62488 not n17585 ; n17585_not
g62489 not n26477 ; n26477_not
g62490 not n17576 ; n17576_not
g62491 not n48518 ; n48518_not
g62492 not n26198 ; n26198_not
g62493 not n41489 ; n41489_not
g62494 not n28367 ; n28367_not
g62495 not n17567 ; n17567_not
g62496 not n48482 ; n48482_not
g62497 not n19358 ; n19358_not
g62498 not n28358 ; n28358_not
g62499 not n26459 ; n26459_not
g62500 not n46349 ; n46349_not
g62501 not n15884 ; n15884_not
g62502 not n28268 ; n28268_not
g62503 not n26846 ; n26846_not
g62504 not n26396 ; n26396_not
g62505 not n31877 ; n31877_not
g62506 not n42299 ; n42299_not
g62507 not n19592 ; n19592_not
g62508 not n36278 ; n36278_not
g62509 not n28925 ; n28925_not
g62510 not n32768 ; n32768_not
g62511 not n34919 ; n34919_not
g62512 not n28259 ; n28259_not
g62513 not n41696 ; n41696_not
g62514 not n35198 ; n35198_not
g62515 not n19637 ; n19637_not
g62516 not n26855 ; n26855_not
g62517 not n29852 ; n29852_not
g62518 not n38861 ; n38861_not
g62519 not n32957 ; n32957_not
g62520 not n28295 ; n28295_not
g62521 not n28907 ; n28907_not
g62522 not n24974 ; n24974_not
g62523 not n44279 ; n44279_not
g62524 not n29249 ; n29249_not
g62525 not n46295 ; n46295_not
g62526 not n41669 ; n41669_not
g62527 not n24965 ; n24965_not
g62528 not n19529 ; n19529_not
g62529 not n17486 ; n17486_not
g62530 not n43757 ; n43757_not
g62531 not n35189 ; n35189_not
g62532 not n19538 ; n19538_not
g62533 not n28286 ; n28286_not
g62534 not n29276 ; n29276_not
g62535 not n26369 ; n26369_not
g62536 not n32966 ; n32966_not
g62537 not n41678 ; n41678_not
g62538 not n19547 ; n19547_not
g62539 not n26378 ; n26378_not
g62540 not n28916 ; n28916_not
g62541 not n18971 ; n18971_not
g62542 not n16298 ; n16298_not
g62543 not n19079 ; n19079_not
g62544 not n44396 ; n44396_not
g62545 not n16379 ; n16379_not
g62546 not n32687 ; n32687_not
g62547 not n28439 ; n28439_not
g62548 not n25478 ; n25478_not
g62549 not n18980 ; n18980_not
g62550 not n34865 ; n34865_not
g62551 not n16199 ; n16199_not
g62552 not n17666 ; n17666_not
g62553 not n26486 ; n26486_not
g62554 not n16289 ; n16289_not
g62555 not n12599 ; n12599_not
g62556 not n46088 ; n46088_not
g62557 not n48590 ; n48590_not
g62558 not n28448 ; n28448_not
g62559 not n29915 ; n29915_not
g62560 not n32696 ; n32696_not
g62561 not n18944 ; n18944_not
g62562 not n48617 ; n48617_not
g62563 not n28277 ; n28277_not
g62564 not n18935 ; n18935_not
g62565 not n28754 ; n28754_not
g62566 not n18953 ; n18953_not
g62567 not n35990 ; n35990_not
g62568 not n18962 ; n18962_not
g62569 not n34856 ; n34856_not
g62570 not n19178 ; n19178_not
g62571 not n26765 ; n26765_not
g62572 not n11969 ; n11969_not
g62573 not n41579 ; n41579_not
g62574 not n25298 ; n25298_not
g62575 not n17657 ; n17657_not
g62576 not n25379 ; n25379_not
g62577 not n17747 ; n17747_not
g62578 not n31886 ; n31886_not
g62579 not n45684 ; n45684_not
g62580 not n28809 ; n28809_not
g62581 not n33957 ; n33957_not
g62582 not n16758 ; n16758_not
g62583 not n41688 ; n41688_not
g62584 not n45693 ; n45693_not
g62585 not n17775 ; n17775_not
g62586 not n37836 ; n37836_not
g62587 not n32868 ; n32868_not
g62588 not n16749 ; n16749_not
g62589 not n17478 ; n17478_not
g62590 not n28818 ; n28818_not
g62591 not n14589 ; n14589_not
g62592 not n28872 ; n28872_not
g62593 not n42885 ; n42885_not
g62594 not n17892 ; n17892_not
g62595 not n20889 ; n20889_not
g62596 not n37863 ; n37863_not
g62597 not n37854 ; n37854_not
g62598 not n41697 ; n41697_not
g62599 not n14886 ; n14886_not
g62600 not n16884 ; n16884_not
g62601 not n45477 ; n45477_not
g62602 not n45189 ; n45189_not
g62603 not n14679 ; n14679_not
g62604 not n27729 ; n27729_not
g62605 not n29547 ; n29547_not
g62606 not n17847 ; n17847_not
g62607 not n47367 ; n47367_not
g62608 not n18189 ; n18189_not
g62609 not n28791 ; n28791_not
g62610 not n45495 ; n45495_not
g62611 not n28980 ; n28980_not
g62612 not n37890 ; n37890_not
g62613 not n32859 ; n32859_not
g62614 not n42795 ; n42795_not
g62615 not n37809 ; n37809_not
g62616 not n28926 ; n28926_not
g62617 not n47349 ; n47349_not
g62618 not n17766 ; n17766_not
g62619 not n37557 ; n37557_not
g62620 not n14868 ; n14868_not
g62621 not n29682 ; n29682_not
g62622 not n38286 ; n38286_not
g62623 not n41679 ; n41679_not
g62624 not n41886 ; n41886_not
g62625 not n42993 ; n42993_not
g62626 not n27675 ; n27675_not
g62627 not n16992 ; n16992_not
g62628 not n28854 ; n28854_not
g62629 not n47169 ; n47169_not
g62630 not n41598 ; n41598_not
g62631 not n16983 ; n16983_not
g62632 not n21897 ; n21897_not
g62633 not n37692 ; n37692_not
g62634 not n28863 ; n28863_not
g62635 not n27792 ; n27792_not
g62636 not n37683 ; n37683_not
g62637 not n42975 ; n42975_not
g62638 not n38079 ; n38079_not
g62639 not n21888 ; n21888_not
g62640 not n47295 ; n47295_not
g62641 not n14499 ; n14499_not
g62642 not n16974 ; n16974_not
g62643 not n21996 ; n21996_not
g62644 not n37584 ; n37584_not
g62645 not n29664 ; n29664_not
g62646 not n29619 ; n29619_not
g62647 not n16776 ; n16776_not
g62648 not n47259 ; n47259_not
g62649 not n21987 ; n21987_not
g62650 not n47268 ; n47268_not
g62651 not n37980 ; n37980_not
g62652 not n21978 ; n21978_not
g62653 not n16767 ; n16767_not
g62654 not n14769 ; n14769_not
g62655 not n21969 ; n21969_not
g62656 not n37728 ; n37728_not
g62657 not n17649 ; n17649_not
g62658 not n37719 ; n37719_not
g62659 not n37746 ; n37746_not
g62660 not n27774 ; n27774_not
g62661 not n29583 ; n29583_not
g62662 not n41787 ; n41787_not
g62663 not n37647 ; n37647_not
g62664 not n41589 ; n41589_not
g62665 not n47196 ; n47196_not
g62666 not n17937 ; n17937_not
g62667 not n28683 ; n28683_not
g62668 not n32985 ; n32985_not
g62669 not n37917 ; n37917_not
g62670 not n42939 ; n42939_not
g62671 not n17946 ; n17946_not
g62672 not n17955 ; n17955_not
g62673 not n17964 ; n17964_not
g62674 not n27819 ; n27819_not
g62675 not n17685 ; n17685_not
g62676 not n17982 ; n17982_not
g62677 not n37656 ; n37656_not
g62678 not n38196 ; n38196_not
g62679 not n17568 ; n17568_not
g62680 not n37665 ; n37665_not
g62681 not n38097 ; n38097_not
g62682 not n47178 ; n47178_not
g62683 not n27747 ; n27747_not
g62684 not n42966 ; n42966_not
g62685 not n17838 ; n17838_not
g62686 not n29592 ; n29592_not
g62687 not n29628 ; n29628_not
g62688 not n21798 ; n21798_not
g62689 not n28845 ; n28845_not
g62690 not n21789 ; n21789_not
g62691 not n17676 ; n17676_not
g62692 not n42948 ; n42948_not
g62693 not n17919 ; n17919_not
g62694 not n27738 ; n27738_not
g62695 not n32994 ; n32994_not
g62696 not n18981 ; n18981_not
g62697 not n19746 ; n19746_not
g62698 not n32499 ; n32499_not
g62699 not n18990 ; n18990_not
g62700 not n15687 ; n15687_not
g62701 not n33696 ; n33696_not
g62702 not n39492 ; n39492_not
g62703 not n39483 ; n39483_not
g62704 not n19809 ; n19809_not
g62705 not n19089 ; n19089_not
g62706 not n46584 ; n46584_not
g62707 not n39519 ; n39519_not
g62708 not n28449 ; n28449_not
g62709 not n18738 ; n18738_not
g62710 not n39528 ; n39528_not
g62711 not n19098 ; n19098_not
g62712 not n39537 ; n39537_not
g62713 not n33399 ; n33399_not
g62714 not n38853 ; n38853_not
g62715 not n19782 ; n19782_not
g62716 not n27972 ; n27972_not
g62717 not n38745 ; n38745_not
g62718 not n39564 ; n39564_not
g62719 not n29196 ; n29196_not
g62720 not n39573 ; n39573_not
g62721 not n19773 ; n19773_not
g62722 not n19197 ; n19197_not
g62723 not n32679 ; n32679_not
g62724 not n39618 ; n39618_not
g62725 not n28395 ; n28395_not
g62726 not n18837 ; n18837_not
g62727 not n42489 ; n42489_not
g62728 not n29097 ; n29097_not
g62729 not n19944 ; n19944_not
g62730 not n27936 ; n27936_not
g62731 not n16569 ; n16569_not
g62732 not n18846 ; n18846_not
g62733 not n27945 ; n27945_not
g62734 not n46674 ; n46674_not
g62735 not n19917 ; n19917_not
g62736 not n38691 ; n38691_not
g62737 not n29367 ; n29367_not
g62738 not n39258 ; n39258_not
g62739 not n39267 ; n39267_not
g62740 not n39168 ; n39168_not
g62741 not n39159 ; n39159_not
g62742 not n29169 ; n29169_not
g62743 not n19827 ; n19827_not
g62744 not n15678 ; n15678_not
g62745 not n19836 ; n19836_not
g62746 not n18936 ; n18936_not
g62747 not n19845 ; n19845_not
g62748 not n18918 ; n18918_not
g62749 not n39393 ; n39393_not
g62750 not n18909 ; n18909_not
g62751 not n39339 ; n39339_not
g62752 not n19683 ; n19683_not
g62753 not n39294 ; n39294_not
g62754 not n18882 ; n18882_not
g62755 not n46665 ; n46665_not
g62756 not n39285 ; n39285_not
g62757 not n19485 ; n19485_not
g62758 not n39807 ; n39807_not
g62759 not n28296 ; n28296_not
g62760 not n28287 ; n28287_not
g62761 not n39843 ; n39843_not
g62762 not n29268 ; n29268_not
g62763 not n19458 ; n19458_not
g62764 not n39825 ; n39825_not
g62765 not n39861 ; n39861_not
g62766 not n28197 ; n28197_not
g62767 not n19548 ; n19548_not
g62768 not n46494 ; n46494_not
g62769 not n39942 ; n39942_not
g62770 not n39951 ; n39951_not
g62771 not n39960 ; n39960_not
g62772 not n39591 ; n39591_not
g62773 not n46467 ; n46467_not
g62774 not n19557 ; n19557_not
g62775 not n19674 ; n19674_not
g62776 not n19575 ; n19575_not
g62777 not n19665 ; n19665_not
g62778 not n46395 ; n46395_not
g62779 not n46458 ; n46458_not
g62780 not n46359 ; n46359_not
g62781 not n29295 ; n29295_not
g62782 not n15849 ; n15849_not
g62783 not n46377 ; n46377_not
g62784 not n15867 ; n15867_not
g62785 not n19692 ; n19692_not
g62786 not n39627 ; n39627_not
g62787 not n46557 ; n46557_not
g62788 not n39645 ; n39645_not
g62789 not n19755 ; n19755_not
g62790 not n28386 ; n28386_not
g62791 not n19269 ; n19269_not
g62792 not n15894 ; n15894_not
g62793 not n46197 ; n46197_not
g62794 not n39681 ; n39681_not
g62795 not n46539 ; n46539_not
g62796 not n19287 ; n19287_not
g62797 not n28377 ; n28377_not
g62798 not n19728 ; n19728_not
g62799 not n38970 ; n38970_not
g62800 not n46278 ; n46278_not
g62801 not n39771 ; n39771_not
g62802 not n39726 ; n39726_not
g62803 not n42399 ; n42399_not
g62804 not n15966 ; n15966_not
g62805 not n33498 ; n33498_not
g62806 not n39735 ; n39735_not
g62807 not n15975 ; n15975_not
g62808 not n15984 ; n15984_not
g62809 not n33597 ; n33597_not
g62810 not n28368 ; n28368_not
g62811 not n14949 ; n14949_not
g62812 not n33876 ; n33876_not
g62813 not n46935 ; n46935_not
g62814 not n18477 ; n18477_not
g62815 not n41967 ; n41967_not
g62816 not n18486 ; n18486_not
g62817 not n45855 ; n45855_not
g62818 not n38556 ; n38556_not
g62819 not n27882 ; n27882_not
g62820 not n38565 ; n38565_not
g62821 not n18495 ; n18495_not
g62822 not n38583 ; n38583_not
g62823 not n38592 ; n38592_not
g62824 not n14976 ; n14976_not
g62825 not n45846 ; n45846_not
g62826 not n14994 ; n14994_not
g62827 not n29493 ; n29493_not
g62828 not n27891 ; n27891_not
g62829 not n33849 ; n33849_not
g62830 not n38619 ; n38619_not
g62831 not n40968 ; n40968_not
g62832 not n28728 ; n28728_not
g62833 not n18549 ; n18549_not
g62834 not n45882 ; n45882_not
g62835 not n29484 ; n29484_not
g62836 not n45918 ; n45918_not
g62837 not n18576 ; n18576_not
g62838 not n38664 ; n38664_not
g62839 not n38529 ; n38529_not
g62840 not n38673 ; n38673_not
g62841 not n46881 ; n46881_not
g62842 not n16875 ; n16875_not
g62843 not n27864 ; n27864_not
g62844 not n27765 ; n27765_not
g62845 not n38367 ; n38367_not
g62846 not n28773 ; n28773_not
g62847 not n46971 ; n46971_not
g62848 not n38376 ; n38376_not
g62849 not n28692 ; n28692_not
g62850 not n16479 ; n16479_not
g62851 not n33885 ; n33885_not
g62852 not n18369 ; n18369_not
g62853 not n16857 ; n16857_not
g62854 not n18378 ; n18378_not
g62855 not n33894 ; n33894_not
g62856 not n16794 ; n16794_not
g62857 not n28944 ; n28944_not
g62858 not n18468 ; n18468_not
g62859 not n18459 ; n18459_not
g62860 not n45837 ; n45837_not
g62861 not n14958 ; n14958_not
g62862 not n41958 ; n41958_not
g62863 not n42768 ; n42768_not
g62864 not n42777 ; n42777_not
g62865 not n41949 ; n41949_not
g62866 not n38466 ; n38466_not
g62867 not n40995 ; n40995_not
g62868 not n38457 ; n38457_not
g62869 not n28764 ; n28764_not
g62870 not n18387 ; n18387_not
g62871 not n38871 ; n38871_not
g62872 not n18675 ; n18675_not
g62873 not n38907 ; n38907_not
g62874 not n38916 ; n38916_not
g62875 not n45891 ; n45891_not
g62876 not n38925 ; n38925_not
g62877 not n28584 ; n28584_not
g62878 not n45954 ; n45954_not
g62879 not n38943 ; n38943_not
g62880 not n38961 ; n38961_not
g62881 not n28593 ; n28593_not
g62882 not n15399 ; n15399_not
g62883 not n17856 ; n17856_not
g62884 not n45972 ; n45972_not
g62885 not n28557 ; n28557_not
g62886 not n18828 ; n18828_not
g62887 not n45990 ; n45990_not
g62888 not n15588 ; n15588_not
g62889 not n19980 ; n19980_not
g62890 not n29385 ; n29385_not
g62891 not n45981 ; n45981_not
g62892 not n40698 ; n40698_not
g62893 not n18792 ; n18792_not
g62894 not n32769 ; n32769_not
g62895 not n39069 ; n39069_not
g62896 not n28566 ; n28566_not
g62897 not n15489 ; n15489_not
g62898 not n30789 ; n30789_not
g62899 not n18747 ; n18747_not
g62900 not n41994 ; n41994_not
g62901 not n38709 ; n38709_not
g62902 not n46872 ; n46872_not
g62903 not n38736 ; n38736_not
g62904 not n18558 ; n18558_not
g62905 not n28953 ; n28953_not
g62906 not n29079 ; n29079_not
g62907 not n29475 ; n29475_not
g62908 not n27909 ; n27909_not
g62909 not n38754 ; n38754_not
g62910 not n38763 ; n38763_not
g62911 not n38772 ; n38772_not
g62912 not n38781 ; n38781_not
g62913 not n28647 ; n28647_not
g62914 not n42588 ; n42588_not
g62915 not n29448 ; n29448_not
g62916 not n46827 ; n46827_not
g62917 not n18666 ; n18666_not
g62918 not n41859 ; n41859_not
g62919 not n38817 ; n38817_not
g62920 not n29088 ; n29088_not
g62921 not n18648 ; n18648_not
g62922 not n27918 ; n27918_not
g62923 not n40797 ; n40797_not
g62924 not n16677 ; n16677_not
g62925 not n46845 ; n46845_not
g62926 not n38790 ; n38790_not
g62927 not n49059 ; n49059_not
g62928 not n27387 ; n27387_not
g62929 not n47619 ; n47619_not
g62930 not n44478 ; n44478_not
g62931 not n25488 ; n25488_not
g62932 not n25749 ; n25749_not
g62933 not n37269 ; n37269_not
g62934 not n25884 ; n25884_not
g62935 not n12798 ; n12798_not
g62936 not n43389 ; n43389_not
g62937 not n49068 ; n49068_not
g62938 not n25956 ; n25956_not
g62939 not n48465 ; n48465_not
g62940 not n47592 ; n47592_not
g62941 not n17577 ; n17577_not
g62942 not n25965 ; n25965_not
g62943 not n29862 ; n29862_not
g62944 not n26982 ; n26982_not
g62945 not n24687 ; n24687_not
g62946 not n36936 ; n36936_not
g62947 not n48654 ; n48654_not
g62948 not n34686 ; n34686_not
g62949 not n48159 ; n48159_not
g62950 not n13896 ; n13896_not
g62951 not n35478 ; n35478_not
g62952 not n35469 ; n35469_not
g62953 not n47673 ; n47673_not
g62954 not n36927 ; n36927_not
g62955 not n36738 ; n36738_not
g62956 not n27369 ; n27369_not
g62957 not n24993 ; n24993_not
g62958 not n27378 ; n27378_not
g62959 not n47664 ; n47664_not
g62960 not n26559 ; n26559_not
g62961 not n43956 ; n43956_not
g62962 not n34884 ; n34884_not
g62963 not n47547 ; n47547_not
g62964 not n47538 ; n47538_not
g62965 not n26676 ; n26676_not
g62966 not n43749 ; n43749_not
g62967 not n27459 ; n27459_not
g62968 not n26496 ; n26496_not
g62969 not n36828 ; n36828_not
g62970 not n24786 ; n24786_not
g62971 not n34569 ; n34569_not
g62972 not n11898 ; n11898_not
g62973 not n24957 ; n24957_not
g62974 not n24948 ; n24948_not
g62975 not n47970 ; n47970_not
g62976 not n43938 ; n43938_not
g62977 not n26838 ; n26838_not
g62978 not n35739 ; n35739_not
g62979 not n35748 ; n35748_not
g62980 not n26928 ; n26928_not
g62981 not n24939 ; n24939_not
g62982 not n47574 ; n47574_not
g62983 not n37296 ; n37296_not
g62984 not n12789 ; n12789_not
g62985 not n26919 ; n26919_not
g62986 not n35397 ; n35397_not
g62987 not n36882 ; n36882_not
g62988 not n25686 ; n25686_not
g62989 not n36639 ; n36639_not
g62990 not n36864 ; n36864_not
g62991 not n27099 ; n27099_not
g62992 not n34587 ; n34587_not
g62993 not n48807 ; n48807_not
g62994 not n36396 ; n36396_not
g62995 not n27198 ; n27198_not
g62996 not n25866 ; n25866_not
g62997 not n23697 ; n23697_not
g62998 not n23886 ; n23886_not
g62999 not n23688 ; n23688_not
g63000 not n47772 ; n47772_not
g63001 not n23679 ; n23679_not
g63002 not n23895 ; n23895_not
g63003 not n31977 ; n31977_not
g63004 not n36099 ; n36099_not
g63005 not n25875 ; n25875_not
g63006 not n34866 ; n34866_not
g63007 not n43587 ; n43587_not
g63008 not n48555 ; n48555_not
g63009 not n34938 ; n34938_not
g63010 not n34389 ; n34389_not
g63011 not n47763 ; n47763_not
g63012 not n43596 ; n43596_not
g63013 not n24597 ; n24597_not
g63014 not n37089 ; n37089_not
g63015 not n23796 ; n23796_not
g63016 not n29763 ; n29763_not
g63017 not n26964 ; n26964_not
g63018 not n48582 ; n48582_not
g63019 not n43965 ; n43965_not
g63020 not n35586 ; n35586_not
g63021 not n26955 ; n26955_not
g63022 not n44487 ; n44487_not
g63023 not n48591 ; n48591_not
g63024 not n35559 ; n35559_not
g63025 not n37098 ; n37098_not
g63026 not n26757 ; n26757_not
g63027 not n23859 ; n23859_not
g63028 not n47781 ; n47781_not
g63029 not n47817 ; n47817_not
g63030 not n43974 ; n43974_not
g63031 not n37188 ; n37188_not
g63032 not n48276 ; n48276_not
g63033 not n44496 ; n44496_not
g63034 not n36963 ; n36963_not
g63035 not n35649 ; n35649_not
g63036 not n36981 ; n36981_not
g63037 not n36954 ; n36954_not
g63038 not n37197 ; n37197_not
g63039 not n26667 ; n26667_not
g63040 not n48645 ; n48645_not
g63041 not n35658 ; n35658_not
g63042 not n13869 ; n13869_not
g63043 not n48177 ; n48177_not
g63044 not n27279 ; n27279_not
g63045 not n23499 ; n23499_not
g63046 not n29727 ; n29727_not
g63047 not n29970 ; n29970_not
g63048 not n23967 ; n23967_not
g63049 not n26973 ; n26973_not
g63050 not n44568 ; n44568_not
g63051 not n48546 ; n48546_not
g63052 not n12888 ; n12888_not
g63053 not n47844 ; n47844_not
g63054 not n48609 ; n48609_not
g63055 not n36990 ; n36990_not
g63056 not n48186 ; n48186_not
g63057 not n23589 ; n23589_not
g63058 not n48852 ; n48852_not
g63059 not n48267 ; n48267_not
g63060 not n34839 ; n34839_not
g63061 not n34659 ; n34659_not
g63062 not n25893 ; n25893_not
g63063 not n25794 ; n25794_not
g63064 not n48843 ; n48843_not
g63065 not n36486 ; n36486_not
g63066 not n36585 ; n36585_not
g63067 not n13986 ; n13986_not
g63068 not n43794 ; n43794_not
g63069 not n25569 ; n25569_not
g63070 not n34758 ; n34758_not
g63071 not n29934 ; n29934_not
g63072 not n36792 ; n36792_not
g63073 not n44199 ; n44199_not
g63074 not n35865 ; n35865_not
g63075 not n22896 ; n22896_not
g63076 not n35829 ; n35829_not
g63077 not n26478 ; n26478_not
g63078 not n43479 ; n43479_not
g63079 not n29808 ; n29808_not
g63080 not n22887 ; n22887_not
g63081 not n34965 ; n34965_not
g63082 not n43677 ; n43677_not
g63083 not n37467 ; n37467_not
g63084 not n26694 ; n26694_not
g63085 not n26874 ; n26874_not
g63086 not n34983 ; n34983_not
g63087 not n13995 ; n13995_not
g63088 not n35973 ; n35973_not
g63089 not n47457 ; n47457_not
g63090 not n25578 ; n25578_not
g63091 not n35298 ; n35298_not
g63092 not n43848 ; n43848_not
g63093 not n24795 ; n24795_not
g63094 not n24885 ; n24885_not
g63095 not n47466 ; n47466_not
g63096 not n26883 ; n26883_not
g63097 not n31959 ; n31959_not
g63098 not n37494 ; n37494_not
g63099 not n35964 ; n35964_not
g63100 not n36297 ; n36297_not
g63101 not n10899 ; n10899_not
g63102 not n26487 ; n26487_not
g63103 not n43875 ; n43875_not
g63104 not n26793 ; n26793_not
g63105 not n36378 ; n36378_not
g63106 not n27567 ; n27567_not
g63107 not n26199 ; n26199_not
g63108 not n48357 ; n48357_not
g63109 not n35289 ; n35289_not
g63110 not n29880 ; n29880_not
g63111 not n31869 ; n31869_not
g63112 not n43857 ; n43857_not
g63113 not n36747 ; n36747_not
g63114 not n35982 ; n35982_not
g63115 not n25497 ; n25497_not
g63116 not n12699 ; n12699_not
g63117 not n47493 ; n47493_not
g63118 not n42597 ; n42597_not
g63119 not n34992 ; n34992_not
g63120 not n26397 ; n26397_not
g63121 not n25596 ; n25596_not
g63122 not n36648 ; n36648_not
g63123 not n47385 ; n47385_not
g63124 not n23994 ; n23994_not
g63125 not n24894 ; n24894_not
g63126 not n36369 ; n36369_not
g63127 not n18856 ; n18856_not
g63128 not n36955 ; n36955_not
g63129 not n39277 ; n39277_not
g63130 not n17857 ; n17857_not
g63131 not n19909 ; n19909_not
g63132 not n31888 ; n31888_not
g63133 not n26749 ; n26749_not
g63134 not n44398 ; n44398_not
g63135 not n23959 ; n23959_not
g63136 not n36883 ; n36883_not
g63137 not n28495 ; n28495_not
g63138 not n18874 ; n18874_not
g63139 not n27928 ; n27928_not
g63140 not n29791 ; n29791_not
g63141 not n18865 ; n18865_not
g63142 not n14995 ; n14995_not
g63143 not n38575 ; n38575_not
g63144 not n35947 ; n35947_not
g63145 not n25777 ; n25777_not
g63146 not n47890 ; n47890_not
g63147 not n48736 ; n48736_not
g63148 not n29395 ; n29395_not
g63149 not n36964 ; n36964_not
g63150 not n39088 ; n39088_not
g63151 not n29980 ; n29980_not
g63152 not n16777 ; n16777_not
g63153 not n36685 ; n36685_not
g63154 not n29188 ; n29188_not
g63155 not n42697 ; n42697_not
g63156 not n48088 ; n48088_not
g63157 not n18388 ; n18388_not
g63158 not n46675 ; n46675_not
g63159 not n30979 ; n30979_not
g63160 not n39196 ; n39196_not
g63161 not n19477 ; n19477_not
g63162 not n44569 ; n44569_not
g63163 not n48871 ; n48871_not
g63164 not n23878 ; n23878_not
g63165 not n38485 ; n38485_not
g63166 not n23869 ; n23869_not
g63167 not n38467 ; n38467_not
g63168 not n15589 ; n15589_not
g63169 not n34867 ; n34867_not
g63170 not n36559 ; n36559_not
g63171 not n31897 ; n31897_not
g63172 not n19963 ; n19963_not
g63173 not n47809 ; n47809_not
g63174 not n45991 ; n45991_not
g63175 not n26569 ; n26569_not
g63176 not n35893 ; n35893_not
g63177 not n35596 ; n35596_not
g63178 not n15769 ; n15769_not
g63179 not n29377 ; n29377_not
g63180 not n38683 ; n38683_not
g63181 not n31699 ; n31699_not
g63182 not n48592 ; n48592_not
g63183 not n31879 ; n31879_not
g63184 not n18748 ; n18748_not
g63185 not n30799 ; n30799_not
g63186 not n28567 ; n28567_not
g63187 not n35587 ; n35587_not
g63188 not n30988 ; n30988_not
g63189 not n23788 ; n23788_not
g63190 not n40987 ; n40987_not
g63191 not n48187 ; n48187_not
g63192 not n36991 ; n36991_not
g63193 not n38548 ; n38548_not
g63194 not n48079 ; n48079_not
g63195 not n29836 ; n29836_not
g63196 not n35875 ; n35875_not
g63197 not n19990 ; n19990_not
g63198 not n46927 ; n46927_not
g63199 not n26992 ; n26992_not
g63200 not n41797 ; n41797_not
g63201 not n14968 ; n14968_not
g63202 not n35884 ; n35884_not
g63203 not n13699 ; n13699_not
g63204 not n36577 ; n36577_not
g63205 not n34957 ; n34957_not
g63206 not n43867 ; n43867_not
g63207 not n42499 ; n42499_not
g63208 not n23896 ; n23896_not
g63209 not n19936 ; n19936_not
g63210 not n38494 ; n38494_not
g63211 not n29368 ; n29368_not
g63212 not n28576 ; n28576_not
g63213 not n16858 ; n16858_not
g63214 not n19972 ; n19972_not
g63215 not n42769 ; n42769_not
g63216 not n38656 ; n38656_not
g63217 not n36865 ; n36865_not
g63218 not n43498 ; n43498_not
g63219 not n25687 ; n25687_not
g63220 not n34498 ; n34498_not
g63221 not n38782 ; n38782_not
g63222 not n27964 ; n27964_not
g63223 not n38818 ; n38818_not
g63224 not n33787 ; n33787_not
g63225 not n38827 ; n38827_not
g63226 not n40789 ; n40789_not
g63227 not n28675 ; n28675_not
g63228 not n12997 ; n12997_not
g63229 not n35767 ; n35767_not
g63230 not n38845 ; n38845_not
g63231 not n39637 ; n39637_not
g63232 not n39394 ; n39394_not
g63233 not n38980 ; n38980_not
g63234 not n41986 ; n41986_not
g63235 not n46747 ; n46747_not
g63236 not n47926 ; n47926_not
g63237 not n18685 ; n18685_not
g63238 not n18676 ; n18676_not
g63239 not n16597 ; n16597_not
g63240 not n43399 ; n43399_not
g63241 not n18577 ; n18577_not
g63242 not n35758 ; n35758_not
g63243 not n18955 ; n18955_not
g63244 not n35749 ; n35749_not
g63245 not n38962 ; n38962_not
g63246 not n28459 ; n28459_not
g63247 not n40897 ; n40897_not
g63248 not n18586 ; n18586_not
g63249 not n35776 ; n35776_not
g63250 not n18937 ; n18937_not
g63251 not n38926 ; n38926_not
g63252 not n38890 ; n38890_not
g63253 not n39349 ; n39349_not
g63254 not n28486 ; n28486_not
g63255 not n41779 ; n41779_not
g63256 not n28639 ; n28639_not
g63257 not n18658 ; n18658_not
g63258 not n35794 ; n35794_not
g63259 not n47962 ; n47962_not
g63260 not n38908 ; n38908_not
g63261 not n39367 ; n39367_not
g63262 not n45946 ; n45946_not
g63263 not n38917 ; n38917_not
g63264 not n19855 ; n19855_not
g63265 not n38791 ; n38791_not
g63266 not n29917 ; n29917_not
g63267 not n39646 ; n39646_not
g63268 not n46819 ; n46819_not
g63269 not n42598 ; n42598_not
g63270 not n35992 ; n35992_not
g63271 not n38863 ; n38863_not
g63272 not n38737 ; n38737_not
g63273 not n45199 ; n45199_not
g63274 not n48781 ; n48781_not
g63275 not n43948 ; n43948_not
g63276 not n38872 ; n38872_not
g63277 not n28648 ; n28648_not
g63278 not n19864 ; n19864_not
g63279 not n38881 ; n38881_not
g63280 not n16687 ; n16687_not
g63281 not n35668 ; n35668_not
g63282 not n23968 ; n23968_not
g63283 not n23977 ; n23977_not
g63284 not n45964 ; n45964_not
g63285 not n39475 ; n39475_not
g63286 not n33697 ; n33697_not
g63287 not n29782 ; n29782_not
g63288 not n19954 ; n19954_not
g63289 not n45838 ; n45838_not
g63290 not n26677 ; n26677_not
g63291 not n34876 ; n34876_not
g63292 not n43894 ; n43894_not
g63293 not n39907 ; n39907_not
g63294 not n38692 ; n38692_not
g63295 not n41887 ; n41887_not
g63296 not n16498 ; n16498_not
g63297 not n40888 ; n40888_not
g63298 not n35866 ; n35866_not
g63299 not n18739 ; n18739_not
g63300 not n39484 ; n39484_not
g63301 not n25759 ; n25759_not
g63302 not n46891 ; n46891_not
g63303 not n41959 ; n41959_not
g63304 not n19882 ; n19882_not
g63305 not n29179 ; n29179_not
g63306 not n38584 ; n38584_not
g63307 not n35938 ; n35938_not
g63308 not n35956 ; n35956_not
g63309 not n16786 ; n16786_not
g63310 not n36676 ; n36676_not
g63311 not n18883 ; n18883_not
g63312 not n45856 ; n45856_not
g63313 not n34489 ; n34489_not
g63314 not n47917 ; n47917_not
g63315 not n46864 ; n46864_not
g63316 not n25678 ; n25678_not
g63317 not n45865 ; n45865_not
g63318 not n38755 ; n38755_not
g63319 not n48808 ; n48808_not
g63320 not n15679 ; n15679_not
g63321 not n25696 ; n25696_not
g63322 not n38773 ; n38773_not
g63323 not n26686 ; n26686_not
g63324 not n28693 ; n28693_not
g63325 not n18487 ; n18487_not
g63326 not n48817 ; n48817_not
g63327 not n46765 ; n46765_not
g63328 not n16759 ; n16759_not
g63329 not n34588 ; n34588_not
g63330 not n35965 ; n35965_not
g63331 not n36793 ; n36793_not
g63332 not n29773 ; n29773_not
g63333 not n35857 ; n35857_not
g63334 not n48835 ; n48835_not
g63335 not n23995 ; n23995_not
g63336 not n18496 ; n18496_not
g63337 not n38728 ; n38728_not
g63338 not n36568 ; n36568_not
g63339 not n47908 ; n47908_not
g63340 not n38953 ; n38953_not
g63341 not n26929 ; n26929_not
g63342 not n37459 ; n37459_not
g63343 not n38665 ; n38665_not
g63344 not n15778 ; n15778_not
g63345 not n29287 ; n29287_not
g63346 not n47296 ; n47296_not
g63347 not n37990 ; n37990_not
g63348 not n21997 ; n21997_not
g63349 not n37288 ; n37288_not
g63350 not n48457 ; n48457_not
g63351 not n33598 ; n33598_not
g63352 not n41599 ; n41599_not
g63353 not n32896 ; n32896_not
g63354 not n29845 ; n29845_not
g63355 not n38449 ; n38449_not
g63356 not n15796 ; n15796_not
g63357 not n19459 ; n19459_not
g63358 not n15958 ; n15958_not
g63359 not n35398 ; n35398_not
g63360 not n37297 ; n37297_not
g63361 not n19369 ; n19369_not
g63362 not n37981 ; n37981_not
g63363 not n19558 ; n19558_not
g63364 not n37819 ; n37819_not
g63365 not n25966 ; n25966_not
g63366 not n29629 ; n29629_not
g63367 not n19729 ; n19729_not
g63368 not n17497 ; n17497_not
g63369 not n17578 ; n17578_not
g63370 not n38089 ; n38089_not
g63371 not n30889 ; n30889_not
g63372 not n19567 ; n19567_not
g63373 not n34687 ; n34687_not
g63374 not n19378 ; n19378_not
g63375 not n27649 ; n27649_not
g63376 not n29926 ; n29926_not
g63377 not n37648 ; n37648_not
g63378 not n21898 ; n21898_not
g63379 not n27694 ; n27694_not
g63380 not n21979 ; n21979_not
g63381 not n27757 ; n27757_not
g63382 not n29728 ; n29728_not
g63383 not n25957 ; n25957_not
g63384 not n37468 ; n37468_not
g63385 not n19387 ; n19387_not
g63386 not n29908 ; n29908_not
g63387 not n32878 ; n32878_not
g63388 not n27784 ; n27784_not
g63389 not n34696 ; n34696_not
g63390 not n29737 ; n29737_not
g63391 not n39943 ; n39943_not
g63392 not n15895 ; n15895_not
g63393 not n39763 ; n39763_not
g63394 not n28972 ; n28972_not
g63395 not n39952 ; n39952_not
g63396 not n28882 ; n28882_not
g63397 not n46387 ; n46387_not
g63398 not n22996 ; n22996_not
g63399 not n39853 ; n39853_not
g63400 not n29458 ; n29458_not
g63401 not n46288 ; n46288_not
g63402 not n25939 ; n25939_not
g63403 not n17587 ; n17587_not
g63404 not n22879 ; n22879_not
g63405 not n37873 ; n37873_not
g63406 not n19684 ; n19684_not
g63407 not n27469 ; n27469_not
g63408 not n30898 ; n30898_not
g63409 not n29647 ; n29647_not
g63410 not n22969 ; n22969_not
g63411 not n17596 ; n17596_not
g63412 not n37378 ; n37378_not
g63413 not n37369 ; n37369_not
g63414 not n37855 ; n37855_not
g63415 not n17695 ; n17695_not
g63416 not n27478 ; n27478_not
g63417 not n27685 ; n27685_not
g63418 not n29278 ; n29278_not
g63419 not n39916 ; n39916_not
g63420 not n47278 ; n47278_not
g63421 not n37936 ; n37936_not
g63422 not n27676 ; n27676_not
g63423 not n15877 ; n15877_not
g63424 not n14698 ; n14698_not
g63425 not n15949 ; n15949_not
g63426 not n37945 ; n37945_not
g63427 not n47557 ; n47557_not
g63428 not n17785 ; n17785_not
g63429 not n39817 ; n39817_not
g63430 not n17794 ; n17794_not
g63431 not n17569 ; n17569_not
g63432 not n37954 ; n37954_not
g63433 not n45298 ; n45298_not
g63434 not n36397 ; n36397_not
g63435 not n19549 ; n19549_not
g63436 not n39844 ; n39844_not
g63437 not n39826 ; n39826_not
g63438 not n16948 ; n16948_not
g63439 not n13969 ; n13969_not
g63440 not n22888 ; n22888_not
g63441 not n43768 ; n43768_not
g63442 not n39835 ; n39835_not
g63443 not n37684 ; n37684_not
g63444 not n29638 ; n29638_not
g63445 not n37927 ; n37927_not
g63446 not n36199 ; n36199_not
g63447 not n15787 ; n15787_not
g63448 not n32599 ; n32599_not
g63449 not n37387 ; n37387_not
g63450 not n27856 ; n27856_not
g63451 not n47359 ; n47359_not
g63452 not n27586 ; n27586_not
g63453 not n34399 ; n34399_not
g63454 not n39466 ; n39466_not
g63455 not n48574 ; n48574_not
g63456 not n34849 ; n34849_not
g63457 not n31789 ; n31789_not
g63458 not n24589 ; n24589_not
g63459 not n29755 ; n29755_not
g63460 not n37774 ; n37774_not
g63461 not n32869 ; n32869_not
g63462 not n14878 ; n14878_not
g63463 not n33949 ; n33949_not
g63464 not n47755 ; n47755_not
g63465 not n48538 ; n48538_not
g63466 not n36496 ; n36496_not
g63467 not n19756 ; n19756_not
g63468 not n48349 ; n48349_not
g63469 not n12898 ; n12898_not
g63470 not n47764 ; n47764_not
g63471 not n28099 ; n28099_not
g63472 not n14869 ; n14869_not
g63473 not n28819 ; n28819_not
g63474 not n15697 ; n15697_not
g63475 not n38386 ; n38386_not
g63476 not n38395 ; n38395_not
g63477 not n39934 ; n39934_not
g63478 not n29818 ; n29818_not
g63479 not n18199 ; n18199_not
g63480 not n48880 ; n48880_not
g63481 not n46963 ; n46963_not
g63482 not n46468 ; n46468_not
g63483 not n22789 ; n22789_not
g63484 not n32689 ; n32689_not
g63485 not n26596 ; n26596_not
g63486 not n29665 ; n29665_not
g63487 not n36298 ; n36298_not
g63488 not n19576 ; n19576_not
g63489 not n29962 ; n29962_not
g63490 not n41869 ; n41869_not
g63491 not n29683 ; n29683_not
g63492 not n13798 ; n13798_not
g63493 not n39592 ; n39592_not
g63494 not n37549 ; n37549_not
g63495 not n38368 ; n38368_not
g63496 not n17398 ; n17398_not
g63497 not n26758 ; n26758_not
g63498 not n14896 ; n14896_not
g63499 not n46369 ; n46369_not
g63500 not n35299 ; n35299_not
g63501 not n38377 ; n38377_not
g63502 not n39583 ; n39583_not
g63503 not n33985 ; n33985_not
g63504 not n24679 ; n24679_not
g63505 not n17884 ; n17884_not
g63506 not n47719 ; n47719_not
g63507 not n36469 ; n36469_not
g63508 not n17479 ; n17479_not
g63509 not n38188 ; n38188_not
g63510 not n37792 ; n37792_not
g63511 not n29575 ; n29575_not
g63512 not n13879 ; n13879_not
g63513 not n29674 ; n29674_not
g63514 not n47728 ; n47728_not
g63515 not n36478 ; n36478_not
g63516 not n48475 ; n48475_not
g63517 not n37666 ; n37666_not
g63518 not n15985 ; n15985_not
g63519 not n28945 ; n28945_not
g63520 not n33994 ; n33994_not
g63521 not n11998 ; n11998_not
g63522 not n39727 ; n39727_not
g63523 not n17938 ; n17938_not
g63524 not n39718 ; n39718_not
g63525 not n47692 ; n47692_not
g63526 not n14779 ; n14779_not
g63527 not n19279 ; n19279_not
g63528 not n29557 ; n29557_not
g63529 not n37585 ; n37585_not
g63530 not n39655 ; n39655_not
g63531 not n17974 ; n17974_not
g63532 not n26785 ; n26785_not
g63533 not n41689 ; n41689_not
g63534 not n43786 ; n43786_not
g63535 not n19693 ; n19693_not
g63536 not n42895 ; n42895_not
g63537 not n28927 ; n28927_not
g63538 not n34669 ; n34669_not
g63539 not n48277 ; n48277_not
g63540 not n37747 ; n37747_not
g63541 not n22699 ; n22699_not
g63542 not n33967 ; n33967_not
g63543 not n28909 ; n28909_not
g63544 not n45658 ; n45658_not
g63545 not n45667 ; n45667_not
g63546 not n29746 ; n29746_not
g63547 not n37594 ; n37594_not
g63548 not n39736 ; n39736_not
g63549 not n48268 ; n48268_not
g63550 not n34796 ; n34796_not
g63551 not n39755 ; n39755_not
g63552 not n39944 ; n39944_not
g63553 not n17849 ; n17849_not
g63554 not n19892 ; n19892_not
g63555 not n24878 ; n24878_not
g63556 not n27947 ; n27947_not
g63557 not n36299 ; n36299_not
g63558 not n29288 ; n29288_not
g63559 not n38855 ; n38855_not
g63560 not n44669 ; n44669_not
g63561 not n19649 ; n19649_not
g63562 not n34679 ; n34679_not
g63563 not n24869 ; n24869_not
g63564 not n26858 ; n26858_not
g63565 not n38963 ; n38963_not
g63566 not n28559 ; n28559_not
g63567 not n39197 ; n39197_not
g63568 not n19676 ; n19676_not
g63569 not n24698 ; n24698_not
g63570 not n19595 ; n19595_not
g63571 not n46397 ; n46397_not
g63572 not n39962 ; n39962_not
g63573 not n28955 ; n28955_not
g63574 not n36668 ; n36668_not
g63575 not n15797 ; n15797_not
g63576 not n48089 ; n48089_not
g63577 not n18866 ; n18866_not
g63578 not n27956 ; n27956_not
g63579 not n38891 ; n38891_not
g63580 not n39980 ; n39980_not
g63581 not n18857 ; n18857_not
g63582 not n27938 ; n27938_not
g63583 not n36695 ; n36695_not
g63584 not n48629 ; n48629_not
g63585 not n19748 ; n19748_not
g63586 not n29189 ; n29189_not
g63587 not n36587 ; n36587_not
g63588 not n28469 ; n28469_not
g63589 not n36596 ; n36596_not
g63590 not n19298 ; n19298_not
g63591 not n26939 ; n26939_not
g63592 not n32699 ; n32699_not
g63593 not n48278 ; n48278_not
g63594 not n19739 ; n19739_not
g63595 not n48494 ; n48494_not
g63596 not n18983 ; n18983_not
g63597 not n48287 ; n48287_not
g63598 not n34877 ; n34877_not
g63599 not n15986 ; n15986_not
g63600 not n34688 ; n34688_not
g63601 not n18974 ; n18974_not
g63602 not n39458 ; n39458_not
g63603 not n38765 ; n38765_not
g63604 not n24986 ; n24986_not
g63605 not n26957 ; n26957_not
g63606 not n39566 ; n39566_not
g63607 not n38837 ; n38837_not
g63608 not n27983 ; n27983_not
g63609 not n19775 ; n19775_not
g63610 not n39557 ; n39557_not
g63611 not n39548 ; n39548_not
g63612 not n42887 ; n42887_not
g63613 not n34859 ; n34859_not
g63614 not n39593 ; n39593_not
g63615 not n19784 ; n19784_not
g63616 not n26948 ; n26948_not
g63617 not n34868 ; n34868_not
g63618 not n48197 ; n48197_not
g63619 not n36578 ; n36578_not
g63620 not n48557 ; n48557_not
g63621 not n19766 ; n19766_not
g63622 not n28397 ; n28397_not
g63623 not n24599 ; n24599_not
g63624 not n26849 ; n26849_not
g63625 not n12899 ; n12899_not
g63626 not n43796 ; n43796_not
g63627 not n19793 ; n19793_not
g63628 not n36497 ; n36497_not
g63629 not n38387 ; n38387_not
g63630 not n36389 ; n36389_not
g63631 not n26894 ; n26894_not
g63632 not n39854 ; n39854_not
g63633 not n28478 ; n28478_not
g63634 not n46748 ; n46748_not
g63635 not n16958 ; n16958_not
g63636 not n46298 ; n46298_not
g63637 not n26984 ; n26984_not
g63638 not n39890 ; n39890_not
g63639 not n46649 ; n46649_not
g63640 not n39737 ; n39737_not
g63641 not n19865 ; n19865_not
g63642 not n29855 ; n29855_not
g63643 not n43499 ; n43499_not
g63644 not n28199 ; n28199_not
g63645 not n46487 ; n46487_not
g63646 not n19874 ; n19874_not
g63647 not n39926 ; n39926_not
g63648 not n39935 ; n39935_not
g63649 not n39764 ; n39764_not
g63650 not n34886 ; n34886_not
g63651 not n18965 ; n18965_not
g63652 not n12989 ; n12989_not
g63653 not n34589 ; n34589_not
g63654 not n19829 ; n19829_not
g63655 not n24968 ; n24968_not
g63656 not n48449 ; n48449_not
g63657 not n18956 ; n18956_not
g63658 not n24779 ; n24779_not
g63659 not n36398 ; n36398_not
g63660 not n39791 ; n39791_not
g63661 not n39638 ; n39638_not
g63662 not n43778 ; n43778_not
g63663 not n39386 ; n39386_not
g63664 not n30998 ; n30998_not
g63665 not n19469 ; n19469_not
g63666 not n19478 ; n19478_not
g63667 not n18947 ; n18947_not
g63668 not n24977 ; n24977_not
g63669 not n28973 ; n28973_not
g63670 not n42896 ; n42896_not
g63671 not n33959 ; n33959_not
g63672 not n47738 ; n47738_not
g63673 not n17894 ; n17894_not
g63674 not n27839 ; n27839_not
g63675 not n42878 ; n42878_not
g63676 not n17867 ; n17867_not
g63677 not n28829 ; n28829_not
g63678 not n45677 ; n45677_not
g63679 not n17984 ; n17984_not
g63680 not n29558 ; n29558_not
g63681 not n40799 ; n40799_not
g63682 not n26579 ; n26579_not
g63683 not n31979 ; n31979_not
g63684 not n45686 ; n45686_not
g63685 not n32888 ; n32888_not
g63686 not n13889 ; n13889_not
g63687 not n47648 ; n47648_not
g63688 not n28847 ; n28847_not
g63689 not n17885 ; n17885_not
g63690 not n38648 ; n38648_not
g63691 not n13898 ; n13898_not
g63692 not n47099 ; n47099_not
g63693 not n33995 ; n33995_not
g63694 not n28838 ; n28838_not
g63695 not n35498 ; n35498_not
g63696 not n16967 ; n16967_not
g63697 not n29747 ; n29747_not
g63698 not n38576 ; n38576_not
g63699 not n38189 ; n38189_not
g63700 not n32879 ; n32879_not
g63701 not n14798 ; n14798_not
g63702 not n16949 ; n16949_not
g63703 not n38396 ; n38396_not
g63704 not n41888 ; n41888_not
g63705 not n42797 ; n42797_not
g63706 not n41897 ; n41897_not
g63707 not n28784 ; n28784_not
g63708 not n23789 ; n23789_not
g63709 not n46955 ; n46955_not
g63710 not n42788 ; n42788_not
g63711 not n27875 ; n27875_not
g63712 not n33887 ; n33887_not
g63713 not n39467 ; n39467_not
g63714 not n16877 ; n16877_not
g63715 not n38459 ; n38459_not
g63716 not n33878 ; n33878_not
g63717 not n38468 ; n38468_not
g63718 not n23879 ; n23879_not
g63719 not n28694 ; n28694_not
g63720 not n29774 ; n29774_not
g63721 not n38477 ; n38477_not
g63722 not n25796 ; n25796_not
g63723 not n20999 ; n20999_not
g63724 not n38297 ; n38297_not
g63725 not n25877 ; n25877_not
g63726 not n47765 ; n47765_not
g63727 not n14879 ; n14879_not
g63728 not n42779 ; n42779_not
g63729 not n46991 ; n46991_not
g63730 not n43976 ; n43976_not
g63731 not n44759 ; n44759_not
g63732 not n47774 ; n47774_not
g63733 not n14888 ; n14888_not
g63734 not n43958 ; n43958_not
g63735 not n27866 ; n27866_not
g63736 not n28991 ; n28991_not
g63737 not n38369 ; n38369_not
g63738 not n26588 ; n26588_not
g63739 not n38378 ; n38378_not
g63740 not n14897 ; n14897_not
g63741 not n16688 ; n16688_not
g63742 not n17579 ; n17579_not
g63743 not n37685 ; n37685_not
g63744 not n13997 ; n13997_not
g63745 not n28937 ; n28937_not
g63746 not n37694 ; n37694_not
g63747 not n27686 ; n27686_not
g63748 not n37739 ; n37739_not
g63749 not n29918 ; n29918_not
g63750 not n37568 ; n37568_not
g63751 not n47459 ; n47459_not
g63752 not n27497 ; n27497_not
g63753 not n28892 ; n28892_not
g63754 not n29657 ; n29657_not
g63755 not n37397 ; n37397_not
g63756 not n17669 ; n17669_not
g63757 not n27578 ; n27578_not
g63758 not n47369 ; n47369_not
g63759 not n47378 ; n47378_not
g63760 not n17399 ; n17399_not
g63761 not n22799 ; n22799_not
g63762 not n37577 ; n37577_not
g63763 not n27596 ; n27596_not
g63764 not n37586 ; n37586_not
g63765 not n47396 ; n47396_not
g63766 not n32969 ; n32969_not
g63767 not n37496 ; n37496_not
g63768 not n29963 ; n29963_not
g63769 not n37478 ; n37478_not
g63770 not n16697 ; n16697_not
g63771 not n27659 ; n27659_not
g63772 not n37658 ; n37658_not
g63773 not n27668 ; n27668_not
g63774 not n32996 ; n32996_not
g63775 not n29639 ; n29639_not
g63776 not n28874 ; n28874_not
g63777 not n37964 ; n37964_not
g63778 not n32897 ; n32897_not
g63779 not n37973 ; n37973_not
g63780 not n37982 ; n37982_not
g63781 not n25976 ; n25976_not
g63782 not n47585 ; n47585_not
g63783 not n28739 ; n28739_not
g63784 not n27389 ; n27389_not
g63785 not n42986 ; n42986_not
g63786 not n38495 ; n38495_not
g63787 not n27785 ; n27785_not
g63788 not n42968 ; n42968_not
g63789 not n25949 ; n25949_not
g63790 not n42977 ; n42977_not
g63791 not n21899 ; n21899_not
g63792 not n29891 ; n29891_not
g63793 not n47639 ; n47639_not
g63794 not n47477 ; n47477_not
g63795 not n29648 ; n29648_not
g63796 not n27488 ; n27488_not
g63797 not n37838 ; n37838_not
g63798 not n47495 ; n47495_not
g63799 not n17696 ; n17696_not
g63800 not n22979 ; n22979_not
g63801 not n37865 ; n37865_not
g63802 not n37874 ; n37874_not
g63803 not n22988 ; n22988_not
g63804 not n25994 ; n25994_not
g63805 not n37892 ; n37892_not
g63806 not n14699 ; n14699_not
g63807 not n47198 ; n47198_not
g63808 not n25985 ; n25985_not
g63809 not n17768 ; n17768_not
g63810 not n37919 ; n37919_not
g63811 not n47189 ; n47189_not
g63812 not n47954 ; n47954_not
g63813 not n39089 ; n39089_not
g63814 not n25598 ; n25598_not
g63815 not n18767 ; n18767_not
g63816 not n18587 ; n18587_not
g63817 not n40988 ; n40988_not
g63818 not n35786 ; n35786_not
g63819 not n45938 ; n45938_not
g63820 not n31988 ; n31988_not
g63821 not n27929 ; n27929_not
g63822 not n36767 ; n36767_not
g63823 not n18776 ; n18776_not
g63824 not n25697 ; n25697_not
g63825 not n19955 ; n19955_not
g63826 not n46856 ; n46856_not
g63827 not n38882 ; n38882_not
g63828 not n41987 ; n41987_not
g63829 not n40898 ; n40898_not
g63830 not n47927 ; n47927_not
g63831 not n39098 ; n39098_not
g63832 not n41996 ; n41996_not
g63833 not n36857 ; n36857_not
g63834 not n36848 ; n36848_not
g63835 not n38828 ; n38828_not
g63836 not n35867 ; n35867_not
g63837 not n43895 ; n43895_not
g63838 not n45965 ; n45965_not
g63839 not n36785 ; n36785_not
g63840 not n46766 ; n46766_not
g63841 not n16589 ; n16589_not
g63842 not n38990 ; n38990_not
g63843 not n32789 ; n32789_not
g63844 not n38909 ; n38909_not
g63845 not n25679 ; n25679_not
g63846 not n18659 ; n18659_not
g63847 not n38927 ; n38927_not
g63848 not n16598 ; n16598_not
g63849 not n46793 ; n46793_not
g63850 not n38936 ; n38936_not
g63851 not n33779 ; n33779_not
g63852 not n48737 ; n48737_not
g63853 not n36776 ; n36776_not
g63854 not n25778 ; n25778_not
g63855 not n36956 ; n36956_not
g63856 not n42698 ; n42698_not
g63857 not n28748 ; n28748_not
g63858 not n19973 ; n19973_not
g63859 not n36758 ; n36758_not
g63860 not n26669 ; n26669_not
g63861 not n36929 ; n36929_not
g63862 not n18794 ; n18794_not
g63863 not n27893 ; n27893_not
g63864 not n36938 ; n36938_not
g63865 not n23969 ; n23969_not
g63866 not n29972 ; n29972_not
g63867 not n25769 ; n25769_not
g63868 not n35678 ; n35678_not
g63869 not n39188 ; n39188_not
g63870 not n48845 ; n48845_not
g63871 not n39179 ; n39179_not
g63872 not n48863 ; n48863_not
g63873 not n38558 ; n38558_not
g63874 not n35894 ; n35894_not
g63875 not n33869 ; n33869_not
g63876 not n46919 ; n46919_not
g63877 not n27884 ; n27884_not
g63878 not n38585 ; n38585_not
g63879 not n46694 ; n46694_not
g63880 not n38594 ; n38594_not
g63881 not n29495 ; n29495_not
g63882 not n48827 ; n48827_not
g63883 not n29459 ; n29459_not
g63884 not n40997 ; n40997_not
g63885 not n18497 ; n18497_not
g63886 not n40979 ; n40979_not
g63887 not n43886 ; n43886_not
g63888 not n29387 ; n29387_not
g63889 not n48836 ; n48836_not
g63890 not n29882 ; n29882_not
g63891 not n38684 ; n38684_not
g63892 not n19982 ; n19982_not
g63893 not n16778 ; n16778_not
g63894 not n24897 ; n24897_not
g63895 not n48783 ; n48783_not
g63896 not n32988 ; n32988_not
g63897 not n43689 ; n43689_not
g63898 not n29856 ; n29856_not
g63899 not n46299 ; n46299_not
g63900 not n32979 ; n32979_not
g63901 not n15888 ; n15888_not
g63902 not n24969 ; n24969_not
g63903 not n18858 ; n18858_not
g63904 not n28884 ; n28884_not
g63905 not n19587 ; n19587_not
g63906 not n25995 ; n25995_not
g63907 not n19668 ; n19668_not
g63908 not n19497 ; n19497_not
g63909 not n16896 ; n16896_not
g63910 not n26499 ; n26499_not
g63911 not n18777 ; n18777_not
g63912 not n43869 ; n43869_not
g63913 not n34797 ; n34797_not
g63914 not n18849 ; n18849_not
g63915 not n48378 ; n48378_not
g63916 not n16995 ; n16995_not
g63917 not n35877 ; n35877_not
g63918 not n39909 ; n39909_not
g63919 not n43698 ; n43698_not
g63920 not n16797 ; n16797_not
g63921 not n28893 ; n28893_not
g63922 not n48396 ; n48396_not
g63923 not n19659 ; n19659_not
g63924 not n29874 ; n29874_not
g63925 not n15897 ; n15897_not
g63926 not n28578 ; n28578_not
g63927 not n17679 ; n17679_not
g63928 not n28938 ; n28938_not
g63929 not n17589 ; n17589_not
g63930 not n43887 ; n43887_not
g63931 not n24888 ; n24888_not
g63932 not n45984 ; n45984_not
g63933 not n17688 ; n17688_not
g63934 not n40989 ; n40989_not
g63935 not n28389 ; n28389_not
g63936 not n35787 ; n35787_not
g63937 not n18489 ; n18489_not
g63938 not n18975 ; n18975_not
g63939 not n28983 ; n28983_not
g63940 not n40998 ; n40998_not
g63941 not n17994 ; n17994_not
g63942 not n26778 ; n26778_not
g63943 not n17976 ; n17976_not
g63944 not n45678 ; n45678_not
g63945 not n17967 ; n17967_not
g63946 not n29865 ; n29865_not
g63947 not n45876 ; n45876_not
g63948 not n41979 ; n41979_not
g63949 not n45894 ; n45894_not
g63950 not n38955 ; n38955_not
g63951 not n19299 ; n19299_not
g63952 not n17958 ; n17958_not
g63953 not n15996 ; n15996_not
g63954 not n43995 ; n43995_not
g63955 not n28767 ; n28767_not
g63956 not n48864 ; n48864_not
g63957 not n25797 ; n25797_not
g63958 not n48855 ; n48855_not
g63959 not n16869 ; n16869_not
g63960 not n35598 ; n35598_not
g63961 not n43968 ; n43968_not
g63962 not n35589 ; n35589_not
g63963 not n16788 ; n16788_not
g63964 not n39738 ; n39738_not
g63965 not n41898 ; n41898_not
g63966 not n48891 ; n48891_not
g63967 not n38883 ; n38883_not
g63968 not n48873 ; n48873_not
g63969 not n18993 ; n18993_not
g63970 not n48567 ; n48567_not
g63971 not n29199 ; n29199_not
g63972 not n45696 ; n45696_not
g63973 not n46839 ; n46839_not
g63974 not n25869 ; n25869_not
g63975 not n43779 ; n43779_not
g63976 not n16599 ; n16599_not
g63977 not n39747 ; n39747_not
g63978 not n18687 ; n18687_not
g63979 not n28866 ; n28866_not
g63980 not n24996 ; n24996_not
g63981 not n18696 ; n18696_not
g63982 not n17778 ; n17778_not
g63983 not n45957 ; n45957_not
g63984 not n28965 ; n28965_not
g63985 not n18894 ; n18894_not
g63986 not n34968 ; n34968_not
g63987 not n25986 ; n25986_not
g63988 not n26688 ; n26688_not
g63989 not n17949 ; n17949_not
g63990 not n28668 ; n28668_not
g63991 not n34896 ; n34896_not
g63992 not n28839 ; n28839_not
g63993 not n18948 ; n18948_not
g63994 not n29973 ; n29973_not
g63995 not n18597 ; n18597_not
g63996 not n48486 ; n48486_not
g63997 not n17895 ; n17895_not
g63998 not n39639 ; n39639_not
g63999 not n15978 ; n15978_not
g64000 not n35985 ; n35985_not
g64001 not n34995 ; n34995_not
g64002 not n28857 ; n28857_not
g64003 not n25959 ; n25959_not
g64004 not n17859 ; n17859_not
g64005 not n25968 ; n25968_not
g64006 not n39288 ; n39288_not
g64007 not n30999 ; n30999_not
g64008 not n36678 ; n36678_not
g64009 not n19884 ; n19884_not
g64010 not n46668 ; n46668_not
g64011 not n36687 ; n36687_not
g64012 not n36696 ; n36696_not
g64013 not n26994 ; n26994_not
g64014 not n38487 ; n38487_not
g64015 not n19983 ; n19983_not
g64016 not n37668 ; n37668_not
g64017 not n39099 ; n39099_not
g64018 not n27669 ; n27669_not
g64019 not n36777 ; n36777_not
g64020 not n36786 ; n36786_not
g64021 not n19938 ; n19938_not
g64022 not n36795 ; n36795_not
g64023 not n38991 ; n38991_not
g64024 not n46785 ; n46785_not
g64025 not n33789 ; n33789_not
g64026 not n47973 ; n47973_not
g64027 not n38892 ; n38892_not
g64028 not n38874 ; n38874_not
g64029 not n38847 ; n38847_not
g64030 not n47955 ; n47955_not
g64031 not n38856 ; n38856_not
g64032 not n38748 ; n38748_not
g64033 not n38775 ; n38775_not
g64034 not n36894 ; n36894_not
g64035 not n37596 ; n37596_not
g64036 not n34689 ; n34689_not
g64037 not n48288 ; n48288_not
g64038 not n24699 ; n24699_not
g64039 not n48279 ; n48279_not
g64040 not n39729 ; n39729_not
g64041 not n39693 ; n39693_not
g64042 not n39684 ; n39684_not
g64043 not n39675 ; n39675_not
g64044 not n36498 ; n36498_not
g64045 not n39648 ; n39648_not
g64046 not n43599 ; n43599_not
g64047 not n39585 ; n39585_not
g64048 not n19767 ; n19767_not
g64049 not n26949 ; n26949_not
g64050 not n29829 ; n29829_not
g64051 not n15699 ; n15699_not
g64052 not n26967 ; n26967_not
g64053 not n46587 ; n46587_not
g64054 not n36588 ; n36588_not
g64055 not n26976 ; n26976_not
g64056 not n39495 ; n39495_not
g64057 not n39486 ; n39486_not
g64058 not n39477 ; n39477_not
g64059 not n39468 ; n39468_not
g64060 not n44499 ; n44499_not
g64061 not n19839 ; n19839_not
g64062 not n19848 ; n19848_not
g64063 not n37488 ; n37488_not
g64064 not n36669 ; n36669_not
g64065 not n39297 ; n39297_not
g64066 not n13989 ; n13989_not
g64067 not n29568 ; n29568_not
g64068 not n14799 ; n14799_not
g64069 not n39864 ; n39864_not
g64070 not n38766 ; n38766_not
g64071 not n33996 ; n33996_not
g64072 not n37398 ; n37398_not
g64073 not n47676 ; n47676_not
g64074 not n29586 ; n29586_not
g64075 not n13899 ; n13899_not
g64076 not n29694 ; n29694_not
g64077 not n27399 ; n27399_not
g64078 not n47595 ; n47595_not
g64079 not n37749 ; n37749_not
g64080 not n37992 ; n37992_not
g64081 not n37974 ; n37974_not
g64082 not n37299 ; n37299_not
g64083 not n37965 ; n37965_not
g64084 not n21999 ; n21999_not
g64085 not n36975 ; n36975_not
g64086 not n47199 ; n47199_not
g64087 not n22998 ; n22998_not
g64088 not n37893 ; n37893_not
g64089 not n37857 ; n37857_not
g64090 not n37884 ; n37884_not
g64091 not n37875 ; n37875_not
g64092 not n37866 ; n37866_not
g64093 not n36966 ; n36966_not
g64094 not n37848 ; n37848_not
g64095 not n38739 ; n38739_not
g64096 not n37695 ; n37695_not
g64097 not n38568 ; n38568_not
g64098 not n38667 ; n38667_not
g64099 not n38694 ; n38694_not
g64100 not n38676 ; n38676_not
g64101 not n47892 ; n47892_not
g64102 not n47874 ; n47874_not
g64103 not n29487 ; n29487_not
g64104 not n36948 ; n36948_not
g64105 not n14997 ; n14997_not
g64106 not n47865 ; n47865_not
g64107 not n47856 ; n47856_not
g64108 not n33798 ; n33798_not
g64109 not n36984 ; n36984_not
g64110 not n47829 ; n47829_not
g64111 not n38469 ; n38469_not
g64112 not n46947 ; n46947_not
g64113 not n23799 ; n23799_not
g64114 not n42789 ; n42789_not
g64115 not n47793 ; n47793_not
g64116 not n22899 ; n22899_not
g64117 not n33897 ; n33897_not
g64118 not n42798 ; n42798_not
g64119 not n38379 ; n38379_not
g64120 not n27858 ; n27858_not
g64121 not n46983 ; n46983_not
g64122 not n27849 ; n27849_not
g64123 not n37758 ; n37758_not
g64124 not n47469 ; n47469_not
g64125 not n29955 ; n29955_not
g64126 not n37767 ; n37767_not
g64127 not n15789 ; n15789_not
g64128 not n37578 ; n37578_not
g64129 not n39954 ; n39954_not
g64130 not n24798 ; n24798_not
g64131 not n27579 ; n27579_not
g64132 not n24789 ; n24789_not
g64133 not n39990 ; n39990_not
g64134 not n46497 ; n46497_not
g64135 not n39846 ; n39846_not
g64136 not n29298 ; n29298_not
g64137 not n39918 ; n39918_not
g64138 not n39981 ; n39981_not
g64139 not n26877 ; n26877_not
g64140 not n39756 ; n39756_not
g64141 not n39891 ; n39891_not
g64142 not n39792 ; n39792_not
g64143 not n39936 ; n39936_not
g64144 not n47389 ; n47389_not
g64145 not n38992 ; n38992_not
g64146 not n38956 ; n38956_not
g64147 not n16699 ; n16699_not
g64148 not n34987 ; n34987_not
g64149 not n37984 ; n37984_not
g64150 not n45958 ; n45958_not
g64151 not n45949 ; n45949_not
g64152 not n46768 ; n46768_not
g64153 not n37975 ; n37975_not
g64154 not n39883 ; n39883_not
g64155 not n37678 ; n37678_not
g64156 not n47947 ; n47947_not
g64157 not n17779 ; n17779_not
g64158 not n34978 ; n34978_not
g64159 not n29929 ; n29929_not
g64160 not n44977 ; n44977_not
g64161 not n38866 ; n38866_not
g64162 not n41998 ; n41998_not
g64163 not n18598 ; n18598_not
g64164 not n47956 ; n47956_not
g64165 not n15898 ; n15898_not
g64166 not n38875 ; n38875_not
g64167 not n35779 ; n35779_not
g64168 not n38884 ; n38884_not
g64169 not n35788 ; n35788_not
g64170 not n47587 ; n47587_not
g64171 not n42997 ; n42997_not
g64172 not n33799 ; n33799_not
g64173 not n25969 ; n25969_not
g64174 not n47983 ; n47983_not
g64175 not n46678 ; n46678_not
g64176 not n39199 ; n39199_not
g64177 not n26986 ; n26986_not
g64178 not n38578 ; n38578_not
g64179 not n27949 ; n27949_not
g64180 not n17788 ; n17788_not
g64181 not n18877 ; n18877_not
g64182 not n38497 ; n38497_not
g64183 not n37948 ; n37948_not
g64184 not n18886 ; n18886_not
g64185 not n35869 ; n35869_not
g64186 not n19867 ; n19867_not
g64187 not n39865 ; n39865_not
g64188 not n39847 ; n39847_not
g64189 not n19858 ; n19858_not
g64190 not n29785 ; n29785_not
g64191 not n19975 ; n19975_not
g64192 not n37957 ; n37957_not
g64193 not n26797 ; n26797_not
g64194 not n35887 ; n35887_not
g64195 not n18796 ; n18796_not
g64196 not n27697 ; n27697_not
g64197 not n28489 ; n28489_not
g64198 not n29794 ; n29794_not
g64199 not n19966 ; n19966_not
g64200 not n32989 ; n32989_not
g64201 not n19948 ; n19948_not
g64202 not n46687 ; n46687_not
g64203 not n35896 ; n35896_not
g64204 not n45994 ; n45994_not
g64205 not n17797 ; n17797_not
g64206 not n19939 ; n19939_not
g64207 not n48892 ; n48892_not
g64208 not n37795 ; n37795_not
g64209 not n47785 ; n47785_not
g64210 not n33898 ; n33898_not
g64211 not n47686 ; n47686_not
g64212 not n39955 ; n39955_not
g64213 not n16879 ; n16879_not
g64214 not n38947 ; n38947_not
g64215 not n48883 ; n48883_not
g64216 not n24799 ; n24799_not
g64217 not n29686 ; n29686_not
g64218 not n29659 ; n29659_not
g64219 not n28984 ; n28984_not
g64220 not n29767 ; n29767_not
g64221 not n17599 ; n17599_not
g64222 not n46939 ; n46939_not
g64223 not n39667 ; n39667_not
g64224 not n33988 ; n33988_not
g64225 not n29578 ; n29578_not
g64226 not n33979 ; n33979_not
g64227 not n17959 ; n17959_not
g64228 not n25888 ; n25888_not
g64229 not n29569 ; n29569_not
g64230 not n17977 ; n17977_not
g64231 not n15799 ; n15799_not
g64232 not n17968 ; n17968_not
g64233 not n47758 ; n47758_not
g64234 not n29695 ; n29695_not
g64235 not n38299 ; n38299_not
g64236 not n43987 ; n43987_not
g64237 not n47767 ; n47767_not
g64238 not n47776 ; n47776_not
g64239 not n46975 ; n46975_not
g64240 not n14899 ; n14899_not
g64241 not n38596 ; n38596_not
g64242 not n37696 ; n37696_not
g64243 not n46876 ; n46876_not
g64244 not n39892 ; n39892_not
g64245 not n19399 ; n19399_not
g64246 not n27796 ; n27796_not
g64247 not n26599 ; n26599_not
g64248 not n36895 ; n36895_not
g64249 not n37687 ; n37687_not
g64250 not n25699 ; n25699_not
g64251 not n38677 ; n38677_not
g64252 not n27589 ; n27589_not
g64253 not n42979 ; n42979_not
g64254 not n38785 ; n38785_not
g64255 not n28678 ; n28678_not
g64256 not n36877 ; n36877_not
g64257 not n47938 ; n47938_not
g64258 not n29776 ; n29776_not
g64259 not n36994 ; n36994_not
g64260 not n19579 ; n19579_not
g64261 not n25798 ; n25798_not
g64262 not n29497 ; n29497_not
g64263 not n38569 ; n38569_not
g64264 not n25789 ; n25789_not
g64265 not n36967 ; n36967_not
g64266 not n36958 ; n36958_not
g64267 not n38938 ; n38938_not
g64268 not n29488 ; n29488_not
g64269 not n38659 ; n38659_not
g64270 not n23989 ; n23989_not
g64271 not n35689 ; n35689_not
g64272 not n38695 ; n38695_not
g64273 not n39568 ; n39568_not
g64274 not n48595 ; n48595_not
g64275 not n19669 ; n19669_not
g64276 not n29299 ; n29299_not
g64277 not n39748 ; n39748_not
g64278 not n29983 ; n29983_not
g64279 not n35977 ; n35977_not
g64280 not n47488 ; n47488_not
g64281 not n36589 ; n36589_not
g64282 not n29866 ; n29866_not
g64283 not n29875 ; n29875_not
g64284 not n39469 ; n39469_not
g64285 not n39874 ; n39874_not
g64286 not n16987 ; n16987_not
g64287 not n29992 ; n29992_not
g64288 not n36598 ; n36598_not
g64289 not n37786 ; n37786_not
g64290 not n28876 ; n28876_not
g64291 not n22999 ; n22999_not
g64292 not n39487 ; n39487_not
g64293 not n39496 ; n39496_not
g64294 not n37858 ; n37858_not
g64295 not n26788 ; n26788_not
g64296 not n29848 ; n29848_not
g64297 not n15988 ; n15988_not
g64298 not n48478 ; n48478_not
g64299 not n15979 ; n15979_not
g64300 not n39784 ; n39784_not
g64301 not n17689 ; n17689_not
g64302 not n39595 ; n39595_not
g64303 not n48559 ; n48559_not
g64304 not n28399 ; n28399_not
g64305 not n39559 ; n39559_not
g64306 not n43798 ; n43798_not
g64307 not n29839 ; n29839_not
g64308 not n17698 ; n17698_not
g64309 not n19849 ; n19849_not
g64310 not n27976 ; n27976_not
g64311 not n29956 ; n29956_not
g64312 not n46579 ; n46579_not
g64313 not n35986 ; n35986_not
g64314 not n34897 ; n34897_not
g64315 not n28687 ; n28687_not
g64316 not n47479 ; n47479_not
g64317 not n37939 ; n37939_not
g64318 not n46895 ; n46895_not
g64319 not n19688 ; n19688_not
g64320 not n28967 ; n28967_not
g64321 not n19769 ; n19769_not
g64322 not n39389 ; n39389_not
g64323 not n38489 ; n38489_not
g64324 not n29984 ; n29984_not
g64325 not n14999 ; n14999_not
g64326 not n34799 ; n34799_not
g64327 not n17969 ; n17969_not
g64328 not n39596 ; n39596_not
g64329 not n43799 ; n43799_not
g64330 not n38588 ; n38588_not
g64331 not n27887 ; n27887_not
g64332 not n39929 ; n39929_not
g64333 not n19499 ; n19499_not
g64334 not n36986 ; n36986_not
g64335 not n29498 ; n29498_not
g64336 not n29669 ; n29669_not
g64337 not n47849 ; n47849_not
g64338 not n19877 ; n19877_not
g64339 not n36887 ; n36887_not
g64340 not n45887 ; n45887_not
g64341 not n38768 ; n38768_not
g64342 not n19778 ; n19778_not
g64343 not n36896 ; n36896_not
g64344 not n35978 ; n35978_not
g64345 not n17789 ; n17789_not
g64346 not n23999 ; n23999_not
g64347 not n48398 ; n48398_not
g64348 not n46868 ; n46868_not
g64349 not n39569 ; n39569_not
g64350 not n47885 ; n47885_not
g64351 not n39857 ; n39857_not
g64352 not n27896 ; n27896_not
g64353 not n19859 ; n19859_not
g64354 not n19679 ; n19679_not
g64355 not n18869 ; n18869_not
g64356 not n47669 ; n47669_not
g64357 not n27779 ; n27779_not
g64358 not n35699 ; n35699_not
g64359 not n39992 ; n39992_not
g64360 not n37949 ; n37949_not
g64361 not n48578 ; n48578_not
g64362 not n39578 ; n39578_not
g64363 not n26888 ; n26888_not
g64364 not n27797 ; n27797_not
g64365 not n27968 ; n27968_not
g64366 not n48983 ; n48983_not
g64367 not n48299 ; n48299_not
g64368 not n33989 ; n33989_not
g64369 not n28895 ; n28895_not
g64370 not n17987 ; n17987_not
g64371 not n39776 ; n39776_not
g64372 not n29678 ; n29678_not
g64373 not n28877 ; n28877_not
g64374 not n39668 ; n39668_not
g64375 not n28886 ; n28886_not
g64376 not n28499 ; n28499_not
g64377 not n28976 ; n28976_not
g64378 not n39794 ; n39794_not
g64379 not n42899 ; n42899_not
g64380 not n39983 ; n39983_not
g64381 not n37778 ; n37778_not
g64382 not n38957 ; n38957_not
g64383 not n39767 ; n39767_not
g64384 not n17978 ; n17978_not
g64385 not n47696 ; n47696_not
g64386 not n25889 ; n25889_not
g64387 not n39956 ; n39956_not
g64388 not n37499 ; n37499_not
g64389 not n27959 ; n27959_not
g64390 not n39848 ; n39848_not
g64391 not n29894 ; n29894_not
g64392 not n26987 ; n26987_not
g64393 not n28778 ; n28778_not
g64394 not n15998 ; n15998_not
g64395 not n27878 ; n27878_not
g64396 not n27977 ; n27977_not
g64397 not n39677 ; n39677_not
g64398 not n29993 ; n29993_not
g64399 not n29588 ; n29588_not
g64400 not n29759 ; n29759_not
g64401 not n45698 ; n45698_not
g64402 not n29966 ; n29966_not
g64403 not n39965 ; n39965_not
g64404 not n45689 ; n45689_not
g64405 not n29849 ; n29849_not
g64406 not n39938 ; n39938_not
g64407 not n16898 ; n16898_not
g64408 not n46967 ; n46967_not
g64409 not n38399 ; n38399_not
g64410 not n28787 ; n28787_not
g64411 not n25988 ; n25988_not
g64412 not n29795 ; n29795_not
g64413 not n18986 ; n18986_not
g64414 not n28958 ; n28958_not
g64415 not n18689 ; n18689_not
g64416 not n38966 ; n38966_not
g64417 not n17798 ; n17798_not
g64418 not n45896 ; n45896_not
g64419 not n32999 ; n32999_not
g64420 not n36689 ; n36689_not
g64421 not n39839 ; n39839_not
g64422 not n46787 ; n46787_not
g64423 not n37994 ; n37994_not
g64424 not n39686 ; n39686_not
g64425 not n28598 ; n28598_not
g64426 not n47975 ; n47975_not
g64427 not n35798 ; n35798_not
g64428 not n25997 ; n25997_not
g64429 not n19796 ; n19796_not
g64430 not n38498 ; n38498_not
g64431 not n26897 ; n26897_not
g64432 not n47588 ; n47588_not
g64433 not n37796 ; n37796_not
g64434 not n35996 ; n35996_not
g64435 not n19976 ; n19976_not
g64436 not n37958 ; n37958_not
g64437 not n26996 ; n26996_not
g64438 not n18968 ; n18968_not
g64439 not n47579 ; n47579_not
g64440 not n18788 ; n18788_not
g64441 not n19994 ; n19994_not
g64442 not n27599 ; n27599_not
g64443 not n18977 ; n18977_not
g64444 not n37967 ; n37967_not
g64445 not n45977 ; n45977_not
g64446 not n29399 ; n29399_not
g64447 not n25979 ; n25979_not
g64448 not n36779 ; n36779_not
g64449 not n45968 ; n45968_not
g64450 not n38948 ; n38948_not
g64451 not n46688 ; n46688_not
g64452 not n29876 ; n29876_not
g64453 not n47597 ; n47597_not
g64454 not n47399 ; n47399_not
g64455 not n38849 ; n38849_not
g64456 not n41999 ; n41999_not
g64457 not n19787 ; n19787_not
g64458 not n42998 ; n42998_not
g64459 not n29687 ; n29687_not
g64460 not n38795 ; n38795_not
g64461 not n27788 ; n27788_not
g64462 not n38777 ; n38777_not
g64463 not n29597 ; n29597_not
g64464 not n18599 ; n18599_not
g64465 not n35997 ; n35997_not
g64466 not n38769 ; n38769_not
g64467 not n36879 ; n36879_not
g64468 not n29895 ; n29895_not
g64469 not n28869 ; n28869_not
g64470 not n26898 ; n26898_not
g64471 not n38949 ; n38949_not
g64472 not n38598 ; n38598_not
g64473 not n17997 ; n17997_not
g64474 not n17889 ; n17889_not
g64475 not n29598 ; n29598_not
g64476 not n46995 ; n46995_not
g64477 not n26799 ; n26799_not
g64478 not n36789 ; n36789_not
g64479 not n37896 ; n37896_not
g64480 not n38994 ; n38994_not
g64481 not n18699 ; n18699_not
g64482 not n47769 ; n47769_not
g64483 not n39993 ; n39993_not
g64484 not n38985 ; n38985_not
g64485 not n38688 ; n38688_not
g64486 not n37878 ; n37878_not
g64487 not n39885 ; n39885_not
g64488 not n27978 ; n27978_not
g64489 not n38877 ; n38877_not
g64490 not n39786 ; n39786_not
g64491 not n36888 ; n36888_not
g64492 not n28968 ; n28968_not
g64493 not n28689 ; n28689_not
g64494 not n37869 ; n37869_not
g64495 not n48984 ; n48984_not
g64496 not n37599 ; n37599_not
g64497 not n39768 ; n39768_not
g64498 not n26979 ; n26979_not
g64499 not n38787 ; n38787_not
g64500 not n19986 ; n19986_not
g64501 not n39867 ; n39867_not
g64502 not n38796 ; n38796_not
g64503 not n19995 ; n19995_not
g64504 not n19689 ; n19689_not
g64505 not n17988 ; n17988_not
g64506 not n39975 ; n39975_not
g64507 not n39588 ; n39588_not
g64508 not n39678 ; n39678_not
g64509 not n47499 ; n47499_not
g64510 not n47859 ; n47859_not
g64511 not n48498 ; n48498_not
g64512 not n37986 ; n37986_not
g64513 not n37698 ; n37698_not
g64514 not n39687 ; n39687_not
g64515 not n38958 ; n38958_not
g64516 not n26988 ; n26988_not
g64517 not n35799 ; n35799_not
g64518 not n39948 ; n39948_not
g64519 not n27897 ; n27897_not
g64520 not n19887 ; n19887_not
g64521 not n47985 ; n47985_not
g64522 not n38895 ; n38895_not
g64523 not n29877 ; n29877_not
g64524 not n38886 ; n38886_not
g64525 not n16998 ; n16998_not
g64526 not n37995 ; n37995_not
g64527 not n46797 ; n46797_not
g64528 not n37779 ; n37779_not
g64529 not n16899 ; n16899_not
g64530 not n19797 ; n19797_not
g64531 not n38679 ; n38679_not
g64532 not n28797 ; n28797_not
g64533 not n24999 ; n24999_not
g64534 not n36798 ; n36798_not
g64535 not n28878 ; n28878_not
g64536 not n38976 ; n38976_not
g64537 not n19788 ; n19788_not
g64538 not n18996 ; n18996_not
g64539 not n39957 ; n39957_not
g64540 not n46959 ; n46959_not
g64541 not n19878 ; n19878_not
g64542 not n28788 ; n28788_not
g64543 not n17899 ; n17899_not
g64544 not n28888 ; n28888_not
g64545 not n29968 ; n29968_not
g64546 not n37978 ; n37978_not
g64547 not n43999 ; n43999_not
g64548 not n39994 ; n39994_not
g64549 not n37789 ; n37789_not
g64550 not n37888 ; n37888_not
g64551 not n26998 ; n26998_not
g64552 not n28699 ; n28699_not
g64553 not n36889 ; n36889_not
g64554 not n39589 ; n39589_not
g64555 not n38788 ; n38788_not
g64556 not n19897 ; n19897_not
g64557 not n18799 ; n18799_not
g64558 not n27988 ; n27988_not
g64559 not n29788 ; n29788_not
g64560 not n48598 ; n48598_not
g64561 not n38869 ; n38869_not
g64562 not n48796 ; n48796_not
g64563 not n34999 ; n34999_not
g64564 not n39697 ; n39697_not
g64565 not n38995 ; n38995_not
g64566 not n39886 ; n39886_not
g64567 not n19798 ; n19798_not
g64568 not n39868 ; n39868_not
g64569 not n29959 ; n29959_not
g64570 not n48787 ; n48787_not
g64571 not n47995 ; n47995_not
g64572 not n39499 ; n39499_not
g64573 not n29977 ; n29977_not
g64574 not n39877 ; n39877_not
g64575 not n38959 ; n38959_not
g64576 not n29887 ; n29887_not
g64577 not n39796 ; n39796_not
g64578 not n29986 ; n29986_not
g64579 not n28897 ; n28897_not
g64580 not n39769 ; n39769_not
g64581 not n46987 ; n46987_not
g64582 not n39895 ; n39895_not
g64583 not n38986 ; n38986_not
g64584 not n39688 ; n39688_not
g64585 not n29797 ; n29797_not
g64586 not n39958 ; n39958_not
g64587 not n19888 ; n19888_not
g64588 not n38968 ; n38968_not
g64589 not n47797 ; n47797_not
g64590 not n36997 ; n36997_not
g64591 not n45997 ; n45997_not
g64592 not n46879 ; n46879_not
g64593 not n38689 ; n38689_not
g64594 not n29779 ; n29779_not
g64595 not n38698 ; n38698_not
g64596 not n39598 ; n39598_not
g64597 not n18989 ; n18989_not
g64598 not n26999 ; n26999_not
g64599 not n27989 ; n27989_not
g64600 not n29789 ; n29789_not
g64601 not n28979 ; n28979_not
g64602 not n37898 ; n37898_not
g64603 not n18899 ; n18899_not
g64604 not n39869 ; n39869_not
g64605 not n27998 ; n27998_not
g64606 not n19898 ; n19898_not
g64607 not n17999 ; n17999_not
g64608 not n39986 ; n39986_not
g64609 not n46979 ; n46979_not
g64610 not n48896 ; n48896_not
g64611 not n39788 ; n39788_not
g64612 not n47789 ; n47789_not
g64613 not n39779 ; n39779_not
g64614 not n28889 ; n28889_not
g64615 not n47897 ; n47897_not
g64616 not n27899 ; n27899_not
g64617 not n29996 ; n29996_not
g64618 not n37799 ; n37799_not
g64619 not n36899 ; n36899_not
g64620 not n38798 ; n38798_not
g64621 not n45899 ; n45899_not
g64622 not n39896 ; n39896_not
g64623 not n38879 ; n38879_not
g64624 not n37889 ; n37889_not
g64625 not n47969 ; n47969_not
g64626 not n38699 ; n38699_not
g64627 not n37988 ; n37988_not
g64628 not n29888 ; n29888_not
g64629 not n47996 ; n47996_not
g64630 not n27999 ; n27999_not
g64631 not n18999 ; n18999_not
g64632 not n39699 ; n39699_not
g64633 not n37899 ; n37899_not
g64634 not n39969 ; n39969_not
g64635 not n39987 ; n39987_not
g64636 not n48897 ; n48897_not
g64637 not n46899 ; n46899_not
g64638 not n39897 ; n39897_not
g64639 not n39888 ; n39888_not
g64640 not n37998 ; n37998_not
g64641 not n19989 ; n19989_not
g64642 not n38988 ; n38988_not
g64643 not n48789 ; n48789_not
g64644 not n48799 ; n48799_not
g64645 not n38899 ; n38899_not
g64646 not n37999 ; n37999_not
g64647 not n39988 ; n39988_not
g64648 not n29989 ; n29989_not
g64649 not n19999 ; n19999_not
g64650 not n39898 ; n39898_not
g64651 not n39997 ; n39997_not
g64652 not n46999 ; n46999_not
g64653 not n29999 ; n29999_not
g64654 not n39999 ; n39999_not
g64655 not pi0100 ; pi0100_not
g64656 not pi0200 ; pi0200_not
g64657 not pi0110 ; pi0110_not
g64658 not pi1100 ; pi1100_not
g64659 not pi0101 ; pi0101_not
g64660 not pi1101 ; pi1101_not
g64661 not pi0210 ; pi0210_not
g64662 not pi0300 ; pi0300_not
g64663 not pi0120 ; pi0120_not
g64664 not pi0102 ; pi0102_not
g64665 not pi0111 ; pi0111_not
g64666 not pi1110 ; pi1110_not
g64667 not pi0201 ; pi0201_not
g64668 not pi0211 ; pi0211_not
g64669 not pi0130 ; pi0130_not
g64670 not pi0103 ; pi0103_not
g64671 not pi0040 ; pi0040_not
g64672 not pi0301 ; pi0301_not
g64673 not pi0121 ; pi0121_not
g64674 not pi1120 ; pi1120_not
g64675 not pi1102 ; pi1102_not
g64676 not pi1111 ; pi1111_not
g64677 not pi0400 ; pi0400_not
g64678 not pi0031 ; pi0031_not
g64679 not pi0202 ; pi0202_not
g64680 not pi0220 ; pi0220_not
g64681 not pi0212 ; pi0212_not
g64682 not pi0230 ; pi0230_not
g64683 not pi0410 ; pi0410_not
g64684 not pi1112 ; pi1112_not
g64685 not pi0113 ; pi0113_not
g64686 not pi0140 ; pi0140_not
g64687 not pi0401 ; pi0401_not
g64688 not pi0032 ; pi0032_not
g64689 not pi0221 ; pi0221_not
g64690 not pi1121 ; pi1121_not
g64691 not pi0500 ; pi0500_not
g64692 not pi1103 ; pi1103_not
g64693 not pi1130 ; pi1130_not
g64694 not pi0104 ; pi0104_not
g64695 not pi0122 ; pi0122_not
g64696 not pi1040 ; pi1040_not
g64697 not pi0050 ; pi0050_not
g64698 not pi0203 ; pi0203_not
g64699 not pi0311 ; pi0311_not
g64700 not pi0041 ; pi0041_not
g64701 not pi0320 ; pi0320_not
g64702 not pi0150 ; pi0150_not
g64703 not pi1131 ; pi1131_not
g64704 not pi0411 ; pi0411_not
g64705 not pi0051 ; pi0051_not
g64706 not pi1104 ; pi1104_not
g64707 not pi0330 ; pi0330_not
g64708 not pi0222 ; pi0222_not
g64709 not pi0024 ; pi0024_not
g64710 not pi0060 ; pi0060_not
g64711 not pi0141 ; pi0141_not
g64712 not pi1113 ; pi1113_not
g64713 not pi0213 ; pi0213_not
g64714 not pi1122 ; pi1122_not
g64715 not pi0321 ; pi0321_not
g64716 not pi0114 ; pi0114_not
g64717 not pi0312 ; pi0312_not
g64718 not pi0123 ; pi0123_not
g64719 not pi0033 ; pi0033_not
g64720 not pi0204 ; pi0204_not
g64721 not pi0105 ; pi0105_not
g64722 not pi0042 ; pi0042_not
g64723 not pi0402 ; pi0402_not
g64724 not pi1050 ; pi1050_not
g64725 not pi0132 ; pi0132_not
g64726 not pi0240 ; pi0240_not
g64727 not pi0214 ; pi0214_not
g64728 not pi0160 ; pi0160_not
g64729 not pi0070 ; pi0070_not
g64730 not pi0151 ; pi0151_not
g64731 not pi0232 ; pi0232_not
g64732 not pi0241 ; pi0241_not
g64733 not pi0223 ; pi0223_not
g64734 not pi1150 ; pi1150_not
g64735 not pi0043 ; pi0043_not
g64736 not pi1114 ; pi1114_not
g64737 not pi0115 ; pi0115_not
g64738 not pi1123 ; pi1123_not
g64739 not pi0250 ; pi0250_not
g64740 not pi0052 ; pi0052_not
g64741 not pi1051 ; pi1051_not
g64742 not pi0700 ; pi0700_not
g64743 not pi1132 ; pi1132_not
g64744 not pi1105 ; pi1105_not
g64745 not pi0034 ; pi0034_not
g64746 not pi0142 ; pi0142_not
g64747 not pi0331 ; pi0331_not
g64748 not pi0601 ; pi0601_not
g64749 not pi0340 ; pi0340_not
g64750 not pi0430 ; pi0430_not
g64751 not pi0502 ; pi0502_not
g64752 not pi0421 ; pi0421_not
g64753 not pi0412 ; pi0412_not
g64754 not pi0205 ; pi0205_not
g64755 not pi0520 ; pi0520_not
g64756 not pi0224 ; pi0224_not
g64757 not pi0215 ; pi0215_not
g64758 not pi0053 ; pi0053_not
g64759 not pi0161 ; pi0161_not
g64760 not pi0152 ; pi0152_not
g64761 not pi0062 ; pi0062_not
g64762 not pi1151 ; pi1151_not
g64763 not pi0044 ; pi0044_not
g64764 not pi0080 ; pi0080_not
g64765 not pi1160 ; pi1160_not
g64766 not pi0116 ; pi0116_not
g64767 not pi0314 ; pi0314_not
g64768 not pi0413 ; pi0413_not
g64769 not pi0404 ; pi0404_not
g64770 not pi0602 ; pi0602_not
g64771 not pi1124 ; pi1124_not
g64772 not pi0071 ; pi0071_not
g64773 not pi0125 ; pi0125_not
g64774 not pi1106 ; pi1106_not
g64775 not pi1142 ; pi1142_not
g64776 not pi0170 ; pi0170_not
g64777 not pi1115 ; pi1115_not
g64778 not pi0332 ; pi0332_not
g64779 not pi0701 ; pi0701_not
g64780 not pi1061 ; pi1061_not
g64781 not pi0233 ; pi0233_not
g64782 not pi0431 ; pi0431_not
g64783 not pi0710 ; pi0710_not
g64784 not pi0107 ; pi0107_not
g64785 not pi0422 ; pi0422_not
g64786 not pi0440 ; pi0440_not
g64787 not pi1133 ; pi1133_not
g64788 not pi0323 ; pi0323_not
g64789 not pi0143 ; pi0143_not
g64790 not pi1070 ; pi1070_not
g64791 not pi0341 ; pi0341_not
g64792 not pi0530 ; pi0530_not
g64793 not pi1043 ; pi1043_not
g64794 not pi0035 ; pi0035_not
g64795 not pi0521 ; pi0521_not
g64796 not pi0350 ; pi0350_not
g64797 not pi0206 ; pi0206_not
g64798 not pi0351 ; pi0351_not
g64799 not pi0207 ; pi0207_not
g64800 not pi0090 ; pi0090_not
g64801 not pi0603 ; pi0603_not
g64802 not pi0252 ; pi0252_not
g64803 not pi0072 ; pi0072_not
g64804 not pi0036 ; pi0036_not
g64805 not pi0630 ; pi0630_not
g64806 not pi0225 ; pi0225_not
g64807 not pi1116 ; pi1116_not
g64808 not pi0216 ; pi0216_not
g64809 not pi0054 ; pi0054_not
g64810 not pi1107 ; pi1107_not
g64811 not pi0243 ; pi0243_not
g64812 not pi1125 ; pi1125_not
g64813 not pi1143 ; pi1143_not
g64814 not pi0333 ; pi0333_not
g64815 not pi0801 ; pi0801_not
g64816 not pi0414 ; pi0414_not
g64817 not pi0540 ; pi0540_not
g64818 not pi0621 ; pi0621_not
g64819 not pi0702 ; pi0702_not
g64820 not pi0432 ; pi0432_not
g64821 not pi0423 ; pi0423_not
g64822 not pi1062 ; pi1062_not
g64823 not pi1044 ; pi1044_not
g64824 not pi0162 ; pi0162_not
g64825 not pi0144 ; pi0144_not
g64826 not pi0171 ; pi0171_not
g64827 not pi1080 ; pi1080_not
g64828 not pi1152 ; pi1152_not
g64829 not pi0081 ; pi0081_not
g64830 not pi0234 ; pi0234_not
g64831 not pi1053 ; pi1053_not
g64832 not pi0126 ; pi0126_not
g64833 not pi0180 ; pi0180_not
g64834 not pi1134 ; pi1134_not
g64835 not po1101 ; po1101_not
g64836 not pi0810 ; pi0810_not
g64837 not pi0153 ; pi0153_not
g64838 not pi0342 ; pi0342_not
g64839 not pi0045 ; pi0045_not
g64840 not pi0441 ; pi0441_not
g64841 not pi0360 ; pi0360_not
g64842 not pi0135 ; pi0135_not
g64843 not pi0504 ; pi0504_not
g64844 not pi0324 ; pi0324_not
g64845 not pi0900 ; pi0900_not
g64846 not pi0450 ; pi0450_not
g64847 not pi0063 ; pi0063_not
g64848 not pi0108 ; pi0108_not
g64849 not pi0315 ; pi0315_not
g64850 not pi0270 ; pi0270_not
g64851 not pi0118 ; pi0118_not
g64852 not pi0208 ; pi0208_not
g64853 not pi0082 ; pi0082_not
g64854 not pi0145 ; pi0145_not
g64855 not pi0460 ; pi0460_not
g64856 not pi0163 ; pi0163_not
g64857 not pi0046 ; pi0046_not
g64858 not pi0091 ; pi0091_not
g64859 not pi0190 ; pi0190_not
g64860 not pi0073 ; pi0073_not
g64861 not pi0316 ; pi0316_not
g64862 not pi0343 ; pi0343_not
g64863 not pi0172 ; pi0172_not
g64864 not pi1054 ; pi1054_not
g64865 not pi0235 ; pi0235_not
g64866 not pi0325 ; pi0325_not
g64867 not pi0910 ; pi0910_not
g64868 not pi0352 ; pi0352_not
g64869 not pi0262 ; pi0262_not
g64870 not pi0055 ; pi0055_not
g64871 not pi1135 ; pi1135_not
g64872 not pi0280 ; pi0280_not
g64873 not pi1153 ; pi1153_not
g64874 not pi0064 ; pi0064_not
g64875 not pi0730 ; pi0730_not
g64876 not pi1144 ; pi1144_not
g64877 not pi0181 ; pi0181_not
g64878 not pi1072 ; pi1072_not
g64879 not pi0136 ; pi0136_not
g64880 not pi0505 ; pi0505_not
g64881 not pi1117 ; pi1117_not
g64882 not pi1036 ; pi1036_not
g64883 not pi0820 ; pi0820_not
g64884 not pi0703 ; pi0703_not
g64885 not pi0442 ; pi0442_not
g64886 not pi0415 ; pi0415_not
g64887 not pi0361 ; pi0361_not
g64888 not pi1108 ; pi1108_not
g64889 not pi1045 ; pi1045_not
g64890 not pi0451 ; pi0451_not
g64891 not pi1126 ; pi1126_not
g64892 not pi0370 ; pi0370_not
g64893 not pi0271 ; pi0271_not
g64894 not pi0334 ; pi0334_not
g64895 not pi0109 ; pi0109_not
g64896 not pi0154 ; pi0154_not
g64897 not pi0523 ; pi0523_not
g64898 not pi1081 ; pi1081_not
g64899 not pi1063 ; pi1063_not
g64900 not pi0550 ; pi0550_not
g64901 not pi0433 ; pi0433_not
g64902 not pi0127 ; pi0127_not
g64903 not pi0253 ; pi0253_not
g64904 not pi0424 ; pi0424_not
g64905 not pi0074 ; pi0074_not
g64906 not pi0182 ; pi0182_not
g64907 not pi0056 ; pi0056_not
g64908 not pi0704 ; pi0704_not
g64909 not pi0164 ; pi0164_not
g64910 not pi0173 ; pi0173_not
g64911 not pi1154 ; pi1154_not
g64912 not pi1055 ; pi1055_not
g64913 not pi0092 ; pi0092_not
g64914 not pi0191 ; pi0191_not
g64915 not pi0047 ; pi0047_not
g64916 not pi1091 ; pi1091_not
g64917 not pi1118 ; pi1118_not
g64918 not pi0038 ; pi0038_not
g64919 not pi0137 ; pi0137_not
g64920 not pi0641 ; pi0641_not
g64921 not pi1163 ; pi1163_not
g64922 not pi0623 ; pi0623_not
g64923 not pi1037 ; pi1037_not
g64924 not pi1109 ; pi1109_not
g64925 not pi0614 ; pi0614_not
g64926 not pi0281 ; pi0281_not
g64927 not pi0146 ; pi0146_not
g64928 not pi1145 ; pi1145_not
g64929 not pi0263 ; pi0263_not
g64930 not pi0830 ; pi0830_not
g64931 not pi0911 ; pi0911_not
g64932 not pi0902 ; pi0902_not
g64933 not pi0290 ; pi0290_not
g64934 not pi1136 ; pi1136_not
g64935 not pi0425 ; pi0425_not
g64936 not pi0407 ; pi0407_not
g64937 not pi0434 ; pi0434_not
g64938 not pi0155 ; pi0155_not
g64939 not pi1127 ; pi1127_not
g64940 not pi0353 ; pi0353_not
g64941 not pi0524 ; pi0524_not
g64942 not pi0533 ; pi0533_not
g64943 not pi0083 ; pi0083_not
g64944 not pi0380 ; pi0380_not
g64945 not pi1082 ; pi1082_not
g64946 not pi0335 ; pi0335_not
g64947 not pi0065 ; pi0065_not
g64948 not pi0443 ; pi0443_not
g64949 not pi0317 ; pi0317_not
g64950 not pi0452 ; pi0452_not
g64951 not pi0209 ; pi0209_not
g64952 not pi0515 ; pi0515_not
g64953 not pi0326 ; pi0326_not
g64954 not pi0218 ; pi0218_not
g64955 not pi0344 ; pi0344_not
g64956 not pi0920 ; pi0920_not
g64957 not pi0416 ; pi0416_not
g64958 not pi1119 ; pi1119_not
g64959 not pi0237 ; pi0237_not
g64960 not pi1146 ; pi1146_not
g64961 not pi0075 ; pi0075_not
g64962 not pi0147 ; pi0147_not
g64963 not pi0444 ; pi0444_not
g64964 not pi0435 ; pi0435_not
g64965 not pi0039 ; pi0039_not
g64966 not pi0138 ; pi0138_not
g64967 not pi1128 ; pi1128_not
g64968 not pi0093 ; pi0093_not
g64969 not pi0174 ; pi0174_not
g64970 not pi0192 ; pi0192_not
g64971 not pi0183 ; pi0183_not
g64972 not pi0219 ; pi0219_not
g64973 not pi0228 ; pi0228_not
g64974 not pi1155 ; pi1155_not
g64975 not pi0084 ; pi0084_not
g64976 not pi0336 ; pi0336_not
g64977 not pi0246 ; pi0246_not
g64978 not pi0048 ; pi0048_not
g64979 not pi0318 ; pi0318_not
g64980 not pi0552 ; pi0552_not
g64981 not pi0129 ; pi0129_not
g64982 not pi0633 ; pi0633_not
g64983 not pi0903 ; pi0903_not
g64984 not pi0057 ; pi0057_not
g64985 not pi0534 ; pi0534_not
g64986 not pi0390 ; pi0390_not
g64987 not pi0156 ; pi0156_not
g64988 not pi0912 ; pi0912_not
g64989 not pi0741 ; pi0741_not
g64990 not pi0408 ; pi0408_not
g64991 not pi0642 ; pi0642_not
g64992 not pi0282 ; pi0282_not
g64993 not pi0264 ; pi0264_not
g64994 not pi0606 ; pi0606_not
g64995 not pi0354 ; pi0354_not
g64996 not pi0453 ; pi0453_not
g64997 not pi0705 ; pi0705_not
g64998 not pi1074 ; pi1074_not
g64999 not pi0660 ; pi0660_not
g65000 not pi0930 ; pi0930_not
g65001 not pi0165 ; pi0165_not
g65002 not pi0291 ; pi0291_not
g65003 not pi0570 ; pi0570_not
g65004 not pi0723 ; pi0723_not
g65005 not pi0345 ; pi0345_not
g65006 not pi0921 ; pi0921_not
g65007 not pi0480 ; pi0480_not
g65008 not pi1065 ; pi1065_not
g65009 not pi1047 ; pi1047_not
g65010 not pi0255 ; pi0255_not
g65011 not pi0273 ; pi0273_not
g65012 not pi0462 ; pi0462_not
g65013 not pi1093 ; pi1093_not
g65014 not pi0913 ; pi0913_not
g65015 not pi0508 ; pi0508_not
g65016 not pi0382 ; pi0382_not
g65017 not pi1147 ; pi1147_not
g65018 not pi0238 ; pi0238_not
g65019 not pi0364 ; pi0364_not
g65020 not pi1156 ; pi1156_not
g65021 not pi0094 ; pi0094_not
g65022 not pi0058 ; pi0058_not
g65023 not pi0337 ; pi0337_not
g65024 not pi0346 ; pi0346_not
g65025 not pi0571 ; pi0571_not
g65026 not pi0625 ; pi0625_not
g65027 not pi0409 ; pi0409_not
g65028 not pi0292 ; pi0292_not
g65029 not pi0841 ; pi0841_not
g65030 not pi0661 ; pi0661_not
g65031 not pi0049 ; pi0049_not
g65032 not pi1084 ; pi1084_not
g65033 not pi0454 ; pi0454_not
g65034 not pi0634 ; pi0634_not
g65035 not pi0391 ; pi0391_not
g65036 not pi0166 ; pi0166_not
g65037 not pi0355 ; pi0355_not
g65038 not pi0274 ; pi0274_not
g65039 not pi0265 ; pi0265_not
g65040 not pi0373 ; pi0373_not
g65041 not pi1129 ; pi1129_not
g65042 not pi0436 ; pi0436_not
g65043 not pi1048 ; pi1048_not
g65044 not pi1039 ; pi1039_not
g65045 not pi0427 ; pi0427_not
g65046 not pi0715 ; pi0715_not
g65047 not pi0940 ; pi0940_not
g65048 not pi0643 ; pi0643_not
g65049 not pi1057 ; pi1057_not
g65050 not pi0706 ; pi0706_not
g65051 not pi0832 ; pi0832_not
g65052 not pi0328 ; pi0328_not
g65053 not pi0553 ; pi0553_not
g65054 not pi0319 ; pi0319_not
g65055 not pi0904 ; pi0904_not
g65056 not pi0067 ; pi0067_not
g65057 not pi0544 ; pi0544_not
g65058 not pi0139 ; pi0139_not
g65059 not pi0850 ; pi0850_not
g65060 not pi0463 ; pi0463_not
g65061 not pi0607 ; pi0607_not
g65062 not pi0193 ; pi0193_not
g65063 not pi0148 ; pi0148_not
g65064 not pi0751 ; pi0751_not
g65065 not pi0157 ; pi0157_not
g65066 not pi0616 ; pi0616_not
g65067 not pi0742 ; pi0742_not
g65068 not pi0724 ; pi0724_not
g65069 not pi0760 ; pi0760_not
g65070 not pi0256 ; pi0256_not
g65071 not pi0184 ; pi0184_not
g65072 not pi0805 ; pi0805_not
g65073 not pi0175 ; pi0175_not
g65074 not pi0644 ; pi0644_not
g65075 not pi0680 ; pi0680_not
g65076 not pi0626 ; pi0626_not
g65077 not pi0239 ; pi0239_not
g65078 not pi0455 ; pi0455_not
g65079 not pi1157 ; pi1157_not
g65080 not pi0347 ; pi0347_not
g65081 not pi0572 ; pi0572_not
g65082 not pi0176 ; pi0176_not
g65083 not pi0545 ; pi0545_not
g65084 not pi0509 ; pi0509_not
g65085 not pi1049 ; pi1049_not
g65086 not pi0383 ; pi0383_not
g65087 not pi0365 ; pi0365_not
g65088 not pi0338 ; pi0338_not
g65089 not pi0428 ; pi0428_not
g65090 not pi0185 ; pi0185_not
g65091 not pi0833 ; pi0833_not
g65092 not pi0761 ; pi0761_not
g65093 not pi0662 ; pi0662_not
g65094 not pi0743 ; pi0743_not
g65095 not pi0464 ; pi0464_not
g65096 not pi0329 ; pi0329_not
g65097 not pi0095 ; pi0095_not
g65098 not pi0068 ; pi0068_not
g65099 not pi0590 ; pi0590_not
g65100 not pi0446 ; pi0446_not
g65101 not pi0248 ; pi0248_not
g65102 not pi0851 ; pi0851_not
g65103 not pi0077 ; pi0077_not
g65104 not pi0059 ; pi0059_not
g65105 not pi0752 ; pi0752_not
g65106 not pi0167 ; pi0167_not
g65107 not pi0725 ; pi0725_not
g65108 not pi0734 ; pi0734_not
g65109 not pi0158 ; pi0158_not
g65110 not pi1067 ; pi1067_not
g65111 not pi1139 ; pi1139_not
g65112 not pi0266 ; pi0266_not
g65113 not pi1076 ; pi1076_not
g65114 not pi0932 ; pi0932_not
g65115 not pi0806 ; pi0806_not
g65116 not pi0086 ; pi0086_not
g65117 not pi0284 ; pi0284_not
g65118 not pi0554 ; pi0554_not
g65119 not pi0563 ; pi0563_not
g65120 not pi0482 ; pi0482_not
g65121 not pi0617 ; pi0617_not
g65122 not pi0770 ; pi0770_not
g65123 not pi0149 ; pi0149_not
g65124 not pi1058 ; pi1058_not
g65125 not pi0518 ; pi0518_not
g65126 not pi0392 ; pi0392_not
g65127 not pi0905 ; pi0905_not
g65128 not pi0608 ; pi0608_not
g65129 not pi1148 ; pi1148_not
g65130 not pi0194 ; pi0194_not
g65131 not pi0293 ; pi0293_not
g65132 not pi0815 ; pi0815_not
g65133 not pi0824 ; pi0824_not
g65134 not pi0257 ; pi0257_not
g65135 not pi0914 ; pi0914_not
g65136 not pi0618 ; pi0618_not
g65137 not pi0609 ; pi0609_not
g65138 not pi0258 ; pi0258_not
g65139 not pi0159 ; pi0159_not
g65140 not pi0753 ; pi0753_not
g65141 not pi0591 ; pi0591_not
g65142 not pi0825 ; pi0825_not
g65143 not pi0249 ; pi0249_not
g65144 not pi0564 ; pi0564_not
g65145 not pi1158 ; pi1158_not
g65146 not pi0555 ; pi0555_not
g65147 not pi0096 ; pi0096_not
g65148 not pi0483 ; pi0483_not
g65149 not pi0069 ; pi0069_not
g65150 not pi0339 ; pi0339_not
g65151 not pi0447 ; pi0447_not
g65152 not pi0366 ; pi0366_not
g65153 not pi0780 ; pi0780_not
g65154 not pi0087 ; pi0087_not
g65155 not pi0168 ; pi0168_not
g65156 not pi0915 ; pi0915_not
g65157 not pi0186 ; pi0186_not
g65158 not pi0429 ; pi0429_not
g65159 not pi1149 ; pi1149_not
g65160 not pi1059 ; pi1059_not
g65161 not pi0726 ; pi0726_not
g65162 not pi0861 ; pi0861_not
g65163 not pi0627 ; pi0627_not
g65164 not pi0177 ; pi0177_not
g65165 not pi0924 ; pi0924_not
g65166 not pi0276 ; pi0276_not
g65167 not pi0933 ; pi0933_not
g65168 not pi0735 ; pi0735_not
g65169 not pi0681 ; pi0681_not
g65170 not pi0690 ; pi0690_not
g65171 not pi0294 ; pi0294_not
g65172 not pi0816 ; pi0816_not
g65173 not pi0438 ; pi0438_not
g65174 not pi0582 ; pi0582_not
g65175 not pi0537 ; pi0537_not
g65176 not pi0456 ; pi0456_not
g65177 not pi0375 ; pi0375_not
g65178 not pi0519 ; pi0519_not
g65179 not pi0906 ; pi0906_not
g65180 not pi0384 ; pi0384_not
g65181 not pi0619 ; pi0619_not
g65182 not pi0592 ; pi0592_not
g65183 not pi0790 ; pi0790_not
g65184 not pi1069 ; pi1069_not
g65185 not pi0628 ; pi0628_not
g65186 not pi0934 ; pi0934_not
g65187 not pi0196 ; pi0196_not
g65188 not pi0745 ; pi0745_not
g65189 not pi0178 ; pi0178_not
g65190 not pi1159 ; pi1159_not
g65191 not pi0295 ; pi0295_not
g65192 not pi0862 ; pi0862_not
g65193 not pi0079 ; pi0079_not
g65194 not pi0097 ; pi0097_not
g65195 not pi0907 ; pi0907_not
g65196 not pi0691 ; pi0691_not
g65197 not pi0169 ; pi0169_not
g65198 not pi0754 ; pi0754_not
g65199 not pi0727 ; pi0727_not
g65200 not pi0709 ; pi0709_not
g65201 not pi0259 ; pi0259_not
g65202 not pi0637 ; pi0637_not
g65203 not pi0736 ; pi0736_not
g65204 not pi0187 ; pi0187_not
g65205 not pi0763 ; pi0763_not
g65206 not pi0781 ; pi0781_not
g65207 not pi0448 ; pi0448_not
g65208 not pi0088 ; pi0088_not
g65209 not pi0385 ; pi0385_not
g65210 not pi0376 ; pi0376_not
g65211 not pi0439 ; pi0439_not
g65212 not pi0772 ; pi0772_not
g65213 not pi0367 ; pi0367_not
g65214 not pi1078 ; pi1078_not
g65215 not pi0547 ; pi0547_not
g65216 not pi1087 ; pi1087_not
g65217 not pi0817 ; pi0817_not
g65218 not pi0286 ; pi0286_not
g65219 not pi0826 ; pi0826_not
g65220 not pi0538 ; pi0538_not
g65221 not pi0565 ; pi0565_not
g65222 not pi0358 ; pi0358_not
g65223 not pi0349 ; pi0349_not
g65224 not pi0916 ; pi0916_not
g65225 not pi0764 ; pi0764_not
g65226 not pi0647 ; pi0647_not
g65227 not po0740 ; po0740_not
g65228 not pi0629 ; pi0629_not
g65229 not pi1196 ; pi1196_not
g65230 not pi0458 ; pi0458_not
g65231 not pi0755 ; pi0755_not
g65232 not pi0665 ; pi0665_not
g65233 not pi0539 ; pi0539_not
g65234 not pi0188 ; pi0188_not
g65235 not pi0944 ; pi0944_not
g65236 not pi0782 ; pi0782_not
g65237 not pi0179 ; pi0179_not
g65238 not pi0746 ; pi0746_not
g65239 not pi0890 ; pi0890_not
g65240 not pi0584 ; pi0584_not
g65241 not pi0089 ; pi0089_not
g65242 not pi0953 ; pi0953_not
g65243 not pi0836 ; pi0836_not
g65244 not pi0197 ; pi0197_not
g65245 not pi0476 ; pi0476_not
g65246 not pi0287 ; pi0287_not
g65247 not pi0917 ; pi0917_not
g65248 not pi0908 ; pi0908_not
g65249 not pi0935 ; pi0935_not
g65250 not pi0359 ; pi0359_not
g65251 not pi0494 ; pi0494_not
g65252 not pi0296 ; pi0296_not
g65253 not pi0737 ; pi0737_not
g65254 not pi0638 ; pi0638_not
g65255 not pi1079 ; pi1079_not
g65256 not pi0980 ; pi0980_not
g65257 not pi0269 ; pi0269_not
g65258 not pi0386 ; pi0386_not
g65259 not pi0683 ; pi0683_not
g65260 not pi0593 ; pi0593_not
g65261 not pi0098 ; pi0098_not
g65262 not pi0557 ; pi0557_not
g65263 not pi0827 ; pi0827_not
g65264 not pi0377 ; pi0377_not
g65265 not pi0495 ; pi0495_not
g65266 not pi0585 ; pi0585_not
g65267 not pi0774 ; pi0774_not
g65268 not pi0792 ; pi0792_not
g65269 not pi0549 ; pi0549_not
g65270 not pi0099 ; pi0099_not
g65271 not po1038 ; po1038_not
g65272 not pi0639 ; pi0639_not
g65273 not pi0648 ; pi0648_not
g65274 not pi0198 ; pi0198_not
g65275 not pi0189 ; pi0189_not
g65276 not pi0927 ; pi0927_not
g65277 not pi0891 ; pi0891_not
g65278 not pi0288 ; pi0288_not
g65279 not pi0468 ; pi0468_not
g65280 not pi0729 ; pi0729_not
g65281 not pi0486 ; pi0486_not
g65282 not po0840 ; po0840_not
g65283 not pi0945 ; pi0945_not
g65284 not pi0567 ; pi0567_not
g65285 not pi1197 ; pi1197_not
g65286 not pi0909 ; pi0909_not
g65287 not pi0738 ; pi0738_not
g65288 not pi0756 ; pi0756_not
g65289 not pi0954 ; pi0954_not
g65290 not pi0828 ; pi0828_not
g65291 not pi0558 ; pi0558_not
g65292 not pi0279 ; pi0279_not
g65293 not pi0459 ; pi0459_not
g65294 not pi0819 ; pi0819_not
g65295 not pi0297 ; pi0297_not
g65296 not pi0846 ; pi0846_not
g65297 not pi0837 ; pi0837_not
g65298 not pi0918 ; pi0918_not
g65299 not pi0775 ; pi0775_not
g65300 not pi0928 ; pi0928_not
g65301 not pi0757 ; pi0757_not
g65302 not pi1198 ; pi1198_not
g65303 not pi0919 ; pi0919_not
g65304 not pi0397 ; pi0397_not
g65305 not po1057 ; po1057_not
g65306 not pi0388 ; pi0388_not
g65307 not pi0199 ; pi0199_not
g65308 not pi0955 ; pi0955_not
g65309 not pi0892 ; pi0892_not
g65310 not pi0289 ; pi0289_not
g65311 not pi0496 ; pi0496_not
g65312 not pi0595 ; pi0595_not
g65313 not pi0379 ; pi0379_not
g65314 not pi0739 ; pi0739_not
g65315 not pi0829 ; pi0829_not
g65316 not pi0766 ; pi0766_not
g65317 not pi0559 ; pi0559_not
g65318 not pi0883 ; pi0883_not
g65319 not pi0478 ; pi0478_not
g65320 not pi0568 ; pi0568_not
g65321 not pi0937 ; pi0937_not
g65322 not pi0973 ; pi0973_not
g65323 not pi0947 ; pi0947_not
g65324 not pi0884 ; pi0884_not
g65325 not pi0695 ; pi0695_not
g65326 not pi0785 ; pi0785_not
g65327 not pi0479 ; pi0479_not
g65328 not pi0767 ; pi0767_not
g65329 not pi0497 ; pi0497_not
g65330 not pi0758 ; pi0758_not
g65331 not pi0299 ; pi0299_not
g65332 not pi0578 ; pi0578_not
g65333 not pi0749 ; pi0749_not
g65334 not pi1199 ; pi1199_not
g65335 not pi0569 ; pi0569_not
g65336 not po1049 ; po1049_not
g65337 not pi0938 ; pi0938_not
g65338 not pi0587 ; pi0587_not
g65339 not pi0686 ; pi0686_not
g65340 not pi0875 ; pi0875_not
g65341 not pi0488 ; pi0488_not
g65342 not pi0398 ; pi0398_not
g65343 not pi0659 ; pi0659_not
g65344 not po0950 ; po0950_not
g65345 not pi0777 ; pi0777_not
g65346 not pi0894 ; pi0894_not
g65347 not pi0489 ; pi0489_not
g65348 not pi0768 ; pi0768_not
g65349 not pi0696 ; pi0696_not
g65350 not pi0759 ; pi0759_not
g65351 not pi0795 ; pi0795_not
g65352 not pi0687 ; pi0687_not
g65353 not pi0948 ; pi0948_not
g65354 not pi0399 ; pi0399_not
g65355 not pi0885 ; pi0885_not
g65356 not pi0939 ; pi0939_not
g65357 not pi0588 ; pi0588_not
g65358 not pi0778 ; pi0778_not
g65359 not pi0787 ; pi0787_not
g65360 not pi0598 ; pi0598_not
g65361 not pi0796 ; pi0796_not
g65362 not po0637 ; po0637_not
g65363 not pi0976 ; pi0976_not
g65364 not pi0958 ; pi0958_not
g65365 not pi0877 ; pi0877_not
g65366 not pi0886 ; pi0886_not
g65367 not pi0895 ; pi0895_not
g65368 not pi0769 ; pi0769_not
g65369 not pi0688 ; pi0688_not
g65370 not po0980 ; po0980_not
g65371 not pi0788 ; pi0788_not
g65372 not pi0698 ; pi0698_not
g65373 not pi0887 ; pi0887_not
g65374 not pi0869 ; pi0869_not
g65375 not pi0599 ; pi0599_not
g65376 not pi0779 ; pi0779_not
g65377 not pi0896 ; pi0896_not
g65378 not pi0878 ; pi0878_not
g65379 not pi0968 ; pi0968_not
g65380 not pi0959 ; pi0959_not
g65381 not pi0789 ; pi0789_not
g65382 not po0954 ; po0954_not
g65383 not po0963 ; po0963_not
g65384 not pi0879 ; pi0879_not
g65385 not pi0699 ; pi0699_not
g65386 not pi0888 ; pi0888_not
g65387 not pi0979 ; pi0979_not
g65388 not pi0889 ; pi0889_not
g65389 not pi0898 ; pi0898_not
g65390 not pi0899 ; pi0899_not
g65391 not pi0999 ; pi0999_not
g65392 not po0978 ; po0978_not
g65393 not po0988 ; po0988_not
