name log2
i a[0]
i a[1]
i a[2]
i a[3]
i a[4]
i a[5]
i a[6]
i a[7]
i a[8]
i a[9]
i a[10]
i a[11]
i a[12]
i a[13]
i a[14]
i a[15]
i a[16]
i a[17]
i a[18]
i a[19]
i a[20]
i a[21]
i a[22]
i a[23]
i a[24]
i a[25]
i a[26]
i a[27]
i a[28]
i a[29]
i a[30]
i a[31]

o result[0]
o result[1]
o result[2]
o result[3]
o result[4]
o result[5]
o result[6]
o result[7]
o result[8]
o result[9]
o result[10]
o result[11]
o result[12]
o result[13]
o result[14]
o result[15]
o result[16]
o result[17]
o result[18]
o result[19]
o result[20]
o result[21]
o result[22]
o result[23]
o result[24]
o result[25]
o result[26]
o result[27]
o result[28]
o result[29]
o result[30]
o result[31]

g1 and a[4] a[5]_not ; n65
g2 and a[4]_not a[5] ; n66
g3 nor n65 n66 ; n67
g4 and a[2] a[3]_not ; n68
g5 and a[2]_not a[3] ; n69
g6 nor n68 n69 ; n70
g7 and n67 n70_not ; n71
g8 and a[29]_not a[30] ; n72
g9 and a[29] a[30]_not ; n73
g10 nor n72 n73 ; n74
g11 and a[31] n74_not ; n75
g12 nor a[24] a[25] ; n76
g13 and a[23]_not a[26] ; n77
g14 and n76 n77 ; n78
g15 and a[27] a[28] ; n79
g16 and n73 n79 ; n80
g17 and n78 n80 ; n81
g18 nor a[27] a[28] ; n82
g19 and n73 n82 ; n83
g20 and a[24] a[25] ; n84
g21 and n77 n84 ; n85
g22 and n83 n85 ; n86
g23 nor a[23] a[26] ; n87
g24 and n76 n87 ; n88
g25 and a[29] a[30] ; n89
g26 and n79 n89 ; n90
g27 and n88 n90 ; n91
g28 and a[23] a[26]_not ; n92
g29 and a[24]_not a[25] ; n93
g30 and n92 n93 ; n94
g31 and n83 n94 ; n95
g32 and n84 n92 ; n96
g33 nor a[29] a[30] ; n97
g34 and n82 n97 ; n98
g35 and n96 n98 ; n99
g36 nor n95 n99 ; n100
g37 and n87 n93 ; n101
g38 and n90 n101 ; n102
g39 and a[27] a[28]_not ; n103
g40 and n89 n103 ; n104
g41 and a[23] a[26] ; n105
g42 and n93 n105 ; n106
g43 and n104 n106 ; n107
g44 nor n102 n107 ; n108
g45 and a[27]_not a[28] ; n109
g46 and n72 n109 ; n110
g47 and n96 n110 ; n111
g48 and a[24] a[25]_not ; n112
g49 and n92 n112 ; n113
g50 and n72 n103 ; n114
g51 and n113 n114 ; n115
g52 nor n111 n115 ; n116
g53 and n82 n89 ; n117
g54 and n94 n117 ; n118
g55 and n83 n106 ; n119
g56 nor n118 n119 ; n120
g57 and n88 n117 ; n121
g58 and n87 n112 ; n122
g59 and n110 n122 ; n123
g60 and n77 n93 ; n124
g61 and n83 n124 ; n125
g62 and n105 n112 ; n126
g63 and n83 n126 ; n127
g64 nor n125 n127 ; n128
g65 and n97 n109 ; n129
g66 and n113 n129 ; n130
g67 and n76 n92 ; n131
g68 and n129 n131 ; n132
g69 nor n130 n132 ; n133
g70 and n72 n82 ; n134
g71 and n113 n134 ; n135
g72 and n110 n126 ; n136
g73 nor n135 n136 ; n137
g74 and n133 n137 ; n138
g75 and n128 n138 ; n139
g76 and n123_not n139 ; n140
g77 and n121_not n140 ; n141
g78 and n98 n126 ; n142
g79 and n79 n97 ; n143
g80 and n122 n143 ; n144
g81 and n78 n143 ; n145
g82 and n104 n126 ; n146
g83 and n78 n117 ; n147
g84 and n77 n112 ; n148
g85 and n117 n148 ; n149
g86 and n114 n124 ; n150
g87 and n114 n122 ; n151
g88 and n101 n134 ; n152
g89 and n72 n79 ; n153
g90 and n126 n153 ; n154
g91 and n117 n124 ; n155
g92 nor n154 n155 ; n156
g93 and n94 n129 ; n157
g94 and n83 n148 ; n158
g95 nor n157 n158 ; n159
g96 and n73 n109 ; n160
g97 and n94 n160 ; n161
g98 and n84 n105 ; n162
g99 and n129 n162 ; n163
g100 and n85 n143 ; n164
g101 and n124 n143 ; n165
g102 and n97 n103 ; n166
g103 and n124 n166 ; n167
g104 and n114 n126 ; n168
g105 and n85 n153 ; n169
g106 and n129 n148 ; n170
g107 and n114 n131 ; n171
g108 nor n170 n171 ; n172
g109 and n88 n143 ; n173
g110 and n89 n109 ; n174
g111 and n106 n174 ; n175
g112 and n84 n87 ; n176
g113 and n117 n176 ; n177
g114 nor n175 n177 ; n178
g115 and n173_not n178 ; n179
g116 and n172 n179 ; n180
g117 and n169_not n180 ; n181
g118 and n168_not n181 ; n182
g119 and n167_not n182 ; n183
g120 and n165_not n183 ; n184
g121 and n164_not n184 ; n185
g122 and n163_not n185 ; n186
g123 and n161_not n186 ; n187
g124 and n80 n124 ; n188
g125 and n106 n114 ; n189
g126 and n122 n153 ; n190
g127 and n98 n162 ; n191
g128 and n101 n166 ; n192
g129 nor n191 n192 ; n193
g130 and n110 n113 ; n194
g131 and n193 n194_not ; n195
g132 and n190_not n195 ; n196
g133 and n189_not n196 ; n197
g134 and n188_not n197 ; n198
g135 and n73 n103 ; n199
g136 and n176 n199 ; n200
g137 and n126 n199 ; n201
g138 nor n200 n201 ; n202
g139 and n126 n174 ; n203
g140 and n202 n203_not ; n204
g141 and n94 n143 ; n205
g142 and n90 n148 ; n206
g143 nor n205 n206 ; n207
g144 and n204 n207 ; n208
g145 and n198 n208 ; n209
g146 and n187 n209 ; n210
g147 and n159 n210 ; n211
g148 and n156 n211 ; n212
g149 and n152_not n212 ; n213
g150 and n151_not n213 ; n214
g151 and n150_not n214 ; n215
g152 and n149_not n215 ; n216
g153 and n147_not n216 ; n217
g154 and n146_not n217 ; n218
g155 and n145_not n218 ; n219
g156 and n144_not n219 ; n220
g157 and n142_not n220 ; n221
g158 and n80 n85 ; n222
g159 and n117 n162 ; n223
g160 and n85 n134 ; n224
g161 and n88 n199 ; n225
g162 and n94 n104 ; n226
g163 nor n225 n226 ; n227
g164 and n90 n122 ; n228
g165 and n78 n153 ; n229
g166 nor n228 n229 ; n230
g167 and n80 n106 ; n231
g168 and n126 n134 ; n232
g169 and n78 n174 ; n233
g170 nor n232 n233 ; n234
g171 and n231_not n234 ; n235
g172 and n85 n110 ; n236
g173 and n148 n199 ; n237
g174 nor n236 n237 ; n238
g175 and n85 n117 ; n239
g176 and n143 n148 ; n240
g177 nor n239 n240 ; n241
g178 and n153 n176 ; n242
g179 and n143 n176 ; n243
g180 nor n242 n243 ; n244
g181 and n98 n124 ; n245
g182 and n126 n166 ; n246
g183 nor n245 n246 ; n247
g184 and n104 n162 ; n248
g185 and n80 n131 ; n249
g186 nor n248 n249 ; n250
g187 and n83 n131 ; n251
g188 and n106 n199 ; n252
g189 nor n251 n252 ; n253
g190 and n114 n176 ; n254
g191 and n106 n134 ; n255
g192 nor n254 n255 ; n256
g193 and n253 n256 ; n257
g194 and n250 n257 ; n258
g195 and n247 n258 ; n259
g196 and n244 n259 ; n260
g197 and n241 n260 ; n261
g198 and n238 n261 ; n262
g199 and n235 n262 ; n263
g200 and n230 n263 ; n264
g201 and n227 n264 ; n265
g202 and n224_not n265 ; n266
g203 and n223_not n266 ; n267
g204 and n222_not n267 ; n268
g205 and n76 n105 ; n269
g206 and n80 n269 ; n270
g207 and n83 n88 ; n271
g208 and n131 n199 ; n272
g209 and n126 n129 ; n273
g210 and n131 n143 ; n274
g211 and n113 n117 ; n275
g212 and n110 n131 ; n276
g213 and n96 n160 ; n277
g214 and n134 n162 ; n278
g215 nor n277 n278 ; n279
g216 and n101 n114 ; n280
g217 and n96 n134 ; n281
g218 nor n280 n281 ; n282
g219 and n98 n131 ; n283
g220 and n134 n148 ; n284
g221 nor n283 n284 ; n285
g222 and n131 n166 ; n286
g223 and n90 n94 ; n287
g224 nor n286 n287 ; n288
g225 and n94 n134 ; n289
g226 and n96 n104 ; n290
g227 nor n289 n290 ; n291
g228 and n104 n131 ; n292
g229 and n83 n162 ; n293
g230 nor n292 n293 ; n294
g231 and n124 n160 ; n295
g232 and n94 n166 ; n296
g233 nor n295 n296 ; n297
g234 and n98 n176 ; n298
g235 and n117 n131 ; n299
g236 nor n298 n299 ; n300
g237 and n110 n176 ; n301
g238 and n90 n124 ; n302
g239 nor n301 n302 ; n303
g240 and n88 n160 ; n304
g241 and n104 n269 ; n305
g242 and n129 n269 ; n306
g243 nor n305 n306 ; n307
g244 and n304_not n307 ; n308
g245 and n303 n308 ; n309
g246 and n300 n309 ; n310
g247 and n297 n310 ; n311
g248 and n294 n311 ; n312
g249 and n291 n312 ; n313
g250 and n288 n313 ; n314
g251 and n285 n314 ; n315
g252 and n282 n315 ; n316
g253 and n279 n316 ; n317
g254 and n276_not n317 ; n318
g255 and n275_not n318 ; n319
g256 and n274_not n319 ; n320
g257 and n273_not n320 ; n321
g258 and n272_not n321 ; n322
g259 and n271_not n322 ; n323
g260 and n270_not n323 ; n324
g261 and n83 n101 ; n325
g262 and n90 n162 ; n326
g263 and n162 n174 ; n327
g264 and n88 n114 ; n328
g265 and n78 n134 ; n329
g266 and n94 n153 ; n330
g267 and n162 n166 ; n331
g268 and n160 n269 ; n332
g269 nor n331 n332 ; n333
g270 and n174 n176 ; n334
g271 and n94 n114 ; n335
g272 nor n334 n335 ; n336
g273 and n80 n101 ; n337
g274 and n85 n199 ; n338
g275 and n101 n174 ; n339
g276 and n113 n160 ; n340
g277 nor n339 n340 ; n341
g278 and n338_not n341 ; n342
g279 and n337_not n342 ; n343
g280 and n336 n343 ; n344
g281 and n333 n344 ; n345
g282 and n330_not n345 ; n346
g283 and n329_not n346 ; n347
g284 and n328_not n347 ; n348
g285 and n327_not n348 ; n349
g286 and n326_not n349 ; n350
g287 and n325_not n350 ; n351
g288 and n122 n174 ; n352
g289 and n134 n176 ; n353
g290 and n124 n134 ; n354
g291 and n134 n269 ; n355
g292 nor n354 n355 ; n356
g293 and n90 n269 ; n357
g294 and n83 n269 ; n358
g295 nor n357 n358 ; n359
g296 and n356 n359 ; n360
g297 and n353_not n360 ; n361
g298 and n352_not n361 ; n362
g299 and n80 n94 ; n363
g300 and n110 n162 ; n364
g301 nor n363 n364 ; n365
g302 and n96 n199 ; n366
g303 and n104 n113 ; n367
g304 and n98 n113 ; n368
g305 nor n367 n368 ; n369
g306 and n366_not n369 ; n370
g307 and n85 n160 ; n371
g308 and n88 n98 ; n372
g309 nor n371 n372 ; n373
g310 and n90 n96 ; n374
g311 and n78 n129 ; n375
g312 nor n374 n375 ; n376
g313 and n373 n376 ; n377
g314 and n370 n377 ; n378
g315 and n365 n378 ; n379
g316 and n362 n379 ; n380
g317 and n351 n380 ; n381
g318 and n324 n381 ; n382
g319 and n268 n382 ; n383
g320 and n221 n383 ; n384
g321 and n141 n384 ; n385
g322 and n120 n385 ; n386
g323 and n116 n386 ; n387
g324 and n108 n387 ; n388
g325 and n100 n388 ; n389
g326 and n91_not n389 ; n390
g327 and n86_not n390 ; n391
g328 and n81_not n391 ; n392
g329 and n85 n129 ; n393
g330 and n124 n129 ; n394
g331 and n90 n113 ; n395
g332 and n78 n104 ; n396
g333 and n106 n110 ; n397
g334 and n131 n153 ; n398
g335 nor n327 n398 ; n399
g336 and n88 n104 ; n400
g337 nor n335 n400 ; n401
g338 and n101 n104 ; n402
g339 and n104 n148 ; n403
g340 nor n402 n403 ; n404
g341 and n375_not n404 ; n405
g342 and n401 n405 ; n406
g343 and n399 n406 ; n407
g344 and n111_not n407 ; n408
g345 and n397_not n408 ; n409
g346 and n177_not n409 ; n410
g347 and n299_not n410 ; n411
g348 and n396_not n411 ; n412
g349 and n395_not n412 ; n413
g350 and n325_not n413 ; n414
g351 and n293_not n414 ; n415
g352 and n78 n90 ; n416
g353 and n117 n122 ; n417
g354 nor n364 n417 ; n418
g355 and n96 n117 ; n419
g356 and n106 n153 ; n420
g357 nor n419 n420 ; n421
g358 and n98 n148 ; n422
g359 nor n146 n422 ; n423
g360 and n101 n143 ; n424
g361 and n166 n269 ; n425
g362 and n114 n148 ; n426
g363 and n110 n148 ; n427
g364 and n80 n176 ; n428
g365 and n80 n148 ; n429
g366 and n148 n166 ; n430
g367 nor n144 n430 ; n431
g368 and n201_not n431 ; n432
g369 and n429_not n432 ; n433
g370 and n428_not n433 ; n434
g371 and n117 n269 ; n435
g372 and n160 n176 ; n436
g373 nor n435 n436 ; n437
g374 and n88 n166 ; n438
g375 nor n371 n438 ; n439
g376 and n437 n439 ; n440
g377 and n434 n440 ; n441
g378 and n427_not n441 ; n442
g379 and n194_not n442 ; n443
g380 and n426_not n443 ; n444
g381 and n280_not n444 ; n445
g382 and n367_not n445 ; n446
g383 and n425_not n446 ; n447
g384 and n424_not n447 ; n448
g385 and n80 n122 ; n449
g386 nor n271 n449 ; n450
g387 and n199 n269 ; n451
g388 and n85 n98 ; n452
g389 and n98 n101 ; n453
g390 nor n452 n453 ; n454
g391 and n289_not n454 ; n455
g392 and n292_not n455 ; n456
g393 and n286_not n456 ; n457
g394 and n225_not n457 ; n458
g395 and n451_not n458 ; n459
g396 and n104 n176 ; n460
g397 and n85 n104 ; n461
g398 and n148 n153 ; n462
g399 nor n461 n462 ; n463
g400 and n460_not n463 ; n464
g401 and n283_not n464 ; n465
g402 and n96 n143 ; n466
g403 nor n233 n466 ; n467
g404 and n106 n129 ; n468
g405 and n94 n110 ; n469
g406 and n94 n199 ; n470
g407 nor n366 n470 ; n471
g408 and n469_not n471 ; n472
g409 and n468_not n472 ; n473
g410 and n101 n160 ; n474
g411 nor n188 n474 ; n475
g412 and n473 n475 ; n476
g413 and n467 n476 ; n477
g414 and n465 n477 ; n478
g415 and n459 n478 ; n479
g416 and n450 n479 ; n480
g417 and n448 n480 ; n481
g418 and n159 n481 ; n482
g419 and n423 n482 ; n483
g420 and n421 n483 ; n484
g421 and n418 n484 ; n485
g422 and n254_not n485 ; n486
g423 and n416_not n486 ; n487
g424 and n337_not n487 ; n488
g425 and n83 n176 ; n489
g426 and n90 n106 ; n490
g427 nor n489 n490 ; n491
g428 and n166 n176 ; n492
g429 and n129 n176 ; n493
g430 nor n167 n493 ; n494
g431 and n85 n174 ; n495
g432 and n78 n166 ; n496
g433 nor n495 n496 ; n497
g434 and n494 n497 ; n498
g435 and n242_not n498 ; n499
g436 and n189_not n499 ; n500
g437 and n290_not n500 ; n501
g438 and n492_not n501 ; n502
g439 and n231_not n502 ; n503
g440 and n143 n162 ; n504
g441 and n96 n166 ; n505
g442 and n96 n174 ; n506
g443 nor n81 n506 ; n507
g444 nor n275 n334 ; n508
g445 and n101 n153 ; n509
g446 nor n135 n509 ; n510
g447 and n114 n269 ; n511
g448 nor n248 n511 ; n512
g449 and n104 n124 ; n513
g450 and n174 n269 ; n514
g451 nor n306 n357 ; n515
g452 and n161_not n515 ; n516
g453 and n332_not n516 ; n517
g454 and n96 n153 ; n518
g455 and n122 n160 ; n519
g456 nor n518 n519 ; n520
g457 and n517 n520 ; n521
g458 and n514_not n521 ; n522
g459 and n513_not n522 ; n523
g460 and n274_not n523 ; n524
g461 and n160 n162 ; n525
g462 nor n272 n525 ; n526
g463 and n104 n122 ; n527
g464 nor n115 n305 ; n528
g465 and n527_not n528 ; n529
g466 nor n127 n223 ; n530
g467 and n101 n199 ; n531
g468 and n148 n160 ; n532
g469 nor n340 n532 ; n533
g470 and n531_not n533 ; n534
g471 and n338_not n534 ; n535
g472 and n78 n98 ; n536
g473 and n98 n122 ; n537
g474 nor n368 n537 ; n538
g475 and n536_not n538 ; n539
g476 and n298_not n539 ; n540
g477 and n358_not n540 ; n541
g478 and n535 n541 ; n542
g479 and n530 n542 ; n543
g480 and n529 n543 ; n544
g481 and n526 n544 ; n545
g482 and n524 n545 ; n546
g483 and n512 n546 ; n547
g484 and n510 n547 ; n548
g485 and n508 n548 ; n549
g486 and n507 n549 ; n550
g487 and n108 n550 ; n551
g488 and n169_not n551 ; n552
g489 and n147_not n552 ; n553
g490 and n505_not n553 ; n554
g491 and n504_not n554 ; n555
g492 and n245_not n555 ; n556
g493 and n88 n134 ; n557
g494 and n88 n110 ; n558
g495 nor n557 n558 ; n559
g496 and n226_not n559 ; n560
g497 and n277_not n560 ; n561
g498 and n80 n162 ; n562
g499 and n85 n166 ; n563
g500 and n78 n160 ; n564
g501 nor n563 n564 ; n565
g502 and n562_not n565 ; n566
g503 and n98 n269 ; n567
g504 and n122 n166 ; n568
g505 and n83 n122 ; n569
g506 nor n568 n569 ; n570
g507 and n88 n174 ; n571
g508 and n570 n571_not ; n572
g509 and n567_not n572 ; n573
g510 and n566 n573 ; n574
g511 and n561 n574 ; n575
g512 and n556 n575 ; n576
g513 and n503 n576 ; n577
g514 and n491 n577 ; n578
g515 and n488 n578 ; n579
g516 and n415 n579 ; n580
g517 and n193 n580 ; n581
g518 and n152_not n581 ; n582
g519 and n302_not n582 ; n583
g520 and n243_not n583 ; n584
g521 and n394_not n584 ; n585
g522 and n393_not n585 ; n586
g523 and n249_not n586 ; n587
g524 nor n392 n587 ; n588
g525 and n96 n129 ; n589
g526 nor n188 n222 ; n590
g527 nor n194 n490 ; n591
g528 and n124 n199 ; n592
g529 nor n228 n592 ; n593
g530 and n117 n126 ; n594
g531 nor n205 n594 ; n595
g532 and n593 n595 ; n596
g533 and n136_not n596 ; n597
g534 and n177_not n597 ; n598
g535 and n394_not n598 ; n599
g536 and n119_not n599 ; n600
g537 and n106 n143 ; n601
g538 and n114 n162 ; n602
g539 and n101 n129 ; n603
g540 nor n493 n603 ; n604
g541 and n359 n604 ; n605
g542 and n602_not n605 ; n606
g543 and n299_not n606 ; n607
g544 and n107_not n607 ; n608
g545 and n243_not n608 ; n609
g546 and n601_not n609 ; n610
g547 and n393_not n610 ; n611
g548 and n470_not n611 ; n612
g549 and n272_not n612 ; n613
g550 and n340_not n613 ; n614
g551 nor n151 n327 ; n615
g552 and n229_not n376 ; n616
g553 and n110 n269 ; n617
g554 nor n171 n617 ; n618
g555 and n124 n174 ; n619
g556 and n131 n134 ; n620
g557 nor n619 n620 ; n621
g558 nor n175 n525 ; n622
g559 and n162 n199 ; n623
g560 nor n135 n152 ; n624
g561 and n335_not n624 ; n625
g562 and n150_not n625 ; n626
g563 and n248_not n626 ; n627
g564 and n164_not n627 ; n628
g565 and n623_not n628 ; n629
g566 and n532_not n629 ; n630
g567 and n86_not n630 ; n631
g568 nor n102 n242 ; n632
g569 and n80 n126 ; n633
g570 nor n424 n633 ; n634
g571 and n154_not n634 ; n635
g572 and n400_not n635 ; n636
g573 and n101 n117 ; n637
g574 nor n571 n637 ; n638
g575 and n90 n126 ; n639
g576 nor n505 n639 ; n640
g577 and n78 n114 ; n641
g578 nor n492 n641 ; n642
g579 and n640 n642 ; n643
g580 and n638 n643 ; n644
g581 and n636 n644 ; n645
g582 and n632 n645 ; n646
g583 and n631 n646 ; n647
g584 and n622 n647 ; n648
g585 and n621 n648 ; n649
g586 and n618 n649 ; n650
g587 and n398_not n650 ; n651
g588 and n149_not n651 ; n652
g589 and n223_not n652 ; n653
g590 nor n123 n125 ; n654
g591 and n80 n113 ; n655
g592 and n94 n174 ; n656
g593 and n113 n199 ; n657
g594 nor n452 n657 ; n658
g595 and n427_not n658 ; n659
g596 and n353_not n659 ; n660
g597 and n426_not n660 ; n661
g598 and n656_not n661 ; n662
g599 and n292_not n662 ; n663
g600 and n655_not n663 ; n664
g601 nor n283 n567 ; n665
g602 and n83 n96 ; n666
g603 and n153 n162 ; n667
g604 nor n281 n667 ; n668
g605 and n430_not n668 ; n669
g606 and n519_not n669 ; n670
g607 and n666_not n670 ; n671
g608 and n106 n160 ; n672
g609 and n143 n269 ; n673
g610 nor n672 n673 ; n674
g611 nor n144 n568 ; n675
g612 and n674 n675 ; n676
g613 and n671 n676 ; n677
g614 and n665 n677 ; n678
g615 and n664 n678 ; n679
g616 and n654 n679 ; n680
g617 and n450 n680 ; n681
g618 and n330_not n681 ; n682
g619 and n419_not n682 ; n683
g620 and n461_not n683 ; n684
g621 and n527_not n684 ; n685
g622 and n422_not n685 ; n686
g623 and n170_not n686 ; n687
g624 and n562_not n687 ; n688
g625 and n113 n143 ; n689
g626 nor n190 n689 ; n690
g627 nor n329 n339 ; n691
g628 nor n420 n536 ; n692
g629 and n468_not n692 ; n693
g630 nor n145 n254 ; n694
g631 and n693 n694 ; n695
g632 and n691 n695 ; n696
g633 and n690 n696 ; n697
g634 and n688 n697 ; n698
g635 and n653 n698 ; n699
g636 and n616 n699 ; n700
g637 and n333 n700 ; n701
g638 and n615 n701 ; n702
g639 and n614 n702 ; n703
g640 and n600 n703 ; n704
g641 and n591 n704 ; n705
g642 and n202 n705 ; n706
g643 and n590 n706 ; n707
g644 and n514_not n707 ; n708
g645 and n326_not n708 ; n709
g646 and n589_not n709 ; n710
g647 nor n587 n710 ; n711
g648 and n78 n199 ; n712
g649 and n122 n134 ; n713
g650 and n126 n143 ; n714
g651 and n90 n131 ; n715
g652 and n113 n166 ; n716
g653 and n137 n462_not ; n717
g654 and n367_not n717 ; n718
g655 and n716_not n718 ; n719
g656 nor n164 n251 ; n720
g657 nor n155 n469 ; n721
g658 and n374_not n721 ; n722
g659 nor n147 n460 ; n723
g660 and n722 n723 ; n724
g661 and n355_not n724 ; n725
g662 and n146_not n725 ; n726
g663 and n286_not n726 ; n727
g664 and n567_not n727 ; n728
g665 and n393_not n728 ; n729
g666 and n338_not n729 ; n730
g667 nor n145 n571 ; n731
g668 nor n371 n474 ; n732
g669 nor n173 n519 ; n733
g670 and n158_not n733 ; n734
g671 nor n536 n656 ; n735
g672 and n734 n735 ; n736
g673 and n732 n736 ; n737
g674 and n242_not n737 ; n738
g675 and n289_not n738 ; n739
g676 and n305_not n739 ; n740
g677 and n248_not n740 ; n741
g678 and n453_not n741 ; n742
g679 and n394_not n742 ; n743
g680 and n95_not n743 ; n744
g681 and n363_not n744 ; n745
g682 and n101 n110 ; n746
g683 nor n206 n302 ; n747
g684 and n746_not n747 ; n748
g685 and n425_not n748 ; n749
g686 and n99_not n749 ; n750
g687 and n592_not n750 ; n751
g688 and n124 n153 ; n752
g689 nor n154 n752 ; n753
g690 and n563_not n753 ; n754
g691 and n193 n490_not ; n755
g692 and n237_not n755 ; n756
g693 and n304_not n756 ; n757
g694 and n754 n757 ; n758
g695 and n751 n758 ; n759
g696 and n745 n759 ; n760
g697 and n731 n760 ; n761
g698 and n730 n761 ; n762
g699 and n720 n762 ; n763
g700 and n719 n763 ; n764
g701 and n227 n764 ; n765
g702 and n203_not n765 ; n766
g703 and n715_not n766 ; n767
g704 and n714_not n767 ; n768
g705 and n165_not n768 ; n769
g706 and n429_not n769 ; n770
g707 and n80 n88 ; n771
g708 nor n451 n771 ; n772
g709 nor n190 n240 ; n773
g710 nor n358 n402 ; n774
g711 nor n364 n427 ; n775
g712 nor n278 n328 ; n776
g713 and n85 n90 ; n777
g714 nor n337 n777 ; n778
g715 and n776 n778 ; n779
g716 and n775 n779 ; n780
g717 and n774 n780 ; n781
g718 and n773 n781 ; n782
g719 and n290_not n782 ; n783
g720 and n357_not n783 ; n784
g721 and n416_not n784 ; n785
g722 and n372_not n785 ; n786
g723 and n271_not n786 ; n787
g724 nor n86 n493 ; n788
g725 nor n470 n667 ; n789
g726 nor n403 n513 ; n790
g727 and n98 n106 ; n791
g728 nor n168 n791 ; n792
g729 nor n161 n245 ; n793
g730 and n792 n793 ; n794
g731 and n790 n794 ; n795
g732 and n789 n795 ; n796
g733 and n622 n796 ; n797
g734 and n177_not n797 ; n798
g735 and n396_not n798 ; n799
g736 and n277_not n799 ; n800
g737 and n788 n800 ; n801
g738 and n449_not n801 ; n802
g739 and n96 n114 ; n803
g740 nor n326 n511 ; n804
g741 nor n495 n514 ; n805
g742 nor n296 n492 ; n806
g743 and n422_not n806 ; n807
g744 and n375_not n807 ; n808
g745 and n113 n174 ; n809
g746 nor n430 n809 ; n810
g747 nor n150 n284 ; n811
g748 nor n149 n417 ; n812
g749 nor n623 n641 ; n813
g750 and n666_not n813 ; n814
g751 nor n169 n620 ; n815
g752 and n672_not n815 ; n816
g753 and n814 n816 ; n817
g754 and n812 n817 ; n818
g755 and n811 n818 ; n819
g756 and n810 n819 ; n820
g757 and n228_not n820 ; n821
g758 and n243_not n821 ; n822
g759 and n366_not n822 ; n823
g760 and n562_not n823 ; n824
g761 and n90 n176 ; n825
g762 nor n246 n420 ; n826
g763 nor n295 n564 ; n827
g764 and n826 n827 ; n828
g765 and n121_not n828 ; n829
g766 and n825_not n829 ; n830
g767 nor n504 n518 ; n831
g768 and n270_not n831 ; n832
g769 and n467 n832 ; n833
g770 and n830 n833 ; n834
g771 and n824 n834 ; n835
g772 and n808 n835 ; n836
g773 and n805 n836 ; n837
g774 and n804 n837 ; n838
g775 and n509_not n838 ; n839
g776 and n557_not n839 ; n840
g777 and n254_not n840 ; n841
g778 and n803_not n841 ; n842
g779 and n280_not n842 ; n843
g780 and n532_not n843 ; n844
g781 and n120 n654 ; n845
g782 and n189_not n845 ; n846
g783 and n88 n153 ; n847
g784 nor n558 n847 ; n848
g785 and n223_not n848 ; n849
g786 and n617_not n849 ; n850
g787 and n353_not n850 ; n851
g788 and n846 n851 ; n852
g789 and n844 n852 ; n853
g790 and n802 n853 ; n854
g791 and n787 n854 ; n855
g792 and n772 n855 ; n856
g793 and n770 n856 ; n857
g794 and n713_not n857 ; n858
g795 and n151_not n858 ; n859
g796 and n299_not n859 ; n860
g797 and n639_not n860 ; n861
g798 and n496_not n861 ; n862
g799 and n142_not n862 ; n863
g800 and n468_not n863 ; n864
g801 and n712_not n864 ; n865
g802 and n489_not n865 ; n866
g803 and n188_not n866 ; n867
g804 nor n710 n867 ; n868
g805 nor n224 n243 ; n869
g806 nor n155 n254 ; n870
g807 and n777_not n870 ; n871
g808 and n304_not n871 ; n872
g809 nor n144 n713 ; n873
g810 nor n236 n272 ; n874
g811 and n80 n96 ; n875
g812 nor n301 n513 ; n876
g813 nor n330 n715 ; n877
g814 and n876 n877 ; n878
g815 and n602_not n878 ; n879
g816 and n205_not n879 ; n880
g817 and n325_not n880 ; n881
g818 and n875_not n881 ; n882
g819 and n78 n83 ; n883
g820 and n106 n117 ; n884
g821 nor n86 n296 ; n885
g822 and n83 n113 ; n886
g823 nor n426 n562 ; n887
g824 nor n326 n637 ; n888
g825 and n496_not n888 ; n889
g826 and n887 n889 ; n890
g827 and n594_not n890 ; n891
g828 and n419_not n891 ; n892
g829 and n417_not n892 ; n893
g830 and n886_not n893 ; n894
g831 and n429_not n894 ; n895
g832 nor n425 n489 ; n896
g833 nor n338 n427 ; n897
g834 and n354_not n719 ; n898
g835 and n393_not n898 ; n899
g836 and n897 n899 ; n900
g837 and n851 n900 ; n901
g838 and n539 n901 ; n902
g839 and n128 n902 ; n903
g840 and n896 n903 ; n904
g841 and n399 n904 ; n905
g842 and n895 n905 ; n906
g843 and n507 n906 ; n907
g844 and n885 n907 ; n908
g845 and n229_not n908 ; n909
g846 and n572 n909 ; n910
g847 and n619_not n910 ; n911
g848 and n884_not n911 ; n912
g849 and n825_not n912 ; n913
g850 and n331_not n913 ; n914
g851 and n883_not n914 ; n915
g852 and n428_not n915 ; n916
g853 nor n242 n335 ; n917
g854 and n771_not n917 ; n918
g855 nor n194 n589 ; n919
g856 and n130_not n919 ; n920
g857 and n633_not n920 ; n921
g858 and n179 n921 ; n922
g859 and n918 n922 ; n923
g860 and n255_not n923 ; n924
g861 and n189_not n924 ; n925
g862 and n328_not n925 ; n926
g863 and n809_not n926 ; n927
g864 and n461_not n927 ; n928
g865 and n395_not n928 ; n929
g866 and n145_not n929 ; n930
g867 and n251_not n930 ; n931
g868 and n88 n129 ; n932
g869 nor n436 n932 ; n933
g870 and n235 n933 ; n934
g871 and n454 n934 ; n935
g872 and n142_not n935 ; n936
g873 nor n119 n438 ; n937
g874 and n281_not n937 ; n938
g875 and n352_not n938 ; n939
g876 and n623_not n939 ; n940
g877 nor n147 n295 ; n941
g878 and n475 n941 ; n942
g879 and n940 n942 ; n943
g880 and n936 n943 ; n944
g881 and n931 n944 ; n945
g882 and n916 n945 ; n946
g883 and n882 n946 ; n947
g884 and n874 n947 ; n948
g885 and n873 n948 ; n949
g886 and n872 n949 ; n950
g887 and n423 n950 ; n951
g888 and n869 n951 ; n952
g889 and n746_not n952 ; n953
g890 and n355_not n953 ; n954
g891 and n400_not n954 ; n955
g892 and n374_not n955 ; n956
g893 and n492_not n956 ; n957
g894 and n158_not n957 ; n958
g895 nor n867 n958 ; n959
g896 nor n111 n254 ; n960
g897 and n94 n98 ; n961
g898 nor n397 n961 ; n962
g899 and n960 n962 ; n963
g900 and n352_not n963 ; n964
g901 and n884_not n964 ; n965
g902 and n102_not n965 ; n966
g903 and n240_not n966 ; n967
g904 nor n81 n337 ; n968
g905 and n276_not n968 ; n969
g906 and n299_not n969 ; n970
g907 and n513_not n970 ; n971
g908 and n165_not n971 ; n972
g909 and n791_not n972 ; n973
g910 and n531_not n973 ; n974
g911 and n489_not n974 ; n975
g912 and n883_not n975 ; n976
g913 nor n394 n429 ; n977
g914 nor n326 n639 ; n978
g915 nor n353 n620 ; n979
g916 and n106 n166 ; n980
g917 nor n203 n286 ; n981
g918 and n366_not n981 ; n982
g919 and n515 n982 ; n983
g920 and n339_not n983 ; n984
g921 and n118_not n984 ; n985
g922 and n980_not n985 ; n986
g923 and n192_not n986 ; n987
g924 and n173_not n987 ; n988
g925 nor n436 n589 ; n989
g926 nor n466 n493 ; n990
g927 nor n149 n617 ; n991
g928 and n825_not n991 ; n992
g929 and n990 n992 ; n993
g930 and n989 n993 ; n994
g931 and n988 n994 ; n995
g932 and n510 n995 ; n996
g933 and n294 n996 ; n997
g934 and n238 n997 ; n998
g935 and n979 n998 ; n999
g936 and n978 n999 ; n1000
g937 and n227 n1000 ; n1001
g938 and n418 n1001 ; n1002
g939 and n746_not n1002 ; n1003
g940 and n177_not n1003 ; n1004
g941 and n689_not n1004 ; n1005
g942 and n164_not n1005 ; n1006
g943 and n338_not n1006 ; n1007
g944 and n125_not n1007 ; n1008
g945 nor n150 n252 ; n1009
g946 and n131 n160 ; n1010
g947 and n113 n153 ; n1011
g948 nor n400 n672 ; n1012
g949 and n427_not n1012 ; n1013
g950 and n1011_not n1013 ; n1014
g951 and n435_not n1014 ; n1015
g952 and n932_not n1015 ; n1016
g953 and n130_not n1016 ; n1017
g954 and n623_not n1017 ; n1018
g955 and n1010_not n1018 ; n1019
g956 and n564_not n1019 ; n1020
g957 nor n190 n224 ; n1021
g958 and n233_not n1021 ; n1022
g959 and n490_not n1022 ; n1023
g960 and n249_not n1023 ; n1024
g961 nor n154 n273 ; n1025
g962 and n405 n1025 ; n1026
g963 and n1024 n1026 ; n1027
g964 and n1020 n1027 ; n1028
g965 and n431 n803_not ; n1029
g966 and n1028 n1029 ; n1030
g967 and n244 n1030 ; n1031
g968 and n1009 n1031 ; n1032
g969 and n747 n1032 ; n1033
g970 and n123_not n1033 ; n1034
g971 and n426_not n1034 ; n1035
g972 and n416_not n1035 ; n1036
g973 and n142_not n1036 ; n1037
g974 and n422_not n1037 ; n1038
g975 and n251_not n1038 ; n1039
g976 nor n304 n557 ; n1040
g977 and n570 n1040 ; n1041
g978 and n847_not n1041 ; n1042
g979 and n152_not n1042 ; n1043
g980 and n171_not n1043 ; n1044
g981 and n136_not n282 ; n1045
g982 nor n167 n246 ; n1046
g983 and n163_not n1046 ; n1047
g984 and n1045 n1047 ; n1048
g985 and n1044 n1048 ; n1049
g986 and n1039 n1049 ; n1050
g987 and n1008 n1050 ; n1051
g988 and n977 n1051 ; n1052
g989 and n622 n1052 ; n1053
g990 and n976 n1053 ; n1054
g991 and n967 n1054 ; n1055
g992 and n885 n1055 ; n1056
g993 and n602_not n1056 ; n1057
g994 and n506_not n1057 ; n1058
g995 and n425_not n1058 ; n1059
g996 and n157_not n1059 ; n1060
g997 nor n958 n1060 ; n1061
g998 and n131 n174 ; n1062
g999 nor n177 n416 ; n1063
g1000 nor n419 n1011 ; n1064
g1001 and n337_not n1064 ; n1065
g1002 and n398_not n1065 ; n1066
g1003 and n400_not n1066 ; n1067
g1004 and n167_not n1067 ; n1068
g1005 and n875_not n1068 ; n1069
g1006 nor n252 n509 ; n1070
g1007 nor n165 n237 ; n1071
g1008 and n110 n124 ; n1072
g1009 nor n155 n1072 ; n1073
g1010 and n1071 n1073 ; n1074
g1011 and n1070 n1074 ; n1075
g1012 and n301_not n1075 ; n1076
g1013 and n641_not n1076 ; n1077
g1014 and n149_not n1077 ; n1078
g1015 and n107_not n1078 ; n1079
g1016 and n173_not n1079 ; n1080
g1017 nor n189 n296 ; n1081
g1018 and n537_not n1081 ; n1082
g1019 and n422_not n1082 ; n1083
g1020 and n451_not n1083 ; n1084
g1021 nor n274 n531 ; n1085
g1022 and n256 n1085 ; n1086
g1023 and n1084 n1086 ; n1087
g1024 and n1080 n1087 ; n1088
g1025 and n1069 n1088 ; n1089
g1026 and n1063 n1089 ; n1090
g1027 and n159 n1090 ; n1091
g1028 and n570 n1091 ; n1092
g1029 and n115_not n1092 ; n1093
g1030 and n1062_not n1093 ; n1094
g1031 and n298_not n1094 ; n1095
g1032 and n589_not n1095 ; n1096
g1033 and n366_not n1096 ; n1097
g1034 and n340_not n1097 ; n1098
g1035 and n371_not n1098 ; n1099
g1036 and n271_not n1099 ; n1100
g1037 and n148 n174 ; n1101
g1038 and n85 n114 ; n1102
g1039 nor n466 n1102 ; n1103
g1040 and n122 n199 ; n1104
g1041 nor n519 n1104 ; n1105
g1042 and n603_not n1105 ; n1106
g1043 and n771_not n1106 ; n1107
g1044 nor n171 n752 ; n1108
g1045 and n712_not n1108 ; n1109
g1046 and n1107 n1109 ; n1110
g1047 and n1103 n1110 ; n1111
g1048 and n136_not n1111 ; n1112
g1049 and n397_not n1112 ; n1113
g1050 and n462_not n1113 ; n1114
g1051 and n847_not n1114 ; n1115
g1052 and n1101_not n1115 ; n1116
g1053 and n435_not n1116 ; n1117
g1054 and n395_not n1117 ; n1118
g1055 and n127_not n1118 ; n1119
g1056 nor n239 n246 ; n1120
g1057 and n273_not n1120 ; n1121
g1058 and n402_not n1121 ; n1122
g1059 and n716_not n1122 ; n1123
g1060 and n144_not n1123 ; n1124
g1061 and n201_not n1124 ; n1125
g1062 and n332_not n1125 ; n1126
g1063 and n126 n160 ; n1127
g1064 nor n883 n1127 ; n1128
g1065 nor n428 n469 ; n1129
g1066 nor n151 n557 ; n1130
g1067 and n506_not n1130 ; n1131
g1068 nor n424 n803 ; n1132
g1069 nor n121 n276 ; n1133
g1070 and n490_not n1133 ; n1134
g1071 and n666_not n1134 ; n1135
g1072 nor n299 n426 ; n1136
g1073 and n673_not n1136 ; n1137
g1074 and n394_not n1137 ; n1138
g1075 nor n205 n292 ; n1139
g1076 and n564_not n1139 ; n1140
g1077 nor n270 n338 ; n1141
g1078 and n275_not n1141 ; n1142
g1079 and n163_not n1142 ; n1143
g1080 and n1140 n1143 ; n1144
g1081 and n1138 n1144 ; n1145
g1082 and n1135 n1145 ; n1146
g1083 and n1132 n1146 ; n1147
g1084 and n936 n1147 ; n1148
g1085 and n1131 n1148 ; n1149
g1086 and n1129 n1149 ; n1150
g1087 and n654 n1150 ; n1151
g1088 and n1128 n1151 ; n1152
g1089 and n637_not n1152 ; n1153
g1090 and n367_not n1153 ; n1154
g1091 nor n304 n1010 ; n1155
g1092 and n773 n979 ; n1156
g1093 and n132_not n1156 ; n1157
g1094 and n655_not n1157 ; n1158
g1095 nor n99 n305 ; n1159
g1096 and n293_not n1159 ; n1160
g1097 nor n191 n468 ; n1161
g1098 and n281_not n1161 ; n1162
g1099 and n714_not n1162 ; n1163
g1100 and n1160 n1163 ; n1164
g1101 and n776 n1164 ; n1165
g1102 and n1158 n1165 ; n1166
g1103 and n1155 n1166 ; n1167
g1104 and n1154 n1167 ; n1168
g1105 and n1126 n1168 ; n1169
g1106 and n1119 n1169 ; n1170
g1107 and n665 n1170 ; n1171
g1108 and n1100 n1171 ; n1172
g1109 and n896 n1172 ; n1173
g1110 and n937 n1173 ; n1174
g1111 and n617_not n1174 ; n1175
g1112 and n495_not n1175 ; n1176
g1113 and n460_not n1176 ; n1177
g1114 and n562_not n1177 ; n1178
g1115 nor n1060 n1178 ; n1179
g1116 nor n135 n657 ; n1180
g1117 nor n152 n505 ; n1181
g1118 nor n81 n329 ; n1182
g1119 nor n419 n435 ; n1183
g1120 and n238 n937 ; n1184
g1121 and n194_not n1184 ; n1185
g1122 and n675 n1185 ; n1186
g1123 and n751 n1186 ; n1187
g1124 and n1155 n1187 ; n1188
g1125 and n787 n1188 ; n1189
g1126 and n1183 n1189 ; n1190
g1127 and n1182 n1190 ; n1191
g1128 and n301_not n1191 ; n1192
g1129 and n136_not n1192 ; n1193
g1130 and n111_not n1193 ; n1194
g1131 and n354_not n1194 ; n1195
g1132 and n224_not n1195 ; n1196
g1133 and n884_not n1196 ; n1197
g1134 and n173_not n1197 ; n1198
g1135 and n164_not n1198 ; n1199
g1136 and n536_not n1199 ; n1200
g1137 and n603_not n1200 ; n1201
g1138 and n655_not n1201 ; n1202
g1139 and n122 n129 ; n1203
g1140 nor n569 n980 ; n1204
g1141 nor n340 n527 ; n1205
g1142 and n875_not n1205 ; n1206
g1143 and n1204 n1206 ; n1207
g1144 and n327_not n1207 ; n1208
g1145 and n228_not n1208 ; n1209
g1146 and n1203_not n1209 ; n1210
g1147 and n325_not n1210 ; n1211
g1148 nor n154 n254 ; n1212
g1149 and n400_not n1212 ; n1213
g1150 and n102_not n1213 ; n1214
g1151 and n331_not n1214 ; n1215
g1152 and n589_not n1215 ; n1216
g1153 nor n167 n563 ; n1217
g1154 and n306_not n1217 ; n1218
g1155 and n251_not n1218 ; n1219
g1156 nor n422 n656 ; n1220
g1157 and n222_not n1220 ; n1221
g1158 and n982 n1221 ; n1222
g1159 and n1219 n1222 ; n1223
g1160 and n1216 n1223 ; n1224
g1161 and n1154 n1224 ; n1225
g1162 and n802 n1225 ; n1226
g1163 and n1211 n1226 ; n1227
g1164 and n1202 n1227 ; n1228
g1165 and n1181 n1228 ; n1229
g1166 and n1180 n1229 ; n1230
g1167 and n518_not n1230 ; n1231
g1168 and n374_not n1231 ; n1232
g1169 and n601_not n1232 ; n1233
g1170 and n200_not n1233 ; n1234
g1171 and n295_not n1234 ; n1235
g1172 nor n1178 n1235 ; n1236
g1173 nor n224 n397 ; n1237
g1174 nor n150 n417 ; n1238
g1175 and n305_not n1238 ; n1239
g1176 and n374_not n1239 ; n1240
g1177 and n590 n1240 ; n1241
g1178 and n402_not n1241 ; n1242
g1179 and n496_not n1242 ; n1243
g1180 and n424_not n1243 ; n1244
g1181 and n277_not n1244 ; n1245
g1182 and n153 n269 ; n1246
g1183 nor n274 n469 ; n1247
g1184 nor n352 n1101 ; n1248
g1185 nor n192 n251 ; n1249
g1186 and n303 n1249 ; n1250
g1187 and n673_not n1250 ; n1251
g1188 nor n371 n504 ; n1252
g1189 nor n368 n771 ; n1253
g1190 nor n255 n562 ; n1254
g1191 nor n99 n249 ; n1255
g1192 and n814 n1255 ; n1256
g1193 and n734 n1256 ; n1257
g1194 and n1254 n1257 ; n1258
g1195 and n1253 n1258 ; n1259
g1196 and n1252 n1259 ; n1260
g1197 and n495_not n1260 ; n1261
g1198 and n296_not n1261 ; n1262
g1199 and n961_not n1262 ; n1263
g1200 and n567_not n1263 ; n1264
g1201 and n244 n980_not ; n1265
g1202 and n537_not n1265 ; n1266
g1203 and n170_not n1266 ; n1267
g1204 and n86_not n1267 ; n1268
g1205 nor n427 n449 ; n1269
g1206 and n329_not n1269 ; n1270
g1207 and n884_not n1270 ; n1271
g1208 nor n154 n514 ; n1272
g1209 and n533 n617_not ; n1273
g1210 and n398_not n1273 ; n1274
g1211 and n1272 n1274 ; n1275
g1212 and n1271 n1275 ; n1276
g1213 and n1103 n1276 ; n1277
g1214 and n1268 n1277 ; n1278
g1215 and n1264 n1278 ; n1279
g1216 and n1251 n1279 ; n1280
g1217 and n235 n1280 ; n1281
g1218 and n285 n1281 ; n1282
g1219 and n1248 n1282 ; n1283
g1220 and n1247 n1283 ; n1284
g1221 and n1246_not n1284 ; n1285
g1222 and n426_not n1285 ; n1286
g1223 and n189_not n1286 ; n1287
g1224 and n460_not n1287 ; n1288
g1225 and n287_not n1288 ; n1289
g1226 and n932_not n1289 ; n1290
g1227 and n569_not n1290 ; n1291
g1228 nor n558 n803 ; n1292
g1229 nor n375 n639 ; n1293
g1230 and n273_not n1293 ; n1294
g1231 and n735 n1294 ; n1295
g1232 and n359 n1295 ; n1296
g1233 and n509_not n1296 ; n1297
g1234 and n190_not n1297 ; n1298
g1235 and n461_not n1298 ; n1299
g1236 and n601_not n1299 ; n1300
g1237 and n191_not n1300 ; n1301
g1238 and n436_not n1301 ; n1302
g1239 and n125_not n1302 ; n1303
g1240 and n81_not n1303 ; n1304
g1241 and n633_not n1304 ; n1305
g1242 and n78 n110 ; n1306
g1243 nor n395 n689 ; n1307
g1244 and n453_not n1307 ; n1308
g1245 and n1306_not n1308 ; n1309
g1246 and n619_not n1309 ; n1310
g1247 and n290_not n1310 ; n1311
g1248 and n331_not n1311 ; n1312
g1249 and n270_not n1312 ; n1313
g1250 nor n394 n396 ; n1314
g1251 and n451_not n1314 ; n1315
g1252 and n1139 n1315 ; n1316
g1253 and n330_not n1316 ; n1317
g1254 and n339_not n1317 ; n1318
g1255 and n146_not n1318 ; n1319
g1256 and n492_not n1319 ; n1320
g1257 and n714_not n1320 ; n1321
g1258 and n304_not n1321 ; n1322
g1259 and n337_not n1322 ; n1323
g1260 nor n518 n568 ; n1324
g1261 and n157_not n1324 ; n1325
g1262 and n470_not n1325 ; n1326
g1263 and n657_not n1326 ; n1327
g1264 and n428_not n1327 ; n1328
g1265 nor n149 n602 ; n1329
g1266 nor n847 n886 ; n1330
g1267 and n237_not n1330 ; n1331
g1268 nor n200 n299 ; n1332
g1269 and n161_not n1332 ; n1333
g1270 and n1331 n1333 ; n1334
g1271 and n1329 n1334 ; n1335
g1272 and n1328 n1335 ; n1336
g1273 and n1323 n1336 ; n1337
g1274 and n731 n1337 ; n1338
g1275 and n1313 n1338 ; n1339
g1276 and n746_not n1339 ; n1340
g1277 and n281_not n1340 ; n1341
g1278 and n335_not n1341 ; n1342
g1279 and n115_not n1342 ; n1343
g1280 and n239_not n1343 ; n1344
g1281 and n226_not n1344 ; n1345
g1282 nor n118 n354 ; n1346
g1283 nor n367 n400 ; n1347
g1284 and n1346 n1347 ; n1348
g1285 and n830 n1348 ; n1349
g1286 and n1345 n1349 ; n1350
g1287 and n1305 n1350 ; n1351
g1288 and n1292 n1351 ; n1352
g1289 and n1291 n1352 ; n1353
g1290 and n1245 n1353 ; n1354
g1291 and n937 n1354 ; n1355
g1292 and n1237 n1355 ; n1356
g1293 and n194_not n1356 ; n1357
g1294 and n328_not n1357 ; n1358
g1295 and n175_not n1358 ; n1359
g1296 and n637_not n1359 ; n1360
g1297 and n422_not n1360 ; n1361
g1298 and n468_not n1361 ; n1362
g1299 and n531_not n1362 ; n1363
g1300 and n366_not n1363 ; n1364
g1301 nor n1235 n1364 ; n1365
g1302 nor n225 n601 ; n1366
g1303 nor n170 n273 ; n1367
g1304 nor n191 n352 ; n1368
g1305 and n272_not n1368 ; n1369
g1306 nor n305 n506 ; n1370
g1307 and n246_not n1370 ; n1371
g1308 and n712_not n1371 ; n1372
g1309 and n1369 n1372 ; n1373
g1310 and n1367 n1373 ; n1374
g1311 and n111_not n1374 ; n1375
g1312 and n147_not n1375 ; n1376
g1313 and n884_not n1376 ; n1377
g1314 and n302_not n1377 ; n1378
g1315 nor n531 n1306 ; n1379
g1316 nor n329 n474 ; n1380
g1317 and n229_not n1380 ; n1381
g1318 and n354_not n1381 ; n1382
g1319 and n296_not n1382 ; n1383
g1320 and n589_not n1383 ; n1384
g1321 nor n330 n803 ; n1385
g1322 and n791_not n1385 ; n1386
g1323 and n372_not n1386 ; n1387
g1324 nor n331 n932 ; n1388
g1325 nor n203 n461 ; n1389
g1326 and n620_not n1389 ; n1390
g1327 and n519_not n1390 ; n1391
g1328 nor n275 n375 ; n1392
g1329 nor n403 n1102 ; n1393
g1330 and n200_not n1393 ; n1394
g1331 and n1392 n1394 ; n1395
g1332 and n846 n1395 ; n1396
g1333 and n1391 n1396 ; n1397
g1334 and n1388 n1397 ; n1398
g1335 and n1387 n1398 ; n1399
g1336 and n1384 n1399 ; n1400
g1337 and n1379 n1400 ; n1401
g1338 and n1180 n1401 ; n1402
g1339 and n1128 n1402 ; n1403
g1340 and n462_not n1403 ; n1404
g1341 and n232_not n1404 ; n1405
g1342 and n223_not n1405 ; n1406
g1343 and n623_not n1406 ; n1407
g1344 nor n107 n715 ; n1408
g1345 nor n633 n961 ; n1409
g1346 and n1408 n1409 ; n1410
g1347 and n789 n1410 ; n1411
g1348 and n752_not n1411 ; n1412
g1349 and n278_not n1412 ; n1413
g1350 and n326_not n1413 ; n1414
g1351 and n490_not n1414 ; n1415
g1352 and n145_not n1415 ; n1416
g1353 and n99_not n1416 ; n1417
g1354 and n672_not n1417 ; n1418
g1355 and n271_not n1418 ; n1419
g1356 nor n367 n496 ; n1420
g1357 and n673_not n1420 ; n1421
g1358 and n86_not n1421 ; n1422
g1359 nor n91 n164 ; n1423
g1360 nor n165 n495 ; n1424
g1361 nor n619 n771 ; n1425
g1362 nor n276 n592 ; n1426
g1363 and n689_not n1426 ; n1427
g1364 and n429_not n1427 ; n1428
g1365 and n1425 n1428 ; n1429
g1366 and n1219 n1429 ; n1430
g1367 and n1424 n1430 ; n1431
g1368 and n1063 n1431 ; n1432
g1369 and n527_not n1432 ; n1433
g1370 and n102_not n1433 ; n1434
g1371 and n231_not n1434 ; n1435
g1372 nor n395 n571 ; n1436
g1373 and n825_not n1436 ; n1437
g1374 nor n289 n1062 ; n1438
g1375 nor n602 n641 ; n1439
g1376 and n150_not n1439 ; n1440
g1377 and n1065 n1440 ; n1441
g1378 and n1438 n1441 ; n1442
g1379 and n1437 n1442 ; n1443
g1380 and n604 n1443 ; n1444
g1381 and n1435 n1444 ; n1445
g1382 and n1139 n1445 ; n1446
g1383 and n896 n1446 ; n1447
g1384 and n827 n1447 ; n1448
g1385 and n1237 n1448 ; n1449
g1386 and n847_not n1449 ; n1450
g1387 and n417_not n1450 ; n1451
g1388 and n228_not n1451 ; n1452
g1389 and n173_not n1452 ; n1453
g1390 and n95_not n1453 ; n1454
g1391 and n454 n1454 ; n1455
g1392 and n639_not n1455 ; n1456
g1393 nor n152 n567 ; n1457
g1394 and n161_not n1457 ; n1458
g1395 and n1456 n1458 ; n1459
g1396 and n1423 n1459 ; n1460
g1397 and n1422 n1460 ; n1461
g1398 and n1419 n1461 ; n1462
g1399 and n1407 n1462 ; n1463
g1400 and n1378 n1463 ; n1464
g1401 and n1366 n1464 ; n1465
g1402 and n1269 n1465 ; n1466
g1403 and n558_not n1466 ; n1467
g1404 and n509_not n1467 ; n1468
g1405 and n149_not n1468 ; n1469
g1406 and n402_not n1469 ; n1470
g1407 and n777_not n1470 ; n1471
g1408 and n132_not n1471 ; n1472
g1409 nor n1364 n1472 ; n1473
g1410 nor n427 n568 ; n1474
g1411 and n283_not n1474 ; n1475
g1412 nor n232 n332 ; n1476
g1413 nor n395 n416 ; n1477
g1414 and n374_not n1477 ; n1478
g1415 nor n496 n746 ; n1479
g1416 nor n249 n655 ; n1480
g1417 and n253 n1384 ; n1481
g1418 and n284_not n1481 ; n1482
g1419 and n715_not n1482 ; n1483
g1420 and n394_not n1483 ; n1484
g1421 and n132_not n1484 ; n1485
g1422 and n470_not n1485 ; n1486
g1423 and n1010_not n1486 ; n1487
g1424 and n158_not n1487 ; n1488
g1425 nor n107 n1011 ; n1489
g1426 and n170_not n1489 ; n1490
g1427 and n435_not n1490 ; n1491
g1428 and n884_not n1491 ; n1492
g1429 and n331_not n1492 ; n1493
g1430 and n157_not n1493 ; n1494
g1431 and n295_not n1494 ; n1495
g1432 and n127_not n1495 ; n1496
g1433 nor n155 n809 ; n1497
g1434 nor n513 n752 ; n1498
g1435 and n425_not n1498 ; n1499
g1436 and n1497 n1499 ; n1500
g1437 and n1496 n1500 ; n1501
g1438 and n1488 n1501 ; n1502
g1439 and n1480 n1502 ; n1503
g1440 and n1479 n1503 ; n1504
g1441 and n1478 n1504 ; n1505
g1442 and n602_not n1505 ; n1506
g1443 and n334_not n1506 ; n1507
g1444 and n173_not n1507 ; n1508
g1445 and n657_not n1508 ; n1509
g1446 and n569_not n1509 ; n1510
g1447 and n270_not n1510 ; n1511
g1448 and n364_not n960 ; n1512
g1449 and n123_not n1512 ; n1513
g1450 and n713_not n1513 ; n1514
g1451 and n327_not n1514 ; n1515
g1452 and n177_not n1515 ; n1516
g1453 and n275_not n1516 ; n1517
g1454 and n825_not n1517 ; n1518
g1455 and n240_not n1518 ; n1519
g1456 and n272_not n1519 ; n1520
g1457 and n771_not n1520 ; n1521
g1458 nor n223 n562 ; n1522
g1459 nor n149 n298 ; n1523
g1460 nor n146 n495 ; n1524
g1461 and n167_not n1524 ; n1525
g1462 and n603_not n1525 ; n1526
g1463 and n489_not n1526 ; n1527
g1464 nor n353 n396 ; n1528
g1465 and n326_not n1528 ; n1529
g1466 and n449_not n1529 ; n1530
g1467 nor n293 n666 ; n1531
g1468 and n1129 n1531 ; n1532
g1469 and n716_not n1532 ; n1533
g1470 and n1331 n1533 ; n1534
g1471 and n1530 n1534 ; n1535
g1472 and n723 n1535 ; n1536
g1473 and n439 n1536 ; n1537
g1474 and n1527 n1537 ; n1538
g1475 and n1105 n1538 ; n1539
g1476 and n1305 n1539 ; n1540
g1477 and n1523 n1540 ; n1541
g1478 and n1426 n1541 ; n1542
g1479 and n590 n1542 ; n1543
g1480 and n1522 n1543 ; n1544
g1481 and n339_not n1544 ; n1545
g1482 and n505_not n1545 ; n1546
g1483 and n306_not n1546 ; n1547
g1484 and n304_not n1547 ; n1548
g1485 and n525_not n1548 ; n1549
g1486 nor n274 n558 ; n1550
g1487 and n202 n282 ; n1551
g1488 and n1550 n1551 ; n1552
g1489 and n980_not n1552 ; n1553
g1490 and n453_not n1553 ; n1554
g1491 and n277_not n1554 ; n1555
g1492 nor n130 n366 ; n1556
g1493 nor n271 n462 ; n1557
g1494 and n1556 n1557 ; n1558
g1495 and n1555 n1558 ; n1559
g1496 and n1549 n1559 ; n1560
g1497 and n1521 n1560 ; n1561
g1498 and n631 n1561 ; n1562
g1499 and n1511 n1562 ; n1563
g1500 and n1476 n1563 ; n1564
g1501 and n1475 n1564 ; n1565
g1502 and n288 n1565 ; n1566
g1503 and n1379 n1566 ; n1567
g1504 and n424_not n1567 ; n1568
g1505 and n205_not n1568 ; n1569
g1506 and n537_not n1569 ; n1570
g1507 and n161_not n1570 ; n1571
g1508 and n429_not n1571 ; n1572
g1509 nor n1472 n1572 ; n1573
g1510 nor n284 n532 ; n1574
g1511 nor n170 n328 ; n1575
g1512 nor n142 n714 ; n1576
g1513 nor n272 n1203 ; n1577
g1514 and n452_not n772 ; n1578
g1515 and n1577 n1578 ; n1579
g1516 and n1181 n1579 ; n1580
g1517 and n873 n1580 ; n1581
g1518 and n235 n1581 ; n1582
g1519 and n617_not n1582 ; n1583
g1520 and n275_not n1583 ; n1584
g1521 and n86_not n1584 ; n1585
g1522 nor n639 n657 ; n1586
g1523 nor n274 n504 ; n1587
g1524 and n201_not n1587 ; n1588
g1525 and n1428 n1588 ; n1589
g1526 and n1586 n1589 ; n1590
g1527 and n1585 n1590 ; n1591
g1528 and n1480 n1591 ; n1592
g1529 and n120 n1592 ; n1593
g1530 and n1576 n1593 ; n1594
g1531 and n731 n1594 ; n1595
g1532 and n156 n1595 ; n1596
g1533 and n254_not n1596 ; n1597
g1534 and n641_not n1597 ; n1598
g1535 and n171_not n1598 ; n1599
g1536 and n287_not n1599 ; n1600
g1537 nor n177 n236 ; n1601
g1538 nor n161 n354 ; n1602
g1539 nor n190 n280 ; n1603
g1540 nor n603 n1011 ; n1604
g1541 and n1603 n1604 ; n1605
g1542 and n294 n1605 ; n1606
g1543 and n400_not n1606 ; n1607
g1544 and n102_not n1607 ; n1608
g1545 and n496_not n1608 ; n1609
g1546 and n246_not n1609 ; n1610
g1547 nor n492 n1010 ; n1611
g1548 and n1246_not n1611 ; n1612
g1549 and n327_not n1612 ; n1613
g1550 and n637_not n1613 ; n1614
g1551 and n438_not n1614 ; n1615
g1552 nor n111 n601 ; n1616
g1553 and n672_not n1616 ; n1617
g1554 nor n329 n620 ; n1618
g1555 and n980_not n1618 ; n1619
g1556 and n337_not n1619 ; n1620
g1557 and n449_not n1620 ; n1621
g1558 and n1617 n1621 ; n1622
g1559 and n1615 n1622 ; n1623
g1560 and n1610 n1623 ; n1624
g1561 and n1602 n1624 ; n1625
g1562 and n301_not n1625 ; n1626
g1563 and n558_not n1626 ; n1627
g1564 and n461_not n1627 ; n1628
g1565 and n91_not n1628 ; n1629
g1566 and n416_not n1629 ; n1630
g1567 and n368_not n1630 ; n1631
g1568 and n468_not n1631 ; n1632
g1569 and n623_not n1632 ; n1633
g1570 and n277_not n1633 ; n1634
g1571 and n489_not n1634 ; n1635
g1572 nor n424 n1306 ; n1636
g1573 and n278_not n1636 ; n1637
g1574 and n619_not n1637 ; n1638
g1575 and n374_not n1638 ; n1639
g1576 and n251_not n1639 ; n1640
g1577 nor n339 n427 ; n1641
g1578 and n273_not n1641 ; n1642
g1579 and n712_not n1642 ; n1643
g1580 nor n228 n777 ; n1644
g1581 and n223_not n1254 ; n1645
g1582 and n331_not n1645 ; n1646
g1583 and n1644 n1646 ; n1647
g1584 and n1643 n1647 ; n1648
g1585 and n1640 n1648 ; n1649
g1586 and n1635 n1649 ; n1650
g1587 and n1601 n1650 ; n1651
g1588 and n1600 n1651 ; n1652
g1589 and n1575 n1652 ; n1653
g1590 and n423 n1653 ; n1654
g1591 and n745 n1654 ; n1655
g1592 and n1248 n1655 ; n1656
g1593 and n1574 n1656 ; n1657
g1594 and n359 n1657 ; n1658
g1595 and n151_not n1658 ; n1659
g1596 and n326_not n1659 ; n1660
g1597 and n568_not n1660 ; n1661
g1598 and n286_not n1661 ; n1662
g1599 and n567_not n1662 ; n1663
g1600 and n1104_not n1663 ; n1664
g1601 and n271_not n1664 ; n1665
g1602 nor n1572 n1665 ; n1666
g1603 nor n132 n249 ; n1667
g1604 nor n91 n462 ; n1668
g1605 and n428_not n788 ; n1669
g1606 and n849 n1669 ; n1670
g1607 and n933 n1670 ; n1671
g1608 and n1475 n1671 ; n1672
g1609 and n1668 n1672 ; n1673
g1610 and n111_not n1673 ; n1674
g1611 and n716_not n1674 ; n1675
g1612 and n425_not n1675 ; n1676
g1613 and n589_not n1676 ; n1677
g1614 and n531_not n1677 ; n1678
g1615 and n231_not n1678 ; n1679
g1616 nor n714 n1104 ; n1680
g1617 and n633_not n1680 ; n1681
g1618 and n303 n1681 ; n1682
g1619 and n790 n1682 ; n1683
g1620 and n364_not n1683 ; n1684
g1621 and n594_not n1684 ; n1685
g1622 and n435_not n1685 ; n1686
g1623 and n290_not n1686 ; n1687
g1624 nor n169 n189 ; n1688
g1625 and n395_not n1688 ; n1689
g1626 and n601_not n1689 ; n1690
g1627 and n393_not n1690 ; n1691
g1628 nor n429 n518 ; n1692
g1629 nor n136 n299 ; n1693
g1630 and n248_not n1693 ; n1694
g1631 and n474_not n1694 ; n1695
g1632 nor n155 n368 ; n1696
g1633 and n363_not n1696 ; n1697
g1634 and n1695 n1697 ; n1698
g1635 and n778 n1698 ; n1699
g1636 and n1692 n1699 ; n1700
g1637 and n1691 n1700 ; n1701
g1638 and n1687 n1701 ; n1702
g1639 and n1679 n1702 ; n1703
g1640 and n1667 n1703 ; n1704
g1641 and n168_not n1704 ; n1705
g1642 and n287_not n1705 ; n1706
g1643 and n372_not n1706 ; n1707
g1644 and n340_not n1707 ; n1708
g1645 nor n466 n536 ; n1709
g1646 and n1329 n1709 ; n1710
g1647 and n1708 n1710 ; n1711
g1648 and n1161 n1711 ; n1712
g1649 and n152_not n1712 ; n1713
g1650 and n289_not n1713 ; n1714
g1651 and n146_not n1714 ; n1715
g1652 and n715_not n1715 ; n1716
g1653 and n206_not n1716 ; n1717
g1654 and n245_not n1717 ; n1718
g1655 and n158_not n1718 ; n1719
g1656 nor n200 n452 ; n1720
g1657 and n519_not n1720 ; n1721
g1658 and n1294 n1721 ; n1722
g1659 and n123_not n1722 ; n1723
g1660 and n1246_not n1723 ; n1724
g1661 and n355_not n1724 ; n1725
g1662 nor n175 n228 ; n1726
g1663 nor n95 n666 ; n1727
g1664 and n194_not n1727 ; n1728
g1665 and n430_not n1728 ; n1729
g1666 and n274_not n1729 ; n1730
g1667 and n489_not n1730 ; n1731
g1668 nor n353 n1072 ; n1732
g1669 and n397_not n1732 ; n1733
g1670 and n163_not n1733 ; n1734
g1671 and n449_not n1734 ; n1735
g1672 and n490_not n1603 ; n1736
g1673 and n251_not n1736 ; n1737
g1674 nor n243 n637 ; n1738
g1675 nor n107 n883 ; n1739
g1676 nor n119 n495 ; n1740
g1677 and n1739 n1740 ; n1741
g1678 and n1738 n1741 ; n1742
g1679 and n1737 n1742 ; n1743
g1680 and n1372 n1743 ; n1744
g1681 and n1735 n1744 ; n1745
g1682 and n1731 n1745 ; n1746
g1683 and n1726 n1746 ; n1747
g1684 and n227 n1747 ; n1748
g1685 and n330_not n1748 ; n1749
g1686 and n426_not n1749 ; n1750
g1687 and n171_not n1750 ; n1751
g1688 and n1101_not n1751 ; n1752
g1689 and n177_not n1752 ; n1753
g1690 and n567_not n1753 ; n1754
g1691 nor n233 n752 ; n1755
g1692 and n144_not n1755 ; n1756
g1693 and n791_not n1756 ; n1757
g1694 and n672_not n1757 ; n1758
g1695 and n655_not n1758 ; n1759
g1696 nor n232 n278 ; n1760
g1697 nor n424 n689 ; n1761
g1698 and n469_not n1761 ; n1762
g1699 and n224_not n1762 ; n1763
g1700 and n1760 n1763 ; n1764
g1701 and n694 n1764 ; n1765
g1702 and n1759 n1765 ; n1766
g1703 and n1754 n1766 ; n1767
g1704 and n774 n1767 ; n1768
g1705 and n1725 n1768 ; n1769
g1706 and n1719 n1769 ; n1770
g1707 and n1182 n1770 ; n1771
g1708 and n590 n1771 ; n1772
g1709 and n135_not n1772 ; n1773
g1710 and n400_not n1773 ; n1774
g1711 and n563_not n1774 ; n1775
g1712 and n504_not n1775 ; n1776
g1713 and n164_not n1776 ; n1777
g1714 and n325_not n1777 ; n1778
g1715 and n875_not n1778 ; n1779
g1716 nor n1665 n1779 ; n1780
g1717 nor n655 n825 ; n1781
g1718 nor n189 n592 ; n1782
g1719 nor n154 n299 ; n1783
g1720 and n1102_not n1783 ; n1784
g1721 nor n163 n1203 ; n1785
g1722 and n1784 n1785 ; n1786
g1723 and n896 n1786 ; n1787
g1724 and n1782 n1787 ; n1788
g1725 and n506_not n1788 ; n1789
g1726 and n1755 n1789 ; n1790
g1727 and n460_not n1790 ; n1791
g1728 and n527_not n1791 ; n1792
g1729 and n331_not n1792 ; n1793
g1730 and n689_not n1793 ; n1794
g1731 nor n352 n514 ; n1795
g1732 and n223_not n1795 ; n1796
g1733 and n513_not n1796 ; n1797
g1734 and n363_not n1797 ; n1798
g1735 nor n335 n619 ; n1799
g1736 and n438_not n1799 ; n1800
g1737 and n1408 n1800 ; n1801
g1738 and n494 n1801 ; n1802
g1739 and n1798 n1802 ; n1803
g1740 and n1020 n1803 ; n1804
g1741 and n515 n1804 ; n1805
g1742 and n193 n1805 ; n1806
g1743 and n136_not n1806 ; n1807
g1744 and n171_not n1807 ; n1808
g1745 and n417_not n1808 ; n1809
g1746 and n296_not n1809 ; n1810
g1747 and n274_not n1810 ; n1811
g1748 and n372_not n1811 ; n1812
g1749 and n886_not n1812 ; n1813
g1750 and n188_not n1813 ; n1814
g1751 nor n469 n641 ; n1815
g1752 and n203_not n1815 ; n1816
g1753 and n305_not n1816 ; n1817
g1754 and n271_not n1817 ; n1818
g1755 and n875_not n1818 ; n1819
g1756 and n454 n508 ; n1820
g1757 and n563_not n1820 ; n1821
g1758 and n1104_not n1821 ; n1822
g1759 and n95_not n1822 ; n1823
g1760 nor n125 n158 ; n1824
g1761 nor n403 n602 ; n1825
g1762 nor n231 n504 ; n1826
g1763 nor n466 n777 ; n1827
g1764 nor n226 n1101 ; n1828
g1765 and n1667 n1828 ; n1829
g1766 and n1827 n1829 ; n1830
g1767 and n591 n1830 ; n1831
g1768 and n1062_not n1831 ; n1832
g1769 and n290_not n1832 ; n1833
g1770 and n505_not n1833 ; n1834
g1771 and n531_not n1834 ; n1835
g1772 and n371_not n1835 ; n1836
g1773 and n569_not n1836 ; n1837
g1774 and n337_not n1837 ; n1838
g1775 nor n121 n536 ; n1839
g1776 and n962 n1839 ; n1840
g1777 and n355_not n1840 ; n1841
g1778 and n150_not n1841 ; n1842
g1779 and n419_not n1842 ; n1843
g1780 and n603_not n1843 ; n1844
g1781 and n1838 n1844 ; n1845
g1782 and n1826 n1845 ; n1846
g1783 and n520 n1846 ; n1847
g1784 and n1576 n1847 ; n1848
g1785 and n826 n1848 ; n1849
g1786 and n1825 n1849 ; n1850
g1787 and n1824 n1850 ; n1851
g1788 and n847_not n1851 ; n1852
g1789 and n329_not n1852 ; n1853
g1790 and n803_not n1853 ; n1854
g1791 and n571_not n1854 ; n1855
g1792 and n495_not n1855 ; n1856
g1793 and n200_not n1856 ; n1857
g1794 and n639_not n1857 ; n1858
g1795 and n492_not n1858 ; n1859
g1796 nor n229 n367 ; n1860
g1797 and n474_not n1860 ; n1861
g1798 and n1859 n1861 ; n1862
g1799 and n776 n1862 ; n1863
g1800 and n1823 n1863 ; n1864
g1801 and n1819 n1864 ; n1865
g1802 and n1814 n1865 ; n1866
g1803 and n1794 n1866 ; n1867
g1804 and n1531 n1867 ; n1868
g1805 and n1781 n1868 ; n1869
g1806 and n533 n1869 ; n1870
g1807 and n282 n1870 ; n1871
g1808 and n399 n1871 ; n1872
g1809 and n1040 n1872 ; n1873
g1810 and n152_not n1873 ; n1874
g1811 and n239_not n1874 ; n1875
g1812 and n287_not n1875 ; n1876
g1813 and n251_not n1876 ; n1877
g1814 nor n1779 n1877 ; n1878
g1815 nor n165 n452 ; n1879
g1816 and n1438 n1879 ; n1880
g1817 and n1247 n1880 ; n1881
g1818 and n398_not n1881 ; n1882
g1819 and n99_not n1882 ; n1883
g1820 and n712_not n1883 ; n1884
g1821 nor n278 n809 ; n1885
g1822 and n884_not n1885 ; n1886
g1823 and n245_not n1886 ; n1887
g1824 and n777_not n1887 ; n1888
g1825 and n283_not n1888 ; n1889
g1826 and n127_not n1889 ; n1890
g1827 nor n136 n287 ; n1891
g1828 and n298_not n1891 ; n1892
g1829 and n201_not n1892 ; n1893
g1830 nor n280 n667 ; n1894
g1831 and n618 n1894 ; n1895
g1832 and n147_not n1895 ; n1896
g1833 nor n158 n511 ; n1897
g1834 and n293_not n1897 ; n1898
g1835 and n1896 n1898 ; n1899
g1836 and n1697 n1899 ; n1900
g1837 and n1345 n1900 ; n1901
g1838 and n1211 n1901 ; n1902
g1839 and n1039 n1902 ; n1903
g1840 and n1601 n1903 ; n1904
g1841 and n1476 n1904 ; n1905
g1842 and n1893 n1905 ; n1906
g1843 and n1890 n1906 ; n1907
g1844 and n1884 n1907 ; n1908
g1845 and n1102_not n1908 ; n1909
g1846 and n594_not n1909 ; n1910
g1847 and n419_not n1910 ; n1911
g1848 and n715_not n1911 ; n1912
g1849 and n592_not n1912 ; n1913
g1850 nor n1877 n1913 ; n1914
g1851 nor n224 n531 ; n1915
g1852 nor n239 n527 ; n1916
g1853 nor n571 n623 ; n1917
g1854 nor n713 n1072 ; n1918
g1855 and n329_not n1918 ; n1919
g1856 and n809_not n1919 ; n1920
g1857 and n302_not n1920 ; n1921
g1858 and n716_not n1921 ; n1922
g1859 and n132_not n1922 ; n1923
g1860 and n252_not n1923 ; n1924
g1861 and n304_not n1924 ; n1925
g1862 nor n232 n752 ; n1926
g1863 and n1102_not n1926 ; n1927
g1864 and n673_not n1927 ; n1928
g1865 and n244 n426_not ; n1929
g1866 and n461_not n1929 ; n1930
g1867 and n372_not n1930 ; n1931
g1868 and n1557 n1931 ; n1932
g1869 and n874 n1932 ; n1933
g1870 and n1426 n1933 ; n1934
g1871 and n641_not n1934 ; n1935
g1872 and n514_not n1935 ; n1936
g1873 and n339_not n1936 ; n1937
g1874 and n273_not n1937 ; n1938
g1875 and n277_not n1938 ; n1939
g1876 and n325_not n1939 ; n1940
g1877 nor n301 n884 ; n1941
g1878 and n374_not n1941 ; n1942
g1879 nor n130 n299 ; n1943
g1880 and n1104_not n1943 ; n1944
g1881 and n989 n1944 ; n1945
g1882 and n1942 n1945 ; n1946
g1883 and n1940 n1946 ; n1947
g1884 and n1928 n1947 ; n1948
g1885 and n977 n1948 ; n1949
g1886 and n538 n1949 ; n1950
g1887 and n118_not n1950 ; n1951
g1888 and n240_not n1951 ; n1952
g1889 and n283_not n1952 ; n1953
g1890 and n791_not n1953 ; n1954
g1891 and n1203_not n1954 ; n1955
g1892 and n1010_not n1955 ; n1956
g1893 and n81_not n1956 ; n1957
g1894 and n222_not n1957 ; n1958
g1895 nor n469 n639 ; n1959
g1896 and n119_not n1959 ; n1960
g1897 and n772 n1960 ; n1961
g1898 and n512 n1961 ; n1962
g1899 and n1183 n1962 ; n1963
g1900 and n896 n1963 ; n1964
g1901 and n617_not n1964 ; n1965
g1902 and n367_not n1965 ; n1966
g1903 and n395_not n1966 ; n1967
g1904 and n525_not n1967 ; n1968
g1905 and n358_not n1968 ; n1969
g1906 and n121_not n221 ; n1970
g1907 and n493_not n1970 ; n1971
g1908 and n418 n1248 ; n1972
g1909 and n95_not n1972 ; n1973
g1910 and n1971 n1973 ; n1974
g1911 and n658 n1974 ; n1975
g1912 and n877 n1975 ; n1976
g1913 and n1969 n1976 ; n1977
g1914 and n1958 n1977 ; n1978
g1915 and n1925 n1978 ; n1979
g1916 and n1917 n1979 ; n1980
g1917 and n1916 n1980 ; n1981
g1918 and n1915 n1981 ; n1982
g1919 and n515 n1982 ; n1983
g1920 and n1574 n1983 ; n1984
g1921 and n558_not n1984 ; n1985
g1922 and n280_not n1985 ; n1986
g1923 and n416_not n1986 ; n1987
g1924 and n296_not n1987 ; n1988
g1925 and n505_not n1988 ; n1989
g1926 and n424_not n1989 ; n1990
g1927 and n293_not n1990 ; n1991
g1928 and n270_not n1991 ; n1992
g1929 nor n1913 n1992 ; n1993
g1930 nor n302 n1102 ; n1994
g1931 nor n168 n397 ; n1995
g1932 and n589_not n1995 ; n1996
g1933 and n1898 n1996 ; n1997
g1934 and n793 n1997 ; n1998
g1935 and n297 n1998 ; n1999
g1936 and n1994 n1999 ; n2000
g1937 and n1101_not n2000 ; n2001
g1938 and n205_not n2001 ; n2002
g1939 and n191_not n2002 ; n2003
g1940 and n1127_not n2003 ; n2004
g1941 and n489_not n2004 ; n2005
g1942 and n875_not n2005 ; n2006
g1943 nor n492 n537 ; n2007
g1944 and n667_not n2007 ; n2008
g1945 and n460_not n2008 ; n2009
g1946 and n130_not n2009 ; n2010
g1947 and n336 n979 ; n2011
g1948 and n372_not n2011 ; n2012
g1949 nor n340 n1011 ; n2013
g1950 nor n165 n240 ; n2014
g1951 and n2013 n2014 ; n2015
g1952 and n1105 n2015 ; n2016
g1953 and n453_not n2016 ; n2017
g1954 nor n355 n509 ; n2018
g1955 and n147_not n2018 ; n2019
g1956 and n371_not n2019 ; n2020
g1957 nor n163 n716 ; n2021
g1958 nor n95 n746 ; n2022
g1959 nor n206 n364 ; n2023
g1960 and n422_not n2023 ; n2024
g1961 and n366_not n2024 ; n2025
g1962 nor n222 n438 ; n2026
g1963 and n1329 n2026 ; n2027
g1964 and n529 n2027 ; n2028
g1965 and n2025 n2028 ; n2029
g1966 and n1691 n2029 ; n2030
g1967 and n2022 n2030 ; n2031
g1968 and n2021 n2031 ; n2032
g1969 and n1330 n2032 ; n2033
g1970 and n1668 n2033 ; n2034
g1971 and n1009 n2034 ; n2035
g1972 and n619_not n2035 ; n2036
g1973 and n192_not n2036 ; n2037
g1974 and n468_not n2037 ; n2038
g1975 and n436_not n2038 ; n2039
g1976 and n569_not n2039 ; n2040
g1977 and n2020 n2040 ; n2041
g1978 and n2017 n2041 ; n2042
g1979 and n1600 n2042 ; n2043
g1980 and n2012 n2043 ; n2044
g1981 and n1183 n2044 ; n2045
g1982 and n2010 n2045 ; n2046
g1983 and n2006 n2046 ; n2047
g1984 and n720 n2047 ; n2048
g1985 and n558_not n2048 ; n2049
g1986 and n284_not n2049 ; n2050
g1987 and n203_not n2050 ; n2051
g1988 and n1795 n2051 ; n2052
g1989 and n290_not n2052 ; n2053
g1990 and n102_not n2053 ; n2054
g1991 and n424_not n2054 ; n2055
g1992 and n470_not n2055 ; n2056
g1993 and n562_not n2056 ; n2057
g1994 nor n1992 n2057 ; n2058
g1995 nor n152 n190 ; n2059
g1996 and n735 n2059 ; n2060
g1997 and n591 n2060 ; n2061
g1998 and n232_not n2061 ; n2062
g1999 and n809_not n2062 ; n2063
g2000 and n496_not n2063 ; n2064
g2001 and n144_not n2064 ; n2065
g2002 and n298_not n2065 ; n2066
g2003 and n337_not n2066 ; n2067
g2004 and n633_not n2067 ; n2068
g2005 and n1248 n1252 ; n2069
g2006 and n289_not n2069 ; n2070
g2007 and n255_not n2070 ; n2071
g2008 and n489_not n2071 ; n2072
g2009 nor n169 n637 ; n2073
g2010 and n248_not n2073 ; n2074
g2011 and n1104_not n2074 ; n2075
g2012 and n1784 n2075 ; n2076
g2013 and n812 n2076 ; n2077
g2014 and n1132 n2077 ; n2078
g2015 and n207 n2078 ; n2079
g2016 and n1085 n2079 ; n2080
g2017 and n918 n2080 ; n2081
g2018 and n2072 n2081 ; n2082
g2019 and n2068 n2082 ; n2083
g2020 and n515 n2083 ; n2084
g2021 and n557_not n2084 ; n2085
g2022 and n419_not n2085 ; n2086
g2023 and n396_not n2086 ; n2087
g2024 and n601_not n2087 ; n2088
g2025 and n364_not n1129 ; n2089
g2026 nor n142 n641 ; n2090
g2027 nor n363 n558 ; n2091
g2028 nor n167 n506 ; n2092
g2029 nor n99 n223 ; n2093
g2030 and n2092 n2093 ; n2094
g2031 and n2091 n2094 ; n2095
g2032 and n2090 n2095 ; n2096
g2033 and n2089 n2096 ; n2097
g2034 and n329_not n2097 ; n2098
g2035 and n150_not n2098 ; n2099
g2036 and n884_not n2099 ; n2100
g2037 and n164_not n2100 ; n2101
g2038 and n372_not n2101 ; n2102
g2039 and n393_not n2102 ; n2103
g2040 and n525_not n2103 ; n2104
g2041 nor n514 n713 ; n2105
g2042 nor n229 n667 ; n2106
g2043 and n426_not n2106 ; n2107
g2044 and n602_not n2107 ; n2108
g2045 and n115_not n2108 ; n2109
g2046 and n334_not n2109 ; n2110
g2047 and n246_not n2110 ; n2111
g2048 and n170_not n2111 ; n2112
g2049 nor n226 n509 ; n2113
g2050 and n1072_not n1128 ; n2114
g2051 and n146_not n2114 ; n2115
g2052 and n2113 n2115 ; n2116
g2053 and n1643 n2116 ; n2117
g2054 and n1879 n2117 ; n2118
g2055 and n1012 n2118 ; n2119
g2056 and n2112 n2119 ; n2120
g2057 and n2021 n2120 ; n2121
g2058 and n1063 n2121 ; n2122
g2059 and n108 n2122 ; n2123
g2060 and n203_not n2123 ; n2124
g2061 and n2105 n2124 ; n2125
g2062 and n594_not n2125 ; n2126
g2063 and n287_not n2126 ; n2127
g2064 nor n397 n527 ; n2128
g2065 and n245_not n2128 ; n2129
g2066 and n567_not n2129 ; n2130
g2067 and n623_not n2130 ; n2131
g2068 and n338_not n2131 ; n2132
g2069 nor n513 n1062 ; n2133
g2070 and n475 n2013 ; n2134
g2071 and n2133 n2134 ; n2135
g2072 and n2132 n2135 ; n2136
g2073 and n2127 n2136 ; n2137
g2074 and n2104 n2137 ; n2138
g2075 and n1251 n2138 ; n2139
g2076 and n120 n2139 ; n2140
g2077 and n2088 n2140 ; n2141
g2078 and n356 n2141 ; n2142
g2079 and n518_not n2142 ; n2143
g2080 and n151_not n2143 ; n2144
g2081 and n155_not n2144 ; n2145
g2082 and n435_not n2145 ; n2146
g2083 and n461_not n2146 ; n2147
g2084 and n326_not n2147 ; n2148
g2085 and n368_not n2148 ; n2149
g2086 and n130_not n2149 ; n2150
g2087 and n569_not n2150 ; n2151
g2088 and n655_not n2151 ; n2152
g2089 nor n2057 n2152 ; n2153
g2090 nor n118 n1072 ; n2154
g2091 and n1328 n2154 ; n2155
g2092 and n1890 n2155 ; n2156
g2093 and n1379 n2156 ; n2157
g2094 and n1128 n2157 ; n2158
g2095 and n2073 n2158 ; n2159
g2096 and n341 n2159 ; n2160
g2097 and n194_not n2160 ; n2161
g2098 and n1246_not n2161 ; n2162
g2099 and n803_not n2162 ; n2163
g2100 and n435_not n2163 ; n2164
g2101 and n357_not n2164 ; n2165
g2102 and n142_not n2165 ; n2166
g2103 and n271_not n2166 ; n2167
g2104 nor n492 n514 ; n2168
g2105 and n525_not n2168 ; n2169
g2106 nor n393 n980 ; n2170
g2107 and n356 n2170 ; n2171
g2108 and n460_not n2171 ; n2172
g2109 and n156 n1893 ; n2173
g2110 and n175_not n2173 ; n2174
g2111 and n747 n773 ; n2175
g2112 and n1141 n2175 ; n2176
g2113 and n1456 n2176 ; n2177
g2114 and n2174 n2177 ; n2178
g2115 and n2172 n2178 ; n2179
g2116 and n757 n2179 ; n2180
g2117 and n671 n2180 ; n2181
g2118 and n2169 n2181 ; n2182
g2119 and n1668 n2182 ; n2183
g2120 and n423 n2183 ; n2184
g2121 and n2167 n2184 ; n2185
g2122 and n1247 n2185 ; n2186
g2123 and n508 n2186 ; n2187
g2124 and n713_not n2187 ; n2188
g2125 and n243_not n2188 ; n2189
g2126 nor n2152 n2189 ; n2190
g2127 nor n157 n276 ; n2191
g2128 nor n144 n1101 ; n2192
g2129 and n2191 n2192 ; n2193
g2130 and n2154 n2193 ; n2194
g2131 and n1825 n2194 ; n2195
g2132 and n1550 n2195 ; n2196
g2133 and n2073 n2196 ; n2197
g2134 and n190_not n2197 ; n2198
g2135 and n278_not n2198 ; n2199
g2136 and n121_not n2199 ; n2200
g2137 and n275_not n2200 ; n2201
g2138 and n173_not n2201 ; n2202
g2139 and n720 n1531 ; n2203
g2140 and n504_not n2203 ; n2204
g2141 and n271_not n2204 ; n2205
g2142 and n95_not n2205 ; n2206
g2143 and n886_not n2206 ; n2207
g2144 and n358_not n2207 ; n2208
g2145 nor n714 n961 ; n2209
g2146 nor n147 n192 ; n2210
g2147 and n2209 n2210 ; n2211
g2148 and n887 n2211 ; n2212
g2149 and n281_not n2212 ; n2213
g2150 and n557_not n2213 ; n2214
g2151 and n571_not n2214 ; n2215
g2152 and n228_not n2215 ; n2216
g2153 and n716_not n2216 ; n2217
g2154 nor n194 n619 ; n2218
g2155 and n825_not n2218 ; n2219
g2156 nor n273 n506 ; n2220
g2157 and n595 n2220 ; n2221
g2158 and n2093 n2221 ; n2222
g2159 and n1069 n2222 ; n2223
g2160 and n354_not n2223 ; n2224
g2161 and n803_not n2224 ; n2225
g2162 and n367_not n2225 ; n2226
g2163 and n146_not n2226 ; n2227
g2164 and n286_not n2227 ; n2228
g2165 and n245_not n2228 ; n2229
g2166 nor n236 n460 ; n2230
g2167 and n133 n2230 ; n2231
g2168 and n1942 n2231 ; n2232
g2169 and n752_not n2232 ; n2233
g2170 and n189_not n2233 ; n2234
g2171 and n417_not n2234 ; n2235
g2172 and n453_not n2235 ; n2236
g2173 and n394_not n2236 ; n2237
g2174 nor n352 n420 ; n2238
g2175 and n505_not n2238 ; n2239
g2176 and n163_not n2239 ; n2240
g2177 nor n107 n563 ; n2241
g2178 and n1763 n2241 ; n2242
g2179 and n2240 n2242 ; n2243
g2180 and n2237 n2243 ; n2244
g2181 and n808 n2244 ; n2245
g2182 and n2229 n2245 ; n2246
g2183 and n1994 n2246 ; n2247
g2184 and n2219 n2247 ; n2248
g2185 and n116 n2248 ; n2249
g2186 and n1389 n2249 ; n2250
g2187 and n136_not n2250 ; n2251
g2188 and n713_not n2251 ; n2252
g2189 and n641_not n2252 ; n2253
g2190 and n292_not n2253 ; n2254
g2191 and n396_not n2254 ; n2255
g2192 and n248_not n2255 ; n2256
g2193 and n290_not n2256 ; n2257
g2194 and n567_not n2257 ; n2258
g2195 and n618 n1827 ; n2259
g2196 and n239_not n2259 ; n2260
g2197 and n513_not n2260 ; n2261
g2198 and n429_not n2261 ; n2262
g2199 nor n746 n809 ; n2263
g2200 and n161_not n202 ; n2264
g2201 and n672_not n2264 ; n2265
g2202 and n526 n732 ; n2266
g2203 and n237_not n2266 ; n2267
g2204 and n2265 n2267 ; n2268
g2205 and n535 n2268 ; n2269
g2206 and n1155 n2269 ; n2270
g2207 and n623_not n2270 ; n2271
g2208 and n712_not n2271 ; n2272
g2209 and n436_not n2272 ; n2273
g2210 and n225_not n2273 ; n2274
g2211 and n158_not n2274 ; n2275
g2212 nor n496 n601 ; n2276
g2213 and n152_not n2276 ; n2277
g2214 and n357_not n2277 ; n2278
g2215 and n2275 n2278 ; n2279
g2216 and n365 n2279 ; n2280
g2217 and n2263 n2280 ; n2281
g2218 and n2262 n2281 ; n2282
g2219 and n1268 n2282 ; n2283
g2220 and n2258 n2283 ; n2284
g2221 and n2217 n2284 ; n2285
g2222 and n2208 n2285 ; n2286
g2223 and n2202 n2286 ; n2287
g2224 and n510 n2287 ; n2288
g2225 and n355_not n2288 ; n2289
g2226 and n255_not n2289 ; n2290
g2227 and n620_not n2290 ; n2291
g2228 nor n2189 n2291 ; n2292
g2229 nor n243 n367 ; n2293
g2230 and n228_not n2293 ; n2294
g2231 and n537_not n2294 ; n2295
g2232 and n470_not n2295 ; n2296
g2233 nor n146 n460 ; n2297
g2234 and n827 n2297 ; n2298
g2235 and n847_not n2298 ; n2299
g2236 and n150_not n2299 ; n2300
g2237 and n290_not n2300 ; n2301
g2238 and n1131 n1476 ; n2302
g2239 and n746_not n2302 ; n2303
g2240 and n1025 n2303 ; n2304
g2241 and n1533 n2304 ; n2305
g2242 and n816 n2305 ; n2306
g2243 and n207 n2306 ; n2307
g2244 and n2091 n2307 ; n2308
g2245 and n2301 n2308 ; n2309
g2246 and n2296 n2309 ; n2310
g2247 and n2169 n2310 ; n2311
g2248 and n1825 n2311 ; n2312
g2249 and n229_not n2312 ; n2313
g2250 and n777_not n2313 ; n2314
g2251 and n287_not n2314 ; n2315
g2252 and n603_not n2315 ; n2316
g2253 and n1104_not n2316 ; n2317
g2254 nor n171 n354 ; n2318
g2255 and n280_not n2318 ; n2319
g2256 and n275_not n2319 ; n2320
g2257 and n292_not n2320 ; n2321
g2258 and n416_not n2321 ; n2322
g2259 and n192_not n2322 ; n2323
g2260 and n164_not n2323 ; n2324
g2261 and n567_not n2324 ; n2325
g2262 and n301_not n437 ; n2326
g2263 and n339_not n2326 ; n2327
g2264 and n357_not n2327 ; n2328
g2265 and n657_not n2328 ; n2329
g2266 and n188_not n2329 ; n2330
g2267 nor n601 n667 ; n2331
g2268 and n337_not n2331 ; n2332
g2269 nor n167 n331 ; n2333
g2270 and n252_not n2333 ; n2334
g2271 and n887 n2334 ; n2335
g2272 and n2332 n2335 ; n2336
g2273 and n632 n2336 ; n2337
g2274 and n2330 n2337 ; n2338
g2275 and n238 n2338 ; n2339
g2276 and n2325 n2339 ; n2340
g2277 and n896 n2340 ; n2341
g2278 and n420_not n2341 ; n2342
g2279 and n353_not n2342 ; n2343
g2280 and n155_not n2343 ; n2344
g2281 and n1127_not n2344 ; n2345
g2282 nor n563 n673 ; n2346
g2283 and n175_not n2346 ; n2347
g2284 nor n468 n961 ; n2348
g2285 nor n589 n1246 ; n2349
g2286 and n1636 n1739 ; n2350
g2287 and n2349 n2350 ; n2351
g2288 and n2348 n2351 ; n2352
g2289 and n241 n2352 ; n2353
g2290 and n1102_not n2353 ; n2354
g2291 and n2347 n2354 ; n2355
g2292 and n327_not n2355 ; n2356
g2293 and n594_not n2356 ; n2357
g2294 and n430_not n2357 ; n2358
g2295 and n1203_not n2358 ; n2359
g2296 and n474_not n2359 ; n2360
g2297 nor n302 n532 ; n2361
g2298 nor n91 n518 ; n2362
g2299 and n142_not n2362 ; n2363
g2300 and n2361 n2363 ; n2364
g2301 and n281_not n2364 ; n2365
g2302 and n147_not n2365 ; n2366
g2303 and n791_not n2366 ; n2367
g2304 and n493_not n2367 ; n2368
g2305 and n358_not n2368 ; n2369
g2306 and n875_not n2369 ; n2370
g2307 nor n328 n569 ; n2371
g2308 and n793 n1839 ; n2372
g2309 and n308 n2372 ; n2373
g2310 and n2371 n2373 ; n2374
g2311 and n2370 n2374 ; n2375
g2312 and n2360 n2375 ; n2376
g2313 and n2345 n2376 ; n2377
g2314 and n2317 n2377 ; n2378
g2315 and n1667 n2378 ; n2379
g2316 and n937 n2379 ; n2380
g2317 and n1252 n2380 ; n2381
g2318 and n462_not n2381 ; n2382
g2319 and n1021 n2382 ; n2383
g2320 and n715_not n2383 ; n2384
g2321 and n157_not n2384 ; n2385
g2322 and n325_not n2385 ; n2386
g2323 and n886_not n2386 ; n2387
g2324 and n231_not n2387 ; n2388
g2325 nor n2291 n2388 ; n2389
g2326 nor n173 n564 ; n2390
g2327 and n362 n2390 ; n2391
g2328 and n1879 n2391 ; n2392
g2329 and n1380 n2392 ; n2393
g2330 and n1761 n2393 ; n2394
g2331 and n123_not n2394 ; n2395
g2332 and n1108 n2395 ; n2396
g2333 and n511_not n2396 ; n2397
g2334 and n118_not n2397 ; n2398
g2335 and n417_not n2398 ; n2399
g2336 and n290_not n2399 ; n2400
g2337 and n777_not n2400 ; n2401
g2338 and n537_not n2401 ; n2402
g2339 and n200_not n2402 ; n2403
g2340 and n272_not n2403 ; n2404
g2341 and n1127_not n2404 ; n2405
g2342 nor n99 n451 ; n2406
g2343 nor n273 n292 ; n2407
g2344 and n883_not n2407 ; n2408
g2345 and n428_not n2408 ; n2409
g2346 nor n147 n271 ; n2410
g2347 and n1324 n2410 ; n2411
g2348 and n639_not n2411 ; n2412
g2349 and n825_not n2412 ; n2413
g2350 and n145_not n2413 ; n2414
g2351 and n240_not n2414 ; n2415
g2352 and n372_not n2415 ; n2416
g2353 and n589_not n2416 ; n2417
g2354 nor n637 n1102 ; n2418
g2355 and n205_not n2418 ; n2419
g2356 and n1203_not n2419 ; n2420
g2357 and n470_not n2420 ; n2421
g2358 and n592_not n2421 ; n2422
g2359 nor n119 n142 ; n2423
g2360 nor n223 n419 ; n2424
g2361 nor n248 n1062 ; n2425
g2362 and n368_not n2425 ; n2426
g2363 and n156 n932_not ; n2427
g2364 and n2426 n2427 ; n2428
g2365 and n2424 n2428 ; n2429
g2366 and n2423 n2429 ; n2430
g2367 and n2422 n2430 ; n2431
g2368 and n1131 n2431 ; n2432
g2369 and n2417 n2432 ; n2433
g2370 and n1247 n2433 ; n2434
g2371 and n236_not n2434 ; n2435
g2372 and n242_not n2435 ; n2436
g2373 and n284_not n2436 ; n2437
g2374 and n130_not n2437 ; n2438
g2375 and n449_not n2438 ; n2439
g2376 and n288 n2439 ; n2440
g2377 and n429_not n2440 ; n2441
g2378 nor n301 n712 ; n2442
g2379 and n791_not n2442 ; n2443
g2380 and n425_not n2443 ; n2444
g2381 and n657_not n2444 ; n2445
g2382 and n2441 n2445 ; n2446
g2383 and n2409 n2446 ; n2447
g2384 and n790 n2447 ; n2448
g2385 and n2040 n2448 ; n2449
g2386 and n665 n2449 ; n2450
g2387 and n604 n2450 ; n2451
g2388 and n2406 n2451 ; n2452
g2389 and n1667 n2452 ; n2453
g2390 and n399 n2453 ; n2454
g2391 and n2068 n2454 ; n2455
g2392 and n2405 n2455 ; n2456
g2393 and n713_not n2456 ; n2457
g2394 and n233_not n2457 ; n2458
g2395 and n461_not n2458 ; n2459
g2396 and n157_not n2459 ; n2460
g2397 and n623_not n2460 ; n2461
g2398 and n338_not n2461 ; n2462
g2399 and n532_not n2462 ; n2463
g2400 and n666_not n2463 ; n2464
g2401 nor n2388 n2464 ; n2465
g2402 nor n255 n617 ; n2466
g2403 nor n305 n451 ; n2467
g2404 nor n366 n689 ; n2468
g2405 and n202 n495_not ; n2469
g2406 and n252_not n2469 ; n2470
g2407 and n990 n2470 ; n2471
g2408 and n899 n2471 ; n2472
g2409 and n2468 n2472 ; n2473
g2410 and n2348 n2473 ; n2474
g2411 and n2467 n2474 ; n2475
g2412 and n193 n2475 ; n2476
g2413 and n2466 n2476 ; n2477
g2414 and n396_not n2477 ; n2478
g2415 and n290_not n2478 ; n2479
g2416 and n283_not n2479 ; n2480
g2417 and n525_not n2480 ; n2481
g2418 and n158_not n2481 ; n2482
g2419 and n655_not n2482 ; n2483
g2420 nor n167 n430 ; n2484
g2421 nor n490 n514 ; n2485
g2422 and n374_not n2485 ; n2486
g2423 and n603_not n2486 ; n2487
g2424 and n365 n1204 ; n2488
g2425 and n300 n2488 ; n2489
g2426 and n2487 n2489 ; n2490
g2427 and n1915 n2490 ; n2491
g2428 and n621 n2491 ; n2492
g2429 and n896 n2492 ; n2493
g2430 and n885 n2493 ; n2494
g2431 and n1072_not n2494 ; n2495
g2432 and n111_not n2495 ; n2496
g2433 and n809_not n2496 ; n2497
g2434 and n121_not n2497 ; n2498
g2435 and n1010_not n2498 ; n2499
g2436 and n771_not n2499 ; n2500
g2437 nor n460 n594 ; n2501
g2438 and n206_not n2501 ; n2502
g2439 and n243_not n2502 ; n2503
g2440 and n657_not n2503 ; n2504
g2441 and n161_not n2504 ; n2505
g2442 and n672_not n2505 ; n2506
g2443 nor n163 n1246 ; n2507
g2444 nor n420 n504 ; n2508
g2445 and n642 n2508 ; n2509
g2446 and n435_not n2509 ; n2510
g2447 and n292_not n2510 ; n2511
g2448 and n519_not n2511 ; n2512
g2449 and n232_not n282 ; n2513
g2450 and n713_not n2513 ; n2514
g2451 and n231_not n2514 ; n2515
g2452 and n351 n2515 ; n2516
g2453 and n2512 n2516 ; n2517
g2454 and n2507 n2517 ; n2518
g2455 and n2439 n2518 ; n2519
g2456 and n2506 n2519 ; n2520
g2457 and n2500 n2520 ; n2521
g2458 and n2484 n2521 ; n2522
g2459 and n720 n2522 ; n2523
g2460 and n2483 n2523 ; n2524
g2461 and n189_not n2524 ; n2525
g2462 and n239_not n2525 ; n2526
g2463 and n417_not n2526 ; n2527
g2464 and n226_not n2527 ; n2528
g2465 and n438_not n2528 ; n2529
g2466 and n563_not n2529 ; n2530
g2467 and n791_not n2530 ; n2531
g2468 and n295_not n2531 ; n2532
g2469 and n293_not n2532 ; n2533
g2470 nor n2464 n2533 ; n2534
g2471 nor n248 n327 ; n2535
g2472 and n91_not n2535 ; n2536
g2473 and n273_not n2536 ; n2537
g2474 and n624 n2537 ; n2538
g2475 and n961_not n2538 ; n2539
g2476 and n130_not n2539 ; n2540
g2477 and n225_not n2540 ; n2541
g2478 and n252_not n2541 ; n2542
g2479 and n95_not n2542 ; n2543
g2480 nor n398 n594 ; n2544
g2481 nor n242 n505 ; n2545
g2482 and n157_not n2545 ; n2546
g2483 and n2427 n2546 ; n2547
g2484 and n2544 n2547 ; n2548
g2485 and n2170 n2548 ; n2549
g2486 and n255_not n2549 ; n2550
g2487 and n619_not n2550 ; n2551
g2488 and n287_not n2551 ; n2552
g2489 and n306_not n2552 ; n2553
g2490 and n371_not n2553 ; n2554
g2491 and n231_not n2554 ; n2555
g2492 nor n239 n633 ; n2556
g2493 and n638 n2556 ; n2557
g2494 and n989 n2557 ; n2558
g2495 and n1879 n2558 ; n2559
g2496 and n844 n2559 ; n2560
g2497 and n1202 n2560 ; n2561
g2498 and n2555 n2561 ; n2562
g2499 and n2543 n2562 ; n2563
g2500 and n1379 n2563 ; n2564
g2501 and n1389 n2564 ; n2565
g2502 and n397_not n2565 ; n2566
g2503 and n752_not n2566 ; n2567
g2504 and n334_not n2567 ; n2568
g2505 and n107_not n2568 ; n2569
g2506 and n716_not n2569 ; n2570
g2507 and n569_not n2570 ; n2571
g2508 nor n2533 n2571 ; n2572
g2509 nor n325 n883 ; n2573
g2510 nor n427 n617 ; n2574
g2511 and n254_not n2574 ; n2575
g2512 and n803_not n2575 ; n2576
g2513 and n228_not n2576 ; n2577
g2514 and n191_not n2577 ; n2578
g2515 and n283_not n2578 ; n2579
g2516 and n366_not n2579 ; n2580
g2517 and n489_not n2580 ; n2581
g2518 nor n363 n875 ; n2582
g2519 nor n509 n623 ; n2583
g2520 nor n398 n468 ; n2584
g2521 and n2090 n2584 ; n2585
g2522 and n847_not n2585 ; n2586
g2523 and n175_not n2586 ; n2587
g2524 and n223_not n2587 ; n2588
g2525 and n568_not n2588 ; n2589
g2526 and n340_not n2589 ; n2590
g2527 and n1127_not n2590 ; n2591
g2528 nor n240 n245 ; n2592
g2529 and n1203_not n2592 ; n2593
g2530 and n873 n1180 ; n2594
g2531 and n95_not n2594 ; n2595
g2532 and n2593 n2595 ; n2596
g2533 and n2349 n2596 ; n2597
g2534 and n1839 n2597 ; n2598
g2535 and n977 n2598 ; n2599
g2536 and n115_not n2599 ; n2600
g2537 and n514_not n2600 ; n2601
g2538 and n435_not n2601 ; n2602
g2539 and n225_not n2602 ; n2603
g2540 and n532_not n2603 ; n2604
g2541 and n81_not n2604 ; n2605
g2542 nor n169 n537 ; n2606
g2543 and n525_not n2606 ; n2607
g2544 nor n461 n504 ; n2608
g2545 and n1800 n2608 ; n2609
g2546 and n2607 n2609 ; n2610
g2547 and n595 n2610 ; n2611
g2548 and n790 n2611 ; n2612
g2549 and n2605 n2612 ; n2613
g2550 and n2591 n2613 ; n2614
g2551 and n1602 n2614 ; n2615
g2552 and n2583 n2615 ; n2616
g2553 and n2582 n2616 ; n2617
g2554 and n364_not n2617 ; n2618
g2555 and n168_not n2618 ; n2619
g2556 and n352_not n2619 ; n2620
g2557 and n118_not n2620 ; n2621
g2558 and n424_not n2621 ; n2622
g2559 and n673_not n2622 ; n2623
g2560 and n511_not n616 ; n2624
g2561 and n130_not n2624 ; n2625
g2562 nor n194 n558 ; n2626
g2563 and n714_not n2626 ; n2627
g2564 and n2625 n2627 ; n2628
g2565 and n2371 n2628 ; n2629
g2566 and n242_not n2629 ; n2630
g2567 and n357_not n2630 ; n2631
g2568 and n712_not n2631 ; n2632
g2569 nor n123 n393 ; n2633
g2570 nor n177 n201 ; n2634
g2571 and n252_not n2634 ; n2635
g2572 and n206_not n2635 ; n2636
g2573 and n358_not n2636 ; n2637
g2574 and n1578 n1828 ; n2638
g2575 and n2637 n2638 ; n2639
g2576 and n1738 n2639 ; n2640
g2577 and n1419 n2640 ; n2641
g2578 and n811 n2641 ; n2642
g2579 and n2633 n2642 ; n2643
g2580 and n933 n2643 ; n2644
g2581 and n2484 n2644 ; n2645
g2582 and n397_not n2645 ; n2646
g2583 and n102_not n2646 ; n2647
g2584 and n237_not n2647 ; n2648
g2585 and n562_not n2648 ; n2649
g2586 and n655_not n2649 ; n2650
g2587 nor n91 n505 ; n2651
g2588 and n282 n2651 ; n2652
g2589 and n527_not n2652 ; n2653
g2590 nor n420 n602 ; n2654
g2591 and n173_not n2654 ; n2655
g2592 and n493_not n2655 ; n2656
g2593 and n2653 n2656 ; n2657
g2594 and n2650 n2657 ; n2658
g2595 and n2632 n2658 ; n2659
g2596 and n2623 n2659 ; n2660
g2597 and n2581 n2660 ; n2661
g2598 and n2573 n2661 ; n2662
g2599 and n159 n2662 ; n2663
g2600 and n979 n2663 ; n2664
g2601 and n720 n2664 ; n2665
g2602 and n1072_not n2665 ; n2666
g2603 and n469_not n2666 ; n2667
g2604 and n518_not n2667 ; n2668
g2605 and n980_not n2668 ; n2669
g2606 and n277_not n2669 ; n2670
g2607 and n564_not n2670 ; n2671
g2608 and n371_not n2671 ; n2672
g2609 and n188_not n2672 ; n2673
g2610 and n231_not n2673 ; n2674
g2611 nor n2571 n2674 ; n2675
g2612 nor n355 n504 ; n2676
g2613 and n240_not n2676 ; n2677
g2614 and n304_not n2677 ; n2678
g2615 and n128 n1121 ; n2679
g2616 and n603_not n2679 ; n2680
g2617 and n1203_not n2680 ; n2681
g2618 and n531_not n2681 ; n2682
g2619 nor n222 n287 ; n2683
g2620 and n115_not n2683 ; n2684
g2621 and n2390 n2684 ; n2685
g2622 and n2133 n2685 ; n2686
g2623 and n1387 n2686 ; n2687
g2624 and n2682 n2687 ; n2688
g2625 and n2325 n2688 ; n2689
g2626 and n1182 n2689 ; n2690
g2627 and n979 n2690 ; n2691
g2628 and n2583 n2691 ; n2692
g2629 and n169_not n2692 ; n2693
g2630 and n396_not n2693 ; n2694
g2631 and n1104_not n2694 ; n2695
g2632 and n883_not n2695 ; n2696
g2633 and n95_not n2696 ; n2697
g2634 nor n422 n525 ; n2698
g2635 nor n571 n809 ; n2699
g2636 and n514_not n2699 ; n2700
g2637 and n339_not n2700 ; n2701
g2638 and n233_not n2701 ; n2702
g2639 and n248_not n2702 ; n2703
g2640 nor n601 n875 ; n2704
g2641 nor n175 n295 ; n2705
g2642 and n1636 n2705 ; n2706
g2643 and n2704 n2706 ; n2707
g2644 and n2507 n2707 ; n2708
g2645 and n1011_not n2708 ; n2709
g2646 and n495_not n2709 ; n2710
g2647 and n118_not n2710 ; n2711
g2648 and n400_not n2711 ; n2712
g2649 and n777_not n2712 ; n2713
g2650 and n394_not n2713 ; n2714
g2651 and n886_not n2714 ; n2715
g2652 and n270_not n2715 ; n2716
g2653 and n453_not n1782 ; n2717
g2654 and n306_not n2717 ; n2718
g2655 and n249_not n2718 ; n2719
g2656 nor n255 n563 ; n2720
g2657 and n86_not n2720 ; n2721
g2658 and n2303 n2721 ; n2722
g2659 and n2230 n2722 ; n2723
g2660 and n2719 n2723 ; n2724
g2661 and n2650 n2724 ; n2725
g2662 and n2716 n2725 ; n2726
g2663 and n2703 n2726 ; n2727
g2664 and n2698 n2727 ; n2728
g2665 and n1183 n2728 ; n2729
g2666 and n2697 n2729 ; n2730
g2667 and n2678 n2730 ; n2731
g2668 and n937 n2731 ; n2732
g2669 and n619_not n2732 ; n2733
g2670 and n639_not n2733 ; n2734
g2671 and n200_not n2734 ; n2735
g2672 and n1010_not n2735 ; n2736
g2673 nor n2674 n2736 ; n2737
g2674 nor n229 n1246 ; n2738
g2675 nor n334 n656 ; n2739
g2676 nor n151 n171 ; n2740
g2677 and n355_not n804 ; n2741
g2678 and n875_not n2741 ; n2742
g2679 and n2740 n2742 ; n2743
g2680 and n2739 n2743 ; n2744
g2681 and n1128 n2744 ; n2745
g2682 and n135_not n2745 ; n2746
g2683 and n809_not n2746 ; n2747
g2684 and n223_not n2747 ; n2748
g2685 and n715_not n2748 ; n2749
g2686 and n438_not n2749 ; n2750
g2687 and n252_not n2750 ; n2751
g2688 nor n436 n567 ; n2752
g2689 and n400_not n520 ; n2753
g2690 and n2752 n2753 ; n2754
g2691 and n2445 n2754 ; n2755
g2692 and n2544 n2755 ; n2756
g2693 and n494 n2756 ; n2757
g2694 nor n152 n617 ; n2758
g2695 and n118_not n2758 ; n2759
g2696 and n1314 n2759 ; n2760
g2697 and n2757 n2760 ; n2761
g2698 and n2751 n2761 ; n2762
g2699 and n2738 n2762 ; n2763
g2700 and n1253 n2763 ; n2764
g2701 and n2651 n2764 ; n2765
g2702 and n507 n2765 ; n2766
g2703 and n254_not n2766 ; n2767
g2704 and n328_not n2767 ; n2768
g2705 and n299_not n2768 ; n2769
g2706 and n568_not n2769 ; n2770
g2707 and n243_not n2770 ; n2771
g2708 and n531_not n2771 ; n2772
g2709 nor n746 n1011 ; n2773
g2710 and n402_not n2773 ; n2774
g2711 and n305_not n2774 ; n2775
g2712 and n825_not n2775 ; n2776
g2713 and n672_not n2776 ; n2777
g2714 and n371_not n2777 ; n2778
g2715 and n566 n1727 ; n2779
g2716 and n426_not n2779 ; n2780
g2717 and n367_not n2780 ; n2781
g2718 and n145_not n2781 ; n2782
g2719 and n418 n492_not ; n2783
g2720 and n245_not n2783 ; n2784
g2721 and n632 n2784 ; n2785
g2722 and n204 n2785 ; n2786
g2723 and n2782 n2786 ; n2787
g2724 and n2778 n2787 ; n2788
g2725 and n1994 n2788 ; n2789
g2726 and n515 n2789 ; n2790
g2727 and n1237 n2790 ; n2791
g2728 and n634 n2791 ; n2792
g2729 and n416_not n2792 ; n2793
g2730 and n714_not n2793 ; n2794
g2731 and n393_not n2794 ; n2795
g2732 and n489_not n2795 ; n2796
g2733 and n1025 n1602 ; n2797
g2734 and n1426 n2797 ; n2798
g2735 and n654 n2798 ; n2799
g2736 and n1072_not n2799 ; n2800
g2737 and n509_not n2800 ; n2801
g2738 and n147_not n2801 ; n2802
g2739 and n130_not n2802 ; n2803
g2740 and n525_not n2803 ; n2804
g2741 and n127_not n2804 ; n2805
g2742 and n655_not n2805 ; n2806
g2743 nor n132 n325 ; n2807
g2744 nor n194 n886 ; n2808
g2745 nor n293 n372 ; n2809
g2746 and n164_not n2073 ; n2810
g2747 and n277_not n2810 ; n2811
g2748 and n1828 n2811 ; n2812
g2749 and n2809 n2812 ; n2813
g2750 and n2808 n2813 ; n2814
g2751 and n2807 n2814 ; n2815
g2752 and n1709 n2815 ; n2816
g2753 and n2806 n2816 ; n2817
g2754 and n2796 n2817 ; n2818
g2755 and n2772 n2818 ; n2819
g2756 and n789 n2819 ; n2820
g2757 and n1577 n2820 ; n2821
g2758 and n1917 n2821 ; n2822
g2759 and n533 n2822 ; n2823
g2760 and n421 n2823 ; n2824
g2761 and n2276 n2824 ; n2825
g2762 and n284_not n2825 ; n2826
g2763 and n146_not n2826 ; n2827
g2764 and n331_not n2827 ; n2828
g2765 and n274_not n2828 ; n2829
g2766 and n2674 n2736_not ; n2830
g2767 and n2829_not n2830 ; n2831
g2768 nor n2737 n2831 ; n2832
g2769 and n2571 n2674 ; n2833
g2770 nor n2675 n2833 ; n2834
g2771 and n2832_not n2834 ; n2835
g2772 nor n2675 n2835 ; n2836
g2773 and n2533 n2571 ; n2837
g2774 nor n2572 n2837 ; n2838
g2775 and n2836_not n2838 ; n2839
g2776 nor n2572 n2839 ; n2840
g2777 and n2464 n2533 ; n2841
g2778 nor n2534 n2841 ; n2842
g2779 and n2840_not n2842 ; n2843
g2780 nor n2534 n2843 ; n2844
g2781 and n2388 n2464 ; n2845
g2782 nor n2465 n2845 ; n2846
g2783 and n2844_not n2846 ; n2847
g2784 nor n2465 n2847 ; n2848
g2785 and n2291 n2388 ; n2849
g2786 nor n2389 n2849 ; n2850
g2787 and n2848_not n2850 ; n2851
g2788 nor n2389 n2851 ; n2852
g2789 and n2189 n2291 ; n2853
g2790 nor n2292 n2853 ; n2854
g2791 and n2852_not n2854 ; n2855
g2792 nor n2292 n2855 ; n2856
g2793 and n2152 n2189 ; n2857
g2794 nor n2190 n2857 ; n2858
g2795 and n2856_not n2858 ; n2859
g2796 nor n2190 n2859 ; n2860
g2797 and n2057 n2152 ; n2861
g2798 nor n2153 n2861 ; n2862
g2799 and n2860_not n2862 ; n2863
g2800 nor n2153 n2863 ; n2864
g2801 and n1992 n2057 ; n2865
g2802 nor n2058 n2865 ; n2866
g2803 and n2864_not n2866 ; n2867
g2804 nor n2058 n2867 ; n2868
g2805 and n1913 n1992 ; n2869
g2806 nor n1993 n2869 ; n2870
g2807 and n2868_not n2870 ; n2871
g2808 nor n1993 n2871 ; n2872
g2809 and n1877 n1913 ; n2873
g2810 nor n1914 n2873 ; n2874
g2811 and n2872_not n2874 ; n2875
g2812 nor n1914 n2875 ; n2876
g2813 and n1779 n1877 ; n2877
g2814 nor n1878 n2877 ; n2878
g2815 and n2876_not n2878 ; n2879
g2816 nor n1878 n2879 ; n2880
g2817 and n1665 n1779 ; n2881
g2818 nor n1780 n2881 ; n2882
g2819 and n2880_not n2882 ; n2883
g2820 nor n1780 n2883 ; n2884
g2821 and n1572 n1665 ; n2885
g2822 nor n1666 n2885 ; n2886
g2823 and n2884_not n2886 ; n2887
g2824 nor n1666 n2887 ; n2888
g2825 and n1472 n1572 ; n2889
g2826 nor n1573 n2889 ; n2890
g2827 and n2888_not n2890 ; n2891
g2828 nor n1573 n2891 ; n2892
g2829 and n1364 n1472 ; n2893
g2830 nor n1473 n2893 ; n2894
g2831 and n2892_not n2894 ; n2895
g2832 nor n1473 n2895 ; n2896
g2833 and n1235 n1364 ; n2897
g2834 nor n1365 n2897 ; n2898
g2835 and n2896_not n2898 ; n2899
g2836 nor n1365 n2899 ; n2900
g2837 and n1178 n1235 ; n2901
g2838 nor n1236 n2901 ; n2902
g2839 and n2900_not n2902 ; n2903
g2840 nor n1236 n2903 ; n2904
g2841 and n1060 n1178 ; n2905
g2842 nor n1179 n2905 ; n2906
g2843 and n2904_not n2906 ; n2907
g2844 nor n1179 n2907 ; n2908
g2845 and n958 n1060 ; n2909
g2846 nor n1061 n2909 ; n2910
g2847 and n2908_not n2910 ; n2911
g2848 nor n1061 n2911 ; n2912
g2849 and n867 n958 ; n2913
g2850 nor n959 n2913 ; n2914
g2851 and n2912_not n2914 ; n2915
g2852 nor n959 n2915 ; n2916
g2853 and n710 n867 ; n2917
g2854 nor n868 n2917 ; n2918
g2855 and n2916_not n2918 ; n2919
g2856 nor n868 n2919 ; n2920
g2857 and n587 n710 ; n2921
g2858 nor n711 n2921 ; n2922
g2859 and n2920_not n2922 ; n2923
g2860 nor n711 n2923 ; n2924
g2861 and n392 n587 ; n2925
g2862 nor n588 n2925 ; n2926
g2863 and n2924_not n2926 ; n2927
g2864 nor n588 n2927 ; n2928
g2865 nor n206 n327 ; n2929
g2866 and n468_not n2929 ; n2930
g2867 and n655_not n2930 ; n2931
g2868 and n2090 n2931 ; n2932
g2869 and n1072_not n2932 ; n2933
g2870 and n557_not n2933 ; n2934
g2871 and n426_not n2934 ; n2935
g2872 and n637_not n2935 ; n2936
g2873 and n306_not n2936 ; n2937
g2874 and n672_not n2937 ; n2938
g2875 and n337_not n2938 ; n2939
g2876 and n771_not n2939 ; n2940
g2877 and n149_not n1556 ; n2941
g2878 and n568_not n2941 ; n2942
g2879 and n99_not n2942 ; n2943
g2880 and n990 n1408 ; n2944
g2881 and n2943 n2944 ; n2945
g2882 and n2940 n2945 ; n2946
g2883 and n2219 n2946 ; n2947
g2884 and n1180 n2947 ; n2948
g2885 and n301_not n2948 ; n2949
g2886 and n276_not n2949 ; n2950
g2887 and n355_not n2950 ; n2951
g2888 and n335_not n2951 ; n2952
g2889 and n639_not n2952 ; n2953
g2890 and n714_not n2953 ; n2954
g2891 and n274_not n2954 ; n2955
g2892 and n240_not n2955 ; n2956
g2893 and n277_not n2956 ; n2957
g2894 and n325_not n2957 ; n2958
g2895 and n2263 n2752 ; n2959
g2896 and n462_not n2959 ; n2960
g2897 and n980_not n2960 ; n2961
g2898 and n713_not n1760 ; n2962
g2899 and n281_not n2962 ; n2963
g2900 and n832 n1423 ; n2964
g2901 and n2230 n2964 ; n2965
g2902 and n2963 n2965 ; n2966
g2903 and n2961 n2966 ; n2967
g2904 and n1916 n2967 ; n2968
g2905 and n2021 n2968 ; n2969
g2906 and n288 n2969 ; n2970
g2907 and n533 n2970 ; n2971
g2908 and n1825 n2971 ; n2972
g2909 and n2466 n2972 ; n2973
g2910 and n594_not n2973 ; n2974
g2911 and n470_not n2974 ; n2975
g2912 and n592_not n2975 ; n2976
g2913 and n666_not n2976 ; n2977
g2914 and n489_not n2977 ; n2978
g2915 and n249_not n2978 ; n2979
g2916 and n171_not n2409 ; n2980
g2917 and n305_not n2980 ; n2981
g2918 and n102_not n2981 ; n2982
g2919 and n331_not n2982 ; n2983
g2920 and n283_not n2983 ; n2984
g2921 and n372_not n2984 ; n2985
g2922 and n1010_not n2985 ; n2986
g2923 and n519_not n2986 ; n2987
g2924 and n634 n1009 ; n2988
g2925 and n289_not n2988 ; n2989
g2926 and n531_not n2989 ; n2990
g2927 and n352_not n421 ; n2991
g2928 and n338_not n2991 ; n2992
g2929 nor n121 n177 ; n2993
g2930 and n398_not n2993 ; n2994
g2931 and n115_not n2994 ; n2995
g2932 and n2113 n2995 ; n2996
g2933 and n2992 n2996 ; n2997
g2934 and n2990 n2997 ; n2998
g2935 and n1823 n2998 ; n2999
g2936 and n2987 n2999 ; n3000
g2937 and n2979 n3000 ; n3001
g2938 and n244 n3001 ; n3002
g2939 and n2958 n3002 ; n3003
g2940 and n590 n3003 ; n3004
g2941 and n1389 n3004 ; n3005
g2942 and n136_not n3005 ; n3006
g2943 and n506_not n3006 ; n3007
g2944 and n357_not n3007 ; n3008
g2945 and n326_not n3008 ; n3009
g2946 and n1203_not n3009 ; n3010
g2947 and n200_not n3010 ; n3011
g2948 and n371_not n3011 ; n3012
g2949 nor n392 n3012 ; n3013
g2950 and n392 n3012 ; n3014
g2951 nor n3013 n3014 ; n3015
g2952 and n2928_not n3015 ; n3016
g2953 and n2928 n3015_not ; n3017
g2954 nor n3016 n3017 ; n3018
g2955 and n75 n3018 ; n3019
g2956 nor a[31] n74 ; n3020
g2957 and n3012_not n3020 ; n3021
g2958 and a[30] n74 ; n3022
g2959 and a[31] n3022 ; n3023
g2960 and n587_not n3023 ; n3024
g2961 and a[30] a[31]_not ; n3025
g2962 and a[30]_not a[31] ; n3026
g2963 nor n3025 n3026 ; n3027
g2964 and n74 n3027_not ; n3028
g2965 and n392_not n3028 ; n3029
g2966 nor n3024 n3029 ; n3030
g2967 and n3021_not n3030 ; n3031
g2968 and n3019_not n3031 ; n3032
g2969 and n275_not n2760 ; n3033
g2970 and n292_not n3033 ; n3034
g2971 and n357_not n3034 ; n3035
g2972 and n274_not n3035 ; n3036
g2973 and n245_not n3036 ; n3037
g2974 and n623_not n3037 ; n3038
g2975 and n489_not n3038 ; n3039
g2976 nor n286 n453 ; n3040
g2977 nor n325 n1127 ; n3041
g2978 nor n188 n656 ; n3042
g2979 nor n190 n527 ; n3043
g2980 nor n400 n713 ; n3044
g2981 and n191_not n3044 ; n3045
g2982 and n3043 n3045 ; n3046
g2983 and n3042 n3046 ; n3047
g2984 and n3041 n3047 ; n3048
g2985 and n3040 n3048 ; n3049
g2986 and n1781 n3049 ; n3050
g2987 and n285 n3050 ; n3051
g2988 and n3039 n3051 ; n3052
g2989 and n533 n3052 ; n3053
g2990 and n1141 n3053 ; n3054
g2991 and n509_not n3054 ; n3055
g2992 and n667_not n3055 ; n3056
g2993 and n563_not n3056 ; n3057
g2994 nor n641 n752 ; n3058
g2995 and n637_not n3058 ; n3059
g2996 and n276_not n3059 ; n3060
g2997 and n397_not n3060 ; n3061
g2998 and n490_not n3061 ; n3062
g2999 and n200_not n3062 ; n3063
g3000 and n161_not n3063 ; n3064
g3001 and n1010_not n3064 ; n3065
g3002 and n1246_not n2633 ; n3066
g3003 and n135_not n3066 ; n3067
g3004 and n562_not n3067 ; n3068
g3005 and n373 n573 ; n3069
g3006 and n1438 n3069 ; n3070
g3007 and n3068 n3070 ; n3071
g3008 and n494 n3071 ; n3072
g3009 and n931 n3072 ; n3073
g3010 and n2317 n3073 ; n3074
g3011 and n2651 n3074 ; n3075
g3012 and n3065 n3075 ; n3076
g3013 and n3057 n3076 ; n3077
g3014 and n804 n3077 ; n3078
g3015 and n427_not n3078 ; n3079
g3016 and n353_not n3079 ; n3080
g3017 and n1102_not n3080 ; n3081
g3018 and n203_not n3081 ; n3082
g3019 and n240_not n3082 ; n3083
g3020 nor n203 n791 ; n3084
g3021 and n532_not n3084 ; n3085
g3022 and n723 n3085 ; n3086
g3023 and n615 n3086 ; n3087
g3024 and n1246_not n3087 ; n3088
g3025 and n135_not n3088 ; n3089
g3026 and n328_not n3089 ; n3090
g3027 and n290_not n3090 ; n3091
g3028 and n961_not n3091 ; n3092
g3029 and n142_not n3092 ; n3093
g3030 and n358_not n3093 ; n3094
g3031 and n497 n3059 ; n3095
g3032 and n3094 n3095 ; n3096
g3033 and n2698 n3096 ; n3097
g3034 and n2573 n3097 ; n3098
g3035 and n1827 n3098 ; n3099
g3036 and n1884 n3099 ; n3100
g3037 and n136_not n3100 ; n3101
g3038 and n177_not n3101 ; n3102
g3039 and n118_not n3102 ; n3103
g3040 and n228_not n3103 ; n3104
g3041 and n287_not n3104 ; n3105
g3042 and n505_not n3105 ; n3106
g3043 and n170_not n3106 ; n3107
g3044 and n666_not n3107 ; n3108
g3045 and n462_not n2191 ; n3109
g3046 and n713_not n3109 ; n3110
g3047 and n281_not n3110 ; n3111
g3048 and n173_not n3111 ; n3112
g3049 and n1203_not n3112 ; n3113
g3050 and n275_not n2347 ; n3114
g3051 and n168_not n968 ; n3115
g3052 and n1333 n3115 ; n3116
g3053 and n3114 n3116 ; n3117
g3054 and n1132 n3117 ; n3118
g3055 and n3113 n3118 ; n3119
g3056 and n1917 n3119 ; n3120
g3057 and n2678 n3120 ; n3121
g3058 and n1781 n3121 ; n3122
g3059 and n1366 n3122 ; n3123
g3060 and n1248 n3123 ; n3124
g3061 and n242_not n3124 ; n3125
g3062 and n191_not n3125 ; n3126
g3063 and n127_not n3126 ; n3127
g3064 and n618 n847_not ; n3128
g3065 and n897 n3128 ; n3129
g3066 and n439 n3129 ; n3130
g3067 and n690 n3130 ; n3131
g3068 and n2091 n3131 ; n3132
g3069 and n1126 n3132 ; n3133
g3070 and n1488 n3133 ; n3134
g3071 and n3127 n3134 ; n3135
g3072 and n512 n3135 ; n3136
g3073 and n3108 n3136 ; n3137
g3074 and n1994 n3137 ; n3138
g3075 and n1237 n3138 ; n3139
g3076 and n341 n3139 ; n3140
g3077 and n1306_not n3140 ; n3141
g3078 and n461_not n3141 ; n3142
g3079 and n403_not n3142 ; n3143
g3080 and n492_not n3143 ; n3144
g3081 and n163_not n3144 ; n3145
g3082 and n271_not n3145 ; n3146
g3083 nor n334 n462 ; n3147
g3084 and n531_not n3147 ; n3148
g3085 and n128 n3148 ; n3149
g3086 and n2467 n3149 ; n3150
g3087 and n505_not n3150 ; n3151
g3088 and n466_not n3151 ; n3152
g3089 and n519_not n3152 ; n3153
g3090 and n251_not n3153 ; n3154
g3091 and n363_not n3154 ; n3155
g3092 and n876 n2808 ; n3156
g3093 and n402_not n3156 ; n3157
g3094 and n460_not n3157 ; n3158
g3095 and n298_not n3158 ; n3159
g3096 nor n325 n803 ; n3160
g3097 and n712_not n747 ; n3161
g3098 and n1010_not n3161 ; n3162
g3099 nor n168 n425 ; n3163
g3100 and n474_not n3163 ; n3164
g3101 and n222_not n3164 ; n3165
g3102 and n2349 n3165 ; n3166
g3103 and n3162 n3166 ; n3167
g3104 and n3160 n3167 ; n3168
g3105 and n665 n3168 ; n3169
g3106 and n2633 n3169 ; n3170
g3107 and n1063 n3170 ; n3171
g3108 and n1139 n3171 ; n3172
g3109 and n804 n3172 ; n3173
g3110 and n3159 n3173 ; n3174
g3111 and n810 n3174 ; n3175
g3112 and n341 n3175 ; n3176
g3113 and n136_not n3176 ; n3177
g3114 and n255_not n3177 ; n3178
g3115 and n656_not n3178 ; n3179
g3116 and n417_not n3179 ; n3180
g3117 and n401 n510 ; n3181
g3118 and n193 n3181 ; n3182
g3119 and n111_not n3182 ; n3183
g3120 and n203_not n3183 ; n3184
g3121 and n368_not n3184 ; n3185
g3122 and n163_not n3185 ; n3186
g3123 and n273_not n3186 ; n3187
g3124 and n237_not n3187 ; n3188
g3125 and n225_not n3188 ; n3189
g3126 and n295_not n3189 ; n3190
g3127 and n270_not n3190 ; n3191
g3128 and n507 n1011_not ; n3192
g3129 nor n276 n330 ; n3193
g3130 and n152_not n3193 ; n3194
g3131 and n3192 n3194 ; n3195
g3132 and n1423 n3195 ; n3196
g3133 and n1555 n3196 ; n3197
g3134 and n3191 n3197 ; n3198
g3135 and n1825 n3198 ; n3199
g3136 and n731 n3199 ; n3200
g3137 and n1252 n3200 ; n3201
g3138 and n514_not n3201 ; n3202
g3139 and n327_not n3202 ; n3203
g3140 and n142_not n3203 ; n3204
g3141 and n99_not n3204 ; n3205
g3142 nor n224 n329 ; n3206
g3143 and n617_not n3206 ; n3207
g3144 and n236_not n3207 ; n3208
g3145 and n420_not n3208 ; n3209
g3146 and n752_not n3209 ; n3210
g3147 and n1101_not n3210 ; n3211
g3148 and n248_not n3211 ; n3212
g3149 and n102_not n3212 ; n3213
g3150 and n825_not n3213 ; n3214
g3151 and n167_not n3214 ; n3215
g3152 and n791_not n3215 ; n3216
g3153 and n338_not n3216 ; n3217
g3154 and n592_not n3217 ; n3218
g3155 and n188_not n3218 ; n3219
g3156 and n674 n1531 ; n3220
g3157 and n130_not n3220 ; n3221
g3158 and n468_not n3221 ; n3222
g3159 and n1127_not n3222 ; n3223
g3160 and n95_not n3223 ; n3224
g3161 and n429_not n3224 ; n3225
g3162 nor n233 n395 ; n3226
g3163 and n2332 n3226 ; n3227
g3164 and n3225 n3227 ; n3228
g3165 and n3219 n3228 ; n3229
g3166 and n3205 n3229 ; n3230
g3167 and n3180 n3230 ; n3231
g3168 and n3155 n3231 ; n3232
g3169 and n120 n3232 ; n3233
g3170 and n621 n3233 ; n3234
g3171 and n1574 n3234 ; n3235
g3172 and n713_not n3235 ; n3236
g3173 and n358_not n3236 ; n3237
g3174 and n158_not n3237 ; n3238
g3175 and n249_not n3238 ; n3239
g3176 nor n3146 n3239 ; n3240
g3177 and n3146 n3239 ; n3241
g3178 nor n3240 n3241 ; n3242
g3179 and a[20]_not n3242 ; n3243
g3180 nor n3240 n3243 ; n3244
g3181 and n3083 n3244_not ; n3245
g3182 and n3083_not n3244 ; n3246
g3183 nor n3245 n3246 ; n3247
g3184 and n3032_not n3247 ; n3248
g3185 nor n3032 n3248 ; n3249
g3186 and n3247 n3248_not ; n3250
g3187 nor n3249 n3250 ; n3251
g3188 nor n173 n226 ; n3252
g3189 and n398_not n2705 ; n3253
g3190 and n154_not n3253 ; n3254
g3191 and n281_not n3254 ; n3255
g3192 and n656_not n3255 ; n3256
g3193 and n637_not n3256 ; n3257
g3194 and n192_not n3257 ; n3258
g3195 and n791_not n3258 ; n3259
g3196 and n255_not n1394 ; n3260
g3197 and n273_not n3260 ; n3261
g3198 and n354_not n539 ; n3262
g3199 and n224_not n3262 ; n3263
g3200 and n666_not n3263 ; n3264
g3201 and n271_not n471 ; n3265
g3202 and n363_not n3265 ; n3266
g3203 and n1063 n1128 ; n3267
g3204 and n225_not n3267 ; n3268
g3205 and n3266 n3268 ; n3269
g3206 and n3264 n3269 ; n3270
g3207 and n2931 n3270 ; n3271
g3208 and n1012 n3271 ; n3272
g3209 and n3261 n3272 ; n3273
g3210 and n3259 n3273 ; n3274
g3211 and n773 n3274 ; n3275
g3212 and n291 n3275 ; n3276
g3213 and n353_not n3276 ; n3277
g3214 and n641_not n3277 ; n3278
g3215 and n352_not n3278 ; n3279
g3216 and n563_not n3279 ; n3280
g3217 and n633_not n3280 ; n3281
g3218 and n188_not n3281 ; n3282
g3219 nor n557 n1246 ; n3283
g3220 and n803_not n3283 ; n3284
g3221 and n334_not n3284 ; n3285
g3222 and n299_not n3285 ; n3286
g3223 and n527_not n3286 ; n3287
g3224 and n639_not n3287 ; n3288
g3225 and n525_not n3288 ; n3289
g3226 and n270_not n3289 ; n3290
g3227 and n280_not n720 ; n3291
g3228 and n715_not n3291 ; n3292
g3229 and n961_not n3292 ; n3293
g3230 and n142_not n3293 ; n3294
g3231 and n932_not n3294 ; n3295
g3232 and n531_not n3295 ; n3296
g3233 and n205_not n2651 ; n3297
g3234 and n222_not n3297 ; n3298
g3235 nor n395 n452 ; n3299
g3236 and n489_not n3299 ; n3300
g3237 and n3298 n3300 ; n3301
g3238 and n3296 n3301 ; n3302
g3239 and n1523 n3302 ; n3303
g3240 and n3290 n3303 ; n3304
g3241 and n1479 n3304 ; n3305
g3242 and n128 n3305 ; n3306
g3243 and n423 n3306 ; n3307
g3244 and n731 n3307 ; n3308
g3245 and n507 n3308 ; n3309
g3246 and n393_not n3309 ; n3310
g3247 and n451_not n3310 ; n3311
g3248 and n231_not n3311 ; n3312
g3249 nor n397 n435 ; n3313
g3250 and n438_not n3313 ; n3314
g3251 and n1071 n3314 ; n3315
g3252 and n1931 n3315 ; n3316
g3253 and n524 n3316 ; n3317
g3254 and n2237 n3317 ; n3318
g3255 and n3312 n3318 ; n3319
g3256 and n3282 n3319 ; n3320
g3257 and n872 n3320 ; n3321
g3258 and n3252 n3321 ; n3322
g3259 and n804 n3322 ; n3323
g3260 and n570 n3323 ; n3324
g3261 and n233_not n3324 ; n3325
g3262 and n594_not n3325 ; n3326
g3263 and n158_not n3326 ; n3327
g3264 and n3146 n3327_not ; n3328
g3265 and n3146_not n3327 ; n3329
g3266 and n2920 n2922_not ; n3330
g3267 nor n2923 n3330 ; n3331
g3268 and n75 n3331 ; n3332
g3269 and n587_not n3020 ; n3333
g3270 and n867_not n3023 ; n3334
g3271 and n710_not n3028 ; n3335
g3272 nor n3334 n3335 ; n3336
g3273 and n3333_not n3336 ; n3337
g3274 and n3332_not n3337 ; n3338
g3275 nor n3328 n3338 ; n3339
g3276 and n3329_not n3339 ; n3340
g3277 nor n3328 n3340 ; n3341
g3278 nor a[20] n3243 ; n3342
g3279 and n3241_not n3244 ; n3343
g3280 nor n3342 n3343 ; n3344
g3281 nor n3341 n3344 ; n3345
g3282 and n2924 n2926_not ; n3346
g3283 nor n2927 n3346 ; n3347
g3284 and n75 n3347 ; n3348
g3285 and n392_not n3020 ; n3349
g3286 and n710_not n3023 ; n3350
g3287 and n587_not n3028 ; n3351
g3288 nor n3350 n3351 ; n3352
g3289 and n3349_not n3352 ; n3353
g3290 and n3348_not n3353 ; n3354
g3291 and n3341 n3344 ; n3355
g3292 nor n3345 n3355 ; n3356
g3293 and n3354_not n3356 ; n3357
g3294 nor n3345 n3357 ; n3358
g3295 nor n3251 n3358 ; n3359
g3296 and n3251 n3358 ; n3360
g3297 nor n3359 n3360 ; n3361
g3298 and a[28] a[29]_not ; n3362
g3299 and a[28]_not a[29] ; n3363
g3300 nor n3362 n3363 ; n3364
g3301 and a[26] a[27]_not ; n3365
g3302 and a[26]_not a[27] ; n3366
g3303 nor n3365 n3366 ; n3367
g3304 nor n3364 n3367 ; n3368
g3305 nor n469 n656 ; n3369
g3306 and n1010_not n3369 ; n3370
g3307 and n2426 n3370 ; n3371
g3308 and n2361 n3371 ; n3372
g3309 and n194_not n3372 ; n3373
g3310 and n746_not n3373 ; n3374
g3311 and n339_not n3374 ; n3375
g3312 and n145_not n3375 ; n3376
g3313 and n567_not n3376 ; n3377
g3314 and n393_not n3377 ; n3378
g3315 nor n146 n536 ; n3379
g3316 and n428_not n3379 ; n3380
g3317 and n301_not n3380 ; n3381
g3318 and n511_not n3381 ; n3382
g3319 and n461_not n3382 ; n3383
g3320 and n563_not n3383 ; n3384
g3321 and n689_not n3384 ; n3385
g3322 and n200_not n3385 ; n3386
g3323 and n1306_not n2508 ; n3387
g3324 and n154_not n3387 ; n3388
g3325 and n417_not n3388 ; n3389
g3326 nor n372 n427 ; n3390
g3327 and n332_not n3390 ; n3391
g3328 and n937 n1181 ; n3392
g3329 and n641_not n3392 ; n3393
g3330 and n1392 n1739 ; n3394
g3331 and n3393 n3394 ; n3395
g3332 and n3391 n3395 ; n3396
g3333 and n3389 n3396 ; n3397
g3334 and n3386 n3397 ; n3398
g3335 and n291 n3398 ; n3399
g3336 and n617_not n3399 ; n3400
g3337 and n135_not n3400 ; n3401
g3338 and n460_not n3401 ; n3402
g3339 and n451_not n3402 ; n3403
g3340 and n337_not n3403 ; n3404
g3341 and n875_not n3404 ; n3405
g3342 and n667_not n2073 ; n3406
g3343 and n752_not n3406 ; n3407
g3344 and n118_not n3407 ; n3408
g3345 nor n254 n335 ; n3409
g3346 and n300 n962 ; n3410
g3347 and n3409 n3410 ; n3411
g3348 and n1072_not n3411 ; n3412
g3349 and n513_not n3412 ; n3413
g3350 and n191_not n3413 ; n3414
g3351 and n712_not n3414 ; n3415
g3352 and n116 n515 ; n3416
g3353 and n1045 n3416 ; n3417
g3354 and n3266 n3417 ; n3418
g3355 and n1388 n3418 ; n3419
g3356 and n1132 n3419 ; n3420
g3357 and n3415 n3420 ; n3421
g3358 and n3408 n3421 ; n3422
g3359 and n1528 n3422 ; n3423
g3360 and n873 n3423 ; n3424
g3361 and n1182 n3424 ; n3425
g3362 and n720 n3425 ; n3426
g3363 and n121_not n3426 ; n3427
g3364 and n305_not n3427 ; n3428
g3365 and n226_not n3428 ; n3429
g3366 and n403_not n3429 ; n3430
g3367 and n206_not n3430 ; n3431
g3368 and n492_not n3431 ; n3432
g3369 and n352_not n1141 ; n3433
g3370 and n537_not n3433 ; n3434
g3371 and n603_not n3434 ; n3435
g3372 nor n568 n716 ; n3436
g3373 and n142_not n3436 ; n3437
g3374 nor n86 n240 ; n3438
g3375 and n3437 n3438 ; n3439
g3376 and n3435 n3439 ; n3440
g3377 and n3225 n3440 ; n3441
g3378 and n3432 n3441 ; n3442
g3379 and n3405 n3442 ; n3443
g3380 and n2740 n3443 ; n3444
g3381 and n3378 n3444 ; n3445
g3382 and n247 n3445 ; n3446
g3383 and n1917 n3446 ; n3447
g3384 and n491 n3447 ; n3448
g3385 and n978 n3448 ; n3449
g3386 and n810 n3449 ; n3450
g3387 and n462_not n3450 ; n3451
g3388 and n777_not n3451 ; n3452
g3389 and n225_not n3452 ; n3453
g3390 and n304_not n3453 ; n3454
g3391 and n295_not n3454 ; n3455
g3392 and n519_not n3455 ; n3456
g3393 and n3364 n3367_not ; n3457
g3394 and n3456_not n3457 ; n3458
g3395 nor n119 n271 ; n3459
g3396 and n254_not n3459 ; n3460
g3397 and n496_not n3460 ; n3461
g3398 and n536_not n3461 ; n3462
g3399 and n712_not n3462 ; n3463
g3400 and n1010_not n3463 ; n3464
g3401 and n792 n2091 ; n3465
g3402 and n1101_not n3465 ; n3466
g3403 and n296_not n3466 ; n3467
g3404 and n980_not n3467 ; n3468
g3405 and n623_not n3468 ; n3469
g3406 and n525_not n3469 ; n3470
g3407 and n331_not n2105 ; n3471
g3408 and n453_not n3471 ; n3472
g3409 and n418 n469_not ; n3473
g3410 and n474_not n3473 ; n3474
g3411 and n754 n3226 ; n3475
g3412 and n3474 n3475 ; n3476
g3413 and n2556 n3476 ; n3477
g3414 and n593 n3477 ; n3478
g3415 and n437 n3478 ; n3479
g3416 and n1601 n3479 ; n3480
g3417 and n3472 n3480 ; n3481
g3418 and n615 n3481 ; n3482
g3419 and n1046 n3482 ; n3483
g3420 and n3470 n3483 ; n3484
g3421 and n1576 n3484 ; n3485
g3422 and n570 n3485 ; n3486
g3423 and n330_not n3486 ; n3487
g3424 and n302_not n3487 ; n3488
g3425 and n164_not n3488 ; n3489
g3426 nor n157 n571 ; n3490
g3427 and n401 n2113 ; n3491
g3428 and n1531 n3491 ; n3492
g3429 and n355_not n3492 ; n3493
g3430 and n284_not n3493 ; n3494
g3431 and n777_not n3494 ; n3495
g3432 and n206_not n3495 ; n3496
g3433 and n237_not n3496 ; n3497
g3434 and n941 n1255 ; n3498
g3435 and n2220 n3498 ; n3499
g3436 and n2007 n3499 ; n3500
g3437 and n3497 n3500 ; n3501
g3438 and n614 n3501 ; n3502
g3439 and n2021 n3502 ; n3503
g3440 and n291 n3503 ; n3504
g3441 and n1269 n3504 ; n3505
g3442 and n617_not n3505 ; n3506
g3443 and n224_not n3506 ; n3507
g3444 and n419_not n3507 ; n3508
g3445 and n3490 n3508 ; n3509
g3446 and n366_not n3509 ; n3510
g3447 nor n248 n426 ; n3511
g3448 and n715_not n3511 ; n3512
g3449 and n968 n1062_not ; n3513
g3450 and n425_not n3513 ; n3514
g3451 and n172 n3514 ; n3515
g3452 and n3512 n3515 ; n3516
g3453 and n2022 n3516 ; n3517
g3454 and n3510 n3517 ; n3518
g3455 and n847_not n3518 ; n3519
g3456 and n961_not n3519 ; n3520
g3457 and n245_not n3520 ; n3521
g3458 nor n121 n145 ; n3522
g3459 and n338_not n3522 ; n3523
g3460 nor n286 n332 ; n3524
g3461 and n3298 n3524 ; n3525
g3462 and n3523 n3525 ; n3526
g3463 and n530 n3526 ; n3527
g3464 and n1586 n3527 ; n3528
g3465 and n465 n3528 ; n3529
g3466 and n3521 n3529 ; n3530
g3467 and n3489 n3530 ; n3531
g3468 and n3464 n3531 ; n3532
g3469 and n1029 n3532 ; n3533
g3470 and n1528 n3533 ; n3534
g3471 and n1254 n3534 ; n3535
g3472 and n591 n3535 ; n3536
g3473 and n334_not n3536 ; n3537
g3474 and n192_not n3537 ; n3538
g3475 and n371_not n3538 ; n3539
g3476 nor n79 n82 ; n3540
g3477 and n3364_not n3367 ; n3541
g3478 and n3540_not n3541 ; n3542
g3479 and n3539_not n3542 ; n3543
g3480 nor n233 n884 ; n3544
g3481 nor n713 n791 ; n3545
g3482 and n375_not n3545 ; n3546
g3483 and n332_not n3546 ; n3547
g3484 and n569_not n3547 ; n3548
g3485 nor n226 n1127 ; n3549
g3486 and n1960 n3549 ; n3550
g3487 and n3548 n3550 ; n3551
g3488 and n2010 n3551 ; n3552
g3489 and n1479 n3552 ; n3553
g3490 and n3544 n3553 ; n3554
g3491 and n1574 n3554 ; n3555
g3492 and n421 n3555 ; n3556
g3493 and n354_not n3556 ; n3557
g3494 and n334_not n3557 ; n3558
g3495 and n623_not n3558 ; n3559
g3496 and n116 n1306_not ; n3560
g3497 and n506_not n3560 ; n3561
g3498 and n326_not n3561 ; n3562
g3499 and n568_not n3562 ; n3563
g3500 and n430_not n3563 ; n3564
g3501 and n422_not n3564 ; n3565
g3502 nor n495 n619 ; n3566
g3503 and n357_not n3566 ; n3567
g3504 and n777_not n3567 ; n3568
g3505 and n490_not n3568 ; n3569
g3506 and n428_not n2582 ; n3570
g3507 and n2267 n3570 ; n3571
g3508 and n2013 n3571 ; n3572
g3509 and n2348 n3572 ; n3573
g3510 and n3569 n3573 ; n3574
g3511 and n462_not n3574 ; n3575
g3512 and n563_not n3575 ; n3576
g3513 and n536_not n3576 ; n3577
g3514 and n132_not n3577 ; n3578
g3515 and n338_not n3578 ; n3579
g3516 and n337_not n3579 ; n3580
g3517 nor n355 n426 ; n3581
g3518 and n396_not n3581 ; n3582
g3519 and n470_not n3582 ; n3583
g3520 and n1330 n1826 ; n3584
g3521 and n398_not n3584 ; n3585
g3522 and n95_not n3585 ; n3586
g3523 and n358_not n3586 ; n3587
g3524 and n3583 n3587 ; n3588
g3525 and n3580 n3588 ; n3589
g3526 and n1928 n3589 ; n3590
g3527 and n3565 n3590 ; n3591
g3528 and n221 n3591 ; n3592
g3529 and n1687 n3592 ; n3593
g3530 and n3559 n3593 ; n3594
g3531 and n236_not n3594 ; n3595
g3532 and n135_not n3595 ; n3596
g3533 and n280_not n3596 ; n3597
g3534 and n1101_not n3597 ; n3598
g3535 and n514_not n3598 ; n3599
g3536 and n305_not n3599 ; n3600
g3537 and n689_not n3600 ; n3601
g3538 and n304_not n3601 ; n3602
g3539 and n86_not n3602 ; n3603
g3540 and n489_not n3603 ; n3604
g3541 and n771_not n3604 ; n3605
g3542 and n3367 n3540 ; n3606
g3543 and n3605_not n3606 ; n3607
g3544 nor n3543 n3607 ; n3608
g3545 and n3458_not n3608 ; n3609
g3546 and n3368_not n3609 ; n3610
g3547 nor n3539 n3605 ; n3611
g3548 nor n3012 n3539 ; n3612
g3549 nor n3013 n3016 ; n3613
g3550 and n3012 n3539 ; n3614
g3551 nor n3612 n3614 ; n3615
g3552 and n3613_not n3615 ; n3616
g3553 nor n3612 n3616 ; n3617
g3554 and n3539 n3605 ; n3618
g3555 nor n3611 n3618 ; n3619
g3556 and n3617_not n3619 ; n3620
g3557 nor n3611 n3620 ; n3621
g3558 nor n3456 n3605 ; n3622
g3559 and n3456 n3605 ; n3623
g3560 nor n3622 n3623 ; n3624
g3561 and n3621_not n3624 ; n3625
g3562 and n3621 n3624_not ; n3626
g3563 nor n3625 n3626 ; n3627
g3564 and n3609 n3627_not ; n3628
g3565 nor n3610 n3628 ; n3629
g3566 and a[29] n3629_not ; n3630
g3567 and a[29]_not n3629 ; n3631
g3568 nor n3630 n3631 ; n3632
g3569 and n3361 n3632_not ; n3633
g3570 nor n3359 n3633 ; n3634
g3571 nor n3245 n3248 ; n3635
g3572 and n619_not n1531 ; n3636
g3573 and n509_not n3226 ; n3637
g3574 and n511_not n3637 ; n3638
g3575 and n1062_not n3638 ; n3639
g3576 and n656_not n3639 ; n3640
g3577 and n149_not n3640 ; n3641
g3578 and n367_not n3641 ; n3642
g3579 and n245_not n3642 ; n3643
g3580 and n81_not n3643 ; n3644
g3581 nor n132 n163 ; n3645
g3582 and n202 n3645 ; n3646
g3583 and n557_not n3646 ; n3647
g3584 and n353_not n3647 ; n3648
g3585 and n175_not n3648 ; n3649
g3586 and n243_not n3649 ; n3650
g3587 and n569_not n3650 ; n3651
g3588 and n1408 n1458 ; n3652
g3589 and n3472 n3652 ; n3653
g3590 and n3252 n3653 ; n3654
g3591 and n398_not n3654 ; n3655
g3592 and n232_not n3655 ; n3656
g3593 and n171_not n3656 ; n3657
g3594 and n299_not n3657 ; n3658
g3595 and n357_not n3658 ; n3659
g3596 and n374_not n3659 ; n3660
g3597 and n368_not n3660 ; n3661
g3598 and n95_not n3661 ; n3662
g3599 and n633_not n3662 ; n3663
g3600 and n3651 n3663 ; n3664
g3601 and n2581 n3664 ; n3665
g3602 and n3644 n3665 ; n3666
g3603 and n241 n3666 ; n3667
g3604 and n136_not n3667 ; n3668
g3605 and n3636 n3668 ; n3669
g3606 and n425_not n3669 ; n3670
g3607 and n274_not n3670 ; n3671
g3608 and n466_not n3671 ; n3672
g3609 and n422_not n3672 ; n3673
g3610 and n338_not n3673 ; n3674
g3611 and n655_not n3674 ; n3675
g3612 nor n229 n1072 ; n3676
g3613 and n275_not n3676 ; n3677
g3614 and n461_not n3677 ; n3678
g3615 and n416_not n3678 ; n3679
g3616 and n1203_not n3679 ; n3680
g3617 and n252_not n3680 ; n3681
g3618 nor n504 n641 ; n3682
g3619 and n306_not n3682 ; n3683
g3620 and n272_not n3683 ; n3684
g3621 and n222_not n3684 ; n3685
g3622 and n493_not n1380 ; n3686
g3623 and n1010_not n3686 ; n3687
g3624 and n2427 n3687 ; n3688
g3625 and n723 n3688 ; n3689
g3626 and n3685 n3689 ; n3690
g3627 and n1323 n3690 ; n3691
g3628 and n3681 n3691 ; n3692
g3629 and n3675 n3692 ; n3693
g3630 and n1915 n3693 ; n3694
g3631 and n1046 n3694 ; n3695
g3632 and n1366 n3695 ; n3696
g3633 and n169_not n3696 ; n3697
g3634 and n847_not n3697 ; n3698
g3635 and n151_not n3698 ; n3699
g3636 and n118_not n3699 ; n3700
g3637 and n206_not n3700 ; n3701
g3638 and n452_not n3701 ; n3702
g3639 and n3083 n3702_not ; n3703
g3640 and n3083_not n3702 ; n3704
g3641 nor n3635 n3704 ; n3705
g3642 and n3703_not n3705 ; n3706
g3643 nor n3635 n3706 ; n3707
g3644 nor n3704 n3706 ; n3708
g3645 and n3703_not n3708 ; n3709
g3646 nor n3707 n3709 ; n3710
g3647 and n3020 n3539_not ; n3711
g3648 and n3012_not n3028 ; n3712
g3649 and n392_not n3023 ; n3713
g3650 and n3613 n3615_not ; n3714
g3651 nor n3616 n3714 ; n3715
g3652 and n75 n3715 ; n3716
g3653 nor n3713 n3716 ; n3717
g3654 and n3712_not n3717 ; n3718
g3655 and n3711_not n3718 ; n3719
g3656 nor n3710 n3719 ; n3720
g3657 nor n3710 n3720 ; n3721
g3658 nor n3719 n3720 ; n3722
g3659 nor n3721 n3722 ; n3723
g3660 nor n3634 n3723 ; n3724
g3661 nor n3634 n3724 ; n3725
g3662 nor n3723 n3724 ; n3726
g3663 nor n3725 n3726 ; n3727
g3664 nor n189 n280 ; n3728
g3665 and n115_not n3728 ; n3729
g3666 and n169_not n3729 ; n3730
g3667 and n149_not n3730 ; n3731
g3668 and n490_not n3731 ; n3732
g3669 and n567_not n3732 ; n3733
g3670 and n558_not n1839 ; n3734
g3671 and n667_not n3734 ; n3735
g3672 and n752_not n3735 ; n3736
g3673 and n557_not n3736 ; n3737
g3674 and n223_not n3737 ; n3738
g3675 and n623_not n3738 ; n3739
g3676 and n640 n895 ; n3740
g3677 and n123_not n3740 ; n3741
g3678 and n150_not n3741 ; n3742
g3679 and n231_not n3742 ; n3743
g3680 and n401 n2556 ; n3744
g3681 and n3743 n3744 ; n3745
g3682 and n3739 n3745 ; n3746
g3683 and n3733 n3746 ; n3747
g3684 and n2582 n3747 ; n3748
g3685 and n720 n3748 ; n3749
g3686 and n1141 n3749 ; n3750
g3687 and n515 n3750 ; n3751
g3688 and n1367 n3751 ; n3752
g3689 and n803_not n3752 ; n3753
g3690 and n511_not n3753 ; n3754
g3691 and n177_not n3754 ; n3755
g3692 and n147_not n3755 ; n3756
g3693 and n425_not n3756 ; n3757
g3694 and n620_not n2293 ; n3758
g3695 and n205_not n3758 ; n3759
g3696 and n161_not n3759 ; n3760
g3697 and n474_not n3760 ; n3761
g3698 and n340_not n3761 ; n3762
g3699 and n436_not n3762 ; n3763
g3700 and n564_not n3763 ; n3764
g3701 and n1392 n3115 ; n3765
g3702 and n590 n3765 ; n3766
g3703 and n118_not n3766 ; n3767
g3704 and n527_not n3767 ; n3768
g3705 and n422_not n747 ; n3769
g3706 and n1010_not n3769 ; n3770
g3707 and n569_not n3770 ; n3771
g3708 and n1784 n3771 ; n3772
g3709 and n3768 n3772 ; n3773
g3710 and n2512 n3773 ; n3774
g3711 and n872 n3774 ; n3775
g3712 and n276_not n3775 ; n3776
g3713 and n602_not n3776 ; n3777
g3714 and n884_not n3777 ; n3778
g3715 and n394_not n3778 ; n3779
g3716 and n325_not n3779 ; n3780
g3717 and n271_not n3780 ; n3781
g3718 and n428_not n3781 ; n3782
g3719 and n1388 n1577 ; n3783
g3720 and n563_not n3783 ; n3784
g3721 and n132_not n3784 ; n3785
g3722 and n225_not n3785 ; n3786
g3723 and n531_not n3786 ; n3787
g3724 and n657_not n3787 ; n3788
g3725 and n1104_not n3788 ; n3789
g3726 and n86_not n3789 ; n3790
g3727 nor n144 n466 ; n3791
g3728 and n191_not n3791 ; n3792
g3729 and n3040 n3792 ; n3793
g3730 and n3790 n3793 ; n3794
g3731 and n3782 n3794 ; n3795
g3732 and n3764 n3795 ; n3796
g3733 and n2740 n3796 ; n3797
g3734 and n937 n3797 ; n3798
g3735 and n3757 n3798 ; n3799
g3736 and n1761 n3799 ; n3800
g3737 and n538 n3800 ; n3801
g3738 and n462_not n3801 ; n3802
g3739 and n402_not n3802 ; n3803
g3740 and n277_not n3803 ; n3804
g3741 and n293_not n3804 ; n3805
g3742 and n3457 n3805_not ; n3806
g3743 and n3542 n3605_not ; n3807
g3744 and n3456_not n3606 ; n3808
g3745 nor n3807 n3808 ; n3809
g3746 and n3806_not n3809 ; n3810
g3747 and n3368_not n3810 ; n3811
g3748 nor n3622 n3625 ; n3812
g3749 nor n3456 n3805 ; n3813
g3750 and n3456 n3805 ; n3814
g3751 nor n3813 n3814 ; n3815
g3752 and n3812_not n3815 ; n3816
g3753 and n3812 n3815_not ; n3817
g3754 nor n3816 n3817 ; n3818
g3755 and n3810 n3818_not ; n3819
g3756 nor n3811 n3819 ; n3820
g3757 and a[29] n3820_not ; n3821
g3758 and a[29]_not n3820 ; n3822
g3759 nor n3821 n3822 ; n3823
g3760 and n3727 n3823 ; n3824
g3761 nor n3727 n3823 ; n3825
g3762 nor n3824 n3825 ; n3826
g3763 nor n286 n438 ; n3827
g3764 and n3437 n3827 ; n3828
g3765 and n245_not n3828 ; n3829
g3766 and n791_not n3829 ; n3830
g3767 and n422_not n3830 ; n3831
g3768 nor n298 n961 ; n3832
g3769 and n3831 n3832 ; n3833
g3770 and n665 n3833 ; n3834
g3771 and n539 n3834 ; n3835
g3772 and n454 n3835 ; n3836
g3773 and n193 n3836 ; n3837
g3774 and n99_not n3837 ; n3838
g3775 and n372_not n3838 ; n3839
g3776 and n772 n1105 ; n3840
g3777 and n471 n3840 ; n3841
g3778 and n827 n3841 ; n3842
g3779 and n657_not n3842 ; n3843
g3780 and n252_not n3843 ; n3844
g3781 and n592_not n3844 ; n3845
g3782 and n277_not n3845 ; n3846
g3783 and n332_not n3846 ; n3847
g3784 and n1127_not n3847 ; n3848
g3785 and n2208 n2573 ; n3849
g3786 and n128 n3849 ; n3850
g3787 and n489_not n3850 ; n3851
g3788 and n119_not n3851 ; n3852
g3789 and n2275 n3852 ; n3853
g3790 and n3848 n3853 ; n3854
g3791 and n86_not n3854 ; n3855
g3792 and n569_not n3855 ; n3856
g3793 and n429_not n590 ; n3857
g3794 and n231_not n3857 ; n3858
g3795 and n624 n3206 ; n3859
g3796 and n2963 n3859 ; n3860
g3797 and n1254 n3860 ; n3861
g3798 and n979 n3861 ; n3862
g3799 and n356 n3862 ; n3863
g3800 and n289_not n3863 ; n3864
g3801 and n284_not n3864 ; n3865
g3802 and n557_not n3865 ; n3866
g3803 and n3858 n3866 ; n3867
g3804 and n633_not n3867 ; n3868
g3805 and n270_not n3868 ; n3869
g3806 and n3570 n3869 ; n3870
g3807 and n1480 n3870 ; n3871
g3808 and n968 n3871 ; n3872
g3809 and n449_not n3872 ; n3873
g3810 and n3856 n3873 ; n3874
g3811 and n3839 n3874 ; n3875
g3812 and n328_not n3875 ; n3876
g3813 and n296_not n3876 ; n3877
g3814 and a[23] a[24]_not ; n3878
g3815 and a[23]_not a[24] ; n3879
g3816 nor n3878 n3879 ; n3880
g3817 and a[25] a[26]_not ; n3881
g3818 and a[25]_not a[26] ; n3882
g3819 nor n3881 n3882 ; n3883
g3820 and n3880_not n3883 ; n3884
g3821 and n3877_not n3884 ; n3885
g3822 nor n127 n277 ; n3886
g3823 and n2390 n3041 ; n3887
g3824 and n2633 n3887 ; n3888
g3825 and n1479 n3888 ; n3889
g3826 and n1824 n3889 ; n3890
g3827 and n3886 n3890 ; n3891
g3828 and n190_not n3891 ; n3892
g3829 and n847_not n3892 ; n3893
g3830 and n777_not n3893 ; n3894
g3831 and n492_not n3894 ; n3895
g3832 and n163_not n3895 ; n3896
g3833 and n170_not n3896 ; n3897
g3834 and n340_not n3897 ; n3898
g3835 and n672_not n3898 ; n3899
g3836 and n436_not n3899 ; n3900
g3837 and n358_not n3900 ; n3901
g3838 nor n111 n505 ; n3902
g3839 and n394_not n3902 ; n3903
g3840 and n375_not n3903 ; n3904
g3841 and n883_not n3904 ; n3905
g3842 and n747 n978 ; n3906
g3843 nor n236 n301 ; n3907
g3844 and n136_not n3907 ; n3908
g3845 and n469_not n3908 ; n3909
g3846 and n1306_not n3909 ; n3910
g3847 and n397_not n3910 ; n3911
g3848 and n398_not n3911 ; n3912
g3849 and n775 n3912 ; n3913
g3850 and n1072_not n3913 ; n3914
g3851 and n517 n3914 ; n3915
g3852 and n3906 n3915 ; n3916
g3853 and n732 n3916 ; n3917
g3854 and n3905 n3917 ; n3918
g3855 and n3901 n3918 ; n3919
g3856 and n1731 n3919 ; n3920
g3857 and n617_not n3920 ; n3921
g3858 and n490_not n3921 ; n3922
g3859 and n425_not n3922 ; n3923
g3860 and n468_not n3923 ; n3924
g3861 and n273_not n3924 ; n3925
g3862 and n295_not n3925 ; n3926
g3863 and n532_not n3926 ; n3927
g3864 and n886_not n3927 ; n3928
g3865 and n569_not n3928 ; n3929
g3866 and n330_not n2738 ; n3930
g3867 and n242_not n3930 ; n3931
g3868 and n2698 n3931 ; n3932
g3869 and n504_not n3932 ; n3933
g3870 and n245_not n3933 ; n3934
g3871 and n142_not n3934 ; n3935
g3872 and n791_not n3935 ; n3936
g3873 and n567_not n3936 ; n3937
g3874 and n271_not n3937 ; n3938
g3875 and n771_not n3938 ; n3939
g3876 and n1440 n3729 ; n3940
g3877 and n3409 n3940 ; n3941
g3878 and n1292 n3941 ; n3942
g3879 and n276_not n3942 ; n3943
g3880 and n168_not n3943 ; n3944
g3881 and n426_not n3944 ; n3945
g3882 and n1102_not n3945 ; n3946
g3883 and n511_not n3946 ; n3947
g3884 and n372_not n1480 ; n3948
g3885 and n449_not n3948 ; n3949
g3886 and n1155 n3949 ; n3950
g3887 and n3947 n3950 ; n3951
g3888 and n2740 n3951 ; n3952
g3889 and n3939 n3952 ; n3953
g3890 and n3929 n3953 ; n3954
g3891 and n1046 n3954 ; n3955
g3892 and n520 n3955 ; n3956
g3893 and n2583 n3956 ; n3957
g3894 and n720 n3957 ; n3958
g3895 and n1011_not n3958 ; n3959
g3896 and n980_not n3959 ; n3960
g3897 and n452_not n3960 ; n3961
g3898 and n536_not n3961 ; n3962
g3899 and n283_not n3962 ; n3963
g3900 and n338_not n3963 ; n3964
g3901 nor n76 n84 ; n3965
g3902 and n3880 n3883_not ; n3966
g3903 and n3965_not n3966 ; n3967
g3904 and n3964_not n3967 ; n3968
g3905 nor n492 n496 ; n3969
g3906 and n430_not n3969 ; n3970
g3907 and n505_not n3970 ; n3971
g3908 and n425_not n3971 ; n3972
g3909 and n2470 n3832 ; n3973
g3910 and n619_not n3973 ; n3974
g3911 and n237_not n3974 ; n3975
g3912 and n712_not n3975 ; n3976
g3913 and n451_not n3976 ; n3977
g3914 and n592_not n3977 ; n3978
g3915 and n1478 n1726 ; n3979
g3916 and n327_not n3979 ; n3980
g3917 and n91_not n3980 ; n3981
g3918 and n715_not n3981 ; n3982
g3919 and n102_not n3982 ; n3983
g3920 and n287_not n3983 ; n3984
g3921 nor n290 n884 ; n3985
g3922 and n147_not n3985 ; n3986
g3923 and n403_not n3986 ; n3987
g3924 and n1347 n3987 ; n3988
g3925 and n155_not n3988 ; n3989
g3926 and n396_not n3989 ; n3990
g3927 and n1916 n2297 ; n3991
g3928 and n149_not n3991 ; n3992
g3929 and n594_not n3992 ; n3993
g3930 and n223_not n3993 ; n3994
g3931 and n402_not n3994 ; n3995
g3932 and n305_not n3995 ; n3996
g3933 and n226_not n3996 ; n3997
g3934 and n3990 n3997 ; n3998
g3935 and n538 n3998 ; n3999
g3936 and n435_not n3999 ; n4000
g3937 and n292_not n4000 ; n4001
g3938 and n283_not n4001 ; n4002
g3939 and n372_not n4002 ; n4003
g3940 and n2133 n2703 ; n4004
g3941 and n2739 n4004 ; n4005
g3942 and n1248 n4005 ; n4006
g3943 and n1389 n4006 ; n4007
g3944 and n506_not n4007 ; n4008
g3945 and n107_not n4008 ; n4009
g3946 and n275_not n2993 ; n4010
g3947 and n417_not n4010 ; n4011
g3948 and n3408 n4011 ; n4012
g3949 and n4009 n4012 ; n4013
g3950 and n4003 n4013 ; n4014
g3951 and n1783 n4014 ; n4015
g3952 and n421 n4015 ; n4016
g3953 and n453_not n4016 ; n4017
g3954 and n3914 n3931 ; n4018
g3955 and n3128 n4018 ; n4019
g3956 and n3947 n4019 ; n4020
g3957 and n123_not n4020 ; n4021
g3958 and n194_not n4021 ; n4022
g3959 and n111_not n4022 ; n4023
g3960 and n746_not n4023 ; n4024
g3961 and n462_not n4024 ; n4025
g3962 and n509_not n4025 ; n4026
g3963 and n1011_not n4026 ; n4027
g3964 and n190_not n4027 ; n4028
g3965 and n518_not n4028 ; n4029
g3966 and n151_not n4029 ; n4030
g3967 and n4017 n4030 ; n4031
g3968 and n3984 n4031 ; n4032
g3969 and n825_not n4032 ; n4033
g3970 and n99_not n4033 ; n4034
g3971 and n1204 n3852 ; n4035
g3972 and n3790 n4035 ; n4036
g3973 and n604 n4036 ; n4037
g3974 and n1046 n4037 ; n4038
g3975 and n159 n4038 ; n4039
g3976 and n130_not n4039 ; n4040
g3977 and n4034 n4040 ; n4041
g3978 and n3978 n4041 ; n4042
g3979 and n3972 n4042 ; n4043
g3980 and n471 n4043 ; n4044
g3981 and n589_not n4044 ; n4045
g3982 and n3880 n3965 ; n4046
g3983 and n4045_not n4046 ; n4047
g3984 nor n3968 n4047 ; n4048
g3985 and n3885_not n4048 ; n4049
g3986 nor n3880 n3883 ; n4050
g3987 nor n3964 n4045 ; n4051
g3988 nor n3805 n3964 ; n4052
g3989 nor n3813 n3816 ; n4053
g3990 and n3805 n3964 ; n4054
g3991 nor n4052 n4054 ; n4055
g3992 and n4053_not n4055 ; n4056
g3993 nor n4052 n4056 ; n4057
g3994 and n3964 n4045 ; n4058
g3995 nor n4051 n4058 ; n4059
g3996 and n4057_not n4059 ; n4060
g3997 nor n4051 n4060 ; n4061
g3998 nor n3877 n4045 ; n4062
g3999 and n3877 n4045 ; n4063
g4000 nor n4062 n4063 ; n4064
g4001 and n4061_not n4064 ; n4065
g4002 and n4061 n4064_not ; n4066
g4003 nor n4065 n4066 ; n4067
g4004 and n4050 n4067 ; n4068
g4005 and n4049 n4068_not ; n4069
g4006 and a[26] n4069_not ; n4070
g4007 and a[26] n4070_not ; n4071
g4008 nor n4069 n4070 ; n4072
g4009 nor n4071 n4072 ; n4073
g4010 and n3826 n4073_not ; n4074
g4011 and n3826 n4074_not ; n4075
g4012 nor n4073 n4074 ; n4076
g4013 nor n4075 n4076 ; n4077
g4014 and n3457 n3605_not ; n4078
g4015 and n3012_not n3542 ; n4079
g4016 and n3539_not n3606 ; n4080
g4017 nor n4079 n4080 ; n4081
g4018 and n4078_not n4081 ; n4082
g4019 and n3617 n3619_not ; n4083
g4020 nor n3620 n4083 ; n4084
g4021 and n3368 n4084 ; n4085
g4022 and n4082 n4085_not ; n4086
g4023 and a[29] n4086_not ; n4087
g4024 nor n4086 n4087 ; n4088
g4025 and a[29] n4087_not ; n4089
g4026 nor n4088 n4089 ; n4090
g4027 nor n3354 n3357 ; n4091
g4028 and n3356 n3357_not ; n4092
g4029 nor n4091 n4092 ; n4093
g4030 nor n4090 n4093 ; n4094
g4031 nor n4090 n4094 ; n4095
g4032 nor n4093 n4094 ; n4096
g4033 nor n4095 n4096 ; n4097
g4034 nor n3338 n3340 ; n4098
g4035 and n3329_not n3341 ; n4099
g4036 nor n4098 n4099 ; n4100
g4037 nor n395 n594 ; n4101
g4038 nor n354 n1011 ; n4102
g4039 and n177_not n4102 ; n4103
g4040 and n367_not n4103 ; n4104
g4041 and n250 n1760 ; n4105
g4042 and n792 n4105 ; n4106
g4043 and n2192 n4106 ; n4107
g4044 and n4104 n4107 ; n4108
g4045 and n2943 n4108 ; n4109
g4046 and n877 n4109 ; n4110
g4047 and n2217 n4110 ; n4111
g4048 and n3405 n4111 ; n4112
g4049 and n3901 n4112 ; n4113
g4050 and n2500 n4113 ; n4114
g4051 and n1183 n4114 ; n4115
g4052 and n507 n4115 ; n4116
g4053 and n4101 n4116 ; n4117
g4054 and n327_not n4117 ; n4118
g4055 and n292_not n4118 ; n4119
g4056 and n286_not n4119 ; n4120
g4057 and n1104_not n4120 ; n4121
g4058 and n395_not n1073 ; n4122
g4059 and n980_not n4122 ; n4123
g4060 and n165_not n4123 ; n4124
g4061 and n932_not n4124 ; n4125
g4062 and n375_not n4125 ; n4126
g4063 and n86_not n4126 ; n4127
g4064 and n1139 n1781 ; n4128
g4065 and n242_not n4128 ; n4129
g4066 and n562_not n4129 ; n4130
g4067 and n402_not n1181 ; n4131
g4068 and n416_not n4131 ; n4132
g4069 and n1045 n4132 ; n4133
g4070 and n812 n4133 ; n4134
g4071 and n1692 n4134 ; n4135
g4072 and n4130 n4135 ; n4136
g4073 and n4127 n4136 ; n4137
g4074 and n491 n4137 ; n4138
g4075 and n1251 n4138 ; n4139
g4076 and n1141 n4139 ; n4140
g4077 and n123_not n4140 ; n4141
g4078 and n334_not n4141 ; n4142
g4079 and n1101_not n4142 ; n4143
g4080 and n594_not n4143 ; n4144
g4081 and n527_not n4144 ; n4145
g4082 and n689_not n4145 ; n4146
g4083 and n200_not n4146 ; n4147
g4084 and n1104_not n4147 ; n4148
g4085 nor n168 n1203 ; n4149
g4086 and n886_not n4149 ; n4150
g4087 and n188_not n4150 ; n4151
g4088 and n279 n589_not ; n4152
g4089 and n394_not n4152 ; n4153
g4090 and n4151 n4153 ; n4154
g4091 and n2371 n4154 ; n4155
g4092 and n3521 n4155 ; n4156
g4093 and n4148 n4156 ; n4157
g4094 and n3408 n4157 ; n4158
g4095 and n773 n4158 ; n4159
g4096 and n235 n4159 ; n4160
g4097 and n454 n4160 ; n4161
g4098 and n1040 n4161 ; n4162
g4099 and n397_not n4162 ; n4163
g4100 and n354_not n4163 ; n4164
g4101 and n1102_not n4164 ; n4165
g4102 and n327_not n4165 ; n4166
g4103 and n403_not n4166 ; n4167
g4104 and n1524 n4167 ; n4168
g4105 and n326_not n4168 ; n4169
g4106 and n438_not n4169 ; n4170
g4107 and n201_not n4170 ; n4171
g4108 nor n4121 n4171 ; n4172
g4109 and n4121 n4171 ; n4173
g4110 nor n4172 n4173 ; n4174
g4111 and a[17]_not n4174 ; n4175
g4112 nor n4172 n4175 ; n4176
g4113 and n3146 n4176_not ; n4177
g4114 and n2916 n2918_not ; n4178
g4115 nor n2919 n4178 ; n4179
g4116 and n75 n4179 ; n4180
g4117 and n710_not n3020 ; n4181
g4118 and n958_not n3023 ; n4182
g4119 and n867_not n3028 ; n4183
g4120 nor n4182 n4183 ; n4184
g4121 and n4181_not n4184 ; n4185
g4122 and n4180_not n4185 ; n4186
g4123 and n3146_not n4176 ; n4187
g4124 nor n4177 n4187 ; n4188
g4125 and n4186_not n4188 ; n4189
g4126 nor n4177 n4189 ; n4190
g4127 nor n4100 n4190 ; n4191
g4128 and n4100 n4190 ; n4192
g4129 nor n4191 n4192 ; n4193
g4130 nor n4186 n4189 ; n4194
g4131 and n4188 n4189_not ; n4195
g4132 nor n4194 n4195 ; n4196
g4133 nor a[17] n4175 ; n4197
g4134 and n4173_not n4176 ; n4198
g4135 nor n4197 n4198 ; n4199
g4136 and n867_not n3020 ; n4200
g4137 and n958_not n3028 ; n4201
g4138 and n1060_not n3023 ; n4202
g4139 and n2912 n2914_not ; n4203
g4140 nor n2915 n4203 ; n4204
g4141 and n75 n4204 ; n4205
g4142 nor n4202 n4205 ; n4206
g4143 and n4201_not n4206 ; n4207
g4144 and n4200_not n4207 ; n4208
g4145 nor n4199 n4208 ; n4209
g4146 and n2348 n2515 ; n4210
g4147 and n977 n4210 ; n4211
g4148 and n2090 n4211 ; n4212
g4149 and n95_not n4212 ; n4213
g4150 and n363_not n4213 ; n4214
g4151 and n449_not n4214 ; n4215
g4152 nor n396 n430 ; n4216
g4153 nor n236 n1127 ; n4217
g4154 and n875_not n4217 ; n4218
g4155 and n3085 n4218 ; n4219
g4156 and n4216 n4219 ; n4220
g4157 and n2132 n4220 ; n4221
g4158 and n2301 n4221 ; n4222
g4159 and n2202 n4222 ; n4223
g4160 and n805 n4223 ; n4224
g4161 and n399 n4224 ; n4225
g4162 and n227 n4225 ; n4226
g4163 and n885 n4226 ; n4227
g4164 and n136_not n4227 ; n4228
g4165 and n667_not n4228 ; n4229
g4166 and n1102_not n4229 ; n4230
g4167 and n189_not n4230 ; n4231
g4168 and n712_not n4231 ; n4232
g4169 and n496_not n2468 ; n4233
g4170 and n883_not n4233 ; n4234
g4171 and n3827 n4234 ; n4235
g4172 and n778 n4235 ; n4236
g4173 and n2017 n4236 ; n4237
g4174 and n2740 n4237 ; n4238
g4175 and n156 n4238 ; n4239
g4176 and n123_not n4239 ; n4240
g4177 and n353_not n4240 ; n4241
g4178 and n115_not n4241 ; n4242
g4179 and n233_not n4242 ; n4243
g4180 and n639_not n4243 ; n4244
g4181 and n425_not n4244 ; n4245
g4182 and n99_not n4245 ; n4246
g4183 and n306_not n4246 ; n4247
g4184 and n541 n2241 ; n4248
g4185 and n2330 n4248 ; n4249
g4186 and n2507 n4249 ; n4250
g4187 and n4247 n4250 ; n4251
g4188 and n4232 n4251 ; n4252
g4189 and n4215 n4252 ; n4253
g4190 and n2635 n4253 ; n4254
g4191 and n2682 n4254 ; n4255
g4192 and n1781 n4255 ; n4256
g4193 and n427_not n4256 ; n4257
g4194 and n461_not n4257 ; n4258
g4195 and n228_not n4258 ; n4259
g4196 and n326_not n4259 ; n4260
g4197 and n395_not n4260 ; n4261
g4198 and n714_not n4261 ; n4262
g4199 and n304_not n4262 ; n4263
g4200 and n666_not n4263 ; n4264
g4201 and n886_not n4264 ; n4265
g4202 and n771_not n4265 ; n4266
g4203 and n4121 n4266_not ; n4267
g4204 and n4121_not n4266 ; n4268
g4205 nor n150 n155 ; n4269
g4206 and n250 n4269 ; n4270
g4207 and n752_not n4270 ; n4271
g4208 and n402_not n4271 ; n4272
g4209 and n430_not n4272 ; n4273
g4210 and n428_not n4273 ; n4274
g4211 nor n276 n419 ; n4275
g4212 and n403_not n4275 ; n4276
g4213 and n424_not n4276 ; n4277
g4214 and n170_not n4277 ; n4278
g4215 and n883_not n4278 ; n4279
g4216 and n1944 n2684 ; n4280
g4217 and n4279 n4280 ; n4281
g4218 and n4215 n4281 ; n4282
g4219 and n4274 n4282 ; n4283
g4220 and n1917 n4283 ; n4284
g4221 and n773 n4284 ; n4285
g4222 and n1237 n4285 ; n4286
g4223 and n278_not n4286 ; n4287
g4224 and n305_not n4287 ; n4288
g4225 and n146_not n4288 ; n4289
g4226 and n102_not n4289 ; n4290
g4227 and n932_not n4290 ; n4291
g4228 and n200_not n4291 ; n4292
g4229 and n371_not n4292 ; n4293
g4230 nor n339 n374 ; n4294
g4231 and n338_not n4294 ; n4295
g4232 nor n99 n330 ; n4296
g4233 and n157_not n4296 ; n4297
g4234 and n470_not n4297 ; n4298
g4235 and n1047 n2637 ; n4299
g4236 and n4218 n4299 ; n4300
g4237 and n4298 n4300 ; n4301
g4238 and n3464 n4301 ; n4302
g4239 and n2738 n4302 ; n4303
g4240 and n4295 n4303 ; n4304
g4241 and n123_not n4304 ; n4305
g4242 and n558_not n4305 ; n4306
g4243 and n149_not n4306 ; n4307
g4244 and n527_not n4307 ; n4308
g4245 and n504_not n4308 ; n4309
g4246 and n273_not n4309 ; n4310
g4247 and n564_not n4310 ; n4311
g4248 nor n135 n452 ; n4312
g4249 and n283_not n4312 ; n4313
g4250 and n941 n4313 ; n4314
g4251 and n1602 n4314 ; n4315
g4252 and n154_not n4315 ; n4316
g4253 and n619_not n4316 ; n4317
g4254 and n121_not n4317 ; n4318
g4255 and n594_not n4318 ; n4319
g4256 and n396_not n4319 ; n4320
g4257 and n777_not n4320 ; n4321
g4258 and n326_not n4321 ; n4322
g4259 and n425_not n4322 ; n4323
g4260 and n298_not n4323 ; n4324
g4261 and n791_not n4324 ; n4325
g4262 nor n274 n426 ; n4326
g4263 and n633_not n4326 ; n4327
g4264 and n2371 n4327 ; n4328
g4265 and n2073 n4328 ; n4329
g4266 and n511_not n4329 ; n4330
g4267 and n656_not n4330 ; n4331
g4268 and n657_not n4331 ; n4332
g4269 nor n192 n509 ; n4333
g4270 and n340_not n4333 ; n4334
g4271 nor n233 n715 ; n4335
g4272 and n3114 n4335 ; n4336
g4273 and n4334 n4336 ; n4337
g4274 and n4332 n4337 ; n4338
g4275 and n2740 n4338 ; n4339
g4276 and n2169 n4339 ; n4340
g4277 and n4325 n4340 ; n4341
g4278 and n4311 n4341 ; n4342
g4279 and n4293 n4342 ; n4343
g4280 and n491 n4343 ; n4344
g4281 and n1182 n4344 ; n4345
g4282 and n118_not n4345 ; n4346
g4283 and n689_not n4346 ; n4347
g4284 and n277_not n4347 ; n4348
g4285 and n672_not n4348 ; n4349
g4286 and n86_not n4349 ; n4350
g4287 and n188_not n4350 ; n4351
g4288 and n1246_not n1669 ; n4352
g4289 and n289_not n4352 ; n4353
g4290 and n461_not n4353 ; n4354
g4291 and n363_not n4354 ; n4355
g4292 and n562_not n4355 ; n4356
g4293 nor n673 n1306 ; n4357
g4294 and n1135 n2334 ; n4358
g4295 and n4357 n4358 ; n4359
g4296 and n1040 n4359 ; n4360
g4297 and n232_not n4360 ; n4361
g4298 and n255_not n4361 ; n4362
g4299 and n203_not n4362 ; n4363
g4300 and n809_not n4363 ; n4364
g4301 and n239_not n4364 ; n4365
g4302 and n372_not n4365 ; n4366
g4303 nor n102 n293 ; n4367
g4304 and n876 n2210 ; n4368
g4305 and n4153 n4368 ; n4369
g4306 and n2013 n4369 ; n4370
g4307 and n2807 n4370 ; n4371
g4308 and n4367 n4371 ; n4372
g4309 and n169_not n4372 ; n4373
g4310 and n190_not n4373 ; n4374
g4311 and n435_not n4374 ; n4375
g4312 and n1272 n4234 ; n4376
g4313 and n439 n4376 ; n4377
g4314 and n4375 n4377 ; n4378
g4315 and n3378 n4378 ; n4379
g4316 and n1550 n4379 ; n4380
g4317 and n427_not n4380 ; n4381
g4318 and n420_not n4381 ; n4382
g4319 and n146_not n4382 ; n4383
g4320 and n296_not n4383 ; n4384
g4321 and n980_not n4384 ; n4385
g4322 and n201_not n4385 ; n4386
g4323 and n271_not n4386 ; n4387
g4324 and n249_not n4387 ; n4388
g4325 and n793 n3296 ; n4389
g4326 and n2296 n4389 ; n4390
g4327 and n615 n4390 ; n4391
g4328 and n1330 n4391 ; n4392
g4329 and n827 n4392 ; n4393
g4330 and n978 n4393 ; n4394
g4331 and n590 n4394 ; n4395
g4332 and n667_not n4395 ; n4396
g4333 and n355_not n4396 ; n4397
g4334 and n152_not n4397 ; n4398
g4335 and n511_not n4398 ; n4399
g4336 and n594_not n4399 ; n4400
g4337 and n637_not n4400 ; n4401
g4338 and n107_not n4401 ; n4402
g4339 and n601_not n4402 ; n4403
g4340 and n603_not n4403 ; n4404
g4341 and n338_not n4404 ; n4405
g4342 and n2014 n3416 ; n4406
g4343 and n1346 n4406 ; n4407
g4344 and n992 n4407 ; n4408
g4345 and n1785 n4408 ; n4409
g4346 and n4405 n4409 ; n4410
g4347 and n4388 n4410 ; n4411
g4348 and n4366 n4411 ; n4412
g4349 and n4356 n4412 ; n4413
g4350 and n774 n4413 ; n4414
g4351 and n2698 n4414 ; n4415
g4352 and n285 n4415 ; n4416
g4353 and n236_not n4416 ; n4417
g4354 and n397_not n4417 ; n4418
g4355 and n335_not n4418 ; n4419
g4356 and n563_not n4419 ; n4420
g4357 and n489_not n4420 ; n4421
g4358 nor n4351 n4421 ; n4422
g4359 and n4351 n4421 ; n4423
g4360 nor n4422 n4423 ; n4424
g4361 and a[14]_not n4424 ; n4425
g4362 nor n4422 n4425 ; n4426
g4363 and n4266 n4426_not ; n4427
g4364 and n2904 n2906_not ; n4428
g4365 nor n2907 n4428 ; n4429
g4366 and n75 n4429 ; n4430
g4367 and n1060_not n3020 ; n4431
g4368 and n1235_not n3023 ; n4432
g4369 and n1178_not n3028 ; n4433
g4370 nor n4432 n4433 ; n4434
g4371 and n4431_not n4434 ; n4435
g4372 and n4430_not n4435 ; n4436
g4373 and n4266_not n4426 ; n4437
g4374 nor n4427 n4437 ; n4438
g4375 and n4436_not n4438 ; n4439
g4376 nor n4427 n4439 ; n4440
g4377 nor n4267 n4440 ; n4441
g4378 and n4268_not n4441 ; n4442
g4379 nor n4267 n4442 ; n4443
g4380 and n4199 n4208 ; n4444
g4381 nor n4209 n4444 ; n4445
g4382 and n4443_not n4445 ; n4446
g4383 nor n4209 n4446 ; n4447
g4384 nor n4196 n4447 ; n4448
g4385 and n4196 n4447 ; n4449
g4386 nor n4448 n4449 ; n4450
g4387 and n3012_not n3457 ; n4451
g4388 and n587_not n3542 ; n4452
g4389 and n392_not n3606 ; n4453
g4390 nor n4452 n4453 ; n4454
g4391 and n4451_not n4454 ; n4455
g4392 and n3368_not n4455 ; n4456
g4393 and n3018_not n4455 ; n4457
g4394 nor n4456 n4457 ; n4458
g4395 and a[29] n4458_not ; n4459
g4396 and a[29]_not n4458 ; n4460
g4397 nor n4459 n4460 ; n4461
g4398 and n4450 n4461_not ; n4462
g4399 nor n4448 n4462 ; n4463
g4400 and n4193 n4463_not ; n4464
g4401 nor n4191 n4464 ; n4465
g4402 nor n4097 n4465 ; n4466
g4403 nor n4094 n4466 ; n4467
g4404 and n3361_not n3632 ; n4468
g4405 nor n3633 n4468 ; n4469
g4406 and n4467_not n4469 ; n4470
g4407 and n3884 n4045_not ; n4471
g4408 and n3805_not n3967 ; n4472
g4409 and n3964_not n4046 ; n4473
g4410 nor n4472 n4473 ; n4474
g4411 and n4471_not n4474 ; n4475
g4412 and n4057 n4059_not ; n4476
g4413 nor n4060 n4476 ; n4477
g4414 and n4050 n4477 ; n4478
g4415 and n4475 n4478_not ; n4479
g4416 and a[26] n4479_not ; n4480
g4417 nor n4479 n4480 ; n4481
g4418 and a[26] n4480_not ; n4482
g4419 nor n4481 n4482 ; n4483
g4420 nor n4467 n4470 ; n4484
g4421 and n4469 n4470_not ; n4485
g4422 nor n4484 n4485 ; n4486
g4423 nor n4483 n4486 ; n4487
g4424 nor n4470 n4487 ; n4488
g4425 and n714_not n2014 ; n4489
g4426 and n243_not n4489 ; n4490
g4427 and n145_not n4490 ; n4491
g4428 and n466_not n4491 ; n4492
g4429 and n205_not n4492 ; n4493
g4430 and n1388 n1785 ; n4494
g4431 and n604 n4494 ; n4495
g4432 and n2170 n4495 ; n4496
g4433 and n173_not n4496 ; n4497
g4434 and n144_not n4497 ; n4498
g4435 and n394_not n4498 ; n4499
g4436 and n306_not n4499 ; n4500
g4437 and n157_not n4500 ; n4501
g4438 and n375_not n4501 ; n4502
g4439 and n133 n4502 ; n4503
g4440 and n4493 n4503 ; n4504
g4441 and n2346 n4504 ; n4505
g4442 and n1046 n4505 ; n4506
g4443 and n1761 n4506 ; n4507
g4444 and n1367 n4507 ; n4508
g4445 and n274_not n4508 ; n4509
g4446 and n589_not n4509 ; n4510
g4447 and n468_not n4510 ; n4511
g4448 and n3972 n4511 ; n4512
g4449 and n296_not n4512 ; n4513
g4450 and n601_not n4513 ; n4514
g4451 and n3839 n4514 ; n4515
g4452 nor n4062 n4065 ; n4516
g4453 nor n3877 n4515 ; n4517
g4454 and n3877 n4515 ; n4518
g4455 nor n4517 n4518 ; n4519
g4456 and n4516_not n4519 ; n4520
g4457 and n3877 n4520_not ; n4521
g4458 nor n4515 n4521 ; n4522
g4459 and a[21]_not a[22] ; n4523
g4460 and a[21] a[22]_not ; n4524
g4461 nor n4523 n4524 ; n4525
g4462 and a[20] a[21]_not ; n4526
g4463 and a[20]_not a[21] ; n4527
g4464 nor n4526 n4527 ; n4528
g4465 and a[22]_not a[23] ; n4529
g4466 and a[22] a[23]_not ; n4530
g4467 nor n4529 n4530 ; n4531
g4468 and n4528 n4531_not ; n4532
g4469 and n4525 n4532 ; n4533
g4470 and n4515_not n4533 ; n4534
g4471 nor n4522 n4534 ; n4535
g4472 nor n4528 n4531 ; n4536
g4473 nor n4534 n4536 ; n4537
g4474 nor n4535 n4537 ; n4538
g4475 and a[23] n4538_not ; n4539
g4476 and a[23]_not n4538 ; n4540
g4477 nor n4539 n4540 ; n4541
g4478 nor n4488 n4541 ; n4542
g4479 and n4488 n4541 ; n4543
g4480 nor n4542 n4543 ; n4544
g4481 and n4077_not n4544 ; n4545
g4482 nor n4077 n4545 ; n4546
g4483 and n4544 n4545_not ; n4547
g4484 nor n4546 n4547 ; n4548
g4485 and n4097 n4465 ; n4549
g4486 nor n4466 n4549 ; n4550
g4487 and n3884 n3964_not ; n4551
g4488 and n3456_not n3967 ; n4552
g4489 and n3805_not n4046 ; n4553
g4490 nor n4552 n4553 ; n4554
g4491 and n4551_not n4554 ; n4555
g4492 and n4050_not n4555 ; n4556
g4493 and n4053 n4055_not ; n4557
g4494 nor n4056 n4557 ; n4558
g4495 and n4555 n4558_not ; n4559
g4496 nor n4556 n4559 ; n4560
g4497 and a[26] n4560_not ; n4561
g4498 and a[26]_not n4560 ; n4562
g4499 nor n4561 n4562 ; n4563
g4500 and n4550 n4563_not ; n4564
g4501 and n3805_not n3884 ; n4565
g4502 and n3605_not n3967 ; n4566
g4503 and n3456_not n4046 ; n4567
g4504 nor n4566 n4567 ; n4568
g4505 and n4565_not n4568 ; n4569
g4506 and n3818 n4050 ; n4570
g4507 and n4569 n4570_not ; n4571
g4508 and a[26] n4571_not ; n4572
g4509 and a[26] n4572_not ; n4573
g4510 nor n4571 n4572 ; n4574
g4511 nor n4573 n4574 ; n4575
g4512 and n4193_not n4463 ; n4576
g4513 nor n4464 n4576 ; n4577
g4514 and n3457 n3539_not ; n4578
g4515 and n392_not n3542 ; n4579
g4516 and n3012_not n3606 ; n4580
g4517 nor n4579 n4580 ; n4581
g4518 and n4578_not n4581 ; n4582
g4519 and n3368_not n4582 ; n4583
g4520 and n3715_not n4582 ; n4584
g4521 nor n4583 n4584 ; n4585
g4522 and a[29] n4585_not ; n4586
g4523 and a[29]_not n4585 ; n4587
g4524 nor n4586 n4587 ; n4588
g4525 and n4577 n4588_not ; n4589
g4526 and n4577_not n4588 ; n4590
g4527 nor n4589 n4590 ; n4591
g4528 and n4575_not n4591 ; n4592
g4529 nor n4589 n4592 ; n4593
g4530 and n4550 n4564_not ; n4594
g4531 nor n4563 n4564 ; n4595
g4532 nor n4594 n4595 ; n4596
g4533 nor n4593 n4596 ; n4597
g4534 nor n4564 n4597 ; n4598
g4535 and n4483 n4485_not ; n4599
g4536 and n4484_not n4599 ; n4600
g4537 nor n4487 n4600 ; n4601
g4538 and n4598_not n4601 ; n4602
g4539 and n3877_not n4533 ; n4603
g4540 and n4525_not n4528 ; n4604
g4541 and n4515_not n4604 ; n4605
g4542 nor n4603 n4605 ; n4606
g4543 nor n4517 n4520 ; n4607
g4544 and n4515 n4607 ; n4608
g4545 nor n4522 n4608 ; n4609
g4546 and n4536 n4609 ; n4610
g4547 and n4606 n4610_not ; n4611
g4548 and a[23] n4611_not ; n4612
g4549 nor n4611 n4612 ; n4613
g4550 and a[23] n4612_not ; n4614
g4551 nor n4613 n4614 ; n4615
g4552 and n4598 n4601_not ; n4616
g4553 nor n4602 n4616 ; n4617
g4554 and n4615_not n4617 ; n4618
g4555 nor n4602 n4618 ; n4619
g4556 and n4548 n4619 ; n4620
g4557 nor n4548 n4619 ; n4621
g4558 nor n4620 n4621 ; n4622
g4559 and n4591 n4592_not ; n4623
g4560 nor n4575 n4592 ; n4624
g4561 nor n4623 n4624 ; n4625
g4562 nor n4440 n4442 ; n4626
g4563 and n4268_not n4443 ; n4627
g4564 nor n4626 n4627 ; n4628
g4565 and n958_not n3020 ; n4629
g4566 and n1060_not n3028 ; n4630
g4567 and n1178_not n3023 ; n4631
g4568 and n2908 n2910_not ; n4632
g4569 nor n2911 n4632 ; n4633
g4570 and n75 n4633 ; n4634
g4571 nor n4631 n4634 ; n4635
g4572 and n4630_not n4635 ; n4636
g4573 and n4629_not n4636 ; n4637
g4574 nor n4628 n4637 ; n4638
g4575 and n587_not n3457 ; n4639
g4576 and n867_not n3542 ; n4640
g4577 and n710_not n3606 ; n4641
g4578 nor n4640 n4641 ; n4642
g4579 and n4639_not n4642 ; n4643
g4580 and n3331 n3368 ; n4644
g4581 and n4643 n4644_not ; n4645
g4582 and a[29] n4645_not ; n4646
g4583 nor n4645 n4646 ; n4647
g4584 and a[29] n4646_not ; n4648
g4585 nor n4647 n4648 ; n4649
g4586 nor n4628 n4638 ; n4650
g4587 nor n4637 n4638 ; n4651
g4588 nor n4650 n4651 ; n4652
g4589 nor n4649 n4652 ; n4653
g4590 nor n4638 n4653 ; n4654
g4591 and n4443 n4445_not ; n4655
g4592 nor n4446 n4655 ; n4656
g4593 and n4654_not n4656 ; n4657
g4594 and n392_not n3457 ; n4658
g4595 and n710_not n3542 ; n4659
g4596 and n587_not n3606 ; n4660
g4597 nor n4659 n4660 ; n4661
g4598 and n4658_not n4661 ; n4662
g4599 and n3347 n3368 ; n4663
g4600 and n4662 n4663_not ; n4664
g4601 and a[29] n4664_not ; n4665
g4602 and a[29] n4665_not ; n4666
g4603 nor n4664 n4665 ; n4667
g4604 nor n4666 n4667 ; n4668
g4605 and n4654 n4656_not ; n4669
g4606 nor n4657 n4669 ; n4670
g4607 and n4668_not n4670 ; n4671
g4608 nor n4657 n4671 ; n4672
g4609 and n4450_not n4461 ; n4673
g4610 nor n4462 n4673 ; n4674
g4611 and n4672_not n4674 ; n4675
g4612 and n4672 n4674_not ; n4676
g4613 nor n4675 n4676 ; n4677
g4614 and n3456_not n3884 ; n4678
g4615 and n3539_not n3967 ; n4679
g4616 and n3605_not n4046 ; n4680
g4617 nor n4679 n4680 ; n4681
g4618 and n4678_not n4681 ; n4682
g4619 and n3627 n4050 ; n4683
g4620 and n4682 n4683_not ; n4684
g4621 and a[26] n4684_not ; n4685
g4622 and a[26] n4685_not ; n4686
g4623 nor n4684 n4685 ; n4687
g4624 nor n4686 n4687 ; n4688
g4625 and n4677 n4688_not ; n4689
g4626 nor n4675 n4689 ; n4690
g4627 nor n4625 n4690 ; n4691
g4628 and n4625 n4690 ; n4692
g4629 nor n4691 n4692 ; n4693
g4630 and n4528_not n4531 ; n4694
g4631 and n3877_not n4694 ; n4695
g4632 and n3964_not n4533 ; n4696
g4633 and n4045_not n4604 ; n4697
g4634 nor n4696 n4697 ; n4698
g4635 and n4695_not n4698 ; n4699
g4636 and n4067 n4536 ; n4700
g4637 and n4699 n4700_not ; n4701
g4638 and a[23] n4701_not ; n4702
g4639 and a[23] n4702_not ; n4703
g4640 nor n4701 n4702 ; n4704
g4641 nor n4703 n4704 ; n4705
g4642 and n4693 n4705_not ; n4706
g4643 nor n4691 n4706 ; n4707
g4644 and n4515_not n4694 ; n4708
g4645 and n4045_not n4533 ; n4709
g4646 and n3877_not n4604 ; n4710
g4647 nor n4709 n4710 ; n4711
g4648 and n4708_not n4711 ; n4712
g4649 and n4536_not n4712 ; n4713
g4650 and n4516 n4519_not ; n4714
g4651 nor n4520 n4714 ; n4715
g4652 and n4712 n4715_not ; n4716
g4653 nor n4713 n4716 ; n4717
g4654 and a[23] n4717_not ; n4718
g4655 and a[23]_not n4717 ; n4719
g4656 nor n4718 n4719 ; n4720
g4657 nor n4707 n4720 ; n4721
g4658 and n4707 n4720 ; n4722
g4659 nor n4721 n4722 ; n4723
g4660 nor n4593 n4597 ; n4724
g4661 nor n4596 n4597 ; n4725
g4662 nor n4724 n4725 ; n4726
g4663 and n4723 n4726_not ; n4727
g4664 nor n4721 n4727 ; n4728
g4665 and n4615 n4617_not ; n4729
g4666 nor n4618 n4729 ; n4730
g4667 and n4728_not n4730 ; n4731
g4668 and n4723 n4727_not ; n4732
g4669 nor n4726 n4727 ; n4733
g4670 nor n4732 n4733 ; n4734
g4671 and n4677 n4689_not ; n4735
g4672 nor n4688 n4689 ; n4736
g4673 nor n4735 n4736 ; n4737
g4674 and n4670 n4671_not ; n4738
g4675 nor n4668 n4671 ; n4739
g4676 nor n4738 n4739 ; n4740
g4677 and n3605_not n3884 ; n4741
g4678 and n3012_not n3967 ; n4742
g4679 and n3539_not n4046 ; n4743
g4680 nor n4742 n4743 ; n4744
g4681 and n4741_not n4744 ; n4745
g4682 and n4050_not n4745 ; n4746
g4683 and n4084_not n4745 ; n4747
g4684 nor n4746 n4747 ; n4748
g4685 and a[26] n4748_not ; n4749
g4686 and a[26]_not n4748 ; n4750
g4687 nor n4749 n4750 ; n4751
g4688 nor n4740 n4751 ; n4752
g4689 nor n4649 n4653 ; n4753
g4690 nor n4652 n4653 ; n4754
g4691 nor n4753 n4754 ; n4755
g4692 nor n4436 n4439 ; n4756
g4693 and n4438 n4439_not ; n4757
g4694 nor n4756 n4757 ; n4758
g4695 nor a[14] n4425 ; n4759
g4696 and n4423_not n4426 ; n4760
g4697 nor n4759 n4760 ; n4761
g4698 and n617_not n3043 ; n4762
g4699 and n154_not n4762 ; n4763
g4700 and n641_not n4763 ; n4764
g4701 and n328_not n4764 ; n4765
g4702 and n394_not n4765 ; n4766
g4703 and n666_not n4766 ; n4767
g4704 and n564_not n3490 ; n4768
g4705 and n886_not n4768 ; n4769
g4706 and n333 n1389 ; n4770
g4707 and n449_not n4770 ; n4771
g4708 and n2361 n4771 ; n4772
g4709 and n4769 n4772 ; n4773
g4710 and n141 n4773 ; n4774
g4711 and n1181 n4774 ; n4775
g4712 and n874 n4775 ; n4776
g4713 and n968 n4776 ; n4777
g4714 and n3252 n4777 ; n4778
g4715 and n1827 n4778 ; n4779
g4716 and n2583 n4779 ; n4780
g4717 and n4101 n4780 ; n4781
g4718 and n169_not n4781 ; n4782
g4719 and n286_not n4782 ; n4783
g4720 and n589_not n4783 ; n4784
g4721 and n252_not n4784 ; n4785
g4722 nor n335 n367 ; n4786
g4723 nor n375 n511 ; n4787
g4724 and n304_not n4787 ; n4788
g4725 and n2154 n4788 ; n4789
g4726 and n1306_not n4789 ; n4790
g4727 and n397_not n4790 ; n4791
g4728 and n189_not n4791 ; n4792
g4729 and n233_not n4792 ; n4793
g4730 and n161_not n4793 ; n4794
g4731 nor n205 n275 ; n4795
g4732 and n961_not n4795 ; n4796
g4733 and n249_not n4796 ; n4797
g4734 and n1761 n4367 ; n4798
g4735 and n715_not n4798 ; n4799
g4736 and n4797 n4799 ; n4800
g4737 and n297 n4800 ; n4801
g4738 and n439 n4801 ; n4802
g4739 and n4794 n4802 ; n4803
g4740 and n4786 n4803 ; n4804
g4741 and n933 n4804 ; n4805
g4742 and n2219 n4805 ; n4806
g4743 and n341 n4806 ; n4807
g4744 and n469_not n4807 ; n4808
g4745 and n276_not n4808 ; n4809
g4746 and n557_not n4809 ; n4810
g4747 and n602_not n4810 ; n4811
g4748 and n150_not n4811 ; n4812
g4749 and n416_not n4812 ; n4813
g4750 and n191_not n4813 ; n4814
g4751 and n791_not n4814 ; n4815
g4752 nor n164 n558 ; n4816
g4753 and n537_not n4816 ; n4817
g4754 and n200_not n4817 ; n4818
g4755 and n672_not n4818 ; n4819
g4756 and n2584 n2721 ; n4820
g4757 and n4819 n4820 ; n4821
g4758 and n1726 n4821 ; n4822
g4759 and n570 n4822 ; n4823
g4760 and n1011_not n4823 ; n4824
g4761 and n290_not n4824 ; n4825
g4762 and n246_not n4825 ; n4826
g4763 and n393_not n4826 ; n4827
g4764 nor n496 n884 ; n4828
g4765 and n1973 n4828 ; n4829
g4766 and n4827 n4829 ; n4830
g4767 and n4815 n4830 ; n4831
g4768 and n1928 n4831 ; n4832
g4769 and n4785 n4832 ; n4833
g4770 and n4767 n4833 ; n4834
g4771 and n1576 n4834 ; n4835
g4772 and n423 n4835 ; n4836
g4773 and n2467 n4836 ; n4837
g4774 and n667_not n4837 ; n4838
g4775 and n91_not n4838 ; n4839
g4776 and n243_not n4839 ; n4840
g4777 and n536_not n4840 ; n4841
g4778 and n283_not n4841 ; n4842
g4779 and n237_not n4842 ; n4843
g4780 and n271_not n4843 ; n4844
g4781 and n4351 n4844_not ; n4845
g4782 and n4351_not n4844 ; n4846
g4783 and n2896 n2898_not ; n4847
g4784 nor n2899 n4847 ; n4848
g4785 and n75 n4848 ; n4849
g4786 and n1235_not n3020 ; n4850
g4787 and n1472_not n3023 ; n4851
g4788 and n1364_not n3028 ; n4852
g4789 nor n4851 n4852 ; n4853
g4790 and n4850_not n4853 ; n4854
g4791 and n4849_not n4854 ; n4855
g4792 nor n4845 n4855 ; n4856
g4793 and n4846_not n4856 ; n4857
g4794 nor n4845 n4857 ; n4858
g4795 nor n4761 n4858 ; n4859
g4796 and n2900 n2902_not ; n4860
g4797 nor n2903 n4860 ; n4861
g4798 and n75 n4861 ; n4862
g4799 and n1178_not n3020 ; n4863
g4800 and n1364_not n3023 ; n4864
g4801 and n1235_not n3028 ; n4865
g4802 nor n4864 n4865 ; n4866
g4803 and n4863_not n4866 ; n4867
g4804 and n4862_not n4867 ; n4868
g4805 and n4761 n4858 ; n4869
g4806 nor n4859 n4869 ; n4870
g4807 and n4868_not n4870 ; n4871
g4808 nor n4859 n4871 ; n4872
g4809 nor n4758 n4872 ; n4873
g4810 and n4758 n4872 ; n4874
g4811 nor n4873 n4874 ; n4875
g4812 and n710_not n3457 ; n4876
g4813 and n958_not n3542 ; n4877
g4814 and n867_not n3606 ; n4878
g4815 nor n4877 n4878 ; n4879
g4816 and n4876_not n4879 ; n4880
g4817 and n3368_not n4880 ; n4881
g4818 and n4179_not n4880 ; n4882
g4819 nor n4881 n4882 ; n4883
g4820 and a[29] n4883_not ; n4884
g4821 and a[29]_not n4883 ; n4885
g4822 nor n4884 n4885 ; n4886
g4823 and n4875 n4886_not ; n4887
g4824 nor n4873 n4887 ; n4888
g4825 nor n4755 n4888 ; n4889
g4826 and n4755 n4888 ; n4890
g4827 nor n4889 n4890 ; n4891
g4828 and n3539_not n3884 ; n4892
g4829 and n392_not n3967 ; n4893
g4830 and n3012_not n4046 ; n4894
g4831 nor n4893 n4894 ; n4895
g4832 and n4892_not n4895 ; n4896
g4833 and n3715 n4050 ; n4897
g4834 and n4896 n4897_not ; n4898
g4835 and a[26] n4898_not ; n4899
g4836 and a[26] n4899_not ; n4900
g4837 nor n4898 n4899 ; n4901
g4838 nor n4900 n4901 ; n4902
g4839 and n4891 n4902_not ; n4903
g4840 nor n4889 n4903 ; n4904
g4841 and n4740 n4751 ; n4905
g4842 nor n4752 n4905 ; n4906
g4843 and n4904_not n4906 ; n4907
g4844 nor n4752 n4907 ; n4908
g4845 nor n4737 n4908 ; n4909
g4846 and n4737 n4908 ; n4910
g4847 nor n4909 n4910 ; n4911
g4848 and n4045_not n4694 ; n4912
g4849 and n3805_not n4533 ; n4913
g4850 and n3964_not n4604 ; n4914
g4851 nor n4913 n4914 ; n4915
g4852 and n4912_not n4915 ; n4916
g4853 and n4477 n4536 ; n4917
g4854 and n4916 n4917_not ; n4918
g4855 and a[23] n4918_not ; n4919
g4856 and a[23] n4919_not ; n4920
g4857 nor n4918 n4919 ; n4921
g4858 nor n4920 n4921 ; n4922
g4859 and n4911 n4922_not ; n4923
g4860 nor n4909 n4923 ; n4924
g4861 and a[18]_not a[19] ; n4925
g4862 and a[18] a[19]_not ; n4926
g4863 nor n4925 n4926 ; n4927
g4864 and a[19] a[20]_not ; n4928
g4865 and a[19]_not a[20] ; n4929
g4866 nor n4928 n4929 ; n4930
g4867 and a[17] a[18]_not ; n4931
g4868 and a[17]_not a[18] ; n4932
g4869 nor n4931 n4932 ; n4933
g4870 and n4930_not n4933 ; n4934
g4871 and n4927 n4934 ; n4935
g4872 and n4515_not n4935 ; n4936
g4873 nor n4522 n4936 ; n4937
g4874 nor n4930 n4933 ; n4938
g4875 nor n4936 n4938 ; n4939
g4876 nor n4937 n4939 ; n4940
g4877 and a[20] n4940_not ; n4941
g4878 and a[20]_not n4940 ; n4942
g4879 nor n4941 n4942 ; n4943
g4880 nor n4924 n4943 ; n4944
g4881 and n4693 n4706_not ; n4945
g4882 nor n4705 n4706 ; n4946
g4883 nor n4945 n4946 ; n4947
g4884 and n4924 n4943 ; n4948
g4885 nor n4944 n4948 ; n4949
g4886 and n4947_not n4949 ; n4950
g4887 nor n4944 n4950 ; n4951
g4888 nor n4734 n4951 ; n4952
g4889 and n4734 n4951 ; n4953
g4890 nor n4952 n4953 ; n4954
g4891 nor n4947 n4950 ; n4955
g4892 and n4949 n4950_not ; n4956
g4893 nor n4955 n4956 ; n4957
g4894 and n4911 n4923_not ; n4958
g4895 nor n4922 n4923 ; n4959
g4896 nor n4958 n4959 ; n4960
g4897 and n3964_not n4694 ; n4961
g4898 and n3456_not n4533 ; n4962
g4899 and n3805_not n4604 ; n4963
g4900 nor n4962 n4963 ; n4964
g4901 and n4961_not n4964 ; n4965
g4902 and n4536 n4558 ; n4966
g4903 and n4965 n4966_not ; n4967
g4904 and a[23] n4967_not ; n4968
g4905 nor n4967 n4968 ; n4969
g4906 and a[23] n4968_not ; n4970
g4907 nor n4969 n4970 ; n4971
g4908 and n4904 n4906_not ; n4972
g4909 nor n4907 n4972 ; n4973
g4910 and n4971_not n4973 ; n4974
g4911 nor n4971 n4974 ; n4975
g4912 and n4973 n4974_not ; n4976
g4913 nor n4975 n4976 ; n4977
g4914 and n4891 n4903_not ; n4978
g4915 nor n4902 n4903 ; n4979
g4916 nor n4978 n4979 ; n4980
g4917 and n867_not n3457 ; n4981
g4918 and n1060_not n3542 ; n4982
g4919 and n958_not n3606 ; n4983
g4920 nor n4982 n4983 ; n4984
g4921 and n4981_not n4984 ; n4985
g4922 and n3368 n4204 ; n4986
g4923 and n4985 n4986_not ; n4987
g4924 and a[29] n4987_not ; n4988
g4925 nor n4987 n4988 ; n4989
g4926 and a[29] n4988_not ; n4990
g4927 nor n4989 n4990 ; n4991
g4928 nor n4868 n4871 ; n4992
g4929 and n4870 n4871_not ; n4993
g4930 nor n4992 n4993 ; n4994
g4931 nor n4991 n4994 ; n4995
g4932 nor n4991 n4995 ; n4996
g4933 nor n4994 n4995 ; n4997
g4934 nor n4996 n4997 ; n4998
g4935 nor n4855 n4857 ; n4999
g4936 and n4846_not n4858 ; n5000
g4937 nor n4999 n5000 ; n5001
g4938 nor n394 n1062 ; n5002
g4939 and n2546 n5002 ; n5003
g4940 and n4357 n5003 ; n5004
g4941 and n3438 n5004 ; n5005
g4942 and n3886 n5005 ; n5006
g4943 and n421 n5006 ; n5007
g4944 and n1237 n5007 ; n5008
g4945 and n305_not n5008 ; n5009
g4946 and n302_not n5009 ; n5010
g4947 and n589_not n5010 ; n5011
g4948 and n468_not n5011 ; n5012
g4949 and n883_not n5012 ; n5013
g4950 and n364_not n1709 ; n5014
g4951 and n121_not n5014 ; n5015
g4952 and n422_not n5015 ; n5016
g4953 and n130_not n5016 ; n5017
g4954 and n325_not n5017 ; n5018
g4955 and n158_not n5018 ; n5019
g4956 nor n170 n825 ; n5020
g4957 and n519_not n5020 ; n5021
g4958 and n1331 n1861 ; n5022
g4959 and n5021 n5022 ; n5023
g4960 and n811 n5023 ; n5024
g4961 and n5019 n5024 ; n5025
g4962 and n3163 n5025 ; n5026
g4963 and n154_not n5026 ; n5027
g4964 and n135_not n5027 ; n5028
g4965 and n1102_not n5028 ; n5029
g4966 and n402_not n5029 ; n5030
g4967 and n290_not n5030 ; n5031
g4968 and n374_not n5031 ; n5032
g4969 and n689_not n5032 ; n5033
g4970 and n231_not n5033 ; n5034
g4971 nor n304 n513 ; n5035
g4972 and n251_not n5035 ; n5036
g4973 nor n339 n398 ; n5037
g4974 and n283_not n5037 ; n5038
g4975 and n979 n2406 ; n5039
g4976 and n1072_not n5039 ; n5040
g4977 and n812 n5040 ; n5041
g4978 and n5038 n5041 ; n5042
g4979 and n5036 n5042 ; n5043
g4980 and n4216 n5043 ; n5044
g4981 and n4332 n5044 ; n5045
g4982 and n1610 n5045 ; n5046
g4983 and n2979 n5046 ; n5047
g4984 and n5034 n5047 ; n5048
g4985 and n5013 n5048 ; n5049
g4986 and n752_not n5049 ; n5050
g4987 and n1101_not n5050 ; n5051
g4988 and n201_not n5051 ; n5052
g4989 and n562_not n5052 ; n5053
g4990 nor n511 n746 ; n5054
g4991 and n283_not n5054 ; n5055
g4992 and n562_not n5055 ; n5056
g4993 and n2608 n3043 ; n5057
g4994 and n5056 n5057 ; n5058
g4995 and n621 n5058 ; n5059
g4996 and n896 n5059 ; n5060
g4997 and n403_not n5060 ; n5061
g4998 and n416_not n5061 ; n5062
g4999 and n144_not n5062 ; n5063
g5000 nor n225 n716 ; n5064
g5001 nor n280 n847 ; n5065
g5002 and n402_not n5065 ; n5066
g5003 and n5064 n5066 ; n5067
g5004 and n1249 n5067 ; n5068
g5005 and n5063 n5068 ; n5069
g5006 and n664 n5069 ; n5070
g5007 and n1668 n5070 ; n5071
g5008 and n1667 n5071 ; n5072
g5009 and n356 n5072 ; n5073
g5010 and n1040 n5073 ; n5074
g5011 and n617_not n5074 ; n5075
g5012 and n169_not n5075 ; n5076
g5013 and n329_not n5076 ; n5077
g5014 and n335_not n5077 ; n5078
g5015 and n803_not n5078 ; n5079
g5016 and n1203_not n5079 ; n5080
g5017 and n375_not n5080 ; n5081
g5018 and n158_not n5081 ; n5082
g5019 nor n298 n825 ; n5083
g5020 and n130_not n5083 ; n5084
g5021 and n493_not n5084 ; n5085
g5022 and n1012 n1107 ; n5086
g5023 and n3663 n5086 ; n5087
g5024 and n789 n5087 ; n5088
g5025 and n811 n5088 ; n5089
g5026 and n3094 n5089 ; n5090
g5027 and n5085 n5090 ; n5091
g5028 and n2170 n5091 ; n5092
g5029 and n5082 n5092 ; n5093
g5030 and n5013 n5093 ; n5094
g5031 and n508 n5094 ; n5095
g5032 and n116 n5095 ; n5096
g5033 and n418 n5096 ; n5097
g5034 and n278_not n5097 ; n5098
g5035 and n506_not n5098 ; n5099
g5036 and n594_not n5099 ; n5100
g5037 and n286_not n5100 ; n5101
g5038 and n424_not n5101 ; n5102
g5039 and n932_not n5102 ; n5103
g5040 and n340_not n5103 ; n5104
g5041 and n337_not n5104 ; n5105
g5042 and n429_not n5105 ; n5106
g5043 nor n5053 n5106 ; n5107
g5044 and n5053 n5106 ; n5108
g5045 nor n5107 n5108 ; n5109
g5046 and a[11]_not n5109 ; n5110
g5047 nor n5107 n5110 ; n5111
g5048 and n4351 n5111_not ; n5112
g5049 and n2892 n2894_not ; n5113
g5050 nor n2895 n5113 ; n5114
g5051 and n75 n5114 ; n5115
g5052 and n1364_not n3020 ; n5116
g5053 and n1572_not n3023 ; n5117
g5054 and n1472_not n3028 ; n5118
g5055 nor n5117 n5118 ; n5119
g5056 and n5116_not n5119 ; n5120
g5057 and n5115_not n5120 ; n5121
g5058 and n4351_not n5111 ; n5122
g5059 nor n5112 n5122 ; n5123
g5060 and n5121_not n5123 ; n5124
g5061 nor n5112 n5124 ; n5125
g5062 nor n5001 n5125 ; n5126
g5063 and n5001 n5125 ; n5127
g5064 nor n5126 n5127 ; n5128
g5065 nor n5121 n5124 ; n5129
g5066 and n5123 n5124_not ; n5130
g5067 nor n5129 n5130 ; n5131
g5068 nor a[11] n5110 ; n5132
g5069 and n5108_not n5111 ; n5133
g5070 nor n5132 n5133 ; n5134
g5071 and n1472_not n3020 ; n5135
g5072 and n1572_not n3028 ; n5136
g5073 and n1665_not n3023 ; n5137
g5074 and n2888 n2890_not ; n5138
g5075 nor n2891 n5138 ; n5139
g5076 and n75 n5139 ; n5140
g5077 nor n5137 n5140 ; n5141
g5078 and n5136_not n5141 ; n5142
g5079 and n5135_not n5142 ; n5143
g5080 nor n5134 n5143 ; n5144
g5081 and n115_not n1183 ; n5145
g5082 and n107_not n5145 ; n5146
g5083 and n205_not n5146 ; n5147
g5084 and n564_not n5147 ; n5148
g5085 and n428_not n1523 ; n5149
g5086 and n270_not n5149 ; n5150
g5087 and n168_not n1330 ; n5151
g5088 and n252_not n5151 ; n5152
g5089 and n5150 n5152 ; n5153
g5090 and n921 n5153 ; n5154
g5091 and n5148 n5154 ; n5155
g5092 and n1635 n5155 ; n5156
g5093 and n3651 n5156 ; n5157
g5094 and n1585 n5157 ; n5158
g5095 and n1915 n5158 ; n5159
g5096 and n2484 n5159 ; n5160
g5097 and n770 n5160 ; n5161
g5098 and n1072_not n5161 ; n5162
g5099 and n514_not n5162 ; n5163
g5100 and n290_not n5163 ; n5164
g5101 and n825_not n5164 ; n5165
g5102 and n673_not n5165 ; n5166
g5103 and n537_not n5166 ; n5167
g5104 and n325_not n5167 ; n5168
g5105 and n5053 n5168_not ; n5169
g5106 and n5053_not n5168 ; n5170
g5107 nor n713 n1101 ; n5171
g5108 and n328_not n1128 ; n5172
g5109 and n287_not n5172 ; n5173
g5110 and n2278 n5173 ; n5174
g5111 and n897 n5174 ; n5175
g5112 and n4356 n5175 ; n5176
g5113 and n512 n5176 ; n5177
g5114 and n654 n5177 ; n5178
g5115 and n356 n5178 ; n5179
g5116 and n3163 n5179 ; n5180
g5117 and n571_not n5180 ; n5181
g5118 and n396_not n5181 ; n5182
g5119 and n226_not n5182 ; n5183
g5120 and n639_not n5183 ; n5184
g5121 and n980_not n5184 ; n5185
g5122 and n200_not n5185 ; n5186
g5123 and n272_not n5186 ; n5187
g5124 and n295_not n5187 ; n5188
g5125 nor n169 n462 ; n5189
g5126 and n286_not n5189 ; n5190
g5127 and n2423 n5190 ; n5191
g5128 and n1011_not n5191 ; n5192
g5129 and n327_not n5192 ; n5193
g5130 and n326_not n2240 ; n5194
g5131 and n673_not n5194 ; n5195
g5132 and n961_not n5195 ; n5196
g5133 and n603_not n5196 ; n5197
g5134 and n366_not n5197 ; n5198
g5135 and n886_not n5198 ; n5199
g5136 nor n175 n453 ; n5200
g5137 and n449_not n5200 ; n5201
g5138 and n236_not n5201 ; n5202
g5139 and n746_not n5202 ; n5203
g5140 and n229_not n5203 ; n5204
g5141 and n150_not n5204 ; n5205
g5142 and n438_not n5205 ; n5206
g5143 and n243_not n5206 ; n5207
g5144 and n372_not n5207 ; n5208
g5145 and n655_not n5208 ; n5209
g5146 and n2297 n4313 ; n5210
g5147 and n593 n5210 ; n5211
g5148 and n1024 n5211 ; n5212
g5149 and n1131 n5212 ; n5213
g5150 and n5209 n5213 ; n5214
g5151 and n5199 n5214 ; n5215
g5152 and n111_not n5215 ; n5216
g5153 and n620_not n5216 ; n5217
g5154 and n417_not n5217 ; n5218
g5155 and n167_not n5218 ; n5219
g5156 and n173_not n5219 ; n5220
g5157 and n623_not n5220 ; n5221
g5158 and n1104_not n5221 ; n5222
g5159 and n474_not n5222 ; n5223
g5160 and n569_not n5223 ; n5224
g5161 and n1085 n2752 ; n5225
g5162 and n1155 n5225 ; n5226
g5163 and n1367 n5226 ; n5227
g5164 and n330_not n5227 ; n5228
g5165 and n298_not n5228 ; n5229
g5166 and n130_not n5229 ; n5230
g5167 and n712_not n5230 ; n5231
g5168 and n532_not n5231 ; n5232
g5169 and n81_not n5232 ; n5233
g5170 and n1732 n2133 ; n5234
g5171 and n232_not n5234 ; n5235
g5172 and n255_not n5235 ; n5236
g5173 and n299_not n5236 ; n5237
g5174 and n527_not n5237 ; n5238
g5175 and n158_not n5238 ; n5239
g5176 and n636 n5066 ; n5240
g5177 and n1819 n5240 ; n5241
g5178 and n5239 n5241 ; n5242
g5179 and n5233 n5242 ; n5243
g5180 and n5224 n5243 ; n5244
g5181 and n5193 n5244 ; n5245
g5182 and n5188 n5245 ; n5246
g5183 and n602_not n5246 ; n5247
g5184 and n5171 n5247 ; n5248
g5185 and n339_not n5248 ; n5249
g5186 and n145_not n5249 ; n5250
g5187 and n201_not n5250 ; n5251
g5188 and n666_not n5251 ; n5252
g5189 and n337_not n5252 ; n5253
g5190 and n429_not n5253 ; n5254
g5191 and n2424 n3040 ; n5255
g5192 and n2021 n5255 ; n5256
g5193 and n364_not n5256 ; n5257
g5194 and n355_not n5257 ; n5258
g5195 and n152_not n5258 ; n5259
g5196 and n115_not n5259 ; n5260
g5197 and n884_not n5260 ; n5261
g5198 and n191_not n5261 ; n5262
g5199 and n1104_not n5262 ; n5263
g5200 and n449_not n5263 ; n5264
g5201 and n634 n937 ; n5265
g5202 and n275_not n5265 ; n5266
g5203 and n240_not n5266 ; n5267
g5204 and n188_not n5267 ; n5268
g5205 and n249_not n5268 ; n5269
g5206 and n202 n513_not ; n5270
g5207 and n428_not n5270 ; n5271
g5208 and n3268 n5271 ; n5272
g5209 and n593 n5272 ; n5273
g5210 and n5269 n5273 ; n5274
g5211 and n5264 n5274 ; n5275
g5212 and n873 n5275 ; n5276
g5213 and n872 n5276 ; n5277
g5214 and n2346 n5277 ; n5278
g5215 and n1575 n5278 ; n5279
g5216 and n621 n5279 ; n5280
g5217 and n1306_not n5280 ; n5281
g5218 and n284_not n5281 ; n5282
g5219 and n425_not n5282 ; n5283
g5220 and n306_not n5283 ; n5284
g5221 and n157_not n5284 ; n5285
g5222 and n519_not n5285 ; n5286
g5223 and n1604 n2508 ; n5287
g5224 and n1103 n5287 ; n5288
g5225 and n665 n5288 ; n5289
g5226 and n123_not n5289 ; n5290
g5227 and n107_not n5290 ; n5291
g5228 and n305_not n5291 ; n5292
g5229 and n287_not n5292 ; n5293
g5230 and n490_not n5293 ; n5294
g5231 and n375_not n5294 ; n5295
g5232 and n277_not n5295 ; n5296
g5233 and n154_not n1248 ; n5297
g5234 and n667_not n5297 ; n5298
g5235 and n278_not n5298 ; n5299
g5236 and n589_not n5299 ; n5300
g5237 and n712_not n5300 ; n5301
g5238 and n338_not n5301 ; n5302
g5239 and n564_not n5302 ; n5303
g5240 and n358_not n5303 ; n5304
g5241 and n2627 n3264 ; n5305
g5242 and n3312 n5305 ; n5306
g5243 and n5304 n5306 ; n5307
g5244 and n1577 n5307 ; n5308
g5245 and n247 n5308 ; n5309
g5246 and n5296 n5309 ; n5310
g5247 and n1254 n5310 ; n5311
g5248 and n615 n5311 ; n5312
g5249 and n5286 n5312 ; n5313
g5250 and n100 n5313 ; n5314
g5251 and n335_not n5314 ; n5315
g5252 and n402_not n5315 ; n5316
g5253 and n825_not n5316 ; n5317
g5254 and n296_not n5317 ; n5318
g5255 and n192_not n5318 ; n5319
g5256 and n429_not n5319 ; n5320
g5257 nor n5254 n5320 ; n5321
g5258 and n5254 n5320 ; n5322
g5259 nor n5321 n5322 ; n5323
g5260 and a[8]_not n5323 ; n5324
g5261 nor n5321 n5324 ; n5325
g5262 and n5053 n5325_not ; n5326
g5263 and n2880 n2882_not ; n5327
g5264 nor n2883 n5327 ; n5328
g5265 and n75 n5328 ; n5329
g5266 and n1665_not n3020 ; n5330
g5267 and n1877_not n3023 ; n5331
g5268 and n1779_not n3028 ; n5332
g5269 nor n5331 n5332 ; n5333
g5270 and n5330_not n5333 ; n5334
g5271 and n5329_not n5334 ; n5335
g5272 and n5053_not n5325 ; n5336
g5273 nor n5326 n5336 ; n5337
g5274 and n5335_not n5337 ; n5338
g5275 nor n5326 n5338 ; n5339
g5276 nor n5169 n5339 ; n5340
g5277 and n5170_not n5340 ; n5341
g5278 nor n5169 n5341 ; n5342
g5279 and n5134 n5143 ; n5343
g5280 nor n5144 n5343 ; n5344
g5281 and n5342_not n5344 ; n5345
g5282 nor n5144 n5345 ; n5346
g5283 nor n5131 n5346 ; n5347
g5284 and n5131 n5346 ; n5348
g5285 nor n5347 n5348 ; n5349
g5286 and n1060_not n3457 ; n5350
g5287 and n1235_not n3542 ; n5351
g5288 and n1178_not n3606 ; n5352
g5289 nor n5351 n5352 ; n5353
g5290 and n5350_not n5353 ; n5354
g5291 and n3368_not n5354 ; n5355
g5292 and n4429_not n5354 ; n5356
g5293 nor n5355 n5356 ; n5357
g5294 and a[29] n5357_not ; n5358
g5295 and a[29]_not n5357 ; n5359
g5296 nor n5358 n5359 ; n5360
g5297 and n5349 n5360_not ; n5361
g5298 nor n5347 n5361 ; n5362
g5299 and n5128 n5362_not ; n5363
g5300 nor n5126 n5363 ; n5364
g5301 nor n4998 n5364 ; n5365
g5302 nor n4995 n5365 ; n5366
g5303 and n4875_not n4886 ; n5367
g5304 nor n4887 n5367 ; n5368
g5305 and n5366_not n5368 ; n5369
g5306 and n5366 n5368_not ; n5370
g5307 nor n5369 n5370 ; n5371
g5308 and n3012_not n3884 ; n5372
g5309 and n587_not n3967 ; n5373
g5310 and n392_not n4046 ; n5374
g5311 nor n5373 n5374 ; n5375
g5312 and n5372_not n5375 ; n5376
g5313 and n3018 n4050 ; n5377
g5314 and n5376 n5377_not ; n5378
g5315 and a[26] n5378_not ; n5379
g5316 and a[26] n5379_not ; n5380
g5317 nor n5378 n5379 ; n5381
g5318 nor n5380 n5381 ; n5382
g5319 and n5371 n5382_not ; n5383
g5320 nor n5369 n5383 ; n5384
g5321 nor n4980 n5384 ; n5385
g5322 and n4980 n5384 ; n5386
g5323 nor n5385 n5386 ; n5387
g5324 and n3805_not n4694 ; n5388
g5325 and n3605_not n4533 ; n5389
g5326 and n3456_not n4604 ; n5390
g5327 nor n5389 n5390 ; n5391
g5328 and n5388_not n5391 ; n5392
g5329 and n3818 n4536 ; n5393
g5330 and n5392 n5393_not ; n5394
g5331 and a[23] n5394_not ; n5395
g5332 and a[23] n5395_not ; n5396
g5333 nor n5394 n5395 ; n5397
g5334 nor n5396 n5397 ; n5398
g5335 and n5387 n5398_not ; n5399
g5336 nor n5385 n5399 ; n5400
g5337 nor n4977 n5400 ; n5401
g5338 nor n4974 n5401 ; n5402
g5339 nor n4960 n5402 ; n5403
g5340 and n4960 n5402 ; n5404
g5341 nor n5403 n5404 ; n5405
g5342 and n3877_not n4935 ; n5406
g5343 and n4927_not n4933 ; n5407
g5344 and n4515_not n5407 ; n5408
g5345 nor n5406 n5408 ; n5409
g5346 and n4609 n4938 ; n5410
g5347 and n5409 n5410_not ; n5411
g5348 and a[20] n5411_not ; n5412
g5349 and a[20] n5412_not ; n5413
g5350 nor n5411 n5412 ; n5414
g5351 nor n5413 n5414 ; n5415
g5352 and n5405 n5415_not ; n5416
g5353 nor n5403 n5416 ; n5417
g5354 nor n4957 n5417 ; n5418
g5355 and n4957 n5417 ; n5419
g5356 nor n5418 n5419 ; n5420
g5357 and n5405 n5416_not ; n5421
g5358 nor n5415 n5416 ; n5422
g5359 nor n5421 n5422 ; n5423
g5360 and n5387 n5399_not ; n5424
g5361 nor n5398 n5399 ; n5425
g5362 nor n5424 n5425 ; n5426
g5363 and n5371 n5383_not ; n5427
g5364 nor n5382 n5383 ; n5428
g5365 nor n5427 n5428 ; n5429
g5366 and n4998 n5364 ; n5430
g5367 nor n5365 n5430 ; n5431
g5368 and n392_not n3884 ; n5432
g5369 and n710_not n3967 ; n5433
g5370 and n587_not n4046 ; n5434
g5371 nor n5433 n5434 ; n5435
g5372 and n5432_not n5435 ; n5436
g5373 and n4050_not n5436 ; n5437
g5374 and n3347_not n5436 ; n5438
g5375 nor n5437 n5438 ; n5439
g5376 and a[26] n5439_not ; n5440
g5377 and a[26]_not n5439 ; n5441
g5378 nor n5440 n5441 ; n5442
g5379 and n5431 n5442_not ; n5443
g5380 and n587_not n3884 ; n5444
g5381 and n867_not n3967 ; n5445
g5382 and n710_not n4046 ; n5446
g5383 nor n5445 n5446 ; n5447
g5384 and n5444_not n5447 ; n5448
g5385 and n3331 n4050 ; n5449
g5386 and n5448 n5449_not ; n5450
g5387 and a[26] n5450_not ; n5451
g5388 and a[26] n5451_not ; n5452
g5389 nor n5450 n5451 ; n5453
g5390 nor n5452 n5453 ; n5454
g5391 and n5128_not n5362 ; n5455
g5392 nor n5363 n5455 ; n5456
g5393 and n958_not n3457 ; n5457
g5394 and n1178_not n3542 ; n5458
g5395 and n1060_not n3606 ; n5459
g5396 nor n5458 n5459 ; n5460
g5397 and n5457_not n5460 ; n5461
g5398 and n3368_not n5461 ; n5462
g5399 and n4633_not n5461 ; n5463
g5400 nor n5462 n5463 ; n5464
g5401 and a[29] n5464_not ; n5465
g5402 and a[29]_not n5464 ; n5466
g5403 nor n5465 n5466 ; n5467
g5404 and n5456 n5467_not ; n5468
g5405 and n5456_not n5467 ; n5469
g5406 nor n5468 n5469 ; n5470
g5407 and n5454_not n5470 ; n5471
g5408 nor n5468 n5471 ; n5472
g5409 and n5431_not n5442 ; n5473
g5410 nor n5443 n5473 ; n5474
g5411 and n5472_not n5474 ; n5475
g5412 nor n5443 n5475 ; n5476
g5413 nor n5429 n5476 ; n5477
g5414 and n5429 n5476 ; n5478
g5415 nor n5477 n5478 ; n5479
g5416 and n3456_not n4694 ; n5480
g5417 and n3539_not n4533 ; n5481
g5418 and n3605_not n4604 ; n5482
g5419 nor n5481 n5482 ; n5483
g5420 and n5480_not n5483 ; n5484
g5421 and n3627 n4536 ; n5485
g5422 and n5484 n5485_not ; n5486
g5423 and a[23] n5486_not ; n5487
g5424 and a[23] n5487_not ; n5488
g5425 nor n5486 n5487 ; n5489
g5426 nor n5488 n5489 ; n5490
g5427 and n5479 n5490_not ; n5491
g5428 nor n5477 n5491 ; n5492
g5429 nor n5426 n5492 ; n5493
g5430 and n5426 n5492 ; n5494
g5431 nor n5493 n5494 ; n5495
g5432 and n4930 n4933_not ; n5496
g5433 and n3877_not n5496 ; n5497
g5434 and n3964_not n4935 ; n5498
g5435 and n4045_not n5407 ; n5499
g5436 nor n5498 n5499 ; n5500
g5437 and n5497_not n5500 ; n5501
g5438 and n4067 n4938 ; n5502
g5439 and n5501 n5502_not ; n5503
g5440 and a[20] n5503_not ; n5504
g5441 and a[20] n5504_not ; n5505
g5442 nor n5503 n5504 ; n5506
g5443 nor n5505 n5506 ; n5507
g5444 and n5495 n5507_not ; n5508
g5445 nor n5493 n5508 ; n5509
g5446 and n4515_not n5496 ; n5510
g5447 and n4045_not n4935 ; n5511
g5448 and n3877_not n5407 ; n5512
g5449 nor n5511 n5512 ; n5513
g5450 and n5510_not n5513 ; n5514
g5451 and n4938_not n5514 ; n5515
g5452 and n4715_not n5514 ; n5516
g5453 nor n5515 n5516 ; n5517
g5454 and a[20] n5517_not ; n5518
g5455 and a[20]_not n5517 ; n5519
g5456 nor n5518 n5519 ; n5520
g5457 nor n5509 n5520 ; n5521
g5458 and n4977 n5400 ; n5522
g5459 nor n5401 n5522 ; n5523
g5460 and n5509 n5520 ; n5524
g5461 nor n5521 n5524 ; n5525
g5462 and n5523 n5525 ; n5526
g5463 nor n5521 n5526 ; n5527
g5464 nor n5423 n5527 ; n5528
g5465 and n5423 n5527 ; n5529
g5466 nor n5528 n5529 ; n5530
g5467 and n5479 n5491_not ; n5531
g5468 nor n5490 n5491 ; n5532
g5469 nor n5531 n5532 ; n5533
g5470 and n3605_not n4694 ; n5534
g5471 and n3012_not n4533 ; n5535
g5472 and n3539_not n4604 ; n5536
g5473 nor n5535 n5536 ; n5537
g5474 and n5534_not n5537 ; n5538
g5475 and n4084 n4536 ; n5539
g5476 and n5538 n5539_not ; n5540
g5477 and a[23] n5540_not ; n5541
g5478 nor n5540 n5541 ; n5542
g5479 and a[23] n5541_not ; n5543
g5480 nor n5542 n5543 ; n5544
g5481 and n5472 n5474_not ; n5545
g5482 nor n5475 n5545 ; n5546
g5483 and n5544_not n5546 ; n5547
g5484 nor n5544 n5547 ; n5548
g5485 and n5546 n5547_not ; n5549
g5486 nor n5548 n5549 ; n5550
g5487 and n5470 n5471_not ; n5551
g5488 nor n5454 n5471 ; n5552
g5489 nor n5551 n5552 ; n5553
g5490 nor n5339 n5341 ; n5554
g5491 and n5170_not n5342 ; n5555
g5492 nor n5554 n5555 ; n5556
g5493 and n1572_not n3020 ; n5557
g5494 and n1665_not n3028 ; n5558
g5495 and n1779_not n3023 ; n5559
g5496 and n2884 n2886_not ; n5560
g5497 nor n2887 n5560 ; n5561
g5498 and n75 n5561 ; n5562
g5499 nor n5559 n5562 ; n5563
g5500 and n5558_not n5563 ; n5564
g5501 and n5557_not n5564 ; n5565
g5502 nor n5556 n5565 ; n5566
g5503 and n1235_not n3457 ; n5567
g5504 and n1472_not n3542 ; n5568
g5505 and n1364_not n3606 ; n5569
g5506 nor n5568 n5569 ; n5570
g5507 and n5567_not n5570 ; n5571
g5508 and n3368 n4848 ; n5572
g5509 and n5571 n5572_not ; n5573
g5510 and a[29] n5573_not ; n5574
g5511 nor n5573 n5574 ; n5575
g5512 and a[29] n5574_not ; n5576
g5513 nor n5575 n5576 ; n5577
g5514 nor n5556 n5566 ; n5578
g5515 nor n5565 n5566 ; n5579
g5516 nor n5578 n5579 ; n5580
g5517 nor n5577 n5580 ; n5581
g5518 nor n5566 n5581 ; n5582
g5519 and n5342 n5344_not ; n5583
g5520 nor n5345 n5583 ; n5584
g5521 and n5582_not n5584 ; n5585
g5522 and n1178_not n3457 ; n5586
g5523 and n1364_not n3542 ; n5587
g5524 and n1235_not n3606 ; n5588
g5525 nor n5587 n5588 ; n5589
g5526 and n5586_not n5589 ; n5590
g5527 and n3368 n4861 ; n5591
g5528 and n5590 n5591_not ; n5592
g5529 and a[29] n5592_not ; n5593
g5530 and a[29] n5593_not ; n5594
g5531 nor n5592 n5593 ; n5595
g5532 nor n5594 n5595 ; n5596
g5533 and n5582 n5584_not ; n5597
g5534 nor n5585 n5597 ; n5598
g5535 and n5596_not n5598 ; n5599
g5536 nor n5585 n5599 ; n5600
g5537 and n5349_not n5360 ; n5601
g5538 nor n5361 n5601 ; n5602
g5539 and n5600_not n5602 ; n5603
g5540 and n5600 n5602_not ; n5604
g5541 nor n5603 n5604 ; n5605
g5542 and n710_not n3884 ; n5606
g5543 and n958_not n3967 ; n5607
g5544 and n867_not n4046 ; n5608
g5545 nor n5607 n5608 ; n5609
g5546 and n5606_not n5609 ; n5610
g5547 and n4050 n4179 ; n5611
g5548 and n5610 n5611_not ; n5612
g5549 and a[26] n5612_not ; n5613
g5550 and a[26] n5613_not ; n5614
g5551 nor n5612 n5613 ; n5615
g5552 nor n5614 n5615 ; n5616
g5553 and n5605 n5616_not ; n5617
g5554 nor n5603 n5617 ; n5618
g5555 nor n5553 n5618 ; n5619
g5556 and n5553 n5618 ; n5620
g5557 nor n5619 n5620 ; n5621
g5558 and n3539_not n4694 ; n5622
g5559 and n392_not n4533 ; n5623
g5560 and n3012_not n4604 ; n5624
g5561 nor n5623 n5624 ; n5625
g5562 and n5622_not n5625 ; n5626
g5563 and n3715 n4536 ; n5627
g5564 and n5626 n5627_not ; n5628
g5565 and a[23] n5628_not ; n5629
g5566 and a[23] n5629_not ; n5630
g5567 nor n5628 n5629 ; n5631
g5568 nor n5630 n5631 ; n5632
g5569 and n5621 n5632_not ; n5633
g5570 nor n5619 n5633 ; n5634
g5571 nor n5550 n5634 ; n5635
g5572 nor n5547 n5635 ; n5636
g5573 nor n5533 n5636 ; n5637
g5574 and n5533 n5636 ; n5638
g5575 nor n5637 n5638 ; n5639
g5576 and n4045_not n5496 ; n5640
g5577 and n3805_not n4935 ; n5641
g5578 and n3964_not n5407 ; n5642
g5579 nor n5641 n5642 ; n5643
g5580 and n5640_not n5643 ; n5644
g5581 and n4477 n4938 ; n5645
g5582 and n5644 n5645_not ; n5646
g5583 and a[20] n5646_not ; n5647
g5584 and a[20] n5647_not ; n5648
g5585 nor n5646 n5647 ; n5649
g5586 nor n5648 n5649 ; n5650
g5587 and n5639 n5650_not ; n5651
g5588 nor n5637 n5651 ; n5652
g5589 and a[15]_not a[16] ; n5653
g5590 and a[15] a[16]_not ; n5654
g5591 nor n5653 n5654 ; n5655
g5592 and a[14] a[15]_not ; n5656
g5593 and a[14]_not a[15] ; n5657
g5594 nor n5656 n5657 ; n5658
g5595 and a[16] a[17]_not ; n5659
g5596 and a[16]_not a[17] ; n5660
g5597 nor n5659 n5660 ; n5661
g5598 and n5658 n5661_not ; n5662
g5599 and n5655 n5662 ; n5663
g5600 and n4515_not n5663 ; n5664
g5601 nor n4522 n5664 ; n5665
g5602 nor n5658 n5661 ; n5666
g5603 nor n5664 n5666 ; n5667
g5604 nor n5665 n5667 ; n5668
g5605 and a[17] n5668_not ; n5669
g5606 and a[17]_not n5668 ; n5670
g5607 nor n5669 n5670 ; n5671
g5608 nor n5652 n5671 ; n5672
g5609 and n5495 n5508_not ; n5673
g5610 nor n5507 n5508 ; n5674
g5611 nor n5673 n5674 ; n5675
g5612 and n5652 n5671 ; n5676
g5613 nor n5672 n5676 ; n5677
g5614 and n5675_not n5677 ; n5678
g5615 nor n5672 n5678 ; n5679
g5616 nor n5523 n5525 ; n5680
g5617 nor n5526 n5680 ; n5681
g5618 and n5679_not n5681 ; n5682
g5619 nor n5675 n5678 ; n5683
g5620 and n5677 n5678_not ; n5684
g5621 nor n5683 n5684 ; n5685
g5622 and n5639 n5651_not ; n5686
g5623 nor n5650 n5651 ; n5687
g5624 nor n5686 n5687 ; n5688
g5625 and n5550 n5634 ; n5689
g5626 nor n5635 n5689 ; n5690
g5627 and n3964_not n5496 ; n5691
g5628 and n3456_not n4935 ; n5692
g5629 and n3805_not n5407 ; n5693
g5630 nor n5692 n5693 ; n5694
g5631 and n5691_not n5694 ; n5695
g5632 and n4938_not n5695 ; n5696
g5633 and n4558_not n5695 ; n5697
g5634 nor n5696 n5697 ; n5698
g5635 and a[20] n5698_not ; n5699
g5636 and a[20]_not n5698 ; n5700
g5637 nor n5699 n5700 ; n5701
g5638 and n5690 n5701_not ; n5702
g5639 and n5621 n5633_not ; n5703
g5640 nor n5632 n5633 ; n5704
g5641 nor n5703 n5704 ; n5705
g5642 and n5605 n5617_not ; n5706
g5643 nor n5616 n5617 ; n5707
g5644 nor n5706 n5707 ; n5708
g5645 and n5598 n5599_not ; n5709
g5646 nor n5596 n5599 ; n5710
g5647 nor n5709 n5710 ; n5711
g5648 and n867_not n3884 ; n5712
g5649 and n1060_not n3967 ; n5713
g5650 and n958_not n4046 ; n5714
g5651 nor n5713 n5714 ; n5715
g5652 and n5712_not n5715 ; n5716
g5653 and n4050_not n5716 ; n5717
g5654 and n4204_not n5716 ; n5718
g5655 nor n5717 n5718 ; n5719
g5656 and a[26] n5719_not ; n5720
g5657 and a[26]_not n5719 ; n5721
g5658 nor n5720 n5721 ; n5722
g5659 nor n5711 n5722 ; n5723
g5660 nor n5577 n5581 ; n5724
g5661 nor n5580 n5581 ; n5725
g5662 nor n5724 n5725 ; n5726
g5663 nor n5335 n5338 ; n5727
g5664 and n5337 n5338_not ; n5728
g5665 nor n5727 n5728 ; n5729
g5666 nor a[8] n5324 ; n5730
g5667 and n5322_not n5325 ; n5731
g5668 nor n5730 n5731 ; n5732
g5669 and n533 n591 ; n5733
g5670 and n296_not n5733 ; n5734
g5671 and n3687 n5734 ; n5735
g5672 and n3583 n5735 ; n5736
g5673 and n1424 n5736 ; n5737
g5674 and n3160 n5737 ; n5738
g5675 and n977 n5738 ; n5739
g5676 and n1575 n5739 ; n5740
g5677 and n469_not n5740 ; n5741
g5678 and n884_not n5741 ; n5742
g5679 and n537_not n5742 ; n5743
g5680 and n1203_not n5743 ; n5744
g5681 and n449_not n5744 ; n5745
g5682 and n655_not n5745 ; n5746
g5683 nor n289 n364 ; n5747
g5684 and n287_not n5747 ; n5748
g5685 and n658 n5748 ; n5749
g5686 and n5269 n5749 ; n5750
g5687 and n824 n5750 ; n5751
g5688 and n5239 n5751 ; n5752
g5689 and n3205 n5752 ; n5753
g5690 and n5746 n5753 ; n5754
g5691 and n2633 n5754 ; n5755
g5692 and n108 n5755 ; n5756
g5693 and n570 n5756 ; n5757
g5694 and n354_not n5757 ; n5758
g5695 and n115_not n5758 ; n5759
g5696 and n177_not n5759 ; n5760
g5697 and n357_not n5760 ; n5761
g5698 and n563_not n5761 ; n5762
g5699 and n173_not n5762 ; n5763
g5700 and n601_not n5763 ; n5764
g5701 and n283_not n5764 ; n5765
g5702 and n5254 n5765_not ; n5766
g5703 and n5254_not n5765 ; n5767
g5704 and n1497 n3524 ; n5768
g5705 and n236_not n5768 ; n5769
g5706 and n504_not n5769 ; n5770
g5707 and n205_not n5770 ; n5771
g5708 and n537_not n5771 ; n5772
g5709 and n666_not n5772 ; n5773
g5710 nor n364 n430 ; n5774
g5711 and n127_not n5774 ; n5775
g5712 nor n281 n328 ; n5776
g5713 and n203_not n5776 ; n5777
g5714 and n5775 n5777 ; n5778
g5715 and n242_not n5778 ; n5779
g5716 and n168_not n5779 ; n5780
g5717 and n884_not n5780 ; n5781
g5718 and n287_not n5781 ; n5782
g5719 and n961_not n5782 ; n5783
g5720 and n86_not n5783 ; n5784
g5721 and n158_not n5784 ; n5785
g5722 nor n451 n932 ; n5786
g5723 and n363_not n5786 ; n5787
g5724 and n136_not n5787 ; n5788
g5725 and n511_not n5788 ; n5789
g5726 and n275_not n5789 ; n5790
g5727 and n228_not n5790 ; n5791
g5728 nor n151 n602 ; n5792
g5729 and n189_not n5792 ; n5793
g5730 and n5791 n5793 ; n5794
g5731 and n5785 n5794 ; n5795
g5732 and n1237 n5795 ; n5796
g5733 and n227 n5796 ; n5797
g5734 and n100 n5797 ; n5798
g5735 and n2758 n5798 ; n5799
g5736 and n620_not n5799 ; n5800
g5737 and n506_not n5800 ; n5801
g5738 and n121_not n5801 ; n5802
g5739 and n527_not n5802 ; n5803
g5740 and n144_not n5803 ; n5804
g5741 and n493_not n5804 ; n5805
g5742 and n1127_not n5805 ; n5806
g5743 nor n330 n449 ; n5807
g5744 and n222_not n5807 ; n5808
g5745 and n2990 n5808 ; n5809
g5746 and n5806 n5809 ; n5810
g5747 and n4388 n5810 ; n5811
g5748 and n616 n5811 ; n5812
g5749 and n5773 n5812 ; n5813
g5750 and n2651 n5813 ; n5814
g5751 and n2940 n5814 ; n5815
g5752 and n520 n5815 ; n5816
g5753 and n847_not n5816 ; n5817
g5754 and n713_not n5817 ; n5818
g5755 and n171_not n5818 ; n5819
g5756 and n460_not n5819 ; n5820
g5757 and n331_not n5820 ; n5821
g5758 and n246_not n5821 ; n5822
g5759 and n623_not n5822 ; n5823
g5760 and n81_not n5823 ; n5824
g5761 and n231_not n5824 ; n5825
g5762 nor a[2] n5825 ; n5826
g5763 and a[2] n5825_not ; n5827
g5764 and a[2]_not n5825 ; n5828
g5765 nor n5827 n5828 ; n5829
g5766 nor a[5] n5829 ; n5830
g5767 nor n5826 n5830 ; n5831
g5768 and n5254 n5831_not ; n5832
g5769 and n2868 n2870_not ; n5833
g5770 nor n2871 n5833 ; n5834
g5771 and n75 n5834 ; n5835
g5772 and n1913_not n3020 ; n5836
g5773 and n2057_not n3023 ; n5837
g5774 and n1992_not n3028 ; n5838
g5775 nor n5837 n5838 ; n5839
g5776 and n5836_not n5839 ; n5840
g5777 and n5835_not n5840 ; n5841
g5778 and n5254_not n5831 ; n5842
g5779 nor n5832 n5842 ; n5843
g5780 and n5841_not n5843 ; n5844
g5781 nor n5832 n5844 ; n5845
g5782 nor n5766 n5845 ; n5846
g5783 and n5767_not n5846 ; n5847
g5784 nor n5766 n5847 ; n5848
g5785 nor n5732 n5848 ; n5849
g5786 and n2876 n2878_not ; n5850
g5787 nor n2879 n5850 ; n5851
g5788 and n75 n5851 ; n5852
g5789 and n1779_not n3020 ; n5853
g5790 and n1913_not n3023 ; n5854
g5791 and n1877_not n3028 ; n5855
g5792 nor n5854 n5855 ; n5856
g5793 and n5853_not n5856 ; n5857
g5794 and n5852_not n5857 ; n5858
g5795 and n5732 n5848 ; n5859
g5796 nor n5849 n5859 ; n5860
g5797 and n5858_not n5860 ; n5861
g5798 nor n5849 n5861 ; n5862
g5799 nor n5729 n5862 ; n5863
g5800 and n5729 n5862 ; n5864
g5801 nor n5863 n5864 ; n5865
g5802 and n1364_not n3457 ; n5866
g5803 and n1572_not n3542 ; n5867
g5804 and n1472_not n3606 ; n5868
g5805 nor n5867 n5868 ; n5869
g5806 and n5866_not n5869 ; n5870
g5807 and n3368_not n5870 ; n5871
g5808 and n5114_not n5870 ; n5872
g5809 nor n5871 n5872 ; n5873
g5810 and a[29] n5873_not ; n5874
g5811 and a[29]_not n5873 ; n5875
g5812 nor n5874 n5875 ; n5876
g5813 and n5865 n5876_not ; n5877
g5814 nor n5863 n5877 ; n5878
g5815 nor n5726 n5878 ; n5879
g5816 and n5726 n5878 ; n5880
g5817 nor n5879 n5880 ; n5881
g5818 and n958_not n3884 ; n5882
g5819 and n1178_not n3967 ; n5883
g5820 and n1060_not n4046 ; n5884
g5821 nor n5883 n5884 ; n5885
g5822 and n5882_not n5885 ; n5886
g5823 and n4050 n4633 ; n5887
g5824 and n5886 n5887_not ; n5888
g5825 and a[26] n5888_not ; n5889
g5826 and a[26] n5889_not ; n5890
g5827 nor n5888 n5889 ; n5891
g5828 nor n5890 n5891 ; n5892
g5829 and n5881 n5892_not ; n5893
g5830 nor n5879 n5893 ; n5894
g5831 and n5711 n5722 ; n5895
g5832 nor n5723 n5895 ; n5896
g5833 and n5894_not n5896 ; n5897
g5834 nor n5723 n5897 ; n5898
g5835 nor n5708 n5898 ; n5899
g5836 and n5708 n5898 ; n5900
g5837 nor n5899 n5900 ; n5901
g5838 and n3012_not n4694 ; n5902
g5839 and n587_not n4533 ; n5903
g5840 and n392_not n4604 ; n5904
g5841 nor n5903 n5904 ; n5905
g5842 and n5902_not n5905 ; n5906
g5843 and n3018 n4536 ; n5907
g5844 and n5906 n5907_not ; n5908
g5845 and a[23] n5908_not ; n5909
g5846 and a[23] n5909_not ; n5910
g5847 nor n5908 n5909 ; n5911
g5848 nor n5910 n5911 ; n5912
g5849 and n5901 n5912_not ; n5913
g5850 nor n5899 n5913 ; n5914
g5851 nor n5705 n5914 ; n5915
g5852 and n5705 n5914 ; n5916
g5853 nor n5915 n5916 ; n5917
g5854 and n3805_not n5496 ; n5918
g5855 and n3605_not n4935 ; n5919
g5856 and n3456_not n5407 ; n5920
g5857 nor n5919 n5920 ; n5921
g5858 and n5918_not n5921 ; n5922
g5859 and n3818 n4938 ; n5923
g5860 and n5922 n5923_not ; n5924
g5861 and a[20] n5924_not ; n5925
g5862 and a[20] n5925_not ; n5926
g5863 nor n5924 n5925 ; n5927
g5864 nor n5926 n5927 ; n5928
g5865 and n5917 n5928_not ; n5929
g5866 nor n5915 n5929 ; n5930
g5867 and n5690_not n5701 ; n5931
g5868 nor n5702 n5931 ; n5932
g5869 and n5930_not n5932 ; n5933
g5870 nor n5702 n5933 ; n5934
g5871 nor n5688 n5934 ; n5935
g5872 and n5688 n5934 ; n5936
g5873 nor n5935 n5936 ; n5937
g5874 and n3877_not n5663 ; n5938
g5875 and n5655_not n5658 ; n5939
g5876 and n4515_not n5939 ; n5940
g5877 nor n5938 n5940 ; n5941
g5878 and n4609 n5666 ; n5942
g5879 and n5941 n5942_not ; n5943
g5880 and a[17] n5943_not ; n5944
g5881 and a[17] n5944_not ; n5945
g5882 nor n5943 n5944 ; n5946
g5883 nor n5945 n5946 ; n5947
g5884 and n5937 n5947_not ; n5948
g5885 nor n5935 n5948 ; n5949
g5886 nor n5685 n5949 ; n5950
g5887 and n5685 n5949 ; n5951
g5888 nor n5950 n5951 ; n5952
g5889 and n5937 n5948_not ; n5953
g5890 nor n5947 n5948 ; n5954
g5891 nor n5953 n5954 ; n5955
g5892 and n5917 n5929_not ; n5956
g5893 nor n5928 n5929 ; n5957
g5894 nor n5956 n5957 ; n5958
g5895 and n5901 n5913_not ; n5959
g5896 nor n5912 n5913 ; n5960
g5897 nor n5959 n5960 ; n5961
g5898 and n392_not n4694 ; n5962
g5899 and n710_not n4533 ; n5963
g5900 and n587_not n4604 ; n5964
g5901 nor n5963 n5964 ; n5965
g5902 and n5962_not n5965 ; n5966
g5903 and n3347 n4536 ; n5967
g5904 and n5966 n5967_not ; n5968
g5905 and a[23] n5968_not ; n5969
g5906 nor n5968 n5969 ; n5970
g5907 and a[23] n5969_not ; n5971
g5908 nor n5970 n5971 ; n5972
g5909 and n5894 n5896_not ; n5973
g5910 nor n5897 n5973 ; n5974
g5911 and n5972_not n5974 ; n5975
g5912 nor n5972 n5975 ; n5976
g5913 and n5974 n5975_not ; n5977
g5914 nor n5976 n5977 ; n5978
g5915 and n5881 n5893_not ; n5979
g5916 nor n5892 n5893 ; n5980
g5917 nor n5979 n5980 ; n5981
g5918 and n1472_not n3457 ; n5982
g5919 and n1665_not n3542 ; n5983
g5920 and n1572_not n3606 ; n5984
g5921 nor n5983 n5984 ; n5985
g5922 and n5982_not n5985 ; n5986
g5923 and n3368 n5139 ; n5987
g5924 and n5986 n5987_not ; n5988
g5925 and a[29] n5988_not ; n5989
g5926 nor n5988 n5989 ; n5990
g5927 and a[29] n5989_not ; n5991
g5928 nor n5990 n5991 ; n5992
g5929 nor n5858 n5861 ; n5993
g5930 and n5860 n5861_not ; n5994
g5931 nor n5993 n5994 ; n5995
g5932 nor n5992 n5995 ; n5996
g5933 nor n5992 n5996 ; n5997
g5934 nor n5995 n5996 ; n5998
g5935 nor n5997 n5998 ; n5999
g5936 nor n5845 n5847 ; n6000
g5937 and n5767_not n5848 ; n6001
g5938 nor n6000 n6001 ; n6002
g5939 and n1877_not n3020 ; n6003
g5940 and n1913_not n3028 ; n6004
g5941 and n1992_not n3023 ; n6005
g5942 and n2872 n2874_not ; n6006
g5943 nor n2875 n6006 ; n6007
g5944 and n75 n6007 ; n6008
g5945 nor n6005 n6008 ; n6009
g5946 and n6004_not n6009 ; n6010
g5947 and n6003_not n6010 ; n6011
g5948 nor n6002 n6011 ; n6012
g5949 nor n5841 n5844 ; n6013
g5950 and n5843 n5844_not ; n6014
g5951 nor n6013 n6014 ; n6015
g5952 and n289_not n2059 ; n6016
g5953 and n620_not n6016 ; n6017
g5954 and n352_not n6017 ; n6018
g5955 and n394_not n6018 ; n6019
g5956 and n603_not n6019 ; n6020
g5957 and n1727 n2705 ; n6021
g5958 and n2556 n6021 ; n6022
g5959 and n330_not n6022 ; n6023
g5960 and n466_not n6023 ; n6024
g5961 and n1680 n6024 ; n6025
g5962 and n270_not n6025 ; n6026
g5963 and n4335 n5152 ; n6027
g5964 and n5056 n6027 ; n6028
g5965 and n1084 n6028 ; n6029
g5966 and n2127 n6029 ; n6030
g5967 and n3580 n6030 ; n6031
g5968 and n6026 n6031 ; n6032
g5969 and n2439 n6032 ; n6033
g5970 and n6020 n6033 ; n6034
g5971 and n1029 n6034 ; n6035
g5972 and n4786 n6035 ; n6036
g5973 and n618 n6036 ; n6037
g5974 and n243_not n6037 ; n6038
g5975 and n519_not n6038 ; n6039
g5976 and n127_not n6039 ; n6040
g5977 and n81_not n6040 ; n6041
g5978 and a[2] n6041_not ; n6042
g5979 and a[2]_not n6041 ; n6043
g5980 and n467 n1611 ; n6044
g5981 and n420_not n6044 ; n6045
g5982 and n1062_not n6045 ; n6046
g5983 and n417_not n6046 ; n6047
g5984 and n400_not n6047 ; n6048
g5985 and n416_not n6048 ; n6049
g5986 and n192_not n6049 ; n6050
g5987 and n563_not n6050 ; n6051
g5988 and n425_not n6051 ; n6052
g5989 and n714_not n6052 ; n6053
g5990 and n243_not n6053 ; n6054
g5991 and n690 n3252 ; n6055
g5992 and n618 n6055 ; n6056
g5993 and n4828 n6056 ; n6057
g5994 and n204 n6057 ; n6058
g5995 and n324 n6058 ; n6059
g5996 and n6054 n6059 ; n6060
g5997 and n2623 n6060 ; n6061
g5998 and n2961 n6061 ; n6062
g5999 and n4274 n6062 ; n6063
g6000 and n604 n6063 ; n6064
g6001 and n454 n6064 ; n6065
g6002 and n423 n6065 ; n6066
g6003 and n731 n6066 ; n6067
g6004 and n1379 n6067 ; n6068
g6005 and n149_not n6068 ; n6069
g6006 and n246_not n6069 ; n6070
g6007 and n791_not n6070 ; n6071
g6008 and n592_not n6071 ; n6072
g6009 and n886_not n6072 ; n6073
g6010 and n449_not n6073 ; n6074
g6011 and a[2] n6074_not ; n6075
g6012 and a[2]_not n6074 ; n6076
g6013 and n1426 n1644 ; n6077
g6014 and n190_not n6077 ; n6078
g6015 and n239_not n6078 ; n6079
g6016 and n637_not n6079 ; n6080
g6017 and n305_not n6080 ; n6081
g6018 and n130_not n6081 ; n6082
g6019 and n1010_not n6082 ; n6083
g6020 nor n295 n395 ; n6084
g6021 and n2593 n5150 ; n6085
g6022 and n1438 n6085 ; n6086
g6023 and n6084 n6086 ; n6087
g6024 and n5193 n6087 ; n6088
g6025 and n1601 n6088 ; n6089
g6026 and n1029 n6089 ; n6090
g6027 and n454 n6090 ; n6091
g6028 and n979 n6091 ; n6092
g6029 and n752_not n6092 ; n6093
g6030 and n224_not n6093 ; n6094
g6031 and n275_not n6094 ; n6095
g6032 and n226_not n6095 ; n6096
g6033 and n451_not n6096 ; n6097
g6034 and n590 n1072_not ; n6098
g6035 and n206_not n6098 ; n6099
g6036 and n714_not n6099 ; n6100
g6037 and n689_not n6100 ; n6101
g6038 and n474_not n6101 ; n6102
g6039 and n111_not n4367 ; n6103
g6040 and n603_not n6103 ; n6104
g6041 and n4269 n6104 ; n6105
g6042 and n2241 n6105 ; n6106
g6043 and n2807 n6106 ; n6107
g6044 and n6102 n6107 ; n6108
g6045 and n2751 n6108 ; n6109
g6046 and n6097 n6109 ; n6110
g6047 and n6083 n6110 ; n6111
g6048 and n333 n6111 ; n6112
g6049 and n1291 n6112 ; n6113
g6050 and n4786 n6113 ; n6114
g6051 and n201_not n6114 ; n6115
g6052 and n564_not n6115 ; n6116
g6053 and n489_not n6116 ; n6117
g6054 and n886_not n6117 ; n6118
g6055 and a[2] n6118_not ; n6119
g6056 and a[2]_not n6118 ; n6120
g6057 and n2852 n2854_not ; n6121
g6058 nor n2855 n6121 ; n6122
g6059 and n75 n6122 ; n6123
g6060 and n2189_not n3020 ; n6124
g6061 and n2388_not n3023 ; n6125
g6062 and n2291_not n3028 ; n6126
g6063 nor n6125 n6126 ; n6127
g6064 and n6124_not n6127 ; n6128
g6065 and n6123_not n6128 ; n6129
g6066 nor n6119 n6129 ; n6130
g6067 and n6120_not n6130 ; n6131
g6068 nor n6119 n6131 ; n6132
g6069 nor n6075 n6132 ; n6133
g6070 and n6076_not n6133 ; n6134
g6071 nor n6075 n6134 ; n6135
g6072 nor n6042 n6135 ; n6136
g6073 and n6043_not n6136 ; n6137
g6074 nor n6042 n6137 ; n6138
g6075 and a[5] n5829 ; n6139
g6076 nor n5830 n6139 ; n6140
g6077 and n6138_not n6140 ; n6141
g6078 and n2864 n2866_not ; n6142
g6079 nor n2867 n6142 ; n6143
g6080 and n75 n6143 ; n6144
g6081 and n1992_not n3020 ; n6145
g6082 and n2152_not n3023 ; n6146
g6083 and n2057_not n3028 ; n6147
g6084 nor n6146 n6147 ; n6148
g6085 and n6145_not n6148 ; n6149
g6086 and n6144_not n6149 ; n6150
g6087 and n6138 n6140_not ; n6151
g6088 nor n6141 n6151 ; n6152
g6089 and n6150_not n6152 ; n6153
g6090 nor n6141 n6153 ; n6154
g6091 nor n6015 n6154 ; n6155
g6092 and n6015 n6154 ; n6156
g6093 nor n6155 n6156 ; n6157
g6094 and n1665_not n3457 ; n6158
g6095 and n1877_not n3542 ; n6159
g6096 and n1779_not n3606 ; n6160
g6097 nor n6159 n6160 ; n6161
g6098 and n6158_not n6161 ; n6162
g6099 and n3368_not n6162 ; n6163
g6100 and n5328_not n6162 ; n6164
g6101 nor n6163 n6164 ; n6165
g6102 and a[29] n6165_not ; n6166
g6103 and a[29]_not n6165 ; n6167
g6104 nor n6166 n6167 ; n6168
g6105 and n6157 n6168_not ; n6169
g6106 nor n6155 n6169 ; n6170
g6107 nor n6002 n6012 ; n6171
g6108 nor n6011 n6012 ; n6172
g6109 nor n6171 n6172 ; n6173
g6110 nor n6170 n6173 ; n6174
g6111 nor n6012 n6174 ; n6175
g6112 nor n5999 n6175 ; n6176
g6113 nor n5996 n6176 ; n6177
g6114 and n5865_not n5876 ; n6178
g6115 nor n5877 n6178 ; n6179
g6116 and n6177_not n6179 ; n6180
g6117 and n6177 n6179_not ; n6181
g6118 nor n6180 n6181 ; n6182
g6119 and n1060_not n3884 ; n6183
g6120 and n1235_not n3967 ; n6184
g6121 and n1178_not n4046 ; n6185
g6122 nor n6184 n6185 ; n6186
g6123 and n6183_not n6186 ; n6187
g6124 and n4050 n4429 ; n6188
g6125 and n6187 n6188_not ; n6189
g6126 and a[26] n6189_not ; n6190
g6127 and a[26] n6190_not ; n6191
g6128 nor n6189 n6190 ; n6192
g6129 nor n6191 n6192 ; n6193
g6130 and n6182 n6193_not ; n6194
g6131 nor n6180 n6194 ; n6195
g6132 nor n5981 n6195 ; n6196
g6133 and n5981 n6195 ; n6197
g6134 nor n6196 n6197 ; n6198
g6135 and n587_not n4694 ; n6199
g6136 and n867_not n4533 ; n6200
g6137 and n710_not n4604 ; n6201
g6138 nor n6200 n6201 ; n6202
g6139 and n6199_not n6202 ; n6203
g6140 and n3331 n4536 ; n6204
g6141 and n6203 n6204_not ; n6205
g6142 and a[23] n6205_not ; n6206
g6143 and a[23] n6206_not ; n6207
g6144 nor n6205 n6206 ; n6208
g6145 nor n6207 n6208 ; n6209
g6146 and n6198 n6209_not ; n6210
g6147 nor n6196 n6210 ; n6211
g6148 nor n5978 n6211 ; n6212
g6149 nor n5975 n6212 ; n6213
g6150 nor n5961 n6213 ; n6214
g6151 and n5961 n6213 ; n6215
g6152 nor n6214 n6215 ; n6216
g6153 and n3456_not n5496 ; n6217
g6154 and n3539_not n4935 ; n6218
g6155 and n3605_not n5407 ; n6219
g6156 nor n6218 n6219 ; n6220
g6157 and n6217_not n6220 ; n6221
g6158 and n3627 n4938 ; n6222
g6159 and n6221 n6222_not ; n6223
g6160 and a[20] n6223_not ; n6224
g6161 and a[20] n6224_not ; n6225
g6162 nor n6223 n6224 ; n6226
g6163 nor n6225 n6226 ; n6227
g6164 and n6216 n6227_not ; n6228
g6165 nor n6214 n6228 ; n6229
g6166 nor n5958 n6229 ; n6230
g6167 and n5958 n6229 ; n6231
g6168 nor n6230 n6231 ; n6232
g6169 and n5658_not n5661 ; n6233
g6170 and n3877_not n6233 ; n6234
g6171 and n3964_not n5663 ; n6235
g6172 and n4045_not n5939 ; n6236
g6173 nor n6235 n6236 ; n6237
g6174 and n6234_not n6237 ; n6238
g6175 and n4067 n5666 ; n6239
g6176 and n6238 n6239_not ; n6240
g6177 and a[17] n6240_not ; n6241
g6178 and a[17] n6241_not ; n6242
g6179 nor n6240 n6241 ; n6243
g6180 nor n6242 n6243 ; n6244
g6181 and n6232 n6244_not ; n6245
g6182 nor n6230 n6245 ; n6246
g6183 and n4515_not n6233 ; n6247
g6184 and n4045_not n5663 ; n6248
g6185 and n3877_not n5939 ; n6249
g6186 nor n6248 n6249 ; n6250
g6187 and n6247_not n6250 ; n6251
g6188 and n5666_not n6251 ; n6252
g6189 and n4715_not n6251 ; n6253
g6190 nor n6252 n6253 ; n6254
g6191 and a[17] n6254_not ; n6255
g6192 and a[17]_not n6254 ; n6256
g6193 nor n6255 n6256 ; n6257
g6194 nor n6246 n6257 ; n6258
g6195 and n6246 n6257 ; n6259
g6196 nor n6258 n6259 ; n6260
g6197 and n5930 n5932_not ; n6261
g6198 nor n5933 n6261 ; n6262
g6199 and n6260 n6262 ; n6263
g6200 nor n6258 n6263 ; n6264
g6201 nor n5955 n6264 ; n6265
g6202 and n5955 n6264 ; n6266
g6203 nor n6265 n6266 ; n6267
g6204 and n6216 n6228_not ; n6268
g6205 nor n6227 n6228 ; n6269
g6206 nor n6268 n6269 ; n6270
g6207 and n5978 n6211 ; n6271
g6208 nor n6212 n6271 ; n6272
g6209 and n3605_not n5496 ; n6273
g6210 and n3012_not n4935 ; n6274
g6211 and n3539_not n5407 ; n6275
g6212 nor n6274 n6275 ; n6276
g6213 and n6273_not n6276 ; n6277
g6214 and n4938_not n6277 ; n6278
g6215 and n4084_not n6277 ; n6279
g6216 nor n6278 n6279 ; n6280
g6217 and a[20] n6280_not ; n6281
g6218 and a[20]_not n6280 ; n6282
g6219 nor n6281 n6282 ; n6283
g6220 and n6272 n6283_not ; n6284
g6221 and n6198 n6210_not ; n6285
g6222 nor n6209 n6210 ; n6286
g6223 nor n6285 n6286 ; n6287
g6224 and n6182 n6194_not ; n6288
g6225 nor n6193 n6194 ; n6289
g6226 nor n6288 n6289 ; n6290
g6227 and n5999 n6175 ; n6291
g6228 nor n6176 n6291 ; n6292
g6229 and n1178_not n3884 ; n6293
g6230 and n1364_not n3967 ; n6294
g6231 and n1235_not n4046 ; n6295
g6232 nor n6294 n6295 ; n6296
g6233 and n6293_not n6296 ; n6297
g6234 and n4050_not n6297 ; n6298
g6235 and n4861_not n6297 ; n6299
g6236 nor n6298 n6299 ; n6300
g6237 and a[26] n6300_not ; n6301
g6238 and a[26]_not n6300 ; n6302
g6239 nor n6301 n6302 ; n6303
g6240 and n6292 n6303_not ; n6304
g6241 nor n6170 n6174 ; n6305
g6242 nor n6173 n6174 ; n6306
g6243 nor n6305 n6306 ; n6307
g6244 and n1572_not n3457 ; n6308
g6245 and n1779_not n3542 ; n6309
g6246 and n1665_not n3606 ; n6310
g6247 nor n6309 n6310 ; n6311
g6248 and n6308_not n6311 ; n6312
g6249 and n3368_not n6312 ; n6313
g6250 and n5561_not n6312 ; n6314
g6251 nor n6313 n6314 ; n6315
g6252 and a[29] n6315_not ; n6316
g6253 and a[29]_not n6315 ; n6317
g6254 nor n6316 n6317 ; n6318
g6255 nor n6307 n6318 ; n6319
g6256 and n6307 n6318 ; n6320
g6257 nor n6319 n6320 ; n6321
g6258 and n1235_not n3884 ; n6322
g6259 and n1472_not n3967 ; n6323
g6260 and n1364_not n4046 ; n6324
g6261 nor n6323 n6324 ; n6325
g6262 and n6322_not n6325 ; n6326
g6263 and n4050 n4848 ; n6327
g6264 and n6326 n6327_not ; n6328
g6265 and a[26] n6328_not ; n6329
g6266 and a[26] n6329_not ; n6330
g6267 nor n6328 n6329 ; n6331
g6268 nor n6330 n6331 ; n6332
g6269 and n6321 n6332_not ; n6333
g6270 nor n6319 n6333 ; n6334
g6271 and n6292_not n6303 ; n6335
g6272 nor n6304 n6335 ; n6336
g6273 and n6334_not n6336 ; n6337
g6274 nor n6304 n6337 ; n6338
g6275 nor n6290 n6338 ; n6339
g6276 and n6290 n6338 ; n6340
g6277 nor n6339 n6340 ; n6341
g6278 and n710_not n4694 ; n6342
g6279 and n958_not n4533 ; n6343
g6280 and n867_not n4604 ; n6344
g6281 nor n6343 n6344 ; n6345
g6282 and n6342_not n6345 ; n6346
g6283 and n4179 n4536 ; n6347
g6284 and n6346 n6347_not ; n6348
g6285 and a[23] n6348_not ; n6349
g6286 and a[23] n6349_not ; n6350
g6287 nor n6348 n6349 ; n6351
g6288 nor n6350 n6351 ; n6352
g6289 and n6341 n6352_not ; n6353
g6290 nor n6339 n6353 ; n6354
g6291 nor n6287 n6354 ; n6355
g6292 and n6287 n6354 ; n6356
g6293 nor n6355 n6356 ; n6357
g6294 and n3539_not n5496 ; n6358
g6295 and n392_not n4935 ; n6359
g6296 and n3012_not n5407 ; n6360
g6297 nor n6359 n6360 ; n6361
g6298 and n6358_not n6361 ; n6362
g6299 and n3715 n4938 ; n6363
g6300 and n6362 n6363_not ; n6364
g6301 and a[20] n6364_not ; n6365
g6302 and a[20] n6365_not ; n6366
g6303 nor n6364 n6365 ; n6367
g6304 nor n6366 n6367 ; n6368
g6305 and n6357 n6368_not ; n6369
g6306 nor n6355 n6369 ; n6370
g6307 and n6272_not n6283 ; n6371
g6308 nor n6284 n6371 ; n6372
g6309 and n6370_not n6372 ; n6373
g6310 nor n6284 n6373 ; n6374
g6311 nor n6270 n6374 ; n6375
g6312 and n6270 n6374 ; n6376
g6313 nor n6375 n6376 ; n6377
g6314 and n4045_not n6233 ; n6378
g6315 and n3805_not n5663 ; n6379
g6316 and n3964_not n5939 ; n6380
g6317 nor n6379 n6380 ; n6381
g6318 and n6378_not n6381 ; n6382
g6319 and n4477 n5666 ; n6383
g6320 and n6382 n6383_not ; n6384
g6321 and a[17] n6384_not ; n6385
g6322 and a[17] n6385_not ; n6386
g6323 nor n6384 n6385 ; n6387
g6324 nor n6386 n6387 ; n6388
g6325 and n6377 n6388_not ; n6389
g6326 nor n6375 n6389 ; n6390
g6327 and a[11] a[12]_not ; n6391
g6328 and a[11]_not a[12] ; n6392
g6329 nor n6391 n6392 ; n6393
g6330 and a[13] a[14]_not ; n6394
g6331 and a[13]_not a[14] ; n6395
g6332 nor n6394 n6395 ; n6396
g6333 nor n6393 n6396 ; n6397
g6334 and a[12]_not a[13] ; n6398
g6335 and a[12] a[13]_not ; n6399
g6336 nor n6398 n6399 ; n6400
g6337 and n6393 n6396_not ; n6401
g6338 and n6400 n6401 ; n6402
g6339 and n4515_not n6402 ; n6403
g6340 nor n6397 n6403 ; n6404
g6341 nor n4522 n6403 ; n6405
g6342 nor n6404 n6405 ; n6406
g6343 and a[14] n6406_not ; n6407
g6344 and a[14]_not n6406 ; n6408
g6345 nor n6407 n6408 ; n6409
g6346 nor n6390 n6409 ; n6410
g6347 and n6232 n6245_not ; n6411
g6348 nor n6244 n6245 ; n6412
g6349 nor n6411 n6412 ; n6413
g6350 and n6390 n6409 ; n6414
g6351 nor n6410 n6414 ; n6415
g6352 and n6413_not n6415 ; n6416
g6353 nor n6410 n6416 ; n6417
g6354 nor n6260 n6262 ; n6418
g6355 nor n6263 n6418 ; n6419
g6356 and n6417_not n6419 ; n6420
g6357 and n6417 n6419_not ; n6421
g6358 nor n6420 n6421 ; n6422
g6359 nor n6413 n6416 ; n6423
g6360 and n6415 n6416_not ; n6424
g6361 nor n6423 n6424 ; n6425
g6362 and n3964_not n6233 ; n6426
g6363 and n3456_not n5663 ; n6427
g6364 and n3805_not n5939 ; n6428
g6365 nor n6427 n6428 ; n6429
g6366 and n6426_not n6429 ; n6430
g6367 and n4558 n5666 ; n6431
g6368 and n6430 n6431_not ; n6432
g6369 and a[17] n6432_not ; n6433
g6370 nor n6432 n6433 ; n6434
g6371 and a[17] n6433_not ; n6435
g6372 nor n6434 n6435 ; n6436
g6373 and n6370 n6372_not ; n6437
g6374 nor n6373 n6437 ; n6438
g6375 and n6436_not n6438 ; n6439
g6376 nor n6436 n6439 ; n6440
g6377 and n6438 n6439_not ; n6441
g6378 nor n6440 n6441 ; n6442
g6379 and n6357 n6369_not ; n6443
g6380 nor n6368 n6369 ; n6444
g6381 nor n6443 n6444 ; n6445
g6382 and n6341 n6353_not ; n6446
g6383 nor n6352 n6353 ; n6447
g6384 nor n6446 n6447 ; n6448
g6385 and n867_not n4694 ; n6449
g6386 and n1060_not n4533 ; n6450
g6387 and n958_not n4604 ; n6451
g6388 nor n6450 n6451 ; n6452
g6389 and n6449_not n6452 ; n6453
g6390 and n4204 n4536 ; n6454
g6391 and n6453 n6454_not ; n6455
g6392 and a[23] n6455_not ; n6456
g6393 nor n6455 n6456 ; n6457
g6394 and a[23] n6456_not ; n6458
g6395 nor n6457 n6458 ; n6459
g6396 and n6334 n6336_not ; n6460
g6397 nor n6337 n6460 ; n6461
g6398 and n6459_not n6461 ; n6462
g6399 nor n6459 n6462 ; n6463
g6400 and n6461 n6462_not ; n6464
g6401 nor n6463 n6464 ; n6465
g6402 and n6321 n6333_not ; n6466
g6403 nor n6332 n6333 ; n6467
g6404 nor n6466 n6467 ; n6468
g6405 and n6152 n6153_not ; n6469
g6406 nor n6150 n6153 ; n6470
g6407 nor n6469 n6470 ; n6471
g6408 nor n6135 n6137 ; n6472
g6409 and n6043_not n6138 ; n6473
g6410 nor n6472 n6473 ; n6474
g6411 and n2057_not n3020 ; n6475
g6412 and n2152_not n3028 ; n6476
g6413 and n2189_not n3023 ; n6477
g6414 and n2860 n2862_not ; n6478
g6415 nor n2863 n6478 ; n6479
g6416 and n75 n6479 ; n6480
g6417 nor n6477 n6480 ; n6481
g6418 and n6476_not n6481 ; n6482
g6419 and n6475_not n6482 ; n6483
g6420 nor n6474 n6483 ; n6484
g6421 nor n6132 n6134 ; n6485
g6422 and n6076_not n6135 ; n6486
g6423 nor n6485 n6486 ; n6487
g6424 and n2152_not n3020 ; n6488
g6425 and n2189_not n3028 ; n6489
g6426 and n2291_not n3023 ; n6490
g6427 and n2856 n2858_not ; n6491
g6428 nor n2859 n6491 ; n6492
g6429 and n75 n6492 ; n6493
g6430 nor n6490 n6493 ; n6494
g6431 and n6489_not n6494 ; n6495
g6432 and n6488_not n6495 ; n6496
g6433 nor n6487 n6496 ; n6497
g6434 nor n6129 n6131 ; n6498
g6435 and n6120_not n6132 ; n6499
g6436 nor n6498 n6499 ; n6500
g6437 and n2608 n4357 ; n6501
g6438 and n4828 n6501 ; n6502
g6439 and n4279 n6502 ; n6503
g6440 and n1794 n6503 ; n6504
g6441 and n1292 n6504 ; n6505
g6442 and n874 n6505 ; n6506
g6443 and n1139 n6506 ; n6507
g6444 and n2993 n6507 ; n6508
g6445 and n116 n6508 ; n6509
g6446 and n617_not n6509 ; n6510
g6447 and n254_not n6510 ; n6511
g6448 and n809_not n6511 ; n6512
g6449 and n368_not n6512 ; n6513
g6450 and n791_not n6513 ; n6514
g6451 and n175_not n5171 ; n6515
g6452 and n206_not n6515 ; n6516
g6453 and n655_not n6516 ; n6517
g6454 nor n123 n518 ; n6518
g6455 and n157_not n6518 ; n6519
g6456 and n270_not n6519 ; n6520
g6457 and n3524 n5775 ; n6521
g6458 and n691 n6521 ; n6522
g6459 and n6520 n6522 ; n6523
g6460 and n6517 n6523 ; n6524
g6461 and n1709 n6524 ; n6525
g6462 and n4405 n6525 ; n6526
g6463 and n4375 n6526 ; n6527
g6464 and n6514 n6527 ; n6528
g6465 and n454 n6528 ; n6529
g6466 and n731 n6529 ; n6530
g6467 and n1478 n6530 ; n6531
g6468 and n136_not n6531 ; n6532
g6469 and n248_not n6532 ; n6533
g6470 and n298_not n6533 ; n6534
g6471 and n273_not n6534 ; n6535
g6472 and n436_not n6535 ; n6536
g6473 and n2291_not n3020 ; n6537
g6474 and n2388_not n3028 ; n6538
g6475 and n2464_not n3023 ; n6539
g6476 and n2848 n2850_not ; n6540
g6477 nor n2851 n6540 ; n6541
g6478 and n75 n6541 ; n6542
g6479 nor n6539 n6542 ; n6543
g6480 and n6538_not n6543 ; n6544
g6481 and n6537_not n6544 ; n6545
g6482 nor n6536 n6545 ; n6546
g6483 nor n278 n396 ; n6547
g6484 and n532_not n6547 ; n6548
g6485 and n5021 n6548 ; n6549
g6486 and n1785 n6549 ; n6550
g6487 and n1586 n6550 ; n6551
g6488 and n4127 n6551 ; n6552
g6489 and n2583 n6552 ; n6553
g6490 and n100 n6553 ; n6554
g6491 and n667_not n6554 ; n6555
g6492 and n641_not n6555 ; n6556
g6493 and n189_not n6556 ; n6557
g6494 and n107_not n6557 ; n6558
g6495 and n777_not n6558 ; n6559
g6496 and n564_not n6559 ; n6560
g6497 and n81_not n6560 ; n6561
g6498 and n423 n1062_not ; n6562
g6499 and n884_not n6562 ; n6563
g6500 and n298_not n6563 ; n6564
g6501 and n525_not n6564 ; n6565
g6502 and n284_not n1128 ; n6566
g6503 and n460_not n6566 ; n6567
g6504 and n1740 n3416 ; n6568
g6505 and n2220 n6568 ; n6569
g6506 and n6567 n6569 ; n6570
g6507 and n1692 n6570 ; n6571
g6508 and n6565 n6571 ; n6572
g6509 and n877 n6572 ; n6573
g6510 and n1709 n6573 ; n6574
g6511 and n268 n6574 ; n6575
g6512 and n4367 n6575 ; n6576
g6513 and n6561 n6576 ; n6577
g6514 and n5063 n6577 ; n6578
g6515 and n450 n6578 ; n6579
g6516 and n1761 n6579 ; n6580
g6517 and n194_not n6580 ; n6581
g6518 and n151_not n6581 ; n6582
g6519 and n275_not n6582 ; n6583
g6520 and n173_not n6583 ; n6584
g6521 and n493_not n6584 ; n6585
g6522 and n200_not n6585 ; n6586
g6523 and n2388_not n3020 ; n6587
g6524 and n2464_not n3028 ; n6588
g6525 and n2533_not n3023 ; n6589
g6526 and n2844 n2846_not ; n6590
g6527 nor n2847 n6590 ; n6591
g6528 and n75 n6591 ; n6592
g6529 nor n6589 n6592 ; n6593
g6530 and n6588_not n6593 ; n6594
g6531 and n6587_not n6594 ; n6595
g6532 nor n6586 n6595 ; n6596
g6533 and n918 n2191 ; n6597
g6534 and n279 n6597 ; n6598
g6535 and n100 n6598 ; n6599
g6536 and n289_not n6599 ; n6600
g6537 and n803_not n6600 ; n6601
g6538 and n246_not n6601 ; n6602
g6539 and n466_not n6602 ; n6603
g6540 and n672_not n6603 ; n6604
g6541 and n328_not n515 ; n6605
g6542 and n396_not n6605 ; n6606
g6543 and n468_not n6606 ; n6607
g6544 and n752_not n1824 ; n6608
g6545 and n716_not n6608 ; n6609
g6546 and n489_not n6609 ; n6610
g6547 and n1424 n1588 ; n6611
g6548 and n6610 n6611 ; n6612
g6549 and n6607 n6612 ; n6613
g6550 and n5148 n6613 ; n6614
g6551 and n720 n6614 ; n6615
g6552 and n634 n6615 ; n6616
g6553 and n398_not n6616 ; n6617
g6554 and n152_not n6617 ; n6618
g6555 and n354_not n6618 ; n6619
g6556 and n777_not n6619 ; n6620
g6557 and n416_not n6620 ; n6621
g6558 and n368_not n6621 ; n6622
g6559 and n932_not n6622 ; n6623
g6560 and n272_not n6623 ; n6624
g6561 and n712_not n6624 ; n6625
g6562 and n558_not n2169 ; n6626
g6563 and n339_not n6626 ; n6627
g6564 and n327_not n6627 ; n6628
g6565 and n172 n1497 ; n6629
g6566 and n6628 n6629 ; n6630
g6567 and n2370 n6630 ; n6631
g6568 and n3768 n6631 ; n6632
g6569 and n5224 n6632 ; n6633
g6570 and n6625 n6633 ; n6634
g6571 and n6604 n6634 ; n6635
g6572 and n353_not n6635 ; n6636
g6573 and n367_not n6636 ; n6637
g6574 and n825_not n6637 ; n6638
g6575 and n191_not n6638 ; n6639
g6576 and n225_not n6639 ; n6640
g6577 and n436_not n6640 ; n6641
g6578 and n2464_not n3020 ; n6642
g6579 and n2533_not n3028 ; n6643
g6580 and n2571_not n3023 ; n6644
g6581 and n2840 n2842_not ; n6645
g6582 nor n2843 n6645 ; n6646
g6583 and n75 n6646 ; n6647
g6584 nor n6644 n6647 ; n6648
g6585 and n6643_not n6648 ; n6649
g6586 and n6642_not n6649 ; n6650
g6587 nor n6641 n6650 ; n6651
g6588 and n3314 n3549 ; n6652
g6589 and n3409 n6652 ; n6653
g6590 and n1105 n6653 ; n6654
g6591 and n1523 n6654 ; n6655
g6592 and n123_not n6655 ; n6656
g6593 and n427_not n6656 ; n6657
g6594 and n329_not n6657 ; n6658
g6595 and n328_not n6658 ; n6659
g6596 and n402_not n6659 ; n6660
g6597 and n430_not n6660 ; n6661
g6598 and n340_not n6661 ; n6662
g6599 nor n358 n518 ; n6663
g6600 and n428_not n6663 ; n6664
g6601 and n827 n6664 ; n6665
g6602 and n306_not n6665 ; n6666
g6603 and n158_not n6666 ; n6667
g6604 nor n161 n531 ; n6668
g6605 and n304_not n6668 ; n6669
g6606 and n222_not n6669 ; n6670
g6607 and n280_not n604 ; n6671
g6608 and n332_not n6671 ; n6672
g6609 and n1578 n6672 ; n6673
g6610 and n4269 n6673 ; n6674
g6611 and n6670 n6674 ; n6675
g6612 and n6667 n6675 ; n6676
g6613 and n2258 n6676 ; n6677
g6614 and n6662 n6677 ; n6678
g6615 and n805 n6678 ; n6679
g6616 and n2573 n6679 ; n6680
g6617 and n1531 n6680 ; n6681
g6618 and n1141 n6681 ; n6682
g6619 and n978 n6682 ; n6683
g6620 and n1161 n6683 ; n6684
g6621 and n353_not n6684 ; n6685
g6622 and n299_not n6685 ; n6686
g6623 and n490_not n6686 ; n6687
g6624 and n568_not n6687 ; n6688
g6625 and n164_not n6688 ; n6689
g6626 and n623_not n6689 ; n6690
g6627 and n2533_not n3020 ; n6691
g6628 and n2571_not n3028 ; n6692
g6629 and n2674_not n3023 ; n6693
g6630 and n2836 n2838_not ; n6694
g6631 nor n2839 n6694 ; n6695
g6632 and n75 n6695 ; n6696
g6633 nor n6693 n6696 ; n6697
g6634 and n6692_not n6697 ; n6698
g6635 and n6691_not n6698 ; n6699
g6636 nor n6690 n6699 ; n6700
g6637 and n300 n301_not ; n6701
g6638 and n1102_not n6701 ; n6702
g6639 and n203_not n6702 ; n6703
g6640 and n326_not n6703 ; n6704
g6641 and n287_not n6704 ; n6705
g6642 nor n145 n164 ; n6706
g6643 and n536_not n6706 ; n6707
g6644 and n1528 n1617 ; n6708
g6645 and n2633 n6708 ; n6709
g6646 and n3886 n6709 ; n6710
g6647 and n715_not n6710 ; n6711
g6648 and n372_not n6711 ; n6712
g6649 and n366_not n6712 ; n6713
g6650 and n633_not n6713 ; n6714
g6651 and n132_not n3581 ; n6715
g6652 and n201_not n6715 ; n6716
g6653 and n557_not n2089 ; n6717
g6654 and n2423 n6717 ; n6718
g6655 and n6716 n6718 ; n6719
g6656 and n897 n6719 ; n6720
g6657 and n1476 n6720 ; n6721
g6658 and n665 n6721 ; n6722
g6659 and n6714 n6722 ; n6723
g6660 and n1531 n6723 ; n6724
g6661 and n826 n6724 ; n6725
g6662 and n227 n6725 ; n6726
g6663 and n518_not n6726 ; n6727
g6664 and n1101_not n6727 ; n6728
g6665 and n192_not n6728 ; n6729
g6666 and n932_not n6729 ; n6730
g6667 and n474_not n6730 ; n6731
g6668 and n532_not n6731 ; n6732
g6669 and n233_not n885 ; n6733
g6670 and n144_not n6733 ; n6734
g6671 and n1221 n6734 ; n6735
g6672 and n1615 n6735 ; n6736
g6673 and n2632 n6736 ; n6737
g6674 and n1454 n6737 ; n6738
g6675 and n6732 n6738 ; n6739
g6676 and n6707 n6739 ; n6740
g6677 and n2021 n6740 ; n6741
g6678 and n6705 n6741 ; n6742
g6679 and n331_not n6742 ; n6743
g6680 and n272_not n6743 ; n6744
g6681 and n451_not n6744 ; n6745
g6682 and n1104_not n6745 ; n6746
g6683 and n562_not n6746 ; n6747
g6684 and n655_not n6747 ; n6748
g6685 and n300 n2704 ; n6749
g6686 and n111_not n6749 ; n6750
g6687 and n1306_not n6750 ; n6751
g6688 and n374_not n6751 ; n6752
g6689 and n563_not n6752 ; n6753
g6690 and n331_not n6753 ; n6754
g6691 and n371_not n6754 ; n6755
g6692 and n5201 n5793 ; n6756
g6693 and n776 n6756 ; n6757
g6694 and n467 n6757 ; n6758
g6695 and n6670 n6758 ; n6759
g6696 and n2738 n6759 ; n6760
g6697 and n873 n6760 ; n6761
g6698 and n2010 n6761 ; n6762
g6699 and n1824 n6762 ; n6763
g6700 and n2073 n6763 ; n6764
g6701 and n716_not n6764 ; n6765
g6702 and n422_not n6765 ; n6766
g6703 and n394_not n6766 ; n6767
g6704 and n603_not n6767 ; n6768
g6705 and n883_not n6768 ; n6769
g6706 and n1127_not n3636 ; n6770
g6707 and n633_not n6770 ; n6771
g6708 and n735 n1586 ; n6772
g6709 and n6771 n6772 ; n6773
g6710 and n4148 n6773 ; n6774
g6711 and n2104 n6774 ; n6775
g6712 and n6769 n6775 ; n6776
g6713 and n6755 n6776 ; n6777
g6714 and n510 n6777 ; n6778
g6715 and n1668 n6778 ; n6779
g6716 and n288 n6779 ; n6780
g6717 and n869 n6780 ; n6781
g6718 and n2466 n6781 ; n6782
g6719 and n810 n6782 ; n6783
g6720 and n236_not n6783 ; n6784
g6721 and n289_not n6784 ; n6785
g6722 and n254_not n6785 ; n6786
g6723 and n511_not n6786 ; n6787
g6724 and n203_not n6787 ; n6788
g6725 and n367_not n6788 ; n6789
g6726 and n777_not n6789 ; n6790
g6727 and n246_not n6790 ; n6791
g6728 and n2674_not n3020 ; n6792
g6729 and n2736_not n3028 ; n6793
g6730 and n2829_not n3023 ; n6794
g6731 and n2736_not n2829 ; n6795
g6732 and n2674 n6795_not ; n6796
g6733 and n2737 n2829 ; n6797
g6734 nor n6796 n6797 ; n6798
g6735 and n75 n6798 ; n6799
g6736 nor n6794 n6799 ; n6800
g6737 and n6793_not n6800 ; n6801
g6738 and n6792_not n6801 ; n6802
g6739 nor n6791 n6802 ; n6803
g6740 and n6748_not n6803 ; n6804
g6741 and n2832 n2834_not ; n6805
g6742 nor n2835 n6805 ; n6806
g6743 and n75 n6806 ; n6807
g6744 and n2571_not n3020 ; n6808
g6745 and n2736_not n3023 ; n6809
g6746 and n2674_not n3028 ; n6810
g6747 nor n6809 n6810 ; n6811
g6748 and n6808_not n6811 ; n6812
g6749 and n6807_not n6812 ; n6813
g6750 and n6748 n6803_not ; n6814
g6751 nor n6804 n6814 ; n6815
g6752 and n6813_not n6815 ; n6816
g6753 nor n6804 n6816 ; n6817
g6754 nor n6690 n6700 ; n6818
g6755 nor n6699 n6700 ; n6819
g6756 nor n6818 n6819 ; n6820
g6757 nor n6817 n6820 ; n6821
g6758 nor n6700 n6821 ; n6822
g6759 nor n6641 n6651 ; n6823
g6760 nor n6650 n6651 ; n6824
g6761 nor n6823 n6824 ; n6825
g6762 nor n6822 n6825 ; n6826
g6763 nor n6651 n6826 ; n6827
g6764 nor n6586 n6596 ; n6828
g6765 nor n6595 n6596 ; n6829
g6766 nor n6828 n6829 ; n6830
g6767 nor n6827 n6830 ; n6831
g6768 nor n6596 n6831 ; n6832
g6769 nor n6536 n6546 ; n6833
g6770 nor n6545 n6546 ; n6834
g6771 nor n6833 n6834 ; n6835
g6772 nor n6832 n6835 ; n6836
g6773 nor n6546 n6836 ; n6837
g6774 nor n6500 n6837 ; n6838
g6775 and n6500 n6837 ; n6839
g6776 nor n6838 n6839 ; n6840
g6777 and n1992_not n3457 ; n6841
g6778 and n2152_not n3542 ; n6842
g6779 and n2057_not n3606 ; n6843
g6780 nor n6842 n6843 ; n6844
g6781 and n6841_not n6844 ; n6845
g6782 and n3368_not n6845 ; n6846
g6783 and n6143_not n6845 ; n6847
g6784 nor n6846 n6847 ; n6848
g6785 and a[29] n6848_not ; n6849
g6786 and a[29]_not n6848 ; n6850
g6787 nor n6849 n6850 ; n6851
g6788 and n6840 n6851_not ; n6852
g6789 nor n6838 n6852 ; n6853
g6790 nor n6487 n6497 ; n6854
g6791 nor n6496 n6497 ; n6855
g6792 nor n6854 n6855 ; n6856
g6793 nor n6853 n6856 ; n6857
g6794 nor n6497 n6857 ; n6858
g6795 nor n6474 n6484 ; n6859
g6796 nor n6483 n6484 ; n6860
g6797 nor n6859 n6860 ; n6861
g6798 nor n6858 n6861 ; n6862
g6799 nor n6484 n6862 ; n6863
g6800 nor n6471 n6863 ; n6864
g6801 and n6471 n6863 ; n6865
g6802 nor n6864 n6865 ; n6866
g6803 and n1779_not n3457 ; n6867
g6804 and n1913_not n3542 ; n6868
g6805 and n1877_not n3606 ; n6869
g6806 nor n6868 n6869 ; n6870
g6807 and n6867_not n6870 ; n6871
g6808 and n3368 n5851 ; n6872
g6809 and n6871 n6872_not ; n6873
g6810 and a[29] n6873_not ; n6874
g6811 and a[29] n6874_not ; n6875
g6812 nor n6873 n6874 ; n6876
g6813 nor n6875 n6876 ; n6877
g6814 and n6866 n6877_not ; n6878
g6815 nor n6864 n6878 ; n6879
g6816 and n6157_not n6168 ; n6880
g6817 nor n6169 n6880 ; n6881
g6818 and n6879_not n6881 ; n6882
g6819 and n6879 n6881_not ; n6883
g6820 nor n6882 n6883 ; n6884
g6821 and n1364_not n3884 ; n6885
g6822 and n1572_not n3967 ; n6886
g6823 and n1472_not n4046 ; n6887
g6824 nor n6886 n6887 ; n6888
g6825 and n6885_not n6888 ; n6889
g6826 and n4050 n5114 ; n6890
g6827 and n6889 n6890_not ; n6891
g6828 and a[26] n6891_not ; n6892
g6829 and a[26] n6892_not ; n6893
g6830 nor n6891 n6892 ; n6894
g6831 nor n6893 n6894 ; n6895
g6832 and n6884 n6895_not ; n6896
g6833 nor n6882 n6896 ; n6897
g6834 nor n6468 n6897 ; n6898
g6835 and n6468 n6897 ; n6899
g6836 nor n6898 n6899 ; n6900
g6837 and n958_not n4694 ; n6901
g6838 and n1178_not n4533 ; n6902
g6839 and n1060_not n4604 ; n6903
g6840 nor n6902 n6903 ; n6904
g6841 and n6901_not n6904 ; n6905
g6842 and n4536 n4633 ; n6906
g6843 and n6905 n6906_not ; n6907
g6844 and a[23] n6907_not ; n6908
g6845 and a[23] n6908_not ; n6909
g6846 nor n6907 n6908 ; n6910
g6847 nor n6909 n6910 ; n6911
g6848 and n6900 n6911_not ; n6912
g6849 nor n6898 n6912 ; n6913
g6850 nor n6465 n6913 ; n6914
g6851 nor n6462 n6914 ; n6915
g6852 nor n6448 n6915 ; n6916
g6853 and n6448 n6915 ; n6917
g6854 nor n6916 n6917 ; n6918
g6855 and n3012_not n5496 ; n6919
g6856 and n587_not n4935 ; n6920
g6857 and n392_not n5407 ; n6921
g6858 nor n6920 n6921 ; n6922
g6859 and n6919_not n6922 ; n6923
g6860 and n3018 n4938 ; n6924
g6861 and n6923 n6924_not ; n6925
g6862 and a[20] n6925_not ; n6926
g6863 and a[20] n6926_not ; n6927
g6864 nor n6925 n6926 ; n6928
g6865 nor n6927 n6928 ; n6929
g6866 and n6918 n6929_not ; n6930
g6867 nor n6916 n6930 ; n6931
g6868 nor n6445 n6931 ; n6932
g6869 and n6445 n6931 ; n6933
g6870 nor n6932 n6933 ; n6934
g6871 and n3805_not n6233 ; n6935
g6872 and n3605_not n5663 ; n6936
g6873 and n3456_not n5939 ; n6937
g6874 nor n6936 n6937 ; n6938
g6875 and n6935_not n6938 ; n6939
g6876 and n3818 n5666 ; n6940
g6877 and n6939 n6940_not ; n6941
g6878 and a[17] n6941_not ; n6942
g6879 and a[17] n6942_not ; n6943
g6880 nor n6941 n6942 ; n6944
g6881 nor n6943 n6944 ; n6945
g6882 and n6934 n6945_not ; n6946
g6883 nor n6932 n6946 ; n6947
g6884 nor n6442 n6947 ; n6948
g6885 nor n6439 n6948 ; n6949
g6886 and n3877_not n6402 ; n6950
g6887 and n6393 n6400_not ; n6951
g6888 and n4515_not n6951 ; n6952
g6889 nor n6950 n6952 ; n6953
g6890 and n6397_not n6953 ; n6954
g6891 and n4609_not n6953 ; n6955
g6892 nor n6954 n6955 ; n6956
g6893 and a[14] n6956_not ; n6957
g6894 and a[14]_not n6956 ; n6958
g6895 nor n6957 n6958 ; n6959
g6896 nor n6949 n6959 ; n6960
g6897 and n6377 n6389_not ; n6961
g6898 nor n6388 n6389 ; n6962
g6899 nor n6961 n6962 ; n6963
g6900 and n6949 n6959 ; n6964
g6901 nor n6960 n6964 ; n6965
g6902 and n6963_not n6965 ; n6966
g6903 nor n6960 n6966 ; n6967
g6904 nor n6425 n6967 ; n6968
g6905 and n6425 n6967 ; n6969
g6906 nor n6968 n6969 ; n6970
g6907 and n6934 n6946_not ; n6971
g6908 nor n6945 n6946 ; n6972
g6909 nor n6971 n6972 ; n6973
g6910 and n6918 n6930_not ; n6974
g6911 nor n6929 n6930 ; n6975
g6912 nor n6974 n6975 ; n6976
g6913 and n6465 n6913 ; n6977
g6914 nor n6914 n6977 ; n6978
g6915 and n392_not n5496 ; n6979
g6916 and n710_not n4935 ; n6980
g6917 and n587_not n5407 ; n6981
g6918 nor n6980 n6981 ; n6982
g6919 and n6979_not n6982 ; n6983
g6920 and n4938_not n6983 ; n6984
g6921 and n3347_not n6983 ; n6985
g6922 nor n6984 n6985 ; n6986
g6923 and a[20] n6986_not ; n6987
g6924 and a[20]_not n6986 ; n6988
g6925 nor n6987 n6988 ; n6989
g6926 and n6978 n6989_not ; n6990
g6927 and n6900 n6912_not ; n6991
g6928 nor n6911 n6912 ; n6992
g6929 nor n6991 n6992 ; n6993
g6930 and n6884 n6896_not ; n6994
g6931 nor n6895 n6896 ; n6995
g6932 nor n6994 n6995 ; n6996
g6933 and n6866 n6878_not ; n6997
g6934 nor n6877 n6878 ; n6998
g6935 nor n6997 n6998 ; n6999
g6936 and n1472_not n3884 ; n7000
g6937 and n1665_not n3967 ; n7001
g6938 and n1572_not n4046 ; n7002
g6939 nor n7001 n7002 ; n7003
g6940 and n7000_not n7003 ; n7004
g6941 and n4050_not n7004 ; n7005
g6942 and n5139_not n7004 ; n7006
g6943 nor n7005 n7006 ; n7007
g6944 and a[26] n7007_not ; n7008
g6945 and a[26]_not n7007 ; n7009
g6946 nor n7008 n7009 ; n7010
g6947 nor n6999 n7010 ; n7011
g6948 nor n6858 n6862 ; n7012
g6949 nor n6861 n6862 ; n7013
g6950 nor n7012 n7013 ; n7014
g6951 and n1877_not n3457 ; n7015
g6952 and n1992_not n3542 ; n7016
g6953 and n1913_not n3606 ; n7017
g6954 nor n7016 n7017 ; n7018
g6955 and n7015_not n7018 ; n7019
g6956 and n3368_not n7019 ; n7020
g6957 and n6007_not n7019 ; n7021
g6958 nor n7020 n7021 ; n7022
g6959 and a[29] n7022_not ; n7023
g6960 and a[29]_not n7022 ; n7024
g6961 nor n7023 n7024 ; n7025
g6962 nor n7014 n7025 ; n7026
g6963 and n7014 n7025 ; n7027
g6964 nor n7026 n7027 ; n7028
g6965 and n1572_not n3884 ; n7029
g6966 and n1779_not n3967 ; n7030
g6967 and n1665_not n4046 ; n7031
g6968 nor n7030 n7031 ; n7032
g6969 and n7029_not n7032 ; n7033
g6970 and n4050 n5561 ; n7034
g6971 and n7033 n7034_not ; n7035
g6972 and a[26] n7035_not ; n7036
g6973 and a[26] n7036_not ; n7037
g6974 nor n7035 n7036 ; n7038
g6975 nor n7037 n7038 ; n7039
g6976 and n7028 n7039_not ; n7040
g6977 nor n7026 n7040 ; n7041
g6978 and n6999 n7010 ; n7042
g6979 nor n7011 n7042 ; n7043
g6980 and n7041_not n7043 ; n7044
g6981 nor n7011 n7044 ; n7045
g6982 nor n6996 n7045 ; n7046
g6983 and n6996 n7045 ; n7047
g6984 nor n7046 n7047 ; n7048
g6985 and n1060_not n4694 ; n7049
g6986 and n1235_not n4533 ; n7050
g6987 and n1178_not n4604 ; n7051
g6988 nor n7050 n7051 ; n7052
g6989 and n7049_not n7052 ; n7053
g6990 and n4429 n4536 ; n7054
g6991 and n7053 n7054_not ; n7055
g6992 and a[23] n7055_not ; n7056
g6993 and a[23] n7056_not ; n7057
g6994 nor n7055 n7056 ; n7058
g6995 nor n7057 n7058 ; n7059
g6996 and n7048 n7059_not ; n7060
g6997 nor n7046 n7060 ; n7061
g6998 nor n6993 n7061 ; n7062
g6999 and n6993 n7061 ; n7063
g7000 nor n7062 n7063 ; n7064
g7001 and n587_not n5496 ; n7065
g7002 and n867_not n4935 ; n7066
g7003 and n710_not n5407 ; n7067
g7004 nor n7066 n7067 ; n7068
g7005 and n7065_not n7068 ; n7069
g7006 and n3331 n4938 ; n7070
g7007 and n7069 n7070_not ; n7071
g7008 and a[20] n7071_not ; n7072
g7009 and a[20] n7072_not ; n7073
g7010 nor n7071 n7072 ; n7074
g7011 nor n7073 n7074 ; n7075
g7012 and n7064 n7075_not ; n7076
g7013 nor n7062 n7076 ; n7077
g7014 and n6978_not n6989 ; n7078
g7015 nor n6990 n7078 ; n7079
g7016 and n7077_not n7079 ; n7080
g7017 nor n6990 n7080 ; n7081
g7018 nor n6976 n7081 ; n7082
g7019 and n6976 n7081 ; n7083
g7020 nor n7082 n7083 ; n7084
g7021 and n3456_not n6233 ; n7085
g7022 and n3539_not n5663 ; n7086
g7023 and n3605_not n5939 ; n7087
g7024 nor n7086 n7087 ; n7088
g7025 and n7085_not n7088 ; n7089
g7026 and n3627 n5666 ; n7090
g7027 and n7089 n7090_not ; n7091
g7028 and a[17] n7091_not ; n7092
g7029 and a[17] n7092_not ; n7093
g7030 nor n7091 n7092 ; n7094
g7031 nor n7093 n7094 ; n7095
g7032 and n7084 n7095_not ; n7096
g7033 nor n7082 n7096 ; n7097
g7034 nor n6973 n7097 ; n7098
g7035 and n6973 n7097 ; n7099
g7036 nor n7098 n7099 ; n7100
g7037 and n6393_not n6396 ; n7101
g7038 and n3877_not n7101 ; n7102
g7039 and n3964_not n6402 ; n7103
g7040 and n4045_not n6951 ; n7104
g7041 nor n7103 n7104 ; n7105
g7042 and n7102_not n7105 ; n7106
g7043 and n4067 n6397 ; n7107
g7044 and n7106 n7107_not ; n7108
g7045 and a[14] n7108_not ; n7109
g7046 and a[14] n7109_not ; n7110
g7047 nor n7108 n7109 ; n7111
g7048 nor n7110 n7111 ; n7112
g7049 and n7100 n7112_not ; n7113
g7050 nor n7098 n7113 ; n7114
g7051 and n4515_not n7101 ; n7115
g7052 and n4045_not n6402 ; n7116
g7053 and n3877_not n6951 ; n7117
g7054 nor n7116 n7117 ; n7118
g7055 and n7115_not n7118 ; n7119
g7056 and n6397_not n7119 ; n7120
g7057 and n4715_not n7119 ; n7121
g7058 nor n7120 n7121 ; n7122
g7059 and a[14] n7122_not ; n7123
g7060 and a[14]_not n7122 ; n7124
g7061 nor n7123 n7124 ; n7125
g7062 nor n7114 n7125 ; n7126
g7063 and n6442 n6947 ; n7127
g7064 nor n6948 n7127 ; n7128
g7065 nor n7114 n7126 ; n7129
g7066 nor n7125 n7126 ; n7130
g7067 nor n7129 n7130 ; n7131
g7068 and n7128 n7131_not ; n7132
g7069 nor n7126 n7132 ; n7133
g7070 and n6963 n6965_not ; n7134
g7071 nor n6966 n7134 ; n7135
g7072 and n7133_not n7135 ; n7136
g7073 and n7084 n7096_not ; n7137
g7074 nor n7095 n7096 ; n7138
g7075 nor n7137 n7138 ; n7139
g7076 and n3605_not n6233 ; n7140
g7077 and n3012_not n5663 ; n7141
g7078 and n3539_not n5939 ; n7142
g7079 nor n7141 n7142 ; n7143
g7080 and n7140_not n7143 ; n7144
g7081 and n4084 n5666 ; n7145
g7082 and n7144 n7145_not ; n7146
g7083 and a[17] n7146_not ; n7147
g7084 nor n7146 n7147 ; n7148
g7085 and a[17] n7147_not ; n7149
g7086 nor n7148 n7149 ; n7150
g7087 and n7077 n7079_not ; n7151
g7088 nor n7080 n7151 ; n7152
g7089 and n7150_not n7152 ; n7153
g7090 nor n7150 n7153 ; n7154
g7091 and n7152 n7153_not ; n7155
g7092 nor n7154 n7155 ; n7156
g7093 and n7064 n7076_not ; n7157
g7094 nor n7075 n7076 ; n7158
g7095 nor n7157 n7158 ; n7159
g7096 and n7048 n7060_not ; n7160
g7097 nor n7059 n7060 ; n7161
g7098 nor n7160 n7161 ; n7162
g7099 and n1178_not n4694 ; n7163
g7100 and n1364_not n4533 ; n7164
g7101 and n1235_not n4604 ; n7165
g7102 nor n7164 n7165 ; n7166
g7103 and n7163_not n7166 ; n7167
g7104 and n4536 n4861 ; n7168
g7105 and n7167 n7168_not ; n7169
g7106 and a[23] n7169_not ; n7170
g7107 nor n7169 n7170 ; n7171
g7108 and a[23] n7170_not ; n7172
g7109 nor n7171 n7172 ; n7173
g7110 and n7041 n7043_not ; n7174
g7111 nor n7044 n7174 ; n7175
g7112 and n7173_not n7175 ; n7176
g7113 nor n7173 n7176 ; n7177
g7114 and n7175 n7176_not ; n7178
g7115 nor n7177 n7178 ; n7179
g7116 and n7028 n7040_not ; n7180
g7117 nor n7039 n7040 ; n7181
g7118 nor n7180 n7181 ; n7182
g7119 nor n6853 n6857 ; n7183
g7120 nor n6856 n6857 ; n7184
g7121 nor n7183 n7184 ; n7185
g7122 and n1913_not n3457 ; n7186
g7123 and n2057_not n3542 ; n7187
g7124 and n1992_not n3606 ; n7188
g7125 nor n7187 n7188 ; n7189
g7126 and n7186_not n7189 ; n7190
g7127 and n3368_not n7190 ; n7191
g7128 and n5834_not n7190 ; n7192
g7129 nor n7191 n7192 ; n7193
g7130 and a[29] n7193_not ; n7194
g7131 and a[29]_not n7193 ; n7195
g7132 nor n7194 n7195 ; n7196
g7133 nor n7185 n7196 ; n7197
g7134 and n7185 n7196 ; n7198
g7135 nor n7197 n7198 ; n7199
g7136 and n1665_not n3884 ; n7200
g7137 and n1877_not n3967 ; n7201
g7138 and n1779_not n4046 ; n7202
g7139 nor n7201 n7202 ; n7203
g7140 and n7200_not n7203 ; n7204
g7141 and n4050 n5328 ; n7205
g7142 and n7204 n7205_not ; n7206
g7143 and a[26] n7206_not ; n7207
g7144 and a[26] n7207_not ; n7208
g7145 nor n7206 n7207 ; n7209
g7146 nor n7208 n7209 ; n7210
g7147 and n7199 n7210_not ; n7211
g7148 nor n7197 n7211 ; n7212
g7149 nor n7182 n7212 ; n7213
g7150 and n7182 n7212 ; n7214
g7151 nor n7213 n7214 ; n7215
g7152 and n1235_not n4694 ; n7216
g7153 and n1472_not n4533 ; n7217
g7154 and n1364_not n4604 ; n7218
g7155 nor n7217 n7218 ; n7219
g7156 and n7216_not n7219 ; n7220
g7157 and n4536 n4848 ; n7221
g7158 and n7220 n7221_not ; n7222
g7159 and a[23] n7222_not ; n7223
g7160 and a[23] n7223_not ; n7224
g7161 nor n7222 n7223 ; n7225
g7162 nor n7224 n7225 ; n7226
g7163 and n7215 n7226_not ; n7227
g7164 nor n7213 n7227 ; n7228
g7165 nor n7179 n7228 ; n7229
g7166 nor n7176 n7229 ; n7230
g7167 nor n7162 n7230 ; n7231
g7168 and n7162 n7230 ; n7232
g7169 nor n7231 n7232 ; n7233
g7170 and n710_not n5496 ; n7234
g7171 and n958_not n4935 ; n7235
g7172 and n867_not n5407 ; n7236
g7173 nor n7235 n7236 ; n7237
g7174 and n7234_not n7237 ; n7238
g7175 and n4179 n4938 ; n7239
g7176 and n7238 n7239_not ; n7240
g7177 and a[20] n7240_not ; n7241
g7178 and a[20] n7241_not ; n7242
g7179 nor n7240 n7241 ; n7243
g7180 nor n7242 n7243 ; n7244
g7181 and n7233 n7244_not ; n7245
g7182 nor n7231 n7245 ; n7246
g7183 nor n7159 n7246 ; n7247
g7184 and n7159 n7246 ; n7248
g7185 nor n7247 n7248 ; n7249
g7186 and n3539_not n6233 ; n7250
g7187 and n392_not n5663 ; n7251
g7188 and n3012_not n5939 ; n7252
g7189 nor n7251 n7252 ; n7253
g7190 and n7250_not n7253 ; n7254
g7191 and n3715 n5666 ; n7255
g7192 and n7254 n7255_not ; n7256
g7193 and a[17] n7256_not ; n7257
g7194 and a[17] n7257_not ; n7258
g7195 nor n7256 n7257 ; n7259
g7196 nor n7258 n7259 ; n7260
g7197 and n7249 n7260_not ; n7261
g7198 nor n7247 n7261 ; n7262
g7199 nor n7156 n7262 ; n7263
g7200 nor n7153 n7263 ; n7264
g7201 nor n7139 n7264 ; n7265
g7202 and n7139 n7264 ; n7266
g7203 nor n7265 n7266 ; n7267
g7204 and n4045_not n7101 ; n7268
g7205 and n3805_not n6402 ; n7269
g7206 and n3964_not n6951 ; n7270
g7207 nor n7269 n7270 ; n7271
g7208 and n7268_not n7271 ; n7272
g7209 and n4477 n6397 ; n7273
g7210 and n7272 n7273_not ; n7274
g7211 and a[14] n7274_not ; n7275
g7212 and a[14] n7275_not ; n7276
g7213 nor n7274 n7275 ; n7277
g7214 nor n7276 n7277 ; n7278
g7215 and n7267 n7278_not ; n7279
g7216 nor n7265 n7279 ; n7280
g7217 and a[9]_not a[10] ; n7281
g7218 and a[9] a[10]_not ; n7282
g7219 nor n7281 n7282 ; n7283
g7220 and a[10] a[11]_not ; n7284
g7221 and a[10]_not a[11] ; n7285
g7222 nor n7284 n7285 ; n7286
g7223 and a[8] a[9]_not ; n7287
g7224 and a[8]_not a[9] ; n7288
g7225 nor n7287 n7288 ; n7289
g7226 and n7286_not n7289 ; n7290
g7227 and n7283 n7290 ; n7291
g7228 and n4515_not n7291 ; n7292
g7229 nor n4522 n7292 ; n7293
g7230 nor n7286 n7289 ; n7294
g7231 nor n7292 n7294 ; n7295
g7232 nor n7293 n7295 ; n7296
g7233 and a[11] n7296_not ; n7297
g7234 and a[11]_not n7296 ; n7298
g7235 nor n7297 n7298 ; n7299
g7236 nor n7280 n7299 ; n7300
g7237 and n7100 n7113_not ; n7301
g7238 nor n7112 n7113 ; n7302
g7239 nor n7301 n7302 ; n7303
g7240 and n7280 n7299 ; n7304
g7241 nor n7300 n7304 ; n7305
g7242 and n7303_not n7305 ; n7306
g7243 nor n7300 n7306 ; n7307
g7244 nor n7128 n7130 ; n7308
g7245 and n7129_not n7308 ; n7309
g7246 nor n7132 n7309 ; n7310
g7247 and n7307_not n7310 ; n7311
g7248 nor n7303 n7306 ; n7312
g7249 and n7305 n7306_not ; n7313
g7250 nor n7312 n7313 ; n7314
g7251 and n7156 n7262 ; n7315
g7252 nor n7263 n7315 ; n7316
g7253 and n3964_not n7101 ; n7317
g7254 and n3456_not n6402 ; n7318
g7255 and n3805_not n6951 ; n7319
g7256 nor n7318 n7319 ; n7320
g7257 and n7317_not n7320 ; n7321
g7258 and n6397_not n7321 ; n7322
g7259 and n4558_not n7321 ; n7323
g7260 nor n7322 n7323 ; n7324
g7261 and a[14] n7324_not ; n7325
g7262 and a[14]_not n7324 ; n7326
g7263 nor n7325 n7326 ; n7327
g7264 and n7316 n7327_not ; n7328
g7265 and n7249 n7261_not ; n7329
g7266 nor n7260 n7261 ; n7330
g7267 nor n7329 n7330 ; n7331
g7268 and n7233 n7245_not ; n7332
g7269 nor n7244 n7245 ; n7333
g7270 nor n7332 n7333 ; n7334
g7271 and n7179 n7228 ; n7335
g7272 nor n7229 n7335 ; n7336
g7273 and n867_not n5496 ; n7337
g7274 and n1060_not n4935 ; n7338
g7275 and n958_not n5407 ; n7339
g7276 nor n7338 n7339 ; n7340
g7277 and n7337_not n7340 ; n7341
g7278 and n4938_not n7341 ; n7342
g7279 and n4204_not n7341 ; n7343
g7280 nor n7342 n7343 ; n7344
g7281 and a[20] n7344_not ; n7345
g7282 and a[20]_not n7344 ; n7346
g7283 nor n7345 n7346 ; n7347
g7284 and n7336 n7347_not ; n7348
g7285 and n7215 n7227_not ; n7349
g7286 nor n7226 n7227 ; n7350
g7287 nor n7349 n7350 ; n7351
g7288 and n7199 n7211_not ; n7352
g7289 nor n7210 n7211 ; n7353
g7290 nor n7352 n7353 ; n7354
g7291 nor n6832 n6836 ; n7355
g7292 nor n6835 n6836 ; n7356
g7293 nor n7355 n7356 ; n7357
g7294 and n2057_not n3457 ; n7358
g7295 and n2189_not n3542 ; n7359
g7296 and n2152_not n3606 ; n7360
g7297 nor n7359 n7360 ; n7361
g7298 and n7358_not n7361 ; n7362
g7299 and n3368_not n7362 ; n7363
g7300 and n6479_not n7362 ; n7364
g7301 nor n7363 n7364 ; n7365
g7302 and a[29] n7365_not ; n7366
g7303 and a[29]_not n7365 ; n7367
g7304 nor n7366 n7367 ; n7368
g7305 nor n7357 n7368 ; n7369
g7306 nor n6827 n6831 ; n7370
g7307 nor n6830 n6831 ; n7371
g7308 nor n7370 n7371 ; n7372
g7309 and n2152_not n3457 ; n7373
g7310 and n2291_not n3542 ; n7374
g7311 and n2189_not n3606 ; n7375
g7312 nor n7374 n7375 ; n7376
g7313 and n7373_not n7376 ; n7377
g7314 and n3368_not n7377 ; n7378
g7315 and n6492_not n7377 ; n7379
g7316 nor n7378 n7379 ; n7380
g7317 and a[29] n7380_not ; n7381
g7318 and a[29]_not n7380 ; n7382
g7319 nor n7381 n7382 ; n7383
g7320 nor n7372 n7383 ; n7384
g7321 and n2189_not n3457 ; n7385
g7322 and n2388_not n3542 ; n7386
g7323 and n2291_not n3606 ; n7387
g7324 nor n7386 n7387 ; n7388
g7325 and n7385_not n7388 ; n7389
g7326 and n3368 n6122 ; n7390
g7327 and n7389 n7390_not ; n7391
g7328 and a[29] n7391_not ; n7392
g7329 nor n7391 n7392 ; n7393
g7330 and a[29] n7392_not ; n7394
g7331 nor n7393 n7394 ; n7395
g7332 nor n6822 n6826 ; n7396
g7333 nor n6825 n6826 ; n7397
g7334 nor n7396 n7397 ; n7398
g7335 nor n7395 n7398 ; n7399
g7336 nor n7395 n7399 ; n7400
g7337 nor n7398 n7399 ; n7401
g7338 nor n7400 n7401 ; n7402
g7339 and n2291_not n3457 ; n7403
g7340 and n2464_not n3542 ; n7404
g7341 and n2388_not n3606 ; n7405
g7342 nor n7404 n7405 ; n7406
g7343 and n7403_not n7406 ; n7407
g7344 and n3368 n6541 ; n7408
g7345 and n7407 n7408_not ; n7409
g7346 and a[29] n7409_not ; n7410
g7347 nor n7409 n7410 ; n7411
g7348 and a[29] n7410_not ; n7412
g7349 nor n7411 n7412 ; n7413
g7350 nor n6817 n6821 ; n7414
g7351 nor n6820 n6821 ; n7415
g7352 nor n7414 n7415 ; n7416
g7353 nor n7413 n7416 ; n7417
g7354 nor n7413 n7417 ; n7418
g7355 nor n7416 n7417 ; n7419
g7356 nor n7418 n7419 ; n7420
g7357 and n2388_not n3457 ; n7421
g7358 and n2533_not n3542 ; n7422
g7359 and n2464_not n3606 ; n7423
g7360 nor n7422 n7423 ; n7424
g7361 and n7421_not n7424 ; n7425
g7362 and n3368 n6591 ; n7426
g7363 and n7425 n7426_not ; n7427
g7364 and a[29] n7427_not ; n7428
g7365 nor n7427 n7428 ; n7429
g7366 and a[29] n7428_not ; n7430
g7367 nor n7429 n7430 ; n7431
g7368 nor n6813 n6816 ; n7432
g7369 and n6815 n6816_not ; n7433
g7370 nor n7432 n7433 ; n7434
g7371 nor n7431 n7434 ; n7435
g7372 nor n7431 n7435 ; n7436
g7373 nor n7434 n7435 ; n7437
g7374 nor n7436 n7437 ; n7438
g7375 and n2464_not n3457 ; n7439
g7376 and n2571_not n3542 ; n7440
g7377 and n2533_not n3606 ; n7441
g7378 nor n7440 n7441 ; n7442
g7379 and n7439_not n7442 ; n7443
g7380 and n3368 n6646 ; n7444
g7381 and n7443 n7444_not ; n7445
g7382 and a[29] n7445_not ; n7446
g7383 nor n7445 n7446 ; n7447
g7384 and a[29] n7446_not ; n7448
g7385 nor n7447 n7448 ; n7449
g7386 nor n6791 n6803 ; n7450
g7387 nor n6802 n6803 ; n7451
g7388 nor n7450 n7451 ; n7452
g7389 nor n7449 n7452 ; n7453
g7390 nor n7449 n7453 ; n7454
g7391 nor n7452 n7453 ; n7455
g7392 nor n7454 n7455 ; n7456
g7393 and n2533_not n3457 ; n7457
g7394 and n2674_not n3542 ; n7458
g7395 and n2571_not n3606 ; n7459
g7396 nor n7458 n7459 ; n7460
g7397 and n7457_not n7460 ; n7461
g7398 and n3368 n6695 ; n7462
g7399 and n7461 n7462_not ; n7463
g7400 and a[29] n7463_not ; n7464
g7401 nor n7463 n7464 ; n7465
g7402 and a[29] n7464_not ; n7466
g7403 nor n7465 n7466 ; n7467
g7404 and n2736 n2829_not ; n7468
g7405 nor n6795 n7468 ; n7469
g7406 and n75 n7469_not ; n7470
g7407 and n2829_not n3028 ; n7471
g7408 and n2736_not n3020 ; n7472
g7409 nor n7471 n7472 ; n7473
g7410 and n7470_not n7473 ; n7474
g7411 nor n7467 n7474 ; n7475
g7412 nor n7467 n7475 ; n7476
g7413 nor n7474 n7475 ; n7477
g7414 nor n7476 n7477 ; n7478
g7415 nor n75 n3020 ; n7479
g7416 nor n2829 n7479 ; n7480
g7417 and n2829_not n3606 ; n7481
g7418 and n2736_not n3457 ; n7482
g7419 nor n7481 n7482 ; n7483
g7420 and n3368 n7469_not ; n7484
g7421 and n7483 n7484_not ; n7485
g7422 and a[29] n7485_not ; n7486
g7423 and a[29] n7486_not ; n7487
g7424 nor n7485 n7486 ; n7488
g7425 nor n7487 n7488 ; n7489
g7426 nor n2829 n3367 ; n7490
g7427 and a[29] n7490_not ; n7491
g7428 and n7489_not n7491 ; n7492
g7429 and n2674_not n3457 ; n7493
g7430 and n2829_not n3542 ; n7494
g7431 and n2736_not n3606 ; n7495
g7432 nor n7494 n7495 ; n7496
g7433 and n7493_not n7496 ; n7497
g7434 and n3368_not n7497 ; n7498
g7435 and n6798_not n7497 ; n7499
g7436 nor n7498 n7499 ; n7500
g7437 and a[29] n7500_not ; n7501
g7438 and a[29]_not n7500 ; n7502
g7439 nor n7501 n7502 ; n7503
g7440 and n7492 n7503_not ; n7504
g7441 and n7480 n7504 ; n7505
g7442 and n2571_not n3457 ; n7506
g7443 and n2736_not n3542 ; n7507
g7444 and n2674_not n3606 ; n7508
g7445 nor n7507 n7508 ; n7509
g7446 and n7506_not n7509 ; n7510
g7447 and n3368 n6806 ; n7511
g7448 and n7510 n7511_not ; n7512
g7449 and a[29] n7512_not ; n7513
g7450 nor n7512 n7513 ; n7514
g7451 and a[29] n7513_not ; n7515
g7452 nor n7514 n7515 ; n7516
g7453 and n7480_not n7504 ; n7517
g7454 and n7480 n7504_not ; n7518
g7455 nor n7517 n7518 ; n7519
g7456 nor n7516 n7519 ; n7520
g7457 nor n7505 n7520 ; n7521
g7458 nor n7478 n7521 ; n7522
g7459 nor n7475 n7522 ; n7523
g7460 nor n7456 n7523 ; n7524
g7461 nor n7453 n7524 ; n7525
g7462 nor n7438 n7525 ; n7526
g7463 nor n7435 n7526 ; n7527
g7464 nor n7420 n7527 ; n7528
g7465 nor n7417 n7528 ; n7529
g7466 nor n7402 n7529 ; n7530
g7467 nor n7399 n7530 ; n7531
g7468 and n7372 n7383 ; n7532
g7469 nor n7384 n7532 ; n7533
g7470 and n7531_not n7533 ; n7534
g7471 nor n7384 n7534 ; n7535
g7472 and n7357 n7368 ; n7536
g7473 nor n7369 n7536 ; n7537
g7474 and n7535_not n7537 ; n7538
g7475 nor n7369 n7538 ; n7539
g7476 and n6840_not n6851 ; n7540
g7477 nor n6852 n7540 ; n7541
g7478 and n7539_not n7541 ; n7542
g7479 and n1779_not n3884 ; n7543
g7480 and n1913_not n3967 ; n7544
g7481 and n1877_not n4046 ; n7545
g7482 nor n7544 n7545 ; n7546
g7483 and n7543_not n7546 ; n7547
g7484 and n4050 n5851 ; n7548
g7485 and n7547 n7548_not ; n7549
g7486 and a[26] n7549_not ; n7550
g7487 nor n7549 n7550 ; n7551
g7488 and a[26] n7550_not ; n7552
g7489 nor n7551 n7552 ; n7553
g7490 and n7539 n7541_not ; n7554
g7491 nor n7542 n7554 ; n7555
g7492 and n7553_not n7555 ; n7556
g7493 nor n7542 n7556 ; n7557
g7494 nor n7354 n7557 ; n7558
g7495 and n7354 n7557 ; n7559
g7496 nor n7558 n7559 ; n7560
g7497 and n1364_not n4694 ; n7561
g7498 and n1572_not n4533 ; n7562
g7499 and n1472_not n4604 ; n7563
g7500 nor n7562 n7563 ; n7564
g7501 and n7561_not n7564 ; n7565
g7502 and n4536 n5114 ; n7566
g7503 and n7565 n7566_not ; n7567
g7504 and a[23] n7567_not ; n7568
g7505 and a[23] n7568_not ; n7569
g7506 nor n7567 n7568 ; n7570
g7507 nor n7569 n7570 ; n7571
g7508 and n7560 n7571_not ; n7572
g7509 nor n7558 n7572 ; n7573
g7510 nor n7351 n7573 ; n7574
g7511 and n7351 n7573 ; n7575
g7512 nor n7574 n7575 ; n7576
g7513 and n958_not n5496 ; n7577
g7514 and n1178_not n4935 ; n7578
g7515 and n1060_not n5407 ; n7579
g7516 nor n7578 n7579 ; n7580
g7517 and n7577_not n7580 ; n7581
g7518 and n4633 n4938 ; n7582
g7519 and n7581 n7582_not ; n7583
g7520 and a[20] n7583_not ; n7584
g7521 and a[20] n7584_not ; n7585
g7522 nor n7583 n7584 ; n7586
g7523 nor n7585 n7586 ; n7587
g7524 and n7576 n7587_not ; n7588
g7525 nor n7574 n7588 ; n7589
g7526 and n7336_not n7347 ; n7590
g7527 nor n7348 n7590 ; n7591
g7528 and n7589_not n7591 ; n7592
g7529 nor n7348 n7592 ; n7593
g7530 nor n7334 n7593 ; n7594
g7531 and n7334 n7593 ; n7595
g7532 nor n7594 n7595 ; n7596
g7533 and n3012_not n6233 ; n7597
g7534 and n587_not n5663 ; n7598
g7535 and n392_not n5939 ; n7599
g7536 nor n7598 n7599 ; n7600
g7537 and n7597_not n7600 ; n7601
g7538 and n3018 n5666 ; n7602
g7539 and n7601 n7602_not ; n7603
g7540 and a[17] n7603_not ; n7604
g7541 and a[17] n7604_not ; n7605
g7542 nor n7603 n7604 ; n7606
g7543 nor n7605 n7606 ; n7607
g7544 and n7596 n7607_not ; n7608
g7545 nor n7594 n7608 ; n7609
g7546 nor n7331 n7609 ; n7610
g7547 and n7331 n7609 ; n7611
g7548 nor n7610 n7611 ; n7612
g7549 and n3805_not n7101 ; n7613
g7550 and n3605_not n6402 ; n7614
g7551 and n3456_not n6951 ; n7615
g7552 nor n7614 n7615 ; n7616
g7553 and n7613_not n7616 ; n7617
g7554 and n3818 n6397 ; n7618
g7555 and n7617 n7618_not ; n7619
g7556 and a[14] n7619_not ; n7620
g7557 and a[14] n7620_not ; n7621
g7558 nor n7619 n7620 ; n7622
g7559 nor n7621 n7622 ; n7623
g7560 and n7612 n7623_not ; n7624
g7561 nor n7610 n7624 ; n7625
g7562 and n7316 n7328_not ; n7626
g7563 nor n7327 n7328 ; n7627
g7564 nor n7626 n7627 ; n7628
g7565 nor n7625 n7628 ; n7629
g7566 nor n7328 n7629 ; n7630
g7567 and n3877_not n7291 ; n7631
g7568 and n7283_not n7289 ; n7632
g7569 and n4515_not n7632 ; n7633
g7570 nor n7631 n7633 ; n7634
g7571 and n7294_not n7634 ; n7635
g7572 and n4609_not n7634 ; n7636
g7573 nor n7635 n7636 ; n7637
g7574 and a[11] n7637_not ; n7638
g7575 and a[11]_not n7637 ; n7639
g7576 nor n7638 n7639 ; n7640
g7577 nor n7630 n7640 ; n7641
g7578 and n7267 n7279_not ; n7642
g7579 nor n7278 n7279 ; n7643
g7580 nor n7642 n7643 ; n7644
g7581 and n7630 n7640 ; n7645
g7582 nor n7641 n7645 ; n7646
g7583 and n7644_not n7646 ; n7647
g7584 nor n7641 n7647 ; n7648
g7585 nor n7314 n7648 ; n7649
g7586 and n7314 n7648 ; n7650
g7587 nor n7649 n7650 ; n7651
g7588 and n7612 n7624_not ; n7652
g7589 nor n7623 n7624 ; n7653
g7590 nor n7652 n7653 ; n7654
g7591 and n7596 n7608_not ; n7655
g7592 nor n7607 n7608 ; n7656
g7593 nor n7655 n7656 ; n7657
g7594 and n392_not n6233 ; n7658
g7595 and n710_not n5663 ; n7659
g7596 and n587_not n5939 ; n7660
g7597 nor n7659 n7660 ; n7661
g7598 and n7658_not n7661 ; n7662
g7599 and n3347 n5666 ; n7663
g7600 and n7662 n7663_not ; n7664
g7601 and a[17] n7664_not ; n7665
g7602 nor n7664 n7665 ; n7666
g7603 and a[17] n7665_not ; n7667
g7604 nor n7666 n7667 ; n7668
g7605 and n7589 n7591_not ; n7669
g7606 nor n7592 n7669 ; n7670
g7607 and n7668_not n7670 ; n7671
g7608 nor n7668 n7671 ; n7672
g7609 and n7670 n7671_not ; n7673
g7610 nor n7672 n7673 ; n7674
g7611 and n7576 n7588_not ; n7675
g7612 nor n7587 n7588 ; n7676
g7613 nor n7675 n7676 ; n7677
g7614 and n7560 n7572_not ; n7678
g7615 nor n7571 n7572 ; n7679
g7616 nor n7678 n7679 ; n7680
g7617 and n7535 n7537_not ; n7681
g7618 nor n7538 n7681 ; n7682
g7619 and n1877_not n3884 ; n7683
g7620 and n1992_not n3967 ; n7684
g7621 and n1913_not n4046 ; n7685
g7622 nor n7684 n7685 ; n7686
g7623 and n7683_not n7686 ; n7687
g7624 and n4050_not n7687 ; n7688
g7625 and n6007_not n7687 ; n7689
g7626 nor n7688 n7689 ; n7690
g7627 and a[26] n7690_not ; n7691
g7628 and a[26]_not n7690 ; n7692
g7629 nor n7691 n7692 ; n7693
g7630 and n7682 n7693_not ; n7694
g7631 and n7531 n7533_not ; n7695
g7632 nor n7534 n7695 ; n7696
g7633 and n1913_not n3884 ; n7697
g7634 and n2057_not n3967 ; n7698
g7635 and n1992_not n4046 ; n7699
g7636 nor n7698 n7699 ; n7700
g7637 and n7697_not n7700 ; n7701
g7638 and n4050_not n7701 ; n7702
g7639 and n5834_not n7701 ; n7703
g7640 nor n7702 n7703 ; n7704
g7641 and a[26] n7704_not ; n7705
g7642 and a[26]_not n7704 ; n7706
g7643 nor n7705 n7706 ; n7707
g7644 and n7696 n7707_not ; n7708
g7645 and n7402 n7529 ; n7709
g7646 nor n7530 n7709 ; n7710
g7647 and n1992_not n3884 ; n7711
g7648 and n2152_not n3967 ; n7712
g7649 and n2057_not n4046 ; n7713
g7650 nor n7712 n7713 ; n7714
g7651 and n7711_not n7714 ; n7715
g7652 and n4050_not n7715 ; n7716
g7653 and n6143_not n7715 ; n7717
g7654 nor n7716 n7717 ; n7718
g7655 and a[26] n7718_not ; n7719
g7656 and a[26]_not n7718 ; n7720
g7657 nor n7719 n7720 ; n7721
g7658 and n7710 n7721_not ; n7722
g7659 and n7420 n7527 ; n7723
g7660 nor n7528 n7723 ; n7724
g7661 and n2057_not n3884 ; n7725
g7662 and n2189_not n3967 ; n7726
g7663 and n2152_not n4046 ; n7727
g7664 nor n7726 n7727 ; n7728
g7665 and n7725_not n7728 ; n7729
g7666 and n4050_not n7729 ; n7730
g7667 and n6479_not n7729 ; n7731
g7668 nor n7730 n7731 ; n7732
g7669 and a[26] n7732_not ; n7733
g7670 and a[26]_not n7732 ; n7734
g7671 nor n7733 n7734 ; n7735
g7672 and n7724 n7735_not ; n7736
g7673 and n7438 n7525 ; n7737
g7674 nor n7526 n7737 ; n7738
g7675 and n2152_not n3884 ; n7739
g7676 and n2291_not n3967 ; n7740
g7677 and n2189_not n4046 ; n7741
g7678 nor n7740 n7741 ; n7742
g7679 and n7739_not n7742 ; n7743
g7680 and n4050_not n7743 ; n7744
g7681 and n6492_not n7743 ; n7745
g7682 nor n7744 n7745 ; n7746
g7683 and a[26] n7746_not ; n7747
g7684 and a[26]_not n7746 ; n7748
g7685 nor n7747 n7748 ; n7749
g7686 and n7738 n7749_not ; n7750
g7687 and n7456 n7523 ; n7751
g7688 nor n7524 n7751 ; n7752
g7689 and n2189_not n3884 ; n7753
g7690 and n2388_not n3967 ; n7754
g7691 and n2291_not n4046 ; n7755
g7692 nor n7754 n7755 ; n7756
g7693 and n7753_not n7756 ; n7757
g7694 and n4050_not n7757 ; n7758
g7695 and n6122_not n7757 ; n7759
g7696 nor n7758 n7759 ; n7760
g7697 and a[26] n7760_not ; n7761
g7698 and a[26]_not n7760 ; n7762
g7699 nor n7761 n7762 ; n7763
g7700 and n7752 n7763_not ; n7764
g7701 nor n7478 n7522 ; n7765
g7702 nor n7521 n7522 ; n7766
g7703 nor n7765 n7766 ; n7767
g7704 and n2291_not n3884 ; n7768
g7705 and n2464_not n3967 ; n7769
g7706 and n2388_not n4046 ; n7770
g7707 nor n7769 n7770 ; n7771
g7708 and n7768_not n7771 ; n7772
g7709 and n4050_not n7772 ; n7773
g7710 and n6541_not n7772 ; n7774
g7711 nor n7773 n7774 ; n7775
g7712 and a[26] n7775_not ; n7776
g7713 and a[26]_not n7775 ; n7777
g7714 nor n7776 n7777 ; n7778
g7715 nor n7767 n7778 ; n7779
g7716 and n2388_not n3884 ; n7780
g7717 and n2533_not n3967 ; n7781
g7718 and n2464_not n4046 ; n7782
g7719 nor n7781 n7782 ; n7783
g7720 and n7780_not n7783 ; n7784
g7721 and n4050 n6591 ; n7785
g7722 and n7784 n7785_not ; n7786
g7723 and a[26] n7786_not ; n7787
g7724 nor n7786 n7787 ; n7788
g7725 and a[26] n7787_not ; n7789
g7726 nor n7788 n7789 ; n7790
g7727 and n7516 n7519 ; n7791
g7728 nor n7520 n7791 ; n7792
g7729 and n7790_not n7792 ; n7793
g7730 nor n7790 n7793 ; n7794
g7731 and n7792 n7793_not ; n7795
g7732 nor n7794 n7795 ; n7796
g7733 and n2464_not n3884 ; n7797
g7734 and n2571_not n3967 ; n7798
g7735 and n2533_not n4046 ; n7799
g7736 nor n7798 n7799 ; n7800
g7737 and n7797_not n7800 ; n7801
g7738 and n4050 n6646 ; n7802
g7739 and n7801 n7802_not ; n7803
g7740 and a[26] n7803_not ; n7804
g7741 nor n7803 n7804 ; n7805
g7742 and a[26] n7804_not ; n7806
g7743 nor n7805 n7806 ; n7807
g7744 and n7492_not n7503 ; n7808
g7745 nor n7504 n7808 ; n7809
g7746 and n7807_not n7809 ; n7810
g7747 nor n7807 n7810 ; n7811
g7748 and n7809 n7810_not ; n7812
g7749 nor n7811 n7812 ; n7813
g7750 and n7489 n7491_not ; n7814
g7751 nor n7492 n7814 ; n7815
g7752 and n2533_not n3884 ; n7816
g7753 and n2674_not n3967 ; n7817
g7754 and n2571_not n4046 ; n7818
g7755 nor n7817 n7818 ; n7819
g7756 and n7816_not n7819 ; n7820
g7757 and n4050_not n7820 ; n7821
g7758 and n6695_not n7820 ; n7822
g7759 nor n7821 n7822 ; n7823
g7760 and a[26] n7823_not ; n7824
g7761 and a[26]_not n7823 ; n7825
g7762 nor n7824 n7825 ; n7826
g7763 and n7815 n7826_not ; n7827
g7764 and n2829_not n4046 ; n7828
g7765 and n2736_not n3884 ; n7829
g7766 nor n7828 n7829 ; n7830
g7767 and n4050 n7469_not ; n7831
g7768 and n7830 n7831_not ; n7832
g7769 and a[26] n7832_not ; n7833
g7770 and a[26] n7833_not ; n7834
g7771 nor n7832 n7833 ; n7835
g7772 nor n7834 n7835 ; n7836
g7773 nor n2829 n3880 ; n7837
g7774 and a[26] n7837_not ; n7838
g7775 and n7836_not n7838 ; n7839
g7776 and n2674_not n3884 ; n7840
g7777 and n2829_not n3967 ; n7841
g7778 and n2736_not n4046 ; n7842
g7779 nor n7841 n7842 ; n7843
g7780 and n7840_not n7843 ; n7844
g7781 and n4050_not n7844 ; n7845
g7782 and n6798_not n7844 ; n7846
g7783 nor n7845 n7846 ; n7847
g7784 and a[26] n7847_not ; n7848
g7785 and a[26]_not n7847 ; n7849
g7786 nor n7848 n7849 ; n7850
g7787 and n7839 n7850_not ; n7851
g7788 and n7490 n7851 ; n7852
g7789 and n7851 n7852_not ; n7853
g7790 and n7490 n7852_not ; n7854
g7791 nor n7853 n7854 ; n7855
g7792 and n2571_not n3884 ; n7856
g7793 and n2736_not n3967 ; n7857
g7794 and n2674_not n4046 ; n7858
g7795 nor n7857 n7858 ; n7859
g7796 and n7856_not n7859 ; n7860
g7797 and n4050 n6806 ; n7861
g7798 and n7860 n7861_not ; n7862
g7799 and a[26] n7862_not ; n7863
g7800 and a[26] n7863_not ; n7864
g7801 nor n7862 n7863 ; n7865
g7802 nor n7864 n7865 ; n7866
g7803 nor n7855 n7866 ; n7867
g7804 nor n7852 n7867 ; n7868
g7805 and n7815_not n7826 ; n7869
g7806 nor n7827 n7869 ; n7870
g7807 and n7868_not n7870 ; n7871
g7808 nor n7827 n7871 ; n7872
g7809 nor n7813 n7872 ; n7873
g7810 nor n7810 n7873 ; n7874
g7811 nor n7796 n7874 ; n7875
g7812 nor n7793 n7875 ; n7876
g7813 nor n7767 n7779 ; n7877
g7814 nor n7778 n7779 ; n7878
g7815 nor n7877 n7878 ; n7879
g7816 nor n7876 n7879 ; n7880
g7817 nor n7779 n7880 ; n7881
g7818 and n7752 n7764_not ; n7882
g7819 nor n7763 n7764 ; n7883
g7820 nor n7882 n7883 ; n7884
g7821 nor n7881 n7884 ; n7885
g7822 nor n7764 n7885 ; n7886
g7823 and n7738 n7750_not ; n7887
g7824 nor n7749 n7750 ; n7888
g7825 nor n7887 n7888 ; n7889
g7826 nor n7886 n7889 ; n7890
g7827 nor n7750 n7890 ; n7891
g7828 and n7724 n7736_not ; n7892
g7829 nor n7735 n7736 ; n7893
g7830 nor n7892 n7893 ; n7894
g7831 nor n7891 n7894 ; n7895
g7832 nor n7736 n7895 ; n7896
g7833 and n7710 n7722_not ; n7897
g7834 nor n7721 n7722 ; n7898
g7835 nor n7897 n7898 ; n7899
g7836 nor n7896 n7899 ; n7900
g7837 nor n7722 n7900 ; n7901
g7838 and n7696 n7708_not ; n7902
g7839 nor n7707 n7708 ; n7903
g7840 nor n7902 n7903 ; n7904
g7841 nor n7901 n7904 ; n7905
g7842 nor n7708 n7905 ; n7906
g7843 and n7682 n7694_not ; n7907
g7844 nor n7693 n7694 ; n7908
g7845 nor n7907 n7908 ; n7909
g7846 nor n7906 n7909 ; n7910
g7847 nor n7694 n7910 ; n7911
g7848 and n7553 n7555_not ; n7912
g7849 nor n7556 n7912 ; n7913
g7850 and n7911_not n7913 ; n7914
g7851 and n1472_not n4694 ; n7915
g7852 and n1665_not n4533 ; n7916
g7853 and n1572_not n4604 ; n7917
g7854 nor n7916 n7917 ; n7918
g7855 and n7915_not n7918 ; n7919
g7856 and n4536 n5139 ; n7920
g7857 and n7919 n7920_not ; n7921
g7858 and a[23] n7921_not ; n7922
g7859 nor n7921 n7922 ; n7923
g7860 and a[23] n7922_not ; n7924
g7861 nor n7923 n7924 ; n7925
g7862 and n7911 n7913_not ; n7926
g7863 nor n7914 n7926 ; n7927
g7864 and n7925_not n7927 ; n7928
g7865 nor n7914 n7928 ; n7929
g7866 nor n7680 n7929 ; n7930
g7867 and n7680 n7929 ; n7931
g7868 nor n7930 n7931 ; n7932
g7869 and n1060_not n5496 ; n7933
g7870 and n1235_not n4935 ; n7934
g7871 and n1178_not n5407 ; n7935
g7872 nor n7934 n7935 ; n7936
g7873 and n7933_not n7936 ; n7937
g7874 and n4429 n4938 ; n7938
g7875 and n7937 n7938_not ; n7939
g7876 and a[20] n7939_not ; n7940
g7877 and a[20] n7940_not ; n7941
g7878 nor n7939 n7940 ; n7942
g7879 nor n7941 n7942 ; n7943
g7880 and n7932 n7943_not ; n7944
g7881 nor n7930 n7944 ; n7945
g7882 nor n7677 n7945 ; n7946
g7883 and n7677 n7945 ; n7947
g7884 nor n7946 n7947 ; n7948
g7885 and n587_not n6233 ; n7949
g7886 and n867_not n5663 ; n7950
g7887 and n710_not n5939 ; n7951
g7888 nor n7950 n7951 ; n7952
g7889 and n7949_not n7952 ; n7953
g7890 and n3331 n5666 ; n7954
g7891 and n7953 n7954_not ; n7955
g7892 and a[17] n7955_not ; n7956
g7893 and a[17] n7956_not ; n7957
g7894 nor n7955 n7956 ; n7958
g7895 nor n7957 n7958 ; n7959
g7896 and n7948 n7959_not ; n7960
g7897 nor n7946 n7960 ; n7961
g7898 nor n7674 n7961 ; n7962
g7899 nor n7671 n7962 ; n7963
g7900 nor n7657 n7963 ; n7964
g7901 and n7657 n7963 ; n7965
g7902 nor n7964 n7965 ; n7966
g7903 and n3456_not n7101 ; n7967
g7904 and n3539_not n6402 ; n7968
g7905 and n3605_not n6951 ; n7969
g7906 nor n7968 n7969 ; n7970
g7907 and n7967_not n7970 ; n7971
g7908 and n3627 n6397 ; n7972
g7909 and n7971 n7972_not ; n7973
g7910 and a[14] n7973_not ; n7974
g7911 and a[14] n7974_not ; n7975
g7912 nor n7973 n7974 ; n7976
g7913 nor n7975 n7976 ; n7977
g7914 and n7966 n7977_not ; n7978
g7915 nor n7964 n7978 ; n7979
g7916 nor n7654 n7979 ; n7980
g7917 and n7654 n7979 ; n7981
g7918 nor n7980 n7981 ; n7982
g7919 and n7286 n7289_not ; n7983
g7920 and n3877_not n7983 ; n7984
g7921 and n3964_not n7291 ; n7985
g7922 and n4045_not n7632 ; n7986
g7923 nor n7985 n7986 ; n7987
g7924 and n7984_not n7987 ; n7988
g7925 and n4067 n7294 ; n7989
g7926 and n7988 n7989_not ; n7990
g7927 and a[11] n7990_not ; n7991
g7928 and a[11] n7991_not ; n7992
g7929 nor n7990 n7991 ; n7993
g7930 nor n7992 n7993 ; n7994
g7931 and n7982 n7994_not ; n7995
g7932 nor n7980 n7995 ; n7996
g7933 and n4515_not n7983 ; n7997
g7934 and n4045_not n7291 ; n7998
g7935 and n3877_not n7632 ; n7999
g7936 nor n7998 n7999 ; n8000
g7937 and n7997_not n8000 ; n8001
g7938 and n7294_not n8001 ; n8002
g7939 and n4715_not n8001 ; n8003
g7940 nor n8002 n8003 ; n8004
g7941 and a[11] n8004_not ; n8005
g7942 and a[11]_not n8004 ; n8006
g7943 nor n8005 n8006 ; n8007
g7944 nor n7996 n8007 ; n8008
g7945 and n7996 n8007 ; n8009
g7946 nor n8008 n8009 ; n8010
g7947 nor n7625 n7629 ; n8011
g7948 nor n7628 n7629 ; n8012
g7949 nor n8011 n8012 ; n8013
g7950 and n8010 n8013_not ; n8014
g7951 nor n8008 n8014 ; n8015
g7952 and n7644 n7646_not ; n8016
g7953 nor n7647 n8016 ; n8017
g7954 and n8015_not n8017 ; n8018
g7955 and n8010 n8014_not ; n8019
g7956 nor n8013 n8014 ; n8020
g7957 nor n8019 n8020 ; n8021
g7958 and n7966 n7978_not ; n8022
g7959 nor n7977 n7978 ; n8023
g7960 nor n8022 n8023 ; n8024
g7961 and n7674 n7961 ; n8025
g7962 nor n7962 n8025 ; n8026
g7963 and n3605_not n7101 ; n8027
g7964 and n3012_not n6402 ; n8028
g7965 and n3539_not n6951 ; n8029
g7966 nor n8028 n8029 ; n8030
g7967 and n8027_not n8030 ; n8031
g7968 and n6397_not n8031 ; n8032
g7969 and n4084_not n8031 ; n8033
g7970 nor n8032 n8033 ; n8034
g7971 and a[14] n8034_not ; n8035
g7972 and a[14]_not n8034 ; n8036
g7973 nor n8035 n8036 ; n8037
g7974 and n8026 n8037_not ; n8038
g7975 and n7948 n7960_not ; n8039
g7976 nor n7959 n7960 ; n8040
g7977 nor n8039 n8040 ; n8041
g7978 and n7932 n7944_not ; n8042
g7979 nor n7943 n7944 ; n8043
g7980 nor n8042 n8043 ; n8044
g7981 and n1572_not n4694 ; n8045
g7982 and n1779_not n4533 ; n8046
g7983 and n1665_not n4604 ; n8047
g7984 nor n8046 n8047 ; n8048
g7985 and n8045_not n8048 ; n8049
g7986 and n4536 n5561 ; n8050
g7987 and n8049 n8050_not ; n8051
g7988 and a[23] n8051_not ; n8052
g7989 nor n8051 n8052 ; n8053
g7990 and a[23] n8052_not ; n8054
g7991 nor n8053 n8054 ; n8055
g7992 nor n7906 n7910 ; n8056
g7993 nor n7909 n7910 ; n8057
g7994 nor n8056 n8057 ; n8058
g7995 nor n8055 n8058 ; n8059
g7996 nor n8055 n8059 ; n8060
g7997 nor n8058 n8059 ; n8061
g7998 nor n8060 n8061 ; n8062
g7999 and n1665_not n4694 ; n8063
g8000 and n1877_not n4533 ; n8064
g8001 and n1779_not n4604 ; n8065
g8002 nor n8064 n8065 ; n8066
g8003 and n8063_not n8066 ; n8067
g8004 and n4536 n5328 ; n8068
g8005 and n8067 n8068_not ; n8069
g8006 and a[23] n8069_not ; n8070
g8007 nor n8069 n8070 ; n8071
g8008 and a[23] n8070_not ; n8072
g8009 nor n8071 n8072 ; n8073
g8010 nor n7901 n7905 ; n8074
g8011 nor n7904 n7905 ; n8075
g8012 nor n8074 n8075 ; n8076
g8013 nor n8073 n8076 ; n8077
g8014 nor n8073 n8077 ; n8078
g8015 nor n8076 n8077 ; n8079
g8016 nor n8078 n8079 ; n8080
g8017 and n1779_not n4694 ; n8081
g8018 and n1913_not n4533 ; n8082
g8019 and n1877_not n4604 ; n8083
g8020 nor n8082 n8083 ; n8084
g8021 and n8081_not n8084 ; n8085
g8022 and n4536 n5851 ; n8086
g8023 and n8085 n8086_not ; n8087
g8024 and a[23] n8087_not ; n8088
g8025 nor n8087 n8088 ; n8089
g8026 and a[23] n8088_not ; n8090
g8027 nor n8089 n8090 ; n8091
g8028 nor n7896 n7900 ; n8092
g8029 nor n7899 n7900 ; n8093
g8030 nor n8092 n8093 ; n8094
g8031 nor n8091 n8094 ; n8095
g8032 nor n8091 n8095 ; n8096
g8033 nor n8094 n8095 ; n8097
g8034 nor n8096 n8097 ; n8098
g8035 and n1877_not n4694 ; n8099
g8036 and n1992_not n4533 ; n8100
g8037 and n1913_not n4604 ; n8101
g8038 nor n8100 n8101 ; n8102
g8039 and n8099_not n8102 ; n8103
g8040 and n4536 n6007 ; n8104
g8041 and n8103 n8104_not ; n8105
g8042 and a[23] n8105_not ; n8106
g8043 nor n8105 n8106 ; n8107
g8044 and a[23] n8106_not ; n8108
g8045 nor n8107 n8108 ; n8109
g8046 nor n7891 n7895 ; n8110
g8047 nor n7894 n7895 ; n8111
g8048 nor n8110 n8111 ; n8112
g8049 nor n8109 n8112 ; n8113
g8050 nor n8109 n8113 ; n8114
g8051 nor n8112 n8113 ; n8115
g8052 nor n8114 n8115 ; n8116
g8053 and n1913_not n4694 ; n8117
g8054 and n2057_not n4533 ; n8118
g8055 and n1992_not n4604 ; n8119
g8056 nor n8118 n8119 ; n8120
g8057 and n8117_not n8120 ; n8121
g8058 and n4536 n5834 ; n8122
g8059 and n8121 n8122_not ; n8123
g8060 and a[23] n8123_not ; n8124
g8061 nor n8123 n8124 ; n8125
g8062 and a[23] n8124_not ; n8126
g8063 nor n8125 n8126 ; n8127
g8064 nor n7886 n7890 ; n8128
g8065 nor n7889 n7890 ; n8129
g8066 nor n8128 n8129 ; n8130
g8067 nor n8127 n8130 ; n8131
g8068 nor n8127 n8131 ; n8132
g8069 nor n8130 n8131 ; n8133
g8070 nor n8132 n8133 ; n8134
g8071 and n1992_not n4694 ; n8135
g8072 and n2152_not n4533 ; n8136
g8073 and n2057_not n4604 ; n8137
g8074 nor n8136 n8137 ; n8138
g8075 and n8135_not n8138 ; n8139
g8076 and n4536 n6143 ; n8140
g8077 and n8139 n8140_not ; n8141
g8078 and a[23] n8141_not ; n8142
g8079 nor n8141 n8142 ; n8143
g8080 and a[23] n8142_not ; n8144
g8081 nor n8143 n8144 ; n8145
g8082 nor n7881 n7885 ; n8146
g8083 nor n7884 n7885 ; n8147
g8084 nor n8146 n8147 ; n8148
g8085 nor n8145 n8148 ; n8149
g8086 nor n8145 n8149 ; n8150
g8087 nor n8148 n8149 ; n8151
g8088 nor n8150 n8151 ; n8152
g8089 and n2057_not n4694 ; n8153
g8090 and n2189_not n4533 ; n8154
g8091 and n2152_not n4604 ; n8155
g8092 nor n8154 n8155 ; n8156
g8093 and n8153_not n8156 ; n8157
g8094 and n4536 n6479 ; n8158
g8095 and n8157 n8158_not ; n8159
g8096 and a[23] n8159_not ; n8160
g8097 nor n8159 n8160 ; n8161
g8098 and a[23] n8160_not ; n8162
g8099 nor n8161 n8162 ; n8163
g8100 nor n7876 n7880 ; n8164
g8101 nor n7879 n7880 ; n8165
g8102 nor n8164 n8165 ; n8166
g8103 nor n8163 n8166 ; n8167
g8104 nor n8163 n8167 ; n8168
g8105 nor n8166 n8167 ; n8169
g8106 nor n8168 n8169 ; n8170
g8107 and n7796 n7874 ; n8171
g8108 nor n7875 n8171 ; n8172
g8109 and n2152_not n4694 ; n8173
g8110 and n2291_not n4533 ; n8174
g8111 and n2189_not n4604 ; n8175
g8112 nor n8174 n8175 ; n8176
g8113 and n8173_not n8176 ; n8177
g8114 and n4536_not n8177 ; n8178
g8115 and n6492_not n8177 ; n8179
g8116 nor n8178 n8179 ; n8180
g8117 and a[23] n8180_not ; n8181
g8118 and a[23]_not n8180 ; n8182
g8119 nor n8181 n8182 ; n8183
g8120 and n8172 n8183_not ; n8184
g8121 and n7813 n7872 ; n8185
g8122 nor n7873 n8185 ; n8186
g8123 and n2189_not n4694 ; n8187
g8124 and n2388_not n4533 ; n8188
g8125 and n2291_not n4604 ; n8189
g8126 nor n8188 n8189 ; n8190
g8127 and n8187_not n8190 ; n8191
g8128 and n4536_not n8191 ; n8192
g8129 and n6122_not n8191 ; n8193
g8130 nor n8192 n8193 ; n8194
g8131 and a[23] n8194_not ; n8195
g8132 and a[23]_not n8194 ; n8196
g8133 nor n8195 n8196 ; n8197
g8134 and n8186 n8197_not ; n8198
g8135 and n2291_not n4694 ; n8199
g8136 and n2464_not n4533 ; n8200
g8137 and n2388_not n4604 ; n8201
g8138 nor n8200 n8201 ; n8202
g8139 and n8199_not n8202 ; n8203
g8140 and n4536 n6541 ; n8204
g8141 and n8203 n8204_not ; n8205
g8142 and a[23] n8205_not ; n8206
g8143 nor n8205 n8206 ; n8207
g8144 and a[23] n8206_not ; n8208
g8145 nor n8207 n8208 ; n8209
g8146 and n7868 n7870_not ; n8210
g8147 nor n7871 n8210 ; n8211
g8148 and n8209_not n8211 ; n8212
g8149 nor n8209 n8212 ; n8213
g8150 and n8211 n8212_not ; n8214
g8151 nor n8213 n8214 ; n8215
g8152 nor n7855 n7867 ; n8216
g8153 nor n7866 n7867 ; n8217
g8154 nor n8216 n8217 ; n8218
g8155 and n2388_not n4694 ; n8219
g8156 and n2533_not n4533 ; n8220
g8157 and n2464_not n4604 ; n8221
g8158 nor n8220 n8221 ; n8222
g8159 and n8219_not n8222 ; n8223
g8160 and n4536_not n8223 ; n8224
g8161 and n6591_not n8223 ; n8225
g8162 nor n8224 n8225 ; n8226
g8163 and a[23] n8226_not ; n8227
g8164 and a[23]_not n8226 ; n8228
g8165 nor n8227 n8228 ; n8229
g8166 nor n8218 n8229 ; n8230
g8167 and n2464_not n4694 ; n8231
g8168 and n2571_not n4533 ; n8232
g8169 and n2533_not n4604 ; n8233
g8170 nor n8232 n8233 ; n8234
g8171 and n8231_not n8234 ; n8235
g8172 and n4536 n6646 ; n8236
g8173 and n8235 n8236_not ; n8237
g8174 and a[23] n8237_not ; n8238
g8175 nor n8237 n8238 ; n8239
g8176 and a[23] n8238_not ; n8240
g8177 nor n8239 n8240 ; n8241
g8178 and n7839_not n7850 ; n8242
g8179 nor n7851 n8242 ; n8243
g8180 and n8241_not n8243 ; n8244
g8181 nor n8241 n8244 ; n8245
g8182 and n8243 n8244_not ; n8246
g8183 nor n8245 n8246 ; n8247
g8184 and n7836 n7838_not ; n8248
g8185 nor n7839 n8248 ; n8249
g8186 and n2533_not n4694 ; n8250
g8187 and n2674_not n4533 ; n8251
g8188 and n2571_not n4604 ; n8252
g8189 nor n8251 n8252 ; n8253
g8190 and n8250_not n8253 ; n8254
g8191 and n4536_not n8254 ; n8255
g8192 and n6695_not n8254 ; n8256
g8193 nor n8255 n8256 ; n8257
g8194 and a[23] n8257_not ; n8258
g8195 and a[23]_not n8257 ; n8259
g8196 nor n8258 n8259 ; n8260
g8197 and n8249 n8260_not ; n8261
g8198 and n2829_not n4604 ; n8262
g8199 and n2736_not n4694 ; n8263
g8200 nor n8262 n8263 ; n8264
g8201 and n4536 n7469_not ; n8265
g8202 and n8264 n8265_not ; n8266
g8203 and a[23] n8266_not ; n8267
g8204 and a[23] n8267_not ; n8268
g8205 nor n8266 n8267 ; n8269
g8206 nor n8268 n8269 ; n8270
g8207 nor n2829 n4528 ; n8271
g8208 and a[23] n8271_not ; n8272
g8209 and n8270_not n8272 ; n8273
g8210 and n2674_not n4694 ; n8274
g8211 and n2829_not n4533 ; n8275
g8212 and n2736_not n4604 ; n8276
g8213 nor n8275 n8276 ; n8277
g8214 and n8274_not n8277 ; n8278
g8215 and n4536_not n8278 ; n8279
g8216 and n6798_not n8278 ; n8280
g8217 nor n8279 n8280 ; n8281
g8218 and a[23] n8281_not ; n8282
g8219 and a[23]_not n8281 ; n8283
g8220 nor n8282 n8283 ; n8284
g8221 and n8273 n8284_not ; n8285
g8222 and n7837 n8285 ; n8286
g8223 and n8285 n8286_not ; n8287
g8224 and n7837 n8286_not ; n8288
g8225 nor n8287 n8288 ; n8289
g8226 and n2571_not n4694 ; n8290
g8227 and n2736_not n4533 ; n8291
g8228 and n2674_not n4604 ; n8292
g8229 nor n8291 n8292 ; n8293
g8230 and n8290_not n8293 ; n8294
g8231 and n4536 n6806 ; n8295
g8232 and n8294 n8295_not ; n8296
g8233 and a[23] n8296_not ; n8297
g8234 and a[23] n8297_not ; n8298
g8235 nor n8296 n8297 ; n8299
g8236 nor n8298 n8299 ; n8300
g8237 nor n8289 n8300 ; n8301
g8238 nor n8286 n8301 ; n8302
g8239 and n8249_not n8260 ; n8303
g8240 nor n8261 n8303 ; n8304
g8241 and n8302_not n8304 ; n8305
g8242 nor n8261 n8305 ; n8306
g8243 nor n8247 n8306 ; n8307
g8244 nor n8244 n8307 ; n8308
g8245 and n8218 n8229 ; n8309
g8246 nor n8230 n8309 ; n8310
g8247 and n8308_not n8310 ; n8311
g8248 nor n8230 n8311 ; n8312
g8249 nor n8215 n8312 ; n8313
g8250 nor n8212 n8313 ; n8314
g8251 and n8186 n8198_not ; n8315
g8252 nor n8197 n8198 ; n8316
g8253 nor n8315 n8316 ; n8317
g8254 nor n8314 n8317 ; n8318
g8255 nor n8198 n8318 ; n8319
g8256 and n8172_not n8183 ; n8320
g8257 nor n8184 n8320 ; n8321
g8258 and n8319_not n8321 ; n8322
g8259 nor n8184 n8322 ; n8323
g8260 nor n8170 n8323 ; n8324
g8261 nor n8167 n8324 ; n8325
g8262 nor n8152 n8325 ; n8326
g8263 nor n8149 n8326 ; n8327
g8264 nor n8134 n8327 ; n8328
g8265 nor n8131 n8328 ; n8329
g8266 nor n8116 n8329 ; n8330
g8267 nor n8113 n8330 ; n8331
g8268 nor n8098 n8331 ; n8332
g8269 nor n8095 n8332 ; n8333
g8270 nor n8080 n8333 ; n8334
g8271 nor n8077 n8334 ; n8335
g8272 nor n8062 n8335 ; n8336
g8273 nor n8059 n8336 ; n8337
g8274 and n7925 n7927_not ; n8338
g8275 nor n7928 n8338 ; n8339
g8276 and n8337_not n8339 ; n8340
g8277 and n1178_not n5496 ; n8341
g8278 and n1364_not n4935 ; n8342
g8279 and n1235_not n5407 ; n8343
g8280 nor n8342 n8343 ; n8344
g8281 and n8341_not n8344 ; n8345
g8282 and n4861 n4938 ; n8346
g8283 and n8345 n8346_not ; n8347
g8284 and a[20] n8347_not ; n8348
g8285 nor n8347 n8348 ; n8349
g8286 and a[20] n8348_not ; n8350
g8287 nor n8349 n8350 ; n8351
g8288 and n8337 n8339_not ; n8352
g8289 nor n8340 n8352 ; n8353
g8290 and n8351_not n8353 ; n8354
g8291 nor n8340 n8354 ; n8355
g8292 nor n8044 n8355 ; n8356
g8293 and n8044 n8355 ; n8357
g8294 nor n8356 n8357 ; n8358
g8295 and n710_not n6233 ; n8359
g8296 and n958_not n5663 ; n8360
g8297 and n867_not n5939 ; n8361
g8298 nor n8360 n8361 ; n8362
g8299 and n8359_not n8362 ; n8363
g8300 and n4179 n5666 ; n8364
g8301 and n8363 n8364_not ; n8365
g8302 and a[17] n8365_not ; n8366
g8303 and a[17] n8366_not ; n8367
g8304 nor n8365 n8366 ; n8368
g8305 nor n8367 n8368 ; n8369
g8306 and n8358 n8369_not ; n8370
g8307 nor n8356 n8370 ; n8371
g8308 nor n8041 n8371 ; n8372
g8309 and n8041 n8371 ; n8373
g8310 nor n8372 n8373 ; n8374
g8311 and n3539_not n7101 ; n8375
g8312 and n392_not n6402 ; n8376
g8313 and n3012_not n6951 ; n8377
g8314 nor n8376 n8377 ; n8378
g8315 and n8375_not n8378 ; n8379
g8316 and n3715 n6397 ; n8380
g8317 and n8379 n8380_not ; n8381
g8318 and a[14] n8381_not ; n8382
g8319 and a[14] n8382_not ; n8383
g8320 nor n8381 n8382 ; n8384
g8321 nor n8383 n8384 ; n8385
g8322 and n8374 n8385_not ; n8386
g8323 nor n8372 n8386 ; n8387
g8324 and n8026_not n8037 ; n8388
g8325 nor n8038 n8388 ; n8389
g8326 and n8387_not n8389 ; n8390
g8327 nor n8038 n8390 ; n8391
g8328 nor n8024 n8391 ; n8392
g8329 and n8024 n8391 ; n8393
g8330 nor n8392 n8393 ; n8394
g8331 and n4045_not n7983 ; n8395
g8332 and n3805_not n7291 ; n8396
g8333 and n3964_not n7632 ; n8397
g8334 nor n8396 n8397 ; n8398
g8335 and n8395_not n8398 ; n8399
g8336 and n4477 n7294 ; n8400
g8337 and n8399 n8400_not ; n8401
g8338 and a[11] n8401_not ; n8402
g8339 and a[11] n8402_not ; n8403
g8340 nor n8401 n8402 ; n8404
g8341 nor n8403 n8404 ; n8405
g8342 and n8394 n8405_not ; n8406
g8343 nor n8392 n8406 ; n8407
g8344 and a[6]_not a[7] ; n8408
g8345 and a[6] a[7]_not ; n8409
g8346 nor n8408 n8409 ; n8410
g8347 and a[7] a[8]_not ; n8411
g8348 and a[7]_not a[8] ; n8412
g8349 nor n8411 n8412 ; n8413
g8350 and a[5] a[6]_not ; n8414
g8351 and a[5]_not a[6] ; n8415
g8352 nor n8414 n8415 ; n8416
g8353 and n8413_not n8416 ; n8417
g8354 and n8410 n8417 ; n8418
g8355 and n4515_not n8418 ; n8419
g8356 nor n4522 n8419 ; n8420
g8357 nor n8413 n8416 ; n8421
g8358 nor n8419 n8421 ; n8422
g8359 nor n8420 n8422 ; n8423
g8360 and a[8] n8423_not ; n8424
g8361 and a[8]_not n8423 ; n8425
g8362 nor n8424 n8425 ; n8426
g8363 nor n8407 n8426 ; n8427
g8364 and n7982 n7995_not ; n8428
g8365 nor n7994 n7995 ; n8429
g8366 nor n8428 n8429 ; n8430
g8367 and n8407 n8426 ; n8431
g8368 nor n8427 n8431 ; n8432
g8369 and n8430_not n8432 ; n8433
g8370 nor n8427 n8433 ; n8434
g8371 nor n8021 n8434 ; n8435
g8372 and n8021 n8434 ; n8436
g8373 nor n8435 n8436 ; n8437
g8374 nor n8430 n8433 ; n8438
g8375 and n8432 n8433_not ; n8439
g8376 nor n8438 n8439 ; n8440
g8377 and n8374 n8386_not ; n8441
g8378 nor n8385 n8386 ; n8442
g8379 nor n8441 n8442 ; n8443
g8380 and n8358 n8370_not ; n8444
g8381 nor n8369 n8370 ; n8445
g8382 nor n8444 n8445 ; n8446
g8383 and n8062 n8335 ; n8447
g8384 nor n8336 n8447 ; n8448
g8385 and n1235_not n5496 ; n8449
g8386 and n1472_not n4935 ; n8450
g8387 and n1364_not n5407 ; n8451
g8388 nor n8450 n8451 ; n8452
g8389 and n8449_not n8452 ; n8453
g8390 and n4938_not n8453 ; n8454
g8391 and n4848_not n8453 ; n8455
g8392 nor n8454 n8455 ; n8456
g8393 and a[20] n8456_not ; n8457
g8394 and a[20]_not n8456 ; n8458
g8395 nor n8457 n8458 ; n8459
g8396 and n8448 n8459_not ; n8460
g8397 and n8080 n8333 ; n8461
g8398 nor n8334 n8461 ; n8462
g8399 and n1364_not n5496 ; n8463
g8400 and n1572_not n4935 ; n8464
g8401 and n1472_not n5407 ; n8465
g8402 nor n8464 n8465 ; n8466
g8403 and n8463_not n8466 ; n8467
g8404 and n4938_not n8467 ; n8468
g8405 and n5114_not n8467 ; n8469
g8406 nor n8468 n8469 ; n8470
g8407 and a[20] n8470_not ; n8471
g8408 and a[20]_not n8470 ; n8472
g8409 nor n8471 n8472 ; n8473
g8410 and n8462 n8473_not ; n8474
g8411 and n8098 n8331 ; n8475
g8412 nor n8332 n8475 ; n8476
g8413 and n1472_not n5496 ; n8477
g8414 and n1665_not n4935 ; n8478
g8415 and n1572_not n5407 ; n8479
g8416 nor n8478 n8479 ; n8480
g8417 and n8477_not n8480 ; n8481
g8418 and n4938_not n8481 ; n8482
g8419 and n5139_not n8481 ; n8483
g8420 nor n8482 n8483 ; n8484
g8421 and a[20] n8484_not ; n8485
g8422 and a[20]_not n8484 ; n8486
g8423 nor n8485 n8486 ; n8487
g8424 and n8476 n8487_not ; n8488
g8425 and n8116 n8329 ; n8489
g8426 nor n8330 n8489 ; n8490
g8427 and n1572_not n5496 ; n8491
g8428 and n1779_not n4935 ; n8492
g8429 and n1665_not n5407 ; n8493
g8430 nor n8492 n8493 ; n8494
g8431 and n8491_not n8494 ; n8495
g8432 and n4938_not n8495 ; n8496
g8433 and n5561_not n8495 ; n8497
g8434 nor n8496 n8497 ; n8498
g8435 and a[20] n8498_not ; n8499
g8436 and a[20]_not n8498 ; n8500
g8437 nor n8499 n8500 ; n8501
g8438 and n8490 n8501_not ; n8502
g8439 and n8134 n8327 ; n8503
g8440 nor n8328 n8503 ; n8504
g8441 and n1665_not n5496 ; n8505
g8442 and n1877_not n4935 ; n8506
g8443 and n1779_not n5407 ; n8507
g8444 nor n8506 n8507 ; n8508
g8445 and n8505_not n8508 ; n8509
g8446 and n4938_not n8509 ; n8510
g8447 and n5328_not n8509 ; n8511
g8448 nor n8510 n8511 ; n8512
g8449 and a[20] n8512_not ; n8513
g8450 and a[20]_not n8512 ; n8514
g8451 nor n8513 n8514 ; n8515
g8452 and n8504 n8515_not ; n8516
g8453 and n8152 n8325 ; n8517
g8454 nor n8326 n8517 ; n8518
g8455 and n1779_not n5496 ; n8519
g8456 and n1913_not n4935 ; n8520
g8457 and n1877_not n5407 ; n8521
g8458 nor n8520 n8521 ; n8522
g8459 and n8519_not n8522 ; n8523
g8460 and n4938_not n8523 ; n8524
g8461 and n5851_not n8523 ; n8525
g8462 nor n8524 n8525 ; n8526
g8463 and a[20] n8526_not ; n8527
g8464 and a[20]_not n8526 ; n8528
g8465 nor n8527 n8528 ; n8529
g8466 and n8518 n8529_not ; n8530
g8467 and n8170 n8323 ; n8531
g8468 nor n8324 n8531 ; n8532
g8469 and n1877_not n5496 ; n8533
g8470 and n1992_not n4935 ; n8534
g8471 and n1913_not n5407 ; n8535
g8472 nor n8534 n8535 ; n8536
g8473 and n8533_not n8536 ; n8537
g8474 and n4938_not n8537 ; n8538
g8475 and n6007_not n8537 ; n8539
g8476 nor n8538 n8539 ; n8540
g8477 and a[20] n8540_not ; n8541
g8478 and a[20]_not n8540 ; n8542
g8479 nor n8541 n8542 ; n8543
g8480 and n8532 n8543_not ; n8544
g8481 and n1913_not n5496 ; n8545
g8482 and n2057_not n4935 ; n8546
g8483 and n1992_not n5407 ; n8547
g8484 nor n8546 n8547 ; n8548
g8485 and n8545_not n8548 ; n8549
g8486 and n4938 n5834 ; n8550
g8487 and n8549 n8550_not ; n8551
g8488 and a[20] n8551_not ; n8552
g8489 nor n8551 n8552 ; n8553
g8490 and a[20] n8552_not ; n8554
g8491 nor n8553 n8554 ; n8555
g8492 and n8319 n8321_not ; n8556
g8493 nor n8322 n8556 ; n8557
g8494 and n8555_not n8557 ; n8558
g8495 nor n8555 n8558 ; n8559
g8496 and n8557 n8558_not ; n8560
g8497 nor n8559 n8560 ; n8561
g8498 and n1992_not n5496 ; n8562
g8499 and n2152_not n4935 ; n8563
g8500 and n2057_not n5407 ; n8564
g8501 nor n8563 n8564 ; n8565
g8502 and n8562_not n8565 ; n8566
g8503 and n4938 n6143 ; n8567
g8504 and n8566 n8567_not ; n8568
g8505 and a[20] n8568_not ; n8569
g8506 nor n8568 n8569 ; n8570
g8507 and a[20] n8569_not ; n8571
g8508 nor n8570 n8571 ; n8572
g8509 nor n8314 n8318 ; n8573
g8510 nor n8317 n8318 ; n8574
g8511 nor n8573 n8574 ; n8575
g8512 nor n8572 n8575 ; n8576
g8513 nor n8572 n8576 ; n8577
g8514 nor n8575 n8576 ; n8578
g8515 nor n8577 n8578 ; n8579
g8516 and n8215 n8312 ; n8580
g8517 nor n8313 n8580 ; n8581
g8518 and n2057_not n5496 ; n8582
g8519 and n2189_not n4935 ; n8583
g8520 and n2152_not n5407 ; n8584
g8521 nor n8583 n8584 ; n8585
g8522 and n8582_not n8585 ; n8586
g8523 and n4938_not n8586 ; n8587
g8524 and n6479_not n8586 ; n8588
g8525 nor n8587 n8588 ; n8589
g8526 and a[20] n8589_not ; n8590
g8527 and a[20]_not n8589 ; n8591
g8528 nor n8590 n8591 ; n8592
g8529 and n8581 n8592_not ; n8593
g8530 and n8308 n8310_not ; n8594
g8531 nor n8311 n8594 ; n8595
g8532 and n2152_not n5496 ; n8596
g8533 and n2291_not n4935 ; n8597
g8534 and n2189_not n5407 ; n8598
g8535 nor n8597 n8598 ; n8599
g8536 and n8596_not n8599 ; n8600
g8537 and n4938_not n8600 ; n8601
g8538 and n6492_not n8600 ; n8602
g8539 nor n8601 n8602 ; n8603
g8540 and a[20] n8603_not ; n8604
g8541 and a[20]_not n8603 ; n8605
g8542 nor n8604 n8605 ; n8606
g8543 and n8595 n8606_not ; n8607
g8544 and n8247 n8306 ; n8608
g8545 nor n8307 n8608 ; n8609
g8546 and n2189_not n5496 ; n8610
g8547 and n2388_not n4935 ; n8611
g8548 and n2291_not n5407 ; n8612
g8549 nor n8611 n8612 ; n8613
g8550 and n8610_not n8613 ; n8614
g8551 and n4938_not n8614 ; n8615
g8552 and n6122_not n8614 ; n8616
g8553 nor n8615 n8616 ; n8617
g8554 and a[20] n8617_not ; n8618
g8555 and a[20]_not n8617 ; n8619
g8556 nor n8618 n8619 ; n8620
g8557 and n8609 n8620_not ; n8621
g8558 and n2291_not n5496 ; n8622
g8559 and n2464_not n4935 ; n8623
g8560 and n2388_not n5407 ; n8624
g8561 nor n8623 n8624 ; n8625
g8562 and n8622_not n8625 ; n8626
g8563 and n4938 n6541 ; n8627
g8564 and n8626 n8627_not ; n8628
g8565 and a[20] n8628_not ; n8629
g8566 nor n8628 n8629 ; n8630
g8567 and a[20] n8629_not ; n8631
g8568 nor n8630 n8631 ; n8632
g8569 and n8302 n8304_not ; n8633
g8570 nor n8305 n8633 ; n8634
g8571 and n8632_not n8634 ; n8635
g8572 nor n8632 n8635 ; n8636
g8573 and n8634 n8635_not ; n8637
g8574 nor n8636 n8637 ; n8638
g8575 nor n8289 n8301 ; n8639
g8576 nor n8300 n8301 ; n8640
g8577 nor n8639 n8640 ; n8641
g8578 and n2388_not n5496 ; n8642
g8579 and n2533_not n4935 ; n8643
g8580 and n2464_not n5407 ; n8644
g8581 nor n8643 n8644 ; n8645
g8582 and n8642_not n8645 ; n8646
g8583 and n4938_not n8646 ; n8647
g8584 and n6591_not n8646 ; n8648
g8585 nor n8647 n8648 ; n8649
g8586 and a[20] n8649_not ; n8650
g8587 and a[20]_not n8649 ; n8651
g8588 nor n8650 n8651 ; n8652
g8589 nor n8641 n8652 ; n8653
g8590 and n2464_not n5496 ; n8654
g8591 and n2571_not n4935 ; n8655
g8592 and n2533_not n5407 ; n8656
g8593 nor n8655 n8656 ; n8657
g8594 and n8654_not n8657 ; n8658
g8595 and n4938 n6646 ; n8659
g8596 and n8658 n8659_not ; n8660
g8597 and a[20] n8660_not ; n8661
g8598 nor n8660 n8661 ; n8662
g8599 and a[20] n8661_not ; n8663
g8600 nor n8662 n8663 ; n8664
g8601 and n8273_not n8284 ; n8665
g8602 nor n8285 n8665 ; n8666
g8603 and n8664_not n8666 ; n8667
g8604 nor n8664 n8667 ; n8668
g8605 and n8666 n8667_not ; n8669
g8606 nor n8668 n8669 ; n8670
g8607 and n8270 n8272_not ; n8671
g8608 nor n8273 n8671 ; n8672
g8609 and n2533_not n5496 ; n8673
g8610 and n2674_not n4935 ; n8674
g8611 and n2571_not n5407 ; n8675
g8612 nor n8674 n8675 ; n8676
g8613 and n8673_not n8676 ; n8677
g8614 and n4938_not n8677 ; n8678
g8615 and n6695_not n8677 ; n8679
g8616 nor n8678 n8679 ; n8680
g8617 and a[20] n8680_not ; n8681
g8618 and a[20]_not n8680 ; n8682
g8619 nor n8681 n8682 ; n8683
g8620 and n8672 n8683_not ; n8684
g8621 and n2829_not n5407 ; n8685
g8622 and n2736_not n5496 ; n8686
g8623 nor n8685 n8686 ; n8687
g8624 and n4938 n7469_not ; n8688
g8625 and n8687 n8688_not ; n8689
g8626 and a[20] n8689_not ; n8690
g8627 and a[20] n8690_not ; n8691
g8628 nor n8689 n8690 ; n8692
g8629 nor n8691 n8692 ; n8693
g8630 nor n2829 n4933 ; n8694
g8631 and a[20] n8694_not ; n8695
g8632 and n8693_not n8695 ; n8696
g8633 and n2674_not n5496 ; n8697
g8634 and n2829_not n4935 ; n8698
g8635 and n2736_not n5407 ; n8699
g8636 nor n8698 n8699 ; n8700
g8637 and n8697_not n8700 ; n8701
g8638 and n4938_not n8701 ; n8702
g8639 and n6798_not n8701 ; n8703
g8640 nor n8702 n8703 ; n8704
g8641 and a[20] n8704_not ; n8705
g8642 and a[20]_not n8704 ; n8706
g8643 nor n8705 n8706 ; n8707
g8644 and n8696 n8707_not ; n8708
g8645 and n8271 n8708 ; n8709
g8646 and n8708 n8709_not ; n8710
g8647 and n8271 n8709_not ; n8711
g8648 nor n8710 n8711 ; n8712
g8649 and n2571_not n5496 ; n8713
g8650 and n2736_not n4935 ; n8714
g8651 and n2674_not n5407 ; n8715
g8652 nor n8714 n8715 ; n8716
g8653 and n8713_not n8716 ; n8717
g8654 and n4938 n6806 ; n8718
g8655 and n8717 n8718_not ; n8719
g8656 and a[20] n8719_not ; n8720
g8657 and a[20] n8720_not ; n8721
g8658 nor n8719 n8720 ; n8722
g8659 nor n8721 n8722 ; n8723
g8660 nor n8712 n8723 ; n8724
g8661 nor n8709 n8724 ; n8725
g8662 and n8672_not n8683 ; n8726
g8663 nor n8684 n8726 ; n8727
g8664 and n8725_not n8727 ; n8728
g8665 nor n8684 n8728 ; n8729
g8666 nor n8670 n8729 ; n8730
g8667 nor n8667 n8730 ; n8731
g8668 and n8641 n8652 ; n8732
g8669 nor n8653 n8732 ; n8733
g8670 and n8731_not n8733 ; n8734
g8671 nor n8653 n8734 ; n8735
g8672 nor n8638 n8735 ; n8736
g8673 nor n8635 n8736 ; n8737
g8674 and n8609 n8621_not ; n8738
g8675 nor n8620 n8621 ; n8739
g8676 nor n8738 n8739 ; n8740
g8677 nor n8737 n8740 ; n8741
g8678 nor n8621 n8741 ; n8742
g8679 and n8595 n8607_not ; n8743
g8680 nor n8606 n8607 ; n8744
g8681 nor n8743 n8744 ; n8745
g8682 nor n8742 n8745 ; n8746
g8683 nor n8607 n8746 ; n8747
g8684 and n8581_not n8592 ; n8748
g8685 nor n8593 n8748 ; n8749
g8686 and n8747_not n8749 ; n8750
g8687 nor n8593 n8750 ; n8751
g8688 nor n8579 n8751 ; n8752
g8689 nor n8576 n8752 ; n8753
g8690 nor n8561 n8753 ; n8754
g8691 nor n8558 n8754 ; n8755
g8692 and n8532 n8544_not ; n8756
g8693 nor n8543 n8544 ; n8757
g8694 nor n8756 n8757 ; n8758
g8695 nor n8755 n8758 ; n8759
g8696 nor n8544 n8759 ; n8760
g8697 and n8518 n8530_not ; n8761
g8698 nor n8529 n8530 ; n8762
g8699 nor n8761 n8762 ; n8763
g8700 nor n8760 n8763 ; n8764
g8701 nor n8530 n8764 ; n8765
g8702 and n8504 n8516_not ; n8766
g8703 nor n8515 n8516 ; n8767
g8704 nor n8766 n8767 ; n8768
g8705 nor n8765 n8768 ; n8769
g8706 nor n8516 n8769 ; n8770
g8707 and n8490 n8502_not ; n8771
g8708 nor n8501 n8502 ; n8772
g8709 nor n8771 n8772 ; n8773
g8710 nor n8770 n8773 ; n8774
g8711 nor n8502 n8774 ; n8775
g8712 and n8476 n8488_not ; n8776
g8713 nor n8487 n8488 ; n8777
g8714 nor n8776 n8777 ; n8778
g8715 nor n8775 n8778 ; n8779
g8716 nor n8488 n8779 ; n8780
g8717 and n8462 n8474_not ; n8781
g8718 nor n8473 n8474 ; n8782
g8719 nor n8781 n8782 ; n8783
g8720 nor n8780 n8783 ; n8784
g8721 nor n8474 n8784 ; n8785
g8722 and n8448 n8460_not ; n8786
g8723 nor n8459 n8460 ; n8787
g8724 nor n8786 n8787 ; n8788
g8725 nor n8785 n8788 ; n8789
g8726 nor n8460 n8789 ; n8790
g8727 and n8351 n8353_not ; n8791
g8728 nor n8354 n8791 ; n8792
g8729 and n8790_not n8792 ; n8793
g8730 and n867_not n6233 ; n8794
g8731 and n1060_not n5663 ; n8795
g8732 and n958_not n5939 ; n8796
g8733 nor n8795 n8796 ; n8797
g8734 and n8794_not n8797 ; n8798
g8735 and n4204 n5666 ; n8799
g8736 and n8798 n8799_not ; n8800
g8737 and a[17] n8800_not ; n8801
g8738 nor n8800 n8801 ; n8802
g8739 and a[17] n8801_not ; n8803
g8740 nor n8802 n8803 ; n8804
g8741 and n8790 n8792_not ; n8805
g8742 nor n8793 n8805 ; n8806
g8743 and n8804_not n8806 ; n8807
g8744 nor n8793 n8807 ; n8808
g8745 nor n8446 n8808 ; n8809
g8746 and n8446 n8808 ; n8810
g8747 nor n8809 n8810 ; n8811
g8748 and n3012_not n7101 ; n8812
g8749 and n587_not n6402 ; n8813
g8750 and n392_not n6951 ; n8814
g8751 nor n8813 n8814 ; n8815
g8752 and n8812_not n8815 ; n8816
g8753 and n3018 n6397 ; n8817
g8754 and n8816 n8817_not ; n8818
g8755 and a[14] n8818_not ; n8819
g8756 and a[14] n8819_not ; n8820
g8757 nor n8818 n8819 ; n8821
g8758 nor n8820 n8821 ; n8822
g8759 and n8811 n8822_not ; n8823
g8760 nor n8809 n8823 ; n8824
g8761 nor n8443 n8824 ; n8825
g8762 and n8443 n8824 ; n8826
g8763 nor n8825 n8826 ; n8827
g8764 and n3805_not n7983 ; n8828
g8765 and n3605_not n7291 ; n8829
g8766 and n3456_not n7632 ; n8830
g8767 nor n8829 n8830 ; n8831
g8768 and n8828_not n8831 ; n8832
g8769 and n3818 n7294 ; n8833
g8770 and n8832 n8833_not ; n8834
g8771 and a[11] n8834_not ; n8835
g8772 and a[11] n8835_not ; n8836
g8773 nor n8834 n8835 ; n8837
g8774 nor n8836 n8837 ; n8838
g8775 and n8827 n8838_not ; n8839
g8776 nor n8825 n8839 ; n8840
g8777 and n3964_not n7983 ; n8841
g8778 and n3456_not n7291 ; n8842
g8779 and n3805_not n7632 ; n8843
g8780 nor n8842 n8843 ; n8844
g8781 and n8841_not n8844 ; n8845
g8782 and n7294_not n8845 ; n8846
g8783 and n4558_not n8845 ; n8847
g8784 nor n8846 n8847 ; n8848
g8785 and a[11] n8848_not ; n8849
g8786 and a[11]_not n8848 ; n8850
g8787 nor n8849 n8850 ; n8851
g8788 nor n8840 n8851 ; n8852
g8789 and n8840 n8851 ; n8853
g8790 nor n8852 n8853 ; n8854
g8791 and n8387 n8389_not ; n8855
g8792 nor n8390 n8855 ; n8856
g8793 and n8854 n8856 ; n8857
g8794 nor n8852 n8857 ; n8858
g8795 and n3877_not n8418 ; n8859
g8796 and n8410_not n8416 ; n8860
g8797 and n4515_not n8860 ; n8861
g8798 nor n8859 n8861 ; n8862
g8799 and n8421_not n8862 ; n8863
g8800 and n4609_not n8862 ; n8864
g8801 nor n8863 n8864 ; n8865
g8802 and a[8] n8865_not ; n8866
g8803 and a[8]_not n8865 ; n8867
g8804 nor n8866 n8867 ; n8868
g8805 nor n8858 n8868 ; n8869
g8806 and n8394 n8406_not ; n8870
g8807 nor n8405 n8406 ; n8871
g8808 nor n8870 n8871 ; n8872
g8809 and n8858 n8868 ; n8873
g8810 nor n8869 n8873 ; n8874
g8811 and n8872_not n8874 ; n8875
g8812 nor n8869 n8875 ; n8876
g8813 nor n8440 n8876 ; n8877
g8814 and n8440 n8876 ; n8878
g8815 nor n8877 n8878 ; n8879
g8816 and n8827 n8839_not ; n8880
g8817 nor n8838 n8839 ; n8881
g8818 nor n8880 n8881 ; n8882
g8819 and n8811 n8823_not ; n8883
g8820 nor n8822 n8823 ; n8884
g8821 nor n8883 n8884 ; n8885
g8822 and n958_not n6233 ; n8886
g8823 and n1178_not n5663 ; n8887
g8824 and n1060_not n5939 ; n8888
g8825 nor n8887 n8888 ; n8889
g8826 and n8886_not n8889 ; n8890
g8827 and n4633 n5666 ; n8891
g8828 and n8890 n8891_not ; n8892
g8829 and a[17] n8892_not ; n8893
g8830 nor n8892 n8893 ; n8894
g8831 and a[17] n8893_not ; n8895
g8832 nor n8894 n8895 ; n8896
g8833 nor n8785 n8789 ; n8897
g8834 nor n8788 n8789 ; n8898
g8835 nor n8897 n8898 ; n8899
g8836 nor n8896 n8899 ; n8900
g8837 nor n8896 n8900 ; n8901
g8838 nor n8899 n8900 ; n8902
g8839 nor n8901 n8902 ; n8903
g8840 and n1060_not n6233 ; n8904
g8841 and n1235_not n5663 ; n8905
g8842 and n1178_not n5939 ; n8906
g8843 nor n8905 n8906 ; n8907
g8844 and n8904_not n8907 ; n8908
g8845 and n4429 n5666 ; n8909
g8846 and n8908 n8909_not ; n8910
g8847 and a[17] n8910_not ; n8911
g8848 nor n8910 n8911 ; n8912
g8849 and a[17] n8911_not ; n8913
g8850 nor n8912 n8913 ; n8914
g8851 nor n8780 n8784 ; n8915
g8852 nor n8783 n8784 ; n8916
g8853 nor n8915 n8916 ; n8917
g8854 nor n8914 n8917 ; n8918
g8855 nor n8914 n8918 ; n8919
g8856 nor n8917 n8918 ; n8920
g8857 nor n8919 n8920 ; n8921
g8858 and n1178_not n6233 ; n8922
g8859 and n1364_not n5663 ; n8923
g8860 and n1235_not n5939 ; n8924
g8861 nor n8923 n8924 ; n8925
g8862 and n8922_not n8925 ; n8926
g8863 and n4861 n5666 ; n8927
g8864 and n8926 n8927_not ; n8928
g8865 and a[17] n8928_not ; n8929
g8866 nor n8928 n8929 ; n8930
g8867 and a[17] n8929_not ; n8931
g8868 nor n8930 n8931 ; n8932
g8869 nor n8775 n8779 ; n8933
g8870 nor n8778 n8779 ; n8934
g8871 nor n8933 n8934 ; n8935
g8872 nor n8932 n8935 ; n8936
g8873 nor n8932 n8936 ; n8937
g8874 nor n8935 n8936 ; n8938
g8875 nor n8937 n8938 ; n8939
g8876 and n1235_not n6233 ; n8940
g8877 and n1472_not n5663 ; n8941
g8878 and n1364_not n5939 ; n8942
g8879 nor n8941 n8942 ; n8943
g8880 and n8940_not n8943 ; n8944
g8881 and n4848 n5666 ; n8945
g8882 and n8944 n8945_not ; n8946
g8883 and a[17] n8946_not ; n8947
g8884 nor n8946 n8947 ; n8948
g8885 and a[17] n8947_not ; n8949
g8886 nor n8948 n8949 ; n8950
g8887 nor n8770 n8774 ; n8951
g8888 nor n8773 n8774 ; n8952
g8889 nor n8951 n8952 ; n8953
g8890 nor n8950 n8953 ; n8954
g8891 nor n8950 n8954 ; n8955
g8892 nor n8953 n8954 ; n8956
g8893 nor n8955 n8956 ; n8957
g8894 and n1364_not n6233 ; n8958
g8895 and n1572_not n5663 ; n8959
g8896 and n1472_not n5939 ; n8960
g8897 nor n8959 n8960 ; n8961
g8898 and n8958_not n8961 ; n8962
g8899 and n5114 n5666 ; n8963
g8900 and n8962 n8963_not ; n8964
g8901 and a[17] n8964_not ; n8965
g8902 nor n8964 n8965 ; n8966
g8903 and a[17] n8965_not ; n8967
g8904 nor n8966 n8967 ; n8968
g8905 nor n8765 n8769 ; n8969
g8906 nor n8768 n8769 ; n8970
g8907 nor n8969 n8970 ; n8971
g8908 nor n8968 n8971 ; n8972
g8909 nor n8968 n8972 ; n8973
g8910 nor n8971 n8972 ; n8974
g8911 nor n8973 n8974 ; n8975
g8912 and n1472_not n6233 ; n8976
g8913 and n1665_not n5663 ; n8977
g8914 and n1572_not n5939 ; n8978
g8915 nor n8977 n8978 ; n8979
g8916 and n8976_not n8979 ; n8980
g8917 and n5139 n5666 ; n8981
g8918 and n8980 n8981_not ; n8982
g8919 and a[17] n8982_not ; n8983
g8920 nor n8982 n8983 ; n8984
g8921 and a[17] n8983_not ; n8985
g8922 nor n8984 n8985 ; n8986
g8923 nor n8760 n8764 ; n8987
g8924 nor n8763 n8764 ; n8988
g8925 nor n8987 n8988 ; n8989
g8926 nor n8986 n8989 ; n8990
g8927 nor n8986 n8990 ; n8991
g8928 nor n8989 n8990 ; n8992
g8929 nor n8991 n8992 ; n8993
g8930 and n1572_not n6233 ; n8994
g8931 and n1779_not n5663 ; n8995
g8932 and n1665_not n5939 ; n8996
g8933 nor n8995 n8996 ; n8997
g8934 and n8994_not n8997 ; n8998
g8935 and n5561 n5666 ; n8999
g8936 and n8998 n8999_not ; n9000
g8937 and a[17] n9000_not ; n9001
g8938 nor n9000 n9001 ; n9002
g8939 and a[17] n9001_not ; n9003
g8940 nor n9002 n9003 ; n9004
g8941 nor n8755 n8759 ; n9005
g8942 nor n8758 n8759 ; n9006
g8943 nor n9005 n9006 ; n9007
g8944 nor n9004 n9007 ; n9008
g8945 nor n9004 n9008 ; n9009
g8946 nor n9007 n9008 ; n9010
g8947 nor n9009 n9010 ; n9011
g8948 and n8561 n8753 ; n9012
g8949 nor n8754 n9012 ; n9013
g8950 and n1665_not n6233 ; n9014
g8951 and n1877_not n5663 ; n9015
g8952 and n1779_not n5939 ; n9016
g8953 nor n9015 n9016 ; n9017
g8954 and n9014_not n9017 ; n9018
g8955 and n5666_not n9018 ; n9019
g8956 and n5328_not n9018 ; n9020
g8957 nor n9019 n9020 ; n9021
g8958 and a[17] n9021_not ; n9022
g8959 and a[17]_not n9021 ; n9023
g8960 nor n9022 n9023 ; n9024
g8961 and n9013 n9024_not ; n9025
g8962 and n8579 n8751 ; n9026
g8963 nor n8752 n9026 ; n9027
g8964 and n1779_not n6233 ; n9028
g8965 and n1913_not n5663 ; n9029
g8966 and n1877_not n5939 ; n9030
g8967 nor n9029 n9030 ; n9031
g8968 and n9028_not n9031 ; n9032
g8969 and n5666_not n9032 ; n9033
g8970 and n5851_not n9032 ; n9034
g8971 nor n9033 n9034 ; n9035
g8972 and a[17] n9035_not ; n9036
g8973 and a[17]_not n9035 ; n9037
g8974 nor n9036 n9037 ; n9038
g8975 and n9027 n9038_not ; n9039
g8976 and n1877_not n6233 ; n9040
g8977 and n1992_not n5663 ; n9041
g8978 and n1913_not n5939 ; n9042
g8979 nor n9041 n9042 ; n9043
g8980 and n9040_not n9043 ; n9044
g8981 and n5666 n6007 ; n9045
g8982 and n9044 n9045_not ; n9046
g8983 and a[17] n9046_not ; n9047
g8984 nor n9046 n9047 ; n9048
g8985 and a[17] n9047_not ; n9049
g8986 nor n9048 n9049 ; n9050
g8987 and n8747 n8749_not ; n9051
g8988 nor n8750 n9051 ; n9052
g8989 and n9050_not n9052 ; n9053
g8990 nor n9050 n9053 ; n9054
g8991 and n9052 n9053_not ; n9055
g8992 nor n9054 n9055 ; n9056
g8993 and n1913_not n6233 ; n9057
g8994 and n2057_not n5663 ; n9058
g8995 and n1992_not n5939 ; n9059
g8996 nor n9058 n9059 ; n9060
g8997 and n9057_not n9060 ; n9061
g8998 and n5666 n5834 ; n9062
g8999 and n9061 n9062_not ; n9063
g9000 and a[17] n9063_not ; n9064
g9001 nor n9063 n9064 ; n9065
g9002 and a[17] n9064_not ; n9066
g9003 nor n9065 n9066 ; n9067
g9004 nor n8742 n8746 ; n9068
g9005 nor n8745 n8746 ; n9069
g9006 nor n9068 n9069 ; n9070
g9007 nor n9067 n9070 ; n9071
g9008 nor n9067 n9071 ; n9072
g9009 nor n9070 n9071 ; n9073
g9010 nor n9072 n9073 ; n9074
g9011 and n1992_not n6233 ; n9075
g9012 and n2152_not n5663 ; n9076
g9013 and n2057_not n5939 ; n9077
g9014 nor n9076 n9077 ; n9078
g9015 and n9075_not n9078 ; n9079
g9016 and n5666 n6143 ; n9080
g9017 and n9079 n9080_not ; n9081
g9018 and a[17] n9081_not ; n9082
g9019 nor n9081 n9082 ; n9083
g9020 and a[17] n9082_not ; n9084
g9021 nor n9083 n9084 ; n9085
g9022 nor n8737 n8741 ; n9086
g9023 nor n8740 n8741 ; n9087
g9024 nor n9086 n9087 ; n9088
g9025 nor n9085 n9088 ; n9089
g9026 nor n9085 n9089 ; n9090
g9027 nor n9088 n9089 ; n9091
g9028 nor n9090 n9091 ; n9092
g9029 and n8638 n8735 ; n9093
g9030 nor n8736 n9093 ; n9094
g9031 and n2057_not n6233 ; n9095
g9032 and n2189_not n5663 ; n9096
g9033 and n2152_not n5939 ; n9097
g9034 nor n9096 n9097 ; n9098
g9035 and n9095_not n9098 ; n9099
g9036 and n5666_not n9099 ; n9100
g9037 and n6479_not n9099 ; n9101
g9038 nor n9100 n9101 ; n9102
g9039 and a[17] n9102_not ; n9103
g9040 and a[17]_not n9102 ; n9104
g9041 nor n9103 n9104 ; n9105
g9042 and n9094 n9105_not ; n9106
g9043 and n8731 n8733_not ; n9107
g9044 nor n8734 n9107 ; n9108
g9045 and n2152_not n6233 ; n9109
g9046 and n2291_not n5663 ; n9110
g9047 and n2189_not n5939 ; n9111
g9048 nor n9110 n9111 ; n9112
g9049 and n9109_not n9112 ; n9113
g9050 and n5666_not n9113 ; n9114
g9051 and n6492_not n9113 ; n9115
g9052 nor n9114 n9115 ; n9116
g9053 and a[17] n9116_not ; n9117
g9054 and a[17]_not n9116 ; n9118
g9055 nor n9117 n9118 ; n9119
g9056 and n9108 n9119_not ; n9120
g9057 and n8670 n8729 ; n9121
g9058 nor n8730 n9121 ; n9122
g9059 and n2189_not n6233 ; n9123
g9060 and n2388_not n5663 ; n9124
g9061 and n2291_not n5939 ; n9125
g9062 nor n9124 n9125 ; n9126
g9063 and n9123_not n9126 ; n9127
g9064 and n5666_not n9127 ; n9128
g9065 and n6122_not n9127 ; n9129
g9066 nor n9128 n9129 ; n9130
g9067 and a[17] n9130_not ; n9131
g9068 and a[17]_not n9130 ; n9132
g9069 nor n9131 n9132 ; n9133
g9070 and n9122 n9133_not ; n9134
g9071 and n2291_not n6233 ; n9135
g9072 and n2464_not n5663 ; n9136
g9073 and n2388_not n5939 ; n9137
g9074 nor n9136 n9137 ; n9138
g9075 and n9135_not n9138 ; n9139
g9076 and n5666 n6541 ; n9140
g9077 and n9139 n9140_not ; n9141
g9078 and a[17] n9141_not ; n9142
g9079 nor n9141 n9142 ; n9143
g9080 and a[17] n9142_not ; n9144
g9081 nor n9143 n9144 ; n9145
g9082 and n8725 n8727_not ; n9146
g9083 nor n8728 n9146 ; n9147
g9084 and n9145_not n9147 ; n9148
g9085 nor n9145 n9148 ; n9149
g9086 and n9147 n9148_not ; n9150
g9087 nor n9149 n9150 ; n9151
g9088 nor n8712 n8724 ; n9152
g9089 nor n8723 n8724 ; n9153
g9090 nor n9152 n9153 ; n9154
g9091 and n2388_not n6233 ; n9155
g9092 and n2533_not n5663 ; n9156
g9093 and n2464_not n5939 ; n9157
g9094 nor n9156 n9157 ; n9158
g9095 and n9155_not n9158 ; n9159
g9096 and n5666_not n9159 ; n9160
g9097 and n6591_not n9159 ; n9161
g9098 nor n9160 n9161 ; n9162
g9099 and a[17] n9162_not ; n9163
g9100 and a[17]_not n9162 ; n9164
g9101 nor n9163 n9164 ; n9165
g9102 nor n9154 n9165 ; n9166
g9103 and n2464_not n6233 ; n9167
g9104 and n2571_not n5663 ; n9168
g9105 and n2533_not n5939 ; n9169
g9106 nor n9168 n9169 ; n9170
g9107 and n9167_not n9170 ; n9171
g9108 and n5666 n6646 ; n9172
g9109 and n9171 n9172_not ; n9173
g9110 and a[17] n9173_not ; n9174
g9111 nor n9173 n9174 ; n9175
g9112 and a[17] n9174_not ; n9176
g9113 nor n9175 n9176 ; n9177
g9114 and n8696_not n8707 ; n9178
g9115 nor n8708 n9178 ; n9179
g9116 and n9177_not n9179 ; n9180
g9117 nor n9177 n9180 ; n9181
g9118 and n9179 n9180_not ; n9182
g9119 nor n9181 n9182 ; n9183
g9120 and n8693 n8695_not ; n9184
g9121 nor n8696 n9184 ; n9185
g9122 and n2533_not n6233 ; n9186
g9123 and n2674_not n5663 ; n9187
g9124 and n2571_not n5939 ; n9188
g9125 nor n9187 n9188 ; n9189
g9126 and n9186_not n9189 ; n9190
g9127 and n5666_not n9190 ; n9191
g9128 and n6695_not n9190 ; n9192
g9129 nor n9191 n9192 ; n9193
g9130 and a[17] n9193_not ; n9194
g9131 and a[17]_not n9193 ; n9195
g9132 nor n9194 n9195 ; n9196
g9133 and n9185 n9196_not ; n9197
g9134 and n2829_not n5939 ; n9198
g9135 and n2736_not n6233 ; n9199
g9136 nor n9198 n9199 ; n9200
g9137 and n5666 n7469_not ; n9201
g9138 and n9200 n9201_not ; n9202
g9139 and a[17] n9202_not ; n9203
g9140 and a[17] n9203_not ; n9204
g9141 nor n9202 n9203 ; n9205
g9142 nor n9204 n9205 ; n9206
g9143 nor n2829 n5658 ; n9207
g9144 and a[17] n9207_not ; n9208
g9145 and n9206_not n9208 ; n9209
g9146 and n2674_not n6233 ; n9210
g9147 and n2829_not n5663 ; n9211
g9148 and n2736_not n5939 ; n9212
g9149 nor n9211 n9212 ; n9213
g9150 and n9210_not n9213 ; n9214
g9151 and n5666_not n9214 ; n9215
g9152 and n6798_not n9214 ; n9216
g9153 nor n9215 n9216 ; n9217
g9154 and a[17] n9217_not ; n9218
g9155 and a[17]_not n9217 ; n9219
g9156 nor n9218 n9219 ; n9220
g9157 and n9209 n9220_not ; n9221
g9158 and n8694 n9221 ; n9222
g9159 and n9221 n9222_not ; n9223
g9160 and n8694 n9222_not ; n9224
g9161 nor n9223 n9224 ; n9225
g9162 and n2571_not n6233 ; n9226
g9163 and n2736_not n5663 ; n9227
g9164 and n2674_not n5939 ; n9228
g9165 nor n9227 n9228 ; n9229
g9166 and n9226_not n9229 ; n9230
g9167 and n5666 n6806 ; n9231
g9168 and n9230 n9231_not ; n9232
g9169 and a[17] n9232_not ; n9233
g9170 and a[17] n9233_not ; n9234
g9171 nor n9232 n9233 ; n9235
g9172 nor n9234 n9235 ; n9236
g9173 nor n9225 n9236 ; n9237
g9174 nor n9222 n9237 ; n9238
g9175 and n9185_not n9196 ; n9239
g9176 nor n9197 n9239 ; n9240
g9177 and n9238_not n9240 ; n9241
g9178 nor n9197 n9241 ; n9242
g9179 nor n9183 n9242 ; n9243
g9180 nor n9180 n9243 ; n9244
g9181 and n9154 n9165 ; n9245
g9182 nor n9166 n9245 ; n9246
g9183 and n9244_not n9246 ; n9247
g9184 nor n9166 n9247 ; n9248
g9185 nor n9151 n9248 ; n9249
g9186 nor n9148 n9249 ; n9250
g9187 and n9122 n9134_not ; n9251
g9188 nor n9133 n9134 ; n9252
g9189 nor n9251 n9252 ; n9253
g9190 nor n9250 n9253 ; n9254
g9191 nor n9134 n9254 ; n9255
g9192 and n9108 n9120_not ; n9256
g9193 nor n9119 n9120 ; n9257
g9194 nor n9256 n9257 ; n9258
g9195 nor n9255 n9258 ; n9259
g9196 nor n9120 n9259 ; n9260
g9197 and n9094_not n9105 ; n9261
g9198 nor n9106 n9261 ; n9262
g9199 and n9260_not n9262 ; n9263
g9200 nor n9106 n9263 ; n9264
g9201 nor n9092 n9264 ; n9265
g9202 nor n9089 n9265 ; n9266
g9203 nor n9074 n9266 ; n9267
g9204 nor n9071 n9267 ; n9268
g9205 nor n9056 n9268 ; n9269
g9206 nor n9053 n9269 ; n9270
g9207 and n9027 n9039_not ; n9271
g9208 nor n9038 n9039 ; n9272
g9209 nor n9271 n9272 ; n9273
g9210 nor n9270 n9273 ; n9274
g9211 nor n9039 n9274 ; n9275
g9212 and n9013_not n9024 ; n9276
g9213 nor n9025 n9276 ; n9277
g9214 and n9275_not n9277 ; n9278
g9215 nor n9025 n9278 ; n9279
g9216 nor n9011 n9279 ; n9280
g9217 nor n9008 n9280 ; n9281
g9218 nor n8993 n9281 ; n9282
g9219 nor n8990 n9282 ; n9283
g9220 nor n8975 n9283 ; n9284
g9221 nor n8972 n9284 ; n9285
g9222 nor n8957 n9285 ; n9286
g9223 nor n8954 n9286 ; n9287
g9224 nor n8939 n9287 ; n9288
g9225 nor n8936 n9288 ; n9289
g9226 nor n8921 n9289 ; n9290
g9227 nor n8918 n9290 ; n9291
g9228 nor n8903 n9291 ; n9292
g9229 nor n8900 n9292 ; n9293
g9230 and n8804 n8806_not ; n9294
g9231 nor n8807 n9294 ; n9295
g9232 and n9293_not n9295 ; n9296
g9233 and n392_not n7101 ; n9297
g9234 and n710_not n6402 ; n9298
g9235 and n587_not n6951 ; n9299
g9236 nor n9298 n9299 ; n9300
g9237 and n9297_not n9300 ; n9301
g9238 and n3347 n6397 ; n9302
g9239 and n9301 n9302_not ; n9303
g9240 and a[14] n9303_not ; n9304
g9241 nor n9303 n9304 ; n9305
g9242 and a[14] n9304_not ; n9306
g9243 nor n9305 n9306 ; n9307
g9244 and n9293 n9295_not ; n9308
g9245 nor n9296 n9308 ; n9309
g9246 and n9307_not n9309 ; n9310
g9247 nor n9296 n9310 ; n9311
g9248 nor n8885 n9311 ; n9312
g9249 and n8885 n9311 ; n9313
g9250 nor n9312 n9313 ; n9314
g9251 and n3456_not n7983 ; n9315
g9252 and n3539_not n7291 ; n9316
g9253 and n3605_not n7632 ; n9317
g9254 nor n9316 n9317 ; n9318
g9255 and n9315_not n9318 ; n9319
g9256 and n3627 n7294 ; n9320
g9257 and n9319 n9320_not ; n9321
g9258 and a[11] n9321_not ; n9322
g9259 and a[11] n9322_not ; n9323
g9260 nor n9321 n9322 ; n9324
g9261 nor n9323 n9324 ; n9325
g9262 and n9314 n9325_not ; n9326
g9263 nor n9312 n9326 ; n9327
g9264 nor n8882 n9327 ; n9328
g9265 and n8882 n9327 ; n9329
g9266 nor n9328 n9329 ; n9330
g9267 and n8413 n8416_not ; n9331
g9268 and n3877_not n9331 ; n9332
g9269 and n3964_not n8418 ; n9333
g9270 and n4045_not n8860 ; n9334
g9271 nor n9333 n9334 ; n9335
g9272 and n9332_not n9335 ; n9336
g9273 and n4067 n8421 ; n9337
g9274 and n9336 n9337_not ; n9338
g9275 and a[8] n9338_not ; n9339
g9276 and a[8] n9339_not ; n9340
g9277 nor n9338 n9339 ; n9341
g9278 nor n9340 n9341 ; n9342
g9279 and n9330 n9342_not ; n9343
g9280 nor n9328 n9343 ; n9344
g9281 and n4515_not n9331 ; n9345
g9282 and n4045_not n8418 ; n9346
g9283 and n3877_not n8860 ; n9347
g9284 nor n9346 n9347 ; n9348
g9285 and n9345_not n9348 ; n9349
g9286 and n8421_not n9349 ; n9350
g9287 and n4715_not n9349 ; n9351
g9288 nor n9350 n9351 ; n9352
g9289 and a[8] n9352_not ; n9353
g9290 and a[8]_not n9352 ; n9354
g9291 nor n9353 n9354 ; n9355
g9292 nor n9344 n9355 ; n9356
g9293 nor n9344 n9356 ; n9357
g9294 nor n9355 n9356 ; n9358
g9295 nor n9357 n9358 ; n9359
g9296 nor n8854 n8856 ; n9360
g9297 nor n8857 n9360 ; n9361
g9298 and n9359_not n9361 ; n9362
g9299 nor n9356 n9362 ; n9363
g9300 and n8872 n8874_not ; n9364
g9301 nor n8875 n9364 ; n9365
g9302 and n9363_not n9365 ; n9366
g9303 and n9314 n9326_not ; n9367
g9304 nor n9325 n9326 ; n9368
g9305 nor n9367 n9368 ; n9369
g9306 and n8903 n9291 ; n9370
g9307 nor n9292 n9370 ; n9371
g9308 and n587_not n7101 ; n9372
g9309 and n867_not n6402 ; n9373
g9310 and n710_not n6951 ; n9374
g9311 nor n9373 n9374 ; n9375
g9312 and n9372_not n9375 ; n9376
g9313 and n6397_not n9376 ; n9377
g9314 and n3331_not n9376 ; n9378
g9315 nor n9377 n9378 ; n9379
g9316 and a[14] n9379_not ; n9380
g9317 and a[14]_not n9379 ; n9381
g9318 nor n9380 n9381 ; n9382
g9319 and n9371 n9382_not ; n9383
g9320 and n8921 n9289 ; n9384
g9321 nor n9290 n9384 ; n9385
g9322 and n710_not n7101 ; n9386
g9323 and n958_not n6402 ; n9387
g9324 and n867_not n6951 ; n9388
g9325 nor n9387 n9388 ; n9389
g9326 and n9386_not n9389 ; n9390
g9327 and n6397_not n9390 ; n9391
g9328 and n4179_not n9390 ; n9392
g9329 nor n9391 n9392 ; n9393
g9330 and a[14] n9393_not ; n9394
g9331 and a[14]_not n9393 ; n9395
g9332 nor n9394 n9395 ; n9396
g9333 and n9385 n9396_not ; n9397
g9334 and n8939 n9287 ; n9398
g9335 nor n9288 n9398 ; n9399
g9336 and n867_not n7101 ; n9400
g9337 and n1060_not n6402 ; n9401
g9338 and n958_not n6951 ; n9402
g9339 nor n9401 n9402 ; n9403
g9340 and n9400_not n9403 ; n9404
g9341 and n6397_not n9404 ; n9405
g9342 and n4204_not n9404 ; n9406
g9343 nor n9405 n9406 ; n9407
g9344 and a[14] n9407_not ; n9408
g9345 and a[14]_not n9407 ; n9409
g9346 nor n9408 n9409 ; n9410
g9347 and n9399 n9410_not ; n9411
g9348 and n8957 n9285 ; n9412
g9349 nor n9286 n9412 ; n9413
g9350 and n958_not n7101 ; n9414
g9351 and n1178_not n6402 ; n9415
g9352 and n1060_not n6951 ; n9416
g9353 nor n9415 n9416 ; n9417
g9354 and n9414_not n9417 ; n9418
g9355 and n6397_not n9418 ; n9419
g9356 and n4633_not n9418 ; n9420
g9357 nor n9419 n9420 ; n9421
g9358 and a[14] n9421_not ; n9422
g9359 and a[14]_not n9421 ; n9423
g9360 nor n9422 n9423 ; n9424
g9361 and n9413 n9424_not ; n9425
g9362 and n8975 n9283 ; n9426
g9363 nor n9284 n9426 ; n9427
g9364 and n1060_not n7101 ; n9428
g9365 and n1235_not n6402 ; n9429
g9366 and n1178_not n6951 ; n9430
g9367 nor n9429 n9430 ; n9431
g9368 and n9428_not n9431 ; n9432
g9369 and n6397_not n9432 ; n9433
g9370 and n4429_not n9432 ; n9434
g9371 nor n9433 n9434 ; n9435
g9372 and a[14] n9435_not ; n9436
g9373 and a[14]_not n9435 ; n9437
g9374 nor n9436 n9437 ; n9438
g9375 and n9427 n9438_not ; n9439
g9376 and n8993 n9281 ; n9440
g9377 nor n9282 n9440 ; n9441
g9378 and n1178_not n7101 ; n9442
g9379 and n1364_not n6402 ; n9443
g9380 and n1235_not n6951 ; n9444
g9381 nor n9443 n9444 ; n9445
g9382 and n9442_not n9445 ; n9446
g9383 and n6397_not n9446 ; n9447
g9384 and n4861_not n9446 ; n9448
g9385 nor n9447 n9448 ; n9449
g9386 and a[14] n9449_not ; n9450
g9387 and a[14]_not n9449 ; n9451
g9388 nor n9450 n9451 ; n9452
g9389 and n9441 n9452_not ; n9453
g9390 and n9011 n9279 ; n9454
g9391 nor n9280 n9454 ; n9455
g9392 and n1235_not n7101 ; n9456
g9393 and n1472_not n6402 ; n9457
g9394 and n1364_not n6951 ; n9458
g9395 nor n9457 n9458 ; n9459
g9396 and n9456_not n9459 ; n9460
g9397 and n6397_not n9460 ; n9461
g9398 and n4848_not n9460 ; n9462
g9399 nor n9461 n9462 ; n9463
g9400 and a[14] n9463_not ; n9464
g9401 and a[14]_not n9463 ; n9465
g9402 nor n9464 n9465 ; n9466
g9403 and n9455 n9466_not ; n9467
g9404 and n1364_not n7101 ; n9468
g9405 and n1572_not n6402 ; n9469
g9406 and n1472_not n6951 ; n9470
g9407 nor n9469 n9470 ; n9471
g9408 and n9468_not n9471 ; n9472
g9409 and n5114 n6397 ; n9473
g9410 and n9472 n9473_not ; n9474
g9411 and a[14] n9474_not ; n9475
g9412 nor n9474 n9475 ; n9476
g9413 and a[14] n9475_not ; n9477
g9414 nor n9476 n9477 ; n9478
g9415 and n9275 n9277_not ; n9479
g9416 nor n9278 n9479 ; n9480
g9417 and n9478_not n9480 ; n9481
g9418 nor n9478 n9481 ; n9482
g9419 and n9480 n9481_not ; n9483
g9420 nor n9482 n9483 ; n9484
g9421 and n1472_not n7101 ; n9485
g9422 and n1665_not n6402 ; n9486
g9423 and n1572_not n6951 ; n9487
g9424 nor n9486 n9487 ; n9488
g9425 and n9485_not n9488 ; n9489
g9426 and n5139 n6397 ; n9490
g9427 and n9489 n9490_not ; n9491
g9428 and a[14] n9491_not ; n9492
g9429 nor n9491 n9492 ; n9493
g9430 and a[14] n9492_not ; n9494
g9431 nor n9493 n9494 ; n9495
g9432 nor n9270 n9274 ; n9496
g9433 nor n9273 n9274 ; n9497
g9434 nor n9496 n9497 ; n9498
g9435 nor n9495 n9498 ; n9499
g9436 nor n9495 n9499 ; n9500
g9437 nor n9498 n9499 ; n9501
g9438 nor n9500 n9501 ; n9502
g9439 and n9056 n9268 ; n9503
g9440 nor n9269 n9503 ; n9504
g9441 and n1572_not n7101 ; n9505
g9442 and n1779_not n6402 ; n9506
g9443 and n1665_not n6951 ; n9507
g9444 nor n9506 n9507 ; n9508
g9445 and n9505_not n9508 ; n9509
g9446 and n6397_not n9509 ; n9510
g9447 and n5561_not n9509 ; n9511
g9448 nor n9510 n9511 ; n9512
g9449 and a[14] n9512_not ; n9513
g9450 and a[14]_not n9512 ; n9514
g9451 nor n9513 n9514 ; n9515
g9452 and n9504 n9515_not ; n9516
g9453 and n9074 n9266 ; n9517
g9454 nor n9267 n9517 ; n9518
g9455 and n1665_not n7101 ; n9519
g9456 and n1877_not n6402 ; n9520
g9457 and n1779_not n6951 ; n9521
g9458 nor n9520 n9521 ; n9522
g9459 and n9519_not n9522 ; n9523
g9460 and n6397_not n9523 ; n9524
g9461 and n5328_not n9523 ; n9525
g9462 nor n9524 n9525 ; n9526
g9463 and a[14] n9526_not ; n9527
g9464 and a[14]_not n9526 ; n9528
g9465 nor n9527 n9528 ; n9529
g9466 and n9518 n9529_not ; n9530
g9467 and n9092 n9264 ; n9531
g9468 nor n9265 n9531 ; n9532
g9469 and n1779_not n7101 ; n9533
g9470 and n1913_not n6402 ; n9534
g9471 and n1877_not n6951 ; n9535
g9472 nor n9534 n9535 ; n9536
g9473 and n9533_not n9536 ; n9537
g9474 and n6397_not n9537 ; n9538
g9475 and n5851_not n9537 ; n9539
g9476 nor n9538 n9539 ; n9540
g9477 and a[14] n9540_not ; n9541
g9478 and a[14]_not n9540 ; n9542
g9479 nor n9541 n9542 ; n9543
g9480 and n9532 n9543_not ; n9544
g9481 and n1877_not n7101 ; n9545
g9482 and n1992_not n6402 ; n9546
g9483 and n1913_not n6951 ; n9547
g9484 nor n9546 n9547 ; n9548
g9485 and n9545_not n9548 ; n9549
g9486 and n6007 n6397 ; n9550
g9487 and n9549 n9550_not ; n9551
g9488 and a[14] n9551_not ; n9552
g9489 nor n9551 n9552 ; n9553
g9490 and a[14] n9552_not ; n9554
g9491 nor n9553 n9554 ; n9555
g9492 and n9260 n9262_not ; n9556
g9493 nor n9263 n9556 ; n9557
g9494 and n9555_not n9557 ; n9558
g9495 nor n9555 n9558 ; n9559
g9496 and n9557 n9558_not ; n9560
g9497 nor n9559 n9560 ; n9561
g9498 and n1913_not n7101 ; n9562
g9499 and n2057_not n6402 ; n9563
g9500 and n1992_not n6951 ; n9564
g9501 nor n9563 n9564 ; n9565
g9502 and n9562_not n9565 ; n9566
g9503 and n5834 n6397 ; n9567
g9504 and n9566 n9567_not ; n9568
g9505 and a[14] n9568_not ; n9569
g9506 nor n9568 n9569 ; n9570
g9507 and a[14] n9569_not ; n9571
g9508 nor n9570 n9571 ; n9572
g9509 nor n9255 n9259 ; n9573
g9510 nor n9258 n9259 ; n9574
g9511 nor n9573 n9574 ; n9575
g9512 nor n9572 n9575 ; n9576
g9513 nor n9572 n9576 ; n9577
g9514 nor n9575 n9576 ; n9578
g9515 nor n9577 n9578 ; n9579
g9516 and n1992_not n7101 ; n9580
g9517 and n2152_not n6402 ; n9581
g9518 and n2057_not n6951 ; n9582
g9519 nor n9581 n9582 ; n9583
g9520 and n9580_not n9583 ; n9584
g9521 and n6143 n6397 ; n9585
g9522 and n9584 n9585_not ; n9586
g9523 and a[14] n9586_not ; n9587
g9524 nor n9586 n9587 ; n9588
g9525 and a[14] n9587_not ; n9589
g9526 nor n9588 n9589 ; n9590
g9527 nor n9250 n9254 ; n9591
g9528 nor n9253 n9254 ; n9592
g9529 nor n9591 n9592 ; n9593
g9530 nor n9590 n9593 ; n9594
g9531 nor n9590 n9594 ; n9595
g9532 nor n9593 n9594 ; n9596
g9533 nor n9595 n9596 ; n9597
g9534 and n9151 n9248 ; n9598
g9535 nor n9249 n9598 ; n9599
g9536 and n2057_not n7101 ; n9600
g9537 and n2189_not n6402 ; n9601
g9538 and n2152_not n6951 ; n9602
g9539 nor n9601 n9602 ; n9603
g9540 and n9600_not n9603 ; n9604
g9541 and n6397_not n9604 ; n9605
g9542 and n6479_not n9604 ; n9606
g9543 nor n9605 n9606 ; n9607
g9544 and a[14] n9607_not ; n9608
g9545 and a[14]_not n9607 ; n9609
g9546 nor n9608 n9609 ; n9610
g9547 and n9599 n9610_not ; n9611
g9548 and n9244 n9246_not ; n9612
g9549 nor n9247 n9612 ; n9613
g9550 and n2152_not n7101 ; n9614
g9551 and n2291_not n6402 ; n9615
g9552 and n2189_not n6951 ; n9616
g9553 nor n9615 n9616 ; n9617
g9554 and n9614_not n9617 ; n9618
g9555 and n6397_not n9618 ; n9619
g9556 and n6492_not n9618 ; n9620
g9557 nor n9619 n9620 ; n9621
g9558 and a[14] n9621_not ; n9622
g9559 and a[14]_not n9621 ; n9623
g9560 nor n9622 n9623 ; n9624
g9561 and n9613 n9624_not ; n9625
g9562 and n9183 n9242 ; n9626
g9563 nor n9243 n9626 ; n9627
g9564 and n2189_not n7101 ; n9628
g9565 and n2388_not n6402 ; n9629
g9566 and n2291_not n6951 ; n9630
g9567 nor n9629 n9630 ; n9631
g9568 and n9628_not n9631 ; n9632
g9569 and n6397_not n9632 ; n9633
g9570 and n6122_not n9632 ; n9634
g9571 nor n9633 n9634 ; n9635
g9572 and a[14] n9635_not ; n9636
g9573 and a[14]_not n9635 ; n9637
g9574 nor n9636 n9637 ; n9638
g9575 and n9627 n9638_not ; n9639
g9576 and n2291_not n7101 ; n9640
g9577 and n2464_not n6402 ; n9641
g9578 and n2388_not n6951 ; n9642
g9579 nor n9641 n9642 ; n9643
g9580 and n9640_not n9643 ; n9644
g9581 and n6397 n6541 ; n9645
g9582 and n9644 n9645_not ; n9646
g9583 and a[14] n9646_not ; n9647
g9584 nor n9646 n9647 ; n9648
g9585 and a[14] n9647_not ; n9649
g9586 nor n9648 n9649 ; n9650
g9587 and n9238 n9240_not ; n9651
g9588 nor n9241 n9651 ; n9652
g9589 and n9650_not n9652 ; n9653
g9590 nor n9650 n9653 ; n9654
g9591 and n9652 n9653_not ; n9655
g9592 nor n9654 n9655 ; n9656
g9593 nor n9225 n9237 ; n9657
g9594 nor n9236 n9237 ; n9658
g9595 nor n9657 n9658 ; n9659
g9596 and n2388_not n7101 ; n9660
g9597 and n2533_not n6402 ; n9661
g9598 and n2464_not n6951 ; n9662
g9599 nor n9661 n9662 ; n9663
g9600 and n9660_not n9663 ; n9664
g9601 and n6397_not n9664 ; n9665
g9602 and n6591_not n9664 ; n9666
g9603 nor n9665 n9666 ; n9667
g9604 and a[14] n9667_not ; n9668
g9605 and a[14]_not n9667 ; n9669
g9606 nor n9668 n9669 ; n9670
g9607 nor n9659 n9670 ; n9671
g9608 and n2464_not n7101 ; n9672
g9609 and n2571_not n6402 ; n9673
g9610 and n2533_not n6951 ; n9674
g9611 nor n9673 n9674 ; n9675
g9612 and n9672_not n9675 ; n9676
g9613 and n6397 n6646 ; n9677
g9614 and n9676 n9677_not ; n9678
g9615 and a[14] n9678_not ; n9679
g9616 nor n9678 n9679 ; n9680
g9617 and a[14] n9679_not ; n9681
g9618 nor n9680 n9681 ; n9682
g9619 and n9209_not n9220 ; n9683
g9620 nor n9221 n9683 ; n9684
g9621 and n9682_not n9684 ; n9685
g9622 nor n9682 n9685 ; n9686
g9623 and n9684 n9685_not ; n9687
g9624 nor n9686 n9687 ; n9688
g9625 and n9206 n9208_not ; n9689
g9626 nor n9209 n9689 ; n9690
g9627 and n2533_not n7101 ; n9691
g9628 and n2674_not n6402 ; n9692
g9629 and n2571_not n6951 ; n9693
g9630 nor n9692 n9693 ; n9694
g9631 and n9691_not n9694 ; n9695
g9632 and n6397_not n9695 ; n9696
g9633 and n6695_not n9695 ; n9697
g9634 nor n9696 n9697 ; n9698
g9635 and a[14] n9698_not ; n9699
g9636 and a[14]_not n9698 ; n9700
g9637 nor n9699 n9700 ; n9701
g9638 and n9690 n9701_not ; n9702
g9639 and n2829_not n6951 ; n9703
g9640 and n2736_not n7101 ; n9704
g9641 nor n9703 n9704 ; n9705
g9642 and n6397 n7469_not ; n9706
g9643 and n9705 n9706_not ; n9707
g9644 and a[14] n9707_not ; n9708
g9645 and a[14] n9708_not ; n9709
g9646 nor n9707 n9708 ; n9710
g9647 nor n9709 n9710 ; n9711
g9648 nor n2829 n6393 ; n9712
g9649 and a[14] n9712_not ; n9713
g9650 and n9711_not n9713 ; n9714
g9651 and n2674_not n7101 ; n9715
g9652 and n2829_not n6402 ; n9716
g9653 and n2736_not n6951 ; n9717
g9654 nor n9716 n9717 ; n9718
g9655 and n9715_not n9718 ; n9719
g9656 and n6397_not n9719 ; n9720
g9657 and n6798_not n9719 ; n9721
g9658 nor n9720 n9721 ; n9722
g9659 and a[14] n9722_not ; n9723
g9660 and a[14]_not n9722 ; n9724
g9661 nor n9723 n9724 ; n9725
g9662 and n9714 n9725_not ; n9726
g9663 and n9207 n9726 ; n9727
g9664 and n9726 n9727_not ; n9728
g9665 and n9207 n9727_not ; n9729
g9666 nor n9728 n9729 ; n9730
g9667 and n2571_not n7101 ; n9731
g9668 and n2736_not n6402 ; n9732
g9669 and n2674_not n6951 ; n9733
g9670 nor n9732 n9733 ; n9734
g9671 and n9731_not n9734 ; n9735
g9672 and n6397 n6806 ; n9736
g9673 and n9735 n9736_not ; n9737
g9674 and a[14] n9737_not ; n9738
g9675 and a[14] n9738_not ; n9739
g9676 nor n9737 n9738 ; n9740
g9677 nor n9739 n9740 ; n9741
g9678 nor n9730 n9741 ; n9742
g9679 nor n9727 n9742 ; n9743
g9680 and n9690_not n9701 ; n9744
g9681 nor n9702 n9744 ; n9745
g9682 and n9743_not n9745 ; n9746
g9683 nor n9702 n9746 ; n9747
g9684 nor n9688 n9747 ; n9748
g9685 nor n9685 n9748 ; n9749
g9686 and n9659 n9670 ; n9750
g9687 nor n9671 n9750 ; n9751
g9688 and n9749_not n9751 ; n9752
g9689 nor n9671 n9752 ; n9753
g9690 nor n9656 n9753 ; n9754
g9691 nor n9653 n9754 ; n9755
g9692 and n9627 n9639_not ; n9756
g9693 nor n9638 n9639 ; n9757
g9694 nor n9756 n9757 ; n9758
g9695 nor n9755 n9758 ; n9759
g9696 nor n9639 n9759 ; n9760
g9697 and n9613 n9625_not ; n9761
g9698 nor n9624 n9625 ; n9762
g9699 nor n9761 n9762 ; n9763
g9700 nor n9760 n9763 ; n9764
g9701 nor n9625 n9764 ; n9765
g9702 and n9599_not n9610 ; n9766
g9703 nor n9611 n9766 ; n9767
g9704 and n9765_not n9767 ; n9768
g9705 nor n9611 n9768 ; n9769
g9706 nor n9597 n9769 ; n9770
g9707 nor n9594 n9770 ; n9771
g9708 nor n9579 n9771 ; n9772
g9709 nor n9576 n9772 ; n9773
g9710 nor n9561 n9773 ; n9774
g9711 nor n9558 n9774 ; n9775
g9712 and n9532 n9544_not ; n9776
g9713 nor n9543 n9544 ; n9777
g9714 nor n9776 n9777 ; n9778
g9715 nor n9775 n9778 ; n9779
g9716 nor n9544 n9779 ; n9780
g9717 and n9518 n9530_not ; n9781
g9718 nor n9529 n9530 ; n9782
g9719 nor n9781 n9782 ; n9783
g9720 nor n9780 n9783 ; n9784
g9721 nor n9530 n9784 ; n9785
g9722 and n9504_not n9515 ; n9786
g9723 nor n9516 n9786 ; n9787
g9724 and n9785_not n9787 ; n9788
g9725 nor n9516 n9788 ; n9789
g9726 nor n9502 n9789 ; n9790
g9727 nor n9499 n9790 ; n9791
g9728 nor n9484 n9791 ; n9792
g9729 nor n9481 n9792 ; n9793
g9730 and n9455 n9467_not ; n9794
g9731 nor n9466 n9467 ; n9795
g9732 nor n9794 n9795 ; n9796
g9733 nor n9793 n9796 ; n9797
g9734 nor n9467 n9797 ; n9798
g9735 and n9441 n9453_not ; n9799
g9736 nor n9452 n9453 ; n9800
g9737 nor n9799 n9800 ; n9801
g9738 nor n9798 n9801 ; n9802
g9739 nor n9453 n9802 ; n9803
g9740 and n9427 n9439_not ; n9804
g9741 nor n9438 n9439 ; n9805
g9742 nor n9804 n9805 ; n9806
g9743 nor n9803 n9806 ; n9807
g9744 nor n9439 n9807 ; n9808
g9745 and n9413 n9425_not ; n9809
g9746 nor n9424 n9425 ; n9810
g9747 nor n9809 n9810 ; n9811
g9748 nor n9808 n9811 ; n9812
g9749 nor n9425 n9812 ; n9813
g9750 and n9399 n9411_not ; n9814
g9751 nor n9410 n9411 ; n9815
g9752 nor n9814 n9815 ; n9816
g9753 nor n9813 n9816 ; n9817
g9754 nor n9411 n9817 ; n9818
g9755 and n9385 n9397_not ; n9819
g9756 nor n9396 n9397 ; n9820
g9757 nor n9819 n9820 ; n9821
g9758 nor n9818 n9821 ; n9822
g9759 nor n9397 n9822 ; n9823
g9760 and n9371 n9383_not ; n9824
g9761 nor n9382 n9383 ; n9825
g9762 nor n9824 n9825 ; n9826
g9763 nor n9823 n9826 ; n9827
g9764 nor n9383 n9827 ; n9828
g9765 and n9307 n9309_not ; n9829
g9766 nor n9310 n9829 ; n9830
g9767 and n9828_not n9830 ; n9831
g9768 and n3605_not n7983 ; n9832
g9769 and n3012_not n7291 ; n9833
g9770 and n3539_not n7632 ; n9834
g9771 nor n9833 n9834 ; n9835
g9772 and n9832_not n9835 ; n9836
g9773 and n4084 n7294 ; n9837
g9774 and n9836 n9837_not ; n9838
g9775 and a[11] n9838_not ; n9839
g9776 nor n9838 n9839 ; n9840
g9777 and a[11] n9839_not ; n9841
g9778 nor n9840 n9841 ; n9842
g9779 and n9828 n9830_not ; n9843
g9780 nor n9831 n9843 ; n9844
g9781 and n9842_not n9844 ; n9845
g9782 nor n9831 n9845 ; n9846
g9783 nor n9369 n9846 ; n9847
g9784 and n9369 n9846 ; n9848
g9785 nor n9847 n9848 ; n9849
g9786 and n4045_not n9331 ; n9850
g9787 and n3805_not n8418 ; n9851
g9788 and n3964_not n8860 ; n9852
g9789 nor n9851 n9852 ; n9853
g9790 and n9850_not n9853 ; n9854
g9791 and n4477 n8421 ; n9855
g9792 and n9854 n9855_not ; n9856
g9793 and a[8] n9856_not ; n9857
g9794 and a[8] n9857_not ; n9858
g9795 nor n9856 n9857 ; n9859
g9796 nor n9858 n9859 ; n9860
g9797 and n9849 n9860_not ; n9861
g9798 nor n9847 n9861 ; n9862
g9799 and a[3]_not a[4] ; n9863
g9800 and a[3] a[4]_not ; n9864
g9801 nor n9863 n9864 ; n9865
g9802 and n67_not n70 ; n9866
g9803 and n9865 n9866 ; n9867
g9804 and n4515_not n9867 ; n9868
g9805 nor n4522 n9868 ; n9869
g9806 nor n67 n70 ; n9870
g9807 nor n9868 n9870 ; n9871
g9808 nor n9869 n9871 ; n9872
g9809 and a[5] n9872_not ; n9873
g9810 and a[5]_not n9872 ; n9874
g9811 nor n9873 n9874 ; n9875
g9812 nor n9862 n9875 ; n9876
g9813 and n9330 n9343_not ; n9877
g9814 nor n9342 n9343 ; n9878
g9815 nor n9877 n9878 ; n9879
g9816 and n9862 n9875 ; n9880
g9817 nor n9876 n9880 ; n9881
g9818 and n9879_not n9881 ; n9882
g9819 nor n9876 n9882 ; n9883
g9820 nor n9358 n9361 ; n9884
g9821 and n9357_not n9884 ; n9885
g9822 nor n9362 n9885 ; n9886
g9823 and n9883_not n9886 ; n9887
g9824 nor n9879 n9882 ; n9888
g9825 and n9881 n9882_not ; n9889
g9826 nor n9888 n9889 ; n9890
g9827 and n3539_not n7983 ; n9891
g9828 and n392_not n7291 ; n9892
g9829 and n3012_not n7632 ; n9893
g9830 nor n9892 n9893 ; n9894
g9831 and n9891_not n9894 ; n9895
g9832 and n3715 n7294 ; n9896
g9833 and n9895 n9896_not ; n9897
g9834 and a[11] n9897_not ; n9898
g9835 nor n9897 n9898 ; n9899
g9836 and a[11] n9898_not ; n9900
g9837 nor n9899 n9900 ; n9901
g9838 nor n9823 n9827 ; n9902
g9839 nor n9826 n9827 ; n9903
g9840 nor n9902 n9903 ; n9904
g9841 nor n9901 n9904 ; n9905
g9842 nor n9901 n9905 ; n9906
g9843 nor n9904 n9905 ; n9907
g9844 nor n9906 n9907 ; n9908
g9845 and n3012_not n7983 ; n9909
g9846 and n587_not n7291 ; n9910
g9847 and n392_not n7632 ; n9911
g9848 nor n9910 n9911 ; n9912
g9849 and n9909_not n9912 ; n9913
g9850 and n3018 n7294 ; n9914
g9851 and n9913 n9914_not ; n9915
g9852 and a[11] n9915_not ; n9916
g9853 nor n9915 n9916 ; n9917
g9854 and a[11] n9916_not ; n9918
g9855 nor n9917 n9918 ; n9919
g9856 nor n9818 n9822 ; n9920
g9857 nor n9821 n9822 ; n9921
g9858 nor n9920 n9921 ; n9922
g9859 nor n9919 n9922 ; n9923
g9860 nor n9919 n9923 ; n9924
g9861 nor n9922 n9923 ; n9925
g9862 nor n9924 n9925 ; n9926
g9863 and n392_not n7983 ; n9927
g9864 and n710_not n7291 ; n9928
g9865 and n587_not n7632 ; n9929
g9866 nor n9928 n9929 ; n9930
g9867 and n9927_not n9930 ; n9931
g9868 and n3347 n7294 ; n9932
g9869 and n9931 n9932_not ; n9933
g9870 and a[11] n9933_not ; n9934
g9871 nor n9933 n9934 ; n9935
g9872 and a[11] n9934_not ; n9936
g9873 nor n9935 n9936 ; n9937
g9874 nor n9813 n9817 ; n9938
g9875 nor n9816 n9817 ; n9939
g9876 nor n9938 n9939 ; n9940
g9877 nor n9937 n9940 ; n9941
g9878 nor n9937 n9941 ; n9942
g9879 nor n9940 n9941 ; n9943
g9880 nor n9942 n9943 ; n9944
g9881 and n587_not n7983 ; n9945
g9882 and n867_not n7291 ; n9946
g9883 and n710_not n7632 ; n9947
g9884 nor n9946 n9947 ; n9948
g9885 and n9945_not n9948 ; n9949
g9886 and n3331 n7294 ; n9950
g9887 and n9949 n9950_not ; n9951
g9888 and a[11] n9951_not ; n9952
g9889 nor n9951 n9952 ; n9953
g9890 and a[11] n9952_not ; n9954
g9891 nor n9953 n9954 ; n9955
g9892 nor n9808 n9812 ; n9956
g9893 nor n9811 n9812 ; n9957
g9894 nor n9956 n9957 ; n9958
g9895 nor n9955 n9958 ; n9959
g9896 nor n9955 n9959 ; n9960
g9897 nor n9958 n9959 ; n9961
g9898 nor n9960 n9961 ; n9962
g9899 and n710_not n7983 ; n9963
g9900 and n958_not n7291 ; n9964
g9901 and n867_not n7632 ; n9965
g9902 nor n9964 n9965 ; n9966
g9903 and n9963_not n9966 ; n9967
g9904 and n4179 n7294 ; n9968
g9905 and n9967 n9968_not ; n9969
g9906 and a[11] n9969_not ; n9970
g9907 nor n9969 n9970 ; n9971
g9908 and a[11] n9970_not ; n9972
g9909 nor n9971 n9972 ; n9973
g9910 nor n9803 n9807 ; n9974
g9911 nor n9806 n9807 ; n9975
g9912 nor n9974 n9975 ; n9976
g9913 nor n9973 n9976 ; n9977
g9914 nor n9973 n9977 ; n9978
g9915 nor n9976 n9977 ; n9979
g9916 nor n9978 n9979 ; n9980
g9917 and n867_not n7983 ; n9981
g9918 and n1060_not n7291 ; n9982
g9919 and n958_not n7632 ; n9983
g9920 nor n9982 n9983 ; n9984
g9921 and n9981_not n9984 ; n9985
g9922 and n4204 n7294 ; n9986
g9923 and n9985 n9986_not ; n9987
g9924 and a[11] n9987_not ; n9988
g9925 nor n9987 n9988 ; n9989
g9926 and a[11] n9988_not ; n9990
g9927 nor n9989 n9990 ; n9991
g9928 nor n9798 n9802 ; n9992
g9929 nor n9801 n9802 ; n9993
g9930 nor n9992 n9993 ; n9994
g9931 nor n9991 n9994 ; n9995
g9932 nor n9991 n9995 ; n9996
g9933 nor n9994 n9995 ; n9997
g9934 nor n9996 n9997 ; n9998
g9935 and n958_not n7983 ; n9999
g9936 and n1178_not n7291 ; n10000
g9937 and n1060_not n7632 ; n10001
g9938 nor n10000 n10001 ; n10002
g9939 and n9999_not n10002 ; n10003
g9940 and n4633 n7294 ; n10004
g9941 and n10003 n10004_not ; n10005
g9942 and a[11] n10005_not ; n10006
g9943 nor n10005 n10006 ; n10007
g9944 and a[11] n10006_not ; n10008
g9945 nor n10007 n10008 ; n10009
g9946 nor n9793 n9797 ; n10010
g9947 nor n9796 n9797 ; n10011
g9948 nor n10010 n10011 ; n10012
g9949 nor n10009 n10012 ; n10013
g9950 nor n10009 n10013 ; n10014
g9951 nor n10012 n10013 ; n10015
g9952 nor n10014 n10015 ; n10016
g9953 and n9484 n9791 ; n10017
g9954 nor n9792 n10017 ; n10018
g9955 and n1060_not n7983 ; n10019
g9956 and n1235_not n7291 ; n10020
g9957 and n1178_not n7632 ; n10021
g9958 nor n10020 n10021 ; n10022
g9959 and n10019_not n10022 ; n10023
g9960 and n7294_not n10023 ; n10024
g9961 and n4429_not n10023 ; n10025
g9962 nor n10024 n10025 ; n10026
g9963 and a[11] n10026_not ; n10027
g9964 and a[11]_not n10026 ; n10028
g9965 nor n10027 n10028 ; n10029
g9966 and n10018 n10029_not ; n10030
g9967 and n9502 n9789 ; n10031
g9968 nor n9790 n10031 ; n10032
g9969 and n1178_not n7983 ; n10033
g9970 and n1364_not n7291 ; n10034
g9971 and n1235_not n7632 ; n10035
g9972 nor n10034 n10035 ; n10036
g9973 and n10033_not n10036 ; n10037
g9974 and n7294_not n10037 ; n10038
g9975 and n4861_not n10037 ; n10039
g9976 nor n10038 n10039 ; n10040
g9977 and a[11] n10040_not ; n10041
g9978 and a[11]_not n10040 ; n10042
g9979 nor n10041 n10042 ; n10043
g9980 and n10032 n10043_not ; n10044
g9981 and n1235_not n7983 ; n10045
g9982 and n1472_not n7291 ; n10046
g9983 and n1364_not n7632 ; n10047
g9984 nor n10046 n10047 ; n10048
g9985 and n10045_not n10048 ; n10049
g9986 and n4848 n7294 ; n10050
g9987 and n10049 n10050_not ; n10051
g9988 and a[11] n10051_not ; n10052
g9989 nor n10051 n10052 ; n10053
g9990 and a[11] n10052_not ; n10054
g9991 nor n10053 n10054 ; n10055
g9992 and n9785 n9787_not ; n10056
g9993 nor n9788 n10056 ; n10057
g9994 and n10055_not n10057 ; n10058
g9995 nor n10055 n10058 ; n10059
g9996 and n10057 n10058_not ; n10060
g9997 nor n10059 n10060 ; n10061
g9998 and n1364_not n7983 ; n10062
g9999 and n1572_not n7291 ; n10063
g10000 and n1472_not n7632 ; n10064
g10001 nor n10063 n10064 ; n10065
g10002 and n10062_not n10065 ; n10066
g10003 and n5114 n7294 ; n10067
g10004 and n10066 n10067_not ; n10068
g10005 and a[11] n10068_not ; n10069
g10006 nor n10068 n10069 ; n10070
g10007 and a[11] n10069_not ; n10071
g10008 nor n10070 n10071 ; n10072
g10009 nor n9780 n9784 ; n10073
g10010 nor n9783 n9784 ; n10074
g10011 nor n10073 n10074 ; n10075
g10012 nor n10072 n10075 ; n10076
g10013 nor n10072 n10076 ; n10077
g10014 nor n10075 n10076 ; n10078
g10015 nor n10077 n10078 ; n10079
g10016 and n1472_not n7983 ; n10080
g10017 and n1665_not n7291 ; n10081
g10018 and n1572_not n7632 ; n10082
g10019 nor n10081 n10082 ; n10083
g10020 and n10080_not n10083 ; n10084
g10021 and n5139 n7294 ; n10085
g10022 and n10084 n10085_not ; n10086
g10023 and a[11] n10086_not ; n10087
g10024 nor n10086 n10087 ; n10088
g10025 and a[11] n10087_not ; n10089
g10026 nor n10088 n10089 ; n10090
g10027 nor n9775 n9779 ; n10091
g10028 nor n9778 n9779 ; n10092
g10029 nor n10091 n10092 ; n10093
g10030 nor n10090 n10093 ; n10094
g10031 nor n10090 n10094 ; n10095
g10032 nor n10093 n10094 ; n10096
g10033 nor n10095 n10096 ; n10097
g10034 and n9561 n9773 ; n10098
g10035 nor n9774 n10098 ; n10099
g10036 and n1572_not n7983 ; n10100
g10037 and n1779_not n7291 ; n10101
g10038 and n1665_not n7632 ; n10102
g10039 nor n10101 n10102 ; n10103
g10040 and n10100_not n10103 ; n10104
g10041 and n7294_not n10104 ; n10105
g10042 and n5561_not n10104 ; n10106
g10043 nor n10105 n10106 ; n10107
g10044 and a[11] n10107_not ; n10108
g10045 and a[11]_not n10107 ; n10109
g10046 nor n10108 n10109 ; n10110
g10047 and n10099 n10110_not ; n10111
g10048 and n9579 n9771 ; n10112
g10049 nor n9772 n10112 ; n10113
g10050 and n1665_not n7983 ; n10114
g10051 and n1877_not n7291 ; n10115
g10052 and n1779_not n7632 ; n10116
g10053 nor n10115 n10116 ; n10117
g10054 and n10114_not n10117 ; n10118
g10055 and n7294_not n10118 ; n10119
g10056 and n5328_not n10118 ; n10120
g10057 nor n10119 n10120 ; n10121
g10058 and a[11] n10121_not ; n10122
g10059 and a[11]_not n10121 ; n10123
g10060 nor n10122 n10123 ; n10124
g10061 and n10113 n10124_not ; n10125
g10062 and n9597 n9769 ; n10126
g10063 nor n9770 n10126 ; n10127
g10064 and n1779_not n7983 ; n10128
g10065 and n1913_not n7291 ; n10129
g10066 and n1877_not n7632 ; n10130
g10067 nor n10129 n10130 ; n10131
g10068 and n10128_not n10131 ; n10132
g10069 and n7294_not n10132 ; n10133
g10070 and n5851_not n10132 ; n10134
g10071 nor n10133 n10134 ; n10135
g10072 and a[11] n10135_not ; n10136
g10073 and a[11]_not n10135 ; n10137
g10074 nor n10136 n10137 ; n10138
g10075 and n10127 n10138_not ; n10139
g10076 and n1877_not n7983 ; n10140
g10077 and n1992_not n7291 ; n10141
g10078 and n1913_not n7632 ; n10142
g10079 nor n10141 n10142 ; n10143
g10080 and n10140_not n10143 ; n10144
g10081 and n6007 n7294 ; n10145
g10082 and n10144 n10145_not ; n10146
g10083 and a[11] n10146_not ; n10147
g10084 nor n10146 n10147 ; n10148
g10085 and a[11] n10147_not ; n10149
g10086 nor n10148 n10149 ; n10150
g10087 and n9765 n9767_not ; n10151
g10088 nor n9768 n10151 ; n10152
g10089 and n10150_not n10152 ; n10153
g10090 nor n10150 n10153 ; n10154
g10091 and n10152 n10153_not ; n10155
g10092 nor n10154 n10155 ; n10156
g10093 and n1913_not n7983 ; n10157
g10094 and n2057_not n7291 ; n10158
g10095 and n1992_not n7632 ; n10159
g10096 nor n10158 n10159 ; n10160
g10097 and n10157_not n10160 ; n10161
g10098 and n5834 n7294 ; n10162
g10099 and n10161 n10162_not ; n10163
g10100 and a[11] n10163_not ; n10164
g10101 nor n10163 n10164 ; n10165
g10102 and a[11] n10164_not ; n10166
g10103 nor n10165 n10166 ; n10167
g10104 nor n9760 n9764 ; n10168
g10105 nor n9763 n9764 ; n10169
g10106 nor n10168 n10169 ; n10170
g10107 nor n10167 n10170 ; n10171
g10108 nor n10167 n10171 ; n10172
g10109 nor n10170 n10171 ; n10173
g10110 nor n10172 n10173 ; n10174
g10111 and n1992_not n7983 ; n10175
g10112 and n2152_not n7291 ; n10176
g10113 and n2057_not n7632 ; n10177
g10114 nor n10176 n10177 ; n10178
g10115 and n10175_not n10178 ; n10179
g10116 and n6143 n7294 ; n10180
g10117 and n10179 n10180_not ; n10181
g10118 and a[11] n10181_not ; n10182
g10119 nor n10181 n10182 ; n10183
g10120 and a[11] n10182_not ; n10184
g10121 nor n10183 n10184 ; n10185
g10122 nor n9755 n9759 ; n10186
g10123 nor n9758 n9759 ; n10187
g10124 nor n10186 n10187 ; n10188
g10125 nor n10185 n10188 ; n10189
g10126 nor n10185 n10189 ; n10190
g10127 nor n10188 n10189 ; n10191
g10128 nor n10190 n10191 ; n10192
g10129 and n9656 n9753 ; n10193
g10130 nor n9754 n10193 ; n10194
g10131 and n2057_not n7983 ; n10195
g10132 and n2189_not n7291 ; n10196
g10133 and n2152_not n7632 ; n10197
g10134 nor n10196 n10197 ; n10198
g10135 and n10195_not n10198 ; n10199
g10136 and n7294_not n10199 ; n10200
g10137 and n6479_not n10199 ; n10201
g10138 nor n10200 n10201 ; n10202
g10139 and a[11] n10202_not ; n10203
g10140 and a[11]_not n10202 ; n10204
g10141 nor n10203 n10204 ; n10205
g10142 and n10194 n10205_not ; n10206
g10143 and n9749 n9751_not ; n10207
g10144 nor n9752 n10207 ; n10208
g10145 and n2152_not n7983 ; n10209
g10146 and n2291_not n7291 ; n10210
g10147 and n2189_not n7632 ; n10211
g10148 nor n10210 n10211 ; n10212
g10149 and n10209_not n10212 ; n10213
g10150 and n7294_not n10213 ; n10214
g10151 and n6492_not n10213 ; n10215
g10152 nor n10214 n10215 ; n10216
g10153 and a[11] n10216_not ; n10217
g10154 and a[11]_not n10216 ; n10218
g10155 nor n10217 n10218 ; n10219
g10156 and n10208 n10219_not ; n10220
g10157 and n9688 n9747 ; n10221
g10158 nor n9748 n10221 ; n10222
g10159 and n2189_not n7983 ; n10223
g10160 and n2388_not n7291 ; n10224
g10161 and n2291_not n7632 ; n10225
g10162 nor n10224 n10225 ; n10226
g10163 and n10223_not n10226 ; n10227
g10164 and n7294_not n10227 ; n10228
g10165 and n6122_not n10227 ; n10229
g10166 nor n10228 n10229 ; n10230
g10167 and a[11] n10230_not ; n10231
g10168 and a[11]_not n10230 ; n10232
g10169 nor n10231 n10232 ; n10233
g10170 and n10222 n10233_not ; n10234
g10171 and n2291_not n7983 ; n10235
g10172 and n2464_not n7291 ; n10236
g10173 and n2388_not n7632 ; n10237
g10174 nor n10236 n10237 ; n10238
g10175 and n10235_not n10238 ; n10239
g10176 and n6541 n7294 ; n10240
g10177 and n10239 n10240_not ; n10241
g10178 and a[11] n10241_not ; n10242
g10179 nor n10241 n10242 ; n10243
g10180 and a[11] n10242_not ; n10244
g10181 nor n10243 n10244 ; n10245
g10182 and n9743 n9745_not ; n10246
g10183 nor n9746 n10246 ; n10247
g10184 and n10245_not n10247 ; n10248
g10185 nor n10245 n10248 ; n10249
g10186 and n10247 n10248_not ; n10250
g10187 nor n10249 n10250 ; n10251
g10188 nor n9730 n9742 ; n10252
g10189 nor n9741 n9742 ; n10253
g10190 nor n10252 n10253 ; n10254
g10191 and n2388_not n7983 ; n10255
g10192 and n2533_not n7291 ; n10256
g10193 and n2464_not n7632 ; n10257
g10194 nor n10256 n10257 ; n10258
g10195 and n10255_not n10258 ; n10259
g10196 and n7294_not n10259 ; n10260
g10197 and n6591_not n10259 ; n10261
g10198 nor n10260 n10261 ; n10262
g10199 and a[11] n10262_not ; n10263
g10200 and a[11]_not n10262 ; n10264
g10201 nor n10263 n10264 ; n10265
g10202 nor n10254 n10265 ; n10266
g10203 and n2464_not n7983 ; n10267
g10204 and n2571_not n7291 ; n10268
g10205 and n2533_not n7632 ; n10269
g10206 nor n10268 n10269 ; n10270
g10207 and n10267_not n10270 ; n10271
g10208 and n6646 n7294 ; n10272
g10209 and n10271 n10272_not ; n10273
g10210 and a[11] n10273_not ; n10274
g10211 nor n10273 n10274 ; n10275
g10212 and a[11] n10274_not ; n10276
g10213 nor n10275 n10276 ; n10277
g10214 and n9714_not n9725 ; n10278
g10215 nor n9726 n10278 ; n10279
g10216 and n10277_not n10279 ; n10280
g10217 nor n10277 n10280 ; n10281
g10218 and n10279 n10280_not ; n10282
g10219 nor n10281 n10282 ; n10283
g10220 and n9711 n9713_not ; n10284
g10221 nor n9714 n10284 ; n10285
g10222 and n2533_not n7983 ; n10286
g10223 and n2674_not n7291 ; n10287
g10224 and n2571_not n7632 ; n10288
g10225 nor n10287 n10288 ; n10289
g10226 and n10286_not n10289 ; n10290
g10227 and n7294_not n10290 ; n10291
g10228 and n6695_not n10290 ; n10292
g10229 nor n10291 n10292 ; n10293
g10230 and a[11] n10293_not ; n10294
g10231 and a[11]_not n10293 ; n10295
g10232 nor n10294 n10295 ; n10296
g10233 and n10285 n10296_not ; n10297
g10234 and n2829_not n7632 ; n10298
g10235 and n2736_not n7983 ; n10299
g10236 nor n10298 n10299 ; n10300
g10237 and n7294 n7469_not ; n10301
g10238 and n10300 n10301_not ; n10302
g10239 and a[11] n10302_not ; n10303
g10240 and a[11] n10303_not ; n10304
g10241 nor n10302 n10303 ; n10305
g10242 nor n10304 n10305 ; n10306
g10243 nor n2829 n7289 ; n10307
g10244 and a[11] n10307_not ; n10308
g10245 and n10306_not n10308 ; n10309
g10246 and n2674_not n7983 ; n10310
g10247 and n2829_not n7291 ; n10311
g10248 and n2736_not n7632 ; n10312
g10249 nor n10311 n10312 ; n10313
g10250 and n10310_not n10313 ; n10314
g10251 and n7294_not n10314 ; n10315
g10252 and n6798_not n10314 ; n10316
g10253 nor n10315 n10316 ; n10317
g10254 and a[11] n10317_not ; n10318
g10255 and a[11]_not n10317 ; n10319
g10256 nor n10318 n10319 ; n10320
g10257 and n10309 n10320_not ; n10321
g10258 and n9712 n10321 ; n10322
g10259 and n10321 n10322_not ; n10323
g10260 and n9712 n10322_not ; n10324
g10261 nor n10323 n10324 ; n10325
g10262 and n2571_not n7983 ; n10326
g10263 and n2736_not n7291 ; n10327
g10264 and n2674_not n7632 ; n10328
g10265 nor n10327 n10328 ; n10329
g10266 and n10326_not n10329 ; n10330
g10267 and n6806 n7294 ; n10331
g10268 and n10330 n10331_not ; n10332
g10269 and a[11] n10332_not ; n10333
g10270 and a[11] n10333_not ; n10334
g10271 nor n10332 n10333 ; n10335
g10272 nor n10334 n10335 ; n10336
g10273 nor n10325 n10336 ; n10337
g10274 nor n10322 n10337 ; n10338
g10275 and n10285_not n10296 ; n10339
g10276 nor n10297 n10339 ; n10340
g10277 and n10338_not n10340 ; n10341
g10278 nor n10297 n10341 ; n10342
g10279 nor n10283 n10342 ; n10343
g10280 nor n10280 n10343 ; n10344
g10281 and n10254 n10265 ; n10345
g10282 nor n10266 n10345 ; n10346
g10283 and n10344_not n10346 ; n10347
g10284 nor n10266 n10347 ; n10348
g10285 nor n10251 n10348 ; n10349
g10286 nor n10248 n10349 ; n10350
g10287 and n10222 n10234_not ; n10351
g10288 nor n10233 n10234 ; n10352
g10289 nor n10351 n10352 ; n10353
g10290 nor n10350 n10353 ; n10354
g10291 nor n10234 n10354 ; n10355
g10292 and n10208 n10220_not ; n10356
g10293 nor n10219 n10220 ; n10357
g10294 nor n10356 n10357 ; n10358
g10295 nor n10355 n10358 ; n10359
g10296 nor n10220 n10359 ; n10360
g10297 and n10194_not n10205 ; n10361
g10298 nor n10206 n10361 ; n10362
g10299 and n10360_not n10362 ; n10363
g10300 nor n10206 n10363 ; n10364
g10301 nor n10192 n10364 ; n10365
g10302 nor n10189 n10365 ; n10366
g10303 nor n10174 n10366 ; n10367
g10304 nor n10171 n10367 ; n10368
g10305 nor n10156 n10368 ; n10369
g10306 nor n10153 n10369 ; n10370
g10307 and n10127 n10139_not ; n10371
g10308 nor n10138 n10139 ; n10372
g10309 nor n10371 n10372 ; n10373
g10310 nor n10370 n10373 ; n10374
g10311 nor n10139 n10374 ; n10375
g10312 and n10113 n10125_not ; n10376
g10313 nor n10124 n10125 ; n10377
g10314 nor n10376 n10377 ; n10378
g10315 nor n10375 n10378 ; n10379
g10316 nor n10125 n10379 ; n10380
g10317 and n10099_not n10110 ; n10381
g10318 nor n10111 n10381 ; n10382
g10319 and n10380_not n10382 ; n10383
g10320 nor n10111 n10383 ; n10384
g10321 nor n10097 n10384 ; n10385
g10322 nor n10094 n10385 ; n10386
g10323 nor n10079 n10386 ; n10387
g10324 nor n10076 n10387 ; n10388
g10325 nor n10061 n10388 ; n10389
g10326 nor n10058 n10389 ; n10390
g10327 and n10032 n10044_not ; n10391
g10328 nor n10043 n10044 ; n10392
g10329 nor n10391 n10392 ; n10393
g10330 nor n10390 n10393 ; n10394
g10331 nor n10044 n10394 ; n10395
g10332 and n10018_not n10029 ; n10396
g10333 nor n10030 n10396 ; n10397
g10334 and n10395_not n10397 ; n10398
g10335 nor n10030 n10398 ; n10399
g10336 nor n10016 n10399 ; n10400
g10337 nor n10013 n10400 ; n10401
g10338 nor n9998 n10401 ; n10402
g10339 nor n9995 n10402 ; n10403
g10340 nor n9980 n10403 ; n10404
g10341 nor n9977 n10404 ; n10405
g10342 nor n9962 n10405 ; n10406
g10343 nor n9959 n10406 ; n10407
g10344 nor n9944 n10407 ; n10408
g10345 nor n9941 n10408 ; n10409
g10346 nor n9926 n10409 ; n10410
g10347 nor n9923 n10410 ; n10411
g10348 nor n9908 n10411 ; n10412
g10349 nor n9905 n10412 ; n10413
g10350 and n9842 n9844_not ; n10414
g10351 nor n9845 n10414 ; n10415
g10352 and n10413_not n10415 ; n10416
g10353 and n3964_not n9331 ; n10417
g10354 and n3456_not n8418 ; n10418
g10355 and n3805_not n8860 ; n10419
g10356 nor n10418 n10419 ; n10420
g10357 and n10417_not n10420 ; n10421
g10358 and n4558 n8421 ; n10422
g10359 and n10421 n10422_not ; n10423
g10360 and a[8] n10423_not ; n10424
g10361 nor n10423 n10424 ; n10425
g10362 and a[8] n10424_not ; n10426
g10363 nor n10425 n10426 ; n10427
g10364 nor n10413 n10416 ; n10428
g10365 and n10415 n10416_not ; n10429
g10366 nor n10428 n10429 ; n10430
g10367 nor n10427 n10430 ; n10431
g10368 nor n10416 n10431 ; n10432
g10369 and n3877_not n9867 ; n10433
g10370 and n70 n9865_not ; n10434
g10371 and n4515_not n10434 ; n10435
g10372 nor n10433 n10435 ; n10436
g10373 and n9870_not n10436 ; n10437
g10374 and n4609_not n10436 ; n10438
g10375 nor n10437 n10438 ; n10439
g10376 and a[5] n10439_not ; n10440
g10377 and a[5]_not n10439 ; n10441
g10378 nor n10440 n10441 ; n10442
g10379 nor n10432 n10442 ; n10443
g10380 and n9849 n9861_not ; n10444
g10381 nor n9860 n9861 ; n10445
g10382 nor n10444 n10445 ; n10446
g10383 and n10432 n10442 ; n10447
g10384 nor n10443 n10447 ; n10448
g10385 and n10446_not n10448 ; n10449
g10386 nor n10443 n10449 ; n10450
g10387 nor n9890 n10450 ; n10451
g10388 and n9890 n10450 ; n10452
g10389 nor n10451 n10452 ; n10453
g10390 and n9908 n10411 ; n10454
g10391 nor n10412 n10454 ; n10455
g10392 and n3805_not n9331 ; n10456
g10393 and n3605_not n8418 ; n10457
g10394 and n3456_not n8860 ; n10458
g10395 nor n10457 n10458 ; n10459
g10396 and n10456_not n10459 ; n10460
g10397 and n8421_not n10460 ; n10461
g10398 and n3818_not n10460 ; n10462
g10399 nor n10461 n10462 ; n10463
g10400 and a[8] n10463_not ; n10464
g10401 and a[8]_not n10463 ; n10465
g10402 nor n10464 n10465 ; n10466
g10403 and n10455 n10466_not ; n10467
g10404 and n9926 n10409 ; n10468
g10405 nor n10410 n10468 ; n10469
g10406 and n3456_not n9331 ; n10470
g10407 and n3539_not n8418 ; n10471
g10408 and n3605_not n8860 ; n10472
g10409 nor n10471 n10472 ; n10473
g10410 and n10470_not n10473 ; n10474
g10411 and n8421_not n10474 ; n10475
g10412 and n3627_not n10474 ; n10476
g10413 nor n10475 n10476 ; n10477
g10414 and a[8] n10477_not ; n10478
g10415 and a[8]_not n10477 ; n10479
g10416 nor n10478 n10479 ; n10480
g10417 and n10469 n10480_not ; n10481
g10418 and n9944 n10407 ; n10482
g10419 nor n10408 n10482 ; n10483
g10420 and n3605_not n9331 ; n10484
g10421 and n3012_not n8418 ; n10485
g10422 and n3539_not n8860 ; n10486
g10423 nor n10485 n10486 ; n10487
g10424 and n10484_not n10487 ; n10488
g10425 and n8421_not n10488 ; n10489
g10426 and n4084_not n10488 ; n10490
g10427 nor n10489 n10490 ; n10491
g10428 and a[8] n10491_not ; n10492
g10429 and a[8]_not n10491 ; n10493
g10430 nor n10492 n10493 ; n10494
g10431 and n10483 n10494_not ; n10495
g10432 and n9962 n10405 ; n10496
g10433 nor n10406 n10496 ; n10497
g10434 and n3539_not n9331 ; n10498
g10435 and n392_not n8418 ; n10499
g10436 and n3012_not n8860 ; n10500
g10437 nor n10499 n10500 ; n10501
g10438 and n10498_not n10501 ; n10502
g10439 and n8421_not n10502 ; n10503
g10440 and n3715_not n10502 ; n10504
g10441 nor n10503 n10504 ; n10505
g10442 and a[8] n10505_not ; n10506
g10443 and a[8]_not n10505 ; n10507
g10444 nor n10506 n10507 ; n10508
g10445 and n10497 n10508_not ; n10509
g10446 and n9980 n10403 ; n10510
g10447 nor n10404 n10510 ; n10511
g10448 and n3012_not n9331 ; n10512
g10449 and n587_not n8418 ; n10513
g10450 and n392_not n8860 ; n10514
g10451 nor n10513 n10514 ; n10515
g10452 and n10512_not n10515 ; n10516
g10453 and n8421_not n10516 ; n10517
g10454 and n3018_not n10516 ; n10518
g10455 nor n10517 n10518 ; n10519
g10456 and a[8] n10519_not ; n10520
g10457 and a[8]_not n10519 ; n10521
g10458 nor n10520 n10521 ; n10522
g10459 and n10511 n10522_not ; n10523
g10460 and n9998 n10401 ; n10524
g10461 nor n10402 n10524 ; n10525
g10462 and n392_not n9331 ; n10526
g10463 and n710_not n8418 ; n10527
g10464 and n587_not n8860 ; n10528
g10465 nor n10527 n10528 ; n10529
g10466 and n10526_not n10529 ; n10530
g10467 and n8421_not n10530 ; n10531
g10468 and n3347_not n10530 ; n10532
g10469 nor n10531 n10532 ; n10533
g10470 and a[8] n10533_not ; n10534
g10471 and a[8]_not n10533 ; n10535
g10472 nor n10534 n10535 ; n10536
g10473 and n10525 n10536_not ; n10537
g10474 and n10016 n10399 ; n10538
g10475 nor n10400 n10538 ; n10539
g10476 and n587_not n9331 ; n10540
g10477 and n867_not n8418 ; n10541
g10478 and n710_not n8860 ; n10542
g10479 nor n10541 n10542 ; n10543
g10480 and n10540_not n10543 ; n10544
g10481 and n8421_not n10544 ; n10545
g10482 and n3331_not n10544 ; n10546
g10483 nor n10545 n10546 ; n10547
g10484 and a[8] n10547_not ; n10548
g10485 and a[8]_not n10547 ; n10549
g10486 nor n10548 n10549 ; n10550
g10487 and n10539 n10550_not ; n10551
g10488 and n710_not n9331 ; n10552
g10489 and n958_not n8418 ; n10553
g10490 and n867_not n8860 ; n10554
g10491 nor n10553 n10554 ; n10555
g10492 and n10552_not n10555 ; n10556
g10493 and n4179 n8421 ; n10557
g10494 and n10556 n10557_not ; n10558
g10495 and a[8] n10558_not ; n10559
g10496 nor n10558 n10559 ; n10560
g10497 and a[8] n10559_not ; n10561
g10498 nor n10560 n10561 ; n10562
g10499 and n10395 n10397_not ; n10563
g10500 nor n10398 n10563 ; n10564
g10501 and n10562_not n10564 ; n10565
g10502 nor n10562 n10565 ; n10566
g10503 and n10564 n10565_not ; n10567
g10504 nor n10566 n10567 ; n10568
g10505 and n867_not n9331 ; n10569
g10506 and n1060_not n8418 ; n10570
g10507 and n958_not n8860 ; n10571
g10508 nor n10570 n10571 ; n10572
g10509 and n10569_not n10572 ; n10573
g10510 and n4204 n8421 ; n10574
g10511 and n10573 n10574_not ; n10575
g10512 and a[8] n10575_not ; n10576
g10513 nor n10575 n10576 ; n10577
g10514 and a[8] n10576_not ; n10578
g10515 nor n10577 n10578 ; n10579
g10516 nor n10390 n10394 ; n10580
g10517 nor n10393 n10394 ; n10581
g10518 nor n10580 n10581 ; n10582
g10519 nor n10579 n10582 ; n10583
g10520 nor n10579 n10583 ; n10584
g10521 nor n10582 n10583 ; n10585
g10522 nor n10584 n10585 ; n10586
g10523 and n10061 n10388 ; n10587
g10524 nor n10389 n10587 ; n10588
g10525 and n958_not n9331 ; n10589
g10526 and n1178_not n8418 ; n10590
g10527 and n1060_not n8860 ; n10591
g10528 nor n10590 n10591 ; n10592
g10529 and n10589_not n10592 ; n10593
g10530 and n8421_not n10593 ; n10594
g10531 and n4633_not n10593 ; n10595
g10532 nor n10594 n10595 ; n10596
g10533 and a[8] n10596_not ; n10597
g10534 and a[8]_not n10596 ; n10598
g10535 nor n10597 n10598 ; n10599
g10536 and n10588 n10599_not ; n10600
g10537 and n10079 n10386 ; n10601
g10538 nor n10387 n10601 ; n10602
g10539 and n1060_not n9331 ; n10603
g10540 and n1235_not n8418 ; n10604
g10541 and n1178_not n8860 ; n10605
g10542 nor n10604 n10605 ; n10606
g10543 and n10603_not n10606 ; n10607
g10544 and n8421_not n10607 ; n10608
g10545 and n4429_not n10607 ; n10609
g10546 nor n10608 n10609 ; n10610
g10547 and a[8] n10610_not ; n10611
g10548 and a[8]_not n10610 ; n10612
g10549 nor n10611 n10612 ; n10613
g10550 and n10602 n10613_not ; n10614
g10551 and n10097 n10384 ; n10615
g10552 nor n10385 n10615 ; n10616
g10553 and n1178_not n9331 ; n10617
g10554 and n1364_not n8418 ; n10618
g10555 and n1235_not n8860 ; n10619
g10556 nor n10618 n10619 ; n10620
g10557 and n10617_not n10620 ; n10621
g10558 and n8421_not n10621 ; n10622
g10559 and n4861_not n10621 ; n10623
g10560 nor n10622 n10623 ; n10624
g10561 and a[8] n10624_not ; n10625
g10562 and a[8]_not n10624 ; n10626
g10563 nor n10625 n10626 ; n10627
g10564 and n10616 n10627_not ; n10628
g10565 and n1235_not n9331 ; n10629
g10566 and n1472_not n8418 ; n10630
g10567 and n1364_not n8860 ; n10631
g10568 nor n10630 n10631 ; n10632
g10569 and n10629_not n10632 ; n10633
g10570 and n4848 n8421 ; n10634
g10571 and n10633 n10634_not ; n10635
g10572 and a[8] n10635_not ; n10636
g10573 nor n10635 n10636 ; n10637
g10574 and a[8] n10636_not ; n10638
g10575 nor n10637 n10638 ; n10639
g10576 and n10380 n10382_not ; n10640
g10577 nor n10383 n10640 ; n10641
g10578 and n10639_not n10641 ; n10642
g10579 nor n10639 n10642 ; n10643
g10580 and n10641 n10642_not ; n10644
g10581 nor n10643 n10644 ; n10645
g10582 and n1364_not n9331 ; n10646
g10583 and n1572_not n8418 ; n10647
g10584 and n1472_not n8860 ; n10648
g10585 nor n10647 n10648 ; n10649
g10586 and n10646_not n10649 ; n10650
g10587 and n5114 n8421 ; n10651
g10588 and n10650 n10651_not ; n10652
g10589 and a[8] n10652_not ; n10653
g10590 nor n10652 n10653 ; n10654
g10591 and a[8] n10653_not ; n10655
g10592 nor n10654 n10655 ; n10656
g10593 nor n10375 n10379 ; n10657
g10594 nor n10378 n10379 ; n10658
g10595 nor n10657 n10658 ; n10659
g10596 nor n10656 n10659 ; n10660
g10597 nor n10656 n10660 ; n10661
g10598 nor n10659 n10660 ; n10662
g10599 nor n10661 n10662 ; n10663
g10600 and n1472_not n9331 ; n10664
g10601 and n1665_not n8418 ; n10665
g10602 and n1572_not n8860 ; n10666
g10603 nor n10665 n10666 ; n10667
g10604 and n10664_not n10667 ; n10668
g10605 and n5139 n8421 ; n10669
g10606 and n10668 n10669_not ; n10670
g10607 and a[8] n10670_not ; n10671
g10608 nor n10670 n10671 ; n10672
g10609 and a[8] n10671_not ; n10673
g10610 nor n10672 n10673 ; n10674
g10611 nor n10370 n10374 ; n10675
g10612 nor n10373 n10374 ; n10676
g10613 nor n10675 n10676 ; n10677
g10614 nor n10674 n10677 ; n10678
g10615 nor n10674 n10678 ; n10679
g10616 nor n10677 n10678 ; n10680
g10617 nor n10679 n10680 ; n10681
g10618 and n10156 n10368 ; n10682
g10619 nor n10369 n10682 ; n10683
g10620 and n1572_not n9331 ; n10684
g10621 and n1779_not n8418 ; n10685
g10622 and n1665_not n8860 ; n10686
g10623 nor n10685 n10686 ; n10687
g10624 and n10684_not n10687 ; n10688
g10625 and n8421_not n10688 ; n10689
g10626 and n5561_not n10688 ; n10690
g10627 nor n10689 n10690 ; n10691
g10628 and a[8] n10691_not ; n10692
g10629 and a[8]_not n10691 ; n10693
g10630 nor n10692 n10693 ; n10694
g10631 and n10683 n10694_not ; n10695
g10632 and n10174 n10366 ; n10696
g10633 nor n10367 n10696 ; n10697
g10634 and n1665_not n9331 ; n10698
g10635 and n1877_not n8418 ; n10699
g10636 and n1779_not n8860 ; n10700
g10637 nor n10699 n10700 ; n10701
g10638 and n10698_not n10701 ; n10702
g10639 and n8421_not n10702 ; n10703
g10640 and n5328_not n10702 ; n10704
g10641 nor n10703 n10704 ; n10705
g10642 and a[8] n10705_not ; n10706
g10643 and a[8]_not n10705 ; n10707
g10644 nor n10706 n10707 ; n10708
g10645 and n10697 n10708_not ; n10709
g10646 and n10192 n10364 ; n10710
g10647 nor n10365 n10710 ; n10711
g10648 and n1779_not n9331 ; n10712
g10649 and n1913_not n8418 ; n10713
g10650 and n1877_not n8860 ; n10714
g10651 nor n10713 n10714 ; n10715
g10652 and n10712_not n10715 ; n10716
g10653 and n8421_not n10716 ; n10717
g10654 and n5851_not n10716 ; n10718
g10655 nor n10717 n10718 ; n10719
g10656 and a[8] n10719_not ; n10720
g10657 and a[8]_not n10719 ; n10721
g10658 nor n10720 n10721 ; n10722
g10659 and n10711 n10722_not ; n10723
g10660 and n1877_not n9331 ; n10724
g10661 and n1992_not n8418 ; n10725
g10662 and n1913_not n8860 ; n10726
g10663 nor n10725 n10726 ; n10727
g10664 and n10724_not n10727 ; n10728
g10665 and n6007 n8421 ; n10729
g10666 and n10728 n10729_not ; n10730
g10667 and a[8] n10730_not ; n10731
g10668 nor n10730 n10731 ; n10732
g10669 and a[8] n10731_not ; n10733
g10670 nor n10732 n10733 ; n10734
g10671 and n10360 n10362_not ; n10735
g10672 nor n10363 n10735 ; n10736
g10673 and n10734_not n10736 ; n10737
g10674 nor n10734 n10737 ; n10738
g10675 and n10736 n10737_not ; n10739
g10676 nor n10738 n10739 ; n10740
g10677 and n1913_not n9331 ; n10741
g10678 and n2057_not n8418 ; n10742
g10679 and n1992_not n8860 ; n10743
g10680 nor n10742 n10743 ; n10744
g10681 and n10741_not n10744 ; n10745
g10682 and n5834 n8421 ; n10746
g10683 and n10745 n10746_not ; n10747
g10684 and a[8] n10747_not ; n10748
g10685 nor n10747 n10748 ; n10749
g10686 and a[8] n10748_not ; n10750
g10687 nor n10749 n10750 ; n10751
g10688 nor n10355 n10359 ; n10752
g10689 nor n10358 n10359 ; n10753
g10690 nor n10752 n10753 ; n10754
g10691 nor n10751 n10754 ; n10755
g10692 nor n10751 n10755 ; n10756
g10693 nor n10754 n10755 ; n10757
g10694 nor n10756 n10757 ; n10758
g10695 and n1992_not n9331 ; n10759
g10696 and n2152_not n8418 ; n10760
g10697 and n2057_not n8860 ; n10761
g10698 nor n10760 n10761 ; n10762
g10699 and n10759_not n10762 ; n10763
g10700 and n6143 n8421 ; n10764
g10701 and n10763 n10764_not ; n10765
g10702 and a[8] n10765_not ; n10766
g10703 nor n10765 n10766 ; n10767
g10704 and a[8] n10766_not ; n10768
g10705 nor n10767 n10768 ; n10769
g10706 nor n10350 n10354 ; n10770
g10707 nor n10353 n10354 ; n10771
g10708 nor n10770 n10771 ; n10772
g10709 nor n10769 n10772 ; n10773
g10710 nor n10769 n10773 ; n10774
g10711 nor n10772 n10773 ; n10775
g10712 nor n10774 n10775 ; n10776
g10713 and n10251 n10348 ; n10777
g10714 nor n10349 n10777 ; n10778
g10715 and n2057_not n9331 ; n10779
g10716 and n2189_not n8418 ; n10780
g10717 and n2152_not n8860 ; n10781
g10718 nor n10780 n10781 ; n10782
g10719 and n10779_not n10782 ; n10783
g10720 and n8421_not n10783 ; n10784
g10721 and n6479_not n10783 ; n10785
g10722 nor n10784 n10785 ; n10786
g10723 and a[8] n10786_not ; n10787
g10724 and a[8]_not n10786 ; n10788
g10725 nor n10787 n10788 ; n10789
g10726 and n10778 n10789_not ; n10790
g10727 and n10344 n10346_not ; n10791
g10728 nor n10347 n10791 ; n10792
g10729 and n2152_not n9331 ; n10793
g10730 and n2291_not n8418 ; n10794
g10731 and n2189_not n8860 ; n10795
g10732 nor n10794 n10795 ; n10796
g10733 and n10793_not n10796 ; n10797
g10734 and n8421_not n10797 ; n10798
g10735 and n6492_not n10797 ; n10799
g10736 nor n10798 n10799 ; n10800
g10737 and a[8] n10800_not ; n10801
g10738 and a[8]_not n10800 ; n10802
g10739 nor n10801 n10802 ; n10803
g10740 and n10792 n10803_not ; n10804
g10741 and n10283 n10342 ; n10805
g10742 nor n10343 n10805 ; n10806
g10743 and n2189_not n9331 ; n10807
g10744 and n2388_not n8418 ; n10808
g10745 and n2291_not n8860 ; n10809
g10746 nor n10808 n10809 ; n10810
g10747 and n10807_not n10810 ; n10811
g10748 and n8421_not n10811 ; n10812
g10749 and n6122_not n10811 ; n10813
g10750 nor n10812 n10813 ; n10814
g10751 and a[8] n10814_not ; n10815
g10752 and a[8]_not n10814 ; n10816
g10753 nor n10815 n10816 ; n10817
g10754 and n10806 n10817_not ; n10818
g10755 and n2291_not n9331 ; n10819
g10756 and n2464_not n8418 ; n10820
g10757 and n2388_not n8860 ; n10821
g10758 nor n10820 n10821 ; n10822
g10759 and n10819_not n10822 ; n10823
g10760 and n6541 n8421 ; n10824
g10761 and n10823 n10824_not ; n10825
g10762 and a[8] n10825_not ; n10826
g10763 nor n10825 n10826 ; n10827
g10764 and a[8] n10826_not ; n10828
g10765 nor n10827 n10828 ; n10829
g10766 and n10338 n10340_not ; n10830
g10767 nor n10341 n10830 ; n10831
g10768 and n10829_not n10831 ; n10832
g10769 nor n10829 n10832 ; n10833
g10770 and n10831 n10832_not ; n10834
g10771 nor n10833 n10834 ; n10835
g10772 nor n10325 n10337 ; n10836
g10773 nor n10336 n10337 ; n10837
g10774 nor n10836 n10837 ; n10838
g10775 and n2388_not n9331 ; n10839
g10776 and n2533_not n8418 ; n10840
g10777 and n2464_not n8860 ; n10841
g10778 nor n10840 n10841 ; n10842
g10779 and n10839_not n10842 ; n10843
g10780 and n8421_not n10843 ; n10844
g10781 and n6591_not n10843 ; n10845
g10782 nor n10844 n10845 ; n10846
g10783 and a[8] n10846_not ; n10847
g10784 and a[8]_not n10846 ; n10848
g10785 nor n10847 n10848 ; n10849
g10786 nor n10838 n10849 ; n10850
g10787 and n2464_not n9331 ; n10851
g10788 and n2571_not n8418 ; n10852
g10789 and n2533_not n8860 ; n10853
g10790 nor n10852 n10853 ; n10854
g10791 and n10851_not n10854 ; n10855
g10792 and n6646 n8421 ; n10856
g10793 and n10855 n10856_not ; n10857
g10794 and a[8] n10857_not ; n10858
g10795 nor n10857 n10858 ; n10859
g10796 and a[8] n10858_not ; n10860
g10797 nor n10859 n10860 ; n10861
g10798 and n10309_not n10320 ; n10862
g10799 nor n10321 n10862 ; n10863
g10800 and n10861_not n10863 ; n10864
g10801 nor n10861 n10864 ; n10865
g10802 and n10863 n10864_not ; n10866
g10803 nor n10865 n10866 ; n10867
g10804 and n10306 n10308_not ; n10868
g10805 nor n10309 n10868 ; n10869
g10806 and n2533_not n9331 ; n10870
g10807 and n2674_not n8418 ; n10871
g10808 and n2571_not n8860 ; n10872
g10809 nor n10871 n10872 ; n10873
g10810 and n10870_not n10873 ; n10874
g10811 and n8421_not n10874 ; n10875
g10812 and n6695_not n10874 ; n10876
g10813 nor n10875 n10876 ; n10877
g10814 and a[8] n10877_not ; n10878
g10815 and a[8]_not n10877 ; n10879
g10816 nor n10878 n10879 ; n10880
g10817 and n10869 n10880_not ; n10881
g10818 and n2829_not n8860 ; n10882
g10819 and n2736_not n9331 ; n10883
g10820 nor n10882 n10883 ; n10884
g10821 and n7469_not n8421 ; n10885
g10822 and n10884 n10885_not ; n10886
g10823 and a[8] n10886_not ; n10887
g10824 and a[8] n10887_not ; n10888
g10825 nor n10886 n10887 ; n10889
g10826 nor n10888 n10889 ; n10890
g10827 nor n2829 n8416 ; n10891
g10828 and a[8] n10891_not ; n10892
g10829 and n10890_not n10892 ; n10893
g10830 and n2674_not n9331 ; n10894
g10831 and n2829_not n8418 ; n10895
g10832 and n2736_not n8860 ; n10896
g10833 nor n10895 n10896 ; n10897
g10834 and n10894_not n10897 ; n10898
g10835 and n8421_not n10898 ; n10899
g10836 and n6798_not n10898 ; n10900
g10837 nor n10899 n10900 ; n10901
g10838 and a[8] n10901_not ; n10902
g10839 and a[8]_not n10901 ; n10903
g10840 nor n10902 n10903 ; n10904
g10841 and n10893 n10904_not ; n10905
g10842 and n10307 n10905 ; n10906
g10843 and n10905 n10906_not ; n10907
g10844 and n10307 n10906_not ; n10908
g10845 nor n10907 n10908 ; n10909
g10846 and n2571_not n9331 ; n10910
g10847 and n2736_not n8418 ; n10911
g10848 and n2674_not n8860 ; n10912
g10849 nor n10911 n10912 ; n10913
g10850 and n10910_not n10913 ; n10914
g10851 and n6806 n8421 ; n10915
g10852 and n10914 n10915_not ; n10916
g10853 and a[8] n10916_not ; n10917
g10854 and a[8] n10917_not ; n10918
g10855 nor n10916 n10917 ; n10919
g10856 nor n10918 n10919 ; n10920
g10857 nor n10909 n10920 ; n10921
g10858 nor n10906 n10921 ; n10922
g10859 and n10869_not n10880 ; n10923
g10860 nor n10881 n10923 ; n10924
g10861 and n10922_not n10924 ; n10925
g10862 nor n10881 n10925 ; n10926
g10863 nor n10867 n10926 ; n10927
g10864 nor n10864 n10927 ; n10928
g10865 and n10838 n10849 ; n10929
g10866 nor n10850 n10929 ; n10930
g10867 and n10928_not n10930 ; n10931
g10868 nor n10850 n10931 ; n10932
g10869 nor n10835 n10932 ; n10933
g10870 nor n10832 n10933 ; n10934
g10871 and n10806 n10818_not ; n10935
g10872 nor n10817 n10818 ; n10936
g10873 nor n10935 n10936 ; n10937
g10874 nor n10934 n10937 ; n10938
g10875 nor n10818 n10938 ; n10939
g10876 and n10792 n10804_not ; n10940
g10877 nor n10803 n10804 ; n10941
g10878 nor n10940 n10941 ; n10942
g10879 nor n10939 n10942 ; n10943
g10880 nor n10804 n10943 ; n10944
g10881 and n10778_not n10789 ; n10945
g10882 nor n10790 n10945 ; n10946
g10883 and n10944_not n10946 ; n10947
g10884 nor n10790 n10947 ; n10948
g10885 nor n10776 n10948 ; n10949
g10886 nor n10773 n10949 ; n10950
g10887 nor n10758 n10950 ; n10951
g10888 nor n10755 n10951 ; n10952
g10889 nor n10740 n10952 ; n10953
g10890 nor n10737 n10953 ; n10954
g10891 and n10711 n10723_not ; n10955
g10892 nor n10722 n10723 ; n10956
g10893 nor n10955 n10956 ; n10957
g10894 nor n10954 n10957 ; n10958
g10895 nor n10723 n10958 ; n10959
g10896 and n10697 n10709_not ; n10960
g10897 nor n10708 n10709 ; n10961
g10898 nor n10960 n10961 ; n10962
g10899 nor n10959 n10962 ; n10963
g10900 nor n10709 n10963 ; n10964
g10901 and n10683_not n10694 ; n10965
g10902 nor n10695 n10965 ; n10966
g10903 and n10964_not n10966 ; n10967
g10904 nor n10695 n10967 ; n10968
g10905 nor n10681 n10968 ; n10969
g10906 nor n10678 n10969 ; n10970
g10907 nor n10663 n10970 ; n10971
g10908 nor n10660 n10971 ; n10972
g10909 nor n10645 n10972 ; n10973
g10910 nor n10642 n10973 ; n10974
g10911 and n10616 n10628_not ; n10975
g10912 nor n10627 n10628 ; n10976
g10913 nor n10975 n10976 ; n10977
g10914 nor n10974 n10977 ; n10978
g10915 nor n10628 n10978 ; n10979
g10916 and n10602 n10614_not ; n10980
g10917 nor n10613 n10614 ; n10981
g10918 nor n10980 n10981 ; n10982
g10919 nor n10979 n10982 ; n10983
g10920 nor n10614 n10983 ; n10984
g10921 and n10588_not n10599 ; n10985
g10922 nor n10600 n10985 ; n10986
g10923 and n10984_not n10986 ; n10987
g10924 nor n10600 n10987 ; n10988
g10925 nor n10586 n10988 ; n10989
g10926 nor n10583 n10989 ; n10990
g10927 nor n10568 n10990 ; n10991
g10928 nor n10565 n10991 ; n10992
g10929 and n10539 n10551_not ; n10993
g10930 nor n10550 n10551 ; n10994
g10931 nor n10993 n10994 ; n10995
g10932 nor n10992 n10995 ; n10996
g10933 nor n10551 n10996 ; n10997
g10934 and n10525 n10537_not ; n10998
g10935 nor n10536 n10537 ; n10999
g10936 nor n10998 n10999 ; n11000
g10937 nor n10997 n11000 ; n11001
g10938 nor n10537 n11001 ; n11002
g10939 and n10511 n10523_not ; n11003
g10940 nor n10522 n10523 ; n11004
g10941 nor n11003 n11004 ; n11005
g10942 nor n11002 n11005 ; n11006
g10943 nor n10523 n11006 ; n11007
g10944 and n10497 n10509_not ; n11008
g10945 nor n10508 n10509 ; n11009
g10946 nor n11008 n11009 ; n11010
g10947 nor n11007 n11010 ; n11011
g10948 nor n10509 n11011 ; n11012
g10949 and n10483 n10495_not ; n11013
g10950 nor n10494 n10495 ; n11014
g10951 nor n11013 n11014 ; n11015
g10952 nor n11012 n11015 ; n11016
g10953 nor n10495 n11016 ; n11017
g10954 and n10469 n10481_not ; n11018
g10955 nor n10480 n10481 ; n11019
g10956 nor n11018 n11019 ; n11020
g10957 nor n11017 n11020 ; n11021
g10958 nor n10481 n11021 ; n11022
g10959 and n10455 n10467_not ; n11023
g10960 nor n10466 n10467 ; n11024
g10961 nor n11023 n11024 ; n11025
g10962 nor n11022 n11025 ; n11026
g10963 nor n10467 n11026 ; n11027
g10964 and n10427 n10429_not ; n11028
g10965 and n10428_not n11028 ; n11029
g10966 nor n10431 n11029 ; n11030
g10967 and n11027_not n11030 ; n11031
g10968 and n71 n4515_not ; n11032
g10969 and n4045_not n9867 ; n11033
g10970 and n3877_not n10434 ; n11034
g10971 nor n11033 n11034 ; n11035
g10972 and n11032_not n11035 ; n11036
g10973 and n4715 n9870 ; n11037
g10974 and n11036 n11037_not ; n11038
g10975 and a[5] n11038_not ; n11039
g10976 nor n11038 n11039 ; n11040
g10977 and a[5] n11039_not ; n11041
g10978 nor n11040 n11041 ; n11042
g10979 nor n11027 n11031 ; n11043
g10980 and n11030 n11031_not ; n11044
g10981 nor n11043 n11044 ; n11045
g10982 nor n11042 n11045 ; n11046
g10983 nor n11031 n11046 ; n11047
g10984 and n10446 n10448_not ; n11048
g10985 nor n10449 n11048 ; n11049
g10986 and n11047_not n11049 ; n11050
g10987 and a[1] a[2]_not ; n11051
g10988 and a[1]_not a[2] ; n11052
g10989 nor n11051 n11052 ; n11053
g10990 nor a[0] a[1] ; n11054
g10991 and n11053_not n11054 ; n11055
g10992 and n4515_not n11055 ; n11056
g10993 and a[0] n11053_not ; n11057
g10994 and n4522 n11057 ; n11058
g10995 nor n11056 n11058 ; n11059
g10996 and a[2] n11059_not ; n11060
g10997 nor n11059 n11060 ; n11061
g10998 and a[2] n11060_not ; n11062
g10999 nor n11061 n11062 ; n11063
g11000 and n71 n3877_not ; n11064
g11001 and n3964_not n9867 ; n11065
g11002 and n4045_not n10434 ; n11066
g11003 nor n11065 n11066 ; n11067
g11004 and n11064_not n11067 ; n11068
g11005 and n4067 n9870 ; n11069
g11006 and n11068 n11069_not ; n11070
g11007 and a[5] n11070_not ; n11071
g11008 and a[5] n11071_not ; n11072
g11009 nor n11070 n11071 ; n11073
g11010 nor n11072 n11073 ; n11074
g11011 nor n11063 n11074 ; n11075
g11012 nor n11063 n11075 ; n11076
g11013 nor n11074 n11075 ; n11077
g11014 nor n11076 n11077 ; n11078
g11015 nor n11022 n11026 ; n11079
g11016 nor n11025 n11026 ; n11080
g11017 nor n11079 n11080 ; n11081
g11018 nor n11078 n11081 ; n11082
g11019 nor n11075 n11082 ; n11083
g11020 and n11042 n11044_not ; n11084
g11021 and n11043_not n11084 ; n11085
g11022 nor n11046 n11085 ; n11086
g11023 and n11083_not n11086 ; n11087
g11024 nor n11078 n11082 ; n11088
g11025 nor n11081 n11082 ; n11089
g11026 nor n11088 n11089 ; n11090
g11027 and n71 n4045_not ; n11091
g11028 and n3805_not n9867 ; n11092
g11029 and n3964_not n10434 ; n11093
g11030 nor n11092 n11093 ; n11094
g11031 and n11091_not n11094 ; n11095
g11032 and n4477 n9870 ; n11096
g11033 and n11095 n11096_not ; n11097
g11034 and a[5] n11097_not ; n11098
g11035 nor n11097 n11098 ; n11099
g11036 and a[5] n11098_not ; n11100
g11037 nor n11099 n11100 ; n11101
g11038 nor n11017 n11021 ; n11102
g11039 nor n11020 n11021 ; n11103
g11040 nor n11102 n11103 ; n11104
g11041 nor n11101 n11104 ; n11105
g11042 nor n11101 n11105 ; n11106
g11043 nor n11104 n11105 ; n11107
g11044 nor n11106 n11107 ; n11108
g11045 and n71 n3964_not ; n11109
g11046 and n3456_not n9867 ; n11110
g11047 and n3805_not n10434 ; n11111
g11048 nor n11110 n11111 ; n11112
g11049 and n11109_not n11112 ; n11113
g11050 and n4558 n9870 ; n11114
g11051 and n11113 n11114_not ; n11115
g11052 and a[5] n11115_not ; n11116
g11053 nor n11115 n11116 ; n11117
g11054 and a[5] n11116_not ; n11118
g11055 nor n11117 n11118 ; n11119
g11056 nor n11012 n11016 ; n11120
g11057 nor n11015 n11016 ; n11121
g11058 nor n11120 n11121 ; n11122
g11059 nor n11119 n11122 ; n11123
g11060 nor n11119 n11123 ; n11124
g11061 nor n11122 n11123 ; n11125
g11062 nor n11124 n11125 ; n11126
g11063 and n71 n3805_not ; n11127
g11064 and n3605_not n9867 ; n11128
g11065 and n3456_not n10434 ; n11129
g11066 nor n11128 n11129 ; n11130
g11067 and n11127_not n11130 ; n11131
g11068 and n3818 n9870 ; n11132
g11069 and n11131 n11132_not ; n11133
g11070 and a[5] n11133_not ; n11134
g11071 nor n11133 n11134 ; n11135
g11072 and a[5] n11134_not ; n11136
g11073 nor n11135 n11136 ; n11137
g11074 nor n11007 n11011 ; n11138
g11075 nor n11010 n11011 ; n11139
g11076 nor n11138 n11139 ; n11140
g11077 nor n11137 n11140 ; n11141
g11078 nor n11137 n11141 ; n11142
g11079 nor n11140 n11141 ; n11143
g11080 nor n11142 n11143 ; n11144
g11081 and n71 n3456_not ; n11145
g11082 and n3539_not n9867 ; n11146
g11083 and n3605_not n10434 ; n11147
g11084 nor n11146 n11147 ; n11148
g11085 and n11145_not n11148 ; n11149
g11086 and n3627 n9870 ; n11150
g11087 and n11149 n11150_not ; n11151
g11088 and a[5] n11151_not ; n11152
g11089 nor n11151 n11152 ; n11153
g11090 and a[5] n11152_not ; n11154
g11091 nor n11153 n11154 ; n11155
g11092 nor n11002 n11006 ; n11156
g11093 nor n11005 n11006 ; n11157
g11094 nor n11156 n11157 ; n11158
g11095 nor n11155 n11158 ; n11159
g11096 nor n11155 n11159 ; n11160
g11097 nor n11158 n11159 ; n11161
g11098 nor n11160 n11161 ; n11162
g11099 and n71 n3605_not ; n11163
g11100 and n3012_not n9867 ; n11164
g11101 and n3539_not n10434 ; n11165
g11102 nor n11164 n11165 ; n11166
g11103 and n11163_not n11166 ; n11167
g11104 and n4084 n9870 ; n11168
g11105 and n11167 n11168_not ; n11169
g11106 and a[5] n11169_not ; n11170
g11107 nor n11169 n11170 ; n11171
g11108 and a[5] n11170_not ; n11172
g11109 nor n11171 n11172 ; n11173
g11110 nor n10997 n11001 ; n11174
g11111 nor n11000 n11001 ; n11175
g11112 nor n11174 n11175 ; n11176
g11113 nor n11173 n11176 ; n11177
g11114 nor n11173 n11177 ; n11178
g11115 nor n11176 n11177 ; n11179
g11116 nor n11178 n11179 ; n11180
g11117 and n71 n3539_not ; n11181
g11118 and n392_not n9867 ; n11182
g11119 and n3012_not n10434 ; n11183
g11120 nor n11182 n11183 ; n11184
g11121 and n11181_not n11184 ; n11185
g11122 and n3715 n9870 ; n11186
g11123 and n11185 n11186_not ; n11187
g11124 and a[5] n11187_not ; n11188
g11125 nor n11187 n11188 ; n11189
g11126 and a[5] n11188_not ; n11190
g11127 nor n11189 n11190 ; n11191
g11128 nor n10992 n10996 ; n11192
g11129 nor n10995 n10996 ; n11193
g11130 nor n11192 n11193 ; n11194
g11131 nor n11191 n11194 ; n11195
g11132 nor n11191 n11195 ; n11196
g11133 nor n11194 n11195 ; n11197
g11134 nor n11196 n11197 ; n11198
g11135 and n10568 n10990 ; n11199
g11136 nor n10991 n11199 ; n11200
g11137 and n71 n3012_not ; n11201
g11138 and n587_not n9867 ; n11202
g11139 and n392_not n10434 ; n11203
g11140 nor n11202 n11203 ; n11204
g11141 and n11201_not n11204 ; n11205
g11142 and n9870_not n11205 ; n11206
g11143 and n3018_not n11205 ; n11207
g11144 nor n11206 n11207 ; n11208
g11145 and a[5] n11208_not ; n11209
g11146 and a[5]_not n11208 ; n11210
g11147 nor n11209 n11210 ; n11211
g11148 and n11200 n11211_not ; n11212
g11149 and n10586 n10988 ; n11213
g11150 nor n10989 n11213 ; n11214
g11151 and n71 n392_not ; n11215
g11152 and n710_not n9867 ; n11216
g11153 and n587_not n10434 ; n11217
g11154 nor n11216 n11217 ; n11218
g11155 and n11215_not n11218 ; n11219
g11156 and n9870_not n11219 ; n11220
g11157 and n3347_not n11219 ; n11221
g11158 nor n11220 n11221 ; n11222
g11159 and a[5] n11222_not ; n11223
g11160 and a[5]_not n11222 ; n11224
g11161 nor n11223 n11224 ; n11225
g11162 and n11214 n11225_not ; n11226
g11163 and n71 n587_not ; n11227
g11164 and n867_not n9867 ; n11228
g11165 and n710_not n10434 ; n11229
g11166 nor n11228 n11229 ; n11230
g11167 and n11227_not n11230 ; n11231
g11168 and n3331 n9870 ; n11232
g11169 and n11231 n11232_not ; n11233
g11170 and a[5] n11233_not ; n11234
g11171 nor n11233 n11234 ; n11235
g11172 and a[5] n11234_not ; n11236
g11173 nor n11235 n11236 ; n11237
g11174 and n10984 n10986_not ; n11238
g11175 nor n10987 n11238 ; n11239
g11176 and n11237_not n11239 ; n11240
g11177 nor n11237 n11240 ; n11241
g11178 and n11239 n11240_not ; n11242
g11179 nor n11241 n11242 ; n11243
g11180 and n71 n710_not ; n11244
g11181 and n958_not n9867 ; n11245
g11182 and n867_not n10434 ; n11246
g11183 nor n11245 n11246 ; n11247
g11184 and n11244_not n11247 ; n11248
g11185 and n4179 n9870 ; n11249
g11186 and n11248 n11249_not ; n11250
g11187 and a[5] n11250_not ; n11251
g11188 nor n11250 n11251 ; n11252
g11189 and a[5] n11251_not ; n11253
g11190 nor n11252 n11253 ; n11254
g11191 nor n10979 n10983 ; n11255
g11192 nor n10982 n10983 ; n11256
g11193 nor n11255 n11256 ; n11257
g11194 nor n11254 n11257 ; n11258
g11195 nor n11254 n11258 ; n11259
g11196 nor n11257 n11258 ; n11260
g11197 nor n11259 n11260 ; n11261
g11198 and n71 n867_not ; n11262
g11199 and n1060_not n9867 ; n11263
g11200 and n958_not n10434 ; n11264
g11201 nor n11263 n11264 ; n11265
g11202 and n11262_not n11265 ; n11266
g11203 and n4204 n9870 ; n11267
g11204 and n11266 n11267_not ; n11268
g11205 and a[5] n11268_not ; n11269
g11206 nor n11268 n11269 ; n11270
g11207 and a[5] n11269_not ; n11271
g11208 nor n11270 n11271 ; n11272
g11209 nor n10974 n10978 ; n11273
g11210 nor n10977 n10978 ; n11274
g11211 nor n11273 n11274 ; n11275
g11212 nor n11272 n11275 ; n11276
g11213 nor n11272 n11276 ; n11277
g11214 nor n11275 n11276 ; n11278
g11215 nor n11277 n11278 ; n11279
g11216 and n10645 n10972 ; n11280
g11217 nor n10973 n11280 ; n11281
g11218 and n71 n958_not ; n11282
g11219 and n1178_not n9867 ; n11283
g11220 and n1060_not n10434 ; n11284
g11221 nor n11283 n11284 ; n11285
g11222 and n11282_not n11285 ; n11286
g11223 and n9870_not n11286 ; n11287
g11224 and n4633_not n11286 ; n11288
g11225 nor n11287 n11288 ; n11289
g11226 and a[5] n11289_not ; n11290
g11227 and a[5]_not n11289 ; n11291
g11228 nor n11290 n11291 ; n11292
g11229 and n11281 n11292_not ; n11293
g11230 and n10663 n10970 ; n11294
g11231 nor n10971 n11294 ; n11295
g11232 and n71 n1060_not ; n11296
g11233 and n1235_not n9867 ; n11297
g11234 and n1178_not n10434 ; n11298
g11235 nor n11297 n11298 ; n11299
g11236 and n11296_not n11299 ; n11300
g11237 and n9870_not n11300 ; n11301
g11238 and n4429_not n11300 ; n11302
g11239 nor n11301 n11302 ; n11303
g11240 and a[5] n11303_not ; n11304
g11241 and a[5]_not n11303 ; n11305
g11242 nor n11304 n11305 ; n11306
g11243 and n11295 n11306_not ; n11307
g11244 and n10681 n10968 ; n11308
g11245 nor n10969 n11308 ; n11309
g11246 and n71 n1178_not ; n11310
g11247 and n1364_not n9867 ; n11311
g11248 and n1235_not n10434 ; n11312
g11249 nor n11311 n11312 ; n11313
g11250 and n11310_not n11313 ; n11314
g11251 and n9870_not n11314 ; n11315
g11252 and n4861_not n11314 ; n11316
g11253 nor n11315 n11316 ; n11317
g11254 and a[5] n11317_not ; n11318
g11255 and a[5]_not n11317 ; n11319
g11256 nor n11318 n11319 ; n11320
g11257 and n11309 n11320_not ; n11321
g11258 and n71 n1235_not ; n11322
g11259 and n1472_not n9867 ; n11323
g11260 and n1364_not n10434 ; n11324
g11261 nor n11323 n11324 ; n11325
g11262 and n11322_not n11325 ; n11326
g11263 and n4848 n9870 ; n11327
g11264 and n11326 n11327_not ; n11328
g11265 and a[5] n11328_not ; n11329
g11266 nor n11328 n11329 ; n11330
g11267 and a[5] n11329_not ; n11331
g11268 nor n11330 n11331 ; n11332
g11269 and n10964 n10966_not ; n11333
g11270 nor n10967 n11333 ; n11334
g11271 and n11332_not n11334 ; n11335
g11272 nor n11332 n11335 ; n11336
g11273 and n11334 n11335_not ; n11337
g11274 nor n11336 n11337 ; n11338
g11275 and n71 n1364_not ; n11339
g11276 and n1572_not n9867 ; n11340
g11277 and n1472_not n10434 ; n11341
g11278 nor n11340 n11341 ; n11342
g11279 and n11339_not n11342 ; n11343
g11280 and n5114 n9870 ; n11344
g11281 and n11343 n11344_not ; n11345
g11282 and a[5] n11345_not ; n11346
g11283 nor n11345 n11346 ; n11347
g11284 and a[5] n11346_not ; n11348
g11285 nor n11347 n11348 ; n11349
g11286 nor n10959 n10963 ; n11350
g11287 nor n10962 n10963 ; n11351
g11288 nor n11350 n11351 ; n11352
g11289 nor n11349 n11352 ; n11353
g11290 nor n11349 n11353 ; n11354
g11291 nor n11352 n11353 ; n11355
g11292 nor n11354 n11355 ; n11356
g11293 and n71 n1472_not ; n11357
g11294 and n1665_not n9867 ; n11358
g11295 and n1572_not n10434 ; n11359
g11296 nor n11358 n11359 ; n11360
g11297 and n11357_not n11360 ; n11361
g11298 and n5139 n9870 ; n11362
g11299 and n11361 n11362_not ; n11363
g11300 and a[5] n11363_not ; n11364
g11301 nor n11363 n11364 ; n11365
g11302 and a[5] n11364_not ; n11366
g11303 nor n11365 n11366 ; n11367
g11304 nor n10954 n10958 ; n11368
g11305 nor n10957 n10958 ; n11369
g11306 nor n11368 n11369 ; n11370
g11307 nor n11367 n11370 ; n11371
g11308 nor n11367 n11371 ; n11372
g11309 nor n11370 n11371 ; n11373
g11310 nor n11372 n11373 ; n11374
g11311 and n10740 n10952 ; n11375
g11312 nor n10953 n11375 ; n11376
g11313 and n71 n1572_not ; n11377
g11314 and n1779_not n9867 ; n11378
g11315 and n1665_not n10434 ; n11379
g11316 nor n11378 n11379 ; n11380
g11317 and n11377_not n11380 ; n11381
g11318 and n9870_not n11381 ; n11382
g11319 and n5561_not n11381 ; n11383
g11320 nor n11382 n11383 ; n11384
g11321 and a[5] n11384_not ; n11385
g11322 and a[5]_not n11384 ; n11386
g11323 nor n11385 n11386 ; n11387
g11324 and n11376 n11387_not ; n11388
g11325 and n10758 n10950 ; n11389
g11326 nor n10951 n11389 ; n11390
g11327 and n71 n1665_not ; n11391
g11328 and n1877_not n9867 ; n11392
g11329 and n1779_not n10434 ; n11393
g11330 nor n11392 n11393 ; n11394
g11331 and n11391_not n11394 ; n11395
g11332 and n9870_not n11395 ; n11396
g11333 and n5328_not n11395 ; n11397
g11334 nor n11396 n11397 ; n11398
g11335 and a[5] n11398_not ; n11399
g11336 and a[5]_not n11398 ; n11400
g11337 nor n11399 n11400 ; n11401
g11338 and n11390 n11401_not ; n11402
g11339 and n10776 n10948 ; n11403
g11340 nor n10949 n11403 ; n11404
g11341 and n71 n1779_not ; n11405
g11342 and n1913_not n9867 ; n11406
g11343 and n1877_not n10434 ; n11407
g11344 nor n11406 n11407 ; n11408
g11345 and n11405_not n11408 ; n11409
g11346 and n9870_not n11409 ; n11410
g11347 and n5851_not n11409 ; n11411
g11348 nor n11410 n11411 ; n11412
g11349 and a[5] n11412_not ; n11413
g11350 and a[5]_not n11412 ; n11414
g11351 nor n11413 n11414 ; n11415
g11352 and n11404 n11415_not ; n11416
g11353 and n71 n1877_not ; n11417
g11354 and n1992_not n9867 ; n11418
g11355 and n1913_not n10434 ; n11419
g11356 nor n11418 n11419 ; n11420
g11357 and n11417_not n11420 ; n11421
g11358 and n6007 n9870 ; n11422
g11359 and n11421 n11422_not ; n11423
g11360 and a[5] n11423_not ; n11424
g11361 nor n11423 n11424 ; n11425
g11362 and a[5] n11424_not ; n11426
g11363 nor n11425 n11426 ; n11427
g11364 and n10944 n10946_not ; n11428
g11365 nor n10947 n11428 ; n11429
g11366 and n11427_not n11429 ; n11430
g11367 nor n11427 n11430 ; n11431
g11368 and n11429 n11430_not ; n11432
g11369 nor n11431 n11432 ; n11433
g11370 and n71 n1913_not ; n11434
g11371 and n2057_not n9867 ; n11435
g11372 and n1992_not n10434 ; n11436
g11373 nor n11435 n11436 ; n11437
g11374 and n11434_not n11437 ; n11438
g11375 and n5834 n9870 ; n11439
g11376 and n11438 n11439_not ; n11440
g11377 and a[5] n11440_not ; n11441
g11378 nor n11440 n11441 ; n11442
g11379 and a[5] n11441_not ; n11443
g11380 nor n11442 n11443 ; n11444
g11381 nor n10939 n10943 ; n11445
g11382 nor n10942 n10943 ; n11446
g11383 nor n11445 n11446 ; n11447
g11384 nor n11444 n11447 ; n11448
g11385 nor n11444 n11448 ; n11449
g11386 nor n11447 n11448 ; n11450
g11387 nor n11449 n11450 ; n11451
g11388 and n71 n1992_not ; n11452
g11389 and n2152_not n9867 ; n11453
g11390 and n2057_not n10434 ; n11454
g11391 nor n11453 n11454 ; n11455
g11392 and n11452_not n11455 ; n11456
g11393 and n6143 n9870 ; n11457
g11394 and n11456 n11457_not ; n11458
g11395 and a[5] n11458_not ; n11459
g11396 nor n11458 n11459 ; n11460
g11397 and a[5] n11459_not ; n11461
g11398 nor n11460 n11461 ; n11462
g11399 nor n10934 n10938 ; n11463
g11400 nor n10937 n10938 ; n11464
g11401 nor n11463 n11464 ; n11465
g11402 nor n11462 n11465 ; n11466
g11403 nor n11462 n11466 ; n11467
g11404 nor n11465 n11466 ; n11468
g11405 nor n11467 n11468 ; n11469
g11406 and n10835 n10932 ; n11470
g11407 nor n10933 n11470 ; n11471
g11408 and n71 n2057_not ; n11472
g11409 and n2189_not n9867 ; n11473
g11410 and n2152_not n10434 ; n11474
g11411 nor n11473 n11474 ; n11475
g11412 and n11472_not n11475 ; n11476
g11413 and n9870_not n11476 ; n11477
g11414 and n6479_not n11476 ; n11478
g11415 nor n11477 n11478 ; n11479
g11416 and a[5] n11479_not ; n11480
g11417 and a[5]_not n11479 ; n11481
g11418 nor n11480 n11481 ; n11482
g11419 and n11471 n11482_not ; n11483
g11420 and n10928 n10930_not ; n11484
g11421 nor n10931 n11484 ; n11485
g11422 and n71 n2152_not ; n11486
g11423 and n2291_not n9867 ; n11487
g11424 and n2189_not n10434 ; n11488
g11425 nor n11487 n11488 ; n11489
g11426 and n11486_not n11489 ; n11490
g11427 and n9870_not n11490 ; n11491
g11428 and n6492_not n11490 ; n11492
g11429 nor n11491 n11492 ; n11493
g11430 and a[5] n11493_not ; n11494
g11431 and a[5]_not n11493 ; n11495
g11432 nor n11494 n11495 ; n11496
g11433 and n11485 n11496_not ; n11497
g11434 and n10867 n10926 ; n11498
g11435 nor n10927 n11498 ; n11499
g11436 and n71 n2189_not ; n11500
g11437 and n2388_not n9867 ; n11501
g11438 and n2291_not n10434 ; n11502
g11439 nor n11501 n11502 ; n11503
g11440 and n11500_not n11503 ; n11504
g11441 and n9870_not n11504 ; n11505
g11442 and n6122_not n11504 ; n11506
g11443 nor n11505 n11506 ; n11507
g11444 and a[5] n11507_not ; n11508
g11445 and a[5]_not n11507 ; n11509
g11446 nor n11508 n11509 ; n11510
g11447 and n11499 n11510_not ; n11511
g11448 and n71 n2291_not ; n11512
g11449 and n2464_not n9867 ; n11513
g11450 and n2388_not n10434 ; n11514
g11451 nor n11513 n11514 ; n11515
g11452 and n11512_not n11515 ; n11516
g11453 and n6541 n9870 ; n11517
g11454 and n11516 n11517_not ; n11518
g11455 and a[5] n11518_not ; n11519
g11456 nor n11518 n11519 ; n11520
g11457 and a[5] n11519_not ; n11521
g11458 nor n11520 n11521 ; n11522
g11459 and n10922 n10924_not ; n11523
g11460 nor n10925 n11523 ; n11524
g11461 and n11522_not n11524 ; n11525
g11462 nor n11522 n11525 ; n11526
g11463 and n11524 n11525_not ; n11527
g11464 nor n11526 n11527 ; n11528
g11465 nor n10909 n10921 ; n11529
g11466 nor n10920 n10921 ; n11530
g11467 nor n11529 n11530 ; n11531
g11468 and n71 n2388_not ; n11532
g11469 and n2533_not n9867 ; n11533
g11470 and n2464_not n10434 ; n11534
g11471 nor n11533 n11534 ; n11535
g11472 and n11532_not n11535 ; n11536
g11473 and n9870_not n11536 ; n11537
g11474 and n6591_not n11536 ; n11538
g11475 nor n11537 n11538 ; n11539
g11476 and a[5] n11539_not ; n11540
g11477 and a[5]_not n11539 ; n11541
g11478 nor n11540 n11541 ; n11542
g11479 nor n11531 n11542 ; n11543
g11480 and n71 n2464_not ; n11544
g11481 and n2571_not n9867 ; n11545
g11482 and n2533_not n10434 ; n11546
g11483 nor n11545 n11546 ; n11547
g11484 and n11544_not n11547 ; n11548
g11485 and n6646 n9870 ; n11549
g11486 and n11548 n11549_not ; n11550
g11487 and a[5] n11550_not ; n11551
g11488 nor n11550 n11551 ; n11552
g11489 and a[5] n11551_not ; n11553
g11490 nor n11552 n11553 ; n11554
g11491 and n10893_not n10904 ; n11555
g11492 nor n10905 n11555 ; n11556
g11493 and n11554_not n11556 ; n11557
g11494 nor n11554 n11557 ; n11558
g11495 and n11556 n11557_not ; n11559
g11496 nor n11558 n11559 ; n11560
g11497 and n10890 n10892_not ; n11561
g11498 nor n10893 n11561 ; n11562
g11499 and n71 n2533_not ; n11563
g11500 and n2674_not n9867 ; n11564
g11501 and n2571_not n10434 ; n11565
g11502 nor n11564 n11565 ; n11566
g11503 and n11563_not n11566 ; n11567
g11504 and n9870_not n11567 ; n11568
g11505 and n6695_not n11567 ; n11569
g11506 nor n11568 n11569 ; n11570
g11507 and a[5] n11570_not ; n11571
g11508 and a[5]_not n11570 ; n11572
g11509 nor n11571 n11572 ; n11573
g11510 and n11562 n11573_not ; n11574
g11511 and n2829_not n10434 ; n11575
g11512 and n71 n2736_not ; n11576
g11513 nor n11575 n11576 ; n11577
g11514 and n7469_not n9870 ; n11578
g11515 and n11577 n11578_not ; n11579
g11516 and a[5] n11579_not ; n11580
g11517 and a[5] n11580_not ; n11581
g11518 nor n11579 n11580 ; n11582
g11519 nor n11581 n11582 ; n11583
g11520 nor n70 n2829 ; n11584
g11521 and a[5] n11584_not ; n11585
g11522 and n11583_not n11585 ; n11586
g11523 and n71 n2674_not ; n11587
g11524 and n2829_not n9867 ; n11588
g11525 and n2736_not n10434 ; n11589
g11526 nor n11588 n11589 ; n11590
g11527 and n11587_not n11590 ; n11591
g11528 and n9870_not n11591 ; n11592
g11529 and n6798_not n11591 ; n11593
g11530 nor n11592 n11593 ; n11594
g11531 and a[5] n11594_not ; n11595
g11532 and a[5]_not n11594 ; n11596
g11533 nor n11595 n11596 ; n11597
g11534 and n11586 n11597_not ; n11598
g11535 and n10891 n11598 ; n11599
g11536 and n11598 n11599_not ; n11600
g11537 and n10891 n11599_not ; n11601
g11538 nor n11600 n11601 ; n11602
g11539 and n71 n2571_not ; n11603
g11540 and n2736_not n9867 ; n11604
g11541 and n2674_not n10434 ; n11605
g11542 nor n11604 n11605 ; n11606
g11543 and n11603_not n11606 ; n11607
g11544 and n6806 n9870 ; n11608
g11545 and n11607 n11608_not ; n11609
g11546 and a[5] n11609_not ; n11610
g11547 and a[5] n11610_not ; n11611
g11548 nor n11609 n11610 ; n11612
g11549 nor n11611 n11612 ; n11613
g11550 nor n11602 n11613 ; n11614
g11551 nor n11599 n11614 ; n11615
g11552 and n11562_not n11573 ; n11616
g11553 nor n11574 n11616 ; n11617
g11554 and n11615_not n11617 ; n11618
g11555 nor n11574 n11618 ; n11619
g11556 nor n11560 n11619 ; n11620
g11557 nor n11557 n11620 ; n11621
g11558 and n11531 n11542 ; n11622
g11559 nor n11543 n11622 ; n11623
g11560 and n11621_not n11623 ; n11624
g11561 nor n11543 n11624 ; n11625
g11562 nor n11528 n11625 ; n11626
g11563 nor n11525 n11626 ; n11627
g11564 and n11499 n11511_not ; n11628
g11565 nor n11510 n11511 ; n11629
g11566 nor n11628 n11629 ; n11630
g11567 nor n11627 n11630 ; n11631
g11568 nor n11511 n11631 ; n11632
g11569 and n11485 n11497_not ; n11633
g11570 nor n11496 n11497 ; n11634
g11571 nor n11633 n11634 ; n11635
g11572 nor n11632 n11635 ; n11636
g11573 nor n11497 n11636 ; n11637
g11574 and n11471_not n11482 ; n11638
g11575 nor n11483 n11638 ; n11639
g11576 and n11637_not n11639 ; n11640
g11577 nor n11483 n11640 ; n11641
g11578 nor n11469 n11641 ; n11642
g11579 nor n11466 n11642 ; n11643
g11580 nor n11451 n11643 ; n11644
g11581 nor n11448 n11644 ; n11645
g11582 nor n11433 n11645 ; n11646
g11583 nor n11430 n11646 ; n11647
g11584 and n11404 n11416_not ; n11648
g11585 nor n11415 n11416 ; n11649
g11586 nor n11648 n11649 ; n11650
g11587 nor n11647 n11650 ; n11651
g11588 nor n11416 n11651 ; n11652
g11589 and n11390 n11402_not ; n11653
g11590 nor n11401 n11402 ; n11654
g11591 nor n11653 n11654 ; n11655
g11592 nor n11652 n11655 ; n11656
g11593 nor n11402 n11656 ; n11657
g11594 and n11376_not n11387 ; n11658
g11595 nor n11388 n11658 ; n11659
g11596 and n11657_not n11659 ; n11660
g11597 nor n11388 n11660 ; n11661
g11598 nor n11374 n11661 ; n11662
g11599 nor n11371 n11662 ; n11663
g11600 nor n11356 n11663 ; n11664
g11601 nor n11353 n11664 ; n11665
g11602 nor n11338 n11665 ; n11666
g11603 nor n11335 n11666 ; n11667
g11604 and n11309 n11321_not ; n11668
g11605 nor n11320 n11321 ; n11669
g11606 nor n11668 n11669 ; n11670
g11607 nor n11667 n11670 ; n11671
g11608 nor n11321 n11671 ; n11672
g11609 and n11295 n11307_not ; n11673
g11610 nor n11306 n11307 ; n11674
g11611 nor n11673 n11674 ; n11675
g11612 nor n11672 n11675 ; n11676
g11613 nor n11307 n11676 ; n11677
g11614 and n11281_not n11292 ; n11678
g11615 nor n11293 n11678 ; n11679
g11616 and n11677_not n11679 ; n11680
g11617 nor n11293 n11680 ; n11681
g11618 nor n11279 n11681 ; n11682
g11619 nor n11276 n11682 ; n11683
g11620 nor n11261 n11683 ; n11684
g11621 nor n11258 n11684 ; n11685
g11622 nor n11243 n11685 ; n11686
g11623 nor n11240 n11686 ; n11687
g11624 and n11214 n11226_not ; n11688
g11625 nor n11225 n11226 ; n11689
g11626 nor n11688 n11689 ; n11690
g11627 nor n11687 n11690 ; n11691
g11628 nor n11226 n11691 ; n11692
g11629 and n11200_not n11211 ; n11693
g11630 nor n11212 n11693 ; n11694
g11631 and n11692_not n11694 ; n11695
g11632 nor n11212 n11695 ; n11696
g11633 nor n11198 n11696 ; n11697
g11634 nor n11195 n11697 ; n11698
g11635 nor n11180 n11698 ; n11699
g11636 nor n11177 n11699 ; n11700
g11637 nor n11162 n11700 ; n11701
g11638 nor n11159 n11701 ; n11702
g11639 nor n11144 n11702 ; n11703
g11640 nor n11141 n11703 ; n11704
g11641 nor n11126 n11704 ; n11705
g11642 nor n11123 n11705 ; n11706
g11643 nor n11108 n11706 ; n11707
g11644 nor n11105 n11707 ; n11708
g11645 nor n11090 n11708 ; n11709
g11646 and n11090 n11708 ; n11710
g11647 nor n11709 n11710 ; n11711
g11648 and n11108 n11706 ; n11712
g11649 nor n11707 n11712 ; n11713
g11650 and n3877_not n11055 ; n11714
g11651 and a[0]_not a[1] ; n11715
g11652 and n4515_not n11715 ; n11716
g11653 nor n11714 n11716 ; n11717
g11654 and n11057_not n11717 ; n11718
g11655 and n4609_not n11717 ; n11719
g11656 nor n11718 n11719 ; n11720
g11657 and a[2] n11720_not ; n11721
g11658 and a[2]_not n11720 ; n11722
g11659 nor n11721 n11722 ; n11723
g11660 and n11713 n11723_not ; n11724
g11661 and n11126 n11704 ; n11725
g11662 nor n11705 n11725 ; n11726
g11663 and a[0] n11053 ; n11727
g11664 and n4515_not n11727 ; n11728
g11665 and n4045_not n11055 ; n11729
g11666 and n3877_not n11715 ; n11730
g11667 nor n11729 n11730 ; n11731
g11668 and n11728_not n11731 ; n11732
g11669 and n11057_not n11732 ; n11733
g11670 and n4715_not n11732 ; n11734
g11671 nor n11733 n11734 ; n11735
g11672 and a[2] n11735_not ; n11736
g11673 and a[2]_not n11735 ; n11737
g11674 nor n11736 n11737 ; n11738
g11675 and n11726 n11738_not ; n11739
g11676 and n11144 n11702 ; n11740
g11677 nor n11703 n11740 ; n11741
g11678 and n3877_not n11727 ; n11742
g11679 and n3964_not n11055 ; n11743
g11680 and n4045_not n11715 ; n11744
g11681 nor n11743 n11744 ; n11745
g11682 and n11742_not n11745 ; n11746
g11683 and n11057_not n11746 ; n11747
g11684 and n4067_not n11746 ; n11748
g11685 nor n11747 n11748 ; n11749
g11686 and a[2] n11749_not ; n11750
g11687 and a[2]_not n11749 ; n11751
g11688 nor n11750 n11751 ; n11752
g11689 and n11741 n11752_not ; n11753
g11690 and n11162 n11700 ; n11754
g11691 nor n11701 n11754 ; n11755
g11692 and n4045_not n11727 ; n11756
g11693 and n3805_not n11055 ; n11757
g11694 and n3964_not n11715 ; n11758
g11695 nor n11757 n11758 ; n11759
g11696 and n11756_not n11759 ; n11760
g11697 and n11057_not n11760 ; n11761
g11698 and n4477_not n11760 ; n11762
g11699 nor n11761 n11762 ; n11763
g11700 and a[2] n11763_not ; n11764
g11701 and a[2]_not n11763 ; n11765
g11702 nor n11764 n11765 ; n11766
g11703 and n11755 n11766_not ; n11767
g11704 and n11180 n11698 ; n11768
g11705 nor n11699 n11768 ; n11769
g11706 and n3964_not n11727 ; n11770
g11707 and n3456_not n11055 ; n11771
g11708 and n3805_not n11715 ; n11772
g11709 nor n11771 n11772 ; n11773
g11710 and n11770_not n11773 ; n11774
g11711 and n11057_not n11774 ; n11775
g11712 and n4558_not n11774 ; n11776
g11713 nor n11775 n11776 ; n11777
g11714 and a[2] n11777_not ; n11778
g11715 and a[2]_not n11777 ; n11779
g11716 nor n11778 n11779 ; n11780
g11717 and n11769 n11780_not ; n11781
g11718 and n11692 n11694_not ; n11782
g11719 nor n11695 n11782 ; n11783
g11720 and n11677 n11679_not ; n11784
g11721 nor n11680 n11784 ; n11785
g11722 and n11657 n11659_not ; n11786
g11723 nor n11660 n11786 ; n11787
g11724 and n11637 n11639_not ; n11788
g11725 nor n11640 n11788 ; n11789
g11726 and n11615 n11617_not ; n11790
g11727 nor n11618 n11790 ; n11791
g11728 and n11586_not n11597 ; n11792
g11729 nor n11598 n11792 ; n11793
g11730 nor n11057 n11727 ; n11794
g11731 nor n2829 n11794 ; n11795
g11732 and a[2] n11057 ; n11796
g11733 and n6798 n11796 ; n11797
g11734 and n2674_not n11727 ; n11798
g11735 and n2829_not n11055 ; n11799
g11736 and n2736_not n11715 ; n11800
g11737 nor n11799 n11800 ; n11801
g11738 and n11798_not n11801 ; n11802
g11739 and a[2] n11802_not ; n11803
g11740 and n7469_not n11796 ; n11804
g11741 and a[2] n11715 ; n11805
g11742 and n2829_not n11805 ; n11806
g11743 and a[2] n11727 ; n11807
g11744 and n2736_not n11807 ; n11808
g11745 and a[2] n11808_not ; n11809
g11746 and n11806_not n11809 ; n11810
g11747 and n11804_not n11810 ; n11811
g11748 and n11803_not n11811 ; n11812
g11749 and n11797_not n11812 ; n11813
g11750 and n11795_not n11813 ; n11814
g11751 and n11584 n11814 ; n11815
g11752 nor n11584 n11814 ; n11816
g11753 and n2571_not n11727 ; n11817
g11754 and n2736_not n11055 ; n11818
g11755 and n2674_not n11715 ; n11819
g11756 nor n11818 n11819 ; n11820
g11757 and n11817_not n11820 ; n11821
g11758 and n6806 n11057 ; n11822
g11759 and n11821 n11822_not ; n11823
g11760 nor a[2] n11823 ; n11824
g11761 and a[2] n11823 ; n11825
g11762 nor n11824 n11825 ; n11826
g11763 nor n11816 n11826 ; n11827
g11764 nor n11815 n11827 ; n11828
g11765 and n2533_not n11727 ; n11829
g11766 and n2674_not n11055 ; n11830
g11767 and n2571_not n11715 ; n11831
g11768 nor n11830 n11831 ; n11832
g11769 and n11829_not n11832 ; n11833
g11770 and n11057_not n11833 ; n11834
g11771 and n6695_not n11833 ; n11835
g11772 nor n11834 n11835 ; n11836
g11773 and a[2] n11836_not ; n11837
g11774 and a[2]_not n11836 ; n11838
g11775 nor n11837 n11838 ; n11839
g11776 and n11828 n11839 ; n11840
g11777 and n11583 n11585_not ; n11841
g11778 nor n11586 n11841 ; n11842
g11779 and n11840_not n11842 ; n11843
g11780 nor n11828 n11839 ; n11844
g11781 nor n11843 n11844 ; n11845
g11782 and n11793 n11845_not ; n11846
g11783 and n11793_not n11845 ; n11847
g11784 and n2464_not n11727 ; n11848
g11785 and n2571_not n11055 ; n11849
g11786 and n2533_not n11715 ; n11850
g11787 nor n11849 n11850 ; n11851
g11788 and n11848_not n11851 ; n11852
g11789 and n6646 n11057 ; n11853
g11790 and n11852 n11853_not ; n11854
g11791 nor a[2] n11854 ; n11855
g11792 and a[2] n11854 ; n11856
g11793 nor n11855 n11856 ; n11857
g11794 nor n11847 n11857 ; n11858
g11795 nor n11846 n11858 ; n11859
g11796 and n2388_not n11727 ; n11860
g11797 and n2533_not n11055 ; n11861
g11798 and n2464_not n11715 ; n11862
g11799 nor n11861 n11862 ; n11863
g11800 and n11860_not n11863 ; n11864
g11801 and n11057_not n11864 ; n11865
g11802 and n6591_not n11864 ; n11866
g11803 nor n11865 n11866 ; n11867
g11804 and a[2] n11867_not ; n11868
g11805 and a[2]_not n11867 ; n11869
g11806 nor n11868 n11869 ; n11870
g11807 nor n11859 n11870 ; n11871
g11808 and n11859 n11870 ; n11872
g11809 and n11602 n11613 ; n11873
g11810 nor n11614 n11873 ; n11874
g11811 and n11872_not n11874 ; n11875
g11812 nor n11871 n11875 ; n11876
g11813 and n11791 n11876_not ; n11877
g11814 and n11791_not n11876 ; n11878
g11815 and n2291_not n11727 ; n11879
g11816 and n2464_not n11055 ; n11880
g11817 and n2388_not n11715 ; n11881
g11818 nor n11880 n11881 ; n11882
g11819 and n11879_not n11882 ; n11883
g11820 and n6541 n11057 ; n11884
g11821 and n11883 n11884_not ; n11885
g11822 nor a[2] n11885 ; n11886
g11823 and a[2] n11885 ; n11887
g11824 nor n11886 n11887 ; n11888
g11825 nor n11878 n11888 ; n11889
g11826 nor n11877 n11889 ; n11890
g11827 and n2189_not n11727 ; n11891
g11828 and n2388_not n11055 ; n11892
g11829 and n2291_not n11715 ; n11893
g11830 nor n11892 n11893 ; n11894
g11831 and n11891_not n11894 ; n11895
g11832 and n11057_not n11895 ; n11896
g11833 and n6122_not n11895 ; n11897
g11834 nor n11896 n11897 ; n11898
g11835 and a[2] n11898_not ; n11899
g11836 and a[2]_not n11898 ; n11900
g11837 nor n11899 n11900 ; n11901
g11838 and n11890 n11901 ; n11902
g11839 and n11560 n11619 ; n11903
g11840 nor n11620 n11903 ; n11904
g11841 and n11902_not n11904 ; n11905
g11842 nor n11890 n11901 ; n11906
g11843 nor n11905 n11906 ; n11907
g11844 and n2152_not n11727 ; n11908
g11845 and n2291_not n11055 ; n11909
g11846 and n2189_not n11715 ; n11910
g11847 nor n11909 n11910 ; n11911
g11848 and n11908_not n11911 ; n11912
g11849 and n11057_not n11912 ; n11913
g11850 and n6492_not n11912 ; n11914
g11851 nor n11913 n11914 ; n11915
g11852 and a[2] n11915_not ; n11916
g11853 and a[2]_not n11915 ; n11917
g11854 nor n11916 n11917 ; n11918
g11855 and n11907 n11918 ; n11919
g11856 and n11621 n11623_not ; n11920
g11857 nor n11624 n11920 ; n11921
g11858 and n11919_not n11921 ; n11922
g11859 nor n11907 n11918 ; n11923
g11860 nor n11922 n11923 ; n11924
g11861 and n2057_not n11727 ; n11925
g11862 and n2189_not n11055 ; n11926
g11863 and n2152_not n11715 ; n11927
g11864 nor n11926 n11927 ; n11928
g11865 and n11925_not n11928 ; n11929
g11866 and n11057_not n11929 ; n11930
g11867 and n6479_not n11929 ; n11931
g11868 nor n11930 n11931 ; n11932
g11869 and a[2] n11932_not ; n11933
g11870 and a[2]_not n11932 ; n11934
g11871 nor n11933 n11934 ; n11935
g11872 and n11924 n11935 ; n11936
g11873 and n11528 n11625 ; n11937
g11874 nor n11626 n11937 ; n11938
g11875 and n11936_not n11938 ; n11939
g11876 nor n11924 n11935 ; n11940
g11877 nor n11939 n11940 ; n11941
g11878 and n11627 n11629_not ; n11942
g11879 and n11628_not n11942 ; n11943
g11880 nor n11631 n11943 ; n11944
g11881 and n11941_not n11944 ; n11945
g11882 and n11941 n11944_not ; n11946
g11883 and n1992_not n11727 ; n11947
g11884 and n2152_not n11055 ; n11948
g11885 and n2057_not n11715 ; n11949
g11886 nor n11948 n11949 ; n11950
g11887 and n11947_not n11950 ; n11951
g11888 and n6143 n11057 ; n11952
g11889 and n11951 n11952_not ; n11953
g11890 nor a[2] n11953 ; n11954
g11891 and a[2] n11953 ; n11955
g11892 nor n11954 n11955 ; n11956
g11893 nor n11946 n11956 ; n11957
g11894 nor n11945 n11957 ; n11958
g11895 and n11632 n11634_not ; n11959
g11896 and n11633_not n11959 ; n11960
g11897 nor n11636 n11960 ; n11961
g11898 and n11958_not n11961 ; n11962
g11899 and n11958 n11961_not ; n11963
g11900 and n1913_not n11727 ; n11964
g11901 and n2057_not n11055 ; n11965
g11902 and n1992_not n11715 ; n11966
g11903 nor n11965 n11966 ; n11967
g11904 and n11964_not n11967 ; n11968
g11905 and n5834 n11057 ; n11969
g11906 and n11968 n11969_not ; n11970
g11907 nor a[2] n11970 ; n11971
g11908 and a[2] n11970 ; n11972
g11909 nor n11971 n11972 ; n11973
g11910 nor n11963 n11973 ; n11974
g11911 nor n11962 n11974 ; n11975
g11912 and n11789 n11975_not ; n11976
g11913 and n11789_not n11975 ; n11977
g11914 and n1877_not n11727 ; n11978
g11915 and n1992_not n11055 ; n11979
g11916 and n1913_not n11715 ; n11980
g11917 nor n11979 n11980 ; n11981
g11918 and n11978_not n11981 ; n11982
g11919 and n6007 n11057 ; n11983
g11920 and n11982 n11983_not ; n11984
g11921 nor a[2] n11984 ; n11985
g11922 and a[2] n11984 ; n11986
g11923 nor n11985 n11986 ; n11987
g11924 nor n11977 n11987 ; n11988
g11925 nor n11976 n11988 ; n11989
g11926 and n1779_not n11727 ; n11990
g11927 and n1913_not n11055 ; n11991
g11928 and n1877_not n11715 ; n11992
g11929 nor n11991 n11992 ; n11993
g11930 and n11990_not n11993 ; n11994
g11931 and n11057_not n11994 ; n11995
g11932 and n5851_not n11994 ; n11996
g11933 nor n11995 n11996 ; n11997
g11934 and a[2] n11997_not ; n11998
g11935 and a[2]_not n11997 ; n11999
g11936 nor n11998 n11999 ; n12000
g11937 and n11989 n12000 ; n12001
g11938 and n11469 n11641 ; n12002
g11939 nor n11642 n12002 ; n12003
g11940 and n12001_not n12003 ; n12004
g11941 nor n11989 n12000 ; n12005
g11942 nor n12004 n12005 ; n12006
g11943 and n1665_not n11727 ; n12007
g11944 and n1877_not n11055 ; n12008
g11945 and n1779_not n11715 ; n12009
g11946 nor n12008 n12009 ; n12010
g11947 and n12007_not n12010 ; n12011
g11948 and n11057_not n12011 ; n12012
g11949 and n5328_not n12011 ; n12013
g11950 nor n12012 n12013 ; n12014
g11951 and a[2] n12014_not ; n12015
g11952 and a[2]_not n12014 ; n12016
g11953 nor n12015 n12016 ; n12017
g11954 and n12006 n12017 ; n12018
g11955 and n11451 n11643 ; n12019
g11956 nor n11644 n12019 ; n12020
g11957 and n12018_not n12020 ; n12021
g11958 nor n12006 n12017 ; n12022
g11959 nor n12021 n12022 ; n12023
g11960 and n1572_not n11727 ; n12024
g11961 and n1779_not n11055 ; n12025
g11962 and n1665_not n11715 ; n12026
g11963 nor n12025 n12026 ; n12027
g11964 and n12024_not n12027 ; n12028
g11965 and n11057_not n12028 ; n12029
g11966 and n5561_not n12028 ; n12030
g11967 nor n12029 n12030 ; n12031
g11968 and a[2] n12031_not ; n12032
g11969 and a[2]_not n12031 ; n12033
g11970 nor n12032 n12033 ; n12034
g11971 and n12023 n12034 ; n12035
g11972 and n11433 n11645 ; n12036
g11973 nor n11646 n12036 ; n12037
g11974 and n12035_not n12037 ; n12038
g11975 nor n12023 n12034 ; n12039
g11976 nor n12038 n12039 ; n12040
g11977 and n11647 n11649_not ; n12041
g11978 and n11648_not n12041 ; n12042
g11979 nor n11651 n12042 ; n12043
g11980 and n12040_not n12043 ; n12044
g11981 and n12040 n12043_not ; n12045
g11982 and n1472_not n11727 ; n12046
g11983 and n1665_not n11055 ; n12047
g11984 and n1572_not n11715 ; n12048
g11985 nor n12047 n12048 ; n12049
g11986 and n12046_not n12049 ; n12050
g11987 and n5139 n11057 ; n12051
g11988 and n12050 n12051_not ; n12052
g11989 nor a[2] n12052 ; n12053
g11990 and a[2] n12052 ; n12054
g11991 nor n12053 n12054 ; n12055
g11992 nor n12045 n12055 ; n12056
g11993 nor n12044 n12056 ; n12057
g11994 and n11652 n11654_not ; n12058
g11995 and n11653_not n12058 ; n12059
g11996 nor n11656 n12059 ; n12060
g11997 and n12057_not n12060 ; n12061
g11998 and n12057 n12060_not ; n12062
g11999 and n1364_not n11727 ; n12063
g12000 and n1572_not n11055 ; n12064
g12001 and n1472_not n11715 ; n12065
g12002 nor n12064 n12065 ; n12066
g12003 and n12063_not n12066 ; n12067
g12004 and n5114 n11057 ; n12068
g12005 and n12067 n12068_not ; n12069
g12006 nor a[2] n12069 ; n12070
g12007 and a[2] n12069 ; n12071
g12008 nor n12070 n12071 ; n12072
g12009 nor n12062 n12072 ; n12073
g12010 nor n12061 n12073 ; n12074
g12011 and n11787 n12074_not ; n12075
g12012 and n11787_not n12074 ; n12076
g12013 and n1235_not n11727 ; n12077
g12014 and n1472_not n11055 ; n12078
g12015 and n1364_not n11715 ; n12079
g12016 nor n12078 n12079 ; n12080
g12017 and n12077_not n12080 ; n12081
g12018 and n4848 n11057 ; n12082
g12019 and n12081 n12082_not ; n12083
g12020 nor a[2] n12083 ; n12084
g12021 and a[2] n12083 ; n12085
g12022 nor n12084 n12085 ; n12086
g12023 nor n12076 n12086 ; n12087
g12024 nor n12075 n12087 ; n12088
g12025 and n1178_not n11727 ; n12089
g12026 and n1364_not n11055 ; n12090
g12027 and n1235_not n11715 ; n12091
g12028 nor n12090 n12091 ; n12092
g12029 and n12089_not n12092 ; n12093
g12030 and n11057_not n12093 ; n12094
g12031 and n4861_not n12093 ; n12095
g12032 nor n12094 n12095 ; n12096
g12033 and a[2] n12096_not ; n12097
g12034 and a[2]_not n12096 ; n12098
g12035 nor n12097 n12098 ; n12099
g12036 and n12088 n12099 ; n12100
g12037 and n11374 n11661 ; n12101
g12038 nor n11662 n12101 ; n12102
g12039 and n12100_not n12102 ; n12103
g12040 nor n12088 n12099 ; n12104
g12041 nor n12103 n12104 ; n12105
g12042 and n1060_not n11727 ; n12106
g12043 and n1235_not n11055 ; n12107
g12044 and n1178_not n11715 ; n12108
g12045 nor n12107 n12108 ; n12109
g12046 and n12106_not n12109 ; n12110
g12047 and n11057_not n12110 ; n12111
g12048 and n4429_not n12110 ; n12112
g12049 nor n12111 n12112 ; n12113
g12050 and a[2] n12113_not ; n12114
g12051 and a[2]_not n12113 ; n12115
g12052 nor n12114 n12115 ; n12116
g12053 and n12105 n12116 ; n12117
g12054 and n11356 n11663 ; n12118
g12055 nor n11664 n12118 ; n12119
g12056 and n12117_not n12119 ; n12120
g12057 nor n12105 n12116 ; n12121
g12058 nor n12120 n12121 ; n12122
g12059 and n958_not n11727 ; n12123
g12060 and n1178_not n11055 ; n12124
g12061 and n1060_not n11715 ; n12125
g12062 nor n12124 n12125 ; n12126
g12063 and n12123_not n12126 ; n12127
g12064 and n11057_not n12127 ; n12128
g12065 and n4633_not n12127 ; n12129
g12066 nor n12128 n12129 ; n12130
g12067 and a[2] n12130_not ; n12131
g12068 and a[2]_not n12130 ; n12132
g12069 nor n12131 n12132 ; n12133
g12070 and n12122 n12133 ; n12134
g12071 and n11338 n11665 ; n12135
g12072 nor n11666 n12135 ; n12136
g12073 and n12134_not n12136 ; n12137
g12074 nor n12122 n12133 ; n12138
g12075 nor n12137 n12138 ; n12139
g12076 and n11667 n11669_not ; n12140
g12077 and n11668_not n12140 ; n12141
g12078 nor n11671 n12141 ; n12142
g12079 and n12139_not n12142 ; n12143
g12080 and n12139 n12142_not ; n12144
g12081 and n867_not n11727 ; n12145
g12082 and n1060_not n11055 ; n12146
g12083 and n958_not n11715 ; n12147
g12084 nor n12146 n12147 ; n12148
g12085 and n12145_not n12148 ; n12149
g12086 and n4204 n11057 ; n12150
g12087 and n12149 n12150_not ; n12151
g12088 nor a[2] n12151 ; n12152
g12089 and a[2] n12151 ; n12153
g12090 nor n12152 n12153 ; n12154
g12091 nor n12144 n12154 ; n12155
g12092 nor n12143 n12155 ; n12156
g12093 and n11672 n11674_not ; n12157
g12094 and n11673_not n12157 ; n12158
g12095 nor n11676 n12158 ; n12159
g12096 and n12156_not n12159 ; n12160
g12097 and n12156 n12159_not ; n12161
g12098 and n710_not n11727 ; n12162
g12099 and n958_not n11055 ; n12163
g12100 and n867_not n11715 ; n12164
g12101 nor n12163 n12164 ; n12165
g12102 and n12162_not n12165 ; n12166
g12103 and n4179 n11057 ; n12167
g12104 and n12166 n12167_not ; n12168
g12105 nor a[2] n12168 ; n12169
g12106 and a[2] n12168 ; n12170
g12107 nor n12169 n12170 ; n12171
g12108 nor n12161 n12171 ; n12172
g12109 nor n12160 n12172 ; n12173
g12110 and n11785 n12173_not ; n12174
g12111 and n11785_not n12173 ; n12175
g12112 and n587_not n11727 ; n12176
g12113 and n867_not n11055 ; n12177
g12114 and n710_not n11715 ; n12178
g12115 nor n12177 n12178 ; n12179
g12116 and n12176_not n12179 ; n12180
g12117 and n3331 n11057 ; n12181
g12118 and n12180 n12181_not ; n12182
g12119 nor a[2] n12182 ; n12183
g12120 and a[2] n12182 ; n12184
g12121 nor n12183 n12184 ; n12185
g12122 nor n12175 n12185 ; n12186
g12123 nor n12174 n12186 ; n12187
g12124 and n392_not n11727 ; n12188
g12125 and n710_not n11055 ; n12189
g12126 and n587_not n11715 ; n12190
g12127 nor n12189 n12190 ; n12191
g12128 and n12188_not n12191 ; n12192
g12129 and n11057_not n12192 ; n12193
g12130 and n3347_not n12192 ; n12194
g12131 nor n12193 n12194 ; n12195
g12132 and a[2] n12195_not ; n12196
g12133 and a[2]_not n12195 ; n12197
g12134 nor n12196 n12197 ; n12198
g12135 and n12187 n12198 ; n12199
g12136 and n11279 n11681 ; n12200
g12137 nor n11682 n12200 ; n12201
g12138 and n12199_not n12201 ; n12202
g12139 nor n12187 n12198 ; n12203
g12140 nor n12202 n12203 ; n12204
g12141 and n3012_not n11727 ; n12205
g12142 and n587_not n11055 ; n12206
g12143 and n392_not n11715 ; n12207
g12144 nor n12206 n12207 ; n12208
g12145 and n12205_not n12208 ; n12209
g12146 and n11057_not n12209 ; n12210
g12147 and n3018_not n12209 ; n12211
g12148 nor n12210 n12211 ; n12212
g12149 and a[2] n12212_not ; n12213
g12150 and a[2]_not n12212 ; n12214
g12151 nor n12213 n12214 ; n12215
g12152 and n12204 n12215 ; n12216
g12153 and n11261 n11683 ; n12217
g12154 nor n11684 n12217 ; n12218
g12155 and n12216_not n12218 ; n12219
g12156 nor n12204 n12215 ; n12220
g12157 nor n12219 n12220 ; n12221
g12158 and n3539_not n11727 ; n12222
g12159 and n392_not n11055 ; n12223
g12160 and n3012_not n11715 ; n12224
g12161 nor n12223 n12224 ; n12225
g12162 and n12222_not n12225 ; n12226
g12163 and n11057_not n12226 ; n12227
g12164 and n3715_not n12226 ; n12228
g12165 nor n12227 n12228 ; n12229
g12166 and a[2] n12229_not ; n12230
g12167 and a[2]_not n12229 ; n12231
g12168 nor n12230 n12231 ; n12232
g12169 and n12221 n12232 ; n12233
g12170 and n11243 n11685 ; n12234
g12171 nor n11686 n12234 ; n12235
g12172 and n12233_not n12235 ; n12236
g12173 nor n12221 n12232 ; n12237
g12174 nor n12236 n12237 ; n12238
g12175 and n11687 n11689_not ; n12239
g12176 and n11688_not n12239 ; n12240
g12177 nor n11691 n12240 ; n12241
g12178 and n12238_not n12241 ; n12242
g12179 and n12238 n12241_not ; n12243
g12180 and n3605_not n11727 ; n12244
g12181 and n3012_not n11055 ; n12245
g12182 and n3539_not n11715 ; n12246
g12183 nor n12245 n12246 ; n12247
g12184 and n12244_not n12247 ; n12248
g12185 and n4084 n11057 ; n12249
g12186 and n12248 n12249_not ; n12250
g12187 nor a[2] n12250 ; n12251
g12188 and a[2] n12250 ; n12252
g12189 nor n12251 n12252 ; n12253
g12190 nor n12243 n12253 ; n12254
g12191 nor n12242 n12254 ; n12255
g12192 and n11783 n12255_not ; n12256
g12193 and n11783_not n12255 ; n12257
g12194 and n3456_not n11727 ; n12258
g12195 and n3539_not n11055 ; n12259
g12196 and n3605_not n11715 ; n12260
g12197 nor n12259 n12260 ; n12261
g12198 and n12258_not n12261 ; n12262
g12199 and n3627 n11057 ; n12263
g12200 and n12262 n12263_not ; n12264
g12201 nor a[2] n12264 ; n12265
g12202 and a[2] n12264 ; n12266
g12203 nor n12265 n12266 ; n12267
g12204 nor n12257 n12267 ; n12268
g12205 nor n12256 n12268 ; n12269
g12206 and n3805_not n11727 ; n12270
g12207 and n3605_not n11055 ; n12271
g12208 and n3456_not n11715 ; n12272
g12209 nor n12271 n12272 ; n12273
g12210 and n12270_not n12273 ; n12274
g12211 and n11057_not n12274 ; n12275
g12212 and n3818_not n12274 ; n12276
g12213 nor n12275 n12276 ; n12277
g12214 and a[2] n12277_not ; n12278
g12215 and a[2]_not n12277 ; n12279
g12216 nor n12278 n12279 ; n12280
g12217 and n12269 n12280 ; n12281
g12218 and n11198 n11696 ; n12282
g12219 nor n11697 n12282 ; n12283
g12220 and n12281_not n12283 ; n12284
g12221 nor n12269 n12280 ; n12285
g12222 nor n12284 n12285 ; n12286
g12223 and n11769 n11781_not ; n12287
g12224 nor n11780 n11781 ; n12288
g12225 nor n12287 n12288 ; n12289
g12226 nor n12286 n12289 ; n12290
g12227 nor n11781 n12290 ; n12291
g12228 and n11755_not n11766 ; n12292
g12229 nor n11767 n12292 ; n12293
g12230 and n12291_not n12293 ; n12294
g12231 nor n11767 n12294 ; n12295
g12232 and n11741_not n11752 ; n12296
g12233 nor n11753 n12296 ; n12297
g12234 and n12295_not n12297 ; n12298
g12235 nor n11753 n12298 ; n12299
g12236 and n11726_not n11738 ; n12300
g12237 nor n11739 n12300 ; n12301
g12238 and n12299_not n12301 ; n12302
g12239 nor n11739 n12302 ; n12303
g12240 and n11713_not n11723 ; n12304
g12241 nor n11724 n12304 ; n12305
g12242 and n12303_not n12305 ; n12306
g12243 nor n11724 n12306 ; n12307
g12244 and n11711 n12307_not ; n12308
g12245 nor n11709 n12308 ; n12309
g12246 and n11083 n11086_not ; n12310
g12247 nor n11087 n12310 ; n12311
g12248 and n12309_not n12311 ; n12312
g12249 nor n11087 n12312 ; n12313
g12250 and n11047 n11049_not ; n12314
g12251 nor n11050 n12314 ; n12315
g12252 and n12313_not n12315 ; n12316
g12253 nor n11050 n12316 ; n12317
g12254 and n10453 n12317_not ; n12318
g12255 nor n10451 n12318 ; n12319
g12256 and n9883 n9886_not ; n12320
g12257 nor n9887 n12320 ; n12321
g12258 and n12319_not n12321 ; n12322
g12259 nor n9887 n12322 ; n12323
g12260 and n9363 n9365_not ; n12324
g12261 nor n9366 n12324 ; n12325
g12262 and n12323_not n12325 ; n12326
g12263 nor n9366 n12326 ; n12327
g12264 and n8879 n12327_not ; n12328
g12265 nor n8877 n12328 ; n12329
g12266 and n8437 n12329_not ; n12330
g12267 nor n8435 n12330 ; n12331
g12268 and n8015 n8017_not ; n12332
g12269 nor n8018 n12332 ; n12333
g12270 and n12331_not n12333 ; n12334
g12271 nor n8018 n12334 ; n12335
g12272 and n7651 n12335_not ; n12336
g12273 nor n7649 n12336 ; n12337
g12274 and n7307 n7310_not ; n12338
g12275 nor n7311 n12338 ; n12339
g12276 and n12337_not n12339 ; n12340
g12277 nor n7311 n12340 ; n12341
g12278 and n7133 n7135_not ; n12342
g12279 nor n7136 n12342 ; n12343
g12280 and n12341_not n12343 ; n12344
g12281 nor n7136 n12344 ; n12345
g12282 and n6970 n12345_not ; n12346
g12283 nor n6968 n12346 ; n12347
g12284 and n6422 n12347_not ; n12348
g12285 nor n6420 n12348 ; n12349
g12286 and n6267 n12349_not ; n12350
g12287 nor n6265 n12350 ; n12351
g12288 and n5952 n12351_not ; n12352
g12289 nor n5950 n12352 ; n12353
g12290 and n5679 n5681_not ; n12354
g12291 nor n5682 n12354 ; n12355
g12292 and n12353_not n12355 ; n12356
g12293 nor n5682 n12356 ; n12357
g12294 and n5530 n12357_not ; n12358
g12295 nor n5528 n12358 ; n12359
g12296 and n5420 n12359_not ; n12360
g12297 nor n5418 n12360 ; n12361
g12298 and n4954 n12361_not ; n12362
g12299 nor n4952 n12362 ; n12363
g12300 and n4728 n4730_not ; n12364
g12301 nor n4731 n12364 ; n12365
g12302 and n12363_not n12365 ; n12366
g12303 nor n4731 n12366 ; n12367
g12304 and n4622 n12367_not ; n12368
g12305 and n4622_not n12367 ; n12369
g12306 nor n12368 n12369 ; n12370
g12307 nor n4621 n12368 ; n12371
g12308 nor n4542 n4545 ; n12372
g12309 and n3457 n3964_not ; n12373
g12310 and n3456_not n3542 ; n12374
g12311 and n3606 n3805_not ; n12375
g12312 nor n12374 n12375 ; n12376
g12313 and n12373_not n12376 ; n12377
g12314 and n3368 n4558 ; n12378
g12315 and n12377 n12378_not ; n12379
g12316 and a[29] n12379_not ; n12380
g12317 and a[29] n12380_not ; n12381
g12318 nor n12379 n12380 ; n12382
g12319 nor n12381 n12382 ; n12383
g12320 nor n3720 n3724 ; n12384
g12321 and n288 n2276 ; n12385
g12322 and n123_not n12385 ; n12386
g12323 and n231_not n12386 ; n12387
g12324 and n495_not n508 ; n12388
g12325 and n367_not n12388 ; n12389
g12326 and n205_not n12389 ; n12390
g12327 and n2584 n12390 ; n12391
g12328 and n12387 n12391 ; n12392
g12329 and n2582 n12392 ; n12393
g12330 and n171_not n12393 ; n12394
g12331 and n121_not n12394 ; n12395
g12332 and n163_not n12395 ; n12396
g12333 nor n400 n1203 ; n12397
g12334 and n1550 n12397 ; n12398
g12335 and n111_not n12398 ; n12399
g12336 and n289_not n12399 ; n12400
g12337 and n426_not n12400 ; n12401
g12338 and n932_not n12401 ; n12402
g12339 and n470_not n12402 ; n12403
g12340 and n271_not n12403 ; n12404
g12341 and n533 n1071 ; n12405
g12342 and n194_not n12405 ; n12406
g12343 and n203_not n12406 ; n12407
g12344 and n147_not n12407 ; n12408
g12345 and n403_not n12408 ; n12409
g12346 and n290_not n2346 ; n12410
g12347 and n452_not n12410 ; n12411
g12348 and n306_not n12411 ; n12412
g12349 and n1644 n12412 ; n12413
g12350 and n12409 n12413 ; n12414
g12351 and n1496 n12414 ; n12415
g12352 and n2961 n12415 ; n12416
g12353 and n811 n12416 ; n12417
g12354 and n774 n12417 ; n12418
g12355 and n1253 n12418 ; n12419
g12356 and n1994 n12419 ; n12420
g12357 and n885 n12420 ; n12421
g12358 and n276_not n12421 ; n12422
g12359 and n847_not n12422 ; n12423
g12360 and n355_not n12423 ; n12424
g12361 and n91_not n12424 ; n12425
g12362 and n424_not n12425 ; n12426
g12363 and n451_not n12426 ; n12427
g12364 and n81_not n12427 ; n12428
g12365 nor n142 n301 ; n12429
g12366 and n564_not n12429 ; n12430
g12367 and n633_not n12430 ; n12431
g12368 and n253 n722 ; n12432
g12369 and n1158 n12432 ; n12433
g12370 and n12431 n12433 ; n12434
g12371 and n12428 n12434 ; n12435
g12372 and n12404 n12435 ; n12436
g12373 and n6769 n12436 ; n12437
g12374 and n12396 n12437 ; n12438
g12375 and n3163 n12438 ; n12439
g12376 and n1306_not n12439 ; n12440
g12377 and n232_not n12440 ; n12441
g12378 and n571_not n12441 ; n12442
g12379 and n656_not n12442 ; n12443
g12380 and n357_not n12443 ; n12444
g12381 and n371_not n12444 ; n12445
g12382 and n119_not n12445 ; n12446
g12383 and n569_not n12446 ; n12447
g12384 and n429_not n12447 ; n12448
g12385 nor n3702 n12448 ; n12449
g12386 and n3702 n12448 ; n12450
g12387 nor n12449 n12450 ; n12451
g12388 and a[23]_not n12451 ; n12452
g12389 nor a[23] n12452 ; n12453
g12390 nor n12449 n12452 ; n12454
g12391 and n12450_not n12454 ; n12455
g12392 nor n12453 n12455 ; n12456
g12393 and n3020 n3605_not ; n12457
g12394 and n3028 n3539_not ; n12458
g12395 and n3012_not n3023 ; n12459
g12396 and n75 n4084 ; n12460
g12397 nor n12459 n12460 ; n12461
g12398 and n12458_not n12461 ; n12462
g12399 and n12457_not n12462 ; n12463
g12400 nor n12456 n12463 ; n12464
g12401 and n12456 n12463 ; n12465
g12402 nor n12464 n12465 ; n12466
g12403 and n3708_not n12466 ; n12467
g12404 and n3708 n12466_not ; n12468
g12405 nor n12467 n12468 ; n12469
g12406 and n12384_not n12469 ; n12470
g12407 and n12384 n12469_not ; n12471
g12408 nor n12470 n12471 ; n12472
g12409 and n12383_not n12472 ; n12473
g12410 and n12472 n12473_not ; n12474
g12411 nor n12383 n12473 ; n12475
g12412 nor n12474 n12475 ; n12476
g12413 nor n3825 n4074 ; n12477
g12414 and n3884 n4515_not ; n12478
g12415 and n3967 n4045_not ; n12479
g12416 and n3877_not n4046 ; n12480
g12417 nor n12479 n12480 ; n12481
g12418 and n12478_not n12481 ; n12482
g12419 and n4050_not n12482 ; n12483
g12420 and n4715_not n12482 ; n12484
g12421 nor n12483 n12484 ; n12485
g12422 and a[26] n12485_not ; n12486
g12423 and a[26]_not n12485 ; n12487
g12424 nor n12486 n12487 ; n12488
g12425 nor n12477 n12488 ; n12489
g12426 nor n12477 n12489 ; n12490
g12427 nor n12488 n12489 ; n12491
g12428 nor n12490 n12491 ; n12492
g12429 nor n12476 n12492 ; n12493
g12430 and n12476 n12491_not ; n12494
g12431 and n12490_not n12494 ; n12495
g12432 nor n12493 n12495 ; n12496
g12433 and n12372_not n12496 ; n12497
g12434 and n12372 n12496_not ; n12498
g12435 nor n12497 n12498 ; n12499
g12436 and n12371_not n12499 ; n12500
g12437 and n12371 n12499_not ; n12501
g12438 nor n12500 n12501 ; n12502
g12439 and n12370 n12502 ; n12503
g12440 and n12363 n12365_not ; n12504
g12441 nor n12366 n12504 ; n12505
g12442 and n12370 n12505 ; n12506
g12443 and n4954_not n12361 ; n12507
g12444 nor n12362 n12507 ; n12508
g12445 and n12505 n12508 ; n12509
g12446 and n5530_not n12357 ; n12510
g12447 nor n12358 n12510 ; n12511
g12448 and n5420_not n12359 ; n12512
g12449 nor n12360 n12512 ; n12513
g12450 and n12511 n12513 ; n12514
g12451 and n12353 n12355_not ; n12515
g12452 nor n12356 n12515 ; n12516
g12453 and n12511 n12516 ; n12517
g12454 and n5952_not n12351 ; n12518
g12455 nor n12352 n12518 ; n12519
g12456 and n12516 n12519 ; n12520
g12457 and n6267_not n12349 ; n12521
g12458 nor n12350 n12521 ; n12522
g12459 and n12519 n12522 ; n12523
g12460 and n6422_not n12347 ; n12524
g12461 nor n12348 n12524 ; n12525
g12462 and n12522 n12525 ; n12526
g12463 and n6970_not n12345 ; n12527
g12464 nor n12346 n12527 ; n12528
g12465 and n12525 n12528 ; n12529
g12466 and n12341 n12343_not ; n12530
g12467 nor n12344 n12530 ; n12531
g12468 and n12528 n12531 ; n12532
g12469 and n12337 n12339_not ; n12533
g12470 nor n12340 n12533 ; n12534
g12471 and n12531 n12534 ; n12535
g12472 and n7651_not n12335 ; n12536
g12473 nor n12336 n12536 ; n12537
g12474 and n12534 n12537 ; n12538
g12475 and n12331 n12333_not ; n12539
g12476 nor n12334 n12539 ; n12540
g12477 and n12537 n12540 ; n12541
g12478 and n8437_not n12329 ; n12542
g12479 nor n12330 n12542 ; n12543
g12480 and n12540 n12543 ; n12544
g12481 and n8879_not n12327 ; n12545
g12482 nor n12328 n12545 ; n12546
g12483 and n12543 n12546 ; n12547
g12484 and n12323 n12325_not ; n12548
g12485 nor n12326 n12548 ; n12549
g12486 and n12546 n12549 ; n12550
g12487 and n12319 n12321_not ; n12551
g12488 nor n12322 n12551 ; n12552
g12489 and n12549 n12552 ; n12553
g12490 and n10453_not n12317 ; n12554
g12491 nor n12318 n12554 ; n12555
g12492 and n12552 n12555 ; n12556
g12493 and n12313 n12315_not ; n12557
g12494 nor n12316 n12557 ; n12558
g12495 and n12555 n12558 ; n12559
g12496 and n12309 n12311_not ; n12560
g12497 nor n12312 n12560 ; n12561
g12498 and n12558 n12561 ; n12562
g12499 and n11711_not n12307 ; n12563
g12500 nor n12308 n12563 ; n12564
g12501 and n12561 n12564 ; n12565
g12502 and n12303 n12305_not ; n12566
g12503 nor n12306 n12566 ; n12567
g12504 and n12564 n12567 ; n12568
g12505 nor n12564 n12567 ; n12569
g12506 and n12299 n12301_not ; n12570
g12507 nor n12302 n12570 ; n12571
g12508 and n12567 n12571 ; n12572
g12509 and n12295 n12297_not ; n12573
g12510 nor n12298 n12573 ; n12574
g12511 and n12571 n12574 ; n12575
g12512 and n12291 n12293_not ; n12576
g12513 nor n12294 n12576 ; n12577
g12514 and n12574 n12577 ; n12578
g12515 nor n12286 n12290 ; n12579
g12516 nor n12289 n12290 ; n12580
g12517 nor n12579 n12580 ; n12581
g12518 and n12577 n12581_not ; n12582
g12519 and n12574_not n12582 ; n12583
g12520 nor n12578 n12583 ; n12584
g12521 nor n12571 n12574 ; n12585
g12522 nor n12575 n12585 ; n12586
g12523 and n12584_not n12586 ; n12587
g12524 nor n12575 n12587 ; n12588
g12525 nor n12567 n12571 ; n12589
g12526 nor n12572 n12589 ; n12590
g12527 and n12588_not n12590 ; n12591
g12528 nor n12572 n12591 ; n12592
g12529 nor n12568 n12592 ; n12593
g12530 and n12569_not n12593 ; n12594
g12531 nor n12568 n12594 ; n12595
g12532 nor n12561 n12564 ; n12596
g12533 nor n12595 n12596 ; n12597
g12534 and n12565_not n12597 ; n12598
g12535 nor n12565 n12598 ; n12599
g12536 nor n12558 n12561 ; n12600
g12537 nor n12562 n12600 ; n12601
g12538 and n12599_not n12601 ; n12602
g12539 nor n12562 n12602 ; n12603
g12540 nor n12555 n12558 ; n12604
g12541 nor n12603 n12604 ; n12605
g12542 and n12559_not n12605 ; n12606
g12543 nor n12559 n12606 ; n12607
g12544 nor n12552 n12555 ; n12608
g12545 nor n12607 n12608 ; n12609
g12546 and n12556_not n12609 ; n12610
g12547 nor n12556 n12610 ; n12611
g12548 nor n12549 n12552 ; n12612
g12549 nor n12553 n12612 ; n12613
g12550 and n12611_not n12613 ; n12614
g12551 nor n12553 n12614 ; n12615
g12552 nor n12546 n12549 ; n12616
g12553 nor n12615 n12616 ; n12617
g12554 and n12550_not n12617 ; n12618
g12555 nor n12550 n12618 ; n12619
g12556 nor n12543 n12546 ; n12620
g12557 nor n12547 n12620 ; n12621
g12558 and n12619_not n12621 ; n12622
g12559 nor n12547 n12622 ; n12623
g12560 nor n12540 n12543 ; n12624
g12561 nor n12623 n12624 ; n12625
g12562 and n12544_not n12625 ; n12626
g12563 nor n12544 n12626 ; n12627
g12564 nor n12537 n12540 ; n12628
g12565 nor n12627 n12628 ; n12629
g12566 and n12541_not n12629 ; n12630
g12567 nor n12541 n12630 ; n12631
g12568 nor n12534 n12537 ; n12632
g12569 nor n12631 n12632 ; n12633
g12570 and n12538_not n12633 ; n12634
g12571 nor n12538 n12634 ; n12635
g12572 nor n12531 n12534 ; n12636
g12573 nor n12535 n12636 ; n12637
g12574 and n12635_not n12637 ; n12638
g12575 nor n12535 n12638 ; n12639
g12576 nor n12528 n12531 ; n12640
g12577 nor n12639 n12640 ; n12641
g12578 and n12532_not n12641 ; n12642
g12579 nor n12532 n12642 ; n12643
g12580 nor n12525 n12528 ; n12644
g12581 nor n12529 n12644 ; n12645
g12582 and n12643_not n12645 ; n12646
g12583 nor n12529 n12646 ; n12647
g12584 nor n12522 n12525 ; n12648
g12585 nor n12526 n12648 ; n12649
g12586 and n12647_not n12649 ; n12650
g12587 nor n12526 n12650 ; n12651
g12588 nor n12519 n12522 ; n12652
g12589 nor n12523 n12652 ; n12653
g12590 and n12651_not n12653 ; n12654
g12591 nor n12523 n12654 ; n12655
g12592 nor n12516 n12519 ; n12656
g12593 nor n12655 n12656 ; n12657
g12594 and n12520_not n12657 ; n12658
g12595 nor n12520 n12658 ; n12659
g12596 nor n12511 n12516 ; n12660
g12597 nor n12659 n12660 ; n12661
g12598 and n12517_not n12661 ; n12662
g12599 nor n12517 n12662 ; n12663
g12600 nor n12511 n12513 ; n12664
g12601 nor n12514 n12664 ; n12665
g12602 and n12663_not n12665 ; n12666
g12603 nor n12514 n12666 ; n12667
g12604 nor n12508 n12513 ; n12668
g12605 and n12508 n12513 ; n12669
g12606 nor n12668 n12669 ; n12670
g12607 and n12667_not n12670 ; n12671
g12608 nor n12669 n12671 ; n12672
g12609 nor n12505 n12508 ; n12673
g12610 nor n12672 n12673 ; n12674
g12611 and n12509_not n12674 ; n12675
g12612 nor n12509 n12675 ; n12676
g12613 nor n12370 n12505 ; n12677
g12614 nor n12676 n12677 ; n12678
g12615 and n12506_not n12678 ; n12679
g12616 nor n12506 n12679 ; n12680
g12617 nor n12370 n12502 ; n12681
g12618 nor n12680 n12681 ; n12682
g12619 and n12503_not n12682 ; n12683
g12620 nor n12503 n12683 ; n12684
g12621 nor n12497 n12500 ; n12685
g12622 nor n12489 n12493 ; n12686
g12623 and n3877_not n3967 ; n12687
g12624 and n4046 n4515_not ; n12688
g12625 nor n12687 n12688 ; n12689
g12626 and n4050 n4609 ; n12690
g12627 and n12689 n12690_not ; n12691
g12628 and a[26] n12691_not ; n12692
g12629 nor n12691 n12692 ; n12693
g12630 and a[26] n12692_not ; n12694
g12631 nor n12693 n12694 ; n12695
g12632 nor n12470 n12473 ; n12696
g12633 and n75 n3627 ; n12697
g12634 and n3020 n3456_not ; n12698
g12635 and n3023 n3539_not ; n12699
g12636 and n3028 n3605_not ; n12700
g12637 nor n12699 n12700 ; n12701
g12638 and n12698_not n12701 ; n12702
g12639 and n12697_not n12702 ; n12703
g12640 nor n169 n194 ; n12704
g12641 and n803_not n12704 ; n12705
g12642 and n1101_not n12705 ; n12706
g12643 and n419_not n12706 ; n12707
g12644 and n394_not n12707 ; n12708
g12645 and n657_not n12708 ; n12709
g12646 and n161_not n12709 ; n12710
g12647 nor n232 n393 ; n12711
g12648 and n201_not n12711 ; n12712
g12649 and n2361 n12712 ; n12713
g12650 and n1879 n12713 ; n12714
g12651 and n6054 n12714 ; n12715
g12652 and n5806 n12715 ; n12716
g12653 and n1549 n12716 ; n12717
g12654 and n2507 n12717 ; n12718
g12655 and n1577 n12718 ; n12719
g12656 and n2573 n12719 ; n12720
g12657 and n12710 n12720 ; n12721
g12658 and n120 n12721 ; n12722
g12659 and n4786 n12722 ; n12723
g12660 and n356 n12723 ; n12724
g12661 and n116 n12724 ; n12725
g12662 and n154_not n12725 ; n12726
g12663 and n715_not n12726 ; n12727
g12664 and n102_not n12727 ; n12728
g12665 and n277_not n12728 ; n12729
g12666 and n270_not n12729 ; n12730
g12667 and n12454_not n12730 ; n12731
g12668 and n12454 n12730_not ; n12732
g12669 nor n12731 n12732 ; n12733
g12670 and n12703_not n12733 ; n12734
g12671 nor n12703 n12734 ; n12735
g12672 and n12733 n12734_not ; n12736
g12673 nor n12735 n12736 ; n12737
g12674 nor n12464 n12467 ; n12738
g12675 and n12737 n12738 ; n12739
g12676 nor n12737 n12738 ; n12740
g12677 nor n12739 n12740 ; n12741
g12678 and n3457 n4045_not ; n12742
g12679 and n3542 n3805_not ; n12743
g12680 and n3606 n3964_not ; n12744
g12681 nor n12743 n12744 ; n12745
g12682 and n12742_not n12745 ; n12746
g12683 and n3368_not n12746 ; n12747
g12684 and n4477_not n12746 ; n12748
g12685 nor n12747 n12748 ; n12749
g12686 and a[29] n12749_not ; n12750
g12687 and a[29]_not n12749 ; n12751
g12688 nor n12750 n12751 ; n12752
g12689 and n12741 n12752_not ; n12753
g12690 and n12741_not n12752 ; n12754
g12691 nor n12753 n12754 ; n12755
g12692 and n12696_not n12755 ; n12756
g12693 nor n12696 n12756 ; n12757
g12694 and n12755 n12756_not ; n12758
g12695 nor n12757 n12758 ; n12759
g12696 nor n12695 n12759 ; n12760
g12697 and n12695 n12758_not ; n12761
g12698 and n12757_not n12761 ; n12762
g12699 nor n12760 n12762 ; n12763
g12700 and n12686_not n12763 ; n12764
g12701 and n12686 n12763_not ; n12765
g12702 nor n12764 n12765 ; n12766
g12703 and n12685_not n12766 ; n12767
g12704 and n12685 n12766_not ; n12768
g12705 nor n12767 n12768 ; n12769
g12706 nor n12502 n12769 ; n12770
g12707 and n12502 n12769 ; n12771
g12708 nor n12770 n12771 ; n12772
g12709 and n12684_not n12772 ; n12773
g12710 nor n12771 n12773 ; n12774
g12711 nor n12764 n12767 ; n12775
g12712 nor n12756 n12760 ; n12776
g12713 and n75 n3818 ; n12777
g12714 and n3020 n3805_not ; n12778
g12715 and n3023 n3605_not ; n12779
g12716 and n3028 n3456_not ; n12780
g12717 nor n12779 n12780 ; n12781
g12718 and n12778_not n12781 ; n12782
g12719 and n12777_not n12782 ; n12783
g12720 nor n224 n305 ; n12784
g12721 and n714_not n12784 ; n12785
g12722 and n653 n12785 ; n12786
g12723 and n2573 n12786 ; n12787
g12724 and n2582 n12787 ; n12788
g12725 and n276_not n12788 ; n12789
g12726 and n460_not n12789 ; n12790
g12727 and n932_not n12790 ; n12791
g12728 and n273_not n12791 ; n12792
g12729 and n225_not n12792 ; n12793
g12730 and n712_not n12793 ; n12794
g12731 and n231_not n12794 ; n12795
g12732 and n561 n5808 ; n12796
g12733 and n1476 n12796 ; n12797
g12734 and n968 n12797 ; n12798
g12735 and n2170 n12798 ; n12799
g12736 and n282 n12799 ; n12800
g12737 and n1247 n12800 ; n12801
g12738 and n206_not n12801 ; n12802
g12739 and n673_not n12802 ; n12803
g12740 and n531_not n12803 ; n12804
g12741 and n1104_not n12804 ; n12805
g12742 nor n462 n667 ; n12806
g12743 and n151_not n12806 ; n12807
g12744 and n1062_not n12807 ; n12808
g12745 and n451_not n12808 ; n12809
g12746 and n125_not n12809 ; n12810
g12747 nor n403 n506 ; n12811
g12748 and n601_not n12811 ; n12812
g12749 and n1527 n12812 ; n12813
g12750 and n12810 n12813 ; n12814
g12751 and n12805 n12814 ; n12815
g12752 and n4794 n12815 ; n12816
g12753 and n202 n12816 ; n12817
g12754 and n190_not n12817 ; n12818
g12755 and n255_not n12818 ; n12819
g12756 and n239_not n12819 ; n12820
g12757 and n121_not n12820 ; n12821
g12758 and n402_not n12821 ; n12822
g12759 and n287_not n12822 ; n12823
g12760 and n302_not n12823 ; n12824
g12761 and n243_not n12824 ; n12825
g12762 and n519_not n12825 ; n12826
g12763 and n271_not n12826 ; n12827
g12764 and n429_not n12827 ; n12828
g12765 nor n334 n435 ; n12829
g12766 and n252_not n12829 ; n12830
g12767 and n3827 n12830 ; n12831
g12768 and n6084 n12831 ; n12832
g12769 and n12828 n12832 ; n12833
g12770 and n12795 n12833 ; n12834
g12771 and n1479 n12834 ; n12835
g12772 and n159 n12835 ; n12836
g12773 and n1667 n12836 ; n12837
g12774 and n570 n12837 ; n12838
g12775 and n284_not n12838 ; n12839
g12776 and n191_not n12839 ; n12840
g12777 and n452_not n12840 ; n12841
g12778 and n474_not n12841 ; n12842
g12779 and n12730_not n12842 ; n12843
g12780 and n12730 n12842_not ; n12844
g12781 nor n12783 n12844 ; n12845
g12782 and n12843_not n12845 ; n12846
g12783 nor n12783 n12846 ; n12847
g12784 nor n12844 n12846 ; n12848
g12785 and n12843_not n12848 ; n12849
g12786 nor n12847 n12849 ; n12850
g12787 nor n12731 n12734 ; n12851
g12788 and n12850 n12851 ; n12852
g12789 nor n12850 n12851 ; n12853
g12790 nor n12852 n12853 ; n12854
g12791 nor n12740 n12753 ; n12855
g12792 and n12854 n12855_not ; n12856
g12793 and n12854_not n12855 ; n12857
g12794 nor n12856 n12857 ; n12858
g12795 and n4050 n4522 ; n12859
g12796 and n3967 n4515_not ; n12860
g12797 nor n12859 n12860 ; n12861
g12798 and a[26] n12861_not ; n12862
g12799 nor n12861 n12862 ; n12863
g12800 and a[26] n12862_not ; n12864
g12801 nor n12863 n12864 ; n12865
g12802 and n3457 n3877_not ; n12866
g12803 and n3542 n3964_not ; n12867
g12804 and n3606 n4045_not ; n12868
g12805 nor n12867 n12868 ; n12869
g12806 and n12866_not n12869 ; n12870
g12807 and n3368 n4067 ; n12871
g12808 and n12870 n12871_not ; n12872
g12809 and a[29] n12872_not ; n12873
g12810 and a[29] n12873_not ; n12874
g12811 nor n12872 n12873 ; n12875
g12812 nor n12874 n12875 ; n12876
g12813 nor n12865 n12876 ; n12877
g12814 nor n12865 n12877 ; n12878
g12815 nor n12876 n12877 ; n12879
g12816 nor n12878 n12879 ; n12880
g12817 and n12858 n12880_not ; n12881
g12818 and n12858_not n12880 ; n12882
g12819 nor n12881 n12882 ; n12883
g12820 and n12776_not n12883 ; n12884
g12821 and n12776 n12883_not ; n12885
g12822 nor n12884 n12885 ; n12886
g12823 and n12775_not n12886 ; n12887
g12824 and n12775 n12886_not ; n12888
g12825 nor n12887 n12888 ; n12889
g12826 nor n12769 n12889 ; n12890
g12827 and n12769 n12889 ; n12891
g12828 nor n12890 n12891 ; n12892
g12829 and n12774_not n12892 ; n12893
g12830 and n12774 n12892_not ; n12894
g12831 nor n12893 n12894 ; n12895
g12832 and n75 n12895 ; n12896
g12833 and n3020 n12889 ; n12897
g12834 and n3023 n12502 ; n12898
g12835 and n3028 n12769 ; n12899
g12836 nor n12898 n12899 ; n12900
g12837 and n12897_not n12900 ; n12901
g12838 and n12896_not n12901 ; n12902
g12839 nor n276 n667 ; n12903
g12840 and n190_not n12903 ; n12904
g12841 and n1101_not n12904 ; n12905
g12842 and n396_not n12905 ; n12906
g12843 and n453_not n12906 ; n12907
g12844 and n422_not n12907 ; n12908
g12845 and n132_not n12908 ; n12909
g12846 and n230 n306_not ; n12910
g12847 and n272_not n12910 ; n12911
g12848 and n1611 n4327 ; n12912
g12849 and n12911 n12912 ; n12913
g12850 and n155_not n12913 ; n12914
g12851 and n402_not n12914 ; n12915
g12852 and n1104_not n12915 ; n12916
g12853 and n883_not n12916 ; n12917
g12854 and n337_not n12917 ; n12918
g12855 and n188_not n12918 ; n12919
g12856 and n239_not n2092 ; n12920
g12857 and n825_not n12920 ; n12921
g12858 and n601_not n12921 ; n12922
g12859 and n567_not n12922 ; n12923
g12860 and n293_not n12923 ; n12924
g12861 and n1994 n6520 ; n12925
g12862 and n1782 n12925 ; n12926
g12863 and n111_not n12926 ; n12927
g12864 and n242_not n12927 ; n12928
g12865 and n327_not n12928 ; n12929
g12866 and n147_not n12929 ; n12930
g12867 and n395_not n12930 ; n12931
g12868 and n86_not n12931 ; n12932
g12869 and n640 n5040 ; n12933
g12870 and n12932 n12933 ; n12934
g12871 and n12924 n12934 ; n12935
g12872 and n2443 n12935 ; n12936
g12873 and n136_not n12936 ; n12937
g12874 and n886_not n12937 ; n12938
g12875 and n358_not n12938 ; n12939
g12876 nor n355 n1011 ; n12940
g12877 and n171_not n12940 ; n12941
g12878 and n373 n12941 ; n12942
g12879 and n1237 n12942 ; n12943
g12880 and n564_not n12943 ; n12944
g12881 and n638 n2230 ; n12945
g12882 and n1249 n12945 ; n12946
g12883 and n2468 n12946 ; n12947
g12884 and n12944 n12947 ; n12948
g12885 and n12939 n12948 ; n12949
g12886 and n2623 n12949 ; n12950
g12887 and n12919 n12950 ; n12951
g12888 and n12909 n12951 ; n12952
g12889 and n1129 n12952 ; n12953
g12890 and n4295 n12953 ; n12954
g12891 and n330_not n12954 ; n12955
g12892 and n254_not n12955 ; n12956
g12893 and n292_not n12956 ; n12957
g12894 and n91_not n12957 ; n12958
g12895 and n2684 n3438 ; n12959
g12896 and n530 n12959 ; n12960
g12897 and n1925 n12960 ; n12961
g12898 and n789 n12961 ; n12962
g12899 and n1254 n12962 ; n12963
g12900 and n1827 n12963 ; n12964
g12901 and n1161 n12964 ; n12965
g12902 and n847_not n12965 ; n12966
g12903 and n619_not n12966 ; n12967
g12904 and n155_not n12967 ; n12968
g12905 and n637_not n12968 ; n12969
g12906 and n980_not n12969 ; n12970
g12907 and n394_not n12970 ; n12971
g12908 and n225_not n12971 ; n12972
g12909 and n332_not n12972 ; n12973
g12910 nor n281 n426 ; n12974
g12911 and n189_not n12974 ; n12975
g12912 and n461_not n12975 ; n12976
g12913 and n231_not n12976 ; n12977
g12914 and n3985 n4334 ; n12978
g12915 and n12977 n12978 ; n12979
g12916 and n1216 n12979 ; n12980
g12917 and n5224 n12980 ; n12981
g12918 and n1969 n12981 ; n12982
g12919 and n12973 n12982 ; n12983
g12920 and n1523 n12983 ; n12984
g12921 and n2633 n12984 ; n12985
g12922 and n1825 n12985 ; n12986
g12923 and n1252 n12986 ; n12987
g12924 and n242_not n12987 ; n12988
g12925 and n355_not n12988 ; n12989
g12926 and n495_not n12989 ; n12990
g12927 and n246_not n12990 ; n12991
g12928 and n6706 n12991 ; n12992
g12929 and n375_not n12992 ; n12993
g12930 and n237_not n12993 ; n12994
g12931 and n564_not n12994 ; n12995
g12932 and n12958 n12995_not ; n12996
g12933 and n12958_not n12995 ; n12997
g12934 and n12684 n12772_not ; n12998
g12935 nor n12773 n12998 ; n12999
g12936 and n75 n12999 ; n13000
g12937 and n3020 n12769 ; n13001
g12938 and n3023 n12370 ; n13002
g12939 and n3028 n12502 ; n13003
g12940 nor n13002 n13003 ; n13004
g12941 and n13001_not n13004 ; n13005
g12942 and n13000_not n13005 ; n13006
g12943 nor n12996 n13006 ; n13007
g12944 and n12997_not n13007 ; n13008
g12945 nor n12996 n13008 ; n13009
g12946 and n169_not n238 ; n13010
g12947 and n514_not n13010 ; n13011
g12948 and n119_not n13011 ; n13012
g12949 nor n353 n847 ; n13013
g12950 and n326_not n13013 ; n13014
g12951 nor n419 n689 ; n13015
g12952 and n493_not n13015 ; n13016
g12953 and n13014 n13016 ; n13017
g12954 and n1693 n13017 ; n13018
g12955 and n13012 n13018 ; n13019
g12956 and n12795 n13019 ; n13020
g12957 and n1511 n13020 ; n13021
g12958 and n2782 n13021 ; n13022
g12959 and n2507 n13022 ; n13023
g12960 and n1827 n13023 ; n13024
g12961 and n1248 n13024 ; n13025
g12962 and n301_not n13025 ; n13026
g12963 and n278_not n13026 ; n13027
g12964 and n115_not n13027 ; n13028
g12965 and n91_not n13028 ; n13029
g12966 and n504_not n13029 ; n13030
g12967 and n436_not n13030 ; n13031
g12968 and n1556 n4151 ; n13032
g12969 and n897 n13032 ; n13033
g12970 and n591 n13033 ; n13034
g12971 and n656_not n13034 ; n13035
g12972 and n594_not n13035 ; n13036
g12973 and n417_not n13036 ; n13037
g12974 and n527_not n13037 ; n13038
g12975 and n165_not n13038 ; n13039
g12976 and n672_not n13039 ; n13040
g12977 and n293_not n13040 ; n13041
g12978 and n2020 n6664 ; n13042
g12979 and n593 n13042 ; n13043
g12980 and n6607 n13043 ; n13044
g12981 and n12828 n13044 ; n13045
g12982 and n13041 n13045 ; n13046
g12983 and n1521 n13046 ; n13047
g12984 and n13031 n13047 ; n13048
g12985 and n1029 n13048 ; n13049
g12986 and n291 n13049 ; n13050
g12987 and n1139 n13050 ; n13051
g12988 and n826 n13051 ; n13052
g12989 and n1389 n13052 ; n13053
g12990 and n341 n13053 ; n13054
g12991 and n1102_not n13054 ; n13055
g12992 and n1127_not n13055 ; n13056
g12993 and n3831 n13056 ; n13057
g12994 and n193 n13057 ; n13058
g12995 and n452_not n13058 ; n13059
g12996 and n1255 n1781 ; n13060
g12997 and n3984 n13060 ; n13061
g12998 and n589_not n13061 ; n13062
g12999 and n449_not n13062 ; n13063
g13000 and n2265 n3906 ; n13064
g13001 and n3580 n13064 ; n13065
g13002 and n5233 n13065 ; n13066
g13003 and n4017 n13066 ; n13067
g13004 and n13063 n13067 ; n13068
g13005 and n4502 n13068 ; n13069
g13006 and n3848 n13069 ; n13070
g13007 and n2738 n13070 ; n13071
g13008 and n2583 n13071 ; n13072
g13009 and n242_not n13072 ; n13073
g13010 and n518_not n13073 ; n13074
g13011 and n3569 n3906 ; n13075
g13012 and n3832 n4034 ; n13076
g13013 and n13075 n13076 ; n13077
g13014 and n3869 n13077 ; n13078
g13015 and n328_not n13078 ; n13079
g13016 and n536_not n13079 ; n13080
g13017 and n567_not n13080 ; n13081
g13018 and n13074 n13081 ; n13082
g13019 and n13059_not n13082 ; n13083
g13020 and n3570 n3832 ; n13084
g13021 and n539 n13084 ; n13085
g13022 and n968 n13085 ; n13086
g13023 and n453_not n13086 ; n13087
g13024 and n3949 n13087 ; n13088
g13025 and n3856 n13088 ; n13089
g13026 and n4493 n13089 ; n13090
g13027 and n665 n13090 ; n13091
g13028 and n1761 n13091 ; n13092
g13029 and n601_not n13092 ; n13093
g13030 and n673_not n13093 ; n13094
g13031 and n99_not n13094 ; n13095
g13032 and n13074 n13095_not ; n13096
g13033 and n13074_not n13095 ; n13097
g13034 and n75 n4522 ; n13098
g13035 and n3023 n4515_not ; n13099
g13036 nor n13098 n13099 ; n13100
g13037 nor n13096 n13100 ; n13101
g13038 and n13097_not n13101 ; n13102
g13039 nor n13096 n13102 ; n13103
g13040 nor n13074 n13081 ; n13104
g13041 nor n13082 n13104 ; n13105
g13042 nor n13103 n13105 ; n13106
g13043 nor n13103 n13106 ; n13107
g13044 nor n13105 n13106 ; n13108
g13045 nor n13107 n13108 ; n13109
g13046 nor n13100 n13102 ; n13110
g13047 and n13097_not n13103 ; n13111
g13048 nor n13110 n13111 ; n13112
g13049 nor n283 n1306 ; n13113
g13050 and n249_not n13113 ; n13114
g13051 and n12397 n13114 ; n13115
g13052 and n4216 n13115 ; n13116
g13053 and n1916 n13116 ; n13117
g13054 and n305_not n13117 ; n13118
g13055 and n403_not n13118 ; n13119
g13056 and n246_not n13119 ; n13120
g13057 and n519_not n13120 ; n13121
g13058 and n125_not n13121 ; n13122
g13059 and n293_not n13122 ; n13123
g13060 and n530 n3570 ; n13124
g13061 and n2740 n13124 ; n13125
g13062 and n232_not n13125 ; n13126
g13063 and n289_not n13126 ; n13127
g13064 and n149_not n13127 ; n13128
g13065 and n226_not n13128 ; n13129
g13066 and n490_not n13129 ; n13130
g13067 and n496_not n13130 ; n13131
g13068 and n157_not n13131 ; n13132
g13069 and n623_not n13132 ; n13133
g13070 and n86_not n13133 ; n13134
g13071 and n771_not n13134 ; n13135
g13072 and n167_not n13135 ; n13136
g13073 and n165_not n13136 ; n13137
g13074 and n158_not n13137 ; n13138
g13075 and n1163 n2544 ; n13139
g13076 and n13138 n13139 ; n13140
g13077 and n1735 n13140 ; n13141
g13078 and n1202 n13141 ; n13142
g13079 and n13123 n13142 ; n13143
g13080 and n5085 n13143 ; n13144
g13081 and n2635 n13144 ; n13145
g13082 and n1366 n13145 ; n13146
g13083 and n730 n13146 ; n13147
g13084 and n1252 n13147 ; n13148
g13085 and n2466 n13148 ; n13149
g13086 and n978 n13149 ; n13150
g13087 and n123_not n13150 ; n13151
g13088 and n847_not n13151 ; n13152
g13089 and n284_not n13152 ; n13153
g13090 and n367_not n13153 ; n13154
g13091 and n292_not n13154 ; n13155
g13092 and n274_not n13155 ; n13156
g13093 and n525_not n13156 ; n13157
g13094 and n672_not n13157 ; n13158
g13095 and n3929 n5064 ; n13159
g13096 and n885 n13159 ; n13160
g13097 and n144_not n13160 ; n13161
g13098 and n1425 n1740 ; n13162
g13099 and n1249 n13162 ; n13163
g13100 and n13161 n13163 ; n13164
g13101 and n13087 n13164 ; n13165
g13102 and n3947 n13165 ; n13166
g13103 and n13063 n13166 ; n13167
g13104 and n4009 n13167 ; n13168
g13105 and n1046 n13168 ; n13169
g13106 and n567_not n13169 ; n13170
g13107 and n525_not n13170 ; n13171
g13108 and n293_not n13171 ; n13172
g13109 nor n13158 n13172 ; n13173
g13110 and n13158 n13172 ; n13174
g13111 nor n13173 n13174 ; n13175
g13112 and a[29]_not n13175 ; n13176
g13113 nor n13173 n13176 ; n13177
g13114 and n13074 n13177_not ; n13178
g13115 and n75 n4609 ; n13179
g13116 and n3023 n3877_not ; n13180
g13117 and n3028 n4515_not ; n13181
g13118 nor n13180 n13181 ; n13182
g13119 and n13179_not n13182 ; n13183
g13120 and n13074_not n13177 ; n13184
g13121 nor n13178 n13184 ; n13185
g13122 and n13183_not n13185 ; n13186
g13123 nor n13178 n13186 ; n13187
g13124 nor n13112 n13187 ; n13188
g13125 and n13112 n13187 ; n13189
g13126 nor n13188 n13189 ; n13190
g13127 nor n13183 n13186 ; n13191
g13128 and n13185 n13186_not ; n13192
g13129 nor n13191 n13192 ; n13193
g13130 nor a[29] n13176 ; n13194
g13131 and n13174_not n13177 ; n13195
g13132 nor n13194 n13195 ; n13196
g13133 and n1138 n3300 ; n13197
g13134 and n775 n13197 ; n13198
g13135 and n288 n13198 ; n13199
g13136 and n471 n13199 ; n13200
g13137 and n1726 n13200 ; n13201
g13138 and n1040 n13201 ; n13202
g13139 and n752_not n13202 ; n13203
g13140 and n354_not n13203 ; n13204
g13141 and n402_not n13204 ; n13205
g13142 and n505_not n13205 ; n13206
g13143 and n466_not n13206 ; n13207
g13144 and n961_not n13207 ; n13208
g13145 and n332_not n13208 ; n13209
g13146 and n95_not n13209 ; n13210
g13147 and n621 n3459 ; n13211
g13148 and n826 n13211 ; n13212
g13149 and n713_not n13212 ; n13213
g13150 and n151_not n13213 ; n13214
g13151 and n328_not n13214 ; n13215
g13152 and n417_not n13215 ; n13216
g13153 and n367_not n13216 ; n13217
g13154 and n91_not n13217 ; n13218
g13155 and n132_not n13218 ; n13219
g13156 and n200_not n13219 ; n13220
g13157 and n655_not n13220 ; n13221
g13158 and n3115 n5787 ; n13222
g13159 and n624 n13222 ; n13223
g13160 and n494 n13223 ; n13224
g13161 and n2987 n13224 ; n13225
g13162 and n13221 n13225 ; n13226
g13163 and n13210 n13226 ; n13227
g13164 and n6707 n13227 ; n13228
g13165 and n4232 n13228 ; n13229
g13166 and n1254 n13229 ; n13230
g13167 and n1531 n13230 ; n13231
g13168 and n224_not n13231 ; n13232
g13169 and n715_not n13232 ; n13233
g13170 and n568_not n13233 ; n13234
g13171 and n492_not n13234 ; n13235
g13172 and n504_not n13235 ; n13236
g13173 and n453_not n13236 ; n13237
g13174 and n170_not n13237 ; n13238
g13175 and n13158 n13238_not ; n13239
g13176 and n13158_not n13238 ; n13240
g13177 and n4797 n12412 ; n13241
g13178 and n1826 n13241 ; n13242
g13179 and n418 n13242 ; n13243
g13180 and n352_not n13243 ; n13244
g13181 and n144_not n13244 ; n13245
g13182 and n325_not n13245 ; n13246
g13183 and n449_not n13246 ; n13247
g13184 nor n146 n713 ; n13248
g13185 and n127_not n13248 ; n13249
g13186 and n691 n13249 ; n13250
g13187 and n6084 n13250 ; n13251
g13188 and n6083 n13251 ; n13252
g13189 and n1292 n13252 ; n13253
g13190 and n3544 n13253 ; n13254
g13191 and n285 n13254 ; n13255
g13192 and n1825 n13255 ; n13256
g13193 and n1366 n13256 ; n13257
g13194 and n236_not n13257 ; n13258
g13195 and n1306_not n13258 ; n13259
g13196 and n1102_not n13259 ; n13260
g13197 and n287_not n13260 ; n13261
g13198 and n490_not n13261 ; n13262
g13199 and n192_not n13262 ; n13263
g13200 and n246_not n13263 ; n13264
g13201 and n666_not n13264 ; n13265
g13202 and n366_not n590 ; n13266
g13203 and n125_not n13266 ; n13267
g13204 and n428_not n13267 ; n13268
g13205 and n3645 n6104 ; n13269
g13206 and n1557 n13269 ; n13270
g13207 and n13268 n13270 ; n13271
g13208 and n2772 n13271 ; n13272
g13209 and n13265 n13272 ; n13273
g13210 and n13247 n13273 ; n13274
g13211 and n2090 n13274 ; n13275
g13212 and n1330 n13275 ; n13276
g13213 and n2406 n13276 ; n13277
g13214 and n156 n13277 ; n13278
g13215 and n279 n13278 ; n13279
g13216 and n232_not n13279 ; n13280
g13217 and n327_not n13280 ; n13281
g13218 and n145_not n13281 ; n13282
g13219 and n165_not n13282 ; n13283
g13220 nor n12730 n13283 ; n13284
g13221 and n12730 n13283 ; n13285
g13222 nor n13284 n13285 ; n13286
g13223 and a[26]_not n13286 ; n13287
g13224 nor n13284 n13287 ; n13288
g13225 and n13238 n13288_not ; n13289
g13226 and n75 n4477 ; n13290
g13227 and n3020 n4045_not ; n13291
g13228 and n3023 n3805_not ; n13292
g13229 and n3028 n3964_not ; n13293
g13230 nor n13292 n13293 ; n13294
g13231 and n13291_not n13294 ; n13295
g13232 and n13290_not n13295 ; n13296
g13233 and n13238_not n13288 ; n13297
g13234 nor n13289 n13297 ; n13298
g13235 and n13296_not n13298 ; n13299
g13236 nor n13289 n13299 ; n13300
g13237 nor n13239 n13300 ; n13301
g13238 and n13240_not n13301 ; n13302
g13239 nor n13239 n13302 ; n13303
g13240 nor n13196 n13303 ; n13304
g13241 and n75 n4715 ; n13305
g13242 and n3020 n4515_not ; n13306
g13243 and n3023 n4045_not ; n13307
g13244 and n3028 n3877_not ; n13308
g13245 nor n13307 n13308 ; n13309
g13246 and n13306_not n13309 ; n13310
g13247 and n13305_not n13310 ; n13311
g13248 and n13196 n13303 ; n13312
g13249 nor n13304 n13312 ; n13313
g13250 and n13311_not n13313 ; n13314
g13251 nor n13304 n13314 ; n13315
g13252 nor n13193 n13315 ; n13316
g13253 and n13193 n13315 ; n13317
g13254 nor n13316 n13317 ; n13318
g13255 and n3542 n4515_not ; n13319
g13256 and n3368 n4522 ; n13320
g13257 nor n13319 n13320 ; n13321
g13258 and a[29] n13321_not ; n13322
g13259 nor n13321 n13322 ; n13323
g13260 and a[29] n13322_not ; n13324
g13261 nor n13323 n13324 ; n13325
g13262 and n75 n4067 ; n13326
g13263 and n3020 n3877_not ; n13327
g13264 and n3023 n3964_not ; n13328
g13265 and n3028 n4045_not ; n13329
g13266 nor n13328 n13329 ; n13330
g13267 and n13327_not n13330 ; n13331
g13268 and n13326_not n13331 ; n13332
g13269 nor n13325 n13332 ; n13333
g13270 nor n13325 n13333 ; n13334
g13271 nor n13332 n13333 ; n13335
g13272 nor n13334 n13335 ; n13336
g13273 nor n13300 n13302 ; n13337
g13274 and n13240_not n13303 ; n13338
g13275 nor n13337 n13338 ; n13339
g13276 nor n13336 n13339 ; n13340
g13277 nor n13333 n13340 ; n13341
g13278 and n13311 n13313_not ; n13342
g13279 nor n13314 n13342 ; n13343
g13280 and n13341_not n13343 ; n13344
g13281 nor n13296 n13299 ; n13345
g13282 and n13298 n13299_not ; n13346
g13283 nor n13345 n13346 ; n13347
g13284 nor a[26] n13287 ; n13348
g13285 and n13285_not n13288 ; n13349
g13286 nor n13348 n13349 ; n13350
g13287 nor n12848 n13350 ; n13351
g13288 and n75 n4558 ; n13352
g13289 and n3020 n3964_not ; n13353
g13290 and n3023 n3456_not ; n13354
g13291 and n3028 n3805_not ; n13355
g13292 nor n13354 n13355 ; n13356
g13293 and n13353_not n13356 ; n13357
g13294 and n13352_not n13357 ; n13358
g13295 and n12848 n13350 ; n13359
g13296 nor n13351 n13359 ; n13360
g13297 and n13358_not n13360 ; n13361
g13298 nor n13351 n13361 ; n13362
g13299 nor n13347 n13362 ; n13363
g13300 and n13347 n13362 ; n13364
g13301 nor n13363 n13364 ; n13365
g13302 and n3542 n3877_not ; n13366
g13303 and n3606 n4515_not ; n13367
g13304 nor n13366 n13367 ; n13368
g13305 and n3368 n4609 ; n13369
g13306 and n13368 n13369_not ; n13370
g13307 and a[29] n13370_not ; n13371
g13308 and a[29] n13371_not ; n13372
g13309 nor n13370 n13371 ; n13373
g13310 nor n13372 n13373 ; n13374
g13311 and n13365 n13374_not ; n13375
g13312 nor n13363 n13375 ; n13376
g13313 and n13336_not n13339 ; n13377
g13314 and n13336 n13339_not ; n13378
g13315 nor n13377 n13378 ; n13379
g13316 nor n13376 n13379 ; n13380
g13317 and n13365 n13375_not ; n13381
g13318 nor n13374 n13375 ; n13382
g13319 nor n13381 n13382 ; n13383
g13320 nor n12853 n12856 ; n13384
g13321 nor n13358 n13361 ; n13385
g13322 and n13360 n13361_not ; n13386
g13323 nor n13385 n13386 ; n13387
g13324 nor n13384 n13387 ; n13388
g13325 nor n13384 n13388 ; n13389
g13326 nor n13387 n13388 ; n13390
g13327 nor n13389 n13390 ; n13391
g13328 and n3457 n4515_not ; n13392
g13329 and n3542 n4045_not ; n13393
g13330 and n3606 n3877_not ; n13394
g13331 nor n13393 n13394 ; n13395
g13332 and n13392_not n13395 ; n13396
g13333 and n3368 n4715 ; n13397
g13334 and n13396 n13397_not ; n13398
g13335 and a[29] n13398_not ; n13399
g13336 and a[29] n13399_not ; n13400
g13337 nor n13398 n13399 ; n13401
g13338 nor n13400 n13401 ; n13402
g13339 nor n13391 n13402 ; n13403
g13340 nor n13388 n13403 ; n13404
g13341 nor n13383 n13404 ; n13405
g13342 and n13383 n13404 ; n13406
g13343 nor n13405 n13406 ; n13407
g13344 nor n13391 n13403 ; n13408
g13345 nor n13402 n13403 ; n13409
g13346 nor n13408 n13409 ; n13410
g13347 nor n12877 n12881 ; n13411
g13348 nor n13410 n13411 ; n13412
g13349 nor n13410 n13412 ; n13413
g13350 nor n13411 n13412 ; n13414
g13351 nor n13413 n13414 ; n13415
g13352 nor n12884 n12887 ; n13416
g13353 nor n13415 n13416 ; n13417
g13354 nor n13412 n13417 ; n13418
g13355 and n13407 n13418_not ; n13419
g13356 nor n13405 n13419 ; n13420
g13357 and n13376 n13379 ; n13421
g13358 nor n13380 n13421 ; n13422
g13359 and n13420_not n13422 ; n13423
g13360 nor n13380 n13423 ; n13424
g13361 and n13341 n13343_not ; n13425
g13362 nor n13344 n13425 ; n13426
g13363 and n13424_not n13426 ; n13427
g13364 nor n13344 n13427 ; n13428
g13365 and n13318 n13428_not ; n13429
g13366 nor n13316 n13429 ; n13430
g13367 and n13190 n13430_not ; n13431
g13368 nor n13188 n13431 ; n13432
g13369 nor n13109 n13432 ; n13433
g13370 nor n13106 n13433 ; n13434
g13371 and n13059 n13082_not ; n13435
g13372 nor n13434 n13435 ; n13436
g13373 and n13083_not n13436 ; n13437
g13374 and n13059_not n13437 ; n13438
g13375 nor n5407 n5496 ; n13439
g13376 and n4935_not n13439 ; n13440
g13377 and n4938_not n13440 ; n13441
g13378 nor n13438 n13441 ; n13442
g13379 and a[20] n13442_not ; n13443
g13380 and a[20]_not n13442 ; n13444
g13381 nor n13443 n13444 ; n13445
g13382 and n336 n5002 ; n13446
g13383 and n2595 n13446 ; n13447
g13384 and n3435 n13447 ; n13448
g13385 and n1894 n13448 ; n13449
g13386 and n1245 n13449 ; n13450
g13387 and n241 n13450 ; n13451
g13388 and n294 n13451 ; n13452
g13389 and n1252 n13452 ; n13453
g13390 and n229_not n13453 ; n13454
g13391 and n232_not n13454 ; n13455
g13392 and n284_not n13455 ; n13456
g13393 and n712_not n13456 ; n13457
g13394 and n562_not n13457 ; n13458
g13395 and n694 n3192 ; n13459
g13396 and n2806 n13459 ; n13460
g13397 and n988 n13460 ; n13461
g13398 and n805 n13461 ; n13462
g13399 and n13458 n13462 ; n13463
g13400 and n1708 n13463 ; n13464
g13401 and n621 n13464 ; n13465
g13402 and n450 n13465 ; n13466
g13403 and n869 n13466 ; n13467
g13404 and n557_not n13467 ; n13468
g13405 and n255_not n13468 ; n13469
g13406 and n252_not n13469 ; n13470
g13407 and n883_not n13470 ; n13471
g13408 and n569_not n13471 ; n13472
g13409 and n771_not n13472 ; n13473
g13410 and n875_not n13473 ; n13474
g13411 and n12958 n13474 ; n13475
g13412 nor n12958 n13474 ; n13476
g13413 nor n13475 n13476 ; n13477
g13414 and n13445 n13477 ; n13478
g13415 nor n13445 n13477 ; n13479
g13416 nor n13478 n13479 ; n13480
g13417 and n13009_not n13480 ; n13481
g13418 and n13009 n13480_not ; n13482
g13419 nor n13481 n13482 ; n13483
g13420 and n12902_not n13483 ; n13484
g13421 nor n13481 n13484 ; n13485
g13422 nor n13476 n13478 ; n13486
g13423 and n13031 n13486_not ; n13487
g13424 and n13031_not n13486 ; n13488
g13425 nor n13487 n13488 ; n13489
g13426 and n13415 n13416 ; n13490
g13427 nor n13417 n13490 ; n13491
g13428 and n3020 n13491 ; n13492
g13429 and n3028 n12889 ; n13493
g13430 and n3023 n12769 ; n13494
g13431 nor n12891 n12893 ; n13495
g13432 and n12889 n13491 ; n13496
g13433 nor n12889 n13491 ; n13497
g13434 nor n13495 n13497 ; n13498
g13435 and n13496_not n13498 ; n13499
g13436 nor n13495 n13499 ; n13500
g13437 nor n13496 n13499 ; n13501
g13438 and n13497_not n13501 ; n13502
g13439 nor n13500 n13502 ; n13503
g13440 and n75 n13503_not ; n13504
g13441 nor n13494 n13504 ; n13505
g13442 and n13493_not n13505 ; n13506
g13443 and n13492_not n13506 ; n13507
g13444 and n13489 n13507_not ; n13508
g13445 and n13489_not n13507 ; n13509
g13446 nor n13508 n13509 ; n13510
g13447 and n13485_not n13510 ; n13511
g13448 and n13485 n13510_not ; n13512
g13449 nor n13511 n13512 ; n13513
g13450 and n13424 n13426_not ; n13514
g13451 nor n13427 n13514 ; n13515
g13452 and n3457 n13515 ; n13516
g13453 and n13407_not n13418 ; n13517
g13454 nor n13419 n13517 ; n13518
g13455 and n3542 n13518 ; n13519
g13456 and n13420 n13422_not ; n13520
g13457 nor n13423 n13520 ; n13521
g13458 and n3606 n13521 ; n13522
g13459 nor n13519 n13522 ; n13523
g13460 and n13516_not n13523 ; n13524
g13461 and n3368_not n13524 ; n13525
g13462 and n13518 n13521 ; n13526
g13463 and n13491 n13518 ; n13527
g13464 nor n13491 n13518 ; n13528
g13465 nor n13527 n13528 ; n13529
g13466 and n13501_not n13529 ; n13530
g13467 nor n13527 n13530 ; n13531
g13468 nor n13518 n13521 ; n13532
g13469 nor n13531 n13532 ; n13533
g13470 and n13526_not n13533 ; n13534
g13471 nor n13526 n13534 ; n13535
g13472 nor n13515 n13521 ; n13536
g13473 and n13515 n13521 ; n13537
g13474 nor n13536 n13537 ; n13538
g13475 and n13535_not n13538 ; n13539
g13476 and n13535 n13538_not ; n13540
g13477 nor n13539 n13540 ; n13541
g13478 and n13524 n13541_not ; n13542
g13479 nor n13525 n13542 ; n13543
g13480 and a[29] n13543_not ; n13544
g13481 and a[29]_not n13543 ; n13545
g13482 nor n13544 n13545 ; n13546
g13483 and n13513 n13546_not ; n13547
g13484 nor n13511 n13547 ; n13548
g13485 nor n13487 n13508 ; n13549
g13486 and n3792 n4788 ; n13550
g13487 and n989 n13550 ; n13551
g13488 and n2371 n13551 ; n13552
g13489 and n3544 n13552 ; n13553
g13490 and n285 n13553 ; n13554
g13491 and n398_not n13554 ; n13555
g13492 and n1062_not n13555 ; n13556
g13493 and n619_not n13556 ; n13557
g13494 and n470_not n13557 ; n13558
g13495 and n271_not n13558 ; n13559
g13496 and n125_not n13559 ; n13560
g13497 and n3549 n5734 ; n13561
g13498 and n12390 n13561 ; n13562
g13499 and n3389 n13562 ; n13563
g13500 and n12939 n13563 ; n13564
g13501 and n13560 n13564 ; n13565
g13502 and n4293 n13565 ; n13566
g13503 and n2021 n13566 ; n13567
g13504 and n896 n13567 ; n13568
g13505 and n3886 n13568 ; n13569
g13506 and n847_not n13569 ; n13570
g13507 and n175_not n13570 ; n13571
g13508 and n286_not n13571 ; n13572
g13509 and n563_not n13572 ; n13573
g13510 and n368_not n13573 ; n13574
g13511 and n13031_not n13574 ; n13575
g13512 and n13031 n13574_not ; n13576
g13513 nor n13549 n13576 ; n13577
g13514 and n13575_not n13577 ; n13578
g13515 nor n13549 n13578 ; n13579
g13516 nor n13575 n13578 ; n13580
g13517 and n13576_not n13580 ; n13581
g13518 nor n13579 n13581 ; n13582
g13519 and n13501 n13529_not ; n13583
g13520 nor n13530 n13583 ; n13584
g13521 and n75 n13584 ; n13585
g13522 and n3020 n13518 ; n13586
g13523 and n3023 n12889 ; n13587
g13524 and n3028 n13491 ; n13588
g13525 nor n13587 n13588 ; n13589
g13526 and n13586_not n13589 ; n13590
g13527 and n13585_not n13590 ; n13591
g13528 nor n13582 n13591 ; n13592
g13529 nor n13582 n13592 ; n13593
g13530 nor n13591 n13592 ; n13594
g13531 nor n13593 n13594 ; n13595
g13532 and n13318_not n13428 ; n13596
g13533 nor n13429 n13596 ; n13597
g13534 and n3457 n13597 ; n13598
g13535 and n3542 n13521 ; n13599
g13536 and n3606 n13515 ; n13600
g13537 nor n13599 n13600 ; n13601
g13538 and n13598_not n13601 ; n13602
g13539 and n3368_not n13602 ; n13603
g13540 nor n13537 n13539 ; n13604
g13541 and n13515 n13597 ; n13605
g13542 nor n13515 n13597 ; n13606
g13543 nor n13604 n13606 ; n13607
g13544 and n13605_not n13607 ; n13608
g13545 nor n13604 n13608 ; n13609
g13546 nor n13605 n13608 ; n13610
g13547 and n13606_not n13610 ; n13611
g13548 nor n13609 n13611 ; n13612
g13549 and n13602 n13612 ; n13613
g13550 nor n13603 n13613 ; n13614
g13551 and a[29] n13614_not ; n13615
g13552 and a[29]_not n13614 ; n13616
g13553 nor n13615 n13616 ; n13617
g13554 nor n13595 n13617 ; n13618
g13555 and n13595 n13617 ; n13619
g13556 nor n13618 n13619 ; n13620
g13557 and n13548_not n13620 ; n13621
g13558 and n13548 n13620_not ; n13622
g13559 nor n13621 n13622 ; n13623
g13560 nor n13434 n13437 ; n13624
g13561 nor n13435 n13437 ; n13625
g13562 and n13083_not n13625 ; n13626
g13563 nor n13624 n13626 ; n13627
g13564 and n3884 n13627_not ; n13628
g13565 and n13190_not n13430 ; n13629
g13566 nor n13431 n13629 ; n13630
g13567 and n3967 n13630 ; n13631
g13568 and n13109 n13432 ; n13632
g13569 nor n13433 n13632 ; n13633
g13570 and n4046 n13633 ; n13634
g13571 nor n13631 n13634 ; n13635
g13572 and n13628_not n13635 ; n13636
g13573 and n13630 n13633 ; n13637
g13574 and n13597 n13630 ; n13638
g13575 nor n13597 n13630 ; n13639
g13576 nor n13638 n13639 ; n13640
g13577 and n13610_not n13640 ; n13641
g13578 nor n13638 n13641 ; n13642
g13579 nor n13630 n13633 ; n13643
g13580 nor n13637 n13643 ; n13644
g13581 and n13642_not n13644 ; n13645
g13582 nor n13637 n13645 ; n13646
g13583 and n13627_not n13633 ; n13647
g13584 and n13627 n13633_not ; n13648
g13585 nor n13646 n13648 ; n13649
g13586 and n13647_not n13649 ; n13650
g13587 nor n13646 n13650 ; n13651
g13588 nor n13647 n13650 ; n13652
g13589 and n13648_not n13652 ; n13653
g13590 nor n13651 n13653 ; n13654
g13591 and n4050 n13654_not ; n13655
g13592 and n13636 n13655_not ; n13656
g13593 and a[26] n13656_not ; n13657
g13594 and a[26] n13657_not ; n13658
g13595 nor n13656 n13657 ; n13659
g13596 nor n13658 n13659 ; n13660
g13597 and n13623 n13660_not ; n13661
g13598 and n13623 n13661_not ; n13662
g13599 nor n13660 n13661 ; n13663
g13600 nor n13662 n13663 ; n13664
g13601 and n13483 n13484_not ; n13665
g13602 nor n12902 n13484 ; n13666
g13603 nor n13665 n13666 ; n13667
g13604 nor n13006 n13008 ; n13668
g13605 and n12997_not n13009 ; n13669
g13606 nor n13668 n13669 ; n13670
g13607 nor n330 n352 ; n13671
g13608 and n1072_not n2809 ; n13672
g13609 and n847_not n13672 ; n13673
g13610 and n557_not n13673 ; n13674
g13611 and n417_not n13674 ; n13675
g13612 and n568_not n13675 ; n13676
g13613 and n205_not n13676 ; n13677
g13614 and n1437 n2220 ; n13678
g13615 and n2487 n13678 ; n13679
g13616 and n2345 n13679 ; n13680
g13617 and n13677 n13680 ; n13681
g13618 and n772 n13681 ; n13682
g13619 and n3108 n13682 ; n13683
g13620 and n5264 n13683 ; n13684
g13621 and n4786 n13684 ; n13685
g13622 and n1824 n13685 ; n13686
g13623 and n2583 n13686 ; n13687
g13624 and n2466 n13687 ; n13688
g13625 and n189_not n13688 ; n13689
g13626 and n13671 n13689 ; n13690
g13627 and n656_not n13690 ; n13691
g13628 and n492_not n13691 ; n13692
g13629 and n201_not n13692 ; n13693
g13630 and n470_not n13693 ; n13694
g13631 and n86_not n13694 ; n13695
g13632 nor n656 n809 ; n13696
g13633 and n145_not n13696 ; n13697
g13634 and n489_not n13697 ; n13698
g13635 and n421 n639_not ; n13699
g13636 and n592_not n13699 ; n13700
g13637 and n2753 n13700 ; n13701
g13638 and n6672 n13701 ; n13702
g13639 and n13138 n13702 ; n13703
g13640 and n13698 n13703 ; n13704
g13641 and n12919 n13704 ; n13705
g13642 and n4815 n13705 ; n13706
g13643 and n2605 n13706 ; n13707
g13644 and n1575 n13707 ; n13708
g13645 and n2406 n13708 ; n13709
g13646 and n202 n13709 ; n13710
g13647 and n1380 n13710 ; n13711
g13648 and n136_not n13711 ; n13712
g13649 and n327_not n13712 ; n13713
g13650 and n393_not n13713 ; n13714
g13651 and n270_not n13714 ; n13715
g13652 nor n13695 n13715 ; n13716
g13653 nor n5939 n6233 ; n13717
g13654 and n5663_not n13717 ; n13718
g13655 and n5666_not n13718 ; n13719
g13656 nor n13438 n13719 ; n13720
g13657 and a[17] n13720_not ; n13721
g13658 and a[17]_not n13720 ; n13722
g13659 nor n13721 n13722 ; n13723
g13660 and n13695 n13715 ; n13724
g13661 nor n13716 n13724 ; n13725
g13662 and n13723 n13725 ; n13726
g13663 nor n13716 n13726 ; n13727
g13664 and n12958 n13727_not ; n13728
g13665 and n12958_not n13727 ; n13729
g13666 nor n13728 n13729 ; n13730
g13667 and n3020 n12502 ; n13731
g13668 and n3028 n12370 ; n13732
g13669 and n3023 n12505 ; n13733
g13670 nor n12680 n12683 ; n13734
g13671 and n12681_not n12684 ; n13735
g13672 nor n13734 n13735 ; n13736
g13673 and n75 n13736_not ; n13737
g13674 nor n13733 n13737 ; n13738
g13675 and n13732_not n13738 ; n13739
g13676 and n13731_not n13739 ; n13740
g13677 and n13730 n13740_not ; n13741
g13678 nor n13728 n13741 ; n13742
g13679 nor n13670 n13742 ; n13743
g13680 and n13670 n13742 ; n13744
g13681 nor n13743 n13744 ; n13745
g13682 nor n12676 n12679 ; n13746
g13683 and n12677_not n12680 ; n13747
g13684 nor n13746 n13747 ; n13748
g13685 and n75 n13748_not ; n13749
g13686 and n3020 n12370 ; n13750
g13687 and n3023 n12508 ; n13751
g13688 and n3028 n12505 ; n13752
g13689 nor n13751 n13752 ; n13753
g13690 and n13750_not n13753 ; n13754
g13691 and n13749_not n13754 ; n13755
g13692 nor n13723 n13725 ; n13756
g13693 nor n13726 n13756 ; n13757
g13694 and n13755_not n13757 ; n13758
g13695 and n1253 n2739 ; n13759
g13696 and n2090 n13759 ; n13760
g13697 and n238 n13760 ; n13761
g13698 and n427_not n13761 ; n13762
g13699 and n335_not n13762 ; n13763
g13700 and n280_not n13763 ; n13764
g13701 and n239_not n13764 ; n13765
g13702 and n460_not n13765 ; n13766
g13703 and n657_not n13766 ; n13767
g13704 and n86_not n13767 ; n13768
g13705 nor n617 n1306 ; n13769
g13706 and n752_not n13769 ; n13770
g13707 and n602_not n13770 ; n13771
g13708 and n286_not n13771 ; n13772
g13709 and n532_not n13772 ; n13773
g13710 nor n130 n144 ; n13774
g13711 and n3160 n13774 ; n13775
g13712 and n13773 n13775 ; n13776
g13713 and n4325 n13776 ; n13777
g13714 and n6020 n13777 ; n13778
g13715 and n1366 n13778 ; n13779
g13716 and n667_not n13779 ; n13780
g13717 and n232_not n13780 ; n13781
g13718 and n495_not n13781 ; n13782
g13719 and n435_not n13782 ; n13783
g13720 and n248_not n13783 ; n13784
g13721 and n91_not n13784 ; n13785
g13722 and n272_not n13785 ; n13786
g13723 and n886_not n13786 ; n13787
g13724 and n2683 n13787 ; n13788
g13725 and n168_not n13788 ; n13789
g13726 and n1308 n13789 ; n13790
g13727 and n1942 n13790 ; n13791
g13728 and n5791 n13791 ; n13792
g13729 and n2796 n13792 ; n13793
g13730 and n13768 n13793 ; n13794
g13731 and n1575 n13794 ; n13795
g13732 and n2484 n13795 ; n13796
g13733 and n159 n13796 ; n13797
g13734 and n1161 n13797 ; n13798
g13735 and n229_not n13798 ; n13799
g13736 and n329_not n13799 ; n13800
g13737 and n353_not n13800 ; n13801
g13738 and n639_not n13801 ; n13802
g13739 and n567_not n13802 ; n13803
g13740 and n712_not n13803 ; n13804
g13741 and n304_not n13804 ; n13805
g13742 and n13695 n13805_not ; n13806
g13743 and n136_not n5082 ; n13807
g13744 and n884_not n13807 ; n13808
g13745 and n5271 n13808 ; n13809
g13746 and n3041 n13809 ; n13810
g13747 and n2716 n13810 ; n13811
g13748 and n3489 n13811 ; n13812
g13749 and n4367 n13812 ; n13813
g13750 and n1080 n13813 ; n13814
g13751 and n518_not n13814 ; n13815
g13752 and n602_not n13815 ; n13816
g13753 and n146_not n13816 ; n13817
g13754 and n888 n13817 ; n13818
g13755 and n673_not n13818 ; n13819
g13756 and n564_not n13819 ; n13820
g13757 and n125_not n13820 ; n13821
g13758 and n423 n1366 ; n13822
g13759 and n151_not n13822 ; n13823
g13760 and n537_not n13823 ; n13824
g13761 and n375_not n13824 ; n13825
g13762 and n222_not n13825 ; n13826
g13763 and n773 n1528 ; n13827
g13764 and n1346 n13827 ; n13828
g13765 and n4298 n13828 ; n13829
g13766 and n3068 n13829 ; n13830
g13767 and n434 n13830 ; n13831
g13768 and n13826 n13831 ; n13832
g13769 and n1814 n13832 ; n13833
g13770 and n6514 n13833 ; n13834
g13771 and n774 n13834 ; n13835
g13772 and n1838 n13835 ; n13836
g13773 and n232_not n13836 ; n13837
g13774 and n637_not n13837 ; n13838
g13775 and n228_not n13838 ; n13839
g13776 and n302_not n13839 ; n13840
g13777 and n298_not n13840 ; n13841
g13778 and n295_not n13841 ; n13842
g13779 and n127_not n13842 ; n13843
g13780 nor n13821 n13843 ; n13844
g13781 nor n6951 n7101 ; n13845
g13782 and n6402_not n13845 ; n13846
g13783 and n6397_not n13846 ; n13847
g13784 nor n13438 n13847 ; n13848
g13785 and a[14] n13848_not ; n13849
g13786 and a[14]_not n13848 ; n13850
g13787 nor n13849 n13850 ; n13851
g13788 and n13821 n13843 ; n13852
g13789 nor n13844 n13852 ; n13853
g13790 and n13851 n13853 ; n13854
g13791 nor n13844 n13854 ; n13855
g13792 and n13805 n13855_not ; n13856
g13793 and n13805_not n13855 ; n13857
g13794 nor n13856 n13857 ; n13858
g13795 and n3020 n12508 ; n13859
g13796 and n3028 n12513 ; n13860
g13797 and n3023 n12511 ; n13861
g13798 and n12667 n12670_not ; n13862
g13799 nor n12671 n13862 ; n13863
g13800 and n75 n13863 ; n13864
g13801 nor n13861 n13864 ; n13865
g13802 and n13860_not n13865 ; n13866
g13803 and n13859_not n13866 ; n13867
g13804 and n13858 n13867_not ; n13868
g13805 nor n13856 n13868 ; n13869
g13806 and n13695_not n13805 ; n13870
g13807 nor n13869 n13870 ; n13871
g13808 and n13806_not n13871 ; n13872
g13809 nor n13806 n13872 ; n13873
g13810 and n13757 n13758_not ; n13874
g13811 nor n13755 n13758 ; n13875
g13812 nor n13874 n13875 ; n13876
g13813 nor n13873 n13876 ; n13877
g13814 nor n13758 n13877 ; n13878
g13815 and n13730_not n13740 ; n13879
g13816 nor n13741 n13879 ; n13880
g13817 and n13878_not n13880 ; n13881
g13818 and n13878 n13880_not ; n13882
g13819 nor n13881 n13882 ; n13883
g13820 and n3457 n13491 ; n13884
g13821 and n3542 n12769 ; n13885
g13822 and n3606 n12889 ; n13886
g13823 nor n13885 n13886 ; n13887
g13824 and n13884_not n13887 ; n13888
g13825 and n3368_not n13888 ; n13889
g13826 and n13503 n13888 ; n13890
g13827 nor n13889 n13890 ; n13891
g13828 and a[29] n13891_not ; n13892
g13829 and a[29]_not n13891 ; n13893
g13830 nor n13892 n13893 ; n13894
g13831 and n13883 n13894_not ; n13895
g13832 nor n13881 n13895 ; n13896
g13833 and n13745 n13896_not ; n13897
g13834 nor n13743 n13897 ; n13898
g13835 nor n13667 n13898 ; n13899
g13836 and n13667 n13898 ; n13900
g13837 nor n13899 n13900 ; n13901
g13838 and n3457 n13521 ; n13902
g13839 and n3542 n13491 ; n13903
g13840 and n3606 n13518 ; n13904
g13841 nor n13903 n13904 ; n13905
g13842 and n13902_not n13905 ; n13906
g13843 nor n13531 n13534 ; n13907
g13844 and n13532_not n13535 ; n13908
g13845 nor n13907 n13908 ; n13909
g13846 and n3368 n13909_not ; n13910
g13847 and n13906 n13910_not ; n13911
g13848 and a[29] n13911_not ; n13912
g13849 and a[29] n13912_not ; n13913
g13850 nor n13911 n13912 ; n13914
g13851 nor n13913 n13914 ; n13915
g13852 and n13901 n13915_not ; n13916
g13853 nor n13899 n13916 ; n13917
g13854 and n13513_not n13546 ; n13918
g13855 nor n13547 n13918 ; n13919
g13856 and n13917_not n13919 ; n13920
g13857 and n13917 n13919_not ; n13921
g13858 nor n13920 n13921 ; n13922
g13859 and n3884 n13633 ; n13923
g13860 and n3967 n13597 ; n13924
g13861 and n4046 n13630 ; n13925
g13862 nor n13924 n13925 ; n13926
g13863 and n13923_not n13926 ; n13927
g13864 and n13642 n13644_not ; n13928
g13865 nor n13645 n13928 ; n13929
g13866 and n4050 n13929 ; n13930
g13867 and n13927 n13930_not ; n13931
g13868 and a[26] n13931_not ; n13932
g13869 and a[26] n13932_not ; n13933
g13870 nor n13931 n13932 ; n13934
g13871 nor n13933 n13934 ; n13935
g13872 and n13922 n13935_not ; n13936
g13873 nor n13920 n13936 ; n13937
g13874 nor n4604 n4694 ; n13938
g13875 nor n13438 n13938 ; n13939
g13876 and n13059 n13625 ; n13940
g13877 nor n13438 n13940 ; n13941
g13878 and n4533 n13941 ; n13942
g13879 nor n13939 n13942 ; n13943
g13880 and n4536_not n13943 ; n13944
g13881 and n13627_not n13941 ; n13945
g13882 and n13627 n13941_not ; n13946
g13883 nor n13945 n13946 ; n13947
g13884 and n13652_not n13947 ; n13948
g13885 nor n13945 n13948 ; n13949
g13886 and n13940 n13949_not ; n13950
g13887 nor n13941 n13950 ; n13951
g13888 and n13943 n13951 ; n13952
g13889 nor n13944 n13952 ; n13953
g13890 and a[23] n13953_not ; n13954
g13891 and a[23]_not n13953 ; n13955
g13892 nor n13954 n13955 ; n13956
g13893 nor n13937 n13956 ; n13957
g13894 and n13937 n13956 ; n13958
g13895 nor n13957 n13958 ; n13959
g13896 and n13664_not n13959 ; n13960
g13897 nor n13664 n13960 ; n13961
g13898 and n13959 n13960_not ; n13962
g13899 nor n13961 n13962 ; n13963
g13900 and n13922 n13936_not ; n13964
g13901 nor n13935 n13936 ; n13965
g13902 nor n13964 n13965 ; n13966
g13903 and n13901 n13916_not ; n13967
g13904 nor n13915 n13916 ; n13968
g13905 nor n13967 n13968 ; n13969
g13906 and n3884 n13630 ; n13970
g13907 and n3967 n13515 ; n13971
g13908 and n4046 n13597 ; n13972
g13909 nor n13971 n13972 ; n13973
g13910 and n13970_not n13973 ; n13974
g13911 and n13610 n13640_not ; n13975
g13912 nor n13641 n13975 ; n13976
g13913 and n4050 n13976 ; n13977
g13914 and n13974 n13977_not ; n13978
g13915 and a[26] n13978_not ; n13979
g13916 and a[26] n13979_not ; n13980
g13917 nor n13978 n13979 ; n13981
g13918 nor n13980 n13981 ; n13982
g13919 nor n13969 n13982 ; n13983
g13920 nor n13969 n13983 ; n13984
g13921 nor n13982 n13983 ; n13985
g13922 nor n13984 n13985 ; n13986
g13923 and n13745_not n13896 ; n13987
g13924 nor n13897 n13987 ; n13988
g13925 and n3457 n13518 ; n13989
g13926 and n3542 n12889 ; n13990
g13927 and n3606 n13491 ; n13991
g13928 nor n13990 n13991 ; n13992
g13929 and n13989_not n13992 ; n13993
g13930 and n3368 n13584 ; n13994
g13931 and n13993 n13994_not ; n13995
g13932 and a[29] n13995_not ; n13996
g13933 and a[29] n13996_not ; n13997
g13934 nor n13995 n13996 ; n13998
g13935 nor n13997 n13998 ; n13999
g13936 and n13988 n13999_not ; n14000
g13937 and n13988 n14000_not ; n14001
g13938 nor n13999 n14000 ; n14002
g13939 nor n14001 n14002 ; n14003
g13940 and n3884 n13597 ; n14004
g13941 and n3967 n13521 ; n14005
g13942 and n4046 n13515 ; n14006
g13943 nor n14005 n14006 ; n14007
g13944 and n14004_not n14007 ; n14008
g13945 and n4050 n13612_not ; n14009
g13946 and n14008 n14009_not ; n14010
g13947 and a[26] n14010_not ; n14011
g13948 and a[26] n14011_not ; n14012
g13949 nor n14010 n14011 ; n14013
g13950 nor n14012 n14013 ; n14014
g13951 nor n14003 n14014 ; n14015
g13952 nor n14000 n14015 ; n14016
g13953 nor n13986 n14016 ; n14017
g13954 nor n13983 n14017 ; n14018
g13955 nor n13966 n14018 ; n14019
g13956 and n13966 n14018 ; n14020
g13957 nor n14019 n14020 ; n14021
g13958 and n4694 n13438_not ; n14022
g13959 and n4533 n13627_not ; n14023
g13960 and n4604 n13941 ; n14024
g13961 nor n14023 n14024 ; n14025
g13962 and n14022_not n14025 ; n14026
g13963 and n13940_not n13949 ; n14027
g13964 nor n13950 n14027 ; n14028
g13965 and n4536 n14028 ; n14029
g13966 and n14026 n14029_not ; n14030
g13967 and a[23] n14030_not ; n14031
g13968 and a[23] n14031_not ; n14032
g13969 nor n14030 n14031 ; n14033
g13970 nor n14032 n14033 ; n14034
g13971 and n14021 n14034_not ; n14035
g13972 nor n14019 n14035 ; n14036
g13973 nor n13963 n14036 ; n14037
g13974 and n13963 n14036 ; n14038
g13975 nor n14037 n14038 ; n14039
g13976 and n14021 n14035_not ; n14040
g13977 nor n14034 n14035 ; n14041
g13978 nor n14040 n14041 ; n14042
g13979 nor n14003 n14015 ; n14043
g13980 nor n14014 n14015 ; n14044
g13981 nor n14043 n14044 ; n14045
g13982 nor n13869 n13872 ; n14046
g13983 and n13870_not n13873 ; n14047
g13984 nor n14046 n14047 ; n14048
g13985 nor n12672 n12675 ; n14049
g13986 and n12673_not n12676 ; n14050
g13987 nor n14049 n14050 ; n14051
g13988 and n75 n14051_not ; n14052
g13989 and n3020 n12505 ; n14053
g13990 and n3023 n12513 ; n14054
g13991 and n3028 n12508 ; n14055
g13992 nor n14054 n14055 ; n14056
g13993 and n14053_not n14056 ; n14057
g13994 and n14052_not n14057 ; n14058
g13995 nor n14048 n14058 ; n14059
g13996 nor n14048 n14059 ; n14060
g13997 nor n14058 n14059 ; n14061
g13998 nor n14060 n14061 ; n14062
g13999 and n3457 n12769 ; n14063
g14000 and n3542 n12370 ; n14064
g14001 and n3606 n12502 ; n14065
g14002 nor n14064 n14065 ; n14066
g14003 and n14063_not n14066 ; n14067
g14004 and n3368_not n14067 ; n14068
g14005 and n12999_not n14067 ; n14069
g14006 nor n14068 n14069 ; n14070
g14007 and a[29] n14070_not ; n14071
g14008 and a[29]_not n14070 ; n14072
g14009 nor n14071 n14072 ; n14073
g14010 nor n14062 n14073 ; n14074
g14011 nor n14059 n14074 ; n14075
g14012 nor n13876 n13877 ; n14076
g14013 nor n13873 n13877 ; n14077
g14014 nor n14076 n14077 ; n14078
g14015 nor n14075 n14078 ; n14079
g14016 nor n14075 n14079 ; n14080
g14017 nor n14078 n14079 ; n14081
g14018 nor n14080 n14081 ; n14082
g14019 and n3457 n12889 ; n14083
g14020 and n3542 n12502 ; n14084
g14021 and n3606 n12769 ; n14085
g14022 nor n14084 n14085 ; n14086
g14023 and n14083_not n14086 ; n14087
g14024 and n3368 n12895 ; n14088
g14025 and n14087 n14088_not ; n14089
g14026 and a[29] n14089_not ; n14090
g14027 and a[29] n14090_not ; n14091
g14028 nor n14089 n14090 ; n14092
g14029 nor n14091 n14092 ; n14093
g14030 nor n14082 n14093 ; n14094
g14031 nor n14079 n14094 ; n14095
g14032 and n13883_not n13894 ; n14096
g14033 nor n13895 n14096 ; n14097
g14034 and n14095_not n14097 ; n14098
g14035 and n14095 n14097_not ; n14099
g14036 nor n14098 n14099 ; n14100
g14037 and n3884 n13515 ; n14101
g14038 and n3967 n13518 ; n14102
g14039 and n4046 n13521 ; n14103
g14040 nor n14102 n14103 ; n14104
g14041 and n14101_not n14104 ; n14105
g14042 and n4050 n13541 ; n14106
g14043 and n14105 n14106_not ; n14107
g14044 and a[26] n14107_not ; n14108
g14045 and a[26] n14108_not ; n14109
g14046 nor n14107 n14108 ; n14110
g14047 nor n14109 n14110 ; n14111
g14048 and n14100 n14111_not ; n14112
g14049 nor n14098 n14112 ; n14113
g14050 nor n14045 n14113 ; n14114
g14051 and n14045 n14113 ; n14115
g14052 nor n14114 n14115 ; n14116
g14053 and n4694 n13627_not ; n14117
g14054 and n4533 n13630 ; n14118
g14055 and n4604 n13633 ; n14119
g14056 nor n14118 n14119 ; n14120
g14057 and n14117_not n14120 ; n14121
g14058 and n4536 n13654_not ; n14122
g14059 and n14121 n14122_not ; n14123
g14060 and a[23] n14123_not ; n14124
g14061 and a[23] n14124_not ; n14125
g14062 nor n14123 n14124 ; n14126
g14063 nor n14125 n14126 ; n14127
g14064 and n14116 n14127_not ; n14128
g14065 nor n14114 n14128 ; n14129
g14066 and n4694 n13941 ; n14130
g14067 and n4533 n13633 ; n14131
g14068 and n4604 n13627_not ; n14132
g14069 nor n14131 n14132 ; n14133
g14070 and n14130_not n14133 ; n14134
g14071 and n13652 n13947_not ; n14135
g14072 nor n13948 n14135 ; n14136
g14073 and n4536 n14136 ; n14137
g14074 and n14134 n14137_not ; n14138
g14075 and a[23] n14138_not ; n14139
g14076 and a[23] n14139_not ; n14140
g14077 nor n14138 n14139 ; n14141
g14078 nor n14140 n14141 ; n14142
g14079 nor n14129 n14142 ; n14143
g14080 and n13986 n14016 ; n14144
g14081 nor n14017 n14144 ; n14145
g14082 nor n14129 n14143 ; n14146
g14083 nor n14142 n14143 ; n14147
g14084 nor n14146 n14147 ; n14148
g14085 and n14145 n14148_not ; n14149
g14086 nor n14143 n14149 ; n14150
g14087 nor n14042 n14150 ; n14151
g14088 nor n14042 n14151 ; n14152
g14089 nor n14150 n14151 ; n14153
g14090 nor n14152 n14153 ; n14154
g14091 and n14100 n14112_not ; n14155
g14092 nor n14111 n14112 ; n14156
g14093 nor n14155 n14156 ; n14157
g14094 nor n14082 n14094 ; n14158
g14095 nor n14093 n14094 ; n14159
g14096 nor n14158 n14159 ; n14160
g14097 and n3884 n13521 ; n14161
g14098 and n3967 n13491 ; n14162
g14099 and n4046 n13518 ; n14163
g14100 nor n14162 n14163 ; n14164
g14101 and n14161_not n14164 ; n14165
g14102 and n4050 n13909_not ; n14166
g14103 and n14165 n14166_not ; n14167
g14104 and a[26] n14167_not ; n14168
g14105 and a[26] n14168_not ; n14169
g14106 nor n14167 n14168 ; n14170
g14107 nor n14169 n14170 ; n14171
g14108 nor n14160 n14171 ; n14172
g14109 nor n14160 n14172 ; n14173
g14110 nor n14171 n14172 ; n14174
g14111 nor n14173 n14174 ; n14175
g14112 and n12663 n12665_not ; n14176
g14113 nor n12666 n14176 ; n14177
g14114 and n75 n14177 ; n14178
g14115 and n3020 n12513 ; n14179
g14116 and n3023 n12516 ; n14180
g14117 and n3028 n12511 ; n14181
g14118 nor n14180 n14181 ; n14182
g14119 and n14179_not n14182 ; n14183
g14120 and n14178_not n14183 ; n14184
g14121 nor n142 n506 ; n14185
g14122 and n422_not n14185 ; n14186
g14123 and n603_not n14186 ; n14187
g14124 and n130_not n14187 ; n14188
g14125 and n332_not n14188 ; n14189
g14126 and n1109 n3523 ; n14190
g14127 and n5777 n14190 ; n14191
g14128 and n14189 n14191 ; n14192
g14129 and n2022 n14192 ; n14193
g14130 and n622 n14193 ; n14194
g14131 and n874 n14194 ; n14195
g14132 and n774 n14195 ; n14196
g14133 and n872 n14196 ; n14197
g14134 and n356 n14197 ; n14198
g14135 and n1306_not n14198 ; n14199
g14136 and n403_not n14199 ; n14200
g14137 and n161_not n14200 ; n14201
g14138 and n655_not n14201 ; n14202
g14139 and n642 n3165 ; n14203
g14140 and n2390 n14203 ; n14204
g14141 and n989 n14204 ; n14205
g14142 and n1782 n14205 ; n14206
g14143 and n1011_not n14206 ; n14207
g14144 and n847_not n14207 ; n14208
g14145 and n331_not n14208 ; n14209
g14146 and n132_not n14209 ; n14210
g14147 and n529 n14210 ; n14211
g14148 and n3681 n14211 ; n14212
g14149 and n2296 n14212 ; n14213
g14150 and n14202 n14213 ; n14214
g14151 and n1046 n14214 ; n14215
g14152 and n450 n14215 ; n14216
g14153 and n937 n14216 ; n14217
g14154 and n2088 n14217 ; n14218
g14155 and n4101 n14218 ; n14219
g14156 and n1522 n14219 ; n14220
g14157 and n136_not n14220 ; n14221
g14158 and n1062_not n14221 ; n14222
g14159 and n302_not n14222 ; n14223
g14160 and n192_not n14223 ; n14224
g14161 and n430_not n14224 ; n14225
g14162 and n201_not n14225 ; n14226
g14163 and n657_not n14226 ; n14227
g14164 and n158_not n14227 ; n14228
g14165 and n13821 n14228_not ; n14229
g14166 and n13821_not n14228 ; n14230
g14167 nor n12659 n12662 ; n14231
g14168 and n12660_not n12663 ; n14232
g14169 nor n14231 n14232 ; n14233
g14170 and n75 n14233_not ; n14234
g14171 and n3020 n12511 ; n14235
g14172 and n3023 n12519 ; n14236
g14173 and n3028 n12516 ; n14237
g14174 nor n14236 n14237 ; n14238
g14175 and n14235_not n14238 ; n14239
g14176 and n14234_not n14239 ; n14240
g14177 nor n14229 n14240 ; n14241
g14178 and n14230_not n14241 ; n14242
g14179 nor n14229 n14242 ; n14243
g14180 nor n13851 n13853 ; n14244
g14181 nor n13854 n14244 ; n14245
g14182 and n14243_not n14245 ; n14246
g14183 and n14243 n14245_not ; n14247
g14184 nor n14246 n14247 ; n14248
g14185 and n14184_not n14248 ; n14249
g14186 nor n14246 n14249 ; n14250
g14187 and n13858_not n13867 ; n14251
g14188 nor n13868 n14251 ; n14252
g14189 and n14250_not n14252 ; n14253
g14190 and n14250 n14252_not ; n14254
g14191 nor n14253 n14254 ; n14255
g14192 and n3457 n12502 ; n14256
g14193 and n3542 n12505 ; n14257
g14194 and n3606 n12370 ; n14258
g14195 nor n14257 n14258 ; n14259
g14196 and n14256_not n14259 ; n14260
g14197 and n3368_not n14260 ; n14261
g14198 and n13736 n14260 ; n14262
g14199 nor n14261 n14262 ; n14263
g14200 and a[29] n14263_not ; n14264
g14201 and a[29]_not n14263 ; n14265
g14202 nor n14264 n14265 ; n14266
g14203 and n14255 n14266_not ; n14267
g14204 nor n14253 n14267 ; n14268
g14205 and n14062 n14073 ; n14269
g14206 nor n14074 n14269 ; n14270
g14207 and n14268_not n14270 ; n14271
g14208 and n14268 n14270_not ; n14272
g14209 nor n14271 n14272 ; n14273
g14210 and n3884 n13518 ; n14274
g14211 and n3967 n12889 ; n14275
g14212 and n4046 n13491 ; n14276
g14213 nor n14275 n14276 ; n14277
g14214 and n14274_not n14277 ; n14278
g14215 and n4050 n13584 ; n14279
g14216 and n14278 n14279_not ; n14280
g14217 and a[26] n14280_not ; n14281
g14218 and a[26] n14281_not ; n14282
g14219 nor n14280 n14281 ; n14283
g14220 nor n14282 n14283 ; n14284
g14221 and n14273 n14284_not ; n14285
g14222 nor n14271 n14285 ; n14286
g14223 nor n14175 n14286 ; n14287
g14224 nor n14172 n14287 ; n14288
g14225 nor n14157 n14288 ; n14289
g14226 and n14157 n14288 ; n14290
g14227 nor n14289 n14290 ; n14291
g14228 and n4694 n13633 ; n14292
g14229 and n4533 n13597 ; n14293
g14230 and n4604 n13630 ; n14294
g14231 nor n14293 n14294 ; n14295
g14232 and n14292_not n14295 ; n14296
g14233 and n4536 n13929 ; n14297
g14234 and n14296 n14297_not ; n14298
g14235 and a[23] n14298_not ; n14299
g14236 and a[23] n14299_not ; n14300
g14237 nor n14298 n14299 ; n14301
g14238 nor n14300 n14301 ; n14302
g14239 and n14291 n14302_not ; n14303
g14240 nor n14289 n14303 ; n14304
g14241 nor n13438 n13439 ; n14305
g14242 and n4935 n13941 ; n14306
g14243 nor n14305 n14306 ; n14307
g14244 and n4938_not n14307 ; n14308
g14245 and n13951 n14307 ; n14309
g14246 nor n14308 n14309 ; n14310
g14247 and a[20] n14310_not ; n14311
g14248 and a[20]_not n14310 ; n14312
g14249 nor n14311 n14312 ; n14313
g14250 nor n14304 n14313 ; n14314
g14251 and n14116 n14128_not ; n14315
g14252 nor n14127 n14128 ; n14316
g14253 nor n14315 n14316 ; n14317
g14254 and n14304 n14313 ; n14318
g14255 nor n14314 n14318 ; n14319
g14256 and n14317_not n14319 ; n14320
g14257 nor n14314 n14320 ; n14321
g14258 and n14145_not n14148 ; n14322
g14259 nor n14149 n14322 ; n14323
g14260 and n14321_not n14323 ; n14324
g14261 nor n14317 n14320 ; n14325
g14262 and n14319 n14320_not ; n14326
g14263 nor n14325 n14326 ; n14327
g14264 and n14291 n14303_not ; n14328
g14265 nor n14302 n14303 ; n14329
g14266 nor n14328 n14329 ; n14330
g14267 and n14175 n14286 ; n14331
g14268 nor n14287 n14331 ; n14332
g14269 and n4694 n13630 ; n14333
g14270 and n4533 n13515 ; n14334
g14271 and n4604 n13597 ; n14335
g14272 nor n14334 n14335 ; n14336
g14273 and n14333_not n14336 ; n14337
g14274 and n4536 n13976 ; n14338
g14275 and n14337 n14338_not ; n14339
g14276 and a[23] n14339_not ; n14340
g14277 and a[23] n14340_not ; n14341
g14278 nor n14339 n14340 ; n14342
g14279 nor n14341 n14342 ; n14343
g14280 and n14332 n14343_not ; n14344
g14281 and n14332 n14344_not ; n14345
g14282 nor n14343 n14344 ; n14346
g14283 nor n14345 n14346 ; n14347
g14284 and n14273 n14285_not ; n14348
g14285 nor n14284 n14285 ; n14349
g14286 nor n14348 n14349 ; n14350
g14287 and n14248 n14249_not ; n14351
g14288 nor n14184 n14249 ; n14352
g14289 nor n14351 n14352 ; n14353
g14290 and n3457 n12370 ; n14354
g14291 and n3542 n12508 ; n14355
g14292 and n3606 n12505 ; n14356
g14293 nor n14355 n14356 ; n14357
g14294 and n14354_not n14357 ; n14358
g14295 and n3368 n13748_not ; n14359
g14296 and n14358 n14359_not ; n14360
g14297 and a[29] n14360_not ; n14361
g14298 and a[29] n14361_not ; n14362
g14299 nor n14360 n14361 ; n14363
g14300 nor n14362 n14363 ; n14364
g14301 nor n14353 n14364 ; n14365
g14302 nor n14353 n14365 ; n14366
g14303 nor n14364 n14365 ; n14367
g14304 nor n14366 n14367 ; n14368
g14305 nor n14240 n14242 ; n14369
g14306 and n14230_not n14243 ; n14370
g14307 nor n14369 n14370 ; n14371
g14308 and n1271 n1602 ; n14372
g14309 and n2698 n14372 ; n14373
g14310 and n123_not n14373 ; n14374
g14311 and n557_not n14374 ; n14375
g14312 and n571_not n14375 ; n14376
g14313 and n513_not n14376 ; n14377
g14314 and n490_not n14377 ; n14378
g14315 and n302_not n14378 ; n14379
g14316 and n191_not n14379 ; n14380
g14317 and n372_not n14380 ; n14381
g14318 and n278_not n5064 ; n14382
g14319 and n248_not n14382 ; n14383
g14320 and n403_not n14383 ; n14384
g14321 and n164_not n14384 ; n14385
g14322 and n366_not n14385 ; n14386
g14323 and n1996 n13114 ; n14387
g14324 and n4130 n14387 ; n14388
g14325 and n2022 n14388 ; n14389
g14326 and n14386 n14389 ; n14390
g14327 and n2772 n14390 ; n14391
g14328 and n6097 n14391 ; n14392
g14329 and n14381 n14392 ; n14393
g14330 and n2583 n14393 ; n14394
g14331 and n1367 n14394 ; n14395
g14332 and n1389 n14395 ; n14396
g14333 and n420_not n14396 ; n14397
g14334 and n281_not n14397 ; n14398
g14335 and n4294 n14398 ; n14399
g14336 and n393_not n14399 ; n14400
g14337 and n272_not n14400 ; n14401
g14338 and n672_not n14401 ; n14402
g14339 and n371_not n14402 ; n14403
g14340 and n1140 n2210 ; n14404
g14341 and n619_not n14404 ; n14405
g14342 and n157_not n14405 ; n14406
g14343 and n125_not n14406 ; n14407
g14344 and n889 n2363 ; n14408
g14345 and n2544 n14408 ; n14409
g14346 and n1085 n14409 ; n14410
g14347 and n5746 n14410 ; n14411
g14348 and n1119 n14411 ; n14412
g14349 and n268 n14412 ; n14413
g14350 and n3405 n14413 ; n14414
g14351 and n3472 n14414 ; n14415
g14352 and n14407 n14415 ; n14416
g14353 and n933 n14416 ; n14417
g14354 and n4295 n14417 ; n14418
g14355 and n168_not n14418 ; n14419
g14356 and n400_not n14419 ; n14420
g14357 and n206_not n14420 ; n14421
g14358 and n145_not n14421 ; n14422
g14359 nor n14403 n14422 ; n14423
g14360 nor n7632 n7983 ; n14424
g14361 and n7291_not n14424 ; n14425
g14362 and n7294_not n14425 ; n14426
g14363 nor n13438 n14426 ; n14427
g14364 and a[11] n14427_not ; n14428
g14365 and a[11]_not n14427 ; n14429
g14366 nor n14428 n14429 ; n14430
g14367 and n14403 n14422 ; n14431
g14368 nor n14423 n14431 ; n14432
g14369 and n14430 n14432 ; n14433
g14370 nor n14423 n14433 ; n14434
g14371 and n13821 n14434_not ; n14435
g14372 and n13821_not n14434 ; n14436
g14373 nor n14435 n14436 ; n14437
g14374 and n3020 n12516 ; n14438
g14375 and n3028 n12519 ; n14439
g14376 and n3023 n12522 ; n14440
g14377 nor n12655 n12658 ; n14441
g14378 and n12656_not n12659 ; n14442
g14379 nor n14441 n14442 ; n14443
g14380 and n75 n14443_not ; n14444
g14381 nor n14440 n14444 ; n14445
g14382 and n14439_not n14445 ; n14446
g14383 and n14438_not n14446 ; n14447
g14384 and n14437 n14447_not ; n14448
g14385 nor n14435 n14448 ; n14449
g14386 nor n14371 n14449 ; n14450
g14387 and n14371 n14449 ; n14451
g14388 nor n14450 n14451 ; n14452
g14389 and n12651 n12653_not ; n14453
g14390 nor n12654 n14453 ; n14454
g14391 and n75 n14454 ; n14455
g14392 and n3020 n12519 ; n14456
g14393 and n3023 n12525 ; n14457
g14394 and n3028 n12522 ; n14458
g14395 nor n14457 n14458 ; n14459
g14396 and n14456_not n14459 ; n14460
g14397 and n14455_not n14460 ; n14461
g14398 nor n14430 n14432 ; n14462
g14399 nor n14433 n14462 ; n14463
g14400 and n14461_not n14463 ; n14464
g14401 and n14463 n14464_not ; n14465
g14402 nor n14461 n14464 ; n14466
g14403 nor n14465 n14466 ; n14467
g14404 and n1204 n2154 ; n14468
g14405 and n665 n14468 ; n14469
g14406 and n617_not n14469 ; n14470
g14407 and n169_not n14470 ; n14471
g14408 and n667_not n14471 ; n14472
g14409 and n402_not n14472 ; n14473
g14410 and n490_not n14473 ; n14474
g14411 and n374_not n14474 ; n14475
g14412 and n132_not n14475 ; n14476
g14413 nor n601 n1101 ; n14477
g14414 and n251_not n14477 ; n14478
g14415 and n270_not n14478 ; n14479
g14416 and n510 n809_not ; n14480
g14417 and n568_not n14480 ; n14481
g14418 and n424_not n14481 ; n14482
g14419 and n1425 n3549 ; n14483
g14420 and n2653 n14483 ; n14484
g14421 and n14482 n14484 ; n14485
g14422 and n198 n14485 ; n14486
g14423 and n1940 n14486 ; n14487
g14424 and n14479 n14487 ; n14488
g14425 and n1292 n14488 ; n14489
g14426 and n1330 n14489 ; n14490
g14427 and n827 n14490 ; n14491
g14428 and n1380 n14491 ; n14492
g14429 and n1269 n14492 ; n14493
g14430 and n397_not n14493 ; n14494
g14431 and n1246_not n14494 ; n14495
g14432 and n278_not n14495 ; n14496
g14433 and n95_not n14496 ; n14497
g14434 and n125_not n14497 ; n14498
g14435 and n674 n1646 ; n14499
g14436 and n3985 n14499 ; n14500
g14437 and n207 n14500 ; n14501
g14438 and n14498 n14501 ; n14502
g14439 and n4247 n14502 ; n14503
g14440 and n14476 n14503 ; n14504
g14441 and n622 n14504 ; n14505
g14442 and n2739 n14505 ; n14506
g14443 and n159 n14506 ; n14507
g14444 and n356 n14507 ; n14508
g14445 and n229_not n14508 ; n14509
g14446 and n620_not n14509 ; n14510
g14447 and n248_not n14510 ; n14511
g14448 and n416_not n14511 ; n14512
g14449 and n237_not n14512 ; n14513
g14450 and n119_not n14513 ; n14514
g14451 and n14403 n14514_not ; n14515
g14452 and n14403_not n14514 ; n14516
g14453 and n118_not n454 ; n14517
g14454 and n165_not n14517 ; n14518
g14455 and n2348 n14518 ; n14519
g14456 and n1576 n14519 ; n14520
g14457 and n571_not n14520 ; n14521
g14458 and n594_not n14521 ; n14522
g14459 and n132_not n14522 ; n14523
g14460 and n1010_not n14523 ; n14524
g14461 and n270_not n14524 ; n14525
g14462 and n343 n13700 ; n14526
g14463 and n1070 n14526 ; n14527
g14464 and n3409 n14527 ; n14528
g14465 and n1062_not n14528 ; n14529
g14466 and n809_not n14529 ; n14530
g14467 and n331_not n14530 ; n14531
g14468 and n689_not n14531 ; n14532
g14469 and n673_not n14532 ; n14533
g14470 and n474_not n14533 ; n14534
g14471 and n497 n1315 ; n14535
g14472 and n4132 n14535 ; n14536
g14473 and n2192 n14536 ; n14537
g14474 and n450 n14537 ; n14538
g14475 and n227 n14538 ; n14539
g14476 and n803_not n14539 ; n14540
g14477 and n435_not n14540 ; n14541
g14478 and n461_not n14541 ; n14542
g14479 and n306_not n14542 ; n14543
g14480 and n237_not n14543 ; n14544
g14481 and n2026 n2995 ; n14545
g14482 and n3512 n14545 ; n14546
g14483 and n2317 n14546 ; n14547
g14484 and n3113 n14547 ; n14548
g14485 and n14544 n14548 ; n14549
g14486 and n14534 n14549 ; n14550
g14487 and n14525 n14550 ; n14551
g14488 and n2633 n14551 ; n14552
g14489 and n2443 n14552 ; n14553
g14490 and n720 n14553 ; n14554
g14491 and n356 n14554 ; n14555
g14492 and n1180 n14555 ; n14556
g14493 and n194_not n14556 ; n14557
g14494 and n334_not n14557 ; n14558
g14495 and n125_not n14558 ; n14559
g14496 nor n594 n716 ; n14560
g14497 and n331_not n14560 ; n14561
g14498 and n1246_not n14561 ; n14562
g14499 and n289_not n14562 ; n14563
g14500 and n527_not n14563 ; n14564
g14501 and n201_not n14564 ; n14565
g14502 and n1695 n2012 ; n14566
g14503 and n1602 n14566 ; n14567
g14504 and n810 n14567 ; n14568
g14505 and n151_not n14568 ; n14569
g14506 and n286_not n14569 ; n14570
g14507 and n496_not n14570 ; n14571
g14508 and n272_not n14571 ; n14572
g14509 and n1896 n2293 ; n14573
g14510 and n693 n14573 ; n14574
g14511 and n5036 n14574 ; n14575
g14512 and n1692 n14575 ; n14576
g14513 and n13265 n14576 ; n14577
g14514 and n14572 n14577 ; n14578
g14515 and n1100 n14578 ; n14579
g14516 and n120 n14579 ; n14580
g14517 and n14565 n14580 ; n14581
g14518 and n359 n14581 ; n14582
g14519 and n427_not n14582 ; n14583
g14520 and n397_not n14583 ; n14584
g14521 and n206_not n14584 ; n14585
g14522 and n505_not n14585 ; n14586
g14523 and n170_not n14586 ; n14587
g14524 and n493_not n14587 ; n14588
g14525 nor n14559 n14588 ; n14589
g14526 nor n8860 n9331 ; n14590
g14527 and n8418_not n14590 ; n14591
g14528 and n8421_not n14591 ; n14592
g14529 nor n13438 n14592 ; n14593
g14530 and a[8] n14593_not ; n14594
g14531 and a[8]_not n14593 ; n14595
g14532 nor n14594 n14595 ; n14596
g14533 and n14559 n14588 ; n14597
g14534 nor n14589 n14597 ; n14598
g14535 and n14596 n14598 ; n14599
g14536 nor n14589 n14599 ; n14600
g14537 and n14403 n14600_not ; n14601
g14538 and n14403_not n14600 ; n14602
g14539 nor n14601 n14602 ; n14603
g14540 and n3020 n12525 ; n14604
g14541 and n3028 n12528 ; n14605
g14542 and n3023 n12531 ; n14606
g14543 and n12643 n12645_not ; n14607
g14544 nor n12646 n14607 ; n14608
g14545 and n75 n14608 ; n14609
g14546 nor n14606 n14609 ; n14610
g14547 and n14605_not n14610 ; n14611
g14548 and n14604_not n14611 ; n14612
g14549 and n14603 n14612_not ; n14613
g14550 nor n14601 n14613 ; n14614
g14551 nor n14515 n14614 ; n14615
g14552 and n14516_not n14615 ; n14616
g14553 nor n14515 n14616 ; n14617
g14554 nor n14467 n14617 ; n14618
g14555 nor n14464 n14618 ; n14619
g14556 and n14437_not n14447 ; n14620
g14557 nor n14448 n14620 ; n14621
g14558 and n14619_not n14621 ; n14622
g14559 and n14619 n14621_not ; n14623
g14560 nor n14622 n14623 ; n14624
g14561 and n3457 n12508 ; n14625
g14562 and n3542 n12511 ; n14626
g14563 and n3606 n12513 ; n14627
g14564 nor n14626 n14627 ; n14628
g14565 and n14625_not n14628 ; n14629
g14566 and n3368_not n14629 ; n14630
g14567 and n13863_not n14629 ; n14631
g14568 nor n14630 n14631 ; n14632
g14569 and a[29] n14632_not ; n14633
g14570 and a[29]_not n14632 ; n14634
g14571 nor n14633 n14634 ; n14635
g14572 and n14624 n14635_not ; n14636
g14573 nor n14622 n14636 ; n14637
g14574 and n14452 n14637_not ; n14638
g14575 nor n14450 n14638 ; n14639
g14576 nor n14368 n14639 ; n14640
g14577 nor n14365 n14640 ; n14641
g14578 and n14255_not n14266 ; n14642
g14579 nor n14267 n14642 ; n14643
g14580 and n14641_not n14643 ; n14644
g14581 and n14641 n14643_not ; n14645
g14582 nor n14644 n14645 ; n14646
g14583 and n3884 n13491 ; n14647
g14584 and n3967 n12769 ; n14648
g14585 and n4046 n12889 ; n14649
g14586 nor n14648 n14649 ; n14650
g14587 and n14647_not n14650 ; n14651
g14588 and n4050 n13503_not ; n14652
g14589 and n14651 n14652_not ; n14653
g14590 and a[26] n14653_not ; n14654
g14591 and a[26] n14654_not ; n14655
g14592 nor n14653 n14654 ; n14656
g14593 nor n14655 n14656 ; n14657
g14594 and n14646 n14657_not ; n14658
g14595 nor n14644 n14658 ; n14659
g14596 nor n14350 n14659 ; n14660
g14597 and n14350 n14659 ; n14661
g14598 nor n14660 n14661 ; n14662
g14599 and n4694 n13597 ; n14663
g14600 and n4533 n13521 ; n14664
g14601 and n4604 n13515 ; n14665
g14602 nor n14664 n14665 ; n14666
g14603 and n14663_not n14666 ; n14667
g14604 and n4536 n13612_not ; n14668
g14605 and n14667 n14668_not ; n14669
g14606 and a[23] n14669_not ; n14670
g14607 and a[23] n14670_not ; n14671
g14608 nor n14669 n14670 ; n14672
g14609 nor n14671 n14672 ; n14673
g14610 and n14662 n14673_not ; n14674
g14611 nor n14660 n14674 ; n14675
g14612 nor n14347 n14675 ; n14676
g14613 nor n14344 n14676 ; n14677
g14614 nor n14330 n14677 ; n14678
g14615 and n14330 n14677 ; n14679
g14616 nor n14678 n14679 ; n14680
g14617 and n5496 n13438_not ; n14681
g14618 and n4935 n13627_not ; n14682
g14619 and n5407 n13941 ; n14683
g14620 nor n14682 n14683 ; n14684
g14621 and n14681_not n14684 ; n14685
g14622 and n4938 n14028 ; n14686
g14623 and n14685 n14686_not ; n14687
g14624 and a[20] n14687_not ; n14688
g14625 and a[20] n14688_not ; n14689
g14626 nor n14687 n14688 ; n14690
g14627 nor n14689 n14690 ; n14691
g14628 and n14680 n14691_not ; n14692
g14629 nor n14678 n14692 ; n14693
g14630 nor n14327 n14693 ; n14694
g14631 and n14327 n14693 ; n14695
g14632 nor n14694 n14695 ; n14696
g14633 and n14680 n14692_not ; n14697
g14634 nor n14691 n14692 ; n14698
g14635 nor n14697 n14698 ; n14699
g14636 and n14662 n14674_not ; n14700
g14637 nor n14673 n14674 ; n14701
g14638 nor n14700 n14701 ; n14702
g14639 and n14646 n14658_not ; n14703
g14640 nor n14657 n14658 ; n14704
g14641 nor n14703 n14704 ; n14705
g14642 and n14368 n14639 ; n14706
g14643 nor n14640 n14706 ; n14707
g14644 and n3884 n12889 ; n14708
g14645 and n3967 n12502 ; n14709
g14646 and n4046 n12769 ; n14710
g14647 nor n14709 n14710 ; n14711
g14648 and n14708_not n14711 ; n14712
g14649 and n4050 n12895 ; n14713
g14650 and n14712 n14713_not ; n14714
g14651 and a[26] n14714_not ; n14715
g14652 and a[26] n14715_not ; n14716
g14653 nor n14714 n14715 ; n14717
g14654 nor n14716 n14717 ; n14718
g14655 and n14707 n14718_not ; n14719
g14656 and n14707 n14719_not ; n14720
g14657 nor n14718 n14719 ; n14721
g14658 nor n14720 n14721 ; n14722
g14659 and n14452_not n14637 ; n14723
g14660 nor n14638 n14723 ; n14724
g14661 and n3457 n12505 ; n14725
g14662 and n3542 n12513 ; n14726
g14663 and n3606 n12508 ; n14727
g14664 nor n14726 n14727 ; n14728
g14665 and n14725_not n14728 ; n14729
g14666 and n3368 n14051_not ; n14730
g14667 and n14729 n14730_not ; n14731
g14668 and a[29] n14731_not ; n14732
g14669 and a[29] n14732_not ; n14733
g14670 nor n14731 n14732 ; n14734
g14671 nor n14733 n14734 ; n14735
g14672 and n14724 n14735_not ; n14736
g14673 and n14724 n14736_not ; n14737
g14674 nor n14735 n14736 ; n14738
g14675 nor n14737 n14738 ; n14739
g14676 and n3884 n12769 ; n14740
g14677 and n3967 n12370 ; n14741
g14678 and n4046 n12502 ; n14742
g14679 nor n14741 n14742 ; n14743
g14680 and n14740_not n14743 ; n14744
g14681 and n4050 n12999 ; n14745
g14682 and n14744 n14745_not ; n14746
g14683 and a[26] n14746_not ; n14747
g14684 and a[26] n14747_not ; n14748
g14685 nor n14746 n14747 ; n14749
g14686 nor n14748 n14749 ; n14750
g14687 nor n14739 n14750 ; n14751
g14688 nor n14736 n14751 ; n14752
g14689 nor n14722 n14752 ; n14753
g14690 nor n14719 n14753 ; n14754
g14691 nor n14705 n14754 ; n14755
g14692 and n14705 n14754 ; n14756
g14693 nor n14755 n14756 ; n14757
g14694 and n4694 n13515 ; n14758
g14695 and n4533 n13518 ; n14759
g14696 and n4604 n13521 ; n14760
g14697 nor n14759 n14760 ; n14761
g14698 and n14758_not n14761 ; n14762
g14699 and n4536 n13541 ; n14763
g14700 and n14762 n14763_not ; n14764
g14701 and a[23] n14764_not ; n14765
g14702 and a[23] n14765_not ; n14766
g14703 nor n14764 n14765 ; n14767
g14704 nor n14766 n14767 ; n14768
g14705 and n14757 n14768_not ; n14769
g14706 nor n14755 n14769 ; n14770
g14707 nor n14702 n14770 ; n14771
g14708 and n14702 n14770 ; n14772
g14709 nor n14771 n14772 ; n14773
g14710 and n5496 n13627_not ; n14774
g14711 and n4935 n13630 ; n14775
g14712 and n5407 n13633 ; n14776
g14713 nor n14775 n14776 ; n14777
g14714 and n14774_not n14777 ; n14778
g14715 and n4938 n13654_not ; n14779
g14716 and n14778 n14779_not ; n14780
g14717 and a[20] n14780_not ; n14781
g14718 and a[20] n14781_not ; n14782
g14719 nor n14780 n14781 ; n14783
g14720 nor n14782 n14783 ; n14784
g14721 and n14773 n14784_not ; n14785
g14722 nor n14771 n14785 ; n14786
g14723 and n5496 n13941 ; n14787
g14724 and n4935 n13633 ; n14788
g14725 and n5407 n13627_not ; n14789
g14726 nor n14788 n14789 ; n14790
g14727 and n14787_not n14790 ; n14791
g14728 and n4938 n14136 ; n14792
g14729 and n14791 n14792_not ; n14793
g14730 and a[20] n14793_not ; n14794
g14731 and a[20] n14794_not ; n14795
g14732 nor n14793 n14794 ; n14796
g14733 nor n14795 n14796 ; n14797
g14734 nor n14786 n14797 ; n14798
g14735 and n14347 n14675 ; n14799
g14736 nor n14676 n14799 ; n14800
g14737 nor n14786 n14798 ; n14801
g14738 nor n14797 n14798 ; n14802
g14739 nor n14801 n14802 ; n14803
g14740 and n14800 n14803_not ; n14804
g14741 nor n14798 n14804 ; n14805
g14742 nor n14699 n14805 ; n14806
g14743 nor n14699 n14806 ; n14807
g14744 nor n14805 n14806 ; n14808
g14745 nor n14807 n14808 ; n14809
g14746 and n14757 n14769_not ; n14810
g14747 nor n14768 n14769 ; n14811
g14748 nor n14810 n14811 ; n14812
g14749 and n14722 n14752 ; n14813
g14750 nor n14753 n14813 ; n14814
g14751 and n4694 n13521 ; n14815
g14752 and n4533 n13491 ; n14816
g14753 and n4604 n13518 ; n14817
g14754 nor n14816 n14817 ; n14818
g14755 and n14815_not n14818 ; n14819
g14756 and n4536 n13909_not ; n14820
g14757 and n14819 n14820_not ; n14821
g14758 and a[23] n14821_not ; n14822
g14759 and a[23] n14822_not ; n14823
g14760 nor n14821 n14822 ; n14824
g14761 nor n14823 n14824 ; n14825
g14762 and n14814 n14825_not ; n14826
g14763 and n14814 n14826_not ; n14827
g14764 nor n14825 n14826 ; n14828
g14765 nor n14827 n14828 ; n14829
g14766 nor n14739 n14751 ; n14830
g14767 nor n14750 n14751 ; n14831
g14768 nor n14830 n14831 ; n14832
g14769 nor n14614 n14616 ; n14833
g14770 and n14516_not n14617 ; n14834
g14771 nor n14833 n14834 ; n14835
g14772 and n12647 n12649_not ; n14836
g14773 nor n12650 n14836 ; n14837
g14774 and n75 n14837 ; n14838
g14775 and n3020 n12522 ; n14839
g14776 and n3023 n12528 ; n14840
g14777 and n3028 n12525 ; n14841
g14778 nor n14840 n14841 ; n14842
g14779 and n14839_not n14842 ; n14843
g14780 and n14838_not n14843 ; n14844
g14781 nor n14835 n14844 ; n14845
g14782 nor n14835 n14845 ; n14846
g14783 nor n14844 n14845 ; n14847
g14784 nor n14846 n14847 ; n14848
g14785 and n3457 n12511 ; n14849
g14786 and n3542 n12519 ; n14850
g14787 and n3606 n12516 ; n14851
g14788 nor n14850 n14851 ; n14852
g14789 and n14849_not n14852 ; n14853
g14790 and n3368_not n14853 ; n14854
g14791 and n14233 n14853 ; n14855
g14792 nor n14854 n14855 ; n14856
g14793 and a[29] n14856_not ; n14857
g14794 and a[29]_not n14856 ; n14858
g14795 nor n14857 n14858 ; n14859
g14796 nor n14848 n14859 ; n14860
g14797 nor n14845 n14860 ; n14861
g14798 nor n14467 n14618 ; n14862
g14799 nor n14617 n14618 ; n14863
g14800 nor n14862 n14863 ; n14864
g14801 nor n14861 n14864 ; n14865
g14802 nor n14861 n14865 ; n14866
g14803 nor n14864 n14865 ; n14867
g14804 nor n14866 n14867 ; n14868
g14805 and n3457 n12513 ; n14869
g14806 and n3542 n12516 ; n14870
g14807 and n3606 n12511 ; n14871
g14808 nor n14870 n14871 ; n14872
g14809 and n14869_not n14872 ; n14873
g14810 and n3368 n14177 ; n14874
g14811 and n14873 n14874_not ; n14875
g14812 and a[29] n14875_not ; n14876
g14813 and a[29] n14876_not ; n14877
g14814 nor n14875 n14876 ; n14878
g14815 nor n14877 n14878 ; n14879
g14816 nor n14868 n14879 ; n14880
g14817 nor n14865 n14880 ; n14881
g14818 and n14624_not n14635 ; n14882
g14819 nor n14636 n14882 ; n14883
g14820 and n14881_not n14883 ; n14884
g14821 and n14881 n14883_not ; n14885
g14822 nor n14884 n14885 ; n14886
g14823 and n3884 n12502 ; n14887
g14824 and n3967 n12505 ; n14888
g14825 and n4046 n12370 ; n14889
g14826 nor n14888 n14889 ; n14890
g14827 and n14887_not n14890 ; n14891
g14828 and n4050 n13736_not ; n14892
g14829 and n14891 n14892_not ; n14893
g14830 and a[26] n14893_not ; n14894
g14831 and a[26] n14894_not ; n14895
g14832 nor n14893 n14894 ; n14896
g14833 nor n14895 n14896 ; n14897
g14834 and n14886 n14897_not ; n14898
g14835 nor n14884 n14898 ; n14899
g14836 nor n14832 n14899 ; n14900
g14837 and n14832 n14899 ; n14901
g14838 nor n14900 n14901 ; n14902
g14839 and n4694 n13518 ; n14903
g14840 and n4533 n12889 ; n14904
g14841 and n4604 n13491 ; n14905
g14842 nor n14904 n14905 ; n14906
g14843 and n14903_not n14906 ; n14907
g14844 and n4536 n13584 ; n14908
g14845 and n14907 n14908_not ; n14909
g14846 and a[23] n14909_not ; n14910
g14847 and a[23] n14910_not ; n14911
g14848 nor n14909 n14910 ; n14912
g14849 nor n14911 n14912 ; n14913
g14850 and n14902 n14913_not ; n14914
g14851 nor n14900 n14914 ; n14915
g14852 nor n14829 n14915 ; n14916
g14853 nor n14826 n14916 ; n14917
g14854 nor n14812 n14917 ; n14918
g14855 and n14812 n14917 ; n14919
g14856 nor n14918 n14919 ; n14920
g14857 and n5496 n13633 ; n14921
g14858 and n4935 n13597 ; n14922
g14859 and n5407 n13630 ; n14923
g14860 nor n14922 n14923 ; n14924
g14861 and n14921_not n14924 ; n14925
g14862 and n4938 n13929 ; n14926
g14863 and n14925 n14926_not ; n14927
g14864 and a[20] n14927_not ; n14928
g14865 and a[20] n14928_not ; n14929
g14866 nor n14927 n14928 ; n14930
g14867 nor n14929 n14930 ; n14931
g14868 and n14920 n14931_not ; n14932
g14869 nor n14918 n14932 ; n14933
g14870 nor n13438 n13717 ; n14934
g14871 and n5663 n13941 ; n14935
g14872 nor n14934 n14935 ; n14936
g14873 and n5666_not n14936 ; n14937
g14874 and n13951 n14936 ; n14938
g14875 nor n14937 n14938 ; n14939
g14876 and a[17] n14939_not ; n14940
g14877 and a[17]_not n14939 ; n14941
g14878 nor n14940 n14941 ; n14942
g14879 nor n14933 n14942 ; n14943
g14880 and n14773 n14785_not ; n14944
g14881 nor n14784 n14785 ; n14945
g14882 nor n14944 n14945 ; n14946
g14883 and n14933 n14942 ; n14947
g14884 nor n14943 n14947 ; n14948
g14885 and n14946_not n14948 ; n14949
g14886 nor n14943 n14949 ; n14950
g14887 and n14800_not n14803 ; n14951
g14888 nor n14804 n14951 ; n14952
g14889 and n14950_not n14952 ; n14953
g14890 nor n14946 n14949 ; n14954
g14891 and n14948 n14949_not ; n14955
g14892 nor n14954 n14955 ; n14956
g14893 and n14920 n14932_not ; n14957
g14894 nor n14931 n14932 ; n14958
g14895 nor n14957 n14958 ; n14959
g14896 and n14829 n14915 ; n14960
g14897 nor n14916 n14960 ; n14961
g14898 and n5496 n13630 ; n14962
g14899 and n4935 n13515 ; n14963
g14900 and n5407 n13597 ; n14964
g14901 nor n14963 n14964 ; n14965
g14902 and n14962_not n14965 ; n14966
g14903 and n4938 n13976 ; n14967
g14904 and n14966 n14967_not ; n14968
g14905 and a[20] n14968_not ; n14969
g14906 and a[20] n14969_not ; n14970
g14907 nor n14968 n14969 ; n14971
g14908 nor n14970 n14971 ; n14972
g14909 and n14961 n14972_not ; n14973
g14910 and n14961 n14973_not ; n14974
g14911 nor n14972 n14973 ; n14975
g14912 nor n14974 n14975 ; n14976
g14913 and n14902 n14914_not ; n14977
g14914 nor n14913 n14914 ; n14978
g14915 nor n14977 n14978 ; n14979
g14916 and n14886 n14898_not ; n14980
g14917 nor n14897 n14898 ; n14981
g14918 nor n14980 n14981 ; n14982
g14919 nor n14868 n14880 ; n14983
g14920 nor n14879 n14880 ; n14984
g14921 nor n14983 n14984 ; n14985
g14922 and n3884 n12370 ; n14986
g14923 and n3967 n12508 ; n14987
g14924 and n4046 n12505 ; n14988
g14925 nor n14987 n14988 ; n14989
g14926 and n14986_not n14989 ; n14990
g14927 and n4050 n13748_not ; n14991
g14928 and n14990 n14991_not ; n14992
g14929 and a[26] n14992_not ; n14993
g14930 and a[26] n14993_not ; n14994
g14931 nor n14992 n14993 ; n14995
g14932 nor n14994 n14995 ; n14996
g14933 nor n14985 n14996 ; n14997
g14934 nor n14985 n14997 ; n14998
g14935 nor n14996 n14997 ; n14999
g14936 nor n14998 n14999 ; n15000
g14937 nor n12639 n12642 ; n15001
g14938 and n12640_not n12643 ; n15002
g14939 nor n15001 n15002 ; n15003
g14940 and n75 n15003_not ; n15004
g14941 and n3020 n12528 ; n15005
g14942 and n3023 n12534 ; n15006
g14943 and n3028 n12531 ; n15007
g14944 nor n15006 n15007 ; n15008
g14945 and n15005_not n15008 ; n15009
g14946 and n15004_not n15009 ; n15010
g14947 and n667_not n1139 ; n15011
g14948 and n886_not n15011 ; n15012
g14949 and n256 n5173 ; n15013
g14950 and n15012 n15013 ; n15014
g14951 and n2093 n15014 ; n15015
g14952 and n1958 n15015 ; n15016
g14953 and n3565 n15016 ; n15017
g14954 and n2738 n15017 ; n15018
g14955 and n187 n15018 ; n15019
g14956 and n2170 n15019 ; n15020
g14957 and n471 n15020 ; n15021
g14958 and n1857 n15021 ; n15022
g14959 and n427_not n15022 ; n15023
g14960 and n289_not n15023 ; n15024
g14961 and n281_not n15024 ; n15025
g14962 and n557_not n15025 ; n15026
g14963 and n237_not n15026 ; n15027
g14964 and n201_not n15027 ; n15028
g14965 and n14559 n15028_not ; n15029
g14966 and n14559_not n15028 ; n15030
g14967 and n11053 n11054 ; n15031
g14968 nor n13438 n15031 ; n15032
g14969 and a[2] n15032_not ; n15033
g14970 and a[2]_not n15032 ; n15034
g14971 nor n15033 n15034 ; n15035
g14972 and n1738 n3645 ; n15036
g14973 and n1070 n15036 ; n15037
g14974 and n3548 n15037 ; n15038
g14975 and n439 n15038 ; n15039
g14976 and n508 n15039 ; n15040
g14977 and n168_not n15040 ; n15041
g14978 and n402_not n15041 ; n15042
g14979 and n961_not n15042 ; n15043
g14980 and n170_not n15043 ; n15044
g14981 and n1010_not n15044 ; n15045
g14982 and n489_not n15045 ; n15046
g14983 and n771_not n15046 ; n15047
g14984 and n2651 n14479 ; n15048
g14985 and n301_not n15048 ; n15049
g14986 and n229_not n15049 ; n15050
g14987 and n3194 n13827 ; n15051
g14988 and n370 n15051 ; n15052
g14989 and n2241 n15052 ; n15053
g14990 and n15050 n15053 ; n15054
g14991 and n12810 n15054 ; n15055
g14992 and n2591 n15055 ; n15056
g14993 and n294 n15056 ; n15057
g14994 and n1781 n15057 ; n15058
g14995 and n15047 n15058 ; n15059
g14996 and n1389 n15059 ; n15060
g14997 and n417_not n15060 ; n15061
g14998 and n137 n3192 ; n15062
g14999 and n6102 n15062 ; n15063
g15000 and n6667 n15063 ; n15064
g15001 and n14381 n15064 ; n15065
g15002 and n12404 n15065 ; n15066
g15003 and n15061 n15066 ; n15067
g15004 and n1523 n15067 ; n15068
g15005 and n247 n15068 ; n15069
g15006 and n3252 n15069 ; n15070
g15007 and n620_not n15070 ; n15071
g15008 and n352_not n15071 ; n15072
g15009 and n118_not n15072 ; n15073
g15010 and n532_not n15073 ; n15074
g15011 and n15035 n15074_not ; n15075
g15012 nor n71 n10434 ; n15076
g15013 and n9867_not n15076 ; n15077
g15014 and n9870_not n15077 ; n15078
g15015 nor n13438 n15078 ; n15079
g15016 and a[5]_not n15079 ; n15080
g15017 and n15035 n15074 ; n15081
g15018 nor n15035 n15074 ; n15082
g15019 nor n15081 n15082 ; n15083
g15020 and a[5] n15079_not ; n15084
g15021 nor n15083 n15084 ; n15085
g15022 and n15080_not n15085 ; n15086
g15023 nor n15075 n15086 ; n15087
g15024 and n14559 n15087_not ; n15088
g15025 and n14559_not n15087 ; n15089
g15026 nor n15088 n15089 ; n15090
g15027 and n3020 n12534 ; n15091
g15028 and n3028 n12537 ; n15092
g15029 and n3023 n12540 ; n15093
g15030 nor n12631 n12634 ; n15094
g15031 and n12632_not n12635 ; n15095
g15032 nor n15094 n15095 ; n15096
g15033 and n75 n15096_not ; n15097
g15034 nor n15093 n15097 ; n15098
g15035 and n15092_not n15098 ; n15099
g15036 and n15091_not n15099 ; n15100
g15037 and n15090 n15100_not ; n15101
g15038 nor n15088 n15101 ; n15102
g15039 nor n15029 n15102 ; n15103
g15040 and n15030_not n15103 ; n15104
g15041 nor n15029 n15104 ; n15105
g15042 nor n14596 n14598 ; n15106
g15043 nor n14599 n15106 ; n15107
g15044 and n15105_not n15107 ; n15108
g15045 and n15105 n15107_not ; n15109
g15046 nor n15108 n15109 ; n15110
g15047 and n15010_not n15110 ; n15111
g15048 nor n15108 n15111 ; n15112
g15049 and n14603_not n14612 ; n15113
g15050 nor n14613 n15113 ; n15114
g15051 and n15112_not n15114 ; n15115
g15052 and n15112 n15114_not ; n15116
g15053 nor n15115 n15116 ; n15117
g15054 and n3457 n12516 ; n15118
g15055 and n3542 n12522 ; n15119
g15056 and n3606 n12519 ; n15120
g15057 nor n15119 n15120 ; n15121
g15058 and n15118_not n15121 ; n15122
g15059 and n3368_not n15122 ; n15123
g15060 and n14443 n15122 ; n15124
g15061 nor n15123 n15124 ; n15125
g15062 and a[29] n15125_not ; n15126
g15063 and a[29]_not n15125 ; n15127
g15064 nor n15126 n15127 ; n15128
g15065 and n15117 n15128_not ; n15129
g15066 nor n15115 n15129 ; n15130
g15067 and n14848 n14859 ; n15131
g15068 nor n14860 n15131 ; n15132
g15069 and n15130_not n15132 ; n15133
g15070 and n15130 n15132_not ; n15134
g15071 nor n15133 n15134 ; n15135
g15072 and n3884 n12505 ; n15136
g15073 and n3967 n12513 ; n15137
g15074 and n4046 n12508 ; n15138
g15075 nor n15137 n15138 ; n15139
g15076 and n15136_not n15139 ; n15140
g15077 and n4050 n14051_not ; n15141
g15078 and n15140 n15141_not ; n15142
g15079 and a[26] n15142_not ; n15143
g15080 and a[26] n15143_not ; n15144
g15081 nor n15142 n15143 ; n15145
g15082 nor n15144 n15145 ; n15146
g15083 and n15135 n15146_not ; n15147
g15084 nor n15133 n15147 ; n15148
g15085 nor n15000 n15148 ; n15149
g15086 nor n14997 n15149 ; n15150
g15087 nor n14982 n15150 ; n15151
g15088 and n14982 n15150 ; n15152
g15089 nor n15151 n15152 ; n15153
g15090 and n4694 n13491 ; n15154
g15091 and n4533 n12769 ; n15155
g15092 and n4604 n12889 ; n15156
g15093 nor n15155 n15156 ; n15157
g15094 and n15154_not n15157 ; n15158
g15095 and n4536 n13503_not ; n15159
g15096 and n15158 n15159_not ; n15160
g15097 and a[23] n15160_not ; n15161
g15098 and a[23] n15161_not ; n15162
g15099 nor n15160 n15161 ; n15163
g15100 nor n15162 n15163 ; n15164
g15101 and n15153 n15164_not ; n15165
g15102 nor n15151 n15165 ; n15166
g15103 nor n14979 n15166 ; n15167
g15104 and n14979 n15166 ; n15168
g15105 nor n15167 n15168 ; n15169
g15106 and n5496 n13597 ; n15170
g15107 and n4935 n13521 ; n15171
g15108 and n5407 n13515 ; n15172
g15109 nor n15171 n15172 ; n15173
g15110 and n15170_not n15173 ; n15174
g15111 and n4938 n13612_not ; n15175
g15112 and n15174 n15175_not ; n15176
g15113 and a[20] n15176_not ; n15177
g15114 and a[20] n15177_not ; n15178
g15115 nor n15176 n15177 ; n15179
g15116 nor n15178 n15179 ; n15180
g15117 and n15169 n15180_not ; n15181
g15118 nor n15167 n15181 ; n15182
g15119 nor n14976 n15182 ; n15183
g15120 nor n14973 n15183 ; n15184
g15121 nor n14959 n15184 ; n15185
g15122 and n14959 n15184 ; n15186
g15123 nor n15185 n15186 ; n15187
g15124 and n6233 n13438_not ; n15188
g15125 and n5663 n13627_not ; n15189
g15126 and n5939 n13941 ; n15190
g15127 nor n15189 n15190 ; n15191
g15128 and n15188_not n15191 ; n15192
g15129 and n5666 n14028 ; n15193
g15130 and n15192 n15193_not ; n15194
g15131 and a[17] n15194_not ; n15195
g15132 and a[17] n15195_not ; n15196
g15133 nor n15194 n15195 ; n15197
g15134 nor n15196 n15197 ; n15198
g15135 and n15187 n15198_not ; n15199
g15136 nor n15185 n15199 ; n15200
g15137 nor n14956 n15200 ; n15201
g15138 and n14956 n15200 ; n15202
g15139 nor n15201 n15202 ; n15203
g15140 and n15187 n15199_not ; n15204
g15141 nor n15198 n15199 ; n15205
g15142 nor n15204 n15205 ; n15206
g15143 and n15169 n15181_not ; n15207
g15144 nor n15180 n15181 ; n15208
g15145 nor n15207 n15208 ; n15209
g15146 and n15153 n15165_not ; n15210
g15147 nor n15164 n15165 ; n15211
g15148 nor n15210 n15211 ; n15212
g15149 and n15000 n15148 ; n15213
g15150 nor n15149 n15213 ; n15214
g15151 and n4694 n12889 ; n15215
g15152 and n4533 n12502 ; n15216
g15153 and n4604 n12769 ; n15217
g15154 nor n15216 n15217 ; n15218
g15155 and n15215_not n15218 ; n15219
g15156 and n4536 n12895 ; n15220
g15157 and n15219 n15220_not ; n15221
g15158 and a[23] n15221_not ; n15222
g15159 and a[23] n15222_not ; n15223
g15160 nor n15221 n15222 ; n15224
g15161 nor n15223 n15224 ; n15225
g15162 and n15214 n15225_not ; n15226
g15163 and n15214 n15226_not ; n15227
g15164 nor n15225 n15226 ; n15228
g15165 nor n15227 n15228 ; n15229
g15166 and n15135 n15147_not ; n15230
g15167 nor n15146 n15147 ; n15231
g15168 nor n15230 n15231 ; n15232
g15169 and n15110 n15111_not ; n15233
g15170 nor n15010 n15111 ; n15234
g15171 nor n15233 n15234 ; n15235
g15172 and n3457 n12519 ; n15236
g15173 and n3542 n12525 ; n15237
g15174 and n3606 n12522 ; n15238
g15175 nor n15237 n15238 ; n15239
g15176 and n15236_not n15239 ; n15240
g15177 and n3368 n14454 ; n15241
g15178 and n15240 n15241_not ; n15242
g15179 and a[29] n15242_not ; n15243
g15180 and a[29] n15243_not ; n15244
g15181 nor n15242 n15243 ; n15245
g15182 nor n15244 n15245 ; n15246
g15183 nor n15235 n15246 ; n15247
g15184 nor n15235 n15247 ; n15248
g15185 nor n15246 n15247 ; n15249
g15186 nor n15248 n15249 ; n15250
g15187 nor n15102 n15104 ; n15251
g15188 and n15030_not n15105 ; n15252
g15189 nor n15251 n15252 ; n15253
g15190 and n12635 n12637_not ; n15254
g15191 nor n12638 n15254 ; n15255
g15192 and n75 n15255 ; n15256
g15193 and n3020 n12531 ; n15257
g15194 and n3023 n12537 ; n15258
g15195 and n3028 n12534 ; n15259
g15196 nor n15258 n15259 ; n15260
g15197 and n15257_not n15260 ; n15261
g15198 and n15256_not n15261 ; n15262
g15199 nor n15253 n15262 ; n15263
g15200 nor n15253 n15263 ; n15264
g15201 nor n15262 n15263 ; n15265
g15202 nor n15264 n15265 ; n15266
g15203 and n1185 n2349 ; n15267
g15204 and n1894 n15267 ; n15268
g15205 and n3743 n15268 ; n15269
g15206 and n3675 n15269 ; n15270
g15207 and n5785 n15270 ; n15271
g15208 and n2778 n15271 ; n15272
g15209 and n1180 n15272 ; n15273
g15210 and n469_not n15273 ; n15274
g15211 and n1101_not n15274 ; n15275
g15212 and n513_not n15275 ; n15276
g15213 and n298_not n15276 ; n15277
g15214 and n372_not n15277 ; n15278
g15215 and n157_not n15278 ; n15279
g15216 and n1104_not n15279 ; n15280
g15217 and n592_not n15280 ; n15281
g15218 and n295_not n15281 ; n15282
g15219 and n525_not n15282 ; n15283
g15220 nor n15035 n15283 ; n15284
g15221 and n634 n13774 ; n15285
g15222 and n328_not n15285 ; n15286
g15223 and n13012 n15286 ; n15287
g15224 and n1709 n15287 ; n15288
g15225 and n15061 n15288 ; n15289
g15226 and n503 n15289 ; n15290
g15227 and n512 n15290 ; n15291
g15228 and n1915 n15291 ; n15292
g15229 and n1183 n15292 ; n15293
g15230 and n285 n15293 ; n15294
g15231 and n730 n15294 ; n15295
g15232 and n1783 n15295 ; n15296
g15233 and n202 n15296 ; n15297
g15234 and n4101 n15297 ; n15298
g15235 and n746_not n15298 ; n15299
g15236 and n239_not n15299 ; n15300
g15237 and n192_not n15300 ; n15301
g15238 and n453_not n15301 ; n15302
g15239 and n883_not n15302 ; n15303
g15240 and n886_not n15303 ; n15304
g15241 and n337_not n15304 ; n15305
g15242 nor n15035 n15305 ; n15306
g15243 and n1557 n2209 ; n15307
g15244 and n420_not n15307 ; n15308
g15245 and n278_not n15308 ; n15309
g15246 and n435_not n15309 ; n15310
g15247 and n589_not n15310 ; n15311
g15248 and n569_not n15311 ; n15312
g15249 and n365 n1329 ; n15313
g15250 and n2468 n15313 ; n15314
g15251 and n12431 n15314 ; n15315
g15252 and n5085 n15315 ; n15316
g15253 and n1725 n15316 ; n15317
g15254 and n15312 n15317 ; n15318
g15255 and n2346 n15318 ; n15319
g15256 and n151_not n15319 ; n15320
g15257 and n275_not n15320 ; n15321
g15258 and n438_not n15321 ; n15322
g15259 and n1203_not n15322 ; n15323
g15260 and n623_not n15323 ; n15324
g15261 and n1692 n15324 ; n15325
g15262 and n354_not n15325 ; n15326
g15263 and n168_not n15326 ; n15327
g15264 and n296_not n15327 ; n15328
g15265 and n1104_not n15328 ; n15329
g15266 and n532_not n15329 ; n15330
g15267 and n1306_not n3380 ; n15331
g15268 and n746_not n15331 ; n15332
g15269 and n232_not n15332 ; n15333
g15270 and n152_not n15333 ; n15334
g15271 and n203_not n15334 ; n15335
g15272 and n245_not n15335 ; n15336
g15273 and n932_not n15336 ; n15337
g15274 and n475 n1530 ; n15338
g15275 and n2809 n15338 ; n15339
g15276 and n1759 n15339 ; n15340
g15277 and n15337 n15340 ; n15341
g15278 and n12973 n15341 ; n15342
g15279 and n15330 n15342 ; n15343
g15280 and n14479 n15343 ; n15344
g15281 and n1237 n15344 ; n15345
g15282 and n111_not n15345 ; n15346
g15283 and n150_not n15346 ; n15347
g15284 and n571_not n15347 ; n15348
g15285 and n118_not n15348 ; n15349
g15286 and n107_not n15349 ; n15350
g15287 and n286_not n15350 ; n15351
g15288 and n592_not n15351 ; n15352
g15289 nor n15035 n15352 ; n15353
g15290 nor n12615 n12618 ; n15354
g15291 and n12616_not n12619 ; n15355
g15292 nor n15354 n15355 ; n15356
g15293 and n75 n15356_not ; n15357
g15294 and n3020 n12546 ; n15358
g15295 and n3023 n12552 ; n15359
g15296 and n3028 n12549 ; n15360
g15297 nor n15359 n15360 ; n15361
g15298 and n15358_not n15361 ; n15362
g15299 and n15357_not n15362 ; n15363
g15300 and n15035 n15352 ; n15364
g15301 nor n15363 n15364 ; n15365
g15302 and n15353_not n15365 ; n15366
g15303 nor n15353 n15366 ; n15367
g15304 and n15035 n15305 ; n15368
g15305 nor n15367 n15368 ; n15369
g15306 and n15306_not n15369 ; n15370
g15307 nor n15306 n15370 ; n15371
g15308 and n15035 n15283 ; n15372
g15309 nor n15371 n15372 ; n15373
g15310 and n15284_not n15373 ; n15374
g15311 nor n15284 n15374 ; n15375
g15312 nor n15083 n15086 ; n15376
g15313 nor n15084 n15086 ; n15377
g15314 and n15080_not n15377 ; n15378
g15315 nor n15376 n15378 ; n15379
g15316 and n15375_not n15379 ; n15380
g15317 and n15375 n15379_not ; n15381
g15318 nor n15380 n15381 ; n15382
g15319 nor n12627 n12630 ; n15383
g15320 and n12628_not n12631 ; n15384
g15321 nor n15383 n15384 ; n15385
g15322 and n75 n15385_not ; n15386
g15323 and n3020 n12537 ; n15387
g15324 and n3023 n12543 ; n15388
g15325 and n3028 n12540 ; n15389
g15326 nor n15388 n15389 ; n15390
g15327 and n15387_not n15390 ; n15391
g15328 and n15386_not n15391 ; n15392
g15329 nor n15382 n15392 ; n15393
g15330 nor n15375 n15379 ; n15394
g15331 nor n15393 n15394 ; n15395
g15332 and n15090_not n15100 ; n15396
g15333 nor n15101 n15396 ; n15397
g15334 and n15395_not n15397 ; n15398
g15335 and n15395 n15397_not ; n15399
g15336 nor n15398 n15399 ; n15400
g15337 and n3457 n12525 ; n15401
g15338 and n3542 n12531 ; n15402
g15339 and n3606 n12528 ; n15403
g15340 nor n15402 n15403 ; n15404
g15341 and n15401_not n15404 ; n15405
g15342 and n3368_not n15405 ; n15406
g15343 and n14608_not n15405 ; n15407
g15344 nor n15406 n15407 ; n15408
g15345 and a[29] n15408_not ; n15409
g15346 and a[29]_not n15408 ; n15410
g15347 nor n15409 n15410 ; n15411
g15348 and n15400 n15411_not ; n15412
g15349 nor n15398 n15412 ; n15413
g15350 nor n15266 n15413 ; n15414
g15351 nor n15263 n15414 ; n15415
g15352 nor n15250 n15415 ; n15416
g15353 nor n15247 n15416 ; n15417
g15354 and n15117_not n15128 ; n15418
g15355 nor n15129 n15418 ; n15419
g15356 and n15417_not n15419 ; n15420
g15357 and n15417 n15419_not ; n15421
g15358 nor n15420 n15421 ; n15422
g15359 and n3884 n12508 ; n15423
g15360 and n3967 n12511 ; n15424
g15361 and n4046 n12513 ; n15425
g15362 nor n15424 n15425 ; n15426
g15363 and n15423_not n15426 ; n15427
g15364 and n4050 n13863 ; n15428
g15365 and n15427 n15428_not ; n15429
g15366 and a[26] n15429_not ; n15430
g15367 and a[26] n15430_not ; n15431
g15368 nor n15429 n15430 ; n15432
g15369 nor n15431 n15432 ; n15433
g15370 and n15422 n15433_not ; n15434
g15371 nor n15420 n15434 ; n15435
g15372 nor n15232 n15435 ; n15436
g15373 and n15232 n15435 ; n15437
g15374 nor n15436 n15437 ; n15438
g15375 and n4694 n12769 ; n15439
g15376 and n4533 n12370 ; n15440
g15377 and n4604 n12502 ; n15441
g15378 nor n15440 n15441 ; n15442
g15379 and n15439_not n15442 ; n15443
g15380 and n4536 n12999 ; n15444
g15381 and n15443 n15444_not ; n15445
g15382 and a[23] n15445_not ; n15446
g15383 and a[23] n15446_not ; n15447
g15384 nor n15445 n15446 ; n15448
g15385 nor n15447 n15448 ; n15449
g15386 and n15438 n15449_not ; n15450
g15387 nor n15436 n15450 ; n15451
g15388 nor n15229 n15451 ; n15452
g15389 nor n15226 n15452 ; n15453
g15390 nor n15212 n15453 ; n15454
g15391 and n15212 n15453 ; n15455
g15392 nor n15454 n15455 ; n15456
g15393 and n5496 n13515 ; n15457
g15394 and n4935 n13518 ; n15458
g15395 and n5407 n13521 ; n15459
g15396 nor n15458 n15459 ; n15460
g15397 and n15457_not n15460 ; n15461
g15398 and n4938 n13541 ; n15462
g15399 and n15461 n15462_not ; n15463
g15400 and a[20] n15463_not ; n15464
g15401 and a[20] n15464_not ; n15465
g15402 nor n15463 n15464 ; n15466
g15403 nor n15465 n15466 ; n15467
g15404 and n15456 n15467_not ; n15468
g15405 nor n15454 n15468 ; n15469
g15406 nor n15209 n15469 ; n15470
g15407 and n15209 n15469 ; n15471
g15408 nor n15470 n15471 ; n15472
g15409 and n6233 n13627_not ; n15473
g15410 and n5663 n13630 ; n15474
g15411 and n5939 n13633 ; n15475
g15412 nor n15474 n15475 ; n15476
g15413 and n15473_not n15476 ; n15477
g15414 and n5666 n13654_not ; n15478
g15415 and n15477 n15478_not ; n15479
g15416 and a[17] n15479_not ; n15480
g15417 and a[17] n15480_not ; n15481
g15418 nor n15479 n15480 ; n15482
g15419 nor n15481 n15482 ; n15483
g15420 and n15472 n15483_not ; n15484
g15421 nor n15470 n15484 ; n15485
g15422 and n6233 n13941 ; n15486
g15423 and n5663 n13633 ; n15487
g15424 and n5939 n13627_not ; n15488
g15425 nor n15487 n15488 ; n15489
g15426 and n15486_not n15489 ; n15490
g15427 and n5666 n14136 ; n15491
g15428 and n15490 n15491_not ; n15492
g15429 and a[17] n15492_not ; n15493
g15430 and a[17] n15493_not ; n15494
g15431 nor n15492 n15493 ; n15495
g15432 nor n15494 n15495 ; n15496
g15433 nor n15485 n15496 ; n15497
g15434 and n14976 n15182 ; n15498
g15435 nor n15183 n15498 ; n15499
g15436 nor n15485 n15497 ; n15500
g15437 nor n15496 n15497 ; n15501
g15438 nor n15500 n15501 ; n15502
g15439 and n15499 n15502_not ; n15503
g15440 nor n15497 n15503 ; n15504
g15441 nor n15206 n15504 ; n15505
g15442 nor n15206 n15505 ; n15506
g15443 nor n15504 n15505 ; n15507
g15444 nor n15506 n15507 ; n15508
g15445 and n15456 n15468_not ; n15509
g15446 nor n15467 n15468 ; n15510
g15447 nor n15509 n15510 ; n15511
g15448 and n15229 n15451 ; n15512
g15449 nor n15452 n15512 ; n15513
g15450 and n5496 n13521 ; n15514
g15451 and n4935 n13491 ; n15515
g15452 and n5407 n13518 ; n15516
g15453 nor n15515 n15516 ; n15517
g15454 and n15514_not n15517 ; n15518
g15455 and n4938 n13909_not ; n15519
g15456 and n15518 n15519_not ; n15520
g15457 and a[20] n15520_not ; n15521
g15458 and a[20] n15521_not ; n15522
g15459 nor n15520 n15521 ; n15523
g15460 nor n15522 n15523 ; n15524
g15461 and n15513 n15524_not ; n15525
g15462 and n15513 n15525_not ; n15526
g15463 nor n15524 n15525 ; n15527
g15464 nor n15526 n15527 ; n15528
g15465 and n15438 n15450_not ; n15529
g15466 nor n15449 n15450 ; n15530
g15467 nor n15529 n15530 ; n15531
g15468 and n15422 n15434_not ; n15532
g15469 nor n15433 n15434 ; n15533
g15470 nor n15532 n15533 ; n15534
g15471 and n15250 n15415 ; n15535
g15472 nor n15416 n15535 ; n15536
g15473 and n3884 n12513 ; n15537
g15474 and n3967 n12516 ; n15538
g15475 and n4046 n12511 ; n15539
g15476 nor n15538 n15539 ; n15540
g15477 and n15537_not n15540 ; n15541
g15478 and n4050 n14177 ; n15542
g15479 and n15541 n15542_not ; n15543
g15480 and a[26] n15543_not ; n15544
g15481 and a[26] n15544_not ; n15545
g15482 nor n15543 n15544 ; n15546
g15483 nor n15545 n15546 ; n15547
g15484 and n15536 n15547_not ; n15548
g15485 and n15536 n15548_not ; n15549
g15486 nor n15547 n15548 ; n15550
g15487 nor n15549 n15550 ; n15551
g15488 and n15266 n15413 ; n15552
g15489 nor n15414 n15552 ; n15553
g15490 and n3457 n12522 ; n15554
g15491 and n3542 n12528 ; n15555
g15492 and n3606 n12525 ; n15556
g15493 nor n15555 n15556 ; n15557
g15494 and n15554_not n15557 ; n15558
g15495 and n3368 n14837 ; n15559
g15496 and n15558 n15559_not ; n15560
g15497 and a[29] n15560_not ; n15561
g15498 and a[29] n15561_not ; n15562
g15499 nor n15560 n15561 ; n15563
g15500 nor n15562 n15563 ; n15564
g15501 and n15553 n15564_not ; n15565
g15502 and n15553 n15565_not ; n15566
g15503 nor n15564 n15565 ; n15567
g15504 nor n15566 n15567 ; n15568
g15505 and n3884 n12511 ; n15569
g15506 and n3967 n12519 ; n15570
g15507 and n4046 n12516 ; n15571
g15508 nor n15570 n15571 ; n15572
g15509 and n15569_not n15572 ; n15573
g15510 and n4050 n14233_not ; n15574
g15511 and n15573 n15574_not ; n15575
g15512 and a[26] n15575_not ; n15576
g15513 and a[26] n15576_not ; n15577
g15514 nor n15575 n15576 ; n15578
g15515 nor n15577 n15578 ; n15579
g15516 nor n15568 n15579 ; n15580
g15517 nor n15565 n15580 ; n15581
g15518 nor n15551 n15581 ; n15582
g15519 nor n15548 n15582 ; n15583
g15520 nor n15534 n15583 ; n15584
g15521 and n15534 n15583 ; n15585
g15522 nor n15584 n15585 ; n15586
g15523 and n4694 n12502 ; n15587
g15524 and n4533 n12505 ; n15588
g15525 and n4604 n12370 ; n15589
g15526 nor n15588 n15589 ; n15590
g15527 and n15587_not n15590 ; n15591
g15528 and n4536 n13736_not ; n15592
g15529 and n15591 n15592_not ; n15593
g15530 and a[23] n15593_not ; n15594
g15531 and a[23] n15594_not ; n15595
g15532 nor n15593 n15594 ; n15596
g15533 nor n15595 n15596 ; n15597
g15534 and n15586 n15597_not ; n15598
g15535 nor n15584 n15598 ; n15599
g15536 nor n15531 n15599 ; n15600
g15537 and n15531 n15599 ; n15601
g15538 nor n15600 n15601 ; n15602
g15539 and n5496 n13518 ; n15603
g15540 and n4935 n12889 ; n15604
g15541 and n5407 n13491 ; n15605
g15542 nor n15604 n15605 ; n15606
g15543 and n15603_not n15606 ; n15607
g15544 and n4938 n13584 ; n15608
g15545 and n15607 n15608_not ; n15609
g15546 and a[20] n15609_not ; n15610
g15547 and a[20] n15610_not ; n15611
g15548 nor n15609 n15610 ; n15612
g15549 nor n15611 n15612 ; n15613
g15550 and n15602 n15613_not ; n15614
g15551 nor n15600 n15614 ; n15615
g15552 nor n15528 n15615 ; n15616
g15553 nor n15525 n15616 ; n15617
g15554 nor n15511 n15617 ; n15618
g15555 and n15511 n15617 ; n15619
g15556 nor n15618 n15619 ; n15620
g15557 and n6233 n13633 ; n15621
g15558 and n5663 n13597 ; n15622
g15559 and n5939 n13630 ; n15623
g15560 nor n15622 n15623 ; n15624
g15561 and n15621_not n15624 ; n15625
g15562 and n5666 n13929 ; n15626
g15563 and n15625 n15626_not ; n15627
g15564 and a[17] n15627_not ; n15628
g15565 and a[17] n15628_not ; n15629
g15566 nor n15627 n15628 ; n15630
g15567 nor n15629 n15630 ; n15631
g15568 and n15620 n15631_not ; n15632
g15569 nor n15618 n15632 ; n15633
g15570 nor n13438 n13845 ; n15634
g15571 and n6402 n13941 ; n15635
g15572 nor n15634 n15635 ; n15636
g15573 and n6397_not n15636 ; n15637
g15574 and n13951 n15636 ; n15638
g15575 nor n15637 n15638 ; n15639
g15576 and a[14] n15639_not ; n15640
g15577 and a[14]_not n15639 ; n15641
g15578 nor n15640 n15641 ; n15642
g15579 nor n15633 n15642 ; n15643
g15580 and n15472 n15484_not ; n15644
g15581 nor n15483 n15484 ; n15645
g15582 nor n15644 n15645 ; n15646
g15583 and n15633 n15642 ; n15647
g15584 nor n15643 n15647 ; n15648
g15585 and n15646_not n15648 ; n15649
g15586 nor n15643 n15649 ; n15650
g15587 and n15499_not n15502 ; n15651
g15588 nor n15503 n15651 ; n15652
g15589 and n15650_not n15652 ; n15653
g15590 nor n15646 n15649 ; n15654
g15591 and n15648 n15649_not ; n15655
g15592 nor n15654 n15655 ; n15656
g15593 and n15620 n15632_not ; n15657
g15594 nor n15631 n15632 ; n15658
g15595 nor n15657 n15658 ; n15659
g15596 and n15528 n15615 ; n15660
g15597 nor n15616 n15660 ; n15661
g15598 and n6233 n13630 ; n15662
g15599 and n5663 n13515 ; n15663
g15600 and n5939 n13597 ; n15664
g15601 nor n15663 n15664 ; n15665
g15602 and n15662_not n15665 ; n15666
g15603 and n5666 n13976 ; n15667
g15604 and n15666 n15667_not ; n15668
g15605 and a[17] n15668_not ; n15669
g15606 and a[17] n15669_not ; n15670
g15607 nor n15668 n15669 ; n15671
g15608 nor n15670 n15671 ; n15672
g15609 and n15661 n15672_not ; n15673
g15610 and n15661 n15673_not ; n15674
g15611 nor n15672 n15673 ; n15675
g15612 nor n15674 n15675 ; n15676
g15613 and n15602 n15614_not ; n15677
g15614 nor n15613 n15614 ; n15678
g15615 nor n15677 n15678 ; n15679
g15616 and n15586 n15598_not ; n15680
g15617 nor n15597 n15598 ; n15681
g15618 nor n15680 n15681 ; n15682
g15619 and n15551 n15581 ; n15683
g15620 nor n15582 n15683 ; n15684
g15621 and n4694 n12370 ; n15685
g15622 and n4533 n12508 ; n15686
g15623 and n4604 n12505 ; n15687
g15624 nor n15686 n15687 ; n15688
g15625 and n15685_not n15688 ; n15689
g15626 and n4536 n13748_not ; n15690
g15627 and n15689 n15690_not ; n15691
g15628 and a[23] n15691_not ; n15692
g15629 and a[23] n15692_not ; n15693
g15630 nor n15691 n15692 ; n15694
g15631 nor n15693 n15694 ; n15695
g15632 and n15684 n15695_not ; n15696
g15633 and n15684 n15696_not ; n15697
g15634 nor n15695 n15696 ; n15698
g15635 nor n15697 n15698 ; n15699
g15636 nor n15568 n15580 ; n15700
g15637 nor n15579 n15580 ; n15701
g15638 nor n15700 n15701 ; n15702
g15639 nor n15371 n15374 ; n15703
g15640 and n15372_not n15375 ; n15704
g15641 nor n15703 n15704 ; n15705
g15642 nor n12623 n12626 ; n15706
g15643 and n12624_not n12627 ; n15707
g15644 nor n15706 n15707 ; n15708
g15645 and n75 n15708_not ; n15709
g15646 and n3020 n12540 ; n15710
g15647 and n3023 n12546 ; n15711
g15648 and n3028 n12543 ; n15712
g15649 nor n15711 n15712 ; n15713
g15650 and n15710_not n15713 ; n15714
g15651 and n15709_not n15714 ; n15715
g15652 nor n15705 n15715 ; n15716
g15653 nor n15705 n15716 ; n15717
g15654 nor n15715 n15716 ; n15718
g15655 nor n15717 n15718 ; n15719
g15656 nor n15367 n15370 ; n15720
g15657 and n15368_not n15371 ; n15721
g15658 nor n15720 n15721 ; n15722
g15659 and n12619 n12621_not ; n15723
g15660 nor n12622 n15723 ; n15724
g15661 and n75 n15724 ; n15725
g15662 and n3020 n12543 ; n15726
g15663 and n3023 n12549 ; n15727
g15664 and n3028 n12546 ; n15728
g15665 nor n15727 n15728 ; n15729
g15666 and n15726_not n15729 ; n15730
g15667 and n15725_not n15730 ; n15731
g15668 nor n15722 n15731 ; n15732
g15669 nor n15722 n15732 ; n15733
g15670 nor n15731 n15732 ; n15734
g15671 nor n15733 n15734 ; n15735
g15672 nor n15363 n15366 ; n15736
g15673 and n15364_not n15367 ; n15737
g15674 nor n15736 n15737 ; n15738
g15675 and n289_not n12830 ; n15739
g15676 and n395_not n15739 ; n15740
g15677 and n173_not n15740 ; n15741
g15678 and n306_not n15741 ; n15742
g15679 and n270_not n15742 ; n15743
g15680 and n2784 n3162 ; n15744
g15681 and n2807 n15744 ; n15745
g15682 and n2262 n15745 ; n15746
g15683 and n2091 n15746 ; n15747
g15684 and n688 n15747 ; n15748
g15685 and n4815 n15748 ; n15749
g15686 and n14386 n15749 ; n15750
g15687 and n15743 n15750 ; n15751
g15688 and n288 n15751 ; n15752
g15689 and n356 n15752 ; n15753
g15690 and n116 n15753 ; n15754
g15691 and n149_not n15754 ; n15755
g15692 and n396_not n15755 ; n15756
g15693 and n167_not n15756 ; n15757
g15694 and n99_not n15757 ; n15758
g15695 and n237_not n15758 ; n15759
g15696 and n3020 n12549 ; n15760
g15697 and n3028 n12552 ; n15761
g15698 and n3023 n12555 ; n15762
g15699 and n12611 n12613_not ; n15763
g15700 nor n12614 n15763 ; n15764
g15701 and n75 n15764 ; n15765
g15702 nor n15762 n15765 ; n15766
g15703 and n15761_not n15766 ; n15767
g15704 and n15760_not n15767 ; n15768
g15705 nor n15759 n15768 ; n15769
g15706 and n1073 n3042 ; n15770
g15707 and n2704 n15770 ; n15771
g15708 and n2808 n15771 ; n15772
g15709 and n2422 n15772 ; n15773
g15710 and n13221 n15773 ; n15774
g15711 and n6026 n15774 ; n15775
g15712 and n1039 n15775 ; n15776
g15713 and n556 n15776 ; n15777
g15714 and n230 n15777 ; n15778
g15715 and n454 n15778 ; n15779
g15716 and n301_not n15779 ; n15780
g15717 and n1101_not n15780 ; n15781
g15718 and n716_not n15781 ; n15782
g15719 and n99_not n15782 ; n15783
g15720 and n86_not n15783 ; n15784
g15721 and n429_not n15784 ; n15785
g15722 and n3020 n12552 ; n15786
g15723 and n3028 n12555 ; n15787
g15724 and n3023 n12558 ; n15788
g15725 nor n12607 n12610 ; n15789
g15726 and n12608_not n12611 ; n15790
g15727 nor n15789 n15790 ; n15791
g15728 and n75 n15791_not ; n15792
g15729 nor n15788 n15792 ; n15793
g15730 and n15787_not n15793 ; n15794
g15731 and n15786_not n15794 ; n15795
g15732 nor n15785 n15795 ; n15796
g15733 and n2607 n3987 ; n15797
g15734 and n1604 n15797 ; n15798
g15735 and n1754 n15798 ; n15799
g15736 and n2555 n15799 ; n15800
g15737 and n15330 n15800 ; n15801
g15738 and n874 n15801 ; n15802
g15739 and n1475 n15802 ; n15803
g15740 and n4295 n15803 ; n15804
g15741 and n1040 n15804 ; n15805
g15742 and n281_not n15805 ; n15806
g15743 and n641_not n15806 ; n15807
g15744 and n170_not n15807 ; n15808
g15745 and n657_not n15808 ; n15809
g15746 and n771_not n15809 ; n15810
g15747 and n3020 n12555 ; n15811
g15748 and n3028 n12558 ; n15812
g15749 and n3023 n12561 ; n15813
g15750 nor n12603 n12606 ; n15814
g15751 and n12604_not n12607 ; n15815
g15752 nor n15814 n15815 ; n15816
g15753 and n75 n15816_not ; n15817
g15754 nor n15813 n15817 ; n15818
g15755 and n15812_not n15818 ; n15819
g15756 and n15811_not n15819 ; n15820
g15757 nor n15810 n15820 ; n15821
g15758 and n202 n877 ; n15822
g15759 and n364_not n15822 ; n15823
g15760 and n339_not n15823 ; n15824
g15761 and n493_not n15824 ; n15825
g15762 and n225_not n15825 ; n15826
g15763 and n1272 n1586 ; n15827
g15764 and n12428 n15827 ; n15828
g15765 and n3219 n15828 ; n15829
g15766 and n3415 n15829 ; n15830
g15767 and n6769 n15830 ; n15831
g15768 and n6707 n15831 ; n15832
g15769 and n1916 n15832 ; n15833
g15770 and n1475 n15833 ; n15834
g15771 and n1531 n15834 ; n15835
g15772 and n15826 n15835 ; n15836
g15773 and n509_not n15836 ; n15837
g15774 and n352_not n15837 ; n15838
g15775 and n461_not n15838 ; n15839
g15776 and n689_not n15839 ; n15840
g15777 and n99_not n15840 ; n15841
g15778 and n277_not n15841 ; n15842
g15779 and n3020 n12558 ; n15843
g15780 and n3028 n12561 ; n15844
g15781 and n3023 n12564 ; n15845
g15782 and n12599 n12601_not ; n15846
g15783 nor n12602 n15846 ; n15847
g15784 and n75 n15847 ; n15848
g15785 nor n15845 n15848 ; n15849
g15786 and n15844_not n15849 ; n15850
g15787 and n15843_not n15850 ; n15851
g15788 nor n15842 n15851 ; n15852
g15789 nor n374 n505 ; n15853
g15790 and n1203_not n15853 ; n15854
g15791 and n1391 n15854 ; n15855
g15792 and n690 n15855 ; n15856
g15793 and n4101 n15856 ; n15857
g15794 and n3159 n15857 ; n15858
g15795 and n6604 n15858 ; n15859
g15796 and n1522 n15859 ; n15860
g15797 and n602_not n15860 ; n15861
g15798 and n239_not n15861 ; n15862
g15799 and n715_not n15862 ; n15863
g15800 and n167_not n15863 ; n15864
g15801 and n338_not n15864 ; n15865
g15802 and n295_not n15865 ; n15866
g15803 and n249_not n15866 ; n15867
g15804 and n2209 n14518 ; n15868
g15805 and n4011 n15868 ; n15869
g15806 and n5190 n15869 ; n15870
g15807 and n6707 n15870 ; n15871
g15808 and n3990 n15871 ; n15872
g15809 and n2573 n15872 ; n15873
g15810 and n937 n15873 ; n15874
g15811 and n193 n15874 ; n15875
g15812 and n570 n15875 ; n15876
g15813 and n518_not n15876 ; n15877
g15814 and n673_not n15877 ; n15878
g15815 and n127_not n15878 ; n15879
g15816 and n358_not n15879 ; n15880
g15817 and n777_not n12711 ; n15881
g15818 and n81_not n15881 ; n15882
g15819 and n1274 n2742 ; n15883
g15820 and n15882 n15883 ; n15884
g15821 and n6517 n15884 ; n15885
g15822 and n14210 n15885 ; n15886
g15823 and n2703 n15886 ; n15887
g15824 and n15880 n15887 ; n15888
g15825 and n1915 n15888 ; n15889
g15826 and n1129 n15889 ; n15890
g15827 and n2583 n15890 ; n15891
g15828 and n202 n15891 ; n15892
g15829 and n15867 n15892 ; n15893
g15830 and n353_not n15893 ; n15894
g15831 and n151_not n15894 ; n15895
g15832 and n495_not n15895 ; n15896
g15833 and n375_not n15896 ; n15897
g15834 and n1104_not n15897 ; n15898
g15835 and n371_not n15898 ; n15899
g15836 and n3020 n12561 ; n15900
g15837 and n3028 n12564 ; n15901
g15838 and n3023 n12567 ; n15902
g15839 nor n12595 n12598 ; n15903
g15840 and n12596_not n12599 ; n15904
g15841 nor n15903 n15904 ; n15905
g15842 and n75 n15905_not ; n15906
g15843 nor n15902 n15906 ; n15907
g15844 and n15901_not n15907 ; n15908
g15845 and n15900_not n15908 ; n15909
g15846 nor n15899 n15909 ; n15910
g15847 and n12812 n13249 ; n15911
g15848 and n14572 n15911 ; n15912
g15849 and n247 n15912 ; n15913
g15850 and n622 n15913 ; n15914
g15851 and n1264 n15914 ; n15915
g15852 and n1183 n15915 ; n15916
g15853 and n1063 n15916 ; n15917
g15854 and n1781 n15917 ; n15918
g15855 and n2467 n15918 ; n15919
g15856 and n634 n15919 ; n15920
g15857 and n355_not n15920 ; n15921
g15858 and n689_not n15921 ; n15922
g15859 and n791_not n15922 ; n15923
g15860 and n394_not n15923 ; n15924
g15861 and n1798 n2442 ; n15925
g15862 and n2022 n15925 ; n15926
g15863 and n12805 n15926 ; n15927
g15864 and n13041 n15927 ; n15928
g15865 and n15924 n15928 ; n15929
g15866 and n731 n15929 ; n15930
g15867 and n978 n15930 ; n15931
g15868 and n236_not n15931 ; n15932
g15869 and n1246_not n15932 ; n15933
g15870 and n602_not n15933 ; n15934
g15871 and n400_not n15934 ; n15935
g15872 and n192_not n15935 ; n15936
g15873 and n537_not n15936 ; n15937
g15874 and n170_not n15937 ; n15938
g15875 and n3020 n12564 ; n15939
g15876 and n3028 n12567 ; n15940
g15877 and n3023 n12571 ; n15941
g15878 nor n12592 n12594 ; n15942
g15879 and n12569_not n12595 ; n15943
g15880 nor n15942 n15943 ; n15944
g15881 and n75 n15944_not ; n15945
g15882 nor n15941 n15945 ; n15946
g15883 and n15940_not n15946 ; n15947
g15884 and n15939_not n15947 ; n15948
g15885 nor n15938 n15948 ; n15949
g15886 and n3160 n3391 ; n15950
g15887 and n1011_not n15950 ; n15951
g15888 and n168_not n15951 ; n15952
g15889 and n492_not n15952 ; n15953
g15890 and n121_not n13671 ; n15954
g15891 and n825_not n15954 ; n15955
g15892 and n173_not n15955 ; n15956
g15893 and n14476 n15956 ; n15957
g15894 and n15953 n15957 ; n15958
g15895 and n471 n15958 ; n15959
g15896 and n1009 n15959 ; n15960
g15897 and n2443 n15960 ; n15961
g15898 and n827 n15961 ; n15962
g15899 and n746_not n15962 ; n15963
g15900 and n154_not n15963 ; n15964
g15901 and n637_not n15964 ; n15965
g15902 and n302_not n15965 ; n15966
g15903 and n274_not n15966 ; n15967
g15904 and n466_not n15967 ; n15968
g15905 and n623_not n15968 ; n15969
g15906 and n363_not n15969 ; n15970
g15907 and n1388 n2192 ; n15971
g15908 and n1693 n15971 ; n15972
g15909 and n4819 n15972 ; n15973
g15910 and n459 n15973 ; n15974
g15911 and n1549 n15974 ; n15975
g15912 and n2360 n15975 ; n15976
g15913 and n1131 n15976 ; n15977
g15914 and n15970 n15977 ; n15978
g15915 and n1253 n15978 ; n15979
g15916 and n135_not n15979 ; n15980
g15917 and n641_not n15980 ; n15981
g15918 and n417_not n15981 ; n15982
g15919 and n496_not n15982 ; n15983
g15920 and n714_not n15983 ; n15984
g15921 and n3020 n12567 ; n15985
g15922 and n3028 n12571 ; n15986
g15923 and n3023 n12574 ; n15987
g15924 and n12588 n12590_not ; n15988
g15925 nor n12591 n15988 ; n15989
g15926 and n75 n15989 ; n15990
g15927 nor n15987 n15990 ; n15991
g15928 and n15986_not n15991 ; n15992
g15929 and n15985_not n15992 ; n15993
g15930 nor n15984 n15993 ; n15994
g15931 and n2625 n3148 ; n15995
g15932 and n595 n15995 ; n15996
g15933 and n6565 n15996 ; n15997
g15934 and n5304 n15997 ; n15998
g15935 and n3205 n15998 ; n15999
g15936 and n13210 n15999 ; n16000
g15937 and n13135 n16000 ; n16001
g15938 and n3912 n16001 ; n16002
g15939 and n1916 n16002 ; n16003
g15940 and n2073 n16003 ; n16004
g15941 and n150_not n16004 ; n16005
g15942 and n563_not n16005 ; n16006
g15943 and n716_not n16006 ; n16007
g15944 and n468_not n16007 ; n16008
g15945 and n3020 n12571 ; n16009
g15946 and n3028 n12574 ; n16010
g15947 and n3023 n12577 ; n16011
g15948 and n12584 n12586_not ; n16012
g15949 nor n12587 n16012 ; n16013
g15950 and n75 n16013 ; n16014
g15951 nor n16011 n16014 ; n16015
g15952 and n16010_not n16015 ; n16016
g15953 and n16009_not n16016 ; n16017
g15954 nor n16008 n16017 ; n16018
g15955 nor n150 n713 ; n16019
g15956 and n589_not n16019 ; n16020
g15957 and n1409 n16020 ; n16021
g15958 and n1103 n16021 ; n16022
g15959 and n877 n16022 ; n16023
g15960 and n808 n16023 ; n16024
g15961 and n1480 n16024 ; n16025
g15962 and n731 n16025 ; n16026
g15963 and n111_not n16026 ; n16027
g15964 and n327_not n16027 ; n16028
g15965 and n430_not n16028 ; n16029
g15966 and n293_not n16029 ; n16030
g15967 and n429_not n16030 ; n16031
g15968 and n2992 n12785 ; n16032
g15969 and n658 n16032 ; n16033
g15970 and n3409 n16033 ; n16034
g15971 and n16031 n16034 ; n16035
g15972 and n14498 n16035 ; n16036
g15973 and n15337 n16036 ; n16037
g15974 and n5085 n16037 ; n16038
g15975 and n1247 n16038 ; n16039
g15976 and n418 n16039 ; n16040
g15977 and n328_not n16040 ; n16041
g15978 and n511_not n16041 ; n16042
g15979 and n147_not n16042 ; n16043
g15980 and n292_not n16043 ; n16044
g15981 and n513_not n16044 ; n16045
g15982 and n395_not n16045 ; n16046
g15983 and n716_not n16046 ; n16047
g15984 and n436_not n16047 ; n16048
g15985 and n222_not n16048 ; n16049
g15986 and n1160 n2191 ; n16050
g15987 and n752_not n16050 ; n16051
g15988 and n239_not n16051 ; n16052
g15989 and n146_not n16052 ; n16053
g15990 and n452_not n16053 ; n16054
g15991 and n161_not n16054 ; n16055
g15992 and n2007 n3128 ; n16056
g15993 and n13268 n16056 ; n16057
g15994 and n3905 n16057 ; n16058
g15995 and n790 n16058 ; n16059
g15996 and n15826 n16059 ; n16060
g15997 and n16055 n16060 ; n16061
g15998 and n282 n16061 ; n16062
g15999 and n827 n16062 ; n16063
g16000 and n107_not n16063 ; n16064
g16001 and n326_not n16064 ; n16065
g16002 and n81_not n16065 ; n16066
g16003 and n231_not n16066 ; n16067
g16004 and n1409 n1644 ; n16068
g16005 and n2441 n16068 ; n16069
g16006 and n2172 n16069 ; n16070
g16007 and n3771 n16070 ; n16071
g16008 and n2072 n16071 ; n16072
g16009 and n6662 n16072 ; n16073
g16010 and n2112 n16073 ; n16074
g16011 and n2346 n16074 ; n16075
g16012 and n16067 n16075 ; n16076
g16013 and n746_not n16076 ; n16077
g16014 and n292_not n16077 ; n16078
g16015 and n192_not n16078 ; n16079
g16016 and n173_not n16079 ; n16080
g16017 and n436_not n16080 ; n16081
g16018 and n3020 n12577 ; n16082
g16019 and n12577 n12581 ; n16083
g16020 nor n12577 n12581 ; n16084
g16021 nor n16083 n16084 ; n16085
g16022 and n75 n16085_not ; n16086
g16023 and n3028 n12581_not ; n16087
g16024 nor n16086 n16087 ; n16088
g16025 and n16082_not n16088 ; n16089
g16026 nor n16081 n16089 ; n16090
g16027 and n16049_not n16090 ; n16091
g16028 and n12574_not n16083 ; n16092
g16029 and n12574 n16083_not ; n16093
g16030 nor n16092 n16093 ; n16094
g16031 and n75 n16094_not ; n16095
g16032 and n3020 n12574 ; n16096
g16033 and n3023 n12581_not ; n16097
g16034 and n3028 n12577 ; n16098
g16035 nor n16097 n16098 ; n16099
g16036 and n16096_not n16099 ; n16100
g16037 and n16095_not n16100 ; n16101
g16038 and n16049 n16090_not ; n16102
g16039 nor n16091 n16102 ; n16103
g16040 and n16101_not n16103 ; n16104
g16041 nor n16091 n16104 ; n16105
g16042 nor n16008 n16018 ; n16106
g16043 nor n16017 n16018 ; n16107
g16044 nor n16106 n16107 ; n16108
g16045 nor n16105 n16108 ; n16109
g16046 nor n16018 n16109 ; n16110
g16047 nor n15984 n15994 ; n16111
g16048 nor n15993 n15994 ; n16112
g16049 nor n16111 n16112 ; n16113
g16050 nor n16110 n16113 ; n16114
g16051 nor n15994 n16114 ; n16115
g16052 nor n15938 n15949 ; n16116
g16053 nor n15948 n15949 ; n16117
g16054 nor n16116 n16117 ; n16118
g16055 nor n16115 n16118 ; n16119
g16056 nor n15949 n16119 ; n16120
g16057 nor n15899 n15910 ; n16121
g16058 nor n15909 n15910 ; n16122
g16059 nor n16121 n16122 ; n16123
g16060 nor n16120 n16123 ; n16124
g16061 nor n15910 n16124 ; n16125
g16062 nor n15842 n15852 ; n16126
g16063 nor n15851 n15852 ; n16127
g16064 nor n16126 n16127 ; n16128
g16065 nor n16125 n16128 ; n16129
g16066 nor n15852 n16129 ; n16130
g16067 nor n15810 n15821 ; n16131
g16068 nor n15820 n15821 ; n16132
g16069 nor n16131 n16132 ; n16133
g16070 nor n16130 n16133 ; n16134
g16071 nor n15821 n16134 ; n16135
g16072 nor n15785 n15796 ; n16136
g16073 nor n15795 n15796 ; n16137
g16074 nor n16136 n16137 ; n16138
g16075 nor n16135 n16138 ; n16139
g16076 nor n15796 n16139 ; n16140
g16077 nor n15759 n15769 ; n16141
g16078 nor n15768 n15769 ; n16142
g16079 nor n16141 n16142 ; n16143
g16080 nor n16140 n16143 ; n16144
g16081 nor n15769 n16144 ; n16145
g16082 nor n15738 n16145 ; n16146
g16083 and n15738 n16145 ; n16147
g16084 nor n16146 n16147 ; n16148
g16085 and n3457 n12537 ; n16149
g16086 and n3542 n12543 ; n16150
g16087 and n3606 n12540 ; n16151
g16088 nor n16150 n16151 ; n16152
g16089 and n16149_not n16152 ; n16153
g16090 and n3368_not n16153 ; n16154
g16091 and n15385 n16153 ; n16155
g16092 nor n16154 n16155 ; n16156
g16093 and a[29] n16156_not ; n16157
g16094 and a[29]_not n16156 ; n16158
g16095 nor n16157 n16158 ; n16159
g16096 and n16148 n16159_not ; n16160
g16097 nor n16146 n16160 ; n16161
g16098 nor n15735 n16161 ; n16162
g16099 nor n15732 n16162 ; n16163
g16100 nor n15719 n16163 ; n16164
g16101 nor n15716 n16164 ; n16165
g16102 and n15382 n15392 ; n16166
g16103 nor n15393 n16166 ; n16167
g16104 and n16165_not n16167 ; n16168
g16105 and n16165 n16167_not ; n16169
g16106 nor n16168 n16169 ; n16170
g16107 and n3457 n12528 ; n16171
g16108 and n3542 n12534 ; n16172
g16109 and n3606 n12531 ; n16173
g16110 nor n16172 n16173 ; n16174
g16111 and n16171_not n16174 ; n16175
g16112 and n3368 n15003_not ; n16176
g16113 and n16175 n16176_not ; n16177
g16114 and a[29] n16177_not ; n16178
g16115 and a[29] n16178_not ; n16179
g16116 nor n16177 n16178 ; n16180
g16117 nor n16179 n16180 ; n16181
g16118 and n16170 n16181_not ; n16182
g16119 nor n16168 n16182 ; n16183
g16120 and n15400_not n15411 ; n16184
g16121 nor n15412 n16184 ; n16185
g16122 and n16183_not n16185 ; n16186
g16123 and n16183 n16185_not ; n16187
g16124 nor n16186 n16187 ; n16188
g16125 and n3884 n12516 ; n16189
g16126 and n3967 n12522 ; n16190
g16127 and n4046 n12519 ; n16191
g16128 nor n16190 n16191 ; n16192
g16129 and n16189_not n16192 ; n16193
g16130 and n4050 n14443_not ; n16194
g16131 and n16193 n16194_not ; n16195
g16132 and a[26] n16195_not ; n16196
g16133 and a[26] n16196_not ; n16197
g16134 nor n16195 n16196 ; n16198
g16135 nor n16197 n16198 ; n16199
g16136 and n16188 n16199_not ; n16200
g16137 nor n16186 n16200 ; n16201
g16138 nor n15702 n16201 ; n16202
g16139 and n15702 n16201 ; n16203
g16140 nor n16202 n16203 ; n16204
g16141 and n4694 n12505 ; n16205
g16142 and n4533 n12513 ; n16206
g16143 and n4604 n12508 ; n16207
g16144 nor n16206 n16207 ; n16208
g16145 and n16205_not n16208 ; n16209
g16146 and n4536 n14051_not ; n16210
g16147 and n16209 n16210_not ; n16211
g16148 and a[23] n16211_not ; n16212
g16149 and a[23] n16212_not ; n16213
g16150 nor n16211 n16212 ; n16214
g16151 nor n16213 n16214 ; n16215
g16152 and n16204 n16215_not ; n16216
g16153 nor n16202 n16216 ; n16217
g16154 nor n15699 n16217 ; n16218
g16155 nor n15696 n16218 ; n16219
g16156 nor n15682 n16219 ; n16220
g16157 and n15682 n16219 ; n16221
g16158 nor n16220 n16221 ; n16222
g16159 and n5496 n13491 ; n16223
g16160 and n4935 n12769 ; n16224
g16161 and n5407 n12889 ; n16225
g16162 nor n16224 n16225 ; n16226
g16163 and n16223_not n16226 ; n16227
g16164 and n4938 n13503_not ; n16228
g16165 and n16227 n16228_not ; n16229
g16166 and a[20] n16229_not ; n16230
g16167 and a[20] n16230_not ; n16231
g16168 nor n16229 n16230 ; n16232
g16169 nor n16231 n16232 ; n16233
g16170 and n16222 n16233_not ; n16234
g16171 nor n16220 n16234 ; n16235
g16172 nor n15679 n16235 ; n16236
g16173 and n15679 n16235 ; n16237
g16174 nor n16236 n16237 ; n16238
g16175 and n6233 n13597 ; n16239
g16176 and n5663 n13521 ; n16240
g16177 and n5939 n13515 ; n16241
g16178 nor n16240 n16241 ; n16242
g16179 and n16239_not n16242 ; n16243
g16180 and n5666 n13612_not ; n16244
g16181 and n16243 n16244_not ; n16245
g16182 and a[17] n16245_not ; n16246
g16183 and a[17] n16246_not ; n16247
g16184 nor n16245 n16246 ; n16248
g16185 nor n16247 n16248 ; n16249
g16186 and n16238 n16249_not ; n16250
g16187 nor n16236 n16250 ; n16251
g16188 nor n15676 n16251 ; n16252
g16189 nor n15673 n16252 ; n16253
g16190 nor n15659 n16253 ; n16254
g16191 and n15659 n16253 ; n16255
g16192 nor n16254 n16255 ; n16256
g16193 and n7101 n13438_not ; n16257
g16194 and n6402 n13627_not ; n16258
g16195 and n6951 n13941 ; n16259
g16196 nor n16258 n16259 ; n16260
g16197 and n16257_not n16260 ; n16261
g16198 and n6397 n14028 ; n16262
g16199 and n16261 n16262_not ; n16263
g16200 and a[14] n16263_not ; n16264
g16201 and a[14] n16264_not ; n16265
g16202 nor n16263 n16264 ; n16266
g16203 nor n16265 n16266 ; n16267
g16204 and n16256 n16267_not ; n16268
g16205 nor n16254 n16268 ; n16269
g16206 nor n15656 n16269 ; n16270
g16207 and n15656 n16269 ; n16271
g16208 nor n16270 n16271 ; n16272
g16209 and n16256 n16268_not ; n16273
g16210 nor n16267 n16268 ; n16274
g16211 nor n16273 n16274 ; n16275
g16212 and n16238 n16250_not ; n16276
g16213 nor n16249 n16250 ; n16277
g16214 nor n16276 n16277 ; n16278
g16215 and n16222 n16234_not ; n16279
g16216 nor n16233 n16234 ; n16280
g16217 nor n16279 n16280 ; n16281
g16218 and n15699 n16217 ; n16282
g16219 nor n16218 n16282 ; n16283
g16220 and n5496 n12889 ; n16284
g16221 and n4935 n12502 ; n16285
g16222 and n5407 n12769 ; n16286
g16223 nor n16285 n16286 ; n16287
g16224 and n16284_not n16287 ; n16288
g16225 and n4938 n12895 ; n16289
g16226 and n16288 n16289_not ; n16290
g16227 and a[20] n16290_not ; n16291
g16228 and a[20] n16291_not ; n16292
g16229 nor n16290 n16291 ; n16293
g16230 nor n16292 n16293 ; n16294
g16231 and n16283 n16294_not ; n16295
g16232 and n16283 n16295_not ; n16296
g16233 nor n16294 n16295 ; n16297
g16234 nor n16296 n16297 ; n16298
g16235 and n16204 n16216_not ; n16299
g16236 nor n16215 n16216 ; n16300
g16237 nor n16299 n16300 ; n16301
g16238 and n16188 n16200_not ; n16302
g16239 nor n16199 n16200 ; n16303
g16240 nor n16302 n16303 ; n16304
g16241 and n16170 n16182_not ; n16305
g16242 nor n16181 n16182 ; n16306
g16243 nor n16305 n16306 ; n16307
g16244 and n3884 n12519 ; n16308
g16245 and n3967 n12525 ; n16309
g16246 and n4046 n12522 ; n16310
g16247 nor n16309 n16310 ; n16311
g16248 and n16308_not n16311 ; n16312
g16249 and n4050 n14454 ; n16313
g16250 and n16312 n16313_not ; n16314
g16251 and a[26] n16314_not ; n16315
g16252 and a[26] n16315_not ; n16316
g16253 nor n16314 n16315 ; n16317
g16254 nor n16316 n16317 ; n16318
g16255 nor n16307 n16318 ; n16319
g16256 nor n16307 n16319 ; n16320
g16257 nor n16318 n16319 ; n16321
g16258 nor n16320 n16321 ; n16322
g16259 and n15719 n16163 ; n16323
g16260 nor n16164 n16323 ; n16324
g16261 and n3457 n12531 ; n16325
g16262 and n3542 n12537 ; n16326
g16263 and n3606 n12534 ; n16327
g16264 nor n16326 n16327 ; n16328
g16265 and n16325_not n16328 ; n16329
g16266 and n3368 n15255 ; n16330
g16267 and n16329 n16330_not ; n16331
g16268 and a[29] n16331_not ; n16332
g16269 and a[29] n16332_not ; n16333
g16270 nor n16331 n16332 ; n16334
g16271 nor n16333 n16334 ; n16335
g16272 and n16324 n16335_not ; n16336
g16273 and n16324 n16336_not ; n16337
g16274 nor n16335 n16336 ; n16338
g16275 nor n16337 n16338 ; n16339
g16276 and n3967 n12528 ; n16340
g16277 and n4046 n12525 ; n16341
g16278 and n3884 n12522 ; n16342
g16279 nor n16341 n16342 ; n16343
g16280 and n16340_not n16343 ; n16344
g16281 and n4050 n14837 ; n16345
g16282 and n16344 n16345_not ; n16346
g16283 and a[26] n16346_not ; n16347
g16284 and a[26] n16347_not ; n16348
g16285 nor n16346 n16347 ; n16349
g16286 nor n16348 n16349 ; n16350
g16287 nor n16339 n16350 ; n16351
g16288 nor n16336 n16351 ; n16352
g16289 nor n16322 n16352 ; n16353
g16290 nor n16319 n16353 ; n16354
g16291 nor n16304 n16354 ; n16355
g16292 and n16304 n16354 ; n16356
g16293 nor n16355 n16356 ; n16357
g16294 and n4694 n12508 ; n16358
g16295 and n4533 n12511 ; n16359
g16296 and n4604 n12513 ; n16360
g16297 nor n16359 n16360 ; n16361
g16298 and n16358_not n16361 ; n16362
g16299 and n4536 n13863 ; n16363
g16300 and n16362 n16363_not ; n16364
g16301 and a[23] n16364_not ; n16365
g16302 and a[23] n16365_not ; n16366
g16303 nor n16364 n16365 ; n16367
g16304 nor n16366 n16367 ; n16368
g16305 and n16357 n16368_not ; n16369
g16306 nor n16355 n16369 ; n16370
g16307 nor n16301 n16370 ; n16371
g16308 and n16301 n16370 ; n16372
g16309 nor n16371 n16372 ; n16373
g16310 and n5496 n12769 ; n16374
g16311 and n4935 n12370 ; n16375
g16312 and n5407 n12502 ; n16376
g16313 nor n16375 n16376 ; n16377
g16314 and n16374_not n16377 ; n16378
g16315 and n4938 n12999 ; n16379
g16316 and n16378 n16379_not ; n16380
g16317 and a[20] n16380_not ; n16381
g16318 and a[20] n16381_not ; n16382
g16319 nor n16380 n16381 ; n16383
g16320 nor n16382 n16383 ; n16384
g16321 and n16373 n16384_not ; n16385
g16322 nor n16371 n16385 ; n16386
g16323 nor n16298 n16386 ; n16387
g16324 nor n16295 n16387 ; n16388
g16325 nor n16281 n16388 ; n16389
g16326 and n16281 n16388 ; n16390
g16327 nor n16389 n16390 ; n16391
g16328 and n6233 n13515 ; n16392
g16329 and n5663 n13518 ; n16393
g16330 and n5939 n13521 ; n16394
g16331 nor n16393 n16394 ; n16395
g16332 and n16392_not n16395 ; n16396
g16333 and n5666 n13541 ; n16397
g16334 and n16396 n16397_not ; n16398
g16335 and a[17] n16398_not ; n16399
g16336 and a[17] n16399_not ; n16400
g16337 nor n16398 n16399 ; n16401
g16338 nor n16400 n16401 ; n16402
g16339 and n16391 n16402_not ; n16403
g16340 nor n16389 n16403 ; n16404
g16341 nor n16278 n16404 ; n16405
g16342 and n16278 n16404 ; n16406
g16343 nor n16405 n16406 ; n16407
g16344 and n7101 n13627_not ; n16408
g16345 and n6402 n13630 ; n16409
g16346 and n6951 n13633 ; n16410
g16347 nor n16409 n16410 ; n16411
g16348 and n16408_not n16411 ; n16412
g16349 and n6397 n13654_not ; n16413
g16350 and n16412 n16413_not ; n16414
g16351 and a[14] n16414_not ; n16415
g16352 and a[14] n16415_not ; n16416
g16353 nor n16414 n16415 ; n16417
g16354 nor n16416 n16417 ; n16418
g16355 and n16407 n16418_not ; n16419
g16356 nor n16405 n16419 ; n16420
g16357 and n7101 n13941 ; n16421
g16358 and n6402 n13633 ; n16422
g16359 and n6951 n13627_not ; n16423
g16360 nor n16422 n16423 ; n16424
g16361 and n16421_not n16424 ; n16425
g16362 and n6397 n14136 ; n16426
g16363 and n16425 n16426_not ; n16427
g16364 and a[14] n16427_not ; n16428
g16365 and a[14] n16428_not ; n16429
g16366 nor n16427 n16428 ; n16430
g16367 nor n16429 n16430 ; n16431
g16368 nor n16420 n16431 ; n16432
g16369 and n15676 n16251 ; n16433
g16370 nor n16252 n16433 ; n16434
g16371 nor n16420 n16432 ; n16435
g16372 nor n16431 n16432 ; n16436
g16373 nor n16435 n16436 ; n16437
g16374 and n16434 n16437_not ; n16438
g16375 nor n16432 n16438 ; n16439
g16376 nor n16275 n16439 ; n16440
g16377 nor n16275 n16440 ; n16441
g16378 nor n16439 n16440 ; n16442
g16379 nor n16441 n16442 ; n16443
g16380 and n16391 n16403_not ; n16444
g16381 nor n16402 n16403 ; n16445
g16382 nor n16444 n16445 ; n16446
g16383 and n16298 n16386 ; n16447
g16384 nor n16387 n16447 ; n16448
g16385 and n6233 n13521 ; n16449
g16386 and n5663 n13491 ; n16450
g16387 and n5939 n13518 ; n16451
g16388 nor n16450 n16451 ; n16452
g16389 and n16449_not n16452 ; n16453
g16390 and n5666 n13909_not ; n16454
g16391 and n16453 n16454_not ; n16455
g16392 and a[17] n16455_not ; n16456
g16393 and a[17] n16456_not ; n16457
g16394 nor n16455 n16456 ; n16458
g16395 nor n16457 n16458 ; n16459
g16396 and n16448 n16459_not ; n16460
g16397 and n16448 n16460_not ; n16461
g16398 nor n16459 n16460 ; n16462
g16399 nor n16461 n16462 ; n16463
g16400 and n16373 n16385_not ; n16464
g16401 nor n16384 n16385 ; n16465
g16402 nor n16464 n16465 ; n16466
g16403 and n16357 n16369_not ; n16467
g16404 nor n16368 n16369 ; n16468
g16405 nor n16467 n16468 ; n16469
g16406 and n16322 n16352 ; n16470
g16407 nor n16353 n16470 ; n16471
g16408 and n4694 n12513 ; n16472
g16409 and n4533 n12516 ; n16473
g16410 and n4604 n12511 ; n16474
g16411 nor n16473 n16474 ; n16475
g16412 and n16472_not n16475 ; n16476
g16413 and n4536 n14177 ; n16477
g16414 and n16476 n16477_not ; n16478
g16415 and a[23] n16478_not ; n16479
g16416 and a[23] n16479_not ; n16480
g16417 nor n16478 n16479 ; n16481
g16418 nor n16480 n16481 ; n16482
g16419 and n16471 n16482_not ; n16483
g16420 and n16471 n16483_not ; n16484
g16421 nor n16482 n16483 ; n16485
g16422 nor n16484 n16485 ; n16486
g16423 nor n16339 n16351 ; n16487
g16424 nor n16350 n16351 ; n16488
g16425 nor n16487 n16488 ; n16489
g16426 and n15735 n16161 ; n16490
g16427 nor n16162 n16490 ; n16491
g16428 and n3457 n12534 ; n16492
g16429 and n3542 n12540 ; n16493
g16430 and n3606 n12537 ; n16494
g16431 nor n16493 n16494 ; n16495
g16432 and n16492_not n16495 ; n16496
g16433 and n3368 n15096_not ; n16497
g16434 and n16496 n16497_not ; n16498
g16435 and a[29] n16498_not ; n16499
g16436 and a[29] n16499_not ; n16500
g16437 nor n16498 n16499 ; n16501
g16438 nor n16500 n16501 ; n16502
g16439 and n16491 n16502_not ; n16503
g16440 and n16491 n16503_not ; n16504
g16441 nor n16502 n16503 ; n16505
g16442 nor n16504 n16505 ; n16506
g16443 and n4046 n12528 ; n16507
g16444 and n3884 n12525 ; n16508
g16445 and n3967 n12531 ; n16509
g16446 nor n16508 n16509 ; n16510
g16447 and n16507_not n16510 ; n16511
g16448 and n4050 n14608 ; n16512
g16449 and n16511 n16512_not ; n16513
g16450 and a[26] n16513_not ; n16514
g16451 and a[26] n16514_not ; n16515
g16452 nor n16513 n16514 ; n16516
g16453 nor n16515 n16516 ; n16517
g16454 nor n16506 n16517 ; n16518
g16455 nor n16503 n16518 ; n16519
g16456 nor n16489 n16519 ; n16520
g16457 and n16489 n16519 ; n16521
g16458 nor n16520 n16521 ; n16522
g16459 and n4694 n12511 ; n16523
g16460 and n4533 n12519 ; n16524
g16461 and n4604 n12516 ; n16525
g16462 nor n16524 n16525 ; n16526
g16463 and n16523_not n16526 ; n16527
g16464 and n4536 n14233_not ; n16528
g16465 and n16527 n16528_not ; n16529
g16466 and a[23] n16529_not ; n16530
g16467 and a[23] n16530_not ; n16531
g16468 nor n16529 n16530 ; n16532
g16469 nor n16531 n16532 ; n16533
g16470 and n16522 n16533_not ; n16534
g16471 nor n16520 n16534 ; n16535
g16472 nor n16486 n16535 ; n16536
g16473 nor n16483 n16536 ; n16537
g16474 nor n16469 n16537 ; n16538
g16475 and n16469 n16537 ; n16539
g16476 nor n16538 n16539 ; n16540
g16477 and n5496 n12502 ; n16541
g16478 and n4935 n12505 ; n16542
g16479 and n5407 n12370 ; n16543
g16480 nor n16542 n16543 ; n16544
g16481 and n16541_not n16544 ; n16545
g16482 and n4938 n13736_not ; n16546
g16483 and n16545 n16546_not ; n16547
g16484 and a[20] n16547_not ; n16548
g16485 and a[20] n16548_not ; n16549
g16486 nor n16547 n16548 ; n16550
g16487 nor n16549 n16550 ; n16551
g16488 and n16540 n16551_not ; n16552
g16489 nor n16538 n16552 ; n16553
g16490 nor n16466 n16553 ; n16554
g16491 and n16466 n16553 ; n16555
g16492 nor n16554 n16555 ; n16556
g16493 and n6233 n13518 ; n16557
g16494 and n5663 n12889 ; n16558
g16495 and n5939 n13491 ; n16559
g16496 nor n16558 n16559 ; n16560
g16497 and n16557_not n16560 ; n16561
g16498 and n5666 n13584 ; n16562
g16499 and n16561 n16562_not ; n16563
g16500 and a[17] n16563_not ; n16564
g16501 and a[17] n16564_not ; n16565
g16502 nor n16563 n16564 ; n16566
g16503 nor n16565 n16566 ; n16567
g16504 and n16556 n16567_not ; n16568
g16505 nor n16554 n16568 ; n16569
g16506 nor n16463 n16569 ; n16570
g16507 nor n16460 n16570 ; n16571
g16508 nor n16446 n16571 ; n16572
g16509 and n16446 n16571 ; n16573
g16510 nor n16572 n16573 ; n16574
g16511 and n7101 n13633 ; n16575
g16512 and n6402 n13597 ; n16576
g16513 and n6951 n13630 ; n16577
g16514 nor n16576 n16577 ; n16578
g16515 and n16575_not n16578 ; n16579
g16516 and n6397 n13929 ; n16580
g16517 and n16579 n16580_not ; n16581
g16518 and a[14] n16581_not ; n16582
g16519 and a[14] n16582_not ; n16583
g16520 nor n16581 n16582 ; n16584
g16521 nor n16583 n16584 ; n16585
g16522 and n16574 n16585_not ; n16586
g16523 nor n16572 n16586 ; n16587
g16524 nor n13438 n14424 ; n16588
g16525 and n7291 n13941 ; n16589
g16526 nor n16588 n16589 ; n16590
g16527 and n7294_not n16590 ; n16591
g16528 and n13951 n16590 ; n16592
g16529 nor n16591 n16592 ; n16593
g16530 and a[11] n16593_not ; n16594
g16531 and a[11]_not n16593 ; n16595
g16532 nor n16594 n16595 ; n16596
g16533 nor n16587 n16596 ; n16597
g16534 and n16407 n16419_not ; n16598
g16535 nor n16418 n16419 ; n16599
g16536 nor n16598 n16599 ; n16600
g16537 and n16587 n16596 ; n16601
g16538 nor n16597 n16601 ; n16602
g16539 and n16600_not n16602 ; n16603
g16540 nor n16597 n16603 ; n16604
g16541 and n16434_not n16437 ; n16605
g16542 nor n16438 n16605 ; n16606
g16543 and n16604_not n16606 ; n16607
g16544 nor n16600 n16603 ; n16608
g16545 and n16602 n16603_not ; n16609
g16546 nor n16608 n16609 ; n16610
g16547 and n16574 n16586_not ; n16611
g16548 nor n16585 n16586 ; n16612
g16549 nor n16611 n16612 ; n16613
g16550 and n16463 n16569 ; n16614
g16551 nor n16570 n16614 ; n16615
g16552 and n7101 n13630 ; n16616
g16553 and n6402 n13515 ; n16617
g16554 and n6951 n13597 ; n16618
g16555 nor n16617 n16618 ; n16619
g16556 and n16616_not n16619 ; n16620
g16557 and n6397 n13976 ; n16621
g16558 and n16620 n16621_not ; n16622
g16559 and a[14] n16622_not ; n16623
g16560 and a[14] n16623_not ; n16624
g16561 nor n16622 n16623 ; n16625
g16562 nor n16624 n16625 ; n16626
g16563 and n16615 n16626_not ; n16627
g16564 and n16615 n16627_not ; n16628
g16565 nor n16626 n16627 ; n16629
g16566 nor n16628 n16629 ; n16630
g16567 and n16556 n16568_not ; n16631
g16568 nor n16567 n16568 ; n16632
g16569 nor n16631 n16632 ; n16633
g16570 and n16540 n16552_not ; n16634
g16571 nor n16551 n16552 ; n16635
g16572 nor n16634 n16635 ; n16636
g16573 and n16486 n16535 ; n16637
g16574 nor n16536 n16637 ; n16638
g16575 and n5496 n12370 ; n16639
g16576 and n4935 n12508 ; n16640
g16577 and n5407 n12505 ; n16641
g16578 nor n16640 n16641 ; n16642
g16579 and n16639_not n16642 ; n16643
g16580 and n4938 n13748_not ; n16644
g16581 and n16643 n16644_not ; n16645
g16582 and a[20] n16645_not ; n16646
g16583 and a[20] n16646_not ; n16647
g16584 nor n16645 n16646 ; n16648
g16585 nor n16647 n16648 ; n16649
g16586 and n16638 n16649_not ; n16650
g16587 and n16638 n16650_not ; n16651
g16588 nor n16649 n16650 ; n16652
g16589 nor n16651 n16652 ; n16653
g16590 and n16522 n16534_not ; n16654
g16591 nor n16533 n16534 ; n16655
g16592 nor n16654 n16655 ; n16656
g16593 nor n16506 n16518 ; n16657
g16594 nor n16517 n16518 ; n16658
g16595 nor n16657 n16658 ; n16659
g16596 nor n16140 n16144 ; n16660
g16597 nor n16143 n16144 ; n16661
g16598 nor n16660 n16661 ; n16662
g16599 and n3457 n12540 ; n16663
g16600 and n3542 n12546 ; n16664
g16601 and n3606 n12543 ; n16665
g16602 nor n16664 n16665 ; n16666
g16603 and n16663_not n16666 ; n16667
g16604 and n3368_not n16667 ; n16668
g16605 and n15708 n16667 ; n16669
g16606 nor n16668 n16669 ; n16670
g16607 and a[29] n16670_not ; n16671
g16608 and a[29]_not n16670 ; n16672
g16609 nor n16671 n16672 ; n16673
g16610 nor n16662 n16673 ; n16674
g16611 nor n16135 n16139 ; n16675
g16612 nor n16138 n16139 ; n16676
g16613 nor n16675 n16676 ; n16677
g16614 and n3457 n12543 ; n16678
g16615 and n3542 n12549 ; n16679
g16616 and n3606 n12546 ; n16680
g16617 nor n16679 n16680 ; n16681
g16618 and n16678_not n16681 ; n16682
g16619 and n3368_not n16682 ; n16683
g16620 and n15724_not n16682 ; n16684
g16621 nor n16683 n16684 ; n16685
g16622 and a[29] n16685_not ; n16686
g16623 and a[29]_not n16685 ; n16687
g16624 nor n16686 n16687 ; n16688
g16625 nor n16677 n16688 ; n16689
g16626 nor n16130 n16134 ; n16690
g16627 nor n16133 n16134 ; n16691
g16628 nor n16690 n16691 ; n16692
g16629 and n3457 n12546 ; n16693
g16630 and n3542 n12552 ; n16694
g16631 and n3606 n12549 ; n16695
g16632 nor n16694 n16695 ; n16696
g16633 and n16693_not n16696 ; n16697
g16634 and n3368_not n16697 ; n16698
g16635 and n15356 n16697 ; n16699
g16636 nor n16698 n16699 ; n16700
g16637 and a[29] n16700_not ; n16701
g16638 and a[29]_not n16700 ; n16702
g16639 nor n16701 n16702 ; n16703
g16640 nor n16692 n16703 ; n16704
g16641 nor n16125 n16129 ; n16705
g16642 nor n16128 n16129 ; n16706
g16643 nor n16705 n16706 ; n16707
g16644 and n3457 n12549 ; n16708
g16645 and n3542 n12555 ; n16709
g16646 and n3606 n12552 ; n16710
g16647 nor n16709 n16710 ; n16711
g16648 and n16708_not n16711 ; n16712
g16649 and n3368_not n16712 ; n16713
g16650 and n15764_not n16712 ; n16714
g16651 nor n16713 n16714 ; n16715
g16652 and a[29] n16715_not ; n16716
g16653 and a[29]_not n16715 ; n16717
g16654 nor n16716 n16717 ; n16718
g16655 nor n16707 n16718 ; n16719
g16656 nor n16120 n16124 ; n16720
g16657 nor n16123 n16124 ; n16721
g16658 nor n16720 n16721 ; n16722
g16659 and n3457 n12552 ; n16723
g16660 and n3542 n12558 ; n16724
g16661 and n3606 n12555 ; n16725
g16662 nor n16724 n16725 ; n16726
g16663 and n16723_not n16726 ; n16727
g16664 and n3368_not n16727 ; n16728
g16665 and n15791 n16727 ; n16729
g16666 nor n16728 n16729 ; n16730
g16667 and a[29] n16730_not ; n16731
g16668 and a[29]_not n16730 ; n16732
g16669 nor n16731 n16732 ; n16733
g16670 nor n16722 n16733 ; n16734
g16671 and n3457 n12555 ; n16735
g16672 and n3542 n12561 ; n16736
g16673 and n3606 n12558 ; n16737
g16674 nor n16736 n16737 ; n16738
g16675 and n16735_not n16738 ; n16739
g16676 and n3368 n15816_not ; n16740
g16677 and n16739 n16740_not ; n16741
g16678 and a[29] n16741_not ; n16742
g16679 nor n16741 n16742 ; n16743
g16680 and a[29] n16742_not ; n16744
g16681 nor n16743 n16744 ; n16745
g16682 nor n16115 n16119 ; n16746
g16683 nor n16118 n16119 ; n16747
g16684 nor n16746 n16747 ; n16748
g16685 nor n16745 n16748 ; n16749
g16686 nor n16745 n16749 ; n16750
g16687 nor n16748 n16749 ; n16751
g16688 nor n16750 n16751 ; n16752
g16689 and n3457 n12558 ; n16753
g16690 and n3542 n12564 ; n16754
g16691 and n3606 n12561 ; n16755
g16692 nor n16754 n16755 ; n16756
g16693 and n16753_not n16756 ; n16757
g16694 and n3368 n15847 ; n16758
g16695 and n16757 n16758_not ; n16759
g16696 and a[29] n16759_not ; n16760
g16697 nor n16759 n16760 ; n16761
g16698 and a[29] n16760_not ; n16762
g16699 nor n16761 n16762 ; n16763
g16700 nor n16110 n16114 ; n16764
g16701 nor n16113 n16114 ; n16765
g16702 nor n16764 n16765 ; n16766
g16703 nor n16763 n16766 ; n16767
g16704 nor n16763 n16767 ; n16768
g16705 nor n16766 n16767 ; n16769
g16706 nor n16768 n16769 ; n16770
g16707 and n3457 n12561 ; n16771
g16708 and n3542 n12567 ; n16772
g16709 and n3606 n12564 ; n16773
g16710 nor n16772 n16773 ; n16774
g16711 and n16771_not n16774 ; n16775
g16712 and n3368 n15905_not ; n16776
g16713 and n16775 n16776_not ; n16777
g16714 and a[29] n16777_not ; n16778
g16715 nor n16777 n16778 ; n16779
g16716 and a[29] n16778_not ; n16780
g16717 nor n16779 n16780 ; n16781
g16718 nor n16105 n16109 ; n16782
g16719 nor n16108 n16109 ; n16783
g16720 nor n16782 n16783 ; n16784
g16721 nor n16781 n16784 ; n16785
g16722 nor n16781 n16785 ; n16786
g16723 nor n16784 n16785 ; n16787
g16724 nor n16786 n16787 ; n16788
g16725 and n3457 n12564 ; n16789
g16726 and n3542 n12571 ; n16790
g16727 and n3606 n12567 ; n16791
g16728 nor n16790 n16791 ; n16792
g16729 and n16789_not n16792 ; n16793
g16730 and n3368 n15944_not ; n16794
g16731 and n16793 n16794_not ; n16795
g16732 and a[29] n16795_not ; n16796
g16733 nor n16795 n16796 ; n16797
g16734 and a[29] n16796_not ; n16798
g16735 nor n16797 n16798 ; n16799
g16736 nor n16101 n16104 ; n16800
g16737 and n16103 n16104_not ; n16801
g16738 nor n16800 n16801 ; n16802
g16739 nor n16799 n16802 ; n16803
g16740 nor n16799 n16803 ; n16804
g16741 nor n16802 n16803 ; n16805
g16742 nor n16804 n16805 ; n16806
g16743 and n3457 n12567 ; n16807
g16744 and n3542 n12574 ; n16808
g16745 and n3606 n12571 ; n16809
g16746 nor n16808 n16809 ; n16810
g16747 and n16807_not n16810 ; n16811
g16748 and n3368 n15989 ; n16812
g16749 and n16811 n16812_not ; n16813
g16750 and a[29] n16813_not ; n16814
g16751 nor n16813 n16814 ; n16815
g16752 and a[29] n16814_not ; n16816
g16753 nor n16815 n16816 ; n16817
g16754 nor n16081 n16090 ; n16818
g16755 nor n16089 n16090 ; n16819
g16756 nor n16818 n16819 ; n16820
g16757 nor n16817 n16820 ; n16821
g16758 nor n16817 n16821 ; n16822
g16759 nor n16820 n16821 ; n16823
g16760 nor n16822 n16823 ; n16824
g16761 nor n7479 n12581 ; n16825
g16762 and n3606 n12581_not ; n16826
g16763 and n3457 n12577 ; n16827
g16764 nor n16826 n16827 ; n16828
g16765 and n3368 n16085_not ; n16829
g16766 and n16828 n16829_not ; n16830
g16767 and a[29] n16830_not ; n16831
g16768 and a[29] n16831_not ; n16832
g16769 nor n16830 n16831 ; n16833
g16770 nor n16832 n16833 ; n16834
g16771 nor n3367 n12581 ; n16835
g16772 and a[29] n16835_not ; n16836
g16773 and n16834_not n16836 ; n16837
g16774 and n3457 n12574 ; n16838
g16775 and n3542 n12581_not ; n16839
g16776 and n3606 n12577 ; n16840
g16777 nor n16839 n16840 ; n16841
g16778 and n16838_not n16841 ; n16842
g16779 and n3368_not n16842 ; n16843
g16780 and n16094 n16842 ; n16844
g16781 nor n16843 n16844 ; n16845
g16782 and a[29] n16845_not ; n16846
g16783 and a[29]_not n16845 ; n16847
g16784 nor n16846 n16847 ; n16848
g16785 and n16837 n16848_not ; n16849
g16786 and n16825 n16849 ; n16850
g16787 and n3457 n12571 ; n16851
g16788 and n3542 n12577 ; n16852
g16789 and n3606 n12574 ; n16853
g16790 nor n16852 n16853 ; n16854
g16791 and n16851_not n16854 ; n16855
g16792 and n3368 n16013 ; n16856
g16793 and n16855 n16856_not ; n16857
g16794 and a[29] n16857_not ; n16858
g16795 nor n16857 n16858 ; n16859
g16796 and a[29] n16858_not ; n16860
g16797 nor n16859 n16860 ; n16861
g16798 and n16825_not n16849 ; n16862
g16799 and n16825 n16849_not ; n16863
g16800 nor n16862 n16863 ; n16864
g16801 nor n16861 n16864 ; n16865
g16802 nor n16850 n16865 ; n16866
g16803 nor n16824 n16866 ; n16867
g16804 nor n16821 n16867 ; n16868
g16805 nor n16806 n16868 ; n16869
g16806 nor n16803 n16869 ; n16870
g16807 nor n16788 n16870 ; n16871
g16808 nor n16785 n16871 ; n16872
g16809 nor n16770 n16872 ; n16873
g16810 nor n16767 n16873 ; n16874
g16811 nor n16752 n16874 ; n16875
g16812 nor n16749 n16875 ; n16876
g16813 and n16722 n16733 ; n16877
g16814 nor n16734 n16877 ; n16878
g16815 and n16876_not n16878 ; n16879
g16816 nor n16734 n16879 ; n16880
g16817 and n16707 n16718 ; n16881
g16818 nor n16719 n16881 ; n16882
g16819 and n16880_not n16882 ; n16883
g16820 nor n16719 n16883 ; n16884
g16821 and n16692 n16703 ; n16885
g16822 nor n16704 n16885 ; n16886
g16823 and n16884_not n16886 ; n16887
g16824 nor n16704 n16887 ; n16888
g16825 and n16677 n16688 ; n16889
g16826 nor n16689 n16889 ; n16890
g16827 and n16888_not n16890 ; n16891
g16828 nor n16689 n16891 ; n16892
g16829 and n16662 n16673 ; n16893
g16830 nor n16674 n16893 ; n16894
g16831 and n16892_not n16894 ; n16895
g16832 nor n16674 n16895 ; n16896
g16833 and n16148_not n16159 ; n16897
g16834 nor n16160 n16897 ; n16898
g16835 and n16896_not n16898 ; n16899
g16836 and n16896 n16898_not ; n16900
g16837 nor n16899 n16900 ; n16901
g16838 and n3884 n12528 ; n16902
g16839 and n3967 n12534 ; n16903
g16840 and n4046 n12531 ; n16904
g16841 nor n16903 n16904 ; n16905
g16842 and n16902_not n16905 ; n16906
g16843 and n4050 n15003_not ; n16907
g16844 and n16906 n16907_not ; n16908
g16845 and a[26] n16908_not ; n16909
g16846 and a[26] n16909_not ; n16910
g16847 nor n16908 n16909 ; n16911
g16848 nor n16910 n16911 ; n16912
g16849 and n16901 n16912_not ; n16913
g16850 nor n16899 n16913 ; n16914
g16851 nor n16659 n16914 ; n16915
g16852 and n16659 n16914 ; n16916
g16853 nor n16915 n16916 ; n16917
g16854 and n4694 n12516 ; n16918
g16855 and n4533 n12522 ; n16919
g16856 and n4604 n12519 ; n16920
g16857 nor n16919 n16920 ; n16921
g16858 and n16918_not n16921 ; n16922
g16859 and n4536 n14443_not ; n16923
g16860 and n16922 n16923_not ; n16924
g16861 and a[23] n16924_not ; n16925
g16862 and a[23] n16925_not ; n16926
g16863 nor n16924 n16925 ; n16927
g16864 nor n16926 n16927 ; n16928
g16865 and n16917 n16928_not ; n16929
g16866 nor n16915 n16929 ; n16930
g16867 nor n16656 n16930 ; n16931
g16868 and n16656 n16930 ; n16932
g16869 nor n16931 n16932 ; n16933
g16870 and n5496 n12505 ; n16934
g16871 and n4935 n12513 ; n16935
g16872 and n5407 n12508 ; n16936
g16873 nor n16935 n16936 ; n16937
g16874 and n16934_not n16937 ; n16938
g16875 and n4938 n14051_not ; n16939
g16876 and n16938 n16939_not ; n16940
g16877 and a[20] n16940_not ; n16941
g16878 and a[20] n16941_not ; n16942
g16879 nor n16940 n16941 ; n16943
g16880 nor n16942 n16943 ; n16944
g16881 and n16933 n16944_not ; n16945
g16882 nor n16931 n16945 ; n16946
g16883 nor n16653 n16946 ; n16947
g16884 nor n16650 n16947 ; n16948
g16885 nor n16636 n16948 ; n16949
g16886 and n16636 n16948 ; n16950
g16887 nor n16949 n16950 ; n16951
g16888 and n6233 n13491 ; n16952
g16889 and n5663 n12769 ; n16953
g16890 and n5939 n12889 ; n16954
g16891 nor n16953 n16954 ; n16955
g16892 and n16952_not n16955 ; n16956
g16893 and n5666 n13503_not ; n16957
g16894 and n16956 n16957_not ; n16958
g16895 and a[17] n16958_not ; n16959
g16896 and a[17] n16959_not ; n16960
g16897 nor n16958 n16959 ; n16961
g16898 nor n16960 n16961 ; n16962
g16899 and n16951 n16962_not ; n16963
g16900 nor n16949 n16963 ; n16964
g16901 nor n16633 n16964 ; n16965
g16902 and n16633 n16964 ; n16966
g16903 nor n16965 n16966 ; n16967
g16904 and n7101 n13597 ; n16968
g16905 and n6402 n13521 ; n16969
g16906 and n6951 n13515 ; n16970
g16907 nor n16969 n16970 ; n16971
g16908 and n16968_not n16971 ; n16972
g16909 and n6397 n13612_not ; n16973
g16910 and n16972 n16973_not ; n16974
g16911 and a[14] n16974_not ; n16975
g16912 and a[14] n16975_not ; n16976
g16913 nor n16974 n16975 ; n16977
g16914 nor n16976 n16977 ; n16978
g16915 and n16967 n16978_not ; n16979
g16916 nor n16965 n16979 ; n16980
g16917 nor n16630 n16980 ; n16981
g16918 nor n16627 n16981 ; n16982
g16919 nor n16613 n16982 ; n16983
g16920 and n16613 n16982 ; n16984
g16921 nor n16983 n16984 ; n16985
g16922 and n7983 n13438_not ; n16986
g16923 and n7291 n13627_not ; n16987
g16924 and n7632 n13941 ; n16988
g16925 nor n16987 n16988 ; n16989
g16926 and n16986_not n16989 ; n16990
g16927 and n7294 n14028 ; n16991
g16928 and n16990 n16991_not ; n16992
g16929 and a[11] n16992_not ; n16993
g16930 and a[11] n16993_not ; n16994
g16931 nor n16992 n16993 ; n16995
g16932 nor n16994 n16995 ; n16996
g16933 and n16985 n16996_not ; n16997
g16934 nor n16983 n16997 ; n16998
g16935 nor n16610 n16998 ; n16999
g16936 and n16610 n16998 ; n17000
g16937 nor n16999 n17000 ; n17001
g16938 and n16985 n16997_not ; n17002
g16939 nor n16996 n16997 ; n17003
g16940 nor n17002 n17003 ; n17004
g16941 and n16967 n16979_not ; n17005
g16942 nor n16978 n16979 ; n17006
g16943 nor n17005 n17006 ; n17007
g16944 and n16951 n16963_not ; n17008
g16945 nor n16962 n16963 ; n17009
g16946 nor n17008 n17009 ; n17010
g16947 and n16653 n16946 ; n17011
g16948 nor n16947 n17011 ; n17012
g16949 and n6233 n12889 ; n17013
g16950 and n5663 n12502 ; n17014
g16951 and n5939 n12769 ; n17015
g16952 nor n17014 n17015 ; n17016
g16953 and n17013_not n17016 ; n17017
g16954 and n5666 n12895 ; n17018
g16955 and n17017 n17018_not ; n17019
g16956 and a[17] n17019_not ; n17020
g16957 and a[17] n17020_not ; n17021
g16958 nor n17019 n17020 ; n17022
g16959 nor n17021 n17022 ; n17023
g16960 and n17012 n17023_not ; n17024
g16961 and n17012 n17024_not ; n17025
g16962 nor n17023 n17024 ; n17026
g16963 nor n17025 n17026 ; n17027
g16964 and n16933 n16945_not ; n17028
g16965 nor n16944 n16945 ; n17029
g16966 nor n17028 n17029 ; n17030
g16967 and n16917 n16929_not ; n17031
g16968 nor n16928 n16929 ; n17032
g16969 nor n17031 n17032 ; n17033
g16970 and n16901 n16913_not ; n17034
g16971 nor n16912 n16913 ; n17035
g16972 nor n17034 n17035 ; n17036
g16973 and n16892 n16894_not ; n17037
g16974 nor n16895 n17037 ; n17038
g16975 and n3884 n12531 ; n17039
g16976 and n3967 n12537 ; n17040
g16977 and n4046 n12534 ; n17041
g16978 nor n17040 n17041 ; n17042
g16979 and n17039_not n17042 ; n17043
g16980 and n4050_not n17043 ; n17044
g16981 and n15255_not n17043 ; n17045
g16982 nor n17044 n17045 ; n17046
g16983 and a[26] n17046_not ; n17047
g16984 and a[26]_not n17046 ; n17048
g16985 nor n17047 n17048 ; n17049
g16986 and n17038 n17049_not ; n17050
g16987 and n16888 n16890_not ; n17051
g16988 nor n16891 n17051 ; n17052
g16989 and n3884 n12534 ; n17053
g16990 and n3967 n12540 ; n17054
g16991 and n4046 n12537 ; n17055
g16992 nor n17054 n17055 ; n17056
g16993 and n17053_not n17056 ; n17057
g16994 and n4050_not n17057 ; n17058
g16995 and n15096 n17057 ; n17059
g16996 nor n17058 n17059 ; n17060
g16997 and a[26] n17060_not ; n17061
g16998 and a[26]_not n17060 ; n17062
g16999 nor n17061 n17062 ; n17063
g17000 and n17052 n17063_not ; n17064
g17001 and n16884 n16886_not ; n17065
g17002 nor n16887 n17065 ; n17066
g17003 and n3884 n12537 ; n17067
g17004 and n3967 n12543 ; n17068
g17005 and n4046 n12540 ; n17069
g17006 nor n17068 n17069 ; n17070
g17007 and n17067_not n17070 ; n17071
g17008 and n4050_not n17071 ; n17072
g17009 and n15385 n17071 ; n17073
g17010 nor n17072 n17073 ; n17074
g17011 and a[26] n17074_not ; n17075
g17012 and a[26]_not n17074 ; n17076
g17013 nor n17075 n17076 ; n17077
g17014 and n17066 n17077_not ; n17078
g17015 and n16880 n16882_not ; n17079
g17016 nor n16883 n17079 ; n17080
g17017 and n3884 n12540 ; n17081
g17018 and n3967 n12546 ; n17082
g17019 and n4046 n12543 ; n17083
g17020 nor n17082 n17083 ; n17084
g17021 and n17081_not n17084 ; n17085
g17022 and n4050_not n17085 ; n17086
g17023 and n15708 n17085 ; n17087
g17024 nor n17086 n17087 ; n17088
g17025 and a[26] n17088_not ; n17089
g17026 and a[26]_not n17088 ; n17090
g17027 nor n17089 n17090 ; n17091
g17028 and n17080 n17091_not ; n17092
g17029 and n16876 n16878_not ; n17093
g17030 nor n16879 n17093 ; n17094
g17031 and n3884 n12543 ; n17095
g17032 and n3967 n12549 ; n17096
g17033 and n4046 n12546 ; n17097
g17034 nor n17096 n17097 ; n17098
g17035 and n17095_not n17098 ; n17099
g17036 and n4050_not n17099 ; n17100
g17037 and n15724_not n17099 ; n17101
g17038 nor n17100 n17101 ; n17102
g17039 and a[26] n17102_not ; n17103
g17040 and a[26]_not n17102 ; n17104
g17041 nor n17103 n17104 ; n17105
g17042 and n17094 n17105_not ; n17106
g17043 and n16752 n16874 ; n17107
g17044 nor n16875 n17107 ; n17108
g17045 and n3884 n12546 ; n17109
g17046 and n3967 n12552 ; n17110
g17047 and n4046 n12549 ; n17111
g17048 nor n17110 n17111 ; n17112
g17049 and n17109_not n17112 ; n17113
g17050 and n4050_not n17113 ; n17114
g17051 and n15356 n17113 ; n17115
g17052 nor n17114 n17115 ; n17116
g17053 and a[26] n17116_not ; n17117
g17054 and a[26]_not n17116 ; n17118
g17055 nor n17117 n17118 ; n17119
g17056 and n17108 n17119_not ; n17120
g17057 and n16770 n16872 ; n17121
g17058 nor n16873 n17121 ; n17122
g17059 and n3967 n12555 ; n17123
g17060 and n4046 n12552 ; n17124
g17061 and n3884 n12549 ; n17125
g17062 nor n17124 n17125 ; n17126
g17063 and n17123_not n17126 ; n17127
g17064 and n4050_not n17127 ; n17128
g17065 and n15764_not n17127 ; n17129
g17066 nor n17128 n17129 ; n17130
g17067 and a[26] n17130_not ; n17131
g17068 and a[26]_not n17130 ; n17132
g17069 nor n17131 n17132 ; n17133
g17070 and n17122 n17133_not ; n17134
g17071 and n16788 n16870 ; n17135
g17072 nor n16871 n17135 ; n17136
g17073 and n3967 n12558 ; n17137
g17074 and n3884 n12552 ; n17138
g17075 and n4046 n12555 ; n17139
g17076 nor n17138 n17139 ; n17140
g17077 and n17137_not n17140 ; n17141
g17078 and n4050_not n17141 ; n17142
g17079 and n15791 n17141 ; n17143
g17080 nor n17142 n17143 ; n17144
g17081 and a[26] n17144_not ; n17145
g17082 and a[26]_not n17144 ; n17146
g17083 nor n17145 n17146 ; n17147
g17084 and n17136 n17147_not ; n17148
g17085 and n16806 n16868 ; n17149
g17086 nor n16869 n17149 ; n17150
g17087 and n4046 n12558 ; n17151
g17088 and n3884 n12555 ; n17152
g17089 and n3967 n12561 ; n17153
g17090 nor n17152 n17153 ; n17154
g17091 and n17151_not n17154 ; n17155
g17092 and n4050_not n17155 ; n17156
g17093 and n15816 n17155 ; n17157
g17094 nor n17156 n17157 ; n17158
g17095 and a[26] n17158_not ; n17159
g17096 and a[26]_not n17158 ; n17160
g17097 nor n17159 n17160 ; n17161
g17098 and n17150 n17161_not ; n17162
g17099 nor n16824 n16867 ; n17163
g17100 nor n16866 n16867 ; n17164
g17101 nor n17163 n17164 ; n17165
g17102 and n3967 n12564 ; n17166
g17103 and n4046 n12561 ; n17167
g17104 and n3884 n12558 ; n17168
g17105 nor n17167 n17168 ; n17169
g17106 and n17166_not n17169 ; n17170
g17107 and n4050_not n17170 ; n17171
g17108 and n15847_not n17170 ; n17172
g17109 nor n17171 n17172 ; n17173
g17110 and a[26] n17173_not ; n17174
g17111 and a[26]_not n17173 ; n17175
g17112 nor n17174 n17175 ; n17176
g17113 nor n17165 n17176 ; n17177
g17114 and n4046 n12564 ; n17178
g17115 and n3884 n12561 ; n17179
g17116 and n3967 n12567 ; n17180
g17117 nor n17179 n17180 ; n17181
g17118 and n17178_not n17181 ; n17182
g17119 and n4050 n15905_not ; n17183
g17120 and n17182 n17183_not ; n17184
g17121 and a[26] n17184_not ; n17185
g17122 nor n17184 n17185 ; n17186
g17123 and a[26] n17185_not ; n17187
g17124 nor n17186 n17187 ; n17188
g17125 and n16861 n16864 ; n17189
g17126 nor n16865 n17189 ; n17190
g17127 and n17188_not n17190 ; n17191
g17128 nor n17188 n17191 ; n17192
g17129 and n17190 n17191_not ; n17193
g17130 nor n17192 n17193 ; n17194
g17131 and n3967 n12571 ; n17195
g17132 and n4046 n12567 ; n17196
g17133 and n3884 n12564 ; n17197
g17134 nor n17196 n17197 ; n17198
g17135 and n17195_not n17198 ; n17199
g17136 and n4050 n15944_not ; n17200
g17137 and n17199 n17200_not ; n17201
g17138 and a[26] n17201_not ; n17202
g17139 nor n17201 n17202 ; n17203
g17140 and a[26] n17202_not ; n17204
g17141 nor n17203 n17204 ; n17205
g17142 and n16837_not n16848 ; n17206
g17143 nor n16849 n17206 ; n17207
g17144 and n17205_not n17207 ; n17208
g17145 nor n17205 n17208 ; n17209
g17146 and n17207 n17208_not ; n17210
g17147 nor n17209 n17210 ; n17211
g17148 and n16834 n16836_not ; n17212
g17149 nor n16837 n17212 ; n17213
g17150 and n3967 n12574 ; n17214
g17151 and n3884 n12567 ; n17215
g17152 and n4046 n12571 ; n17216
g17153 nor n17215 n17216 ; n17217
g17154 and n17214_not n17217 ; n17218
g17155 and n4050_not n17218 ; n17219
g17156 and n15989_not n17218 ; n17220
g17157 nor n17219 n17220 ; n17221
g17158 and a[26] n17221_not ; n17222
g17159 and a[26]_not n17221 ; n17223
g17160 nor n17222 n17223 ; n17224
g17161 and n17213 n17224_not ; n17225
g17162 and n3884 n12577 ; n17226
g17163 and n4046 n12581_not ; n17227
g17164 nor n17226 n17227 ; n17228
g17165 and n4050 n16085_not ; n17229
g17166 and n17228 n17229_not ; n17230
g17167 and a[26] n17230_not ; n17231
g17168 and a[26] n17231_not ; n17232
g17169 nor n17230 n17231 ; n17233
g17170 nor n17232 n17233 ; n17234
g17171 nor n3880 n12581 ; n17235
g17172 and a[26] n17235_not ; n17236
g17173 and n17234_not n17236 ; n17237
g17174 and n3967 n12581_not ; n17238
g17175 and n3884 n12574 ; n17239
g17176 and n4046 n12577 ; n17240
g17177 nor n17239 n17240 ; n17241
g17178 and n17238_not n17241 ; n17242
g17179 and n4050_not n17242 ; n17243
g17180 and n16094 n17242 ; n17244
g17181 nor n17243 n17244 ; n17245
g17182 and a[26] n17245_not ; n17246
g17183 and a[26]_not n17245 ; n17247
g17184 nor n17246 n17247 ; n17248
g17185 and n17237 n17248_not ; n17249
g17186 and n16835 n17249 ; n17250
g17187 and n17249 n17250_not ; n17251
g17188 and n16835 n17250_not ; n17252
g17189 nor n17251 n17252 ; n17253
g17190 and n3967 n12577 ; n17254
g17191 and n3884 n12571 ; n17255
g17192 and n4046 n12574 ; n17256
g17193 nor n17255 n17256 ; n17257
g17194 and n17254_not n17257 ; n17258
g17195 and n4050 n16013 ; n17259
g17196 and n17258 n17259_not ; n17260
g17197 and a[26] n17260_not ; n17261
g17198 and a[26] n17261_not ; n17262
g17199 nor n17260 n17261 ; n17263
g17200 nor n17262 n17263 ; n17264
g17201 nor n17253 n17264 ; n17265
g17202 nor n17250 n17265 ; n17266
g17203 and n17213_not n17224 ; n17267
g17204 nor n17225 n17267 ; n17268
g17205 and n17266_not n17268 ; n17269
g17206 nor n17225 n17269 ; n17270
g17207 nor n17211 n17270 ; n17271
g17208 nor n17208 n17271 ; n17272
g17209 nor n17194 n17272 ; n17273
g17210 nor n17191 n17273 ; n17274
g17211 nor n17165 n17177 ; n17275
g17212 nor n17176 n17177 ; n17276
g17213 nor n17275 n17276 ; n17277
g17214 nor n17274 n17277 ; n17278
g17215 nor n17177 n17278 ; n17279
g17216 and n17150 n17162_not ; n17280
g17217 nor n17161 n17162 ; n17281
g17218 nor n17280 n17281 ; n17282
g17219 nor n17279 n17282 ; n17283
g17220 nor n17162 n17283 ; n17284
g17221 and n17136 n17148_not ; n17285
g17222 nor n17147 n17148 ; n17286
g17223 nor n17285 n17286 ; n17287
g17224 nor n17284 n17287 ; n17288
g17225 nor n17148 n17288 ; n17289
g17226 and n17122 n17134_not ; n17290
g17227 nor n17133 n17134 ; n17291
g17228 nor n17290 n17291 ; n17292
g17229 nor n17289 n17292 ; n17293
g17230 nor n17134 n17293 ; n17294
g17231 and n17108 n17120_not ; n17295
g17232 nor n17119 n17120 ; n17296
g17233 nor n17295 n17296 ; n17297
g17234 nor n17294 n17297 ; n17298
g17235 nor n17120 n17298 ; n17299
g17236 and n17094 n17106_not ; n17300
g17237 nor n17105 n17106 ; n17301
g17238 nor n17300 n17301 ; n17302
g17239 nor n17299 n17302 ; n17303
g17240 nor n17106 n17303 ; n17304
g17241 and n17080 n17092_not ; n17305
g17242 nor n17091 n17092 ; n17306
g17243 nor n17305 n17306 ; n17307
g17244 nor n17304 n17307 ; n17308
g17245 nor n17092 n17308 ; n17309
g17246 and n17066 n17078_not ; n17310
g17247 nor n17077 n17078 ; n17311
g17248 nor n17310 n17311 ; n17312
g17249 nor n17309 n17312 ; n17313
g17250 nor n17078 n17313 ; n17314
g17251 and n17052 n17064_not ; n17315
g17252 nor n17063 n17064 ; n17316
g17253 nor n17315 n17316 ; n17317
g17254 nor n17314 n17317 ; n17318
g17255 nor n17064 n17318 ; n17319
g17256 and n17038_not n17049 ; n17320
g17257 nor n17050 n17320 ; n17321
g17258 and n17319_not n17321 ; n17322
g17259 nor n17050 n17322 ; n17323
g17260 nor n17036 n17323 ; n17324
g17261 and n17036 n17323 ; n17325
g17262 nor n17324 n17325 ; n17326
g17263 and n4694 n12519 ; n17327
g17264 and n4533 n12525 ; n17328
g17265 and n4604 n12522 ; n17329
g17266 nor n17328 n17329 ; n17330
g17267 and n17327_not n17330 ; n17331
g17268 and n4536 n14454 ; n17332
g17269 and n17331 n17332_not ; n17333
g17270 and a[23] n17333_not ; n17334
g17271 and a[23] n17334_not ; n17335
g17272 nor n17333 n17334 ; n17336
g17273 nor n17335 n17336 ; n17337
g17274 and n17326 n17337_not ; n17338
g17275 nor n17324 n17338 ; n17339
g17276 nor n17033 n17339 ; n17340
g17277 and n17033 n17339 ; n17341
g17278 nor n17340 n17341 ; n17342
g17279 and n5496 n12508 ; n17343
g17280 and n4935 n12511 ; n17344
g17281 and n5407 n12513 ; n17345
g17282 nor n17344 n17345 ; n17346
g17283 and n17343_not n17346 ; n17347
g17284 and n4938 n13863 ; n17348
g17285 and n17347 n17348_not ; n17349
g17286 and a[20] n17349_not ; n17350
g17287 and a[20] n17350_not ; n17351
g17288 nor n17349 n17350 ; n17352
g17289 nor n17351 n17352 ; n17353
g17290 and n17342 n17353_not ; n17354
g17291 nor n17340 n17354 ; n17355
g17292 nor n17030 n17355 ; n17356
g17293 and n17030 n17355 ; n17357
g17294 nor n17356 n17357 ; n17358
g17295 and n6233 n12769 ; n17359
g17296 and n5663 n12370 ; n17360
g17297 and n5939 n12502 ; n17361
g17298 nor n17360 n17361 ; n17362
g17299 and n17359_not n17362 ; n17363
g17300 and n5666 n12999 ; n17364
g17301 and n17363 n17364_not ; n17365
g17302 and a[17] n17365_not ; n17366
g17303 and a[17] n17366_not ; n17367
g17304 nor n17365 n17366 ; n17368
g17305 nor n17367 n17368 ; n17369
g17306 and n17358 n17369_not ; n17370
g17307 nor n17356 n17370 ; n17371
g17308 nor n17027 n17371 ; n17372
g17309 nor n17024 n17372 ; n17373
g17310 nor n17010 n17373 ; n17374
g17311 and n17010 n17373 ; n17375
g17312 nor n17374 n17375 ; n17376
g17313 and n7101 n13515 ; n17377
g17314 and n6402 n13518 ; n17378
g17315 and n6951 n13521 ; n17379
g17316 nor n17378 n17379 ; n17380
g17317 and n17377_not n17380 ; n17381
g17318 and n6397 n13541 ; n17382
g17319 and n17381 n17382_not ; n17383
g17320 and a[14] n17383_not ; n17384
g17321 and a[14] n17384_not ; n17385
g17322 nor n17383 n17384 ; n17386
g17323 nor n17385 n17386 ; n17387
g17324 and n17376 n17387_not ; n17388
g17325 nor n17374 n17388 ; n17389
g17326 nor n17007 n17389 ; n17390
g17327 and n17007 n17389 ; n17391
g17328 nor n17390 n17391 ; n17392
g17329 and n7983 n13627_not ; n17393
g17330 and n7291 n13630 ; n17394
g17331 and n7632 n13633 ; n17395
g17332 nor n17394 n17395 ; n17396
g17333 and n17393_not n17396 ; n17397
g17334 and n7294 n13654_not ; n17398
g17335 and n17397 n17398_not ; n17399
g17336 and a[11] n17399_not ; n17400
g17337 and a[11] n17400_not ; n17401
g17338 nor n17399 n17400 ; n17402
g17339 nor n17401 n17402 ; n17403
g17340 and n17392 n17403_not ; n17404
g17341 nor n17390 n17404 ; n17405
g17342 and n7983 n13941 ; n17406
g17343 and n7291 n13633 ; n17407
g17344 and n7632 n13627_not ; n17408
g17345 nor n17407 n17408 ; n17409
g17346 and n17406_not n17409 ; n17410
g17347 and n7294 n14136 ; n17411
g17348 and n17410 n17411_not ; n17412
g17349 and a[11] n17412_not ; n17413
g17350 and a[11] n17413_not ; n17414
g17351 nor n17412 n17413 ; n17415
g17352 nor n17414 n17415 ; n17416
g17353 nor n17405 n17416 ; n17417
g17354 and n16630 n16980 ; n17418
g17355 nor n16981 n17418 ; n17419
g17356 nor n17405 n17417 ; n17420
g17357 nor n17416 n17417 ; n17421
g17358 nor n17420 n17421 ; n17422
g17359 and n17419 n17422_not ; n17423
g17360 nor n17417 n17423 ; n17424
g17361 nor n17004 n17424 ; n17425
g17362 nor n17004 n17425 ; n17426
g17363 nor n17424 n17425 ; n17427
g17364 nor n17426 n17427 ; n17428
g17365 and n17376 n17388_not ; n17429
g17366 nor n17387 n17388 ; n17430
g17367 nor n17429 n17430 ; n17431
g17368 and n17027 n17371 ; n17432
g17369 nor n17372 n17432 ; n17433
g17370 and n7101 n13521 ; n17434
g17371 and n6402 n13491 ; n17435
g17372 and n6951 n13518 ; n17436
g17373 nor n17435 n17436 ; n17437
g17374 and n17434_not n17437 ; n17438
g17375 and n6397 n13909_not ; n17439
g17376 and n17438 n17439_not ; n17440
g17377 and a[14] n17440_not ; n17441
g17378 and a[14] n17441_not ; n17442
g17379 nor n17440 n17441 ; n17443
g17380 nor n17442 n17443 ; n17444
g17381 and n17433 n17444_not ; n17445
g17382 and n17433 n17445_not ; n17446
g17383 nor n17444 n17445 ; n17447
g17384 nor n17446 n17447 ; n17448
g17385 and n17358 n17370_not ; n17449
g17386 nor n17369 n17370 ; n17450
g17387 nor n17449 n17450 ; n17451
g17388 and n17342 n17354_not ; n17452
g17389 nor n17353 n17354 ; n17453
g17390 nor n17452 n17453 ; n17454
g17391 and n17326 n17338_not ; n17455
g17392 nor n17337 n17338 ; n17456
g17393 nor n17455 n17456 ; n17457
g17394 and n4694 n12522 ; n17458
g17395 and n4533 n12528 ; n17459
g17396 and n4604 n12525 ; n17460
g17397 nor n17459 n17460 ; n17461
g17398 and n17458_not n17461 ; n17462
g17399 and n4536 n14837 ; n17463
g17400 and n17462 n17463_not ; n17464
g17401 and a[23] n17464_not ; n17465
g17402 nor n17464 n17465 ; n17466
g17403 and a[23] n17465_not ; n17467
g17404 nor n17466 n17467 ; n17468
g17405 and n17319 n17321_not ; n17469
g17406 nor n17322 n17469 ; n17470
g17407 and n17468_not n17470 ; n17471
g17408 nor n17468 n17471 ; n17472
g17409 and n17470 n17471_not ; n17473
g17410 nor n17472 n17473 ; n17474
g17411 and n4694 n12525 ; n17475
g17412 and n4533 n12531 ; n17476
g17413 and n4604 n12528 ; n17477
g17414 nor n17476 n17477 ; n17478
g17415 and n17475_not n17478 ; n17479
g17416 and n4536 n14608 ; n17480
g17417 and n17479 n17480_not ; n17481
g17418 and a[23] n17481_not ; n17482
g17419 nor n17481 n17482 ; n17483
g17420 and a[23] n17482_not ; n17484
g17421 nor n17483 n17484 ; n17485
g17422 nor n17314 n17318 ; n17486
g17423 nor n17317 n17318 ; n17487
g17424 nor n17486 n17487 ; n17488
g17425 nor n17485 n17488 ; n17489
g17426 nor n17485 n17489 ; n17490
g17427 nor n17488 n17489 ; n17491
g17428 nor n17490 n17491 ; n17492
g17429 and n4694 n12528 ; n17493
g17430 and n4533 n12534 ; n17494
g17431 and n4604 n12531 ; n17495
g17432 nor n17494 n17495 ; n17496
g17433 and n17493_not n17496 ; n17497
g17434 and n4536 n15003_not ; n17498
g17435 and n17497 n17498_not ; n17499
g17436 and a[23] n17499_not ; n17500
g17437 nor n17499 n17500 ; n17501
g17438 and a[23] n17500_not ; n17502
g17439 nor n17501 n17502 ; n17503
g17440 nor n17309 n17313 ; n17504
g17441 nor n17312 n17313 ; n17505
g17442 nor n17504 n17505 ; n17506
g17443 nor n17503 n17506 ; n17507
g17444 nor n17503 n17507 ; n17508
g17445 nor n17506 n17507 ; n17509
g17446 nor n17508 n17509 ; n17510
g17447 and n4694 n12531 ; n17511
g17448 and n4533 n12537 ; n17512
g17449 and n4604 n12534 ; n17513
g17450 nor n17512 n17513 ; n17514
g17451 and n17511_not n17514 ; n17515
g17452 and n4536 n15255 ; n17516
g17453 and n17515 n17516_not ; n17517
g17454 and a[23] n17517_not ; n17518
g17455 nor n17517 n17518 ; n17519
g17456 and a[23] n17518_not ; n17520
g17457 nor n17519 n17520 ; n17521
g17458 nor n17304 n17308 ; n17522
g17459 nor n17307 n17308 ; n17523
g17460 nor n17522 n17523 ; n17524
g17461 nor n17521 n17524 ; n17525
g17462 nor n17521 n17525 ; n17526
g17463 nor n17524 n17525 ; n17527
g17464 nor n17526 n17527 ; n17528
g17465 and n4694 n12534 ; n17529
g17466 and n4533 n12540 ; n17530
g17467 and n4604 n12537 ; n17531
g17468 nor n17530 n17531 ; n17532
g17469 and n17529_not n17532 ; n17533
g17470 and n4536 n15096_not ; n17534
g17471 and n17533 n17534_not ; n17535
g17472 and a[23] n17535_not ; n17536
g17473 nor n17535 n17536 ; n17537
g17474 and a[23] n17536_not ; n17538
g17475 nor n17537 n17538 ; n17539
g17476 nor n17299 n17303 ; n17540
g17477 nor n17302 n17303 ; n17541
g17478 nor n17540 n17541 ; n17542
g17479 nor n17539 n17542 ; n17543
g17480 nor n17539 n17543 ; n17544
g17481 nor n17542 n17543 ; n17545
g17482 nor n17544 n17545 ; n17546
g17483 and n4694 n12537 ; n17547
g17484 and n4533 n12543 ; n17548
g17485 and n4604 n12540 ; n17549
g17486 nor n17548 n17549 ; n17550
g17487 and n17547_not n17550 ; n17551
g17488 and n4536 n15385_not ; n17552
g17489 and n17551 n17552_not ; n17553
g17490 and a[23] n17553_not ; n17554
g17491 nor n17553 n17554 ; n17555
g17492 and a[23] n17554_not ; n17556
g17493 nor n17555 n17556 ; n17557
g17494 nor n17294 n17298 ; n17558
g17495 nor n17297 n17298 ; n17559
g17496 nor n17558 n17559 ; n17560
g17497 nor n17557 n17560 ; n17561
g17498 nor n17557 n17561 ; n17562
g17499 nor n17560 n17561 ; n17563
g17500 nor n17562 n17563 ; n17564
g17501 and n4694 n12540 ; n17565
g17502 and n4533 n12546 ; n17566
g17503 and n4604 n12543 ; n17567
g17504 nor n17566 n17567 ; n17568
g17505 and n17565_not n17568 ; n17569
g17506 and n4536 n15708_not ; n17570
g17507 and n17569 n17570_not ; n17571
g17508 and a[23] n17571_not ; n17572
g17509 nor n17571 n17572 ; n17573
g17510 and a[23] n17572_not ; n17574
g17511 nor n17573 n17574 ; n17575
g17512 nor n17289 n17293 ; n17576
g17513 nor n17292 n17293 ; n17577
g17514 nor n17576 n17577 ; n17578
g17515 nor n17575 n17578 ; n17579
g17516 nor n17575 n17579 ; n17580
g17517 nor n17578 n17579 ; n17581
g17518 nor n17580 n17581 ; n17582
g17519 and n4694 n12543 ; n17583
g17520 and n4533 n12549 ; n17584
g17521 and n4604 n12546 ; n17585
g17522 nor n17584 n17585 ; n17586
g17523 and n17583_not n17586 ; n17587
g17524 and n4536 n15724 ; n17588
g17525 and n17587 n17588_not ; n17589
g17526 and a[23] n17589_not ; n17590
g17527 nor n17589 n17590 ; n17591
g17528 and a[23] n17590_not ; n17592
g17529 nor n17591 n17592 ; n17593
g17530 nor n17284 n17288 ; n17594
g17531 nor n17287 n17288 ; n17595
g17532 nor n17594 n17595 ; n17596
g17533 nor n17593 n17596 ; n17597
g17534 nor n17593 n17597 ; n17598
g17535 nor n17596 n17597 ; n17599
g17536 nor n17598 n17599 ; n17600
g17537 and n4694 n12546 ; n17601
g17538 and n4533 n12552 ; n17602
g17539 and n4604 n12549 ; n17603
g17540 nor n17602 n17603 ; n17604
g17541 and n17601_not n17604 ; n17605
g17542 and n4536 n15356_not ; n17606
g17543 and n17605 n17606_not ; n17607
g17544 and a[23] n17607_not ; n17608
g17545 nor n17607 n17608 ; n17609
g17546 and a[23] n17608_not ; n17610
g17547 nor n17609 n17610 ; n17611
g17548 nor n17279 n17283 ; n17612
g17549 nor n17282 n17283 ; n17613
g17550 nor n17612 n17613 ; n17614
g17551 nor n17611 n17614 ; n17615
g17552 nor n17611 n17615 ; n17616
g17553 nor n17614 n17615 ; n17617
g17554 nor n17616 n17617 ; n17618
g17555 and n4694 n12549 ; n17619
g17556 and n4533 n12555 ; n17620
g17557 and n4604 n12552 ; n17621
g17558 nor n17620 n17621 ; n17622
g17559 and n17619_not n17622 ; n17623
g17560 and n4536 n15764 ; n17624
g17561 and n17623 n17624_not ; n17625
g17562 and a[23] n17625_not ; n17626
g17563 nor n17625 n17626 ; n17627
g17564 and a[23] n17626_not ; n17628
g17565 nor n17627 n17628 ; n17629
g17566 nor n17274 n17278 ; n17630
g17567 nor n17277 n17278 ; n17631
g17568 nor n17630 n17631 ; n17632
g17569 nor n17629 n17632 ; n17633
g17570 nor n17629 n17633 ; n17634
g17571 nor n17632 n17633 ; n17635
g17572 nor n17634 n17635 ; n17636
g17573 and n17194 n17272 ; n17637
g17574 nor n17273 n17637 ; n17638
g17575 and n4694 n12552 ; n17639
g17576 and n4533 n12558 ; n17640
g17577 and n4604 n12555 ; n17641
g17578 nor n17640 n17641 ; n17642
g17579 and n17639_not n17642 ; n17643
g17580 and n4536_not n17643 ; n17644
g17581 and n15791 n17643 ; n17645
g17582 nor n17644 n17645 ; n17646
g17583 and a[23] n17646_not ; n17647
g17584 and a[23]_not n17646 ; n17648
g17585 nor n17647 n17648 ; n17649
g17586 and n17638 n17649_not ; n17650
g17587 and n17211 n17270 ; n17651
g17588 nor n17271 n17651 ; n17652
g17589 and n4694 n12555 ; n17653
g17590 and n4533 n12561 ; n17654
g17591 and n4604 n12558 ; n17655
g17592 nor n17654 n17655 ; n17656
g17593 and n17653_not n17656 ; n17657
g17594 and n4536_not n17657 ; n17658
g17595 and n15816 n17657 ; n17659
g17596 nor n17658 n17659 ; n17660
g17597 and a[23] n17660_not ; n17661
g17598 and a[23]_not n17660 ; n17662
g17599 nor n17661 n17662 ; n17663
g17600 and n17652 n17663_not ; n17664
g17601 and n4694 n12558 ; n17665
g17602 and n4533 n12564 ; n17666
g17603 and n4604 n12561 ; n17667
g17604 nor n17666 n17667 ; n17668
g17605 and n17665_not n17668 ; n17669
g17606 and n4536 n15847 ; n17670
g17607 and n17669 n17670_not ; n17671
g17608 and a[23] n17671_not ; n17672
g17609 nor n17671 n17672 ; n17673
g17610 and a[23] n17672_not ; n17674
g17611 nor n17673 n17674 ; n17675
g17612 and n17266 n17268_not ; n17676
g17613 nor n17269 n17676 ; n17677
g17614 and n17675_not n17677 ; n17678
g17615 nor n17675 n17678 ; n17679
g17616 and n17677 n17678_not ; n17680
g17617 nor n17679 n17680 ; n17681
g17618 nor n17253 n17265 ; n17682
g17619 nor n17264 n17265 ; n17683
g17620 nor n17682 n17683 ; n17684
g17621 and n4694 n12561 ; n17685
g17622 and n4533 n12567 ; n17686
g17623 and n4604 n12564 ; n17687
g17624 nor n17686 n17687 ; n17688
g17625 and n17685_not n17688 ; n17689
g17626 and n4536_not n17689 ; n17690
g17627 and n15905 n17689 ; n17691
g17628 nor n17690 n17691 ; n17692
g17629 and a[23] n17692_not ; n17693
g17630 and a[23]_not n17692 ; n17694
g17631 nor n17693 n17694 ; n17695
g17632 nor n17684 n17695 ; n17696
g17633 and n4694 n12564 ; n17697
g17634 and n4533 n12571 ; n17698
g17635 and n4604 n12567 ; n17699
g17636 nor n17698 n17699 ; n17700
g17637 and n17697_not n17700 ; n17701
g17638 and n4536 n15944_not ; n17702
g17639 and n17701 n17702_not ; n17703
g17640 and a[23] n17703_not ; n17704
g17641 nor n17703 n17704 ; n17705
g17642 and a[23] n17704_not ; n17706
g17643 nor n17705 n17706 ; n17707
g17644 and n17237_not n17248 ; n17708
g17645 nor n17249 n17708 ; n17709
g17646 and n17707_not n17709 ; n17710
g17647 nor n17707 n17710 ; n17711
g17648 and n17709 n17710_not ; n17712
g17649 nor n17711 n17712 ; n17713
g17650 and n17234 n17236_not ; n17714
g17651 nor n17237 n17714 ; n17715
g17652 and n4694 n12567 ; n17716
g17653 and n4533 n12574 ; n17717
g17654 and n4604 n12571 ; n17718
g17655 nor n17717 n17718 ; n17719
g17656 and n17716_not n17719 ; n17720
g17657 and n4536_not n17720 ; n17721
g17658 and n15989_not n17720 ; n17722
g17659 nor n17721 n17722 ; n17723
g17660 and a[23] n17723_not ; n17724
g17661 and a[23]_not n17723 ; n17725
g17662 nor n17724 n17725 ; n17726
g17663 and n17715 n17726_not ; n17727
g17664 and n4604 n12581_not ; n17728
g17665 and n4694 n12577 ; n17729
g17666 nor n17728 n17729 ; n17730
g17667 and n4536 n16085_not ; n17731
g17668 and n17730 n17731_not ; n17732
g17669 and a[23] n17732_not ; n17733
g17670 and a[23] n17733_not ; n17734
g17671 nor n17732 n17733 ; n17735
g17672 nor n17734 n17735 ; n17736
g17673 nor n4528 n12581 ; n17737
g17674 and a[23] n17737_not ; n17738
g17675 and n17736_not n17738 ; n17739
g17676 and n4694 n12574 ; n17740
g17677 and n4533 n12581_not ; n17741
g17678 and n4604 n12577 ; n17742
g17679 nor n17741 n17742 ; n17743
g17680 and n17740_not n17743 ; n17744
g17681 and n4536_not n17744 ; n17745
g17682 and n16094 n17744 ; n17746
g17683 nor n17745 n17746 ; n17747
g17684 and a[23] n17747_not ; n17748
g17685 and a[23]_not n17747 ; n17749
g17686 nor n17748 n17749 ; n17750
g17687 and n17739 n17750_not ; n17751
g17688 and n17235 n17751 ; n17752
g17689 and n17751 n17752_not ; n17753
g17690 and n17235 n17752_not ; n17754
g17691 nor n17753 n17754 ; n17755
g17692 and n4694 n12571 ; n17756
g17693 and n4533 n12577 ; n17757
g17694 and n4604 n12574 ; n17758
g17695 nor n17757 n17758 ; n17759
g17696 and n17756_not n17759 ; n17760
g17697 and n4536 n16013 ; n17761
g17698 and n17760 n17761_not ; n17762
g17699 and a[23] n17762_not ; n17763
g17700 and a[23] n17763_not ; n17764
g17701 nor n17762 n17763 ; n17765
g17702 nor n17764 n17765 ; n17766
g17703 nor n17755 n17766 ; n17767
g17704 nor n17752 n17767 ; n17768
g17705 and n17715_not n17726 ; n17769
g17706 nor n17727 n17769 ; n17770
g17707 and n17768_not n17770 ; n17771
g17708 nor n17727 n17771 ; n17772
g17709 nor n17713 n17772 ; n17773
g17710 nor n17710 n17773 ; n17774
g17711 and n17684 n17695 ; n17775
g17712 nor n17696 n17775 ; n17776
g17713 and n17774_not n17776 ; n17777
g17714 nor n17696 n17777 ; n17778
g17715 nor n17681 n17778 ; n17779
g17716 nor n17678 n17779 ; n17780
g17717 and n17652 n17664_not ; n17781
g17718 nor n17663 n17664 ; n17782
g17719 nor n17781 n17782 ; n17783
g17720 nor n17780 n17783 ; n17784
g17721 nor n17664 n17784 ; n17785
g17722 and n17638_not n17649 ; n17786
g17723 nor n17650 n17786 ; n17787
g17724 and n17785_not n17787 ; n17788
g17725 nor n17650 n17788 ; n17789
g17726 nor n17636 n17789 ; n17790
g17727 nor n17633 n17790 ; n17791
g17728 nor n17618 n17791 ; n17792
g17729 nor n17615 n17792 ; n17793
g17730 nor n17600 n17793 ; n17794
g17731 nor n17597 n17794 ; n17795
g17732 nor n17582 n17795 ; n17796
g17733 nor n17579 n17796 ; n17797
g17734 nor n17564 n17797 ; n17798
g17735 nor n17561 n17798 ; n17799
g17736 nor n17546 n17799 ; n17800
g17737 nor n17543 n17800 ; n17801
g17738 nor n17528 n17801 ; n17802
g17739 nor n17525 n17802 ; n17803
g17740 nor n17510 n17803 ; n17804
g17741 nor n17507 n17804 ; n17805
g17742 nor n17492 n17805 ; n17806
g17743 nor n17489 n17806 ; n17807
g17744 nor n17474 n17807 ; n17808
g17745 nor n17471 n17808 ; n17809
g17746 nor n17457 n17809 ; n17810
g17747 and n17457 n17809 ; n17811
g17748 nor n17810 n17811 ; n17812
g17749 and n5496 n12513 ; n17813
g17750 and n4935 n12516 ; n17814
g17751 and n5407 n12511 ; n17815
g17752 nor n17814 n17815 ; n17816
g17753 and n17813_not n17816 ; n17817
g17754 and n4938 n14177 ; n17818
g17755 and n17817 n17818_not ; n17819
g17756 and a[20] n17819_not ; n17820
g17757 and a[20] n17820_not ; n17821
g17758 nor n17819 n17820 ; n17822
g17759 nor n17821 n17822 ; n17823
g17760 and n17812 n17823_not ; n17824
g17761 nor n17810 n17824 ; n17825
g17762 nor n17454 n17825 ; n17826
g17763 and n17454 n17825 ; n17827
g17764 nor n17826 n17827 ; n17828
g17765 and n6233 n12502 ; n17829
g17766 and n5663 n12505 ; n17830
g17767 and n5939 n12370 ; n17831
g17768 nor n17830 n17831 ; n17832
g17769 and n17829_not n17832 ; n17833
g17770 and n5666 n13736_not ; n17834
g17771 and n17833 n17834_not ; n17835
g17772 and a[17] n17835_not ; n17836
g17773 and a[17] n17836_not ; n17837
g17774 nor n17835 n17836 ; n17838
g17775 nor n17837 n17838 ; n17839
g17776 and n17828 n17839_not ; n17840
g17777 nor n17826 n17840 ; n17841
g17778 nor n17451 n17841 ; n17842
g17779 and n17451 n17841 ; n17843
g17780 nor n17842 n17843 ; n17844
g17781 and n7101 n13518 ; n17845
g17782 and n6402 n12889 ; n17846
g17783 and n6951 n13491 ; n17847
g17784 nor n17846 n17847 ; n17848
g17785 and n17845_not n17848 ; n17849
g17786 and n6397 n13584 ; n17850
g17787 and n17849 n17850_not ; n17851
g17788 and a[14] n17851_not ; n17852
g17789 and a[14] n17852_not ; n17853
g17790 nor n17851 n17852 ; n17854
g17791 nor n17853 n17854 ; n17855
g17792 and n17844 n17855_not ; n17856
g17793 nor n17842 n17856 ; n17857
g17794 nor n17448 n17857 ; n17858
g17795 nor n17445 n17858 ; n17859
g17796 nor n17431 n17859 ; n17860
g17797 and n17431 n17859 ; n17861
g17798 nor n17860 n17861 ; n17862
g17799 and n7983 n13633 ; n17863
g17800 and n7291 n13597 ; n17864
g17801 and n7632 n13630 ; n17865
g17802 nor n17864 n17865 ; n17866
g17803 and n17863_not n17866 ; n17867
g17804 and n7294 n13929 ; n17868
g17805 and n17867 n17868_not ; n17869
g17806 and a[11] n17869_not ; n17870
g17807 and a[11] n17870_not ; n17871
g17808 nor n17869 n17870 ; n17872
g17809 nor n17871 n17872 ; n17873
g17810 and n17862 n17873_not ; n17874
g17811 nor n17860 n17874 ; n17875
g17812 nor n13438 n14590 ; n17876
g17813 and n8418 n13941 ; n17877
g17814 nor n17876 n17877 ; n17878
g17815 and n8421_not n17878 ; n17879
g17816 and n13951 n17878 ; n17880
g17817 nor n17879 n17880 ; n17881
g17818 and a[8] n17881_not ; n17882
g17819 and a[8]_not n17881 ; n17883
g17820 nor n17882 n17883 ; n17884
g17821 nor n17875 n17884 ; n17885
g17822 and n17392 n17404_not ; n17886
g17823 nor n17403 n17404 ; n17887
g17824 nor n17886 n17887 ; n17888
g17825 and n17875 n17884 ; n17889
g17826 nor n17885 n17889 ; n17890
g17827 and n17888_not n17890 ; n17891
g17828 nor n17885 n17891 ; n17892
g17829 and n17419_not n17422 ; n17893
g17830 nor n17423 n17893 ; n17894
g17831 and n17892_not n17894 ; n17895
g17832 nor n17888 n17891 ; n17896
g17833 and n17890 n17891_not ; n17897
g17834 nor n17896 n17897 ; n17898
g17835 and n17862 n17874_not ; n17899
g17836 nor n17873 n17874 ; n17900
g17837 nor n17899 n17900 ; n17901
g17838 and n17448 n17857 ; n17902
g17839 nor n17858 n17902 ; n17903
g17840 and n7983 n13630 ; n17904
g17841 and n7291 n13515 ; n17905
g17842 and n7632 n13597 ; n17906
g17843 nor n17905 n17906 ; n17907
g17844 and n17904_not n17907 ; n17908
g17845 and n7294 n13976 ; n17909
g17846 and n17908 n17909_not ; n17910
g17847 and a[11] n17910_not ; n17911
g17848 and a[11] n17911_not ; n17912
g17849 nor n17910 n17911 ; n17913
g17850 nor n17912 n17913 ; n17914
g17851 and n17903 n17914_not ; n17915
g17852 and n17903 n17915_not ; n17916
g17853 nor n17914 n17915 ; n17917
g17854 nor n17916 n17917 ; n17918
g17855 and n17844 n17856_not ; n17919
g17856 nor n17855 n17856 ; n17920
g17857 nor n17919 n17920 ; n17921
g17858 and n17828 n17840_not ; n17922
g17859 nor n17839 n17840 ; n17923
g17860 nor n17922 n17923 ; n17924
g17861 and n17812 n17824_not ; n17925
g17862 nor n17823 n17824 ; n17926
g17863 nor n17925 n17926 ; n17927
g17864 and n17474 n17807 ; n17928
g17865 nor n17808 n17928 ; n17929
g17866 and n5496 n12511 ; n17930
g17867 and n4935 n12519 ; n17931
g17868 and n5407 n12516 ; n17932
g17869 nor n17931 n17932 ; n17933
g17870 and n17930_not n17933 ; n17934
g17871 and n4938_not n17934 ; n17935
g17872 and n14233 n17934 ; n17936
g17873 nor n17935 n17936 ; n17937
g17874 and a[20] n17937_not ; n17938
g17875 and a[20]_not n17937 ; n17939
g17876 nor n17938 n17939 ; n17940
g17877 and n17929 n17940_not ; n17941
g17878 and n17492 n17805 ; n17942
g17879 nor n17806 n17942 ; n17943
g17880 and n5496 n12516 ; n17944
g17881 and n4935 n12522 ; n17945
g17882 and n5407 n12519 ; n17946
g17883 nor n17945 n17946 ; n17947
g17884 and n17944_not n17947 ; n17948
g17885 and n4938_not n17948 ; n17949
g17886 and n14443 n17948 ; n17950
g17887 nor n17949 n17950 ; n17951
g17888 and a[20] n17951_not ; n17952
g17889 and a[20]_not n17951 ; n17953
g17890 nor n17952 n17953 ; n17954
g17891 and n17943 n17954_not ; n17955
g17892 and n17510 n17803 ; n17956
g17893 nor n17804 n17956 ; n17957
g17894 and n5496 n12519 ; n17958
g17895 and n4935 n12525 ; n17959
g17896 and n5407 n12522 ; n17960
g17897 nor n17959 n17960 ; n17961
g17898 and n17958_not n17961 ; n17962
g17899 and n4938_not n17962 ; n17963
g17900 and n14454_not n17962 ; n17964
g17901 nor n17963 n17964 ; n17965
g17902 and a[20] n17965_not ; n17966
g17903 and a[20]_not n17965 ; n17967
g17904 nor n17966 n17967 ; n17968
g17905 and n17957 n17968_not ; n17969
g17906 and n17528 n17801 ; n17970
g17907 nor n17802 n17970 ; n17971
g17908 and n5496 n12522 ; n17972
g17909 and n4935 n12528 ; n17973
g17910 and n5407 n12525 ; n17974
g17911 nor n17973 n17974 ; n17975
g17912 and n17972_not n17975 ; n17976
g17913 and n4938_not n17976 ; n17977
g17914 and n14837_not n17976 ; n17978
g17915 nor n17977 n17978 ; n17979
g17916 and a[20] n17979_not ; n17980
g17917 and a[20]_not n17979 ; n17981
g17918 nor n17980 n17981 ; n17982
g17919 and n17971 n17982_not ; n17983
g17920 and n17546 n17799 ; n17984
g17921 nor n17800 n17984 ; n17985
g17922 and n5496 n12525 ; n17986
g17923 and n4935 n12531 ; n17987
g17924 and n5407 n12528 ; n17988
g17925 nor n17987 n17988 ; n17989
g17926 and n17986_not n17989 ; n17990
g17927 and n4938_not n17990 ; n17991
g17928 and n14608_not n17990 ; n17992
g17929 nor n17991 n17992 ; n17993
g17930 and a[20] n17993_not ; n17994
g17931 and a[20]_not n17993 ; n17995
g17932 nor n17994 n17995 ; n17996
g17933 and n17985 n17996_not ; n17997
g17934 and n17564 n17797 ; n17998
g17935 nor n17798 n17998 ; n17999
g17936 and n5496 n12528 ; n18000
g17937 and n4935 n12534 ; n18001
g17938 and n5407 n12531 ; n18002
g17939 nor n18001 n18002 ; n18003
g17940 and n18000_not n18003 ; n18004
g17941 and n4938_not n18004 ; n18005
g17942 and n15003 n18004 ; n18006
g17943 nor n18005 n18006 ; n18007
g17944 and a[20] n18007_not ; n18008
g17945 and a[20]_not n18007 ; n18009
g17946 nor n18008 n18009 ; n18010
g17947 and n17999 n18010_not ; n18011
g17948 and n17582 n17795 ; n18012
g17949 nor n17796 n18012 ; n18013
g17950 and n5496 n12531 ; n18014
g17951 and n4935 n12537 ; n18015
g17952 and n5407 n12534 ; n18016
g17953 nor n18015 n18016 ; n18017
g17954 and n18014_not n18017 ; n18018
g17955 and n4938_not n18018 ; n18019
g17956 and n15255_not n18018 ; n18020
g17957 nor n18019 n18020 ; n18021
g17958 and a[20] n18021_not ; n18022
g17959 and a[20]_not n18021 ; n18023
g17960 nor n18022 n18023 ; n18024
g17961 and n18013 n18024_not ; n18025
g17962 and n17600 n17793 ; n18026
g17963 nor n17794 n18026 ; n18027
g17964 and n5496 n12534 ; n18028
g17965 and n4935 n12540 ; n18029
g17966 and n5407 n12537 ; n18030
g17967 nor n18029 n18030 ; n18031
g17968 and n18028_not n18031 ; n18032
g17969 and n4938_not n18032 ; n18033
g17970 and n15096 n18032 ; n18034
g17971 nor n18033 n18034 ; n18035
g17972 and a[20] n18035_not ; n18036
g17973 and a[20]_not n18035 ; n18037
g17974 nor n18036 n18037 ; n18038
g17975 and n18027 n18038_not ; n18039
g17976 and n17618 n17791 ; n18040
g17977 nor n17792 n18040 ; n18041
g17978 and n5496 n12537 ; n18042
g17979 and n4935 n12543 ; n18043
g17980 and n5407 n12540 ; n18044
g17981 nor n18043 n18044 ; n18045
g17982 and n18042_not n18045 ; n18046
g17983 and n4938_not n18046 ; n18047
g17984 and n15385 n18046 ; n18048
g17985 nor n18047 n18048 ; n18049
g17986 and a[20] n18049_not ; n18050
g17987 and a[20]_not n18049 ; n18051
g17988 nor n18050 n18051 ; n18052
g17989 and n18041 n18052_not ; n18053
g17990 and n17636 n17789 ; n18054
g17991 nor n17790 n18054 ; n18055
g17992 and n5496 n12540 ; n18056
g17993 and n4935 n12546 ; n18057
g17994 and n5407 n12543 ; n18058
g17995 nor n18057 n18058 ; n18059
g17996 and n18056_not n18059 ; n18060
g17997 and n4938_not n18060 ; n18061
g17998 and n15708 n18060 ; n18062
g17999 nor n18061 n18062 ; n18063
g18000 and a[20] n18063_not ; n18064
g18001 and a[20]_not n18063 ; n18065
g18002 nor n18064 n18065 ; n18066
g18003 and n18055 n18066_not ; n18067
g18004 and n5496 n12543 ; n18068
g18005 and n4935 n12549 ; n18069
g18006 and n5407 n12546 ; n18070
g18007 nor n18069 n18070 ; n18071
g18008 and n18068_not n18071 ; n18072
g18009 and n4938 n15724 ; n18073
g18010 and n18072 n18073_not ; n18074
g18011 and a[20] n18074_not ; n18075
g18012 nor n18074 n18075 ; n18076
g18013 and a[20] n18075_not ; n18077
g18014 nor n18076 n18077 ; n18078
g18015 and n17785 n17787_not ; n18079
g18016 nor n17788 n18079 ; n18080
g18017 and n18078_not n18080 ; n18081
g18018 nor n18078 n18081 ; n18082
g18019 and n18080 n18081_not ; n18083
g18020 nor n18082 n18083 ; n18084
g18021 and n5496 n12546 ; n18085
g18022 and n4935 n12552 ; n18086
g18023 and n5407 n12549 ; n18087
g18024 nor n18086 n18087 ; n18088
g18025 and n18085_not n18088 ; n18089
g18026 and n4938 n15356_not ; n18090
g18027 and n18089 n18090_not ; n18091
g18028 and a[20] n18091_not ; n18092
g18029 nor n18091 n18092 ; n18093
g18030 and a[20] n18092_not ; n18094
g18031 nor n18093 n18094 ; n18095
g18032 nor n17780 n17784 ; n18096
g18033 nor n17783 n17784 ; n18097
g18034 nor n18096 n18097 ; n18098
g18035 nor n18095 n18098 ; n18099
g18036 nor n18095 n18099 ; n18100
g18037 nor n18098 n18099 ; n18101
g18038 nor n18100 n18101 ; n18102
g18039 and n17681 n17778 ; n18103
g18040 nor n17779 n18103 ; n18104
g18041 and n5496 n12549 ; n18105
g18042 and n4935 n12555 ; n18106
g18043 and n5407 n12552 ; n18107
g18044 nor n18106 n18107 ; n18108
g18045 and n18105_not n18108 ; n18109
g18046 and n4938_not n18109 ; n18110
g18047 and n15764_not n18109 ; n18111
g18048 nor n18110 n18111 ; n18112
g18049 and a[20] n18112_not ; n18113
g18050 and a[20]_not n18112 ; n18114
g18051 nor n18113 n18114 ; n18115
g18052 and n18104 n18115_not ; n18116
g18053 and n17774 n17776_not ; n18117
g18054 nor n17777 n18117 ; n18118
g18055 and n5496 n12552 ; n18119
g18056 and n4935 n12558 ; n18120
g18057 and n5407 n12555 ; n18121
g18058 nor n18120 n18121 ; n18122
g18059 and n18119_not n18122 ; n18123
g18060 and n4938_not n18123 ; n18124
g18061 and n15791 n18123 ; n18125
g18062 nor n18124 n18125 ; n18126
g18063 and a[20] n18126_not ; n18127
g18064 and a[20]_not n18126 ; n18128
g18065 nor n18127 n18128 ; n18129
g18066 and n18118 n18129_not ; n18130
g18067 and n17713 n17772 ; n18131
g18068 nor n17773 n18131 ; n18132
g18069 and n5496 n12555 ; n18133
g18070 and n4935 n12561 ; n18134
g18071 and n5407 n12558 ; n18135
g18072 nor n18134 n18135 ; n18136
g18073 and n18133_not n18136 ; n18137
g18074 and n4938_not n18137 ; n18138
g18075 and n15816 n18137 ; n18139
g18076 nor n18138 n18139 ; n18140
g18077 and a[20] n18140_not ; n18141
g18078 and a[20]_not n18140 ; n18142
g18079 nor n18141 n18142 ; n18143
g18080 and n18132 n18143_not ; n18144
g18081 and n5496 n12558 ; n18145
g18082 and n4935 n12564 ; n18146
g18083 and n5407 n12561 ; n18147
g18084 nor n18146 n18147 ; n18148
g18085 and n18145_not n18148 ; n18149
g18086 and n4938 n15847 ; n18150
g18087 and n18149 n18150_not ; n18151
g18088 and a[20] n18151_not ; n18152
g18089 nor n18151 n18152 ; n18153
g18090 and a[20] n18152_not ; n18154
g18091 nor n18153 n18154 ; n18155
g18092 and n17768 n17770_not ; n18156
g18093 nor n17771 n18156 ; n18157
g18094 and n18155_not n18157 ; n18158
g18095 nor n18155 n18158 ; n18159
g18096 and n18157 n18158_not ; n18160
g18097 nor n18159 n18160 ; n18161
g18098 nor n17755 n17767 ; n18162
g18099 nor n17766 n17767 ; n18163
g18100 nor n18162 n18163 ; n18164
g18101 and n5496 n12561 ; n18165
g18102 and n4935 n12567 ; n18166
g18103 and n5407 n12564 ; n18167
g18104 nor n18166 n18167 ; n18168
g18105 and n18165_not n18168 ; n18169
g18106 and n4938_not n18169 ; n18170
g18107 and n15905 n18169 ; n18171
g18108 nor n18170 n18171 ; n18172
g18109 and a[20] n18172_not ; n18173
g18110 and a[20]_not n18172 ; n18174
g18111 nor n18173 n18174 ; n18175
g18112 nor n18164 n18175 ; n18176
g18113 and n5496 n12564 ; n18177
g18114 and n4935 n12571 ; n18178
g18115 and n5407 n12567 ; n18179
g18116 nor n18178 n18179 ; n18180
g18117 and n18177_not n18180 ; n18181
g18118 and n4938 n15944_not ; n18182
g18119 and n18181 n18182_not ; n18183
g18120 and a[20] n18183_not ; n18184
g18121 nor n18183 n18184 ; n18185
g18122 and a[20] n18184_not ; n18186
g18123 nor n18185 n18186 ; n18187
g18124 and n17739_not n17750 ; n18188
g18125 nor n17751 n18188 ; n18189
g18126 and n18187_not n18189 ; n18190
g18127 nor n18187 n18190 ; n18191
g18128 and n18189 n18190_not ; n18192
g18129 nor n18191 n18192 ; n18193
g18130 and n17736 n17738_not ; n18194
g18131 nor n17739 n18194 ; n18195
g18132 and n5496 n12567 ; n18196
g18133 and n4935 n12574 ; n18197
g18134 and n5407 n12571 ; n18198
g18135 nor n18197 n18198 ; n18199
g18136 and n18196_not n18199 ; n18200
g18137 and n4938_not n18200 ; n18201
g18138 and n15989_not n18200 ; n18202
g18139 nor n18201 n18202 ; n18203
g18140 and a[20] n18203_not ; n18204
g18141 and a[20]_not n18203 ; n18205
g18142 nor n18204 n18205 ; n18206
g18143 and n18195 n18206_not ; n18207
g18144 and n5407 n12581_not ; n18208
g18145 and n5496 n12577 ; n18209
g18146 nor n18208 n18209 ; n18210
g18147 and n4938 n16085_not ; n18211
g18148 and n18210 n18211_not ; n18212
g18149 and a[20] n18212_not ; n18213
g18150 and a[20] n18213_not ; n18214
g18151 nor n18212 n18213 ; n18215
g18152 nor n18214 n18215 ; n18216
g18153 nor n4933 n12581 ; n18217
g18154 and a[20] n18217_not ; n18218
g18155 and n18216_not n18218 ; n18219
g18156 and n5496 n12574 ; n18220
g18157 and n4935 n12581_not ; n18221
g18158 and n5407 n12577 ; n18222
g18159 nor n18221 n18222 ; n18223
g18160 and n18220_not n18223 ; n18224
g18161 and n4938_not n18224 ; n18225
g18162 and n16094 n18224 ; n18226
g18163 nor n18225 n18226 ; n18227
g18164 and a[20] n18227_not ; n18228
g18165 and a[20]_not n18227 ; n18229
g18166 nor n18228 n18229 ; n18230
g18167 and n18219 n18230_not ; n18231
g18168 and n17737 n18231 ; n18232
g18169 and n18231 n18232_not ; n18233
g18170 and n17737 n18232_not ; n18234
g18171 nor n18233 n18234 ; n18235
g18172 and n5496 n12571 ; n18236
g18173 and n4935 n12577 ; n18237
g18174 and n5407 n12574 ; n18238
g18175 nor n18237 n18238 ; n18239
g18176 and n18236_not n18239 ; n18240
g18177 and n4938 n16013 ; n18241
g18178 and n18240 n18241_not ; n18242
g18179 and a[20] n18242_not ; n18243
g18180 and a[20] n18243_not ; n18244
g18181 nor n18242 n18243 ; n18245
g18182 nor n18244 n18245 ; n18246
g18183 nor n18235 n18246 ; n18247
g18184 nor n18232 n18247 ; n18248
g18185 and n18195_not n18206 ; n18249
g18186 nor n18207 n18249 ; n18250
g18187 and n18248_not n18250 ; n18251
g18188 nor n18207 n18251 ; n18252
g18189 nor n18193 n18252 ; n18253
g18190 nor n18190 n18253 ; n18254
g18191 and n18164 n18175 ; n18255
g18192 nor n18176 n18255 ; n18256
g18193 and n18254_not n18256 ; n18257
g18194 nor n18176 n18257 ; n18258
g18195 nor n18161 n18258 ; n18259
g18196 nor n18158 n18259 ; n18260
g18197 and n18132 n18144_not ; n18261
g18198 nor n18143 n18144 ; n18262
g18199 nor n18261 n18262 ; n18263
g18200 nor n18260 n18263 ; n18264
g18201 nor n18144 n18264 ; n18265
g18202 and n18118 n18130_not ; n18266
g18203 nor n18129 n18130 ; n18267
g18204 nor n18266 n18267 ; n18268
g18205 nor n18265 n18268 ; n18269
g18206 nor n18130 n18269 ; n18270
g18207 and n18104_not n18115 ; n18271
g18208 nor n18116 n18271 ; n18272
g18209 and n18270_not n18272 ; n18273
g18210 nor n18116 n18273 ; n18274
g18211 nor n18102 n18274 ; n18275
g18212 nor n18099 n18275 ; n18276
g18213 nor n18084 n18276 ; n18277
g18214 nor n18081 n18277 ; n18278
g18215 and n18055 n18067_not ; n18279
g18216 nor n18066 n18067 ; n18280
g18217 nor n18279 n18280 ; n18281
g18218 nor n18278 n18281 ; n18282
g18219 nor n18067 n18282 ; n18283
g18220 and n18041 n18053_not ; n18284
g18221 nor n18052 n18053 ; n18285
g18222 nor n18284 n18285 ; n18286
g18223 nor n18283 n18286 ; n18287
g18224 nor n18053 n18287 ; n18288
g18225 and n18027 n18039_not ; n18289
g18226 nor n18038 n18039 ; n18290
g18227 nor n18289 n18290 ; n18291
g18228 nor n18288 n18291 ; n18292
g18229 nor n18039 n18292 ; n18293
g18230 and n18013 n18025_not ; n18294
g18231 nor n18024 n18025 ; n18295
g18232 nor n18294 n18295 ; n18296
g18233 nor n18293 n18296 ; n18297
g18234 nor n18025 n18297 ; n18298
g18235 and n17999 n18011_not ; n18299
g18236 nor n18010 n18011 ; n18300
g18237 nor n18299 n18300 ; n18301
g18238 nor n18298 n18301 ; n18302
g18239 nor n18011 n18302 ; n18303
g18240 and n17985 n17997_not ; n18304
g18241 nor n17996 n17997 ; n18305
g18242 nor n18304 n18305 ; n18306
g18243 nor n18303 n18306 ; n18307
g18244 nor n17997 n18307 ; n18308
g18245 and n17971 n17983_not ; n18309
g18246 nor n17982 n17983 ; n18310
g18247 nor n18309 n18310 ; n18311
g18248 nor n18308 n18311 ; n18312
g18249 nor n17983 n18312 ; n18313
g18250 and n17957 n17969_not ; n18314
g18251 nor n17968 n17969 ; n18315
g18252 nor n18314 n18315 ; n18316
g18253 nor n18313 n18316 ; n18317
g18254 nor n17969 n18317 ; n18318
g18255 and n17943 n17955_not ; n18319
g18256 nor n17954 n17955 ; n18320
g18257 nor n18319 n18320 ; n18321
g18258 nor n18318 n18321 ; n18322
g18259 nor n17955 n18322 ; n18323
g18260 and n17929_not n17940 ; n18324
g18261 nor n17941 n18324 ; n18325
g18262 and n18323_not n18325 ; n18326
g18263 nor n17941 n18326 ; n18327
g18264 nor n17927 n18327 ; n18328
g18265 and n17927 n18327 ; n18329
g18266 nor n18328 n18329 ; n18330
g18267 and n6233 n12370 ; n18331
g18268 and n5663 n12508 ; n18332
g18269 and n5939 n12505 ; n18333
g18270 nor n18332 n18333 ; n18334
g18271 and n18331_not n18334 ; n18335
g18272 and n5666 n13748_not ; n18336
g18273 and n18335 n18336_not ; n18337
g18274 and a[17] n18337_not ; n18338
g18275 and a[17] n18338_not ; n18339
g18276 nor n18337 n18338 ; n18340
g18277 nor n18339 n18340 ; n18341
g18278 and n18330 n18341_not ; n18342
g18279 nor n18328 n18342 ; n18343
g18280 nor n17924 n18343 ; n18344
g18281 and n17924 n18343 ; n18345
g18282 nor n18344 n18345 ; n18346
g18283 and n7101 n13491 ; n18347
g18284 and n6402 n12769 ; n18348
g18285 and n6951 n12889 ; n18349
g18286 nor n18348 n18349 ; n18350
g18287 and n18347_not n18350 ; n18351
g18288 and n6397 n13503_not ; n18352
g18289 and n18351 n18352_not ; n18353
g18290 and a[14] n18353_not ; n18354
g18291 and a[14] n18354_not ; n18355
g18292 nor n18353 n18354 ; n18356
g18293 nor n18355 n18356 ; n18357
g18294 and n18346 n18357_not ; n18358
g18295 nor n18344 n18358 ; n18359
g18296 nor n17921 n18359 ; n18360
g18297 and n17921 n18359 ; n18361
g18298 nor n18360 n18361 ; n18362
g18299 and n7983 n13597 ; n18363
g18300 and n7291 n13521 ; n18364
g18301 and n7632 n13515 ; n18365
g18302 nor n18364 n18365 ; n18366
g18303 and n18363_not n18366 ; n18367
g18304 and n7294 n13612_not ; n18368
g18305 and n18367 n18368_not ; n18369
g18306 and a[11] n18369_not ; n18370
g18307 and a[11] n18370_not ; n18371
g18308 nor n18369 n18370 ; n18372
g18309 nor n18371 n18372 ; n18373
g18310 and n18362 n18373_not ; n18374
g18311 nor n18360 n18374 ; n18375
g18312 nor n17918 n18375 ; n18376
g18313 nor n17915 n18376 ; n18377
g18314 nor n17901 n18377 ; n18378
g18315 and n17901 n18377 ; n18379
g18316 nor n18378 n18379 ; n18380
g18317 and n9331 n13438_not ; n18381
g18318 and n8418 n13627_not ; n18382
g18319 and n8860 n13941 ; n18383
g18320 nor n18382 n18383 ; n18384
g18321 and n18381_not n18384 ; n18385
g18322 and n8421 n14028 ; n18386
g18323 and n18385 n18386_not ; n18387
g18324 and a[8] n18387_not ; n18388
g18325 and a[8] n18388_not ; n18389
g18326 nor n18387 n18388 ; n18390
g18327 nor n18389 n18390 ; n18391
g18328 and n18380 n18391_not ; n18392
g18329 nor n18378 n18392 ; n18393
g18330 nor n17898 n18393 ; n18394
g18331 and n17898 n18393 ; n18395
g18332 nor n18394 n18395 ; n18396
g18333 and n18380 n18392_not ; n18397
g18334 nor n18391 n18392 ; n18398
g18335 nor n18397 n18398 ; n18399
g18336 and n18362 n18374_not ; n18400
g18337 nor n18373 n18374 ; n18401
g18338 nor n18400 n18401 ; n18402
g18339 and n18346 n18358_not ; n18403
g18340 nor n18357 n18358 ; n18404
g18341 nor n18403 n18404 ; n18405
g18342 and n18330 n18342_not ; n18406
g18343 nor n18341 n18342 ; n18407
g18344 nor n18406 n18407 ; n18408
g18345 and n6233 n12505 ; n18409
g18346 and n5663 n12513 ; n18410
g18347 and n5939 n12508 ; n18411
g18348 nor n18410 n18411 ; n18412
g18349 and n18409_not n18412 ; n18413
g18350 and n5666 n14051_not ; n18414
g18351 and n18413 n18414_not ; n18415
g18352 and a[17] n18415_not ; n18416
g18353 nor n18415 n18416 ; n18417
g18354 and a[17] n18416_not ; n18418
g18355 nor n18417 n18418 ; n18419
g18356 and n18323 n18325_not ; n18420
g18357 nor n18326 n18420 ; n18421
g18358 and n18419_not n18421 ; n18422
g18359 nor n18419 n18422 ; n18423
g18360 and n18421 n18422_not ; n18424
g18361 nor n18423 n18424 ; n18425
g18362 and n6233 n12508 ; n18426
g18363 and n5663 n12511 ; n18427
g18364 and n5939 n12513 ; n18428
g18365 nor n18427 n18428 ; n18429
g18366 and n18426_not n18429 ; n18430
g18367 and n5666 n13863 ; n18431
g18368 and n18430 n18431_not ; n18432
g18369 and a[17] n18432_not ; n18433
g18370 nor n18432 n18433 ; n18434
g18371 and a[17] n18433_not ; n18435
g18372 nor n18434 n18435 ; n18436
g18373 nor n18318 n18322 ; n18437
g18374 nor n18321 n18322 ; n18438
g18375 nor n18437 n18438 ; n18439
g18376 nor n18436 n18439 ; n18440
g18377 nor n18436 n18440 ; n18441
g18378 nor n18439 n18440 ; n18442
g18379 nor n18441 n18442 ; n18443
g18380 and n6233 n12513 ; n18444
g18381 and n5663 n12516 ; n18445
g18382 and n5939 n12511 ; n18446
g18383 nor n18445 n18446 ; n18447
g18384 and n18444_not n18447 ; n18448
g18385 and n5666 n14177 ; n18449
g18386 and n18448 n18449_not ; n18450
g18387 and a[17] n18450_not ; n18451
g18388 nor n18450 n18451 ; n18452
g18389 and a[17] n18451_not ; n18453
g18390 nor n18452 n18453 ; n18454
g18391 nor n18313 n18317 ; n18455
g18392 nor n18316 n18317 ; n18456
g18393 nor n18455 n18456 ; n18457
g18394 nor n18454 n18457 ; n18458
g18395 nor n18454 n18458 ; n18459
g18396 nor n18457 n18458 ; n18460
g18397 nor n18459 n18460 ; n18461
g18398 and n6233 n12511 ; n18462
g18399 and n5663 n12519 ; n18463
g18400 and n5939 n12516 ; n18464
g18401 nor n18463 n18464 ; n18465
g18402 and n18462_not n18465 ; n18466
g18403 and n5666 n14233_not ; n18467
g18404 and n18466 n18467_not ; n18468
g18405 and a[17] n18468_not ; n18469
g18406 nor n18468 n18469 ; n18470
g18407 and a[17] n18469_not ; n18471
g18408 nor n18470 n18471 ; n18472
g18409 nor n18308 n18312 ; n18473
g18410 nor n18311 n18312 ; n18474
g18411 nor n18473 n18474 ; n18475
g18412 nor n18472 n18475 ; n18476
g18413 nor n18472 n18476 ; n18477
g18414 nor n18475 n18476 ; n18478
g18415 nor n18477 n18478 ; n18479
g18416 and n6233 n12516 ; n18480
g18417 and n5663 n12522 ; n18481
g18418 and n5939 n12519 ; n18482
g18419 nor n18481 n18482 ; n18483
g18420 and n18480_not n18483 ; n18484
g18421 and n5666 n14443_not ; n18485
g18422 and n18484 n18485_not ; n18486
g18423 and a[17] n18486_not ; n18487
g18424 nor n18486 n18487 ; n18488
g18425 and a[17] n18487_not ; n18489
g18426 nor n18488 n18489 ; n18490
g18427 nor n18303 n18307 ; n18491
g18428 nor n18306 n18307 ; n18492
g18429 nor n18491 n18492 ; n18493
g18430 nor n18490 n18493 ; n18494
g18431 nor n18490 n18494 ; n18495
g18432 nor n18493 n18494 ; n18496
g18433 nor n18495 n18496 ; n18497
g18434 and n6233 n12519 ; n18498
g18435 and n5663 n12525 ; n18499
g18436 and n5939 n12522 ; n18500
g18437 nor n18499 n18500 ; n18501
g18438 and n18498_not n18501 ; n18502
g18439 and n5666 n14454 ; n18503
g18440 and n18502 n18503_not ; n18504
g18441 and a[17] n18504_not ; n18505
g18442 nor n18504 n18505 ; n18506
g18443 and a[17] n18505_not ; n18507
g18444 nor n18506 n18507 ; n18508
g18445 nor n18298 n18302 ; n18509
g18446 nor n18301 n18302 ; n18510
g18447 nor n18509 n18510 ; n18511
g18448 nor n18508 n18511 ; n18512
g18449 nor n18508 n18512 ; n18513
g18450 nor n18511 n18512 ; n18514
g18451 nor n18513 n18514 ; n18515
g18452 and n6233 n12522 ; n18516
g18453 and n5663 n12528 ; n18517
g18454 and n5939 n12525 ; n18518
g18455 nor n18517 n18518 ; n18519
g18456 and n18516_not n18519 ; n18520
g18457 and n5666 n14837 ; n18521
g18458 and n18520 n18521_not ; n18522
g18459 and a[17] n18522_not ; n18523
g18460 nor n18522 n18523 ; n18524
g18461 and a[17] n18523_not ; n18525
g18462 nor n18524 n18525 ; n18526
g18463 nor n18293 n18297 ; n18527
g18464 nor n18296 n18297 ; n18528
g18465 nor n18527 n18528 ; n18529
g18466 nor n18526 n18529 ; n18530
g18467 nor n18526 n18530 ; n18531
g18468 nor n18529 n18530 ; n18532
g18469 nor n18531 n18532 ; n18533
g18470 and n6233 n12525 ; n18534
g18471 and n5663 n12531 ; n18535
g18472 and n5939 n12528 ; n18536
g18473 nor n18535 n18536 ; n18537
g18474 and n18534_not n18537 ; n18538
g18475 and n5666 n14608 ; n18539
g18476 and n18538 n18539_not ; n18540
g18477 and a[17] n18540_not ; n18541
g18478 nor n18540 n18541 ; n18542
g18479 and a[17] n18541_not ; n18543
g18480 nor n18542 n18543 ; n18544
g18481 nor n18288 n18292 ; n18545
g18482 nor n18291 n18292 ; n18546
g18483 nor n18545 n18546 ; n18547
g18484 nor n18544 n18547 ; n18548
g18485 nor n18544 n18548 ; n18549
g18486 nor n18547 n18548 ; n18550
g18487 nor n18549 n18550 ; n18551
g18488 and n6233 n12528 ; n18552
g18489 and n5663 n12534 ; n18553
g18490 and n5939 n12531 ; n18554
g18491 nor n18553 n18554 ; n18555
g18492 and n18552_not n18555 ; n18556
g18493 and n5666 n15003_not ; n18557
g18494 and n18556 n18557_not ; n18558
g18495 and a[17] n18558_not ; n18559
g18496 nor n18558 n18559 ; n18560
g18497 and a[17] n18559_not ; n18561
g18498 nor n18560 n18561 ; n18562
g18499 nor n18283 n18287 ; n18563
g18500 nor n18286 n18287 ; n18564
g18501 nor n18563 n18564 ; n18565
g18502 nor n18562 n18565 ; n18566
g18503 nor n18562 n18566 ; n18567
g18504 nor n18565 n18566 ; n18568
g18505 nor n18567 n18568 ; n18569
g18506 and n6233 n12531 ; n18570
g18507 and n5663 n12537 ; n18571
g18508 and n5939 n12534 ; n18572
g18509 nor n18571 n18572 ; n18573
g18510 and n18570_not n18573 ; n18574
g18511 and n5666 n15255 ; n18575
g18512 and n18574 n18575_not ; n18576
g18513 and a[17] n18576_not ; n18577
g18514 nor n18576 n18577 ; n18578
g18515 and a[17] n18577_not ; n18579
g18516 nor n18578 n18579 ; n18580
g18517 nor n18278 n18282 ; n18581
g18518 nor n18281 n18282 ; n18582
g18519 nor n18581 n18582 ; n18583
g18520 nor n18580 n18583 ; n18584
g18521 nor n18580 n18584 ; n18585
g18522 nor n18583 n18584 ; n18586
g18523 nor n18585 n18586 ; n18587
g18524 and n18084 n18276 ; n18588
g18525 nor n18277 n18588 ; n18589
g18526 and n6233 n12534 ; n18590
g18527 and n5663 n12540 ; n18591
g18528 and n5939 n12537 ; n18592
g18529 nor n18591 n18592 ; n18593
g18530 and n18590_not n18593 ; n18594
g18531 and n5666_not n18594 ; n18595
g18532 and n15096 n18594 ; n18596
g18533 nor n18595 n18596 ; n18597
g18534 and a[17] n18597_not ; n18598
g18535 and a[17]_not n18597 ; n18599
g18536 nor n18598 n18599 ; n18600
g18537 and n18589 n18600_not ; n18601
g18538 and n18102 n18274 ; n18602
g18539 nor n18275 n18602 ; n18603
g18540 and n6233 n12537 ; n18604
g18541 and n5663 n12543 ; n18605
g18542 and n5939 n12540 ; n18606
g18543 nor n18605 n18606 ; n18607
g18544 and n18604_not n18607 ; n18608
g18545 and n5666_not n18608 ; n18609
g18546 and n15385 n18608 ; n18610
g18547 nor n18609 n18610 ; n18611
g18548 and a[17] n18611_not ; n18612
g18549 and a[17]_not n18611 ; n18613
g18550 nor n18612 n18613 ; n18614
g18551 and n18603 n18614_not ; n18615
g18552 and n6233 n12540 ; n18616
g18553 and n5663 n12546 ; n18617
g18554 and n5939 n12543 ; n18618
g18555 nor n18617 n18618 ; n18619
g18556 and n18616_not n18619 ; n18620
g18557 and n5666 n15708_not ; n18621
g18558 and n18620 n18621_not ; n18622
g18559 and a[17] n18622_not ; n18623
g18560 nor n18622 n18623 ; n18624
g18561 and a[17] n18623_not ; n18625
g18562 nor n18624 n18625 ; n18626
g18563 and n18270 n18272_not ; n18627
g18564 nor n18273 n18627 ; n18628
g18565 and n18626_not n18628 ; n18629
g18566 nor n18626 n18629 ; n18630
g18567 and n18628 n18629_not ; n18631
g18568 nor n18630 n18631 ; n18632
g18569 and n6233 n12543 ; n18633
g18570 and n5663 n12549 ; n18634
g18571 and n5939 n12546 ; n18635
g18572 nor n18634 n18635 ; n18636
g18573 and n18633_not n18636 ; n18637
g18574 and n5666 n15724 ; n18638
g18575 and n18637 n18638_not ; n18639
g18576 and a[17] n18639_not ; n18640
g18577 nor n18639 n18640 ; n18641
g18578 and a[17] n18640_not ; n18642
g18579 nor n18641 n18642 ; n18643
g18580 nor n18265 n18269 ; n18644
g18581 nor n18268 n18269 ; n18645
g18582 nor n18644 n18645 ; n18646
g18583 nor n18643 n18646 ; n18647
g18584 nor n18643 n18647 ; n18648
g18585 nor n18646 n18647 ; n18649
g18586 nor n18648 n18649 ; n18650
g18587 and n6233 n12546 ; n18651
g18588 and n5663 n12552 ; n18652
g18589 and n5939 n12549 ; n18653
g18590 nor n18652 n18653 ; n18654
g18591 and n18651_not n18654 ; n18655
g18592 and n5666 n15356_not ; n18656
g18593 and n18655 n18656_not ; n18657
g18594 and a[17] n18657_not ; n18658
g18595 nor n18657 n18658 ; n18659
g18596 and a[17] n18658_not ; n18660
g18597 nor n18659 n18660 ; n18661
g18598 nor n18260 n18264 ; n18662
g18599 nor n18263 n18264 ; n18663
g18600 nor n18662 n18663 ; n18664
g18601 nor n18661 n18664 ; n18665
g18602 nor n18661 n18665 ; n18666
g18603 nor n18664 n18665 ; n18667
g18604 nor n18666 n18667 ; n18668
g18605 and n18161 n18258 ; n18669
g18606 nor n18259 n18669 ; n18670
g18607 and n6233 n12549 ; n18671
g18608 and n5663 n12555 ; n18672
g18609 and n5939 n12552 ; n18673
g18610 nor n18672 n18673 ; n18674
g18611 and n18671_not n18674 ; n18675
g18612 and n5666_not n18675 ; n18676
g18613 and n15764_not n18675 ; n18677
g18614 nor n18676 n18677 ; n18678
g18615 and a[17] n18678_not ; n18679
g18616 and a[17]_not n18678 ; n18680
g18617 nor n18679 n18680 ; n18681
g18618 and n18670 n18681_not ; n18682
g18619 and n18254 n18256_not ; n18683
g18620 nor n18257 n18683 ; n18684
g18621 and n6233 n12552 ; n18685
g18622 and n5663 n12558 ; n18686
g18623 and n5939 n12555 ; n18687
g18624 nor n18686 n18687 ; n18688
g18625 and n18685_not n18688 ; n18689
g18626 and n5666_not n18689 ; n18690
g18627 and n15791 n18689 ; n18691
g18628 nor n18690 n18691 ; n18692
g18629 and a[17] n18692_not ; n18693
g18630 and a[17]_not n18692 ; n18694
g18631 nor n18693 n18694 ; n18695
g18632 and n18684 n18695_not ; n18696
g18633 and n18193 n18252 ; n18697
g18634 nor n18253 n18697 ; n18698
g18635 and n6233 n12555 ; n18699
g18636 and n5663 n12561 ; n18700
g18637 and n5939 n12558 ; n18701
g18638 nor n18700 n18701 ; n18702
g18639 and n18699_not n18702 ; n18703
g18640 and n5666_not n18703 ; n18704
g18641 and n15816 n18703 ; n18705
g18642 nor n18704 n18705 ; n18706
g18643 and a[17] n18706_not ; n18707
g18644 and a[17]_not n18706 ; n18708
g18645 nor n18707 n18708 ; n18709
g18646 and n18698 n18709_not ; n18710
g18647 and n6233 n12558 ; n18711
g18648 and n5663 n12564 ; n18712
g18649 and n5939 n12561 ; n18713
g18650 nor n18712 n18713 ; n18714
g18651 and n18711_not n18714 ; n18715
g18652 and n5666 n15847 ; n18716
g18653 and n18715 n18716_not ; n18717
g18654 and a[17] n18717_not ; n18718
g18655 nor n18717 n18718 ; n18719
g18656 and a[17] n18718_not ; n18720
g18657 nor n18719 n18720 ; n18721
g18658 and n18248 n18250_not ; n18722
g18659 nor n18251 n18722 ; n18723
g18660 and n18721_not n18723 ; n18724
g18661 nor n18721 n18724 ; n18725
g18662 and n18723 n18724_not ; n18726
g18663 nor n18725 n18726 ; n18727
g18664 nor n18235 n18247 ; n18728
g18665 nor n18246 n18247 ; n18729
g18666 nor n18728 n18729 ; n18730
g18667 and n6233 n12561 ; n18731
g18668 and n5663 n12567 ; n18732
g18669 and n5939 n12564 ; n18733
g18670 nor n18732 n18733 ; n18734
g18671 and n18731_not n18734 ; n18735
g18672 and n5666_not n18735 ; n18736
g18673 and n15905 n18735 ; n18737
g18674 nor n18736 n18737 ; n18738
g18675 and a[17] n18738_not ; n18739
g18676 and a[17]_not n18738 ; n18740
g18677 nor n18739 n18740 ; n18741
g18678 nor n18730 n18741 ; n18742
g18679 and n6233 n12564 ; n18743
g18680 and n5663 n12571 ; n18744
g18681 and n5939 n12567 ; n18745
g18682 nor n18744 n18745 ; n18746
g18683 and n18743_not n18746 ; n18747
g18684 and n5666 n15944_not ; n18748
g18685 and n18747 n18748_not ; n18749
g18686 and a[17] n18749_not ; n18750
g18687 nor n18749 n18750 ; n18751
g18688 and a[17] n18750_not ; n18752
g18689 nor n18751 n18752 ; n18753
g18690 and n18219_not n18230 ; n18754
g18691 nor n18231 n18754 ; n18755
g18692 and n18753_not n18755 ; n18756
g18693 nor n18753 n18756 ; n18757
g18694 and n18755 n18756_not ; n18758
g18695 nor n18757 n18758 ; n18759
g18696 and n18216 n18218_not ; n18760
g18697 nor n18219 n18760 ; n18761
g18698 and n6233 n12567 ; n18762
g18699 and n5663 n12574 ; n18763
g18700 and n5939 n12571 ; n18764
g18701 nor n18763 n18764 ; n18765
g18702 and n18762_not n18765 ; n18766
g18703 and n5666_not n18766 ; n18767
g18704 and n15989_not n18766 ; n18768
g18705 nor n18767 n18768 ; n18769
g18706 and a[17] n18769_not ; n18770
g18707 and a[17]_not n18769 ; n18771
g18708 nor n18770 n18771 ; n18772
g18709 and n18761 n18772_not ; n18773
g18710 and n5939 n12581_not ; n18774
g18711 and n6233 n12577 ; n18775
g18712 nor n18774 n18775 ; n18776
g18713 and n5666 n16085_not ; n18777
g18714 and n18776 n18777_not ; n18778
g18715 and a[17] n18778_not ; n18779
g18716 and a[17] n18779_not ; n18780
g18717 nor n18778 n18779 ; n18781
g18718 nor n18780 n18781 ; n18782
g18719 nor n5658 n12581 ; n18783
g18720 and a[17] n18783_not ; n18784
g18721 and n18782_not n18784 ; n18785
g18722 and n6233 n12574 ; n18786
g18723 and n5663 n12581_not ; n18787
g18724 and n5939 n12577 ; n18788
g18725 nor n18787 n18788 ; n18789
g18726 and n18786_not n18789 ; n18790
g18727 and n5666_not n18790 ; n18791
g18728 and n16094 n18790 ; n18792
g18729 nor n18791 n18792 ; n18793
g18730 and a[17] n18793_not ; n18794
g18731 and a[17]_not n18793 ; n18795
g18732 nor n18794 n18795 ; n18796
g18733 and n18785 n18796_not ; n18797
g18734 and n18217 n18797 ; n18798
g18735 and n18797 n18798_not ; n18799
g18736 and n18217 n18798_not ; n18800
g18737 nor n18799 n18800 ; n18801
g18738 and n6233 n12571 ; n18802
g18739 and n5663 n12577 ; n18803
g18740 and n5939 n12574 ; n18804
g18741 nor n18803 n18804 ; n18805
g18742 and n18802_not n18805 ; n18806
g18743 and n5666 n16013 ; n18807
g18744 and n18806 n18807_not ; n18808
g18745 and a[17] n18808_not ; n18809
g18746 and a[17] n18809_not ; n18810
g18747 nor n18808 n18809 ; n18811
g18748 nor n18810 n18811 ; n18812
g18749 nor n18801 n18812 ; n18813
g18750 nor n18798 n18813 ; n18814
g18751 and n18761_not n18772 ; n18815
g18752 nor n18773 n18815 ; n18816
g18753 and n18814_not n18816 ; n18817
g18754 nor n18773 n18817 ; n18818
g18755 nor n18759 n18818 ; n18819
g18756 nor n18756 n18819 ; n18820
g18757 and n18730 n18741 ; n18821
g18758 nor n18742 n18821 ; n18822
g18759 and n18820_not n18822 ; n18823
g18760 nor n18742 n18823 ; n18824
g18761 nor n18727 n18824 ; n18825
g18762 nor n18724 n18825 ; n18826
g18763 and n18698 n18710_not ; n18827
g18764 nor n18709 n18710 ; n18828
g18765 nor n18827 n18828 ; n18829
g18766 nor n18826 n18829 ; n18830
g18767 nor n18710 n18830 ; n18831
g18768 and n18684 n18696_not ; n18832
g18769 nor n18695 n18696 ; n18833
g18770 nor n18832 n18833 ; n18834
g18771 nor n18831 n18834 ; n18835
g18772 nor n18696 n18835 ; n18836
g18773 and n18670_not n18681 ; n18837
g18774 nor n18682 n18837 ; n18838
g18775 and n18836_not n18838 ; n18839
g18776 nor n18682 n18839 ; n18840
g18777 nor n18668 n18840 ; n18841
g18778 nor n18665 n18841 ; n18842
g18779 nor n18650 n18842 ; n18843
g18780 nor n18647 n18843 ; n18844
g18781 nor n18632 n18844 ; n18845
g18782 nor n18629 n18845 ; n18846
g18783 and n18603 n18615_not ; n18847
g18784 nor n18614 n18615 ; n18848
g18785 nor n18847 n18848 ; n18849
g18786 nor n18846 n18849 ; n18850
g18787 nor n18615 n18850 ; n18851
g18788 and n18589_not n18600 ; n18852
g18789 nor n18601 n18852 ; n18853
g18790 and n18851_not n18853 ; n18854
g18791 nor n18601 n18854 ; n18855
g18792 nor n18587 n18855 ; n18856
g18793 nor n18584 n18856 ; n18857
g18794 nor n18569 n18857 ; n18858
g18795 nor n18566 n18858 ; n18859
g18796 nor n18551 n18859 ; n18860
g18797 nor n18548 n18860 ; n18861
g18798 nor n18533 n18861 ; n18862
g18799 nor n18530 n18862 ; n18863
g18800 nor n18515 n18863 ; n18864
g18801 nor n18512 n18864 ; n18865
g18802 nor n18497 n18865 ; n18866
g18803 nor n18494 n18866 ; n18867
g18804 nor n18479 n18867 ; n18868
g18805 nor n18476 n18868 ; n18869
g18806 nor n18461 n18869 ; n18870
g18807 nor n18458 n18870 ; n18871
g18808 nor n18443 n18871 ; n18872
g18809 nor n18440 n18872 ; n18873
g18810 nor n18425 n18873 ; n18874
g18811 nor n18422 n18874 ; n18875
g18812 nor n18408 n18875 ; n18876
g18813 and n18408 n18875 ; n18877
g18814 nor n18876 n18877 ; n18878
g18815 and n7101 n12889 ; n18879
g18816 and n6402 n12502 ; n18880
g18817 and n6951 n12769 ; n18881
g18818 nor n18880 n18881 ; n18882
g18819 and n18879_not n18882 ; n18883
g18820 and n6397 n12895 ; n18884
g18821 and n18883 n18884_not ; n18885
g18822 and a[14] n18885_not ; n18886
g18823 and a[14] n18886_not ; n18887
g18824 nor n18885 n18886 ; n18888
g18825 nor n18887 n18888 ; n18889
g18826 and n18878 n18889_not ; n18890
g18827 nor n18876 n18890 ; n18891
g18828 nor n18405 n18891 ; n18892
g18829 and n18405 n18891 ; n18893
g18830 nor n18892 n18893 ; n18894
g18831 and n7983 n13515 ; n18895
g18832 and n7291 n13518 ; n18896
g18833 and n7632 n13521 ; n18897
g18834 nor n18896 n18897 ; n18898
g18835 and n18895_not n18898 ; n18899
g18836 and n7294 n13541 ; n18900
g18837 and n18899 n18900_not ; n18901
g18838 and a[11] n18901_not ; n18902
g18839 and a[11] n18902_not ; n18903
g18840 nor n18901 n18902 ; n18904
g18841 nor n18903 n18904 ; n18905
g18842 and n18894 n18905_not ; n18906
g18843 nor n18892 n18906 ; n18907
g18844 nor n18402 n18907 ; n18908
g18845 and n18402 n18907 ; n18909
g18846 nor n18908 n18909 ; n18910
g18847 and n9331 n13627_not ; n18911
g18848 and n8418 n13630 ; n18912
g18849 and n8860 n13633 ; n18913
g18850 nor n18912 n18913 ; n18914
g18851 and n18911_not n18914 ; n18915
g18852 and n8421 n13654_not ; n18916
g18853 and n18915 n18916_not ; n18917
g18854 and a[8] n18917_not ; n18918
g18855 and a[8] n18918_not ; n18919
g18856 nor n18917 n18918 ; n18920
g18857 nor n18919 n18920 ; n18921
g18858 and n18910 n18921_not ; n18922
g18859 nor n18908 n18922 ; n18923
g18860 and n9331 n13941 ; n18924
g18861 and n8418 n13633 ; n18925
g18862 and n8860 n13627_not ; n18926
g18863 nor n18925 n18926 ; n18927
g18864 and n18924_not n18927 ; n18928
g18865 and n8421 n14136 ; n18929
g18866 and n18928 n18929_not ; n18930
g18867 and a[8] n18930_not ; n18931
g18868 and a[8] n18931_not ; n18932
g18869 nor n18930 n18931 ; n18933
g18870 nor n18932 n18933 ; n18934
g18871 nor n18923 n18934 ; n18935
g18872 nor n18923 n18935 ; n18936
g18873 nor n18934 n18935 ; n18937
g18874 nor n18936 n18937 ; n18938
g18875 and n17918 n18375 ; n18939
g18876 nor n18376 n18939 ; n18940
g18877 and n18938_not n18940 ; n18941
g18878 nor n18935 n18941 ; n18942
g18879 nor n18399 n18942 ; n18943
g18880 nor n18399 n18943 ; n18944
g18881 nor n18942 n18943 ; n18945
g18882 nor n18944 n18945 ; n18946
g18883 and n18894 n18906_not ; n18947
g18884 nor n18905 n18906 ; n18948
g18885 nor n18947 n18948 ; n18949
g18886 and n18878 n18890_not ; n18950
g18887 nor n18889 n18890 ; n18951
g18888 nor n18950 n18951 ; n18952
g18889 and n18425 n18873 ; n18953
g18890 nor n18874 n18953 ; n18954
g18891 and n7101 n12769 ; n18955
g18892 and n6402 n12370 ; n18956
g18893 and n6951 n12502 ; n18957
g18894 nor n18956 n18957 ; n18958
g18895 and n18955_not n18958 ; n18959
g18896 and n6397_not n18959 ; n18960
g18897 and n12999_not n18959 ; n18961
g18898 nor n18960 n18961 ; n18962
g18899 and a[14] n18962_not ; n18963
g18900 and a[14]_not n18962 ; n18964
g18901 nor n18963 n18964 ; n18965
g18902 and n18954 n18965_not ; n18966
g18903 and n18443 n18871 ; n18967
g18904 nor n18872 n18967 ; n18968
g18905 and n7101 n12502 ; n18969
g18906 and n6402 n12505 ; n18970
g18907 and n6951 n12370 ; n18971
g18908 nor n18970 n18971 ; n18972
g18909 and n18969_not n18972 ; n18973
g18910 and n6397_not n18973 ; n18974
g18911 and n13736 n18973 ; n18975
g18912 nor n18974 n18975 ; n18976
g18913 and a[14] n18976_not ; n18977
g18914 and a[14]_not n18976 ; n18978
g18915 nor n18977 n18978 ; n18979
g18916 and n18968 n18979_not ; n18980
g18917 and n18461 n18869 ; n18981
g18918 nor n18870 n18981 ; n18982
g18919 and n7101 n12370 ; n18983
g18920 and n6402 n12508 ; n18984
g18921 and n6951 n12505 ; n18985
g18922 nor n18984 n18985 ; n18986
g18923 and n18983_not n18986 ; n18987
g18924 and n6397_not n18987 ; n18988
g18925 and n13748 n18987 ; n18989
g18926 nor n18988 n18989 ; n18990
g18927 and a[14] n18990_not ; n18991
g18928 and a[14]_not n18990 ; n18992
g18929 nor n18991 n18992 ; n18993
g18930 and n18982 n18993_not ; n18994
g18931 and n18479 n18867 ; n18995
g18932 nor n18868 n18995 ; n18996
g18933 and n7101 n12505 ; n18997
g18934 and n6402 n12513 ; n18998
g18935 and n6951 n12508 ; n18999
g18936 nor n18998 n18999 ; n19000
g18937 and n18997_not n19000 ; n19001
g18938 and n6397_not n19001 ; n19002
g18939 and n14051 n19001 ; n19003
g18940 nor n19002 n19003 ; n19004
g18941 and a[14] n19004_not ; n19005
g18942 and a[14]_not n19004 ; n19006
g18943 nor n19005 n19006 ; n19007
g18944 and n18996 n19007_not ; n19008
g18945 and n18497 n18865 ; n19009
g18946 nor n18866 n19009 ; n19010
g18947 and n7101 n12508 ; n19011
g18948 and n6402 n12511 ; n19012
g18949 and n6951 n12513 ; n19013
g18950 nor n19012 n19013 ; n19014
g18951 and n19011_not n19014 ; n19015
g18952 and n6397_not n19015 ; n19016
g18953 and n13863_not n19015 ; n19017
g18954 nor n19016 n19017 ; n19018
g18955 and a[14] n19018_not ; n19019
g18956 and a[14]_not n19018 ; n19020
g18957 nor n19019 n19020 ; n19021
g18958 and n19010 n19021_not ; n19022
g18959 and n18515 n18863 ; n19023
g18960 nor n18864 n19023 ; n19024
g18961 and n7101 n12513 ; n19025
g18962 and n6402 n12516 ; n19026
g18963 and n6951 n12511 ; n19027
g18964 nor n19026 n19027 ; n19028
g18965 and n19025_not n19028 ; n19029
g18966 and n6397_not n19029 ; n19030
g18967 and n14177_not n19029 ; n19031
g18968 nor n19030 n19031 ; n19032
g18969 and a[14] n19032_not ; n19033
g18970 and a[14]_not n19032 ; n19034
g18971 nor n19033 n19034 ; n19035
g18972 and n19024 n19035_not ; n19036
g18973 and n18533 n18861 ; n19037
g18974 nor n18862 n19037 ; n19038
g18975 and n7101 n12511 ; n19039
g18976 and n6402 n12519 ; n19040
g18977 and n6951 n12516 ; n19041
g18978 nor n19040 n19041 ; n19042
g18979 and n19039_not n19042 ; n19043
g18980 and n6397_not n19043 ; n19044
g18981 and n14233 n19043 ; n19045
g18982 nor n19044 n19045 ; n19046
g18983 and a[14] n19046_not ; n19047
g18984 and a[14]_not n19046 ; n19048
g18985 nor n19047 n19048 ; n19049
g18986 and n19038 n19049_not ; n19050
g18987 and n18551 n18859 ; n19051
g18988 nor n18860 n19051 ; n19052
g18989 and n7101 n12516 ; n19053
g18990 and n6402 n12522 ; n19054
g18991 and n6951 n12519 ; n19055
g18992 nor n19054 n19055 ; n19056
g18993 and n19053_not n19056 ; n19057
g18994 and n6397_not n19057 ; n19058
g18995 and n14443 n19057 ; n19059
g18996 nor n19058 n19059 ; n19060
g18997 and a[14] n19060_not ; n19061
g18998 and a[14]_not n19060 ; n19062
g18999 nor n19061 n19062 ; n19063
g19000 and n19052 n19063_not ; n19064
g19001 and n18569 n18857 ; n19065
g19002 nor n18858 n19065 ; n19066
g19003 and n7101 n12519 ; n19067
g19004 and n6402 n12525 ; n19068
g19005 and n6951 n12522 ; n19069
g19006 nor n19068 n19069 ; n19070
g19007 and n19067_not n19070 ; n19071
g19008 and n6397_not n19071 ; n19072
g19009 and n14454_not n19071 ; n19073
g19010 nor n19072 n19073 ; n19074
g19011 and a[14] n19074_not ; n19075
g19012 and a[14]_not n19074 ; n19076
g19013 nor n19075 n19076 ; n19077
g19014 and n19066 n19077_not ; n19078
g19015 and n18587 n18855 ; n19079
g19016 nor n18856 n19079 ; n19080
g19017 and n7101 n12522 ; n19081
g19018 and n6402 n12528 ; n19082
g19019 and n6951 n12525 ; n19083
g19020 nor n19082 n19083 ; n19084
g19021 and n19081_not n19084 ; n19085
g19022 and n6397_not n19085 ; n19086
g19023 and n14837_not n19085 ; n19087
g19024 nor n19086 n19087 ; n19088
g19025 and a[14] n19088_not ; n19089
g19026 and a[14]_not n19088 ; n19090
g19027 nor n19089 n19090 ; n19091
g19028 and n19080 n19091_not ; n19092
g19029 and n7101 n12525 ; n19093
g19030 and n6402 n12531 ; n19094
g19031 and n6951 n12528 ; n19095
g19032 nor n19094 n19095 ; n19096
g19033 and n19093_not n19096 ; n19097
g19034 and n6397 n14608 ; n19098
g19035 and n19097 n19098_not ; n19099
g19036 and a[14] n19099_not ; n19100
g19037 nor n19099 n19100 ; n19101
g19038 and a[14] n19100_not ; n19102
g19039 nor n19101 n19102 ; n19103
g19040 and n18851 n18853_not ; n19104
g19041 nor n18854 n19104 ; n19105
g19042 and n19103_not n19105 ; n19106
g19043 nor n19103 n19106 ; n19107
g19044 and n19105 n19106_not ; n19108
g19045 nor n19107 n19108 ; n19109
g19046 and n7101 n12528 ; n19110
g19047 and n6402 n12534 ; n19111
g19048 and n6951 n12531 ; n19112
g19049 nor n19111 n19112 ; n19113
g19050 and n19110_not n19113 ; n19114
g19051 and n6397 n15003_not ; n19115
g19052 and n19114 n19115_not ; n19116
g19053 and a[14] n19116_not ; n19117
g19054 nor n19116 n19117 ; n19118
g19055 and a[14] n19117_not ; n19119
g19056 nor n19118 n19119 ; n19120
g19057 nor n18846 n18850 ; n19121
g19058 nor n18849 n18850 ; n19122
g19059 nor n19121 n19122 ; n19123
g19060 nor n19120 n19123 ; n19124
g19061 nor n19120 n19124 ; n19125
g19062 nor n19123 n19124 ; n19126
g19063 nor n19125 n19126 ; n19127
g19064 and n18632 n18844 ; n19128
g19065 nor n18845 n19128 ; n19129
g19066 and n7101 n12531 ; n19130
g19067 and n6402 n12537 ; n19131
g19068 and n6951 n12534 ; n19132
g19069 nor n19131 n19132 ; n19133
g19070 and n19130_not n19133 ; n19134
g19071 and n6397_not n19134 ; n19135
g19072 and n15255_not n19134 ; n19136
g19073 nor n19135 n19136 ; n19137
g19074 and a[14] n19137_not ; n19138
g19075 and a[14]_not n19137 ; n19139
g19076 nor n19138 n19139 ; n19140
g19077 and n19129 n19140_not ; n19141
g19078 and n18650 n18842 ; n19142
g19079 nor n18843 n19142 ; n19143
g19080 and n7101 n12534 ; n19144
g19081 and n6402 n12540 ; n19145
g19082 and n6951 n12537 ; n19146
g19083 nor n19145 n19146 ; n19147
g19084 and n19144_not n19147 ; n19148
g19085 and n6397_not n19148 ; n19149
g19086 and n15096 n19148 ; n19150
g19087 nor n19149 n19150 ; n19151
g19088 and a[14] n19151_not ; n19152
g19089 and a[14]_not n19151 ; n19153
g19090 nor n19152 n19153 ; n19154
g19091 and n19143 n19154_not ; n19155
g19092 and n18668 n18840 ; n19156
g19093 nor n18841 n19156 ; n19157
g19094 and n7101 n12537 ; n19158
g19095 and n6402 n12543 ; n19159
g19096 and n6951 n12540 ; n19160
g19097 nor n19159 n19160 ; n19161
g19098 and n19158_not n19161 ; n19162
g19099 and n6397_not n19162 ; n19163
g19100 and n15385 n19162 ; n19164
g19101 nor n19163 n19164 ; n19165
g19102 and a[14] n19165_not ; n19166
g19103 and a[14]_not n19165 ; n19167
g19104 nor n19166 n19167 ; n19168
g19105 and n19157 n19168_not ; n19169
g19106 and n7101 n12540 ; n19170
g19107 and n6402 n12546 ; n19171
g19108 and n6951 n12543 ; n19172
g19109 nor n19171 n19172 ; n19173
g19110 and n19170_not n19173 ; n19174
g19111 and n6397 n15708_not ; n19175
g19112 and n19174 n19175_not ; n19176
g19113 and a[14] n19176_not ; n19177
g19114 nor n19176 n19177 ; n19178
g19115 and a[14] n19177_not ; n19179
g19116 nor n19178 n19179 ; n19180
g19117 and n18836 n18838_not ; n19181
g19118 nor n18839 n19181 ; n19182
g19119 and n19180_not n19182 ; n19183
g19120 nor n19180 n19183 ; n19184
g19121 and n19182 n19183_not ; n19185
g19122 nor n19184 n19185 ; n19186
g19123 and n7101 n12543 ; n19187
g19124 and n6402 n12549 ; n19188
g19125 and n6951 n12546 ; n19189
g19126 nor n19188 n19189 ; n19190
g19127 and n19187_not n19190 ; n19191
g19128 and n6397 n15724 ; n19192
g19129 and n19191 n19192_not ; n19193
g19130 and a[14] n19193_not ; n19194
g19131 nor n19193 n19194 ; n19195
g19132 and a[14] n19194_not ; n19196
g19133 nor n19195 n19196 ; n19197
g19134 nor n18831 n18835 ; n19198
g19135 nor n18834 n18835 ; n19199
g19136 nor n19198 n19199 ; n19200
g19137 nor n19197 n19200 ; n19201
g19138 nor n19197 n19201 ; n19202
g19139 nor n19200 n19201 ; n19203
g19140 nor n19202 n19203 ; n19204
g19141 and n7101 n12546 ; n19205
g19142 and n6402 n12552 ; n19206
g19143 and n6951 n12549 ; n19207
g19144 nor n19206 n19207 ; n19208
g19145 and n19205_not n19208 ; n19209
g19146 and n6397 n15356_not ; n19210
g19147 and n19209 n19210_not ; n19211
g19148 and a[14] n19211_not ; n19212
g19149 nor n19211 n19212 ; n19213
g19150 and a[14] n19212_not ; n19214
g19151 nor n19213 n19214 ; n19215
g19152 nor n18826 n18830 ; n19216
g19153 nor n18829 n18830 ; n19217
g19154 nor n19216 n19217 ; n19218
g19155 nor n19215 n19218 ; n19219
g19156 nor n19215 n19219 ; n19220
g19157 nor n19218 n19219 ; n19221
g19158 nor n19220 n19221 ; n19222
g19159 and n18727 n18824 ; n19223
g19160 nor n18825 n19223 ; n19224
g19161 and n7101 n12549 ; n19225
g19162 and n6402 n12555 ; n19226
g19163 and n6951 n12552 ; n19227
g19164 nor n19226 n19227 ; n19228
g19165 and n19225_not n19228 ; n19229
g19166 and n6397_not n19229 ; n19230
g19167 and n15764_not n19229 ; n19231
g19168 nor n19230 n19231 ; n19232
g19169 and a[14] n19232_not ; n19233
g19170 and a[14]_not n19232 ; n19234
g19171 nor n19233 n19234 ; n19235
g19172 and n19224 n19235_not ; n19236
g19173 and n18820 n18822_not ; n19237
g19174 nor n18823 n19237 ; n19238
g19175 and n7101 n12552 ; n19239
g19176 and n6402 n12558 ; n19240
g19177 and n6951 n12555 ; n19241
g19178 nor n19240 n19241 ; n19242
g19179 and n19239_not n19242 ; n19243
g19180 and n6397_not n19243 ; n19244
g19181 and n15791 n19243 ; n19245
g19182 nor n19244 n19245 ; n19246
g19183 and a[14] n19246_not ; n19247
g19184 and a[14]_not n19246 ; n19248
g19185 nor n19247 n19248 ; n19249
g19186 and n19238 n19249_not ; n19250
g19187 and n18759 n18818 ; n19251
g19188 nor n18819 n19251 ; n19252
g19189 and n7101 n12555 ; n19253
g19190 and n6402 n12561 ; n19254
g19191 and n6951 n12558 ; n19255
g19192 nor n19254 n19255 ; n19256
g19193 and n19253_not n19256 ; n19257
g19194 and n6397_not n19257 ; n19258
g19195 and n15816 n19257 ; n19259
g19196 nor n19258 n19259 ; n19260
g19197 and a[14] n19260_not ; n19261
g19198 and a[14]_not n19260 ; n19262
g19199 nor n19261 n19262 ; n19263
g19200 and n19252 n19263_not ; n19264
g19201 and n7101 n12558 ; n19265
g19202 and n6402 n12564 ; n19266
g19203 and n6951 n12561 ; n19267
g19204 nor n19266 n19267 ; n19268
g19205 and n19265_not n19268 ; n19269
g19206 and n6397 n15847 ; n19270
g19207 and n19269 n19270_not ; n19271
g19208 and a[14] n19271_not ; n19272
g19209 nor n19271 n19272 ; n19273
g19210 and a[14] n19272_not ; n19274
g19211 nor n19273 n19274 ; n19275
g19212 and n18814 n18816_not ; n19276
g19213 nor n18817 n19276 ; n19277
g19214 and n19275_not n19277 ; n19278
g19215 nor n19275 n19278 ; n19279
g19216 and n19277 n19278_not ; n19280
g19217 nor n19279 n19280 ; n19281
g19218 nor n18801 n18813 ; n19282
g19219 nor n18812 n18813 ; n19283
g19220 nor n19282 n19283 ; n19284
g19221 and n7101 n12561 ; n19285
g19222 and n6402 n12567 ; n19286
g19223 and n6951 n12564 ; n19287
g19224 nor n19286 n19287 ; n19288
g19225 and n19285_not n19288 ; n19289
g19226 and n6397_not n19289 ; n19290
g19227 and n15905 n19289 ; n19291
g19228 nor n19290 n19291 ; n19292
g19229 and a[14] n19292_not ; n19293
g19230 and a[14]_not n19292 ; n19294
g19231 nor n19293 n19294 ; n19295
g19232 nor n19284 n19295 ; n19296
g19233 and n7101 n12564 ; n19297
g19234 and n6402 n12571 ; n19298
g19235 and n6951 n12567 ; n19299
g19236 nor n19298 n19299 ; n19300
g19237 and n19297_not n19300 ; n19301
g19238 and n6397 n15944_not ; n19302
g19239 and n19301 n19302_not ; n19303
g19240 and a[14] n19303_not ; n19304
g19241 nor n19303 n19304 ; n19305
g19242 and a[14] n19304_not ; n19306
g19243 nor n19305 n19306 ; n19307
g19244 and n18785_not n18796 ; n19308
g19245 nor n18797 n19308 ; n19309
g19246 and n19307_not n19309 ; n19310
g19247 nor n19307 n19310 ; n19311
g19248 and n19309 n19310_not ; n19312
g19249 nor n19311 n19312 ; n19313
g19250 and n18782 n18784_not ; n19314
g19251 nor n18785 n19314 ; n19315
g19252 and n7101 n12567 ; n19316
g19253 and n6402 n12574 ; n19317
g19254 and n6951 n12571 ; n19318
g19255 nor n19317 n19318 ; n19319
g19256 and n19316_not n19319 ; n19320
g19257 and n6397_not n19320 ; n19321
g19258 and n15989_not n19320 ; n19322
g19259 nor n19321 n19322 ; n19323
g19260 and a[14] n19323_not ; n19324
g19261 and a[14]_not n19323 ; n19325
g19262 nor n19324 n19325 ; n19326
g19263 and n19315 n19326_not ; n19327
g19264 and n6951 n12581_not ; n19328
g19265 and n7101 n12577 ; n19329
g19266 nor n19328 n19329 ; n19330
g19267 and n6397 n16085_not ; n19331
g19268 and n19330 n19331_not ; n19332
g19269 and a[14] n19332_not ; n19333
g19270 and a[14] n19333_not ; n19334
g19271 nor n19332 n19333 ; n19335
g19272 nor n19334 n19335 ; n19336
g19273 nor n6393 n12581 ; n19337
g19274 and a[14] n19337_not ; n19338
g19275 and n19336_not n19338 ; n19339
g19276 and n7101 n12574 ; n19340
g19277 and n6402 n12581_not ; n19341
g19278 and n6951 n12577 ; n19342
g19279 nor n19341 n19342 ; n19343
g19280 and n19340_not n19343 ; n19344
g19281 and n6397_not n19344 ; n19345
g19282 and n16094 n19344 ; n19346
g19283 nor n19345 n19346 ; n19347
g19284 and a[14] n19347_not ; n19348
g19285 and a[14]_not n19347 ; n19349
g19286 nor n19348 n19349 ; n19350
g19287 and n19339 n19350_not ; n19351
g19288 and n18783 n19351 ; n19352
g19289 and n19351 n19352_not ; n19353
g19290 and n18783 n19352_not ; n19354
g19291 nor n19353 n19354 ; n19355
g19292 and n7101 n12571 ; n19356
g19293 and n6402 n12577 ; n19357
g19294 and n6951 n12574 ; n19358
g19295 nor n19357 n19358 ; n19359
g19296 and n19356_not n19359 ; n19360
g19297 and n6397 n16013 ; n19361
g19298 and n19360 n19361_not ; n19362
g19299 and a[14] n19362_not ; n19363
g19300 and a[14] n19363_not ; n19364
g19301 nor n19362 n19363 ; n19365
g19302 nor n19364 n19365 ; n19366
g19303 nor n19355 n19366 ; n19367
g19304 nor n19352 n19367 ; n19368
g19305 and n19315_not n19326 ; n19369
g19306 nor n19327 n19369 ; n19370
g19307 and n19368_not n19370 ; n19371
g19308 nor n19327 n19371 ; n19372
g19309 nor n19313 n19372 ; n19373
g19310 nor n19310 n19373 ; n19374
g19311 and n19284 n19295 ; n19375
g19312 nor n19296 n19375 ; n19376
g19313 and n19374_not n19376 ; n19377
g19314 nor n19296 n19377 ; n19378
g19315 nor n19281 n19378 ; n19379
g19316 nor n19278 n19379 ; n19380
g19317 and n19252 n19264_not ; n19381
g19318 nor n19263 n19264 ; n19382
g19319 nor n19381 n19382 ; n19383
g19320 nor n19380 n19383 ; n19384
g19321 nor n19264 n19384 ; n19385
g19322 and n19238 n19250_not ; n19386
g19323 nor n19249 n19250 ; n19387
g19324 nor n19386 n19387 ; n19388
g19325 nor n19385 n19388 ; n19389
g19326 nor n19250 n19389 ; n19390
g19327 and n19224_not n19235 ; n19391
g19328 nor n19236 n19391 ; n19392
g19329 and n19390_not n19392 ; n19393
g19330 nor n19236 n19393 ; n19394
g19331 nor n19222 n19394 ; n19395
g19332 nor n19219 n19395 ; n19396
g19333 nor n19204 n19396 ; n19397
g19334 nor n19201 n19397 ; n19398
g19335 nor n19186 n19398 ; n19399
g19336 nor n19183 n19399 ; n19400
g19337 and n19157 n19169_not ; n19401
g19338 nor n19168 n19169 ; n19402
g19339 nor n19401 n19402 ; n19403
g19340 nor n19400 n19403 ; n19404
g19341 nor n19169 n19404 ; n19405
g19342 and n19143 n19155_not ; n19406
g19343 nor n19154 n19155 ; n19407
g19344 nor n19406 n19407 ; n19408
g19345 nor n19405 n19408 ; n19409
g19346 nor n19155 n19409 ; n19410
g19347 and n19129_not n19140 ; n19411
g19348 nor n19141 n19411 ; n19412
g19349 and n19410_not n19412 ; n19413
g19350 nor n19141 n19413 ; n19414
g19351 nor n19127 n19414 ; n19415
g19352 nor n19124 n19415 ; n19416
g19353 nor n19109 n19416 ; n19417
g19354 nor n19106 n19417 ; n19418
g19355 and n19080 n19092_not ; n19419
g19356 nor n19091 n19092 ; n19420
g19357 nor n19419 n19420 ; n19421
g19358 nor n19418 n19421 ; n19422
g19359 nor n19092 n19422 ; n19423
g19360 and n19066 n19078_not ; n19424
g19361 nor n19077 n19078 ; n19425
g19362 nor n19424 n19425 ; n19426
g19363 nor n19423 n19426 ; n19427
g19364 nor n19078 n19427 ; n19428
g19365 and n19052 n19064_not ; n19429
g19366 nor n19063 n19064 ; n19430
g19367 nor n19429 n19430 ; n19431
g19368 nor n19428 n19431 ; n19432
g19369 nor n19064 n19432 ; n19433
g19370 and n19038 n19050_not ; n19434
g19371 nor n19049 n19050 ; n19435
g19372 nor n19434 n19435 ; n19436
g19373 nor n19433 n19436 ; n19437
g19374 nor n19050 n19437 ; n19438
g19375 and n19024 n19036_not ; n19439
g19376 nor n19035 n19036 ; n19440
g19377 nor n19439 n19440 ; n19441
g19378 nor n19438 n19441 ; n19442
g19379 nor n19036 n19442 ; n19443
g19380 and n19010 n19022_not ; n19444
g19381 nor n19021 n19022 ; n19445
g19382 nor n19444 n19445 ; n19446
g19383 nor n19443 n19446 ; n19447
g19384 nor n19022 n19447 ; n19448
g19385 and n18996 n19008_not ; n19449
g19386 nor n19007 n19008 ; n19450
g19387 nor n19449 n19450 ; n19451
g19388 nor n19448 n19451 ; n19452
g19389 nor n19008 n19452 ; n19453
g19390 and n18982 n18994_not ; n19454
g19391 nor n18993 n18994 ; n19455
g19392 nor n19454 n19455 ; n19456
g19393 nor n19453 n19456 ; n19457
g19394 nor n18994 n19457 ; n19458
g19395 and n18968 n18980_not ; n19459
g19396 nor n18979 n18980 ; n19460
g19397 nor n19459 n19460 ; n19461
g19398 nor n19458 n19461 ; n19462
g19399 nor n18980 n19462 ; n19463
g19400 and n18954_not n18965 ; n19464
g19401 nor n18966 n19464 ; n19465
g19402 and n19463_not n19465 ; n19466
g19403 nor n18966 n19466 ; n19467
g19404 nor n18952 n19467 ; n19468
g19405 and n18952 n19467 ; n19469
g19406 nor n19468 n19469 ; n19470
g19407 and n7983 n13521 ; n19471
g19408 and n7291 n13491 ; n19472
g19409 and n7632 n13518 ; n19473
g19410 nor n19472 n19473 ; n19474
g19411 and n19471_not n19474 ; n19475
g19412 and n7294 n13909_not ; n19476
g19413 and n19475 n19476_not ; n19477
g19414 and a[11] n19477_not ; n19478
g19415 and a[11] n19478_not ; n19479
g19416 nor n19477 n19478 ; n19480
g19417 nor n19479 n19480 ; n19481
g19418 and n19470 n19481_not ; n19482
g19419 nor n19468 n19482 ; n19483
g19420 nor n18949 n19483 ; n19484
g19421 and n18949 n19483 ; n19485
g19422 nor n19484 n19485 ; n19486
g19423 and n9331 n13633 ; n19487
g19424 and n8418 n13597 ; n19488
g19425 and n8860 n13630 ; n19489
g19426 nor n19488 n19489 ; n19490
g19427 and n19487_not n19490 ; n19491
g19428 and n8421 n13929 ; n19492
g19429 and n19491 n19492_not ; n19493
g19430 and a[8] n19493_not ; n19494
g19431 and a[8] n19494_not ; n19495
g19432 nor n19493 n19494 ; n19496
g19433 nor n19495 n19496 ; n19497
g19434 and n19486 n19497_not ; n19498
g19435 nor n19484 n19498 ; n19499
g19436 nor n13438 n15076 ; n19500
g19437 and n9867 n13941 ; n19501
g19438 nor n19500 n19501 ; n19502
g19439 and n9870_not n19502 ; n19503
g19440 and n13951 n19502 ; n19504
g19441 nor n19503 n19504 ; n19505
g19442 and a[5] n19505_not ; n19506
g19443 and a[5]_not n19505 ; n19507
g19444 nor n19506 n19507 ; n19508
g19445 nor n19499 n19508 ; n19509
g19446 and n18910 n18922_not ; n19510
g19447 nor n18921 n18922 ; n19511
g19448 nor n19510 n19511 ; n19512
g19449 and n19499 n19508 ; n19513
g19450 nor n19509 n19513 ; n19514
g19451 and n19512_not n19514 ; n19515
g19452 nor n19509 n19515 ; n19516
g19453 and n18938 n18940_not ; n19517
g19454 nor n18941 n19517 ; n19518
g19455 and n19516_not n19518 ; n19519
g19456 nor n19512 n19515 ; n19520
g19457 and n19514 n19515_not ; n19521
g19458 nor n19520 n19521 ; n19522
g19459 and n19486 n19498_not ; n19523
g19460 nor n19497 n19498 ; n19524
g19461 nor n19523 n19524 ; n19525
g19462 and n19470 n19482_not ; n19526
g19463 nor n19481 n19482 ; n19527
g19464 nor n19526 n19527 ; n19528
g19465 and n7983 n13518 ; n19529
g19466 and n7291 n12889 ; n19530
g19467 and n7632 n13491 ; n19531
g19468 nor n19530 n19531 ; n19532
g19469 and n19529_not n19532 ; n19533
g19470 and n7294 n13584 ; n19534
g19471 and n19533 n19534_not ; n19535
g19472 and a[11] n19535_not ; n19536
g19473 nor n19535 n19536 ; n19537
g19474 and a[11] n19536_not ; n19538
g19475 nor n19537 n19538 ; n19539
g19476 and n19463 n19465_not ; n19540
g19477 nor n19466 n19540 ; n19541
g19478 and n19539_not n19541 ; n19542
g19479 nor n19539 n19542 ; n19543
g19480 and n19541 n19542_not ; n19544
g19481 nor n19543 n19544 ; n19545
g19482 and n7983 n13491 ; n19546
g19483 and n7291 n12769 ; n19547
g19484 and n7632 n12889 ; n19548
g19485 nor n19547 n19548 ; n19549
g19486 and n19546_not n19549 ; n19550
g19487 and n7294 n13503_not ; n19551
g19488 and n19550 n19551_not ; n19552
g19489 and a[11] n19552_not ; n19553
g19490 nor n19552 n19553 ; n19554
g19491 and a[11] n19553_not ; n19555
g19492 nor n19554 n19555 ; n19556
g19493 nor n19458 n19462 ; n19557
g19494 nor n19461 n19462 ; n19558
g19495 nor n19557 n19558 ; n19559
g19496 nor n19556 n19559 ; n19560
g19497 nor n19556 n19560 ; n19561
g19498 nor n19559 n19560 ; n19562
g19499 nor n19561 n19562 ; n19563
g19500 and n7983 n12889 ; n19564
g19501 and n7291 n12502 ; n19565
g19502 and n7632 n12769 ; n19566
g19503 nor n19565 n19566 ; n19567
g19504 and n19564_not n19567 ; n19568
g19505 and n7294 n12895 ; n19569
g19506 and n19568 n19569_not ; n19570
g19507 and a[11] n19570_not ; n19571
g19508 nor n19570 n19571 ; n19572
g19509 and a[11] n19571_not ; n19573
g19510 nor n19572 n19573 ; n19574
g19511 nor n19453 n19457 ; n19575
g19512 nor n19456 n19457 ; n19576
g19513 nor n19575 n19576 ; n19577
g19514 nor n19574 n19577 ; n19578
g19515 nor n19574 n19578 ; n19579
g19516 nor n19577 n19578 ; n19580
g19517 nor n19579 n19580 ; n19581
g19518 and n7983 n12769 ; n19582
g19519 and n7291 n12370 ; n19583
g19520 and n7632 n12502 ; n19584
g19521 nor n19583 n19584 ; n19585
g19522 and n19582_not n19585 ; n19586
g19523 and n7294 n12999 ; n19587
g19524 and n19586 n19587_not ; n19588
g19525 and a[11] n19588_not ; n19589
g19526 nor n19588 n19589 ; n19590
g19527 and a[11] n19589_not ; n19591
g19528 nor n19590 n19591 ; n19592
g19529 nor n19448 n19452 ; n19593
g19530 nor n19451 n19452 ; n19594
g19531 nor n19593 n19594 ; n19595
g19532 nor n19592 n19595 ; n19596
g19533 nor n19592 n19596 ; n19597
g19534 nor n19595 n19596 ; n19598
g19535 nor n19597 n19598 ; n19599
g19536 and n7983 n12502 ; n19600
g19537 and n7291 n12505 ; n19601
g19538 and n7632 n12370 ; n19602
g19539 nor n19601 n19602 ; n19603
g19540 and n19600_not n19603 ; n19604
g19541 and n7294 n13736_not ; n19605
g19542 and n19604 n19605_not ; n19606
g19543 and a[11] n19606_not ; n19607
g19544 nor n19606 n19607 ; n19608
g19545 and a[11] n19607_not ; n19609
g19546 nor n19608 n19609 ; n19610
g19547 nor n19443 n19447 ; n19611
g19548 nor n19446 n19447 ; n19612
g19549 nor n19611 n19612 ; n19613
g19550 nor n19610 n19613 ; n19614
g19551 nor n19610 n19614 ; n19615
g19552 nor n19613 n19614 ; n19616
g19553 nor n19615 n19616 ; n19617
g19554 and n7983 n12370 ; n19618
g19555 and n7291 n12508 ; n19619
g19556 and n7632 n12505 ; n19620
g19557 nor n19619 n19620 ; n19621
g19558 and n19618_not n19621 ; n19622
g19559 and n7294 n13748_not ; n19623
g19560 and n19622 n19623_not ; n19624
g19561 and a[11] n19624_not ; n19625
g19562 nor n19624 n19625 ; n19626
g19563 and a[11] n19625_not ; n19627
g19564 nor n19626 n19627 ; n19628
g19565 nor n19438 n19442 ; n19629
g19566 nor n19441 n19442 ; n19630
g19567 nor n19629 n19630 ; n19631
g19568 nor n19628 n19631 ; n19632
g19569 nor n19628 n19632 ; n19633
g19570 nor n19631 n19632 ; n19634
g19571 nor n19633 n19634 ; n19635
g19572 and n7983 n12505 ; n19636
g19573 and n7291 n12513 ; n19637
g19574 and n7632 n12508 ; n19638
g19575 nor n19637 n19638 ; n19639
g19576 and n19636_not n19639 ; n19640
g19577 and n7294 n14051_not ; n19641
g19578 and n19640 n19641_not ; n19642
g19579 and a[11] n19642_not ; n19643
g19580 nor n19642 n19643 ; n19644
g19581 and a[11] n19643_not ; n19645
g19582 nor n19644 n19645 ; n19646
g19583 nor n19433 n19437 ; n19647
g19584 nor n19436 n19437 ; n19648
g19585 nor n19647 n19648 ; n19649
g19586 nor n19646 n19649 ; n19650
g19587 nor n19646 n19650 ; n19651
g19588 nor n19649 n19650 ; n19652
g19589 nor n19651 n19652 ; n19653
g19590 and n7983 n12508 ; n19654
g19591 and n7291 n12511 ; n19655
g19592 and n7632 n12513 ; n19656
g19593 nor n19655 n19656 ; n19657
g19594 and n19654_not n19657 ; n19658
g19595 and n7294 n13863 ; n19659
g19596 and n19658 n19659_not ; n19660
g19597 and a[11] n19660_not ; n19661
g19598 nor n19660 n19661 ; n19662
g19599 and a[11] n19661_not ; n19663
g19600 nor n19662 n19663 ; n19664
g19601 nor n19428 n19432 ; n19665
g19602 nor n19431 n19432 ; n19666
g19603 nor n19665 n19666 ; n19667
g19604 nor n19664 n19667 ; n19668
g19605 nor n19664 n19668 ; n19669
g19606 nor n19667 n19668 ; n19670
g19607 nor n19669 n19670 ; n19671
g19608 and n7983 n12513 ; n19672
g19609 and n7291 n12516 ; n19673
g19610 and n7632 n12511 ; n19674
g19611 nor n19673 n19674 ; n19675
g19612 and n19672_not n19675 ; n19676
g19613 and n7294 n14177 ; n19677
g19614 and n19676 n19677_not ; n19678
g19615 and a[11] n19678_not ; n19679
g19616 nor n19678 n19679 ; n19680
g19617 and a[11] n19679_not ; n19681
g19618 nor n19680 n19681 ; n19682
g19619 nor n19423 n19427 ; n19683
g19620 nor n19426 n19427 ; n19684
g19621 nor n19683 n19684 ; n19685
g19622 nor n19682 n19685 ; n19686
g19623 nor n19682 n19686 ; n19687
g19624 nor n19685 n19686 ; n19688
g19625 nor n19687 n19688 ; n19689
g19626 and n7983 n12511 ; n19690
g19627 and n7291 n12519 ; n19691
g19628 and n7632 n12516 ; n19692
g19629 nor n19691 n19692 ; n19693
g19630 and n19690_not n19693 ; n19694
g19631 and n7294 n14233_not ; n19695
g19632 and n19694 n19695_not ; n19696
g19633 and a[11] n19696_not ; n19697
g19634 nor n19696 n19697 ; n19698
g19635 and a[11] n19697_not ; n19699
g19636 nor n19698 n19699 ; n19700
g19637 nor n19418 n19422 ; n19701
g19638 nor n19421 n19422 ; n19702
g19639 nor n19701 n19702 ; n19703
g19640 nor n19700 n19703 ; n19704
g19641 nor n19700 n19704 ; n19705
g19642 nor n19703 n19704 ; n19706
g19643 nor n19705 n19706 ; n19707
g19644 and n19109 n19416 ; n19708
g19645 nor n19417 n19708 ; n19709
g19646 and n7983 n12516 ; n19710
g19647 and n7291 n12522 ; n19711
g19648 and n7632 n12519 ; n19712
g19649 nor n19711 n19712 ; n19713
g19650 and n19710_not n19713 ; n19714
g19651 and n7294_not n19714 ; n19715
g19652 and n14443 n19714 ; n19716
g19653 nor n19715 n19716 ; n19717
g19654 and a[11] n19717_not ; n19718
g19655 and a[11]_not n19717 ; n19719
g19656 nor n19718 n19719 ; n19720
g19657 and n19709 n19720_not ; n19721
g19658 and n19127 n19414 ; n19722
g19659 nor n19415 n19722 ; n19723
g19660 and n7983 n12519 ; n19724
g19661 and n7291 n12525 ; n19725
g19662 and n7632 n12522 ; n19726
g19663 nor n19725 n19726 ; n19727
g19664 and n19724_not n19727 ; n19728
g19665 and n7294_not n19728 ; n19729
g19666 and n14454_not n19728 ; n19730
g19667 nor n19729 n19730 ; n19731
g19668 and a[11] n19731_not ; n19732
g19669 and a[11]_not n19731 ; n19733
g19670 nor n19732 n19733 ; n19734
g19671 and n19723 n19734_not ; n19735
g19672 and n7983 n12522 ; n19736
g19673 and n7291 n12528 ; n19737
g19674 and n7632 n12525 ; n19738
g19675 nor n19737 n19738 ; n19739
g19676 and n19736_not n19739 ; n19740
g19677 and n7294 n14837 ; n19741
g19678 and n19740 n19741_not ; n19742
g19679 and a[11] n19742_not ; n19743
g19680 nor n19742 n19743 ; n19744
g19681 and a[11] n19743_not ; n19745
g19682 nor n19744 n19745 ; n19746
g19683 and n19410 n19412_not ; n19747
g19684 nor n19413 n19747 ; n19748
g19685 and n19746_not n19748 ; n19749
g19686 nor n19746 n19749 ; n19750
g19687 and n19748 n19749_not ; n19751
g19688 nor n19750 n19751 ; n19752
g19689 and n7983 n12525 ; n19753
g19690 and n7291 n12531 ; n19754
g19691 and n7632 n12528 ; n19755
g19692 nor n19754 n19755 ; n19756
g19693 and n19753_not n19756 ; n19757
g19694 and n7294 n14608 ; n19758
g19695 and n19757 n19758_not ; n19759
g19696 and a[11] n19759_not ; n19760
g19697 nor n19759 n19760 ; n19761
g19698 and a[11] n19760_not ; n19762
g19699 nor n19761 n19762 ; n19763
g19700 nor n19405 n19409 ; n19764
g19701 nor n19408 n19409 ; n19765
g19702 nor n19764 n19765 ; n19766
g19703 nor n19763 n19766 ; n19767
g19704 nor n19763 n19767 ; n19768
g19705 nor n19766 n19767 ; n19769
g19706 nor n19768 n19769 ; n19770
g19707 and n7983 n12528 ; n19771
g19708 and n7291 n12534 ; n19772
g19709 and n7632 n12531 ; n19773
g19710 nor n19772 n19773 ; n19774
g19711 and n19771_not n19774 ; n19775
g19712 and n7294 n15003_not ; n19776
g19713 and n19775 n19776_not ; n19777
g19714 and a[11] n19777_not ; n19778
g19715 nor n19777 n19778 ; n19779
g19716 and a[11] n19778_not ; n19780
g19717 nor n19779 n19780 ; n19781
g19718 nor n19400 n19404 ; n19782
g19719 nor n19403 n19404 ; n19783
g19720 nor n19782 n19783 ; n19784
g19721 nor n19781 n19784 ; n19785
g19722 nor n19781 n19785 ; n19786
g19723 nor n19784 n19785 ; n19787
g19724 nor n19786 n19787 ; n19788
g19725 and n19186 n19398 ; n19789
g19726 nor n19399 n19789 ; n19790
g19727 and n7983 n12531 ; n19791
g19728 and n7291 n12537 ; n19792
g19729 and n7632 n12534 ; n19793
g19730 nor n19792 n19793 ; n19794
g19731 and n19791_not n19794 ; n19795
g19732 and n7294_not n19795 ; n19796
g19733 and n15255_not n19795 ; n19797
g19734 nor n19796 n19797 ; n19798
g19735 and a[11] n19798_not ; n19799
g19736 and a[11]_not n19798 ; n19800
g19737 nor n19799 n19800 ; n19801
g19738 and n19790 n19801_not ; n19802
g19739 and n19204 n19396 ; n19803
g19740 nor n19397 n19803 ; n19804
g19741 and n7983 n12534 ; n19805
g19742 and n7291 n12540 ; n19806
g19743 and n7632 n12537 ; n19807
g19744 nor n19806 n19807 ; n19808
g19745 and n19805_not n19808 ; n19809
g19746 and n7294_not n19809 ; n19810
g19747 and n15096 n19809 ; n19811
g19748 nor n19810 n19811 ; n19812
g19749 and a[11] n19812_not ; n19813
g19750 and a[11]_not n19812 ; n19814
g19751 nor n19813 n19814 ; n19815
g19752 and n19804 n19815_not ; n19816
g19753 and n19222 n19394 ; n19817
g19754 nor n19395 n19817 ; n19818
g19755 and n7983 n12537 ; n19819
g19756 and n7291 n12543 ; n19820
g19757 and n7632 n12540 ; n19821
g19758 nor n19820 n19821 ; n19822
g19759 and n19819_not n19822 ; n19823
g19760 and n7294_not n19823 ; n19824
g19761 and n15385 n19823 ; n19825
g19762 nor n19824 n19825 ; n19826
g19763 and a[11] n19826_not ; n19827
g19764 and a[11]_not n19826 ; n19828
g19765 nor n19827 n19828 ; n19829
g19766 and n19818 n19829_not ; n19830
g19767 and n7983 n12540 ; n19831
g19768 and n7291 n12546 ; n19832
g19769 and n7632 n12543 ; n19833
g19770 nor n19832 n19833 ; n19834
g19771 and n19831_not n19834 ; n19835
g19772 and n7294 n15708_not ; n19836
g19773 and n19835 n19836_not ; n19837
g19774 and a[11] n19837_not ; n19838
g19775 nor n19837 n19838 ; n19839
g19776 and a[11] n19838_not ; n19840
g19777 nor n19839 n19840 ; n19841
g19778 and n19390 n19392_not ; n19842
g19779 nor n19393 n19842 ; n19843
g19780 and n19841_not n19843 ; n19844
g19781 nor n19841 n19844 ; n19845
g19782 and n19843 n19844_not ; n19846
g19783 nor n19845 n19846 ; n19847
g19784 and n7983 n12543 ; n19848
g19785 and n7291 n12549 ; n19849
g19786 and n7632 n12546 ; n19850
g19787 nor n19849 n19850 ; n19851
g19788 and n19848_not n19851 ; n19852
g19789 and n7294 n15724 ; n19853
g19790 and n19852 n19853_not ; n19854
g19791 and a[11] n19854_not ; n19855
g19792 nor n19854 n19855 ; n19856
g19793 and a[11] n19855_not ; n19857
g19794 nor n19856 n19857 ; n19858
g19795 nor n19385 n19389 ; n19859
g19796 nor n19388 n19389 ; n19860
g19797 nor n19859 n19860 ; n19861
g19798 nor n19858 n19861 ; n19862
g19799 nor n19858 n19862 ; n19863
g19800 nor n19861 n19862 ; n19864
g19801 nor n19863 n19864 ; n19865
g19802 and n7983 n12546 ; n19866
g19803 and n7291 n12552 ; n19867
g19804 and n7632 n12549 ; n19868
g19805 nor n19867 n19868 ; n19869
g19806 and n19866_not n19869 ; n19870
g19807 and n7294 n15356_not ; n19871
g19808 and n19870 n19871_not ; n19872
g19809 and a[11] n19872_not ; n19873
g19810 nor n19872 n19873 ; n19874
g19811 and a[11] n19873_not ; n19875
g19812 nor n19874 n19875 ; n19876
g19813 nor n19380 n19384 ; n19877
g19814 nor n19383 n19384 ; n19878
g19815 nor n19877 n19878 ; n19879
g19816 nor n19876 n19879 ; n19880
g19817 nor n19876 n19880 ; n19881
g19818 nor n19879 n19880 ; n19882
g19819 nor n19881 n19882 ; n19883
g19820 and n19281 n19378 ; n19884
g19821 nor n19379 n19884 ; n19885
g19822 and n7983 n12549 ; n19886
g19823 and n7291 n12555 ; n19887
g19824 and n7632 n12552 ; n19888
g19825 nor n19887 n19888 ; n19889
g19826 and n19886_not n19889 ; n19890
g19827 and n7294_not n19890 ; n19891
g19828 and n15764_not n19890 ; n19892
g19829 nor n19891 n19892 ; n19893
g19830 and a[11] n19893_not ; n19894
g19831 and a[11]_not n19893 ; n19895
g19832 nor n19894 n19895 ; n19896
g19833 and n19885 n19896_not ; n19897
g19834 and n19374 n19376_not ; n19898
g19835 nor n19377 n19898 ; n19899
g19836 and n7983 n12552 ; n19900
g19837 and n7291 n12558 ; n19901
g19838 and n7632 n12555 ; n19902
g19839 nor n19901 n19902 ; n19903
g19840 and n19900_not n19903 ; n19904
g19841 and n7294_not n19904 ; n19905
g19842 and n15791 n19904 ; n19906
g19843 nor n19905 n19906 ; n19907
g19844 and a[11] n19907_not ; n19908
g19845 and a[11]_not n19907 ; n19909
g19846 nor n19908 n19909 ; n19910
g19847 and n19899 n19910_not ; n19911
g19848 and n19313 n19372 ; n19912
g19849 nor n19373 n19912 ; n19913
g19850 and n7983 n12555 ; n19914
g19851 and n7291 n12561 ; n19915
g19852 and n7632 n12558 ; n19916
g19853 nor n19915 n19916 ; n19917
g19854 and n19914_not n19917 ; n19918
g19855 and n7294_not n19918 ; n19919
g19856 and n15816 n19918 ; n19920
g19857 nor n19919 n19920 ; n19921
g19858 and a[11] n19921_not ; n19922
g19859 and a[11]_not n19921 ; n19923
g19860 nor n19922 n19923 ; n19924
g19861 and n19913 n19924_not ; n19925
g19862 and n7983 n12558 ; n19926
g19863 and n7291 n12564 ; n19927
g19864 and n7632 n12561 ; n19928
g19865 nor n19927 n19928 ; n19929
g19866 and n19926_not n19929 ; n19930
g19867 and n7294 n15847 ; n19931
g19868 and n19930 n19931_not ; n19932
g19869 and a[11] n19932_not ; n19933
g19870 nor n19932 n19933 ; n19934
g19871 and a[11] n19933_not ; n19935
g19872 nor n19934 n19935 ; n19936
g19873 and n19368 n19370_not ; n19937
g19874 nor n19371 n19937 ; n19938
g19875 and n19936_not n19938 ; n19939
g19876 nor n19936 n19939 ; n19940
g19877 and n19938 n19939_not ; n19941
g19878 nor n19940 n19941 ; n19942
g19879 nor n19355 n19367 ; n19943
g19880 nor n19366 n19367 ; n19944
g19881 nor n19943 n19944 ; n19945
g19882 and n7983 n12561 ; n19946
g19883 and n7291 n12567 ; n19947
g19884 and n7632 n12564 ; n19948
g19885 nor n19947 n19948 ; n19949
g19886 and n19946_not n19949 ; n19950
g19887 and n7294_not n19950 ; n19951
g19888 and n15905 n19950 ; n19952
g19889 nor n19951 n19952 ; n19953
g19890 and a[11] n19953_not ; n19954
g19891 and a[11]_not n19953 ; n19955
g19892 nor n19954 n19955 ; n19956
g19893 nor n19945 n19956 ; n19957
g19894 and n7983 n12564 ; n19958
g19895 and n7291 n12571 ; n19959
g19896 and n7632 n12567 ; n19960
g19897 nor n19959 n19960 ; n19961
g19898 and n19958_not n19961 ; n19962
g19899 and n7294 n15944_not ; n19963
g19900 and n19962 n19963_not ; n19964
g19901 and a[11] n19964_not ; n19965
g19902 nor n19964 n19965 ; n19966
g19903 and a[11] n19965_not ; n19967
g19904 nor n19966 n19967 ; n19968
g19905 and n19339_not n19350 ; n19969
g19906 nor n19351 n19969 ; n19970
g19907 and n19968_not n19970 ; n19971
g19908 nor n19968 n19971 ; n19972
g19909 and n19970 n19971_not ; n19973
g19910 nor n19972 n19973 ; n19974
g19911 and n19336 n19338_not ; n19975
g19912 nor n19339 n19975 ; n19976
g19913 and n7983 n12567 ; n19977
g19914 and n7291 n12574 ; n19978
g19915 and n7632 n12571 ; n19979
g19916 nor n19978 n19979 ; n19980
g19917 and n19977_not n19980 ; n19981
g19918 and n7294_not n19981 ; n19982
g19919 and n15989_not n19981 ; n19983
g19920 nor n19982 n19983 ; n19984
g19921 and a[11] n19984_not ; n19985
g19922 and a[11]_not n19984 ; n19986
g19923 nor n19985 n19986 ; n19987
g19924 and n19976 n19987_not ; n19988
g19925 and n7632 n12581_not ; n19989
g19926 and n7983 n12577 ; n19990
g19927 nor n19989 n19990 ; n19991
g19928 and n7294 n16085_not ; n19992
g19929 and n19991 n19992_not ; n19993
g19930 and a[11] n19993_not ; n19994
g19931 and a[11] n19994_not ; n19995
g19932 nor n19993 n19994 ; n19996
g19933 nor n19995 n19996 ; n19997
g19934 nor n7289 n12581 ; n19998
g19935 and a[11] n19998_not ; n19999
g19936 and n19997_not n19999 ; n20000
g19937 and n7983 n12574 ; n20001
g19938 and n7291 n12581_not ; n20002
g19939 and n7632 n12577 ; n20003
g19940 nor n20002 n20003 ; n20004
g19941 and n20001_not n20004 ; n20005
g19942 and n7294_not n20005 ; n20006
g19943 and n16094 n20005 ; n20007
g19944 nor n20006 n20007 ; n20008
g19945 and a[11] n20008_not ; n20009
g19946 and a[11]_not n20008 ; n20010
g19947 nor n20009 n20010 ; n20011
g19948 and n20000 n20011_not ; n20012
g19949 and n19337 n20012 ; n20013
g19950 and n20012 n20013_not ; n20014
g19951 and n19337 n20013_not ; n20015
g19952 nor n20014 n20015 ; n20016
g19953 and n7983 n12571 ; n20017
g19954 and n7291 n12577 ; n20018
g19955 and n7632 n12574 ; n20019
g19956 nor n20018 n20019 ; n20020
g19957 and n20017_not n20020 ; n20021
g19958 and n7294 n16013 ; n20022
g19959 and n20021 n20022_not ; n20023
g19960 and a[11] n20023_not ; n20024
g19961 and a[11] n20024_not ; n20025
g19962 nor n20023 n20024 ; n20026
g19963 nor n20025 n20026 ; n20027
g19964 nor n20016 n20027 ; n20028
g19965 nor n20013 n20028 ; n20029
g19966 and n19976_not n19987 ; n20030
g19967 nor n19988 n20030 ; n20031
g19968 and n20029_not n20031 ; n20032
g19969 nor n19988 n20032 ; n20033
g19970 nor n19974 n20033 ; n20034
g19971 nor n19971 n20034 ; n20035
g19972 and n19945 n19956 ; n20036
g19973 nor n19957 n20036 ; n20037
g19974 and n20035_not n20037 ; n20038
g19975 nor n19957 n20038 ; n20039
g19976 nor n19942 n20039 ; n20040
g19977 nor n19939 n20040 ; n20041
g19978 and n19913 n19925_not ; n20042
g19979 nor n19924 n19925 ; n20043
g19980 nor n20042 n20043 ; n20044
g19981 nor n20041 n20044 ; n20045
g19982 nor n19925 n20045 ; n20046
g19983 and n19899 n19911_not ; n20047
g19984 nor n19910 n19911 ; n20048
g19985 nor n20047 n20048 ; n20049
g19986 nor n20046 n20049 ; n20050
g19987 nor n19911 n20050 ; n20051
g19988 and n19885_not n19896 ; n20052
g19989 nor n19897 n20052 ; n20053
g19990 and n20051_not n20053 ; n20054
g19991 nor n19897 n20054 ; n20055
g19992 nor n19883 n20055 ; n20056
g19993 nor n19880 n20056 ; n20057
g19994 nor n19865 n20057 ; n20058
g19995 nor n19862 n20058 ; n20059
g19996 nor n19847 n20059 ; n20060
g19997 nor n19844 n20060 ; n20061
g19998 and n19818 n19830_not ; n20062
g19999 nor n19829 n19830 ; n20063
g20000 nor n20062 n20063 ; n20064
g20001 nor n20061 n20064 ; n20065
g20002 nor n19830 n20065 ; n20066
g20003 and n19804 n19816_not ; n20067
g20004 nor n19815 n19816 ; n20068
g20005 nor n20067 n20068 ; n20069
g20006 nor n20066 n20069 ; n20070
g20007 nor n19816 n20070 ; n20071
g20008 and n19790_not n19801 ; n20072
g20009 nor n19802 n20072 ; n20073
g20010 and n20071_not n20073 ; n20074
g20011 nor n19802 n20074 ; n20075
g20012 nor n19788 n20075 ; n20076
g20013 nor n19785 n20076 ; n20077
g20014 nor n19770 n20077 ; n20078
g20015 nor n19767 n20078 ; n20079
g20016 nor n19752 n20079 ; n20080
g20017 nor n19749 n20080 ; n20081
g20018 and n19723 n19735_not ; n20082
g20019 nor n19734 n19735 ; n20083
g20020 nor n20082 n20083 ; n20084
g20021 nor n20081 n20084 ; n20085
g20022 nor n19735 n20085 ; n20086
g20023 and n19709_not n19720 ; n20087
g20024 nor n19721 n20087 ; n20088
g20025 and n20086_not n20088 ; n20089
g20026 nor n19721 n20089 ; n20090
g20027 nor n19707 n20090 ; n20091
g20028 nor n19704 n20091 ; n20092
g20029 nor n19689 n20092 ; n20093
g20030 nor n19686 n20093 ; n20094
g20031 nor n19671 n20094 ; n20095
g20032 nor n19668 n20095 ; n20096
g20033 nor n19653 n20096 ; n20097
g20034 nor n19650 n20097 ; n20098
g20035 nor n19635 n20098 ; n20099
g20036 nor n19632 n20099 ; n20100
g20037 nor n19617 n20100 ; n20101
g20038 nor n19614 n20101 ; n20102
g20039 nor n19599 n20102 ; n20103
g20040 nor n19596 n20103 ; n20104
g20041 nor n19581 n20104 ; n20105
g20042 nor n19578 n20105 ; n20106
g20043 nor n19563 n20106 ; n20107
g20044 nor n19560 n20107 ; n20108
g20045 nor n19545 n20108 ; n20109
g20046 nor n19542 n20109 ; n20110
g20047 nor n19528 n20110 ; n20111
g20048 and n19528 n20110 ; n20112
g20049 nor n20111 n20112 ; n20113
g20050 and n9331 n13630 ; n20114
g20051 and n8418 n13515 ; n20115
g20052 and n8860 n13597 ; n20116
g20053 nor n20115 n20116 ; n20117
g20054 and n20114_not n20117 ; n20118
g20055 and n8421 n13976 ; n20119
g20056 and n20118 n20119_not ; n20120
g20057 and a[8] n20120_not ; n20121
g20058 and a[8] n20121_not ; n20122
g20059 nor n20120 n20121 ; n20123
g20060 nor n20122 n20123 ; n20124
g20061 and n20113 n20124_not ; n20125
g20062 nor n20111 n20125 ; n20126
g20063 nor n19525 n20126 ; n20127
g20064 and n19525 n20126 ; n20128
g20065 nor n20127 n20128 ; n20129
g20066 and n71 n13438_not ; n20130
g20067 and n9867 n13627_not ; n20131
g20068 and n10434 n13941 ; n20132
g20069 nor n20131 n20132 ; n20133
g20070 and n20130_not n20133 ; n20134
g20071 and n9870 n14028 ; n20135
g20072 and n20134 n20135_not ; n20136
g20073 and a[5] n20136_not ; n20137
g20074 and a[5] n20137_not ; n20138
g20075 nor n20136 n20137 ; n20139
g20076 nor n20138 n20139 ; n20140
g20077 and n20129 n20140_not ; n20141
g20078 nor n20127 n20141 ; n20142
g20079 nor n19522 n20142 ; n20143
g20080 and n19522 n20142 ; n20144
g20081 nor n20143 n20144 ; n20145
g20082 and n20129 n20141_not ; n20146
g20083 nor n20140 n20141 ; n20147
g20084 nor n20146 n20147 ; n20148
g20085 and n20113 n20125_not ; n20149
g20086 nor n20124 n20125 ; n20150
g20087 nor n20149 n20150 ; n20151
g20088 and n19545 n20108 ; n20152
g20089 nor n20109 n20152 ; n20153
g20090 and n9331 n13597 ; n20154
g20091 and n8418 n13521 ; n20155
g20092 and n8860 n13515 ; n20156
g20093 nor n20155 n20156 ; n20157
g20094 and n20154_not n20157 ; n20158
g20095 and n8421_not n20158 ; n20159
g20096 and n13612 n20158 ; n20160
g20097 nor n20159 n20160 ; n20161
g20098 and a[8] n20161_not ; n20162
g20099 and a[8]_not n20161 ; n20163
g20100 nor n20162 n20163 ; n20164
g20101 and n20153 n20164_not ; n20165
g20102 and n19563 n20106 ; n20166
g20103 nor n20107 n20166 ; n20167
g20104 and n9331 n13515 ; n20168
g20105 and n8418 n13518 ; n20169
g20106 and n8860 n13521 ; n20170
g20107 nor n20169 n20170 ; n20171
g20108 and n20168_not n20171 ; n20172
g20109 and n8421_not n20172 ; n20173
g20110 and n13541_not n20172 ; n20174
g20111 nor n20173 n20174 ; n20175
g20112 and a[8] n20175_not ; n20176
g20113 and a[8]_not n20175 ; n20177
g20114 nor n20176 n20177 ; n20178
g20115 and n20167 n20178_not ; n20179
g20116 and n19581 n20104 ; n20180
g20117 nor n20105 n20180 ; n20181
g20118 and n9331 n13521 ; n20182
g20119 and n8418 n13491 ; n20183
g20120 and n8860 n13518 ; n20184
g20121 nor n20183 n20184 ; n20185
g20122 and n20182_not n20185 ; n20186
g20123 and n8421_not n20186 ; n20187
g20124 and n13909 n20186 ; n20188
g20125 nor n20187 n20188 ; n20189
g20126 and a[8] n20189_not ; n20190
g20127 and a[8]_not n20189 ; n20191
g20128 nor n20190 n20191 ; n20192
g20129 and n20181 n20192_not ; n20193
g20130 and n19599 n20102 ; n20194
g20131 nor n20103 n20194 ; n20195
g20132 and n9331 n13518 ; n20196
g20133 and n8418 n12889 ; n20197
g20134 and n8860 n13491 ; n20198
g20135 nor n20197 n20198 ; n20199
g20136 and n20196_not n20199 ; n20200
g20137 and n8421_not n20200 ; n20201
g20138 and n13584_not n20200 ; n20202
g20139 nor n20201 n20202 ; n20203
g20140 and a[8] n20203_not ; n20204
g20141 and a[8]_not n20203 ; n20205
g20142 nor n20204 n20205 ; n20206
g20143 and n20195 n20206_not ; n20207
g20144 and n19617 n20100 ; n20208
g20145 nor n20101 n20208 ; n20209
g20146 and n9331 n13491 ; n20210
g20147 and n8418 n12769 ; n20211
g20148 and n8860 n12889 ; n20212
g20149 nor n20211 n20212 ; n20213
g20150 and n20210_not n20213 ; n20214
g20151 and n8421_not n20214 ; n20215
g20152 and n13503 n20214 ; n20216
g20153 nor n20215 n20216 ; n20217
g20154 and a[8] n20217_not ; n20218
g20155 and a[8]_not n20217 ; n20219
g20156 nor n20218 n20219 ; n20220
g20157 and n20209 n20220_not ; n20221
g20158 and n19635 n20098 ; n20222
g20159 nor n20099 n20222 ; n20223
g20160 and n9331 n12889 ; n20224
g20161 and n8418 n12502 ; n20225
g20162 and n8860 n12769 ; n20226
g20163 nor n20225 n20226 ; n20227
g20164 and n20224_not n20227 ; n20228
g20165 and n8421_not n20228 ; n20229
g20166 and n12895_not n20228 ; n20230
g20167 nor n20229 n20230 ; n20231
g20168 and a[8] n20231_not ; n20232
g20169 and a[8]_not n20231 ; n20233
g20170 nor n20232 n20233 ; n20234
g20171 and n20223 n20234_not ; n20235
g20172 and n19653 n20096 ; n20236
g20173 nor n20097 n20236 ; n20237
g20174 and n9331 n12769 ; n20238
g20175 and n8418 n12370 ; n20239
g20176 and n8860 n12502 ; n20240
g20177 nor n20239 n20240 ; n20241
g20178 and n20238_not n20241 ; n20242
g20179 and n8421_not n20242 ; n20243
g20180 and n12999_not n20242 ; n20244
g20181 nor n20243 n20244 ; n20245
g20182 and a[8] n20245_not ; n20246
g20183 and a[8]_not n20245 ; n20247
g20184 nor n20246 n20247 ; n20248
g20185 and n20237 n20248_not ; n20249
g20186 and n19671 n20094 ; n20250
g20187 nor n20095 n20250 ; n20251
g20188 and n9331 n12502 ; n20252
g20189 and n8418 n12505 ; n20253
g20190 and n8860 n12370 ; n20254
g20191 nor n20253 n20254 ; n20255
g20192 and n20252_not n20255 ; n20256
g20193 and n8421_not n20256 ; n20257
g20194 and n13736 n20256 ; n20258
g20195 nor n20257 n20258 ; n20259
g20196 and a[8] n20259_not ; n20260
g20197 and a[8]_not n20259 ; n20261
g20198 nor n20260 n20261 ; n20262
g20199 and n20251 n20262_not ; n20263
g20200 and n19689 n20092 ; n20264
g20201 nor n20093 n20264 ; n20265
g20202 and n9331 n12370 ; n20266
g20203 and n8418 n12508 ; n20267
g20204 and n8860 n12505 ; n20268
g20205 nor n20267 n20268 ; n20269
g20206 and n20266_not n20269 ; n20270
g20207 and n8421_not n20270 ; n20271
g20208 and n13748 n20270 ; n20272
g20209 nor n20271 n20272 ; n20273
g20210 and a[8] n20273_not ; n20274
g20211 and a[8]_not n20273 ; n20275
g20212 nor n20274 n20275 ; n20276
g20213 and n20265 n20276_not ; n20277
g20214 and n19707 n20090 ; n20278
g20215 nor n20091 n20278 ; n20279
g20216 and n9331 n12505 ; n20280
g20217 and n8418 n12513 ; n20281
g20218 and n8860 n12508 ; n20282
g20219 nor n20281 n20282 ; n20283
g20220 and n20280_not n20283 ; n20284
g20221 and n8421_not n20284 ; n20285
g20222 and n14051 n20284 ; n20286
g20223 nor n20285 n20286 ; n20287
g20224 and a[8] n20287_not ; n20288
g20225 and a[8]_not n20287 ; n20289
g20226 nor n20288 n20289 ; n20290
g20227 and n20279 n20290_not ; n20291
g20228 and n9331 n12508 ; n20292
g20229 and n8418 n12511 ; n20293
g20230 and n8860 n12513 ; n20294
g20231 nor n20293 n20294 ; n20295
g20232 and n20292_not n20295 ; n20296
g20233 and n8421 n13863 ; n20297
g20234 and n20296 n20297_not ; n20298
g20235 and a[8] n20298_not ; n20299
g20236 nor n20298 n20299 ; n20300
g20237 and a[8] n20299_not ; n20301
g20238 nor n20300 n20301 ; n20302
g20239 and n20086 n20088_not ; n20303
g20240 nor n20089 n20303 ; n20304
g20241 and n20302_not n20304 ; n20305
g20242 nor n20302 n20305 ; n20306
g20243 and n20304 n20305_not ; n20307
g20244 nor n20306 n20307 ; n20308
g20245 and n9331 n12513 ; n20309
g20246 and n8418 n12516 ; n20310
g20247 and n8860 n12511 ; n20311
g20248 nor n20310 n20311 ; n20312
g20249 and n20309_not n20312 ; n20313
g20250 and n8421 n14177 ; n20314
g20251 and n20313 n20314_not ; n20315
g20252 and a[8] n20315_not ; n20316
g20253 nor n20315 n20316 ; n20317
g20254 and a[8] n20316_not ; n20318
g20255 nor n20317 n20318 ; n20319
g20256 nor n20081 n20085 ; n20320
g20257 nor n20084 n20085 ; n20321
g20258 nor n20320 n20321 ; n20322
g20259 nor n20319 n20322 ; n20323
g20260 nor n20319 n20323 ; n20324
g20261 nor n20322 n20323 ; n20325
g20262 nor n20324 n20325 ; n20326
g20263 and n19752 n20079 ; n20327
g20264 nor n20080 n20327 ; n20328
g20265 and n9331 n12511 ; n20329
g20266 and n8418 n12519 ; n20330
g20267 and n8860 n12516 ; n20331
g20268 nor n20330 n20331 ; n20332
g20269 and n20329_not n20332 ; n20333
g20270 and n8421_not n20333 ; n20334
g20271 and n14233 n20333 ; n20335
g20272 nor n20334 n20335 ; n20336
g20273 and a[8] n20336_not ; n20337
g20274 and a[8]_not n20336 ; n20338
g20275 nor n20337 n20338 ; n20339
g20276 and n20328 n20339_not ; n20340
g20277 and n19770 n20077 ; n20341
g20278 nor n20078 n20341 ; n20342
g20279 and n9331 n12516 ; n20343
g20280 and n8418 n12522 ; n20344
g20281 and n8860 n12519 ; n20345
g20282 nor n20344 n20345 ; n20346
g20283 and n20343_not n20346 ; n20347
g20284 and n8421_not n20347 ; n20348
g20285 and n14443 n20347 ; n20349
g20286 nor n20348 n20349 ; n20350
g20287 and a[8] n20350_not ; n20351
g20288 and a[8]_not n20350 ; n20352
g20289 nor n20351 n20352 ; n20353
g20290 and n20342 n20353_not ; n20354
g20291 and n19788 n20075 ; n20355
g20292 nor n20076 n20355 ; n20356
g20293 and n9331 n12519 ; n20357
g20294 and n8418 n12525 ; n20358
g20295 and n8860 n12522 ; n20359
g20296 nor n20358 n20359 ; n20360
g20297 and n20357_not n20360 ; n20361
g20298 and n8421_not n20361 ; n20362
g20299 and n14454_not n20361 ; n20363
g20300 nor n20362 n20363 ; n20364
g20301 and a[8] n20364_not ; n20365
g20302 and a[8]_not n20364 ; n20366
g20303 nor n20365 n20366 ; n20367
g20304 and n20356 n20367_not ; n20368
g20305 and n9331 n12522 ; n20369
g20306 and n8418 n12528 ; n20370
g20307 and n8860 n12525 ; n20371
g20308 nor n20370 n20371 ; n20372
g20309 and n20369_not n20372 ; n20373
g20310 and n8421 n14837 ; n20374
g20311 and n20373 n20374_not ; n20375
g20312 and a[8] n20375_not ; n20376
g20313 nor n20375 n20376 ; n20377
g20314 and a[8] n20376_not ; n20378
g20315 nor n20377 n20378 ; n20379
g20316 and n20071 n20073_not ; n20380
g20317 nor n20074 n20380 ; n20381
g20318 and n20379_not n20381 ; n20382
g20319 nor n20379 n20382 ; n20383
g20320 and n20381 n20382_not ; n20384
g20321 nor n20383 n20384 ; n20385
g20322 and n9331 n12525 ; n20386
g20323 and n8418 n12531 ; n20387
g20324 and n8860 n12528 ; n20388
g20325 nor n20387 n20388 ; n20389
g20326 and n20386_not n20389 ; n20390
g20327 and n8421 n14608 ; n20391
g20328 and n20390 n20391_not ; n20392
g20329 and a[8] n20392_not ; n20393
g20330 nor n20392 n20393 ; n20394
g20331 and a[8] n20393_not ; n20395
g20332 nor n20394 n20395 ; n20396
g20333 nor n20066 n20070 ; n20397
g20334 nor n20069 n20070 ; n20398
g20335 nor n20397 n20398 ; n20399
g20336 nor n20396 n20399 ; n20400
g20337 nor n20396 n20400 ; n20401
g20338 nor n20399 n20400 ; n20402
g20339 nor n20401 n20402 ; n20403
g20340 and n9331 n12528 ; n20404
g20341 and n8418 n12534 ; n20405
g20342 and n8860 n12531 ; n20406
g20343 nor n20405 n20406 ; n20407
g20344 and n20404_not n20407 ; n20408
g20345 and n8421 n15003_not ; n20409
g20346 and n20408 n20409_not ; n20410
g20347 and a[8] n20410_not ; n20411
g20348 nor n20410 n20411 ; n20412
g20349 and a[8] n20411_not ; n20413
g20350 nor n20412 n20413 ; n20414
g20351 nor n20061 n20065 ; n20415
g20352 nor n20064 n20065 ; n20416
g20353 nor n20415 n20416 ; n20417
g20354 nor n20414 n20417 ; n20418
g20355 nor n20414 n20418 ; n20419
g20356 nor n20417 n20418 ; n20420
g20357 nor n20419 n20420 ; n20421
g20358 and n19847 n20059 ; n20422
g20359 nor n20060 n20422 ; n20423
g20360 and n9331 n12531 ; n20424
g20361 and n8418 n12537 ; n20425
g20362 and n8860 n12534 ; n20426
g20363 nor n20425 n20426 ; n20427
g20364 and n20424_not n20427 ; n20428
g20365 and n8421_not n20428 ; n20429
g20366 and n15255_not n20428 ; n20430
g20367 nor n20429 n20430 ; n20431
g20368 and a[8] n20431_not ; n20432
g20369 and a[8]_not n20431 ; n20433
g20370 nor n20432 n20433 ; n20434
g20371 and n20423 n20434_not ; n20435
g20372 and n19865 n20057 ; n20436
g20373 nor n20058 n20436 ; n20437
g20374 and n9331 n12534 ; n20438
g20375 and n8418 n12540 ; n20439
g20376 and n8860 n12537 ; n20440
g20377 nor n20439 n20440 ; n20441
g20378 and n20438_not n20441 ; n20442
g20379 and n8421_not n20442 ; n20443
g20380 and n15096 n20442 ; n20444
g20381 nor n20443 n20444 ; n20445
g20382 and a[8] n20445_not ; n20446
g20383 and a[8]_not n20445 ; n20447
g20384 nor n20446 n20447 ; n20448
g20385 and n20437 n20448_not ; n20449
g20386 and n19883 n20055 ; n20450
g20387 nor n20056 n20450 ; n20451
g20388 and n9331 n12537 ; n20452
g20389 and n8418 n12543 ; n20453
g20390 and n8860 n12540 ; n20454
g20391 nor n20453 n20454 ; n20455
g20392 and n20452_not n20455 ; n20456
g20393 and n8421_not n20456 ; n20457
g20394 and n15385 n20456 ; n20458
g20395 nor n20457 n20458 ; n20459
g20396 and a[8] n20459_not ; n20460
g20397 and a[8]_not n20459 ; n20461
g20398 nor n20460 n20461 ; n20462
g20399 and n20451 n20462_not ; n20463
g20400 and n9331 n12540 ; n20464
g20401 and n8418 n12546 ; n20465
g20402 and n8860 n12543 ; n20466
g20403 nor n20465 n20466 ; n20467
g20404 and n20464_not n20467 ; n20468
g20405 and n8421 n15708_not ; n20469
g20406 and n20468 n20469_not ; n20470
g20407 and a[8] n20470_not ; n20471
g20408 nor n20470 n20471 ; n20472
g20409 and a[8] n20471_not ; n20473
g20410 nor n20472 n20473 ; n20474
g20411 and n20051 n20053_not ; n20475
g20412 nor n20054 n20475 ; n20476
g20413 and n20474_not n20476 ; n20477
g20414 nor n20474 n20477 ; n20478
g20415 and n20476 n20477_not ; n20479
g20416 nor n20478 n20479 ; n20480
g20417 and n9331 n12543 ; n20481
g20418 and n8418 n12549 ; n20482
g20419 and n8860 n12546 ; n20483
g20420 nor n20482 n20483 ; n20484
g20421 and n20481_not n20484 ; n20485
g20422 and n8421 n15724 ; n20486
g20423 and n20485 n20486_not ; n20487
g20424 and a[8] n20487_not ; n20488
g20425 nor n20487 n20488 ; n20489
g20426 and a[8] n20488_not ; n20490
g20427 nor n20489 n20490 ; n20491
g20428 nor n20046 n20050 ; n20492
g20429 nor n20049 n20050 ; n20493
g20430 nor n20492 n20493 ; n20494
g20431 nor n20491 n20494 ; n20495
g20432 nor n20491 n20495 ; n20496
g20433 nor n20494 n20495 ; n20497
g20434 nor n20496 n20497 ; n20498
g20435 and n9331 n12546 ; n20499
g20436 and n8418 n12552 ; n20500
g20437 and n8860 n12549 ; n20501
g20438 nor n20500 n20501 ; n20502
g20439 and n20499_not n20502 ; n20503
g20440 and n8421 n15356_not ; n20504
g20441 and n20503 n20504_not ; n20505
g20442 and a[8] n20505_not ; n20506
g20443 nor n20505 n20506 ; n20507
g20444 and a[8] n20506_not ; n20508
g20445 nor n20507 n20508 ; n20509
g20446 nor n20041 n20045 ; n20510
g20447 nor n20044 n20045 ; n20511
g20448 nor n20510 n20511 ; n20512
g20449 nor n20509 n20512 ; n20513
g20450 nor n20509 n20513 ; n20514
g20451 nor n20512 n20513 ; n20515
g20452 nor n20514 n20515 ; n20516
g20453 and n19942 n20039 ; n20517
g20454 nor n20040 n20517 ; n20518
g20455 and n9331 n12549 ; n20519
g20456 and n8418 n12555 ; n20520
g20457 and n8860 n12552 ; n20521
g20458 nor n20520 n20521 ; n20522
g20459 and n20519_not n20522 ; n20523
g20460 and n8421_not n20523 ; n20524
g20461 and n15764_not n20523 ; n20525
g20462 nor n20524 n20525 ; n20526
g20463 and a[8] n20526_not ; n20527
g20464 and a[8]_not n20526 ; n20528
g20465 nor n20527 n20528 ; n20529
g20466 and n20518 n20529_not ; n20530
g20467 and n20035 n20037_not ; n20531
g20468 nor n20038 n20531 ; n20532
g20469 and n9331 n12552 ; n20533
g20470 and n8418 n12558 ; n20534
g20471 and n8860 n12555 ; n20535
g20472 nor n20534 n20535 ; n20536
g20473 and n20533_not n20536 ; n20537
g20474 and n8421_not n20537 ; n20538
g20475 and n15791 n20537 ; n20539
g20476 nor n20538 n20539 ; n20540
g20477 and a[8] n20540_not ; n20541
g20478 and a[8]_not n20540 ; n20542
g20479 nor n20541 n20542 ; n20543
g20480 and n20532 n20543_not ; n20544
g20481 and n19974 n20033 ; n20545
g20482 nor n20034 n20545 ; n20546
g20483 and n9331 n12555 ; n20547
g20484 and n8418 n12561 ; n20548
g20485 and n8860 n12558 ; n20549
g20486 nor n20548 n20549 ; n20550
g20487 and n20547_not n20550 ; n20551
g20488 and n8421_not n20551 ; n20552
g20489 and n15816 n20551 ; n20553
g20490 nor n20552 n20553 ; n20554
g20491 and a[8] n20554_not ; n20555
g20492 and a[8]_not n20554 ; n20556
g20493 nor n20555 n20556 ; n20557
g20494 and n20546 n20557_not ; n20558
g20495 and n9331 n12558 ; n20559
g20496 and n8418 n12564 ; n20560
g20497 and n8860 n12561 ; n20561
g20498 nor n20560 n20561 ; n20562
g20499 and n20559_not n20562 ; n20563
g20500 and n8421 n15847 ; n20564
g20501 and n20563 n20564_not ; n20565
g20502 and a[8] n20565_not ; n20566
g20503 nor n20565 n20566 ; n20567
g20504 and a[8] n20566_not ; n20568
g20505 nor n20567 n20568 ; n20569
g20506 and n20029 n20031_not ; n20570
g20507 nor n20032 n20570 ; n20571
g20508 and n20569_not n20571 ; n20572
g20509 nor n20569 n20572 ; n20573
g20510 and n20571 n20572_not ; n20574
g20511 nor n20573 n20574 ; n20575
g20512 nor n20016 n20028 ; n20576
g20513 nor n20027 n20028 ; n20577
g20514 nor n20576 n20577 ; n20578
g20515 and n9331 n12561 ; n20579
g20516 and n8418 n12567 ; n20580
g20517 and n8860 n12564 ; n20581
g20518 nor n20580 n20581 ; n20582
g20519 and n20579_not n20582 ; n20583
g20520 and n8421_not n20583 ; n20584
g20521 and n15905 n20583 ; n20585
g20522 nor n20584 n20585 ; n20586
g20523 and a[8] n20586_not ; n20587
g20524 and a[8]_not n20586 ; n20588
g20525 nor n20587 n20588 ; n20589
g20526 nor n20578 n20589 ; n20590
g20527 and n9331 n12564 ; n20591
g20528 and n8418 n12571 ; n20592
g20529 and n8860 n12567 ; n20593
g20530 nor n20592 n20593 ; n20594
g20531 and n20591_not n20594 ; n20595
g20532 and n8421 n15944_not ; n20596
g20533 and n20595 n20596_not ; n20597
g20534 and a[8] n20597_not ; n20598
g20535 nor n20597 n20598 ; n20599
g20536 and a[8] n20598_not ; n20600
g20537 nor n20599 n20600 ; n20601
g20538 and n20000_not n20011 ; n20602
g20539 nor n20012 n20602 ; n20603
g20540 and n20601_not n20603 ; n20604
g20541 nor n20601 n20604 ; n20605
g20542 and n20603 n20604_not ; n20606
g20543 nor n20605 n20606 ; n20607
g20544 and n19997 n19999_not ; n20608
g20545 nor n20000 n20608 ; n20609
g20546 and n9331 n12567 ; n20610
g20547 and n8418 n12574 ; n20611
g20548 and n8860 n12571 ; n20612
g20549 nor n20611 n20612 ; n20613
g20550 and n20610_not n20613 ; n20614
g20551 and n8421_not n20614 ; n20615
g20552 and n15989_not n20614 ; n20616
g20553 nor n20615 n20616 ; n20617
g20554 and a[8] n20617_not ; n20618
g20555 and a[8]_not n20617 ; n20619
g20556 nor n20618 n20619 ; n20620
g20557 and n20609 n20620_not ; n20621
g20558 and n8860 n12581_not ; n20622
g20559 and n9331 n12577 ; n20623
g20560 nor n20622 n20623 ; n20624
g20561 and n8421 n16085_not ; n20625
g20562 and n20624 n20625_not ; n20626
g20563 and a[8] n20626_not ; n20627
g20564 and a[8] n20627_not ; n20628
g20565 nor n20626 n20627 ; n20629
g20566 nor n20628 n20629 ; n20630
g20567 nor n8416 n12581 ; n20631
g20568 and a[8] n20631_not ; n20632
g20569 and n20630_not n20632 ; n20633
g20570 and n9331 n12574 ; n20634
g20571 and n8418 n12581_not ; n20635
g20572 and n8860 n12577 ; n20636
g20573 nor n20635 n20636 ; n20637
g20574 and n20634_not n20637 ; n20638
g20575 and n8421_not n20638 ; n20639
g20576 and n16094 n20638 ; n20640
g20577 nor n20639 n20640 ; n20641
g20578 and a[8] n20641_not ; n20642
g20579 and a[8]_not n20641 ; n20643
g20580 nor n20642 n20643 ; n20644
g20581 and n20633 n20644_not ; n20645
g20582 and n19998 n20645 ; n20646
g20583 and n20645 n20646_not ; n20647
g20584 and n19998 n20646_not ; n20648
g20585 nor n20647 n20648 ; n20649
g20586 and n9331 n12571 ; n20650
g20587 and n8418 n12577 ; n20651
g20588 and n8860 n12574 ; n20652
g20589 nor n20651 n20652 ; n20653
g20590 and n20650_not n20653 ; n20654
g20591 and n8421 n16013 ; n20655
g20592 and n20654 n20655_not ; n20656
g20593 and a[8] n20656_not ; n20657
g20594 and a[8] n20657_not ; n20658
g20595 nor n20656 n20657 ; n20659
g20596 nor n20658 n20659 ; n20660
g20597 nor n20649 n20660 ; n20661
g20598 nor n20646 n20661 ; n20662
g20599 and n20609_not n20620 ; n20663
g20600 nor n20621 n20663 ; n20664
g20601 and n20662_not n20664 ; n20665
g20602 nor n20621 n20665 ; n20666
g20603 nor n20607 n20666 ; n20667
g20604 nor n20604 n20667 ; n20668
g20605 and n20578 n20589 ; n20669
g20606 nor n20590 n20669 ; n20670
g20607 and n20668_not n20670 ; n20671
g20608 nor n20590 n20671 ; n20672
g20609 nor n20575 n20672 ; n20673
g20610 nor n20572 n20673 ; n20674
g20611 and n20546 n20558_not ; n20675
g20612 nor n20557 n20558 ; n20676
g20613 nor n20675 n20676 ; n20677
g20614 nor n20674 n20677 ; n20678
g20615 nor n20558 n20678 ; n20679
g20616 and n20532 n20544_not ; n20680
g20617 nor n20543 n20544 ; n20681
g20618 nor n20680 n20681 ; n20682
g20619 nor n20679 n20682 ; n20683
g20620 nor n20544 n20683 ; n20684
g20621 and n20518_not n20529 ; n20685
g20622 nor n20530 n20685 ; n20686
g20623 and n20684_not n20686 ; n20687
g20624 nor n20530 n20687 ; n20688
g20625 nor n20516 n20688 ; n20689
g20626 nor n20513 n20689 ; n20690
g20627 nor n20498 n20690 ; n20691
g20628 nor n20495 n20691 ; n20692
g20629 nor n20480 n20692 ; n20693
g20630 nor n20477 n20693 ; n20694
g20631 and n20451 n20463_not ; n20695
g20632 nor n20462 n20463 ; n20696
g20633 nor n20695 n20696 ; n20697
g20634 nor n20694 n20697 ; n20698
g20635 nor n20463 n20698 ; n20699
g20636 and n20437 n20449_not ; n20700
g20637 nor n20448 n20449 ; n20701
g20638 nor n20700 n20701 ; n20702
g20639 nor n20699 n20702 ; n20703
g20640 nor n20449 n20703 ; n20704
g20641 and n20423_not n20434 ; n20705
g20642 nor n20435 n20705 ; n20706
g20643 and n20704_not n20706 ; n20707
g20644 nor n20435 n20707 ; n20708
g20645 nor n20421 n20708 ; n20709
g20646 nor n20418 n20709 ; n20710
g20647 nor n20403 n20710 ; n20711
g20648 nor n20400 n20711 ; n20712
g20649 nor n20385 n20712 ; n20713
g20650 nor n20382 n20713 ; n20714
g20651 and n20356 n20368_not ; n20715
g20652 nor n20367 n20368 ; n20716
g20653 nor n20715 n20716 ; n20717
g20654 nor n20714 n20717 ; n20718
g20655 nor n20368 n20718 ; n20719
g20656 and n20342 n20354_not ; n20720
g20657 nor n20353 n20354 ; n20721
g20658 nor n20720 n20721 ; n20722
g20659 nor n20719 n20722 ; n20723
g20660 nor n20354 n20723 ; n20724
g20661 and n20328_not n20339 ; n20725
g20662 nor n20340 n20725 ; n20726
g20663 and n20724_not n20726 ; n20727
g20664 nor n20340 n20727 ; n20728
g20665 nor n20326 n20728 ; n20729
g20666 nor n20323 n20729 ; n20730
g20667 nor n20308 n20730 ; n20731
g20668 nor n20305 n20731 ; n20732
g20669 and n20279 n20291_not ; n20733
g20670 nor n20290 n20291 ; n20734
g20671 nor n20733 n20734 ; n20735
g20672 nor n20732 n20735 ; n20736
g20673 nor n20291 n20736 ; n20737
g20674 and n20265 n20277_not ; n20738
g20675 nor n20276 n20277 ; n20739
g20676 nor n20738 n20739 ; n20740
g20677 nor n20737 n20740 ; n20741
g20678 nor n20277 n20741 ; n20742
g20679 and n20251 n20263_not ; n20743
g20680 nor n20262 n20263 ; n20744
g20681 nor n20743 n20744 ; n20745
g20682 nor n20742 n20745 ; n20746
g20683 nor n20263 n20746 ; n20747
g20684 and n20237 n20249_not ; n20748
g20685 nor n20248 n20249 ; n20749
g20686 nor n20748 n20749 ; n20750
g20687 nor n20747 n20750 ; n20751
g20688 nor n20249 n20751 ; n20752
g20689 and n20223 n20235_not ; n20753
g20690 nor n20234 n20235 ; n20754
g20691 nor n20753 n20754 ; n20755
g20692 nor n20752 n20755 ; n20756
g20693 nor n20235 n20756 ; n20757
g20694 and n20209 n20221_not ; n20758
g20695 nor n20220 n20221 ; n20759
g20696 nor n20758 n20759 ; n20760
g20697 nor n20757 n20760 ; n20761
g20698 nor n20221 n20761 ; n20762
g20699 and n20195 n20207_not ; n20763
g20700 nor n20206 n20207 ; n20764
g20701 nor n20763 n20764 ; n20765
g20702 nor n20762 n20765 ; n20766
g20703 nor n20207 n20766 ; n20767
g20704 and n20181 n20193_not ; n20768
g20705 nor n20192 n20193 ; n20769
g20706 nor n20768 n20769 ; n20770
g20707 nor n20767 n20770 ; n20771
g20708 nor n20193 n20771 ; n20772
g20709 and n20167 n20179_not ; n20773
g20710 nor n20178 n20179 ; n20774
g20711 nor n20773 n20774 ; n20775
g20712 nor n20772 n20775 ; n20776
g20713 nor n20179 n20776 ; n20777
g20714 and n20153_not n20164 ; n20778
g20715 nor n20165 n20778 ; n20779
g20716 and n20777_not n20779 ; n20780
g20717 nor n20165 n20780 ; n20781
g20718 nor n20151 n20781 ; n20782
g20719 and n20151 n20781 ; n20783
g20720 nor n20782 n20783 ; n20784
g20721 and n71 n13941 ; n20785
g20722 and n9867 n13633 ; n20786
g20723 and n10434 n13627_not ; n20787
g20724 nor n20786 n20787 ; n20788
g20725 and n20785_not n20788 ; n20789
g20726 and n9870 n14136 ; n20790
g20727 and n20789 n20790_not ; n20791
g20728 and a[5] n20791_not ; n20792
g20729 and a[5] n20792_not ; n20793
g20730 nor n20791 n20792 ; n20794
g20731 nor n20793 n20794 ; n20795
g20732 and n20784 n20795_not ; n20796
g20733 nor n20782 n20796 ; n20797
g20734 nor n20148 n20797 ; n20798
g20735 and n20148 n20797 ; n20799
g20736 nor n20798 n20799 ; n20800
g20737 and n20784 n20796_not ; n20801
g20738 nor n20795 n20796 ; n20802
g20739 nor n20801 n20802 ; n20803
g20740 and n71 n13627_not ; n20804
g20741 and n9867 n13630 ; n20805
g20742 and n10434 n13633 ; n20806
g20743 nor n20805 n20806 ; n20807
g20744 and n20804_not n20807 ; n20808
g20745 and n9870 n13654_not ; n20809
g20746 and n20808 n20809_not ; n20810
g20747 and a[5] n20810_not ; n20811
g20748 nor n20810 n20811 ; n20812
g20749 and a[5] n20811_not ; n20813
g20750 nor n20812 n20813 ; n20814
g20751 and n20777 n20779_not ; n20815
g20752 nor n20780 n20815 ; n20816
g20753 and n20814_not n20816 ; n20817
g20754 nor n20814 n20817 ; n20818
g20755 and n20816 n20817_not ; n20819
g20756 nor n20818 n20819 ; n20820
g20757 nor n11715 n11727 ; n20821
g20758 nor n13438 n20821 ; n20822
g20759 and n11055 n13941 ; n20823
g20760 nor n20822 n20823 ; n20824
g20761 and n11057 n13951_not ; n20825
g20762 and n20824 n20825_not ; n20826
g20763 and a[2] n20826_not ; n20827
g20764 and a[2] n20827_not ; n20828
g20765 nor n20826 n20827 ; n20829
g20766 nor n20828 n20829 ; n20830
g20767 nor n20820 n20830 ; n20831
g20768 nor n20817 n20831 ; n20832
g20769 nor n20803 n20832 ; n20833
g20770 and n20803 n20832 ; n20834
g20771 nor n20833 n20834 ; n20835
g20772 nor n20820 n20831 ; n20836
g20773 nor n20830 n20831 ; n20837
g20774 nor n20836 n20837 ; n20838
g20775 and n71 n13633 ; n20839
g20776 and n9867 n13597 ; n20840
g20777 and n10434 n13630 ; n20841
g20778 nor n20840 n20841 ; n20842
g20779 and n20839_not n20842 ; n20843
g20780 and n9870 n13929 ; n20844
g20781 and n20843 n20844_not ; n20845
g20782 and a[5] n20845_not ; n20846
g20783 nor n20845 n20846 ; n20847
g20784 and a[5] n20846_not ; n20848
g20785 nor n20847 n20848 ; n20849
g20786 nor n20772 n20776 ; n20850
g20787 nor n20775 n20776 ; n20851
g20788 nor n20850 n20851 ; n20852
g20789 nor n20849 n20852 ; n20853
g20790 nor n20849 n20853 ; n20854
g20791 nor n20852 n20853 ; n20855
g20792 nor n20854 n20855 ; n20856
g20793 and n71 n13630 ; n20857
g20794 and n9867 n13515 ; n20858
g20795 and n10434 n13597 ; n20859
g20796 nor n20858 n20859 ; n20860
g20797 and n20857_not n20860 ; n20861
g20798 and n9870 n13976 ; n20862
g20799 and n20861 n20862_not ; n20863
g20800 and a[5] n20863_not ; n20864
g20801 nor n20863 n20864 ; n20865
g20802 and a[5] n20864_not ; n20866
g20803 nor n20865 n20866 ; n20867
g20804 nor n20767 n20771 ; n20868
g20805 nor n20770 n20771 ; n20869
g20806 nor n20868 n20869 ; n20870
g20807 nor n20867 n20870 ; n20871
g20808 nor n20867 n20871 ; n20872
g20809 nor n20870 n20871 ; n20873
g20810 nor n20872 n20873 ; n20874
g20811 and n71 n13597 ; n20875
g20812 and n9867 n13521 ; n20876
g20813 and n10434 n13515 ; n20877
g20814 nor n20876 n20877 ; n20878
g20815 and n20875_not n20878 ; n20879
g20816 and n9870 n13612_not ; n20880
g20817 and n20879 n20880_not ; n20881
g20818 and a[5] n20881_not ; n20882
g20819 nor n20881 n20882 ; n20883
g20820 and a[5] n20882_not ; n20884
g20821 nor n20883 n20884 ; n20885
g20822 nor n20762 n20766 ; n20886
g20823 nor n20765 n20766 ; n20887
g20824 nor n20886 n20887 ; n20888
g20825 nor n20885 n20888 ; n20889
g20826 nor n20885 n20889 ; n20890
g20827 nor n20888 n20889 ; n20891
g20828 nor n20890 n20891 ; n20892
g20829 and n71 n13515 ; n20893
g20830 and n9867 n13518 ; n20894
g20831 and n10434 n13521 ; n20895
g20832 nor n20894 n20895 ; n20896
g20833 and n20893_not n20896 ; n20897
g20834 and n9870 n13541 ; n20898
g20835 and n20897 n20898_not ; n20899
g20836 and a[5] n20899_not ; n20900
g20837 nor n20899 n20900 ; n20901
g20838 and a[5] n20900_not ; n20902
g20839 nor n20901 n20902 ; n20903
g20840 nor n20757 n20761 ; n20904
g20841 nor n20760 n20761 ; n20905
g20842 nor n20904 n20905 ; n20906
g20843 nor n20903 n20906 ; n20907
g20844 nor n20903 n20907 ; n20908
g20845 nor n20906 n20907 ; n20909
g20846 nor n20908 n20909 ; n20910
g20847 and n71 n13521 ; n20911
g20848 and n9867 n13491 ; n20912
g20849 and n10434 n13518 ; n20913
g20850 nor n20912 n20913 ; n20914
g20851 and n20911_not n20914 ; n20915
g20852 and n9870 n13909_not ; n20916
g20853 and n20915 n20916_not ; n20917
g20854 and a[5] n20917_not ; n20918
g20855 nor n20917 n20918 ; n20919
g20856 and a[5] n20918_not ; n20920
g20857 nor n20919 n20920 ; n20921
g20858 nor n20752 n20756 ; n20922
g20859 nor n20755 n20756 ; n20923
g20860 nor n20922 n20923 ; n20924
g20861 nor n20921 n20924 ; n20925
g20862 nor n20921 n20925 ; n20926
g20863 nor n20924 n20925 ; n20927
g20864 nor n20926 n20927 ; n20928
g20865 and n71 n13518 ; n20929
g20866 and n9867 n12889 ; n20930
g20867 and n10434 n13491 ; n20931
g20868 nor n20930 n20931 ; n20932
g20869 and n20929_not n20932 ; n20933
g20870 and n9870 n13584 ; n20934
g20871 and n20933 n20934_not ; n20935
g20872 and a[5] n20935_not ; n20936
g20873 nor n20935 n20936 ; n20937
g20874 and a[5] n20936_not ; n20938
g20875 nor n20937 n20938 ; n20939
g20876 nor n20747 n20751 ; n20940
g20877 nor n20750 n20751 ; n20941
g20878 nor n20940 n20941 ; n20942
g20879 nor n20939 n20942 ; n20943
g20880 nor n20939 n20943 ; n20944
g20881 nor n20942 n20943 ; n20945
g20882 nor n20944 n20945 ; n20946
g20883 and n71 n13491 ; n20947
g20884 and n9867 n12769 ; n20948
g20885 and n10434 n12889 ; n20949
g20886 nor n20948 n20949 ; n20950
g20887 and n20947_not n20950 ; n20951
g20888 and n9870 n13503_not ; n20952
g20889 and n20951 n20952_not ; n20953
g20890 and a[5] n20953_not ; n20954
g20891 nor n20953 n20954 ; n20955
g20892 and a[5] n20954_not ; n20956
g20893 nor n20955 n20956 ; n20957
g20894 nor n20742 n20746 ; n20958
g20895 nor n20745 n20746 ; n20959
g20896 nor n20958 n20959 ; n20960
g20897 nor n20957 n20960 ; n20961
g20898 nor n20957 n20961 ; n20962
g20899 nor n20960 n20961 ; n20963
g20900 nor n20962 n20963 ; n20964
g20901 and n71 n12889 ; n20965
g20902 and n9867 n12502 ; n20966
g20903 and n10434 n12769 ; n20967
g20904 nor n20966 n20967 ; n20968
g20905 and n20965_not n20968 ; n20969
g20906 and n9870 n12895 ; n20970
g20907 and n20969 n20970_not ; n20971
g20908 and a[5] n20971_not ; n20972
g20909 nor n20971 n20972 ; n20973
g20910 and a[5] n20972_not ; n20974
g20911 nor n20973 n20974 ; n20975
g20912 nor n20737 n20741 ; n20976
g20913 nor n20740 n20741 ; n20977
g20914 nor n20976 n20977 ; n20978
g20915 nor n20975 n20978 ; n20979
g20916 nor n20975 n20979 ; n20980
g20917 nor n20978 n20979 ; n20981
g20918 nor n20980 n20981 ; n20982
g20919 and n71 n12769 ; n20983
g20920 and n9867 n12370 ; n20984
g20921 and n10434 n12502 ; n20985
g20922 nor n20984 n20985 ; n20986
g20923 and n20983_not n20986 ; n20987
g20924 and n9870 n12999 ; n20988
g20925 and n20987 n20988_not ; n20989
g20926 and a[5] n20989_not ; n20990
g20927 nor n20989 n20990 ; n20991
g20928 and a[5] n20990_not ; n20992
g20929 nor n20991 n20992 ; n20993
g20930 nor n20732 n20736 ; n20994
g20931 nor n20735 n20736 ; n20995
g20932 nor n20994 n20995 ; n20996
g20933 nor n20993 n20996 ; n20997
g20934 nor n20993 n20997 ; n20998
g20935 nor n20996 n20997 ; n20999
g20936 nor n20998 n20999 ; n21000
g20937 and n20308 n20730 ; n21001
g20938 nor n20731 n21001 ; n21002
g20939 and n71 n12502 ; n21003
g20940 and n9867 n12505 ; n21004
g20941 and n10434 n12370 ; n21005
g20942 nor n21004 n21005 ; n21006
g20943 and n21003_not n21006 ; n21007
g20944 and n9870_not n21007 ; n21008
g20945 and n13736 n21007 ; n21009
g20946 nor n21008 n21009 ; n21010
g20947 and a[5] n21010_not ; n21011
g20948 and a[5]_not n21010 ; n21012
g20949 nor n21011 n21012 ; n21013
g20950 and n21002 n21013_not ; n21014
g20951 and n20326 n20728 ; n21015
g20952 nor n20729 n21015 ; n21016
g20953 and n71 n12370 ; n21017
g20954 and n9867 n12508 ; n21018
g20955 and n10434 n12505 ; n21019
g20956 nor n21018 n21019 ; n21020
g20957 and n21017_not n21020 ; n21021
g20958 and n9870_not n21021 ; n21022
g20959 and n13748 n21021 ; n21023
g20960 nor n21022 n21023 ; n21024
g20961 and a[5] n21024_not ; n21025
g20962 and a[5]_not n21024 ; n21026
g20963 nor n21025 n21026 ; n21027
g20964 and n21016 n21027_not ; n21028
g20965 and n71 n12505 ; n21029
g20966 and n9867 n12513 ; n21030
g20967 and n10434 n12508 ; n21031
g20968 nor n21030 n21031 ; n21032
g20969 and n21029_not n21032 ; n21033
g20970 and n9870 n14051_not ; n21034
g20971 and n21033 n21034_not ; n21035
g20972 and a[5] n21035_not ; n21036
g20973 nor n21035 n21036 ; n21037
g20974 and a[5] n21036_not ; n21038
g20975 nor n21037 n21038 ; n21039
g20976 and n20724 n20726_not ; n21040
g20977 nor n20727 n21040 ; n21041
g20978 and n21039_not n21041 ; n21042
g20979 nor n21039 n21042 ; n21043
g20980 and n21041 n21042_not ; n21044
g20981 nor n21043 n21044 ; n21045
g20982 and n71 n12508 ; n21046
g20983 and n9867 n12511 ; n21047
g20984 and n10434 n12513 ; n21048
g20985 nor n21047 n21048 ; n21049
g20986 and n21046_not n21049 ; n21050
g20987 and n9870 n13863 ; n21051
g20988 and n21050 n21051_not ; n21052
g20989 and a[5] n21052_not ; n21053
g20990 nor n21052 n21053 ; n21054
g20991 and a[5] n21053_not ; n21055
g20992 nor n21054 n21055 ; n21056
g20993 nor n20719 n20723 ; n21057
g20994 nor n20722 n20723 ; n21058
g20995 nor n21057 n21058 ; n21059
g20996 nor n21056 n21059 ; n21060
g20997 nor n21056 n21060 ; n21061
g20998 nor n21059 n21060 ; n21062
g20999 nor n21061 n21062 ; n21063
g21000 and n71 n12513 ; n21064
g21001 and n9867 n12516 ; n21065
g21002 and n10434 n12511 ; n21066
g21003 nor n21065 n21066 ; n21067
g21004 and n21064_not n21067 ; n21068
g21005 and n9870 n14177 ; n21069
g21006 and n21068 n21069_not ; n21070
g21007 and a[5] n21070_not ; n21071
g21008 nor n21070 n21071 ; n21072
g21009 and a[5] n21071_not ; n21073
g21010 nor n21072 n21073 ; n21074
g21011 nor n20714 n20718 ; n21075
g21012 nor n20717 n20718 ; n21076
g21013 nor n21075 n21076 ; n21077
g21014 nor n21074 n21077 ; n21078
g21015 nor n21074 n21078 ; n21079
g21016 nor n21077 n21078 ; n21080
g21017 nor n21079 n21080 ; n21081
g21018 and n20385 n20712 ; n21082
g21019 nor n20713 n21082 ; n21083
g21020 and n71 n12511 ; n21084
g21021 and n9867 n12519 ; n21085
g21022 and n10434 n12516 ; n21086
g21023 nor n21085 n21086 ; n21087
g21024 and n21084_not n21087 ; n21088
g21025 and n9870_not n21088 ; n21089
g21026 and n14233 n21088 ; n21090
g21027 nor n21089 n21090 ; n21091
g21028 and a[5] n21091_not ; n21092
g21029 and a[5]_not n21091 ; n21093
g21030 nor n21092 n21093 ; n21094
g21031 and n21083 n21094_not ; n21095
g21032 and n20403 n20710 ; n21096
g21033 nor n20711 n21096 ; n21097
g21034 and n71 n12516 ; n21098
g21035 and n9867 n12522 ; n21099
g21036 and n10434 n12519 ; n21100
g21037 nor n21099 n21100 ; n21101
g21038 and n21098_not n21101 ; n21102
g21039 and n9870_not n21102 ; n21103
g21040 and n14443 n21102 ; n21104
g21041 nor n21103 n21104 ; n21105
g21042 and a[5] n21105_not ; n21106
g21043 and a[5]_not n21105 ; n21107
g21044 nor n21106 n21107 ; n21108
g21045 and n21097 n21108_not ; n21109
g21046 and n20421 n20708 ; n21110
g21047 nor n20709 n21110 ; n21111
g21048 and n71 n12519 ; n21112
g21049 and n9867 n12525 ; n21113
g21050 and n10434 n12522 ; n21114
g21051 nor n21113 n21114 ; n21115
g21052 and n21112_not n21115 ; n21116
g21053 and n9870_not n21116 ; n21117
g21054 and n14454_not n21116 ; n21118
g21055 nor n21117 n21118 ; n21119
g21056 and a[5] n21119_not ; n21120
g21057 and a[5]_not n21119 ; n21121
g21058 nor n21120 n21121 ; n21122
g21059 and n21111 n21122_not ; n21123
g21060 and n71 n12522 ; n21124
g21061 and n9867 n12528 ; n21125
g21062 and n10434 n12525 ; n21126
g21063 nor n21125 n21126 ; n21127
g21064 and n21124_not n21127 ; n21128
g21065 and n9870 n14837 ; n21129
g21066 and n21128 n21129_not ; n21130
g21067 and a[5] n21130_not ; n21131
g21068 nor n21130 n21131 ; n21132
g21069 and a[5] n21131_not ; n21133
g21070 nor n21132 n21133 ; n21134
g21071 and n20704 n20706_not ; n21135
g21072 nor n20707 n21135 ; n21136
g21073 and n21134_not n21136 ; n21137
g21074 nor n21134 n21137 ; n21138
g21075 and n21136 n21137_not ; n21139
g21076 nor n21138 n21139 ; n21140
g21077 and n71 n12525 ; n21141
g21078 and n9867 n12531 ; n21142
g21079 and n10434 n12528 ; n21143
g21080 nor n21142 n21143 ; n21144
g21081 and n21141_not n21144 ; n21145
g21082 and n9870 n14608 ; n21146
g21083 and n21145 n21146_not ; n21147
g21084 and a[5] n21147_not ; n21148
g21085 nor n21147 n21148 ; n21149
g21086 and a[5] n21148_not ; n21150
g21087 nor n21149 n21150 ; n21151
g21088 nor n20699 n20703 ; n21152
g21089 nor n20702 n20703 ; n21153
g21090 nor n21152 n21153 ; n21154
g21091 nor n21151 n21154 ; n21155
g21092 nor n21151 n21155 ; n21156
g21093 nor n21154 n21155 ; n21157
g21094 nor n21156 n21157 ; n21158
g21095 and n71 n12528 ; n21159
g21096 and n9867 n12534 ; n21160
g21097 and n10434 n12531 ; n21161
g21098 nor n21160 n21161 ; n21162
g21099 and n21159_not n21162 ; n21163
g21100 and n9870 n15003_not ; n21164
g21101 and n21163 n21164_not ; n21165
g21102 and a[5] n21165_not ; n21166
g21103 nor n21165 n21166 ; n21167
g21104 and a[5] n21166_not ; n21168
g21105 nor n21167 n21168 ; n21169
g21106 nor n20694 n20698 ; n21170
g21107 nor n20697 n20698 ; n21171
g21108 nor n21170 n21171 ; n21172
g21109 nor n21169 n21172 ; n21173
g21110 nor n21169 n21173 ; n21174
g21111 nor n21172 n21173 ; n21175
g21112 nor n21174 n21175 ; n21176
g21113 and n20480 n20692 ; n21177
g21114 nor n20693 n21177 ; n21178
g21115 and n71 n12531 ; n21179
g21116 and n9867 n12537 ; n21180
g21117 and n10434 n12534 ; n21181
g21118 nor n21180 n21181 ; n21182
g21119 and n21179_not n21182 ; n21183
g21120 and n9870_not n21183 ; n21184
g21121 and n15255_not n21183 ; n21185
g21122 nor n21184 n21185 ; n21186
g21123 and a[5] n21186_not ; n21187
g21124 and a[5]_not n21186 ; n21188
g21125 nor n21187 n21188 ; n21189
g21126 and n21178 n21189_not ; n21190
g21127 and n20498 n20690 ; n21191
g21128 nor n20691 n21191 ; n21192
g21129 and n71 n12534 ; n21193
g21130 and n9867 n12540 ; n21194
g21131 and n10434 n12537 ; n21195
g21132 nor n21194 n21195 ; n21196
g21133 and n21193_not n21196 ; n21197
g21134 and n9870_not n21197 ; n21198
g21135 and n15096 n21197 ; n21199
g21136 nor n21198 n21199 ; n21200
g21137 and a[5] n21200_not ; n21201
g21138 and a[5]_not n21200 ; n21202
g21139 nor n21201 n21202 ; n21203
g21140 and n21192 n21203_not ; n21204
g21141 and n20516 n20688 ; n21205
g21142 nor n20689 n21205 ; n21206
g21143 and n71 n12537 ; n21207
g21144 and n9867 n12543 ; n21208
g21145 and n10434 n12540 ; n21209
g21146 nor n21208 n21209 ; n21210
g21147 and n21207_not n21210 ; n21211
g21148 and n9870_not n21211 ; n21212
g21149 and n15385 n21211 ; n21213
g21150 nor n21212 n21213 ; n21214
g21151 and a[5] n21214_not ; n21215
g21152 and a[5]_not n21214 ; n21216
g21153 nor n21215 n21216 ; n21217
g21154 and n21206 n21217_not ; n21218
g21155 and n71 n12540 ; n21219
g21156 and n9867 n12546 ; n21220
g21157 and n10434 n12543 ; n21221
g21158 nor n21220 n21221 ; n21222
g21159 and n21219_not n21222 ; n21223
g21160 and n9870 n15708_not ; n21224
g21161 and n21223 n21224_not ; n21225
g21162 and a[5] n21225_not ; n21226
g21163 nor n21225 n21226 ; n21227
g21164 and a[5] n21226_not ; n21228
g21165 nor n21227 n21228 ; n21229
g21166 and n20684 n20686_not ; n21230
g21167 nor n20687 n21230 ; n21231
g21168 and n21229_not n21231 ; n21232
g21169 nor n21229 n21232 ; n21233
g21170 and n21231 n21232_not ; n21234
g21171 nor n21233 n21234 ; n21235
g21172 and n71 n12543 ; n21236
g21173 and n9867 n12549 ; n21237
g21174 and n10434 n12546 ; n21238
g21175 nor n21237 n21238 ; n21239
g21176 and n21236_not n21239 ; n21240
g21177 and n9870 n15724 ; n21241
g21178 and n21240 n21241_not ; n21242
g21179 and a[5] n21242_not ; n21243
g21180 nor n21242 n21243 ; n21244
g21181 and a[5] n21243_not ; n21245
g21182 nor n21244 n21245 ; n21246
g21183 nor n20679 n20683 ; n21247
g21184 nor n20682 n20683 ; n21248
g21185 nor n21247 n21248 ; n21249
g21186 nor n21246 n21249 ; n21250
g21187 nor n21246 n21250 ; n21251
g21188 nor n21249 n21250 ; n21252
g21189 nor n21251 n21252 ; n21253
g21190 and n71 n12546 ; n21254
g21191 and n9867 n12552 ; n21255
g21192 and n10434 n12549 ; n21256
g21193 nor n21255 n21256 ; n21257
g21194 and n21254_not n21257 ; n21258
g21195 and n9870 n15356_not ; n21259
g21196 and n21258 n21259_not ; n21260
g21197 and a[5] n21260_not ; n21261
g21198 nor n21260 n21261 ; n21262
g21199 and a[5] n21261_not ; n21263
g21200 nor n21262 n21263 ; n21264
g21201 nor n20674 n20678 ; n21265
g21202 nor n20677 n20678 ; n21266
g21203 nor n21265 n21266 ; n21267
g21204 nor n21264 n21267 ; n21268
g21205 nor n21264 n21268 ; n21269
g21206 nor n21267 n21268 ; n21270
g21207 nor n21269 n21270 ; n21271
g21208 and n20575 n20672 ; n21272
g21209 nor n20673 n21272 ; n21273
g21210 and n71 n12549 ; n21274
g21211 and n9867 n12555 ; n21275
g21212 and n10434 n12552 ; n21276
g21213 nor n21275 n21276 ; n21277
g21214 and n21274_not n21277 ; n21278
g21215 and n9870_not n21278 ; n21279
g21216 and n15764_not n21278 ; n21280
g21217 nor n21279 n21280 ; n21281
g21218 and a[5] n21281_not ; n21282
g21219 and a[5]_not n21281 ; n21283
g21220 nor n21282 n21283 ; n21284
g21221 and n21273 n21284_not ; n21285
g21222 and n20668 n20670_not ; n21286
g21223 nor n20671 n21286 ; n21287
g21224 and n71 n12552 ; n21288
g21225 and n9867 n12558 ; n21289
g21226 and n10434 n12555 ; n21290
g21227 nor n21289 n21290 ; n21291
g21228 and n21288_not n21291 ; n21292
g21229 and n9870_not n21292 ; n21293
g21230 and n15791 n21292 ; n21294
g21231 nor n21293 n21294 ; n21295
g21232 and a[5] n21295_not ; n21296
g21233 and a[5]_not n21295 ; n21297
g21234 nor n21296 n21297 ; n21298
g21235 and n21287 n21298_not ; n21299
g21236 and n20607 n20666 ; n21300
g21237 nor n20667 n21300 ; n21301
g21238 and n71 n12555 ; n21302
g21239 and n9867 n12561 ; n21303
g21240 and n10434 n12558 ; n21304
g21241 nor n21303 n21304 ; n21305
g21242 and n21302_not n21305 ; n21306
g21243 and n9870_not n21306 ; n21307
g21244 and n15816 n21306 ; n21308
g21245 nor n21307 n21308 ; n21309
g21246 and a[5] n21309_not ; n21310
g21247 and a[5]_not n21309 ; n21311
g21248 nor n21310 n21311 ; n21312
g21249 and n21301 n21312_not ; n21313
g21250 and n71 n12558 ; n21314
g21251 and n9867 n12564 ; n21315
g21252 and n10434 n12561 ; n21316
g21253 nor n21315 n21316 ; n21317
g21254 and n21314_not n21317 ; n21318
g21255 and n9870 n15847 ; n21319
g21256 and n21318 n21319_not ; n21320
g21257 and a[5] n21320_not ; n21321
g21258 nor n21320 n21321 ; n21322
g21259 and a[5] n21321_not ; n21323
g21260 nor n21322 n21323 ; n21324
g21261 and n20662 n20664_not ; n21325
g21262 nor n20665 n21325 ; n21326
g21263 and n21324_not n21326 ; n21327
g21264 nor n21324 n21327 ; n21328
g21265 and n21326 n21327_not ; n21329
g21266 nor n21328 n21329 ; n21330
g21267 nor n20649 n20661 ; n21331
g21268 nor n20660 n20661 ; n21332
g21269 nor n21331 n21332 ; n21333
g21270 and n71 n12561 ; n21334
g21271 and n9867 n12567 ; n21335
g21272 and n10434 n12564 ; n21336
g21273 nor n21335 n21336 ; n21337
g21274 and n21334_not n21337 ; n21338
g21275 and n9870_not n21338 ; n21339
g21276 and n15905 n21338 ; n21340
g21277 nor n21339 n21340 ; n21341
g21278 and a[5] n21341_not ; n21342
g21279 and a[5]_not n21341 ; n21343
g21280 nor n21342 n21343 ; n21344
g21281 nor n21333 n21344 ; n21345
g21282 and n71 n12564 ; n21346
g21283 and n9867 n12571 ; n21347
g21284 and n10434 n12567 ; n21348
g21285 nor n21347 n21348 ; n21349
g21286 and n21346_not n21349 ; n21350
g21287 and n9870 n15944_not ; n21351
g21288 and n21350 n21351_not ; n21352
g21289 and a[5] n21352_not ; n21353
g21290 nor n21352 n21353 ; n21354
g21291 and a[5] n21353_not ; n21355
g21292 nor n21354 n21355 ; n21356
g21293 and n20633_not n20644 ; n21357
g21294 nor n20645 n21357 ; n21358
g21295 and n21356_not n21358 ; n21359
g21296 nor n21356 n21359 ; n21360
g21297 and n21358 n21359_not ; n21361
g21298 nor n21360 n21361 ; n21362
g21299 and n20630 n20632_not ; n21363
g21300 nor n20633 n21363 ; n21364
g21301 and n71 n12567 ; n21365
g21302 and n9867 n12574 ; n21366
g21303 and n10434 n12571 ; n21367
g21304 nor n21366 n21367 ; n21368
g21305 and n21365_not n21368 ; n21369
g21306 and n9870_not n21369 ; n21370
g21307 and n15989_not n21369 ; n21371
g21308 nor n21370 n21371 ; n21372
g21309 and a[5] n21372_not ; n21373
g21310 and a[5]_not n21372 ; n21374
g21311 nor n21373 n21374 ; n21375
g21312 and n21364 n21375_not ; n21376
g21313 and n10434 n12581_not ; n21377
g21314 and n71 n12577 ; n21378
g21315 nor n21377 n21378 ; n21379
g21316 and n9870 n16085_not ; n21380
g21317 and n21379 n21380_not ; n21381
g21318 and a[5] n21381_not ; n21382
g21319 and a[5] n21382_not ; n21383
g21320 nor n21381 n21382 ; n21384
g21321 nor n21383 n21384 ; n21385
g21322 nor n70 n12581 ; n21386
g21323 and a[5] n21386_not ; n21387
g21324 and n21385_not n21387 ; n21388
g21325 and n71 n12574 ; n21389
g21326 and n9867 n12581_not ; n21390
g21327 and n10434 n12577 ; n21391
g21328 nor n21390 n21391 ; n21392
g21329 and n21389_not n21392 ; n21393
g21330 and n9870_not n21393 ; n21394
g21331 and n16094 n21393 ; n21395
g21332 nor n21394 n21395 ; n21396
g21333 and a[5] n21396_not ; n21397
g21334 and a[5]_not n21396 ; n21398
g21335 nor n21397 n21398 ; n21399
g21336 and n21388 n21399_not ; n21400
g21337 and n20631 n21400 ; n21401
g21338 and n21400 n21401_not ; n21402
g21339 and n20631 n21401_not ; n21403
g21340 nor n21402 n21403 ; n21404
g21341 and n71 n12571 ; n21405
g21342 and n9867 n12577 ; n21406
g21343 and n10434 n12574 ; n21407
g21344 nor n21406 n21407 ; n21408
g21345 and n21405_not n21408 ; n21409
g21346 and n9870 n16013 ; n21410
g21347 and n21409 n21410_not ; n21411
g21348 and a[5] n21411_not ; n21412
g21349 and a[5] n21412_not ; n21413
g21350 nor n21411 n21412 ; n21414
g21351 nor n21413 n21414 ; n21415
g21352 nor n21404 n21415 ; n21416
g21353 nor n21401 n21416 ; n21417
g21354 and n21364_not n21375 ; n21418
g21355 nor n21376 n21418 ; n21419
g21356 and n21417_not n21419 ; n21420
g21357 nor n21376 n21420 ; n21421
g21358 nor n21362 n21421 ; n21422
g21359 nor n21359 n21422 ; n21423
g21360 and n21333 n21344 ; n21424
g21361 nor n21345 n21424 ; n21425
g21362 and n21423_not n21425 ; n21426
g21363 nor n21345 n21426 ; n21427
g21364 nor n21330 n21427 ; n21428
g21365 nor n21327 n21428 ; n21429
g21366 and n21301 n21313_not ; n21430
g21367 nor n21312 n21313 ; n21431
g21368 nor n21430 n21431 ; n21432
g21369 nor n21429 n21432 ; n21433
g21370 nor n21313 n21433 ; n21434
g21371 and n21287 n21299_not ; n21435
g21372 nor n21298 n21299 ; n21436
g21373 nor n21435 n21436 ; n21437
g21374 nor n21434 n21437 ; n21438
g21375 nor n21299 n21438 ; n21439
g21376 and n21273_not n21284 ; n21440
g21377 nor n21285 n21440 ; n21441
g21378 and n21439_not n21441 ; n21442
g21379 nor n21285 n21442 ; n21443
g21380 nor n21271 n21443 ; n21444
g21381 nor n21268 n21444 ; n21445
g21382 nor n21253 n21445 ; n21446
g21383 nor n21250 n21446 ; n21447
g21384 nor n21235 n21447 ; n21448
g21385 nor n21232 n21448 ; n21449
g21386 and n21206 n21218_not ; n21450
g21387 nor n21217 n21218 ; n21451
g21388 nor n21450 n21451 ; n21452
g21389 nor n21449 n21452 ; n21453
g21390 nor n21218 n21453 ; n21454
g21391 and n21192 n21204_not ; n21455
g21392 nor n21203 n21204 ; n21456
g21393 nor n21455 n21456 ; n21457
g21394 nor n21454 n21457 ; n21458
g21395 nor n21204 n21458 ; n21459
g21396 and n21178_not n21189 ; n21460
g21397 nor n21190 n21460 ; n21461
g21398 and n21459_not n21461 ; n21462
g21399 nor n21190 n21462 ; n21463
g21400 nor n21176 n21463 ; n21464
g21401 nor n21173 n21464 ; n21465
g21402 nor n21158 n21465 ; n21466
g21403 nor n21155 n21466 ; n21467
g21404 nor n21140 n21467 ; n21468
g21405 nor n21137 n21468 ; n21469
g21406 and n21111 n21123_not ; n21470
g21407 nor n21122 n21123 ; n21471
g21408 nor n21470 n21471 ; n21472
g21409 nor n21469 n21472 ; n21473
g21410 nor n21123 n21473 ; n21474
g21411 and n21097 n21109_not ; n21475
g21412 nor n21108 n21109 ; n21476
g21413 nor n21475 n21476 ; n21477
g21414 nor n21474 n21477 ; n21478
g21415 nor n21109 n21478 ; n21479
g21416 and n21083_not n21094 ; n21480
g21417 nor n21095 n21480 ; n21481
g21418 and n21479_not n21481 ; n21482
g21419 nor n21095 n21482 ; n21483
g21420 nor n21081 n21483 ; n21484
g21421 nor n21078 n21484 ; n21485
g21422 nor n21063 n21485 ; n21486
g21423 nor n21060 n21486 ; n21487
g21424 nor n21045 n21487 ; n21488
g21425 nor n21042 n21488 ; n21489
g21426 and n21016 n21028_not ; n21490
g21427 nor n21027 n21028 ; n21491
g21428 nor n21490 n21491 ; n21492
g21429 nor n21489 n21492 ; n21493
g21430 nor n21028 n21493 ; n21494
g21431 and n21002_not n21013 ; n21495
g21432 nor n21014 n21495 ; n21496
g21433 and n21494_not n21496 ; n21497
g21434 nor n21014 n21497 ; n21498
g21435 nor n21000 n21498 ; n21499
g21436 nor n20997 n21499 ; n21500
g21437 nor n20982 n21500 ; n21501
g21438 nor n20979 n21501 ; n21502
g21439 nor n20964 n21502 ; n21503
g21440 nor n20961 n21503 ; n21504
g21441 nor n20946 n21504 ; n21505
g21442 nor n20943 n21505 ; n21506
g21443 nor n20928 n21506 ; n21507
g21444 nor n20925 n21507 ; n21508
g21445 nor n20910 n21508 ; n21509
g21446 nor n20907 n21509 ; n21510
g21447 nor n20892 n21510 ; n21511
g21448 nor n20889 n21511 ; n21512
g21449 nor n20874 n21512 ; n21513
g21450 nor n20871 n21513 ; n21514
g21451 nor n20856 n21514 ; n21515
g21452 nor n20853 n21515 ; n21516
g21453 nor n20838 n21516 ; n21517
g21454 and n20838 n21516 ; n21518
g21455 nor n21517 n21518 ; n21519
g21456 and n20856 n21514 ; n21520
g21457 nor n21515 n21520 ; n21521
g21458 and n11727 n13438_not ; n21522
g21459 and n11055 n13627_not ; n21523
g21460 and n11715 n13941 ; n21524
g21461 nor n21523 n21524 ; n21525
g21462 and n21522_not n21525 ; n21526
g21463 and n11057_not n21526 ; n21527
g21464 and n14028_not n21526 ; n21528
g21465 nor n21527 n21528 ; n21529
g21466 and a[2] n21529_not ; n21530
g21467 and a[2]_not n21529 ; n21531
g21468 nor n21530 n21531 ; n21532
g21469 and n21521 n21532_not ; n21533
g21470 and n20874 n21512 ; n21534
g21471 nor n21513 n21534 ; n21535
g21472 and n11727 n13941 ; n21536
g21473 and n11055 n13633 ; n21537
g21474 and n11715 n13627_not ; n21538
g21475 nor n21537 n21538 ; n21539
g21476 and n21536_not n21539 ; n21540
g21477 and n11057_not n21540 ; n21541
g21478 and n14136_not n21540 ; n21542
g21479 nor n21541 n21542 ; n21543
g21480 and a[2] n21543_not ; n21544
g21481 and a[2]_not n21543 ; n21545
g21482 nor n21544 n21545 ; n21546
g21483 and n21535 n21546_not ; n21547
g21484 and n20892 n21510 ; n21548
g21485 nor n21511 n21548 ; n21549
g21486 and n11727 n13627_not ; n21550
g21487 and n11055 n13630 ; n21551
g21488 and n11715 n13633 ; n21552
g21489 nor n21551 n21552 ; n21553
g21490 and n21550_not n21553 ; n21554
g21491 and n11057_not n21554 ; n21555
g21492 and n13654 n21554 ; n21556
g21493 nor n21555 n21556 ; n21557
g21494 and a[2] n21557_not ; n21558
g21495 and a[2]_not n21557 ; n21559
g21496 nor n21558 n21559 ; n21560
g21497 and n21549 n21560_not ; n21561
g21498 and n20910 n21508 ; n21562
g21499 nor n21509 n21562 ; n21563
g21500 and n11727 n13633 ; n21564
g21501 and n11055 n13597 ; n21565
g21502 and n11715 n13630 ; n21566
g21503 nor n21565 n21566 ; n21567
g21504 and n21564_not n21567 ; n21568
g21505 and n11057_not n21568 ; n21569
g21506 and n13929_not n21568 ; n21570
g21507 nor n21569 n21570 ; n21571
g21508 and a[2] n21571_not ; n21572
g21509 and a[2]_not n21571 ; n21573
g21510 nor n21572 n21573 ; n21574
g21511 and n21563 n21574_not ; n21575
g21512 and n20928 n21506 ; n21576
g21513 nor n21507 n21576 ; n21577
g21514 and n11727 n13630 ; n21578
g21515 and n11055 n13515 ; n21579
g21516 and n11715 n13597 ; n21580
g21517 nor n21579 n21580 ; n21581
g21518 and n21578_not n21581 ; n21582
g21519 and n11057_not n21582 ; n21583
g21520 and n13976_not n21582 ; n21584
g21521 nor n21583 n21584 ; n21585
g21522 and a[2] n21585_not ; n21586
g21523 and a[2]_not n21585 ; n21587
g21524 nor n21586 n21587 ; n21588
g21525 and n21577 n21588_not ; n21589
g21526 and n20946 n21504 ; n21590
g21527 nor n21505 n21590 ; n21591
g21528 and n11727 n13597 ; n21592
g21529 and n11055 n13521 ; n21593
g21530 and n11715 n13515 ; n21594
g21531 nor n21593 n21594 ; n21595
g21532 and n21592_not n21595 ; n21596
g21533 and n11057_not n21596 ; n21597
g21534 and n13612 n21596 ; n21598
g21535 nor n21597 n21598 ; n21599
g21536 and a[2] n21599_not ; n21600
g21537 and a[2]_not n21599 ; n21601
g21538 nor n21600 n21601 ; n21602
g21539 and n21591 n21602_not ; n21603
g21540 and n20964 n21502 ; n21604
g21541 nor n21503 n21604 ; n21605
g21542 and n11727 n13515 ; n21606
g21543 and n11055 n13518 ; n21607
g21544 and n11715 n13521 ; n21608
g21545 nor n21607 n21608 ; n21609
g21546 and n21606_not n21609 ; n21610
g21547 and n11057_not n21610 ; n21611
g21548 and n13541_not n21610 ; n21612
g21549 nor n21611 n21612 ; n21613
g21550 and a[2] n21613_not ; n21614
g21551 and a[2]_not n21613 ; n21615
g21552 nor n21614 n21615 ; n21616
g21553 and n21605 n21616_not ; n21617
g21554 and n20982 n21500 ; n21618
g21555 nor n21501 n21618 ; n21619
g21556 and n11727 n13521 ; n21620
g21557 and n11055 n13491 ; n21621
g21558 and n11715 n13518 ; n21622
g21559 nor n21621 n21622 ; n21623
g21560 and n21620_not n21623 ; n21624
g21561 and n11057_not n21624 ; n21625
g21562 and n13909 n21624 ; n21626
g21563 nor n21625 n21626 ; n21627
g21564 and a[2] n21627_not ; n21628
g21565 and a[2]_not n21627 ; n21629
g21566 nor n21628 n21629 ; n21630
g21567 and n21619 n21630_not ; n21631
g21568 and n21000 n21498 ; n21632
g21569 nor n21499 n21632 ; n21633
g21570 and n11727 n13518 ; n21634
g21571 and n11055 n12889 ; n21635
g21572 and n11715 n13491 ; n21636
g21573 nor n21635 n21636 ; n21637
g21574 and n21634_not n21637 ; n21638
g21575 and n11057_not n21638 ; n21639
g21576 and n13584_not n21638 ; n21640
g21577 nor n21639 n21640 ; n21641
g21578 and a[2] n21641_not ; n21642
g21579 and a[2]_not n21641 ; n21643
g21580 nor n21642 n21643 ; n21644
g21581 and n21633 n21644_not ; n21645
g21582 and n21494 n21496_not ; n21646
g21583 nor n21497 n21646 ; n21647
g21584 and n21479 n21481_not ; n21648
g21585 nor n21482 n21648 ; n21649
g21586 and n21459 n21461_not ; n21650
g21587 nor n21462 n21650 ; n21651
g21588 and n21439 n21441_not ; n21652
g21589 nor n21442 n21652 ; n21653
g21590 and n21417 n21419_not ; n21654
g21591 nor n21420 n21654 ; n21655
g21592 and n21388_not n21399 ; n21656
g21593 nor n21400 n21656 ; n21657
g21594 nor n11794 n12581 ; n21658
g21595 and n11796 n16094_not ; n21659
g21596 and n11727 n12574 ; n21660
g21597 and n11055 n12581_not ; n21661
g21598 and n11715 n12577 ; n21662
g21599 nor n21661 n21662 ; n21663
g21600 and n21660_not n21663 ; n21664
g21601 and a[2] n21664_not ; n21665
g21602 and n11796 n16085_not ; n21666
g21603 and n11805 n12581_not ; n21667
g21604 and n11807 n12577 ; n21668
g21605 and a[2] n21668_not ; n21669
g21606 and n21667_not n21669 ; n21670
g21607 and n21666_not n21670 ; n21671
g21608 and n21665_not n21671 ; n21672
g21609 and n21659_not n21672 ; n21673
g21610 and n21658_not n21673 ; n21674
g21611 and n21386 n21674 ; n21675
g21612 nor n21386 n21674 ; n21676
g21613 and n11727 n12571 ; n21677
g21614 and n11055 n12577 ; n21678
g21615 and n11715 n12574 ; n21679
g21616 nor n21678 n21679 ; n21680
g21617 and n21677_not n21680 ; n21681
g21618 and n11057 n16013 ; n21682
g21619 and n21681 n21682_not ; n21683
g21620 nor a[2] n21683 ; n21684
g21621 and a[2] n21683 ; n21685
g21622 nor n21684 n21685 ; n21686
g21623 nor n21676 n21686 ; n21687
g21624 nor n21675 n21687 ; n21688
g21625 and n11727 n12567 ; n21689
g21626 and n11055 n12574 ; n21690
g21627 and n11715 n12571 ; n21691
g21628 nor n21690 n21691 ; n21692
g21629 and n21689_not n21692 ; n21693
g21630 and n11057_not n21693 ; n21694
g21631 and n15989_not n21693 ; n21695
g21632 nor n21694 n21695 ; n21696
g21633 and a[2] n21696_not ; n21697
g21634 and a[2]_not n21696 ; n21698
g21635 nor n21697 n21698 ; n21699
g21636 and n21688 n21699 ; n21700
g21637 and n21385 n21387_not ; n21701
g21638 nor n21388 n21701 ; n21702
g21639 and n21700_not n21702 ; n21703
g21640 nor n21688 n21699 ; n21704
g21641 nor n21703 n21704 ; n21705
g21642 and n21657 n21705_not ; n21706
g21643 and n21657_not n21705 ; n21707
g21644 and n11727 n12564 ; n21708
g21645 and n11055 n12571 ; n21709
g21646 and n11715 n12567 ; n21710
g21647 nor n21709 n21710 ; n21711
g21648 and n21708_not n21711 ; n21712
g21649 and n11057 n15944_not ; n21713
g21650 and n21712 n21713_not ; n21714
g21651 nor a[2] n21714 ; n21715
g21652 and a[2] n21714 ; n21716
g21653 nor n21715 n21716 ; n21717
g21654 nor n21707 n21717 ; n21718
g21655 nor n21706 n21718 ; n21719
g21656 and n11727 n12561 ; n21720
g21657 and n11055 n12567 ; n21721
g21658 and n11715 n12564 ; n21722
g21659 nor n21721 n21722 ; n21723
g21660 and n21720_not n21723 ; n21724
g21661 and n11057_not n21724 ; n21725
g21662 and n15905 n21724 ; n21726
g21663 nor n21725 n21726 ; n21727
g21664 and a[2] n21727_not ; n21728
g21665 and a[2]_not n21727 ; n21729
g21666 nor n21728 n21729 ; n21730
g21667 nor n21719 n21730 ; n21731
g21668 and n21719 n21730 ; n21732
g21669 and n21404 n21415 ; n21733
g21670 nor n21416 n21733 ; n21734
g21671 and n21732_not n21734 ; n21735
g21672 nor n21731 n21735 ; n21736
g21673 and n21655 n21736_not ; n21737
g21674 and n21655_not n21736 ; n21738
g21675 and n11727 n12558 ; n21739
g21676 and n11055 n12564 ; n21740
g21677 and n11715 n12561 ; n21741
g21678 nor n21740 n21741 ; n21742
g21679 and n21739_not n21742 ; n21743
g21680 and n11057 n15847 ; n21744
g21681 and n21743 n21744_not ; n21745
g21682 nor a[2] n21745 ; n21746
g21683 and a[2] n21745 ; n21747
g21684 nor n21746 n21747 ; n21748
g21685 nor n21738 n21748 ; n21749
g21686 nor n21737 n21749 ; n21750
g21687 and n11727 n12555 ; n21751
g21688 and n11055 n12561 ; n21752
g21689 and n11715 n12558 ; n21753
g21690 nor n21752 n21753 ; n21754
g21691 and n21751_not n21754 ; n21755
g21692 and n11057_not n21755 ; n21756
g21693 and n15816 n21755 ; n21757
g21694 nor n21756 n21757 ; n21758
g21695 and a[2] n21758_not ; n21759
g21696 and a[2]_not n21758 ; n21760
g21697 nor n21759 n21760 ; n21761
g21698 and n21750 n21761 ; n21762
g21699 and n21362 n21421 ; n21763
g21700 nor n21422 n21763 ; n21764
g21701 and n21762_not n21764 ; n21765
g21702 nor n21750 n21761 ; n21766
g21703 nor n21765 n21766 ; n21767
g21704 and n11727 n12552 ; n21768
g21705 and n11055 n12558 ; n21769
g21706 and n11715 n12555 ; n21770
g21707 nor n21769 n21770 ; n21771
g21708 and n21768_not n21771 ; n21772
g21709 and n11057_not n21772 ; n21773
g21710 and n15791 n21772 ; n21774
g21711 nor n21773 n21774 ; n21775
g21712 and a[2] n21775_not ; n21776
g21713 and a[2]_not n21775 ; n21777
g21714 nor n21776 n21777 ; n21778
g21715 and n21767 n21778 ; n21779
g21716 and n21423 n21425_not ; n21780
g21717 nor n21426 n21780 ; n21781
g21718 and n21779_not n21781 ; n21782
g21719 nor n21767 n21778 ; n21783
g21720 nor n21782 n21783 ; n21784
g21721 and n11727 n12549 ; n21785
g21722 and n11055 n12555 ; n21786
g21723 and n11715 n12552 ; n21787
g21724 nor n21786 n21787 ; n21788
g21725 and n21785_not n21788 ; n21789
g21726 and n11057_not n21789 ; n21790
g21727 and n15764_not n21789 ; n21791
g21728 nor n21790 n21791 ; n21792
g21729 and a[2] n21792_not ; n21793
g21730 and a[2]_not n21792 ; n21794
g21731 nor n21793 n21794 ; n21795
g21732 and n21784 n21795 ; n21796
g21733 and n21330 n21427 ; n21797
g21734 nor n21428 n21797 ; n21798
g21735 and n21796_not n21798 ; n21799
g21736 nor n21784 n21795 ; n21800
g21737 nor n21799 n21800 ; n21801
g21738 and n21429 n21431_not ; n21802
g21739 and n21430_not n21802 ; n21803
g21740 nor n21433 n21803 ; n21804
g21741 and n21801_not n21804 ; n21805
g21742 and n21801 n21804_not ; n21806
g21743 and n11727 n12546 ; n21807
g21744 and n11055 n12552 ; n21808
g21745 and n11715 n12549 ; n21809
g21746 nor n21808 n21809 ; n21810
g21747 and n21807_not n21810 ; n21811
g21748 and n11057 n15356_not ; n21812
g21749 and n21811 n21812_not ; n21813
g21750 nor a[2] n21813 ; n21814
g21751 and a[2] n21813 ; n21815
g21752 nor n21814 n21815 ; n21816
g21753 nor n21806 n21816 ; n21817
g21754 nor n21805 n21817 ; n21818
g21755 and n21434 n21436_not ; n21819
g21756 and n21435_not n21819 ; n21820
g21757 nor n21438 n21820 ; n21821
g21758 and n21818_not n21821 ; n21822
g21759 and n21818 n21821_not ; n21823
g21760 and n11727 n12543 ; n21824
g21761 and n11055 n12549 ; n21825
g21762 and n11715 n12546 ; n21826
g21763 nor n21825 n21826 ; n21827
g21764 and n21824_not n21827 ; n21828
g21765 and n11057 n15724 ; n21829
g21766 and n21828 n21829_not ; n21830
g21767 nor a[2] n21830 ; n21831
g21768 and a[2] n21830 ; n21832
g21769 nor n21831 n21832 ; n21833
g21770 nor n21823 n21833 ; n21834
g21771 nor n21822 n21834 ; n21835
g21772 and n21653 n21835_not ; n21836
g21773 and n21653_not n21835 ; n21837
g21774 and n11727 n12540 ; n21838
g21775 and n11055 n12546 ; n21839
g21776 and n11715 n12543 ; n21840
g21777 nor n21839 n21840 ; n21841
g21778 and n21838_not n21841 ; n21842
g21779 and n11057 n15708_not ; n21843
g21780 and n21842 n21843_not ; n21844
g21781 nor a[2] n21844 ; n21845
g21782 and a[2] n21844 ; n21846
g21783 nor n21845 n21846 ; n21847
g21784 nor n21837 n21847 ; n21848
g21785 nor n21836 n21848 ; n21849
g21786 and n11727 n12537 ; n21850
g21787 and n11055 n12543 ; n21851
g21788 and n11715 n12540 ; n21852
g21789 nor n21851 n21852 ; n21853
g21790 and n21850_not n21853 ; n21854
g21791 and n11057_not n21854 ; n21855
g21792 and n15385 n21854 ; n21856
g21793 nor n21855 n21856 ; n21857
g21794 and a[2] n21857_not ; n21858
g21795 and a[2]_not n21857 ; n21859
g21796 nor n21858 n21859 ; n21860
g21797 and n21849 n21860 ; n21861
g21798 and n21271 n21443 ; n21862
g21799 nor n21444 n21862 ; n21863
g21800 and n21861_not n21863 ; n21864
g21801 nor n21849 n21860 ; n21865
g21802 nor n21864 n21865 ; n21866
g21803 and n11727 n12534 ; n21867
g21804 and n11055 n12540 ; n21868
g21805 and n11715 n12537 ; n21869
g21806 nor n21868 n21869 ; n21870
g21807 and n21867_not n21870 ; n21871
g21808 and n11057_not n21871 ; n21872
g21809 and n15096 n21871 ; n21873
g21810 nor n21872 n21873 ; n21874
g21811 and a[2] n21874_not ; n21875
g21812 and a[2]_not n21874 ; n21876
g21813 nor n21875 n21876 ; n21877
g21814 and n21866 n21877 ; n21878
g21815 and n21253 n21445 ; n21879
g21816 nor n21446 n21879 ; n21880
g21817 and n21878_not n21880 ; n21881
g21818 nor n21866 n21877 ; n21882
g21819 nor n21881 n21882 ; n21883
g21820 and n11727 n12531 ; n21884
g21821 and n11055 n12537 ; n21885
g21822 and n11715 n12534 ; n21886
g21823 nor n21885 n21886 ; n21887
g21824 and n21884_not n21887 ; n21888
g21825 and n11057_not n21888 ; n21889
g21826 and n15255_not n21888 ; n21890
g21827 nor n21889 n21890 ; n21891
g21828 and a[2] n21891_not ; n21892
g21829 and a[2]_not n21891 ; n21893
g21830 nor n21892 n21893 ; n21894
g21831 and n21883 n21894 ; n21895
g21832 and n21235 n21447 ; n21896
g21833 nor n21448 n21896 ; n21897
g21834 and n21895_not n21897 ; n21898
g21835 nor n21883 n21894 ; n21899
g21836 nor n21898 n21899 ; n21900
g21837 and n21449 n21451_not ; n21901
g21838 and n21450_not n21901 ; n21902
g21839 nor n21453 n21902 ; n21903
g21840 and n21900_not n21903 ; n21904
g21841 and n21900 n21903_not ; n21905
g21842 and n11727 n12528 ; n21906
g21843 and n11055 n12534 ; n21907
g21844 and n11715 n12531 ; n21908
g21845 nor n21907 n21908 ; n21909
g21846 and n21906_not n21909 ; n21910
g21847 and n11057 n15003_not ; n21911
g21848 and n21910 n21911_not ; n21912
g21849 nor a[2] n21912 ; n21913
g21850 and a[2] n21912 ; n21914
g21851 nor n21913 n21914 ; n21915
g21852 nor n21905 n21915 ; n21916
g21853 nor n21904 n21916 ; n21917
g21854 and n21454 n21456_not ; n21918
g21855 and n21455_not n21918 ; n21919
g21856 nor n21458 n21919 ; n21920
g21857 and n21917_not n21920 ; n21921
g21858 and n21917 n21920_not ; n21922
g21859 and n11727 n12525 ; n21923
g21860 and n11055 n12531 ; n21924
g21861 and n11715 n12528 ; n21925
g21862 nor n21924 n21925 ; n21926
g21863 and n21923_not n21926 ; n21927
g21864 and n11057 n14608 ; n21928
g21865 and n21927 n21928_not ; n21929
g21866 nor a[2] n21929 ; n21930
g21867 and a[2] n21929 ; n21931
g21868 nor n21930 n21931 ; n21932
g21869 nor n21922 n21932 ; n21933
g21870 nor n21921 n21933 ; n21934
g21871 and n21651 n21934_not ; n21935
g21872 and n21651_not n21934 ; n21936
g21873 and n11727 n12522 ; n21937
g21874 and n11055 n12528 ; n21938
g21875 and n11715 n12525 ; n21939
g21876 nor n21938 n21939 ; n21940
g21877 and n21937_not n21940 ; n21941
g21878 and n11057 n14837 ; n21942
g21879 and n21941 n21942_not ; n21943
g21880 nor a[2] n21943 ; n21944
g21881 and a[2] n21943 ; n21945
g21882 nor n21944 n21945 ; n21946
g21883 nor n21936 n21946 ; n21947
g21884 nor n21935 n21947 ; n21948
g21885 and n11727 n12519 ; n21949
g21886 and n11055 n12525 ; n21950
g21887 and n11715 n12522 ; n21951
g21888 nor n21950 n21951 ; n21952
g21889 and n21949_not n21952 ; n21953
g21890 and n11057_not n21953 ; n21954
g21891 and n14454_not n21953 ; n21955
g21892 nor n21954 n21955 ; n21956
g21893 and a[2] n21956_not ; n21957
g21894 and a[2]_not n21956 ; n21958
g21895 nor n21957 n21958 ; n21959
g21896 and n21948 n21959 ; n21960
g21897 and n21176 n21463 ; n21961
g21898 nor n21464 n21961 ; n21962
g21899 and n21960_not n21962 ; n21963
g21900 nor n21948 n21959 ; n21964
g21901 nor n21963 n21964 ; n21965
g21902 and n11727 n12516 ; n21966
g21903 and n11055 n12522 ; n21967
g21904 and n11715 n12519 ; n21968
g21905 nor n21967 n21968 ; n21969
g21906 and n21966_not n21969 ; n21970
g21907 and n11057_not n21970 ; n21971
g21908 and n14443 n21970 ; n21972
g21909 nor n21971 n21972 ; n21973
g21910 and a[2] n21973_not ; n21974
g21911 and a[2]_not n21973 ; n21975
g21912 nor n21974 n21975 ; n21976
g21913 and n21965 n21976 ; n21977
g21914 and n21158 n21465 ; n21978
g21915 nor n21466 n21978 ; n21979
g21916 and n21977_not n21979 ; n21980
g21917 nor n21965 n21976 ; n21981
g21918 nor n21980 n21981 ; n21982
g21919 and n11727 n12511 ; n21983
g21920 and n11055 n12519 ; n21984
g21921 and n11715 n12516 ; n21985
g21922 nor n21984 n21985 ; n21986
g21923 and n21983_not n21986 ; n21987
g21924 and n11057_not n21987 ; n21988
g21925 and n14233 n21987 ; n21989
g21926 nor n21988 n21989 ; n21990
g21927 and a[2] n21990_not ; n21991
g21928 and a[2]_not n21990 ; n21992
g21929 nor n21991 n21992 ; n21993
g21930 and n21982 n21993 ; n21994
g21931 and n21140 n21467 ; n21995
g21932 nor n21468 n21995 ; n21996
g21933 and n21994_not n21996 ; n21997
g21934 nor n21982 n21993 ; n21998
g21935 nor n21997 n21998 ; n21999
g21936 and n21469 n21471_not ; n22000
g21937 and n21470_not n22000 ; n22001
g21938 nor n21473 n22001 ; n22002
g21939 and n21999_not n22002 ; n22003
g21940 and n21999 n22002_not ; n22004
g21941 and n11727 n12513 ; n22005
g21942 and n11055 n12516 ; n22006
g21943 and n11715 n12511 ; n22007
g21944 nor n22006 n22007 ; n22008
g21945 and n22005_not n22008 ; n22009
g21946 and n11057 n14177 ; n22010
g21947 and n22009 n22010_not ; n22011
g21948 nor a[2] n22011 ; n22012
g21949 and a[2] n22011 ; n22013
g21950 nor n22012 n22013 ; n22014
g21951 nor n22004 n22014 ; n22015
g21952 nor n22003 n22015 ; n22016
g21953 and n21474 n21476_not ; n22017
g21954 and n21475_not n22017 ; n22018
g21955 nor n21478 n22018 ; n22019
g21956 and n22016_not n22019 ; n22020
g21957 and n22016 n22019_not ; n22021
g21958 and n11727 n12508 ; n22022
g21959 and n11055 n12511 ; n22023
g21960 and n11715 n12513 ; n22024
g21961 nor n22023 n22024 ; n22025
g21962 and n22022_not n22025 ; n22026
g21963 and n11057 n13863 ; n22027
g21964 and n22026 n22027_not ; n22028
g21965 nor a[2] n22028 ; n22029
g21966 and a[2] n22028 ; n22030
g21967 nor n22029 n22030 ; n22031
g21968 nor n22021 n22031 ; n22032
g21969 nor n22020 n22032 ; n22033
g21970 and n21649 n22033_not ; n22034
g21971 and n21649_not n22033 ; n22035
g21972 and n11727 n12505 ; n22036
g21973 and n11055 n12513 ; n22037
g21974 and n11715 n12508 ; n22038
g21975 nor n22037 n22038 ; n22039
g21976 and n22036_not n22039 ; n22040
g21977 and n11057 n14051_not ; n22041
g21978 and n22040 n22041_not ; n22042
g21979 nor a[2] n22042 ; n22043
g21980 and a[2] n22042 ; n22044
g21981 nor n22043 n22044 ; n22045
g21982 nor n22035 n22045 ; n22046
g21983 nor n22034 n22046 ; n22047
g21984 and n11727 n12370 ; n22048
g21985 and n11055 n12508 ; n22049
g21986 and n11715 n12505 ; n22050
g21987 nor n22049 n22050 ; n22051
g21988 and n22048_not n22051 ; n22052
g21989 and n11057_not n22052 ; n22053
g21990 and n13748 n22052 ; n22054
g21991 nor n22053 n22054 ; n22055
g21992 and a[2] n22055_not ; n22056
g21993 and a[2]_not n22055 ; n22057
g21994 nor n22056 n22057 ; n22058
g21995 and n22047 n22058 ; n22059
g21996 and n21081 n21483 ; n22060
g21997 nor n21484 n22060 ; n22061
g21998 and n22059_not n22061 ; n22062
g21999 nor n22047 n22058 ; n22063
g22000 nor n22062 n22063 ; n22064
g22001 and n11727 n12502 ; n22065
g22002 and n11055 n12505 ; n22066
g22003 and n11715 n12370 ; n22067
g22004 nor n22066 n22067 ; n22068
g22005 and n22065_not n22068 ; n22069
g22006 and n11057_not n22069 ; n22070
g22007 and n13736 n22069 ; n22071
g22008 nor n22070 n22071 ; n22072
g22009 and a[2] n22072_not ; n22073
g22010 and a[2]_not n22072 ; n22074
g22011 nor n22073 n22074 ; n22075
g22012 and n22064 n22075 ; n22076
g22013 and n21063 n21485 ; n22077
g22014 nor n21486 n22077 ; n22078
g22015 and n22076_not n22078 ; n22079
g22016 nor n22064 n22075 ; n22080
g22017 nor n22079 n22080 ; n22081
g22018 and n11727 n12769 ; n22082
g22019 and n11055 n12370 ; n22083
g22020 and n11715 n12502 ; n22084
g22021 nor n22083 n22084 ; n22085
g22022 and n22082_not n22085 ; n22086
g22023 and n11057_not n22086 ; n22087
g22024 and n12999_not n22086 ; n22088
g22025 nor n22087 n22088 ; n22089
g22026 and a[2] n22089_not ; n22090
g22027 and a[2]_not n22089 ; n22091
g22028 nor n22090 n22091 ; n22092
g22029 and n22081 n22092 ; n22093
g22030 and n21045 n21487 ; n22094
g22031 nor n21488 n22094 ; n22095
g22032 and n22093_not n22095 ; n22096
g22033 nor n22081 n22092 ; n22097
g22034 nor n22096 n22097 ; n22098
g22035 and n21489 n21491_not ; n22099
g22036 and n21490_not n22099 ; n22100
g22037 nor n21493 n22100 ; n22101
g22038 and n22098_not n22101 ; n22102
g22039 and n22098 n22101_not ; n22103
g22040 and n11727 n12889 ; n22104
g22041 and n11055 n12502 ; n22105
g22042 and n11715 n12769 ; n22106
g22043 nor n22105 n22106 ; n22107
g22044 and n22104_not n22107 ; n22108
g22045 and n11057 n12895 ; n22109
g22046 and n22108 n22109_not ; n22110
g22047 nor a[2] n22110 ; n22111
g22048 and a[2] n22110 ; n22112
g22049 nor n22111 n22112 ; n22113
g22050 nor n22103 n22113 ; n22114
g22051 nor n22102 n22114 ; n22115
g22052 and n21647 n22115_not ; n22116
g22053 and n21647_not n22115 ; n22117
g22054 and n11727 n13491 ; n22118
g22055 and n11055 n12769 ; n22119
g22056 and n11715 n12889 ; n22120
g22057 nor n22119 n22120 ; n22121
g22058 and n22118_not n22121 ; n22122
g22059 and n11057 n13503_not ; n22123
g22060 and n22122 n22123_not ; n22124
g22061 nor a[2] n22124 ; n22125
g22062 and a[2] n22124 ; n22126
g22063 nor n22125 n22126 ; n22127
g22064 nor n22117 n22127 ; n22128
g22065 nor n22116 n22128 ; n22129
g22066 and n21633 n21645_not ; n22130
g22067 nor n21644 n21645 ; n22131
g22068 nor n22130 n22131 ; n22132
g22069 nor n22129 n22132 ; n22133
g22070 nor n21645 n22133 ; n22134
g22071 and n21619_not n21630 ; n22135
g22072 nor n21631 n22135 ; n22136
g22073 and n22134_not n22136 ; n22137
g22074 nor n21631 n22137 ; n22138
g22075 and n21605_not n21616 ; n22139
g22076 nor n21617 n22139 ; n22140
g22077 and n22138_not n22140 ; n22141
g22078 nor n21617 n22141 ; n22142
g22079 and n21591_not n21602 ; n22143
g22080 nor n21603 n22143 ; n22144
g22081 and n22142_not n22144 ; n22145
g22082 nor n21603 n22145 ; n22146
g22083 and n21577_not n21588 ; n22147
g22084 nor n21589 n22147 ; n22148
g22085 and n22146_not n22148 ; n22149
g22086 nor n21589 n22149 ; n22150
g22087 and n21563_not n21574 ; n22151
g22088 nor n21575 n22151 ; n22152
g22089 and n22150_not n22152 ; n22153
g22090 nor n21575 n22153 ; n22154
g22091 and n21549_not n21560 ; n22155
g22092 nor n21561 n22155 ; n22156
g22093 and n22154_not n22156 ; n22157
g22094 nor n21561 n22157 ; n22158
g22095 and n21535_not n21546 ; n22159
g22096 nor n21547 n22159 ; n22160
g22097 and n22158_not n22160 ; n22161
g22098 nor n21547 n22161 ; n22162
g22099 and n21521_not n21532 ; n22163
g22100 nor n21533 n22163 ; n22164
g22101 and n22162_not n22164 ; n22165
g22102 nor n21533 n22165 ; n22166
g22103 and n21519 n22166_not ; n22167
g22104 nor n21517 n22167 ; n22168
g22105 and n20835 n22168_not ; n22169
g22106 nor n20833 n22169 ; n22170
g22107 and n20800 n22170_not ; n22171
g22108 nor n20798 n22171 ; n22172
g22109 and n20145 n22172_not ; n22173
g22110 nor n20143 n22173 ; n22174
g22111 and n19516 n19518_not ; n22175
g22112 nor n19519 n22175 ; n22176
g22113 and n22174_not n22176 ; n22177
g22114 nor n19519 n22177 ; n22178
g22115 nor n18946 n22178 ; n22179
g22116 nor n18943 n22179 ; n22180
g22117 and n18396 n22180_not ; n22181
g22118 nor n18394 n22181 ; n22182
g22119 and n17892 n17894_not ; n22183
g22120 nor n17895 n22183 ; n22184
g22121 and n22182_not n22184 ; n22185
g22122 nor n17895 n22185 ; n22186
g22123 nor n17428 n22186 ; n22187
g22124 nor n17425 n22187 ; n22188
g22125 and n17001 n22188_not ; n22189
g22126 nor n16999 n22189 ; n22190
g22127 and n16604 n16606_not ; n22191
g22128 nor n16607 n22191 ; n22192
g22129 and n22190_not n22192 ; n22193
g22130 nor n16607 n22193 ; n22194
g22131 nor n16443 n22194 ; n22195
g22132 nor n16440 n22195 ; n22196
g22133 and n16272 n22196_not ; n22197
g22134 nor n16270 n22197 ; n22198
g22135 and n15650 n15652_not ; n22199
g22136 nor n15653 n22199 ; n22200
g22137 and n22198_not n22200 ; n22201
g22138 nor n15653 n22201 ; n22202
g22139 nor n15508 n22202 ; n22203
g22140 nor n15505 n22203 ; n22204
g22141 and n15203 n22204_not ; n22205
g22142 nor n15201 n22205 ; n22206
g22143 and n14950 n14952_not ; n22207
g22144 nor n14953 n22207 ; n22208
g22145 and n22206_not n22208 ; n22209
g22146 nor n14953 n22209 ; n22210
g22147 nor n14809 n22210 ; n22211
g22148 nor n14806 n22211 ; n22212
g22149 and n14696 n22212_not ; n22213
g22150 nor n14694 n22213 ; n22214
g22151 and n14321 n14323_not ; n22215
g22152 nor n14324 n22215 ; n22216
g22153 and n22214_not n22216 ; n22217
g22154 nor n14324 n22217 ; n22218
g22155 nor n14154 n22218 ; n22219
g22156 nor n14151 n22219 ; n22220
g22157 and n14039 n22220_not ; n22221
g22158 nor n14037 n22221 ; n22222
g22159 nor n13957 n13960 ; n22223
g22160 nor n13621 n13661 ; n22224
g22161 and n3884 n13941 ; n22225
g22162 and n3967 n13633 ; n22226
g22163 and n4046 n13627_not ; n22227
g22164 nor n22226 n22227 ; n22228
g22165 and n22225_not n22228 ; n22229
g22166 and n4050 n14136 ; n22230
g22167 and n22229 n22230_not ; n22231
g22168 and a[26] n22231_not ; n22232
g22169 and a[26] n22232_not ; n22233
g22170 nor n22231 n22232 ; n22234
g22171 nor n22233 n22234 ; n22235
g22172 nor n22224 n22235 ; n22236
g22173 nor n22224 n22236 ; n22237
g22174 nor n22235 n22236 ; n22238
g22175 nor n22237 n22238 ; n22239
g22176 and n75 n13909_not ; n22240
g22177 and n3020 n13521 ; n22241
g22178 and n3023 n13491 ; n22242
g22179 and n3028 n13518 ; n22243
g22180 nor n22242 n22243 ; n22244
g22181 and n22241_not n22244 ; n22245
g22182 and n22240_not n22245 ; n22246
g22183 and n4533_not n13938 ; n22247
g22184 and n4536_not n22247 ; n22248
g22185 nor n13438 n22248 ; n22249
g22186 and a[23] n22249_not ; n22250
g22187 and a[23]_not n22249 ; n22251
g22188 nor n22250 n22251 ; n22252
g22189 and n303 n3042 ; n22253
g22190 and n6567 n22253 ; n22254
g22191 and n4827 n22254 ; n22255
g22192 and n16031 n22255 ; n22256
g22193 and n13787 n22256 ; n22257
g22194 and n14534 n22257 ; n22258
g22195 and n774 n22258 ; n22259
g22196 and n471 n22259 ; n22260
g22197 and n3733 n22260 ; n22261
g22198 and n1269 n22261 ; n22262
g22199 and n847_not n22262 ; n22263
g22200 and n367_not n22263 ; n22264
g22201 and n226_not n22264 ; n22265
g22202 and n306_not n22265 ; n22266
g22203 and n158_not n22266 ; n22267
g22204 and n270_not n22267 ; n22268
g22205 and n13574 n22268 ; n22269
g22206 nor n13574 n22268 ; n22270
g22207 nor n22269 n22270 ; n22271
g22208 and n22252 n22271 ; n22272
g22209 nor n22252 n22271 ; n22273
g22210 nor n22272 n22273 ; n22274
g22211 and n13580_not n22274 ; n22275
g22212 and n13580 n22274_not ; n22276
g22213 nor n22275 n22276 ; n22277
g22214 and n22246_not n22277 ; n22278
g22215 and n22277 n22278_not ; n22279
g22216 nor n22246 n22278 ; n22280
g22217 nor n22279 n22280 ; n22281
g22218 nor n13592 n13618 ; n22282
g22219 and n22281 n22282 ; n22283
g22220 nor n22281 n22282 ; n22284
g22221 nor n22283 n22284 ; n22285
g22222 and n3457 n13630 ; n22286
g22223 and n3542 n13515 ; n22287
g22224 and n3606 n13597 ; n22288
g22225 nor n22287 n22288 ; n22289
g22226 and n22286_not n22289 ; n22290
g22227 and n3368 n13976 ; n22291
g22228 and n22290 n22291_not ; n22292
g22229 and a[29] n22292_not ; n22293
g22230 and a[29] n22293_not ; n22294
g22231 nor n22292 n22293 ; n22295
g22232 nor n22294 n22295 ; n22296
g22233 and n22285 n22296_not ; n22297
g22234 and n22285 n22297_not ; n22298
g22235 nor n22296 n22297 ; n22299
g22236 nor n22298 n22299 ; n22300
g22237 and n22239_not n22300 ; n22301
g22238 and n22239 n22300_not ; n22302
g22239 nor n22301 n22302 ; n22303
g22240 nor n22223 n22303 ; n22304
g22241 and n22223 n22303 ; n22305
g22242 nor n22304 n22305 ; n22306
g22243 and n22222_not n22306 ; n22307
g22244 and n22222 n22306_not ; n22308
g22245 nor n22307 n22308 ; n22309
g22246 and n71 n22309 ; n22310
g22247 and n14154 n22218 ; n22311
g22248 nor n22219 n22311 ; n22312
g22249 and n9867 n22312 ; n22313
g22250 and n14039_not n22220 ; n22314
g22251 nor n22221 n22314 ; n22315
g22252 and n10434 n22315 ; n22316
g22253 nor n22313 n22316 ; n22317
g22254 and n22310_not n22317 ; n22318
g22255 and n22214 n22216_not ; n22319
g22256 nor n22217 n22319 ; n22320
g22257 and n22312 n22320 ; n22321
g22258 and n14696_not n22212 ; n22322
g22259 nor n22213 n22322 ; n22323
g22260 and n22320 n22323 ; n22324
g22261 and n14809 n22210 ; n22325
g22262 nor n22211 n22325 ; n22326
g22263 and n22323 n22326 ; n22327
g22264 and n22206 n22208_not ; n22328
g22265 nor n22209 n22328 ; n22329
g22266 and n22326 n22329 ; n22330
g22267 and n15203_not n22204 ; n22331
g22268 nor n22205 n22331 ; n22332
g22269 and n22329 n22332 ; n22333
g22270 and n15508 n22202 ; n22334
g22271 nor n22203 n22334 ; n22335
g22272 and n22332 n22335 ; n22336
g22273 and n22198 n22200_not ; n22337
g22274 nor n22201 n22337 ; n22338
g22275 and n22335 n22338 ; n22339
g22276 and n16272_not n22196 ; n22340
g22277 nor n22197 n22340 ; n22341
g22278 and n22338 n22341 ; n22342
g22279 and n16443 n22194 ; n22343
g22280 nor n22195 n22343 ; n22344
g22281 and n22341 n22344 ; n22345
g22282 and n22190 n22192_not ; n22346
g22283 nor n22193 n22346 ; n22347
g22284 and n22344 n22347 ; n22348
g22285 and n17001_not n22188 ; n22349
g22286 nor n22189 n22349 ; n22350
g22287 and n22347 n22350 ; n22351
g22288 and n17428 n22186 ; n22352
g22289 nor n22187 n22352 ; n22353
g22290 and n22350 n22353 ; n22354
g22291 and n22182 n22184_not ; n22355
g22292 nor n22185 n22355 ; n22356
g22293 and n22353 n22356 ; n22357
g22294 and n18396_not n22180 ; n22358
g22295 nor n22181 n22358 ; n22359
g22296 and n22356 n22359 ; n22360
g22297 and n18946 n22178 ; n22361
g22298 nor n22179 n22361 ; n22362
g22299 and n22359 n22362 ; n22363
g22300 and n22174 n22176_not ; n22364
g22301 nor n22177 n22364 ; n22365
g22302 and n22362 n22365 ; n22366
g22303 and n20145_not n22172 ; n22367
g22304 nor n22173 n22367 ; n22368
g22305 and n22365 n22368 ; n22369
g22306 and n20800_not n22170 ; n22370
g22307 nor n22171 n22370 ; n22371
g22308 and n22368 n22371 ; n22372
g22309 and n20835_not n22168 ; n22373
g22310 nor n22169 n22373 ; n22374
g22311 and n22371 n22374 ; n22375
g22312 and n21519_not n22166 ; n22376
g22313 nor n22167 n22376 ; n22377
g22314 and n22374 n22377 ; n22378
g22315 and n22162 n22164_not ; n22379
g22316 nor n22165 n22379 ; n22380
g22317 and n22377 n22380 ; n22381
g22318 nor n22377 n22380 ; n22382
g22319 and n22158 n22160_not ; n22383
g22320 nor n22161 n22383 ; n22384
g22321 and n22380 n22384 ; n22385
g22322 and n22154 n22156_not ; n22386
g22323 nor n22157 n22386 ; n22387
g22324 and n22384 n22387 ; n22388
g22325 and n22150 n22152_not ; n22389
g22326 nor n22153 n22389 ; n22390
g22327 and n22387 n22390 ; n22391
g22328 and n22146 n22148_not ; n22392
g22329 nor n22149 n22392 ; n22393
g22330 and n22390 n22393 ; n22394
g22331 and n22142 n22144_not ; n22395
g22332 nor n22145 n22395 ; n22396
g22333 and n22393 n22396 ; n22397
g22334 and n22138 n22140_not ; n22398
g22335 nor n22141 n22398 ; n22399
g22336 and n22396 n22399 ; n22400
g22337 and n22134 n22136_not ; n22401
g22338 nor n22137 n22401 ; n22402
g22339 and n22399 n22402 ; n22403
g22340 nor n22129 n22133 ; n22404
g22341 nor n22132 n22133 ; n22405
g22342 nor n22404 n22405 ; n22406
g22343 and n22402 n22406_not ; n22407
g22344 and n22399_not n22407 ; n22408
g22345 nor n22403 n22408 ; n22409
g22346 nor n22396 n22399 ; n22410
g22347 nor n22400 n22410 ; n22411
g22348 and n22409_not n22411 ; n22412
g22349 nor n22400 n22412 ; n22413
g22350 nor n22393 n22396 ; n22414
g22351 nor n22397 n22414 ; n22415
g22352 and n22413_not n22415 ; n22416
g22353 nor n22397 n22416 ; n22417
g22354 nor n22390 n22393 ; n22418
g22355 nor n22394 n22418 ; n22419
g22356 and n22417_not n22419 ; n22420
g22357 nor n22394 n22420 ; n22421
g22358 nor n22387 n22390 ; n22422
g22359 nor n22391 n22422 ; n22423
g22360 and n22421_not n22423 ; n22424
g22361 nor n22391 n22424 ; n22425
g22362 nor n22384 n22387 ; n22426
g22363 nor n22388 n22426 ; n22427
g22364 and n22425_not n22427 ; n22428
g22365 nor n22388 n22428 ; n22429
g22366 nor n22380 n22384 ; n22430
g22367 nor n22385 n22430 ; n22431
g22368 and n22429_not n22431 ; n22432
g22369 nor n22385 n22432 ; n22433
g22370 nor n22381 n22433 ; n22434
g22371 and n22382_not n22434 ; n22435
g22372 nor n22381 n22435 ; n22436
g22373 nor n22374 n22377 ; n22437
g22374 nor n22378 n22437 ; n22438
g22375 and n22436_not n22438 ; n22439
g22376 nor n22378 n22439 ; n22440
g22377 nor n22371 n22374 ; n22441
g22378 nor n22375 n22441 ; n22442
g22379 and n22440_not n22442 ; n22443
g22380 nor n22375 n22443 ; n22444
g22381 nor n22368 n22371 ; n22445
g22382 nor n22372 n22445 ; n22446
g22383 and n22444_not n22446 ; n22447
g22384 nor n22372 n22447 ; n22448
g22385 nor n22365 n22368 ; n22449
g22386 nor n22448 n22449 ; n22450
g22387 and n22369_not n22450 ; n22451
g22388 nor n22369 n22451 ; n22452
g22389 nor n22362 n22365 ; n22453
g22390 nor n22452 n22453 ; n22454
g22391 and n22366_not n22454 ; n22455
g22392 nor n22366 n22455 ; n22456
g22393 nor n22359 n22362 ; n22457
g22394 nor n22363 n22457 ; n22458
g22395 and n22456_not n22458 ; n22459
g22396 nor n22363 n22459 ; n22460
g22397 nor n22356 n22359 ; n22461
g22398 nor n22460 n22461 ; n22462
g22399 and n22360_not n22462 ; n22463
g22400 nor n22360 n22463 ; n22464
g22401 nor n22353 n22356 ; n22465
g22402 nor n22464 n22465 ; n22466
g22403 and n22357_not n22466 ; n22467
g22404 nor n22357 n22467 ; n22468
g22405 nor n22350 n22353 ; n22469
g22406 nor n22354 n22469 ; n22470
g22407 and n22468_not n22470 ; n22471
g22408 nor n22354 n22471 ; n22472
g22409 nor n22347 n22350 ; n22473
g22410 nor n22472 n22473 ; n22474
g22411 and n22351_not n22474 ; n22475
g22412 nor n22351 n22475 ; n22476
g22413 nor n22344 n22347 ; n22477
g22414 nor n22476 n22477 ; n22478
g22415 and n22348_not n22478 ; n22479
g22416 nor n22348 n22479 ; n22480
g22417 nor n22341 n22344 ; n22481
g22418 nor n22345 n22481 ; n22482
g22419 and n22480_not n22482 ; n22483
g22420 nor n22345 n22483 ; n22484
g22421 nor n22338 n22341 ; n22485
g22422 nor n22484 n22485 ; n22486
g22423 and n22342_not n22486 ; n22487
g22424 nor n22342 n22487 ; n22488
g22425 nor n22335 n22338 ; n22489
g22426 nor n22488 n22489 ; n22490
g22427 and n22339_not n22490 ; n22491
g22428 nor n22339 n22491 ; n22492
g22429 nor n22332 n22335 ; n22493
g22430 nor n22336 n22493 ; n22494
g22431 and n22492_not n22494 ; n22495
g22432 nor n22336 n22495 ; n22496
g22433 nor n22329 n22332 ; n22497
g22434 nor n22496 n22497 ; n22498
g22435 and n22333_not n22498 ; n22499
g22436 nor n22333 n22499 ; n22500
g22437 nor n22326 n22329 ; n22501
g22438 nor n22500 n22501 ; n22502
g22439 and n22330_not n22502 ; n22503
g22440 nor n22330 n22503 ; n22504
g22441 nor n22323 n22326 ; n22505
g22442 nor n22327 n22505 ; n22506
g22443 and n22504_not n22506 ; n22507
g22444 nor n22327 n22507 ; n22508
g22445 nor n22320 n22323 ; n22509
g22446 nor n22508 n22509 ; n22510
g22447 and n22324_not n22510 ; n22511
g22448 nor n22324 n22511 ; n22512
g22449 nor n22312 n22320 ; n22513
g22450 nor n22512 n22513 ; n22514
g22451 and n22321_not n22514 ; n22515
g22452 nor n22321 n22515 ; n22516
g22453 nor n22312 n22315 ; n22517
g22454 and n22312 n22315 ; n22518
g22455 nor n22517 n22518 ; n22519
g22456 and n22516_not n22519 ; n22520
g22457 nor n22518 n22520 ; n22521
g22458 and n22309 n22315 ; n22522
g22459 nor n22309 n22315 ; n22523
g22460 nor n22521 n22523 ; n22524
g22461 and n22522_not n22524 ; n22525
g22462 nor n22521 n22525 ; n22526
g22463 nor n22522 n22525 ; n22527
g22464 and n22523_not n22527 ; n22528
g22465 nor n22526 n22528 ; n22529
g22466 and n9870 n22529_not ; n22530
g22467 and n22318 n22530_not ; n22531
g22468 and a[5] n22531_not ; n22532
g22469 nor n22531 n22532 ; n22533
g22470 and a[5] n22532_not ; n22534
g22471 nor n22533 n22534 ; n22535
g22472 and n7983 n22332 ; n22536
g22473 and n7291 n22338 ; n22537
g22474 and n7632 n22335 ; n22538
g22475 nor n22537 n22538 ; n22539
g22476 and n22536_not n22539 ; n22540
g22477 and n22492 n22494_not ; n22541
g22478 nor n22495 n22541 ; n22542
g22479 and n7294 n22542 ; n22543
g22480 and n22540 n22543_not ; n22544
g22481 and a[11] n22544_not ; n22545
g22482 nor n22544 n22545 ; n22546
g22483 and a[11] n22545_not ; n22547
g22484 nor n22546 n22547 ; n22548
g22485 and n6233 n22353 ; n22549
g22486 and n5663 n22359 ; n22550
g22487 and n5939 n22356 ; n22551
g22488 nor n22550 n22551 ; n22552
g22489 and n22549_not n22552 ; n22553
g22490 nor n22464 n22467 ; n22554
g22491 and n22465_not n22468 ; n22555
g22492 nor n22554 n22555 ; n22556
g22493 and n5666 n22556_not ; n22557
g22494 and n22553 n22557_not ; n22558
g22495 and a[17] n22558_not ; n22559
g22496 nor n22558 n22559 ; n22560
g22497 and a[17] n22559_not ; n22561
g22498 nor n22560 n22561 ; n22562
g22499 and n4694 n22374 ; n22563
g22500 and n4533 n22380 ; n22564
g22501 and n4604 n22377 ; n22565
g22502 nor n22564 n22565 ; n22566
g22503 and n22563_not n22566 ; n22567
g22504 and n22436 n22438_not ; n22568
g22505 nor n22439 n22568 ; n22569
g22506 and n4536 n22569 ; n22570
g22507 and n22567 n22570_not ; n22571
g22508 and a[23] n22571_not ; n22572
g22509 nor n22571 n22572 ; n22573
g22510 and a[23] n22572_not ; n22574
g22511 nor n22573 n22574 ; n22575
g22512 and n3884 n22387 ; n22576
g22513 and n3967 n22393 ; n22577
g22514 and n4046 n22390 ; n22578
g22515 nor n22577 n22578 ; n22579
g22516 and n22576_not n22579 ; n22580
g22517 and n22421 n22423_not ; n22581
g22518 nor n22424 n22581 ; n22582
g22519 and n4050 n22582 ; n22583
g22520 and n22580 n22583_not ; n22584
g22521 and a[26] n22584_not ; n22585
g22522 nor n22584 n22585 ; n22586
g22523 and a[26] n22585_not ; n22587
g22524 nor n22586 n22587 ; n22588
g22525 and n3457 n22396 ; n22589
g22526 and n3542 n22402 ; n22590
g22527 and n3606 n22399 ; n22591
g22528 nor n22590 n22591 ; n22592
g22529 and n22589_not n22592 ; n22593
g22530 and n22409 n22411_not ; n22594
g22531 nor n22412 n22594 ; n22595
g22532 and n3368 n22595 ; n22596
g22533 and n22593 n22596_not ; n22597
g22534 and a[29] n22597_not ; n22598
g22535 nor n22597 n22598 ; n22599
g22536 and a[29] n22598_not ; n22600
g22537 nor n22599 n22600 ; n22601
g22538 nor n3367 n22406 ; n22602
g22539 and a[29] n22602_not ; n22603
g22540 and n3606 n22406_not ; n22604
g22541 and n3457 n22402 ; n22605
g22542 nor n22604 n22605 ; n22606
g22543 and n22402 n22406 ; n22607
g22544 nor n22402 n22406 ; n22608
g22545 nor n22607 n22608 ; n22609
g22546 and n3368 n22609_not ; n22610
g22547 and n22606 n22610_not ; n22611
g22548 and a[29] n22611_not ; n22612
g22549 and a[29] n22612_not ; n22613
g22550 nor n22611 n22612 ; n22614
g22551 nor n22613 n22614 ; n22615
g22552 and n22603 n22615_not ; n22616
g22553 and n3457 n22399 ; n22617
g22554 and n3542 n22406_not ; n22618
g22555 and n3606 n22402 ; n22619
g22556 nor n22618 n22619 ; n22620
g22557 and n22617_not n22620 ; n22621
g22558 and n3368_not n22621 ; n22622
g22559 and n22399_not n22607 ; n22623
g22560 and n22399 n22607_not ; n22624
g22561 nor n22623 n22624 ; n22625
g22562 and n22621 n22625 ; n22626
g22563 nor n22622 n22626 ; n22627
g22564 and a[29] n22627_not ; n22628
g22565 and a[29]_not n22627 ; n22629
g22566 nor n22628 n22629 ; n22630
g22567 and n22616 n22630_not ; n22631
g22568 nor n7479 n22406 ; n22632
g22569 and n22631 n22632_not ; n22633
g22570 and n22631_not n22632 ; n22634
g22571 nor n22633 n22634 ; n22635
g22572 nor n22601 n22635 ; n22636
g22573 and n22601 n22635 ; n22637
g22574 nor n22636 n22637 ; n22638
g22575 and n22588_not n22638 ; n22639
g22576 nor n22588 n22639 ; n22640
g22577 and n22638 n22639_not ; n22641
g22578 nor n22640 n22641 ; n22642
g22579 and n3884 n22390 ; n22643
g22580 and n3967 n22396 ; n22644
g22581 and n4046 n22393 ; n22645
g22582 nor n22644 n22645 ; n22646
g22583 and n22643_not n22646 ; n22647
g22584 and n22417 n22419_not ; n22648
g22585 nor n22420 n22648 ; n22649
g22586 and n4050 n22649 ; n22650
g22587 and n22647 n22650_not ; n22651
g22588 and a[26] n22651_not ; n22652
g22589 nor n22651 n22652 ; n22653
g22590 and a[26] n22652_not ; n22654
g22591 nor n22653 n22654 ; n22655
g22592 and n22616_not n22630 ; n22656
g22593 nor n22631 n22656 ; n22657
g22594 and n22655_not n22657 ; n22658
g22595 nor n22655 n22658 ; n22659
g22596 and n22657 n22658_not ; n22660
g22597 nor n22659 n22660 ; n22661
g22598 and n22603_not n22615 ; n22662
g22599 nor n22616 n22662 ; n22663
g22600 and n3884 n22393 ; n22664
g22601 and n3967 n22399 ; n22665
g22602 and n4046 n22396 ; n22666
g22603 nor n22665 n22666 ; n22667
g22604 and n22664_not n22667 ; n22668
g22605 and n4050_not n22668 ; n22669
g22606 and n22413 n22415_not ; n22670
g22607 nor n22416 n22670 ; n22671
g22608 and n22668 n22671_not ; n22672
g22609 nor n22669 n22672 ; n22673
g22610 and a[26] n22673_not ; n22674
g22611 and a[26]_not n22673 ; n22675
g22612 nor n22674 n22675 ; n22676
g22613 and n22663 n22676_not ; n22677
g22614 nor n3880 n22406 ; n22678
g22615 and a[26] n22678_not ; n22679
g22616 and n4046 n22406_not ; n22680
g22617 and n3884 n22402 ; n22681
g22618 nor n22680 n22681 ; n22682
g22619 and n4050 n22609_not ; n22683
g22620 and n22682 n22683_not ; n22684
g22621 and a[26] n22684_not ; n22685
g22622 and a[26] n22685_not ; n22686
g22623 nor n22684 n22685 ; n22687
g22624 nor n22686 n22687 ; n22688
g22625 and n22679 n22688_not ; n22689
g22626 and n3884 n22399 ; n22690
g22627 and n3967 n22406_not ; n22691
g22628 and n4046 n22402 ; n22692
g22629 nor n22691 n22692 ; n22693
g22630 and n22690_not n22693 ; n22694
g22631 and n4050_not n22694 ; n22695
g22632 and n22625 n22694 ; n22696
g22633 nor n22695 n22696 ; n22697
g22634 and a[26] n22697_not ; n22698
g22635 and a[26]_not n22697 ; n22699
g22636 nor n22698 n22699 ; n22700
g22637 and n22689 n22700_not ; n22701
g22638 and n22602 n22701 ; n22702
g22639 and n22701 n22702_not ; n22703
g22640 and n22602 n22702_not ; n22704
g22641 nor n22703 n22704 ; n22705
g22642 and n3884 n22396 ; n22706
g22643 and n3967 n22402 ; n22707
g22644 and n4046 n22399 ; n22708
g22645 nor n22707 n22708 ; n22709
g22646 and n22706_not n22709 ; n22710
g22647 and n4050 n22595 ; n22711
g22648 and n22710 n22711_not ; n22712
g22649 and a[26] n22712_not ; n22713
g22650 and a[26] n22713_not ; n22714
g22651 nor n22712 n22713 ; n22715
g22652 nor n22714 n22715 ; n22716
g22653 nor n22705 n22716 ; n22717
g22654 nor n22702 n22717 ; n22718
g22655 and n22663_not n22676 ; n22719
g22656 nor n22677 n22719 ; n22720
g22657 and n22718_not n22720 ; n22721
g22658 nor n22677 n22721 ; n22722
g22659 nor n22661 n22722 ; n22723
g22660 nor n22658 n22723 ; n22724
g22661 nor n22642 n22724 ; n22725
g22662 nor n22639 n22725 ; n22726
g22663 and n3457 n22393 ; n22727
g22664 and n3542 n22399 ; n22728
g22665 and n3606 n22396 ; n22729
g22666 nor n22728 n22729 ; n22730
g22667 and n22727_not n22730 ; n22731
g22668 and n3368 n22671 ; n22732
g22669 and n22731 n22732_not ; n22733
g22670 and a[29] n22733_not ; n22734
g22671 nor n22733 n22734 ; n22735
g22672 and a[29] n22734_not ; n22736
g22673 nor n22735 n22736 ; n22737
g22674 and n437 n2091 ; n22738
g22675 and n885 n22738 ; n22739
g22676 and n108 n22739 ; n22740
g22677 and n1367 n22740 ; n22741
g22678 and n462_not n22741 ; n22742
g22679 and n149_not n22742 ; n22743
g22680 and n228_not n22743 ; n22744
g22681 and n416_not n22744 ; n22745
g22682 and n980_not n22745 ; n22746
g22683 and n791_not n22746 ; n22747
g22684 and n712_not n22747 ; n22748
g22685 and n3206 n3858 ; n22749
g22686 and n2809 n22749 ; n22750
g22687 and n4104 n22750 ; n22751
g22688 and n14189 n22751 ; n22752
g22689 and n804 n22752 ; n22753
g22690 and n3163 n22753 ; n22754
g22691 and n2276 n22754 ; n22755
g22692 and n634 n22755 ; n22756
g22693 and n418 n22756 ; n22757
g22694 and n538 n22757 ; n22758
g22695 and n490_not n22758 ; n22759
g22696 and n589_not n22759 ; n22760
g22697 and n163_not n22760 ; n22761
g22698 and n451_not n22761 ; n22762
g22699 and n735 n2075 ; n22763
g22700 and n1044 n22763 ; n22764
g22701 and n15956 n22764 ; n22765
g22702 and n22762 n22765 ; n22766
g22703 and n22748 n22766 ; n22767
g22704 and n15867 n22767 ; n22768
g22705 and n1161 n22768 ; n22769
g22706 and n1269 n22769 ; n22770
g22707 and n1180 n22770 ; n22771
g22708 and n810 n22771 ; n22772
g22709 and n1128 n22772 ; n22773
g22710 and n341 n22773 ; n22774
g22711 and n397_not n22774 ; n22775
g22712 and n189_not n22775 ; n22776
g22713 and n331_not n22776 ; n22777
g22714 and n144_not n22777 ; n22778
g22715 and n366_not n22778 ; n22779
g22716 and n3020 n22402 ; n22780
g22717 and n75 n22609_not ; n22781
g22718 and n3028 n22406_not ; n22782
g22719 nor n22781 n22782 ; n22783
g22720 and n22780_not n22783 ; n22784
g22721 nor n22779 n22784 ; n22785
g22722 nor n22779 n22785 ; n22786
g22723 nor n22784 n22785 ; n22787
g22724 nor n22786 n22787 ; n22788
g22725 nor n22737 n22788 ; n22789
g22726 nor n22737 n22789 ; n22790
g22727 nor n22788 n22789 ; n22791
g22728 nor n22790 n22791 ; n22792
g22729 and n22631 n22632 ; n22793
g22730 nor n22636 n22793 ; n22794
g22731 nor n22792 n22794 ; n22795
g22732 nor n22792 n22795 ; n22796
g22733 nor n22794 n22795 ; n22797
g22734 nor n22796 n22797 ; n22798
g22735 and n3884 n22384 ; n22799
g22736 and n3967 n22390 ; n22800
g22737 and n4046 n22387 ; n22801
g22738 nor n22800 n22801 ; n22802
g22739 and n22799_not n22802 ; n22803
g22740 and n4050_not n22803 ; n22804
g22741 and n22425 n22427_not ; n22805
g22742 nor n22428 n22805 ; n22806
g22743 and n22803 n22806_not ; n22807
g22744 nor n22804 n22807 ; n22808
g22745 and a[26] n22808_not ; n22809
g22746 and a[26]_not n22808 ; n22810
g22747 nor n22809 n22810 ; n22811
g22748 nor n22798 n22811 ; n22812
g22749 nor n22798 n22812 ; n22813
g22750 nor n22811 n22812 ; n22814
g22751 nor n22813 n22814 ; n22815
g22752 nor n22726 n22815 ; n22816
g22753 nor n22726 n22816 ; n22817
g22754 nor n22815 n22816 ; n22818
g22755 nor n22817 n22818 ; n22819
g22756 nor n22575 n22819 ; n22820
g22757 nor n22575 n22820 ; n22821
g22758 nor n22819 n22820 ; n22822
g22759 nor n22821 n22822 ; n22823
g22760 and n22642 n22724 ; n22824
g22761 nor n22725 n22824 ; n22825
g22762 and n4694 n22377 ; n22826
g22763 and n4533 n22384 ; n22827
g22764 and n4604 n22380 ; n22828
g22765 nor n22827 n22828 ; n22829
g22766 and n22826_not n22829 ; n22830
g22767 and n4536_not n22830 ; n22831
g22768 nor n22433 n22435 ; n22832
g22769 and n22382_not n22436 ; n22833
g22770 nor n22832 n22833 ; n22834
g22771 and n22830 n22834 ; n22835
g22772 nor n22831 n22835 ; n22836
g22773 and a[23] n22836_not ; n22837
g22774 and a[23]_not n22836 ; n22838
g22775 nor n22837 n22838 ; n22839
g22776 and n22825 n22839_not ; n22840
g22777 and n22661 n22722 ; n22841
g22778 nor n22723 n22841 ; n22842
g22779 and n4694 n22380 ; n22843
g22780 and n4533 n22387 ; n22844
g22781 and n4604 n22384 ; n22845
g22782 nor n22844 n22845 ; n22846
g22783 and n22843_not n22846 ; n22847
g22784 and n4536_not n22847 ; n22848
g22785 and n22429 n22431_not ; n22849
g22786 nor n22432 n22849 ; n22850
g22787 and n22847 n22850_not ; n22851
g22788 nor n22848 n22851 ; n22852
g22789 and a[23] n22852_not ; n22853
g22790 and a[23]_not n22852 ; n22854
g22791 nor n22853 n22854 ; n22855
g22792 and n22842 n22855_not ; n22856
g22793 and n4694 n22384 ; n22857
g22794 and n4533 n22390 ; n22858
g22795 and n4604 n22387 ; n22859
g22796 nor n22858 n22859 ; n22860
g22797 and n22857_not n22860 ; n22861
g22798 and n4536 n22806 ; n22862
g22799 and n22861 n22862_not ; n22863
g22800 and a[23] n22863_not ; n22864
g22801 nor n22863 n22864 ; n22865
g22802 and a[23] n22864_not ; n22866
g22803 nor n22865 n22866 ; n22867
g22804 and n22718 n22720_not ; n22868
g22805 nor n22721 n22868 ; n22869
g22806 and n22867_not n22869 ; n22870
g22807 nor n22867 n22870 ; n22871
g22808 and n22869 n22870_not ; n22872
g22809 nor n22871 n22872 ; n22873
g22810 nor n22705 n22717 ; n22874
g22811 nor n22716 n22717 ; n22875
g22812 nor n22874 n22875 ; n22876
g22813 and n4694 n22387 ; n22877
g22814 and n4533 n22393 ; n22878
g22815 and n4604 n22390 ; n22879
g22816 nor n22878 n22879 ; n22880
g22817 and n22877_not n22880 ; n22881
g22818 and n4536_not n22881 ; n22882
g22819 and n22582_not n22881 ; n22883
g22820 nor n22882 n22883 ; n22884
g22821 and a[23] n22884_not ; n22885
g22822 and a[23]_not n22884 ; n22886
g22823 nor n22885 n22886 ; n22887
g22824 nor n22876 n22887 ; n22888
g22825 and n4694 n22390 ; n22889
g22826 and n4533 n22396 ; n22890
g22827 and n4604 n22393 ; n22891
g22828 nor n22890 n22891 ; n22892
g22829 and n22889_not n22892 ; n22893
g22830 and n4536 n22649 ; n22894
g22831 and n22893 n22894_not ; n22895
g22832 and a[23] n22895_not ; n22896
g22833 nor n22895 n22896 ; n22897
g22834 and a[23] n22896_not ; n22898
g22835 nor n22897 n22898 ; n22899
g22836 and n22689_not n22700 ; n22900
g22837 nor n22701 n22900 ; n22901
g22838 and n22899_not n22901 ; n22902
g22839 nor n22899 n22902 ; n22903
g22840 and n22901 n22902_not ; n22904
g22841 nor n22903 n22904 ; n22905
g22842 and n22679_not n22688 ; n22906
g22843 nor n22689 n22906 ; n22907
g22844 and n4694 n22393 ; n22908
g22845 and n4533 n22399 ; n22909
g22846 and n4604 n22396 ; n22910
g22847 nor n22909 n22910 ; n22911
g22848 and n22908_not n22911 ; n22912
g22849 and n4536_not n22912 ; n22913
g22850 and n22671_not n22912 ; n22914
g22851 nor n22913 n22914 ; n22915
g22852 and a[23] n22915_not ; n22916
g22853 and a[23]_not n22915 ; n22917
g22854 nor n22916 n22917 ; n22918
g22855 and n22907 n22918_not ; n22919
g22856 nor n4528 n22406 ; n22920
g22857 and a[23] n22920_not ; n22921
g22858 and n4604 n22406_not ; n22922
g22859 and n4694 n22402 ; n22923
g22860 nor n22922 n22923 ; n22924
g22861 and n4536 n22609_not ; n22925
g22862 and n22924 n22925_not ; n22926
g22863 and a[23] n22926_not ; n22927
g22864 and a[23] n22927_not ; n22928
g22865 nor n22926 n22927 ; n22929
g22866 nor n22928 n22929 ; n22930
g22867 and n22921 n22930_not ; n22931
g22868 and n4694 n22399 ; n22932
g22869 and n4533 n22406_not ; n22933
g22870 and n4604 n22402 ; n22934
g22871 nor n22933 n22934 ; n22935
g22872 and n22932_not n22935 ; n22936
g22873 and n4536_not n22936 ; n22937
g22874 and n22625 n22936 ; n22938
g22875 nor n22937 n22938 ; n22939
g22876 and a[23] n22939_not ; n22940
g22877 and a[23]_not n22939 ; n22941
g22878 nor n22940 n22941 ; n22942
g22879 and n22931 n22942_not ; n22943
g22880 and n22678 n22943 ; n22944
g22881 and n22943 n22944_not ; n22945
g22882 and n22678 n22944_not ; n22946
g22883 nor n22945 n22946 ; n22947
g22884 and n4694 n22396 ; n22948
g22885 and n4533 n22402 ; n22949
g22886 and n4604 n22399 ; n22950
g22887 nor n22949 n22950 ; n22951
g22888 and n22948_not n22951 ; n22952
g22889 and n4536 n22595 ; n22953
g22890 and n22952 n22953_not ; n22954
g22891 and a[23] n22954_not ; n22955
g22892 and a[23] n22955_not ; n22956
g22893 nor n22954 n22955 ; n22957
g22894 nor n22956 n22957 ; n22958
g22895 nor n22947 n22958 ; n22959
g22896 nor n22944 n22959 ; n22960
g22897 and n22907_not n22918 ; n22961
g22898 nor n22919 n22961 ; n22962
g22899 and n22960_not n22962 ; n22963
g22900 nor n22919 n22963 ; n22964
g22901 nor n22905 n22964 ; n22965
g22902 nor n22902 n22965 ; n22966
g22903 and n22876 n22887 ; n22967
g22904 nor n22888 n22967 ; n22968
g22905 and n22966_not n22968 ; n22969
g22906 nor n22888 n22969 ; n22970
g22907 nor n22873 n22970 ; n22971
g22908 nor n22870 n22971 ; n22972
g22909 and n22842 n22856_not ; n22973
g22910 nor n22855 n22856 ; n22974
g22911 nor n22973 n22974 ; n22975
g22912 nor n22972 n22975 ; n22976
g22913 nor n22856 n22976 ; n22977
g22914 and n22825_not n22839 ; n22978
g22915 nor n22840 n22978 ; n22979
g22916 and n22977_not n22979 ; n22980
g22917 nor n22840 n22980 ; n22981
g22918 and n22823 n22981 ; n22982
g22919 nor n22823 n22981 ; n22983
g22920 nor n22982 n22983 ; n22984
g22921 and n5496 n22365 ; n22985
g22922 and n4935 n22371 ; n22986
g22923 and n5407 n22368 ; n22987
g22924 nor n22986 n22987 ; n22988
g22925 and n22985_not n22988 ; n22989
g22926 and n4938_not n22989 ; n22990
g22927 nor n22448 n22451 ; n22991
g22928 and n22449_not n22452 ; n22992
g22929 nor n22991 n22992 ; n22993
g22930 and n22989 n22993 ; n22994
g22931 nor n22990 n22994 ; n22995
g22932 and a[20] n22995_not ; n22996
g22933 and a[20]_not n22995 ; n22997
g22934 nor n22996 n22997 ; n22998
g22935 and n22984 n22998_not ; n22999
g22936 and n5496 n22368 ; n23000
g22937 and n4935 n22374 ; n23001
g22938 and n5407 n22371 ; n23002
g22939 nor n23001 n23002 ; n23003
g22940 and n23000_not n23003 ; n23004
g22941 and n22444 n22446_not ; n23005
g22942 nor n22447 n23005 ; n23006
g22943 and n4938 n23006 ; n23007
g22944 and n23004 n23007_not ; n23008
g22945 and a[20] n23008_not ; n23009
g22946 nor n23008 n23009 ; n23010
g22947 and a[20] n23009_not ; n23011
g22948 nor n23010 n23011 ; n23012
g22949 and n22977 n22979_not ; n23013
g22950 nor n22980 n23013 ; n23014
g22951 and n23012_not n23014 ; n23015
g22952 nor n23012 n23015 ; n23016
g22953 and n23014 n23015_not ; n23017
g22954 nor n23016 n23017 ; n23018
g22955 and n5496 n22371 ; n23019
g22956 and n4935 n22377 ; n23020
g22957 and n5407 n22374 ; n23021
g22958 nor n23020 n23021 ; n23022
g22959 and n23019_not n23022 ; n23023
g22960 and n22440 n22442_not ; n23024
g22961 nor n22443 n23024 ; n23025
g22962 and n4938 n23025 ; n23026
g22963 and n23023 n23026_not ; n23027
g22964 and a[20] n23027_not ; n23028
g22965 nor n23027 n23028 ; n23029
g22966 and a[20] n23028_not ; n23030
g22967 nor n23029 n23030 ; n23031
g22968 nor n22972 n22976 ; n23032
g22969 nor n22975 n22976 ; n23033
g22970 nor n23032 n23033 ; n23034
g22971 nor n23031 n23034 ; n23035
g22972 nor n23031 n23035 ; n23036
g22973 nor n23034 n23035 ; n23037
g22974 nor n23036 n23037 ; n23038
g22975 and n22873 n22970 ; n23039
g22976 nor n22971 n23039 ; n23040
g22977 and n5496 n22374 ; n23041
g22978 and n4935 n22380 ; n23042
g22979 and n5407 n22377 ; n23043
g22980 nor n23042 n23043 ; n23044
g22981 and n23041_not n23044 ; n23045
g22982 and n4938_not n23045 ; n23046
g22983 and n22569_not n23045 ; n23047
g22984 nor n23046 n23047 ; n23048
g22985 and a[20] n23048_not ; n23049
g22986 and a[20]_not n23048 ; n23050
g22987 nor n23049 n23050 ; n23051
g22988 and n23040 n23051_not ; n23052
g22989 and n22966 n22968_not ; n23053
g22990 nor n22969 n23053 ; n23054
g22991 and n5496 n22377 ; n23055
g22992 and n4935 n22384 ; n23056
g22993 and n5407 n22380 ; n23057
g22994 nor n23056 n23057 ; n23058
g22995 and n23055_not n23058 ; n23059
g22996 and n4938_not n23059 ; n23060
g22997 and n22834 n23059 ; n23061
g22998 nor n23060 n23061 ; n23062
g22999 and a[20] n23062_not ; n23063
g23000 and a[20]_not n23062 ; n23064
g23001 nor n23063 n23064 ; n23065
g23002 and n23054 n23065_not ; n23066
g23003 and n22905 n22964 ; n23067
g23004 nor n22965 n23067 ; n23068
g23005 and n5496 n22380 ; n23069
g23006 and n4935 n22387 ; n23070
g23007 and n5407 n22384 ; n23071
g23008 nor n23070 n23071 ; n23072
g23009 and n23069_not n23072 ; n23073
g23010 and n4938_not n23073 ; n23074
g23011 and n22850_not n23073 ; n23075
g23012 nor n23074 n23075 ; n23076
g23013 and a[20] n23076_not ; n23077
g23014 and a[20]_not n23076 ; n23078
g23015 nor n23077 n23078 ; n23079
g23016 and n23068 n23079_not ; n23080
g23017 and n5496 n22384 ; n23081
g23018 and n4935 n22390 ; n23082
g23019 and n5407 n22387 ; n23083
g23020 nor n23082 n23083 ; n23084
g23021 and n23081_not n23084 ; n23085
g23022 and n4938 n22806 ; n23086
g23023 and n23085 n23086_not ; n23087
g23024 and a[20] n23087_not ; n23088
g23025 nor n23087 n23088 ; n23089
g23026 and a[20] n23088_not ; n23090
g23027 nor n23089 n23090 ; n23091
g23028 and n22960 n22962_not ; n23092
g23029 nor n22963 n23092 ; n23093
g23030 and n23091_not n23093 ; n23094
g23031 nor n23091 n23094 ; n23095
g23032 and n23093 n23094_not ; n23096
g23033 nor n23095 n23096 ; n23097
g23034 nor n22947 n22959 ; n23098
g23035 nor n22958 n22959 ; n23099
g23036 nor n23098 n23099 ; n23100
g23037 and n5496 n22387 ; n23101
g23038 and n4935 n22393 ; n23102
g23039 and n5407 n22390 ; n23103
g23040 nor n23102 n23103 ; n23104
g23041 and n23101_not n23104 ; n23105
g23042 and n4938_not n23105 ; n23106
g23043 and n22582_not n23105 ; n23107
g23044 nor n23106 n23107 ; n23108
g23045 and a[20] n23108_not ; n23109
g23046 and a[20]_not n23108 ; n23110
g23047 nor n23109 n23110 ; n23111
g23048 nor n23100 n23111 ; n23112
g23049 and n5496 n22390 ; n23113
g23050 and n4935 n22396 ; n23114
g23051 and n5407 n22393 ; n23115
g23052 nor n23114 n23115 ; n23116
g23053 and n23113_not n23116 ; n23117
g23054 and n4938 n22649 ; n23118
g23055 and n23117 n23118_not ; n23119
g23056 and a[20] n23119_not ; n23120
g23057 nor n23119 n23120 ; n23121
g23058 and a[20] n23120_not ; n23122
g23059 nor n23121 n23122 ; n23123
g23060 and n22931_not n22942 ; n23124
g23061 nor n22943 n23124 ; n23125
g23062 and n23123_not n23125 ; n23126
g23063 nor n23123 n23126 ; n23127
g23064 and n23125 n23126_not ; n23128
g23065 nor n23127 n23128 ; n23129
g23066 and n22921_not n22930 ; n23130
g23067 nor n22931 n23130 ; n23131
g23068 and n5496 n22393 ; n23132
g23069 and n4935 n22399 ; n23133
g23070 and n5407 n22396 ; n23134
g23071 nor n23133 n23134 ; n23135
g23072 and n23132_not n23135 ; n23136
g23073 and n4938_not n23136 ; n23137
g23074 and n22671_not n23136 ; n23138
g23075 nor n23137 n23138 ; n23139
g23076 and a[20] n23139_not ; n23140
g23077 and a[20]_not n23139 ; n23141
g23078 nor n23140 n23141 ; n23142
g23079 and n23131 n23142_not ; n23143
g23080 and n5407 n22406_not ; n23144
g23081 and n5496 n22402 ; n23145
g23082 nor n23144 n23145 ; n23146
g23083 and n4938 n22609_not ; n23147
g23084 and n23146 n23147_not ; n23148
g23085 and a[20] n23148_not ; n23149
g23086 and a[20] n23149_not ; n23150
g23087 nor n23148 n23149 ; n23151
g23088 nor n23150 n23151 ; n23152
g23089 nor n4933 n22406 ; n23153
g23090 and a[20] n23153_not ; n23154
g23091 and n23152_not n23154 ; n23155
g23092 and n5496 n22399 ; n23156
g23093 and n4935 n22406_not ; n23157
g23094 and n5407 n22402 ; n23158
g23095 nor n23157 n23158 ; n23159
g23096 and n23156_not n23159 ; n23160
g23097 and n4938_not n23160 ; n23161
g23098 and n22625 n23160 ; n23162
g23099 nor n23161 n23162 ; n23163
g23100 and a[20] n23163_not ; n23164
g23101 and a[20]_not n23163 ; n23165
g23102 nor n23164 n23165 ; n23166
g23103 and n23155 n23166_not ; n23167
g23104 and n22920 n23167 ; n23168
g23105 and n23167 n23168_not ; n23169
g23106 and n22920 n23168_not ; n23170
g23107 nor n23169 n23170 ; n23171
g23108 and n5496 n22396 ; n23172
g23109 and n4935 n22402 ; n23173
g23110 and n5407 n22399 ; n23174
g23111 nor n23173 n23174 ; n23175
g23112 and n23172_not n23175 ; n23176
g23113 and n4938 n22595 ; n23177
g23114 and n23176 n23177_not ; n23178
g23115 and a[20] n23178_not ; n23179
g23116 and a[20] n23179_not ; n23180
g23117 nor n23178 n23179 ; n23181
g23118 nor n23180 n23181 ; n23182
g23119 nor n23171 n23182 ; n23183
g23120 nor n23168 n23183 ; n23184
g23121 and n23131_not n23142 ; n23185
g23122 nor n23143 n23185 ; n23186
g23123 and n23184_not n23186 ; n23187
g23124 nor n23143 n23187 ; n23188
g23125 nor n23129 n23188 ; n23189
g23126 nor n23126 n23189 ; n23190
g23127 and n23100 n23111 ; n23191
g23128 nor n23112 n23191 ; n23192
g23129 and n23190_not n23192 ; n23193
g23130 nor n23112 n23193 ; n23194
g23131 nor n23097 n23194 ; n23195
g23132 nor n23094 n23195 ; n23196
g23133 and n23068 n23080_not ; n23197
g23134 nor n23079 n23080 ; n23198
g23135 nor n23197 n23198 ; n23199
g23136 nor n23196 n23199 ; n23200
g23137 nor n23080 n23200 ; n23201
g23138 and n23054 n23066_not ; n23202
g23139 nor n23065 n23066 ; n23203
g23140 nor n23202 n23203 ; n23204
g23141 nor n23201 n23204 ; n23205
g23142 nor n23066 n23205 ; n23206
g23143 and n23040_not n23051 ; n23207
g23144 nor n23052 n23207 ; n23208
g23145 and n23206_not n23208 ; n23209
g23146 nor n23052 n23209 ; n23210
g23147 nor n23038 n23210 ; n23211
g23148 nor n23035 n23211 ; n23212
g23149 nor n23018 n23212 ; n23213
g23150 nor n23015 n23213 ; n23214
g23151 and n22984 n22999_not ; n23215
g23152 nor n22998 n22999 ; n23216
g23153 nor n23215 n23216 ; n23217
g23154 nor n23214 n23217 ; n23218
g23155 nor n22999 n23218 ; n23219
g23156 and n4694 n22371 ; n23220
g23157 and n4533 n22377 ; n23221
g23158 and n4604 n22374 ; n23222
g23159 nor n23221 n23222 ; n23223
g23160 and n23220_not n23223 ; n23224
g23161 and n4536 n23025 ; n23225
g23162 and n23224 n23225_not ; n23226
g23163 and a[23] n23226_not ; n23227
g23164 nor n23226 n23227 ; n23228
g23165 and a[23] n23227_not ; n23229
g23166 nor n23228 n23229 ; n23230
g23167 nor n22812 n22816 ; n23231
g23168 and n3457 n22390 ; n23232
g23169 and n3542 n22396 ; n23233
g23170 and n3606 n22393 ; n23234
g23171 nor n23233 n23234 ; n23235
g23172 and n23232_not n23235 ; n23236
g23173 and n3368 n22649 ; n23237
g23174 and n23236 n23237_not ; n23238
g23175 and a[29] n23238_not ; n23239
g23176 nor n23238 n23239 ; n23240
g23177 and a[29] n23239_not ; n23241
g23178 nor n23240 n23241 ; n23242
g23179 and n75 n22625_not ; n23243
g23180 and n3020 n22399 ; n23244
g23181 and n3023 n22406_not ; n23245
g23182 and n3028 n22402 ; n23246
g23183 nor n23245 n23246 ; n23247
g23184 and n23244_not n23247 ; n23248
g23185 and n23243_not n23248 ; n23249
g23186 nor n233 n332 ; n23250
g23187 and n86_not n23250 ; n23251
g23188 and n13774 n23251 ; n23252
g23189 and n3041 n23252 ; n23253
g23190 and n12387 n23253 ; n23254
g23191 and n732 n23254 ; n23255
g23192 and n3261 n23255 ; n23256
g23193 and n6625 n23256 ; n23257
g23194 and n5209 n23257 ; n23258
g23195 and n967 n23258 ; n23259
g23196 and n294 n23259 ; n23260
g23197 and n1129 n23260 ; n23261
g23198 and n731 n23261 ; n23262
g23199 and n15867 n23262 ; n23263
g23200 and n420_not n23263 ; n23264
g23201 and n280_not n23264 ; n23265
g23202 and n228_not n23265 ; n23266
g23203 and n980_not n23266 ; n23267
g23204 and n673_not n23267 ; n23268
g23205 and n567_not n23268 ; n23269
g23206 and n22785 n23269_not ; n23270
g23207 and n22785_not n23269 ; n23271
g23208 nor n23270 n23271 ; n23272
g23209 and n23249_not n23272 ; n23273
g23210 nor n23249 n23273 ; n23274
g23211 and n23272 n23273_not ; n23275
g23212 nor n23274 n23275 ; n23276
g23213 nor n23242 n23276 ; n23277
g23214 nor n23242 n23277 ; n23278
g23215 nor n23276 n23277 ; n23279
g23216 nor n23278 n23279 ; n23280
g23217 nor n22789 n22795 ; n23281
g23218 and n23280 n23281 ; n23282
g23219 nor n23280 n23281 ; n23283
g23220 nor n23282 n23283 ; n23284
g23221 and n3884 n22380 ; n23285
g23222 and n3967 n22387 ; n23286
g23223 and n4046 n22384 ; n23287
g23224 nor n23286 n23287 ; n23288
g23225 and n23285_not n23288 ; n23289
g23226 and n4050_not n23289 ; n23290
g23227 and n22850_not n23289 ; n23291
g23228 nor n23290 n23291 ; n23292
g23229 and a[26] n23292_not ; n23293
g23230 and a[26]_not n23292 ; n23294
g23231 nor n23293 n23294 ; n23295
g23232 and n23284 n23295_not ; n23296
g23233 and n23284 n23296_not ; n23297
g23234 nor n23295 n23296 ; n23298
g23235 nor n23297 n23298 ; n23299
g23236 nor n23231 n23299 ; n23300
g23237 nor n23231 n23300 ; n23301
g23238 nor n23299 n23300 ; n23302
g23239 nor n23301 n23302 ; n23303
g23240 nor n23230 n23303 ; n23304
g23241 nor n23230 n23304 ; n23305
g23242 nor n23303 n23304 ; n23306
g23243 nor n23305 n23306 ; n23307
g23244 nor n22820 n22983 ; n23308
g23245 and n23307 n23308 ; n23309
g23246 nor n23307 n23308 ; n23310
g23247 nor n23309 n23310 ; n23311
g23248 and n5496 n22362 ; n23312
g23249 and n4935 n22368 ; n23313
g23250 and n5407 n22365 ; n23314
g23251 nor n23313 n23314 ; n23315
g23252 and n23312_not n23315 ; n23316
g23253 and n4938_not n23316 ; n23317
g23254 nor n22452 n22455 ; n23318
g23255 and n22453_not n22456 ; n23319
g23256 nor n23318 n23319 ; n23320
g23257 and n23316 n23320 ; n23321
g23258 nor n23317 n23321 ; n23322
g23259 and a[20] n23322_not ; n23323
g23260 and a[20]_not n23322 ; n23324
g23261 nor n23323 n23324 ; n23325
g23262 and n23311 n23325_not ; n23326
g23263 and n23311 n23326_not ; n23327
g23264 nor n23325 n23326 ; n23328
g23265 nor n23327 n23328 ; n23329
g23266 nor n23219 n23329 ; n23330
g23267 nor n23219 n23330 ; n23331
g23268 nor n23329 n23330 ; n23332
g23269 nor n23331 n23332 ; n23333
g23270 nor n22562 n23333 ; n23334
g23271 nor n22562 n23334 ; n23335
g23272 nor n23333 n23334 ; n23336
g23273 nor n23335 n23336 ; n23337
g23274 and n6233 n22356 ; n23338
g23275 and n5663 n22362 ; n23339
g23276 and n5939 n22359 ; n23340
g23277 nor n23339 n23340 ; n23341
g23278 and n23338_not n23341 ; n23342
g23279 nor n22460 n22463 ; n23343
g23280 and n22461_not n22464 ; n23344
g23281 nor n23343 n23344 ; n23345
g23282 and n5666 n23345_not ; n23346
g23283 and n23342 n23346_not ; n23347
g23284 and a[17] n23347_not ; n23348
g23285 nor n23347 n23348 ; n23349
g23286 and a[17] n23348_not ; n23350
g23287 nor n23349 n23350 ; n23351
g23288 nor n23214 n23218 ; n23352
g23289 nor n23217 n23218 ; n23353
g23290 nor n23352 n23353 ; n23354
g23291 nor n23351 n23354 ; n23355
g23292 nor n23351 n23355 ; n23356
g23293 nor n23354 n23355 ; n23357
g23294 nor n23356 n23357 ; n23358
g23295 and n23018 n23212 ; n23359
g23296 nor n23213 n23359 ; n23360
g23297 and n6233 n22359 ; n23361
g23298 and n5663 n22365 ; n23362
g23299 and n5939 n22362 ; n23363
g23300 nor n23362 n23363 ; n23364
g23301 and n23361_not n23364 ; n23365
g23302 and n5666_not n23365 ; n23366
g23303 and n22456 n22458_not ; n23367
g23304 nor n22459 n23367 ; n23368
g23305 and n23365 n23368_not ; n23369
g23306 nor n23366 n23369 ; n23370
g23307 and a[17] n23370_not ; n23371
g23308 and a[17]_not n23370 ; n23372
g23309 nor n23371 n23372 ; n23373
g23310 and n23360 n23373_not ; n23374
g23311 and n23038 n23210 ; n23375
g23312 nor n23211 n23375 ; n23376
g23313 and n6233 n22362 ; n23377
g23314 and n5663 n22368 ; n23378
g23315 and n5939 n22365 ; n23379
g23316 nor n23378 n23379 ; n23380
g23317 and n23377_not n23380 ; n23381
g23318 and n5666_not n23381 ; n23382
g23319 and n23320 n23381 ; n23383
g23320 nor n23382 n23383 ; n23384
g23321 and a[17] n23384_not ; n23385
g23322 and a[17]_not n23384 ; n23386
g23323 nor n23385 n23386 ; n23387
g23324 and n23376 n23387_not ; n23388
g23325 and n6233 n22365 ; n23389
g23326 and n5663 n22371 ; n23390
g23327 and n5939 n22368 ; n23391
g23328 nor n23390 n23391 ; n23392
g23329 and n23389_not n23392 ; n23393
g23330 and n5666 n22993_not ; n23394
g23331 and n23393 n23394_not ; n23395
g23332 and a[17] n23395_not ; n23396
g23333 nor n23395 n23396 ; n23397
g23334 and a[17] n23396_not ; n23398
g23335 nor n23397 n23398 ; n23399
g23336 and n23206 n23208_not ; n23400
g23337 nor n23209 n23400 ; n23401
g23338 and n23399_not n23401 ; n23402
g23339 nor n23399 n23402 ; n23403
g23340 and n23401 n23402_not ; n23404
g23341 nor n23403 n23404 ; n23405
g23342 and n6233 n22368 ; n23406
g23343 and n5663 n22374 ; n23407
g23344 and n5939 n22371 ; n23408
g23345 nor n23407 n23408 ; n23409
g23346 and n23406_not n23409 ; n23410
g23347 and n5666 n23006 ; n23411
g23348 and n23410 n23411_not ; n23412
g23349 and a[17] n23412_not ; n23413
g23350 nor n23412 n23413 ; n23414
g23351 and a[17] n23413_not ; n23415
g23352 nor n23414 n23415 ; n23416
g23353 nor n23201 n23205 ; n23417
g23354 nor n23204 n23205 ; n23418
g23355 nor n23417 n23418 ; n23419
g23356 nor n23416 n23419 ; n23420
g23357 nor n23416 n23420 ; n23421
g23358 nor n23419 n23420 ; n23422
g23359 nor n23421 n23422 ; n23423
g23360 and n6233 n22371 ; n23424
g23361 and n5663 n22377 ; n23425
g23362 and n5939 n22374 ; n23426
g23363 nor n23425 n23426 ; n23427
g23364 and n23424_not n23427 ; n23428
g23365 and n5666 n23025 ; n23429
g23366 and n23428 n23429_not ; n23430
g23367 and a[17] n23430_not ; n23431
g23368 nor n23430 n23431 ; n23432
g23369 and a[17] n23431_not ; n23433
g23370 nor n23432 n23433 ; n23434
g23371 nor n23196 n23200 ; n23435
g23372 nor n23199 n23200 ; n23436
g23373 nor n23435 n23436 ; n23437
g23374 nor n23434 n23437 ; n23438
g23375 nor n23434 n23438 ; n23439
g23376 nor n23437 n23438 ; n23440
g23377 nor n23439 n23440 ; n23441
g23378 and n23097 n23194 ; n23442
g23379 nor n23195 n23442 ; n23443
g23380 and n6233 n22374 ; n23444
g23381 and n5663 n22380 ; n23445
g23382 and n5939 n22377 ; n23446
g23383 nor n23445 n23446 ; n23447
g23384 and n23444_not n23447 ; n23448
g23385 and n5666_not n23448 ; n23449
g23386 and n22569_not n23448 ; n23450
g23387 nor n23449 n23450 ; n23451
g23388 and a[17] n23451_not ; n23452
g23389 and a[17]_not n23451 ; n23453
g23390 nor n23452 n23453 ; n23454
g23391 and n23443 n23454_not ; n23455
g23392 and n23190 n23192_not ; n23456
g23393 nor n23193 n23456 ; n23457
g23394 and n6233 n22377 ; n23458
g23395 and n5663 n22384 ; n23459
g23396 and n5939 n22380 ; n23460
g23397 nor n23459 n23460 ; n23461
g23398 and n23458_not n23461 ; n23462
g23399 and n5666_not n23462 ; n23463
g23400 and n22834 n23462 ; n23464
g23401 nor n23463 n23464 ; n23465
g23402 and a[17] n23465_not ; n23466
g23403 and a[17]_not n23465 ; n23467
g23404 nor n23466 n23467 ; n23468
g23405 and n23457 n23468_not ; n23469
g23406 and n23129 n23188 ; n23470
g23407 nor n23189 n23470 ; n23471
g23408 and n6233 n22380 ; n23472
g23409 and n5663 n22387 ; n23473
g23410 and n5939 n22384 ; n23474
g23411 nor n23473 n23474 ; n23475
g23412 and n23472_not n23475 ; n23476
g23413 and n5666_not n23476 ; n23477
g23414 and n22850_not n23476 ; n23478
g23415 nor n23477 n23478 ; n23479
g23416 and a[17] n23479_not ; n23480
g23417 and a[17]_not n23479 ; n23481
g23418 nor n23480 n23481 ; n23482
g23419 and n23471 n23482_not ; n23483
g23420 and n6233 n22384 ; n23484
g23421 and n5663 n22390 ; n23485
g23422 and n5939 n22387 ; n23486
g23423 nor n23485 n23486 ; n23487
g23424 and n23484_not n23487 ; n23488
g23425 and n5666 n22806 ; n23489
g23426 and n23488 n23489_not ; n23490
g23427 and a[17] n23490_not ; n23491
g23428 nor n23490 n23491 ; n23492
g23429 and a[17] n23491_not ; n23493
g23430 nor n23492 n23493 ; n23494
g23431 and n23184 n23186_not ; n23495
g23432 nor n23187 n23495 ; n23496
g23433 and n23494_not n23496 ; n23497
g23434 nor n23494 n23497 ; n23498
g23435 and n23496 n23497_not ; n23499
g23436 nor n23498 n23499 ; n23500
g23437 nor n23171 n23183 ; n23501
g23438 nor n23182 n23183 ; n23502
g23439 nor n23501 n23502 ; n23503
g23440 and n6233 n22387 ; n23504
g23441 and n5663 n22393 ; n23505
g23442 and n5939 n22390 ; n23506
g23443 nor n23505 n23506 ; n23507
g23444 and n23504_not n23507 ; n23508
g23445 and n5666_not n23508 ; n23509
g23446 and n22582_not n23508 ; n23510
g23447 nor n23509 n23510 ; n23511
g23448 and a[17] n23511_not ; n23512
g23449 and a[17]_not n23511 ; n23513
g23450 nor n23512 n23513 ; n23514
g23451 nor n23503 n23514 ; n23515
g23452 and n6233 n22390 ; n23516
g23453 and n5663 n22396 ; n23517
g23454 and n5939 n22393 ; n23518
g23455 nor n23517 n23518 ; n23519
g23456 and n23516_not n23519 ; n23520
g23457 and n5666 n22649 ; n23521
g23458 and n23520 n23521_not ; n23522
g23459 and a[17] n23522_not ; n23523
g23460 nor n23522 n23523 ; n23524
g23461 and a[17] n23523_not ; n23525
g23462 nor n23524 n23525 ; n23526
g23463 and n23155_not n23166 ; n23527
g23464 nor n23167 n23527 ; n23528
g23465 and n23526_not n23528 ; n23529
g23466 nor n23526 n23529 ; n23530
g23467 and n23528 n23529_not ; n23531
g23468 nor n23530 n23531 ; n23532
g23469 and n23152 n23154_not ; n23533
g23470 nor n23155 n23533 ; n23534
g23471 and n6233 n22393 ; n23535
g23472 and n5663 n22399 ; n23536
g23473 and n5939 n22396 ; n23537
g23474 nor n23536 n23537 ; n23538
g23475 and n23535_not n23538 ; n23539
g23476 and n5666_not n23539 ; n23540
g23477 and n22671_not n23539 ; n23541
g23478 nor n23540 n23541 ; n23542
g23479 and a[17] n23542_not ; n23543
g23480 and a[17]_not n23542 ; n23544
g23481 nor n23543 n23544 ; n23545
g23482 and n23534 n23545_not ; n23546
g23483 and n5939 n22406_not ; n23547
g23484 and n6233 n22402 ; n23548
g23485 nor n23547 n23548 ; n23549
g23486 and n5666 n22609_not ; n23550
g23487 and n23549 n23550_not ; n23551
g23488 and a[17] n23551_not ; n23552
g23489 and a[17] n23552_not ; n23553
g23490 nor n23551 n23552 ; n23554
g23491 nor n23553 n23554 ; n23555
g23492 nor n5658 n22406 ; n23556
g23493 and a[17] n23556_not ; n23557
g23494 and n23555_not n23557 ; n23558
g23495 and n6233 n22399 ; n23559
g23496 and n5663 n22406_not ; n23560
g23497 and n5939 n22402 ; n23561
g23498 nor n23560 n23561 ; n23562
g23499 and n23559_not n23562 ; n23563
g23500 and n5666_not n23563 ; n23564
g23501 and n22625 n23563 ; n23565
g23502 nor n23564 n23565 ; n23566
g23503 and a[17] n23566_not ; n23567
g23504 and a[17]_not n23566 ; n23568
g23505 nor n23567 n23568 ; n23569
g23506 and n23558 n23569_not ; n23570
g23507 and n23153 n23570 ; n23571
g23508 and n23570 n23571_not ; n23572
g23509 and n23153 n23571_not ; n23573
g23510 nor n23572 n23573 ; n23574
g23511 and n6233 n22396 ; n23575
g23512 and n5663 n22402 ; n23576
g23513 and n5939 n22399 ; n23577
g23514 nor n23576 n23577 ; n23578
g23515 and n23575_not n23578 ; n23579
g23516 and n5666 n22595 ; n23580
g23517 and n23579 n23580_not ; n23581
g23518 and a[17] n23581_not ; n23582
g23519 and a[17] n23582_not ; n23583
g23520 nor n23581 n23582 ; n23584
g23521 nor n23583 n23584 ; n23585
g23522 nor n23574 n23585 ; n23586
g23523 nor n23571 n23586 ; n23587
g23524 and n23534_not n23545 ; n23588
g23525 nor n23546 n23588 ; n23589
g23526 and n23587_not n23589 ; n23590
g23527 nor n23546 n23590 ; n23591
g23528 nor n23532 n23591 ; n23592
g23529 nor n23529 n23592 ; n23593
g23530 and n23503 n23514 ; n23594
g23531 nor n23515 n23594 ; n23595
g23532 and n23593_not n23595 ; n23596
g23533 nor n23515 n23596 ; n23597
g23534 nor n23500 n23597 ; n23598
g23535 nor n23497 n23598 ; n23599
g23536 and n23471 n23483_not ; n23600
g23537 nor n23482 n23483 ; n23601
g23538 nor n23600 n23601 ; n23602
g23539 nor n23599 n23602 ; n23603
g23540 nor n23483 n23603 ; n23604
g23541 and n23457 n23469_not ; n23605
g23542 nor n23468 n23469 ; n23606
g23543 nor n23605 n23606 ; n23607
g23544 nor n23604 n23607 ; n23608
g23545 nor n23469 n23608 ; n23609
g23546 and n23443_not n23454 ; n23610
g23547 nor n23455 n23610 ; n23611
g23548 and n23609_not n23611 ; n23612
g23549 nor n23455 n23612 ; n23613
g23550 nor n23441 n23613 ; n23614
g23551 nor n23438 n23614 ; n23615
g23552 nor n23423 n23615 ; n23616
g23553 nor n23420 n23616 ; n23617
g23554 nor n23405 n23617 ; n23618
g23555 nor n23402 n23618 ; n23619
g23556 and n23376 n23388_not ; n23620
g23557 nor n23387 n23388 ; n23621
g23558 nor n23620 n23621 ; n23622
g23559 nor n23619 n23622 ; n23623
g23560 nor n23388 n23623 ; n23624
g23561 and n23360_not n23373 ; n23625
g23562 nor n23374 n23625 ; n23626
g23563 and n23624_not n23626 ; n23627
g23564 nor n23374 n23627 ; n23628
g23565 nor n23358 n23628 ; n23629
g23566 nor n23355 n23629 ; n23630
g23567 and n23337 n23630 ; n23631
g23568 nor n23337 n23630 ; n23632
g23569 nor n23631 n23632 ; n23633
g23570 and n7101 n22344 ; n23634
g23571 and n6402 n22350 ; n23635
g23572 and n6951 n22347 ; n23636
g23573 nor n23635 n23636 ; n23637
g23574 and n23634_not n23637 ; n23638
g23575 and n6397_not n23638 ; n23639
g23576 nor n22476 n22479 ; n23640
g23577 and n22477_not n22480 ; n23641
g23578 nor n23640 n23641 ; n23642
g23579 and n23638 n23642 ; n23643
g23580 nor n23639 n23643 ; n23644
g23581 and a[14] n23644_not ; n23645
g23582 and a[14]_not n23644 ; n23646
g23583 nor n23645 n23646 ; n23647
g23584 and n23633 n23647_not ; n23648
g23585 and n23358 n23628 ; n23649
g23586 nor n23629 n23649 ; n23650
g23587 and n7101 n22347 ; n23651
g23588 and n6402 n22353 ; n23652
g23589 and n6951 n22350 ; n23653
g23590 nor n23652 n23653 ; n23654
g23591 and n23651_not n23654 ; n23655
g23592 and n6397_not n23655 ; n23656
g23593 nor n22472 n22475 ; n23657
g23594 and n22473_not n22476 ; n23658
g23595 nor n23657 n23658 ; n23659
g23596 and n23655 n23659 ; n23660
g23597 nor n23656 n23660 ; n23661
g23598 and a[14] n23661_not ; n23662
g23599 and a[14]_not n23661 ; n23663
g23600 nor n23662 n23663 ; n23664
g23601 and n23650 n23664_not ; n23665
g23602 and n7101 n22350 ; n23666
g23603 and n6402 n22356 ; n23667
g23604 and n6951 n22353 ; n23668
g23605 nor n23667 n23668 ; n23669
g23606 and n23666_not n23669 ; n23670
g23607 and n22468 n22470_not ; n23671
g23608 nor n22471 n23671 ; n23672
g23609 and n6397 n23672 ; n23673
g23610 and n23670 n23673_not ; n23674
g23611 and a[14] n23674_not ; n23675
g23612 nor n23674 n23675 ; n23676
g23613 and a[14] n23675_not ; n23677
g23614 nor n23676 n23677 ; n23678
g23615 and n23624 n23626_not ; n23679
g23616 nor n23627 n23679 ; n23680
g23617 and n23678_not n23680 ; n23681
g23618 nor n23678 n23681 ; n23682
g23619 and n23680 n23681_not ; n23683
g23620 nor n23682 n23683 ; n23684
g23621 and n7101 n22353 ; n23685
g23622 and n6402 n22359 ; n23686
g23623 and n6951 n22356 ; n23687
g23624 nor n23686 n23687 ; n23688
g23625 and n23685_not n23688 ; n23689
g23626 and n6397 n22556_not ; n23690
g23627 and n23689 n23690_not ; n23691
g23628 and a[14] n23691_not ; n23692
g23629 nor n23691 n23692 ; n23693
g23630 and a[14] n23692_not ; n23694
g23631 nor n23693 n23694 ; n23695
g23632 nor n23619 n23623 ; n23696
g23633 nor n23622 n23623 ; n23697
g23634 nor n23696 n23697 ; n23698
g23635 nor n23695 n23698 ; n23699
g23636 nor n23695 n23699 ; n23700
g23637 nor n23698 n23699 ; n23701
g23638 nor n23700 n23701 ; n23702
g23639 and n23405 n23617 ; n23703
g23640 nor n23618 n23703 ; n23704
g23641 and n7101 n22356 ; n23705
g23642 and n6402 n22362 ; n23706
g23643 and n6951 n22359 ; n23707
g23644 nor n23706 n23707 ; n23708
g23645 and n23705_not n23708 ; n23709
g23646 and n6397_not n23709 ; n23710
g23647 and n23345 n23709 ; n23711
g23648 nor n23710 n23711 ; n23712
g23649 and a[14] n23712_not ; n23713
g23650 and a[14]_not n23712 ; n23714
g23651 nor n23713 n23714 ; n23715
g23652 and n23704 n23715_not ; n23716
g23653 and n23423 n23615 ; n23717
g23654 nor n23616 n23717 ; n23718
g23655 and n7101 n22359 ; n23719
g23656 and n6402 n22365 ; n23720
g23657 and n6951 n22362 ; n23721
g23658 nor n23720 n23721 ; n23722
g23659 and n23719_not n23722 ; n23723
g23660 and n6397_not n23723 ; n23724
g23661 and n23368_not n23723 ; n23725
g23662 nor n23724 n23725 ; n23726
g23663 and a[14] n23726_not ; n23727
g23664 and a[14]_not n23726 ; n23728
g23665 nor n23727 n23728 ; n23729
g23666 and n23718 n23729_not ; n23730
g23667 and n23441 n23613 ; n23731
g23668 nor n23614 n23731 ; n23732
g23669 and n7101 n22362 ; n23733
g23670 and n6402 n22368 ; n23734
g23671 and n6951 n22365 ; n23735
g23672 nor n23734 n23735 ; n23736
g23673 and n23733_not n23736 ; n23737
g23674 and n6397_not n23737 ; n23738
g23675 and n23320 n23737 ; n23739
g23676 nor n23738 n23739 ; n23740
g23677 and a[14] n23740_not ; n23741
g23678 and a[14]_not n23740 ; n23742
g23679 nor n23741 n23742 ; n23743
g23680 and n23732 n23743_not ; n23744
g23681 and n7101 n22365 ; n23745
g23682 and n6402 n22371 ; n23746
g23683 and n6951 n22368 ; n23747
g23684 nor n23746 n23747 ; n23748
g23685 and n23745_not n23748 ; n23749
g23686 and n6397 n22993_not ; n23750
g23687 and n23749 n23750_not ; n23751
g23688 and a[14] n23751_not ; n23752
g23689 nor n23751 n23752 ; n23753
g23690 and a[14] n23752_not ; n23754
g23691 nor n23753 n23754 ; n23755
g23692 and n23609 n23611_not ; n23756
g23693 nor n23612 n23756 ; n23757
g23694 and n23755_not n23757 ; n23758
g23695 nor n23755 n23758 ; n23759
g23696 and n23757 n23758_not ; n23760
g23697 nor n23759 n23760 ; n23761
g23698 and n7101 n22368 ; n23762
g23699 and n6402 n22374 ; n23763
g23700 and n6951 n22371 ; n23764
g23701 nor n23763 n23764 ; n23765
g23702 and n23762_not n23765 ; n23766
g23703 and n6397 n23006 ; n23767
g23704 and n23766 n23767_not ; n23768
g23705 and a[14] n23768_not ; n23769
g23706 nor n23768 n23769 ; n23770
g23707 and a[14] n23769_not ; n23771
g23708 nor n23770 n23771 ; n23772
g23709 nor n23604 n23608 ; n23773
g23710 nor n23607 n23608 ; n23774
g23711 nor n23773 n23774 ; n23775
g23712 nor n23772 n23775 ; n23776
g23713 nor n23772 n23776 ; n23777
g23714 nor n23775 n23776 ; n23778
g23715 nor n23777 n23778 ; n23779
g23716 and n7101 n22371 ; n23780
g23717 and n6402 n22377 ; n23781
g23718 and n6951 n22374 ; n23782
g23719 nor n23781 n23782 ; n23783
g23720 and n23780_not n23783 ; n23784
g23721 and n6397 n23025 ; n23785
g23722 and n23784 n23785_not ; n23786
g23723 and a[14] n23786_not ; n23787
g23724 nor n23786 n23787 ; n23788
g23725 and a[14] n23787_not ; n23789
g23726 nor n23788 n23789 ; n23790
g23727 nor n23599 n23603 ; n23791
g23728 nor n23602 n23603 ; n23792
g23729 nor n23791 n23792 ; n23793
g23730 nor n23790 n23793 ; n23794
g23731 nor n23790 n23794 ; n23795
g23732 nor n23793 n23794 ; n23796
g23733 nor n23795 n23796 ; n23797
g23734 and n23500 n23597 ; n23798
g23735 nor n23598 n23798 ; n23799
g23736 and n7101 n22374 ; n23800
g23737 and n6402 n22380 ; n23801
g23738 and n6951 n22377 ; n23802
g23739 nor n23801 n23802 ; n23803
g23740 and n23800_not n23803 ; n23804
g23741 and n6397_not n23804 ; n23805
g23742 and n22569_not n23804 ; n23806
g23743 nor n23805 n23806 ; n23807
g23744 and a[14] n23807_not ; n23808
g23745 and a[14]_not n23807 ; n23809
g23746 nor n23808 n23809 ; n23810
g23747 and n23799 n23810_not ; n23811
g23748 and n23593 n23595_not ; n23812
g23749 nor n23596 n23812 ; n23813
g23750 and n7101 n22377 ; n23814
g23751 and n6402 n22384 ; n23815
g23752 and n6951 n22380 ; n23816
g23753 nor n23815 n23816 ; n23817
g23754 and n23814_not n23817 ; n23818
g23755 and n6397_not n23818 ; n23819
g23756 and n22834 n23818 ; n23820
g23757 nor n23819 n23820 ; n23821
g23758 and a[14] n23821_not ; n23822
g23759 and a[14]_not n23821 ; n23823
g23760 nor n23822 n23823 ; n23824
g23761 and n23813 n23824_not ; n23825
g23762 and n23532 n23591 ; n23826
g23763 nor n23592 n23826 ; n23827
g23764 and n7101 n22380 ; n23828
g23765 and n6402 n22387 ; n23829
g23766 and n6951 n22384 ; n23830
g23767 nor n23829 n23830 ; n23831
g23768 and n23828_not n23831 ; n23832
g23769 and n6397_not n23832 ; n23833
g23770 and n22850_not n23832 ; n23834
g23771 nor n23833 n23834 ; n23835
g23772 and a[14] n23835_not ; n23836
g23773 and a[14]_not n23835 ; n23837
g23774 nor n23836 n23837 ; n23838
g23775 and n23827 n23838_not ; n23839
g23776 and n7101 n22384 ; n23840
g23777 and n6402 n22390 ; n23841
g23778 and n6951 n22387 ; n23842
g23779 nor n23841 n23842 ; n23843
g23780 and n23840_not n23843 ; n23844
g23781 and n6397 n22806 ; n23845
g23782 and n23844 n23845_not ; n23846
g23783 and a[14] n23846_not ; n23847
g23784 nor n23846 n23847 ; n23848
g23785 and a[14] n23847_not ; n23849
g23786 nor n23848 n23849 ; n23850
g23787 and n23587 n23589_not ; n23851
g23788 nor n23590 n23851 ; n23852
g23789 and n23850_not n23852 ; n23853
g23790 nor n23850 n23853 ; n23854
g23791 and n23852 n23853_not ; n23855
g23792 nor n23854 n23855 ; n23856
g23793 nor n23574 n23586 ; n23857
g23794 nor n23585 n23586 ; n23858
g23795 nor n23857 n23858 ; n23859
g23796 and n7101 n22387 ; n23860
g23797 and n6402 n22393 ; n23861
g23798 and n6951 n22390 ; n23862
g23799 nor n23861 n23862 ; n23863
g23800 and n23860_not n23863 ; n23864
g23801 and n6397_not n23864 ; n23865
g23802 and n22582_not n23864 ; n23866
g23803 nor n23865 n23866 ; n23867
g23804 and a[14] n23867_not ; n23868
g23805 and a[14]_not n23867 ; n23869
g23806 nor n23868 n23869 ; n23870
g23807 nor n23859 n23870 ; n23871
g23808 and n7101 n22390 ; n23872
g23809 and n6402 n22396 ; n23873
g23810 and n6951 n22393 ; n23874
g23811 nor n23873 n23874 ; n23875
g23812 and n23872_not n23875 ; n23876
g23813 and n6397 n22649 ; n23877
g23814 and n23876 n23877_not ; n23878
g23815 and a[14] n23878_not ; n23879
g23816 nor n23878 n23879 ; n23880
g23817 and a[14] n23879_not ; n23881
g23818 nor n23880 n23881 ; n23882
g23819 and n23558_not n23569 ; n23883
g23820 nor n23570 n23883 ; n23884
g23821 and n23882_not n23884 ; n23885
g23822 nor n23882 n23885 ; n23886
g23823 and n23884 n23885_not ; n23887
g23824 nor n23886 n23887 ; n23888
g23825 and n23555 n23557_not ; n23889
g23826 nor n23558 n23889 ; n23890
g23827 and n7101 n22393 ; n23891
g23828 and n6402 n22399 ; n23892
g23829 and n6951 n22396 ; n23893
g23830 nor n23892 n23893 ; n23894
g23831 and n23891_not n23894 ; n23895
g23832 and n6397_not n23895 ; n23896
g23833 and n22671_not n23895 ; n23897
g23834 nor n23896 n23897 ; n23898
g23835 and a[14] n23898_not ; n23899
g23836 and a[14]_not n23898 ; n23900
g23837 nor n23899 n23900 ; n23901
g23838 and n23890 n23901_not ; n23902
g23839 and n6951 n22406_not ; n23903
g23840 and n7101 n22402 ; n23904
g23841 nor n23903 n23904 ; n23905
g23842 and n6397 n22609_not ; n23906
g23843 and n23905 n23906_not ; n23907
g23844 and a[14] n23907_not ; n23908
g23845 and a[14] n23908_not ; n23909
g23846 nor n23907 n23908 ; n23910
g23847 nor n23909 n23910 ; n23911
g23848 nor n6393 n22406 ; n23912
g23849 and a[14] n23912_not ; n23913
g23850 and n23911_not n23913 ; n23914
g23851 and n7101 n22399 ; n23915
g23852 and n6402 n22406_not ; n23916
g23853 and n6951 n22402 ; n23917
g23854 nor n23916 n23917 ; n23918
g23855 and n23915_not n23918 ; n23919
g23856 and n6397_not n23919 ; n23920
g23857 and n22625 n23919 ; n23921
g23858 nor n23920 n23921 ; n23922
g23859 and a[14] n23922_not ; n23923
g23860 and a[14]_not n23922 ; n23924
g23861 nor n23923 n23924 ; n23925
g23862 and n23914 n23925_not ; n23926
g23863 and n23556 n23926 ; n23927
g23864 and n23926 n23927_not ; n23928
g23865 and n23556 n23927_not ; n23929
g23866 nor n23928 n23929 ; n23930
g23867 and n7101 n22396 ; n23931
g23868 and n6402 n22402 ; n23932
g23869 and n6951 n22399 ; n23933
g23870 nor n23932 n23933 ; n23934
g23871 and n23931_not n23934 ; n23935
g23872 and n6397 n22595 ; n23936
g23873 and n23935 n23936_not ; n23937
g23874 and a[14] n23937_not ; n23938
g23875 and a[14] n23938_not ; n23939
g23876 nor n23937 n23938 ; n23940
g23877 nor n23939 n23940 ; n23941
g23878 nor n23930 n23941 ; n23942
g23879 nor n23927 n23942 ; n23943
g23880 and n23890_not n23901 ; n23944
g23881 nor n23902 n23944 ; n23945
g23882 and n23943_not n23945 ; n23946
g23883 nor n23902 n23946 ; n23947
g23884 nor n23888 n23947 ; n23948
g23885 nor n23885 n23948 ; n23949
g23886 and n23859 n23870 ; n23950
g23887 nor n23871 n23950 ; n23951
g23888 and n23949_not n23951 ; n23952
g23889 nor n23871 n23952 ; n23953
g23890 nor n23856 n23953 ; n23954
g23891 nor n23853 n23954 ; n23955
g23892 and n23827 n23839_not ; n23956
g23893 nor n23838 n23839 ; n23957
g23894 nor n23956 n23957 ; n23958
g23895 nor n23955 n23958 ; n23959
g23896 nor n23839 n23959 ; n23960
g23897 and n23813 n23825_not ; n23961
g23898 nor n23824 n23825 ; n23962
g23899 nor n23961 n23962 ; n23963
g23900 nor n23960 n23963 ; n23964
g23901 nor n23825 n23964 ; n23965
g23902 and n23799_not n23810 ; n23966
g23903 nor n23811 n23966 ; n23967
g23904 and n23965_not n23967 ; n23968
g23905 nor n23811 n23968 ; n23969
g23906 nor n23797 n23969 ; n23970
g23907 nor n23794 n23970 ; n23971
g23908 nor n23779 n23971 ; n23972
g23909 nor n23776 n23972 ; n23973
g23910 nor n23761 n23973 ; n23974
g23911 nor n23758 n23974 ; n23975
g23912 and n23732 n23744_not ; n23976
g23913 nor n23743 n23744 ; n23977
g23914 nor n23976 n23977 ; n23978
g23915 nor n23975 n23978 ; n23979
g23916 nor n23744 n23979 ; n23980
g23917 and n23718 n23730_not ; n23981
g23918 nor n23729 n23730 ; n23982
g23919 nor n23981 n23982 ; n23983
g23920 nor n23980 n23983 ; n23984
g23921 nor n23730 n23984 ; n23985
g23922 and n23704_not n23715 ; n23986
g23923 nor n23716 n23986 ; n23987
g23924 and n23985_not n23987 ; n23988
g23925 nor n23716 n23988 ; n23989
g23926 nor n23702 n23989 ; n23990
g23927 nor n23699 n23990 ; n23991
g23928 nor n23684 n23991 ; n23992
g23929 nor n23681 n23992 ; n23993
g23930 and n23650 n23665_not ; n23994
g23931 nor n23664 n23665 ; n23995
g23932 nor n23994 n23995 ; n23996
g23933 nor n23993 n23996 ; n23997
g23934 nor n23665 n23997 ; n23998
g23935 and n23633 n23648_not ; n23999
g23936 nor n23647 n23648 ; n24000
g23937 nor n23999 n24000 ; n24001
g23938 nor n23998 n24001 ; n24002
g23939 nor n23648 n24002 ; n24003
g23940 and n6233 n22350 ; n24004
g23941 and n5663 n22356 ; n24005
g23942 and n5939 n22353 ; n24006
g23943 nor n24005 n24006 ; n24007
g23944 and n24004_not n24007 ; n24008
g23945 and n5666 n23672 ; n24009
g23946 and n24008 n24009_not ; n24010
g23947 and a[17] n24010_not ; n24011
g23948 nor n24010 n24011 ; n24012
g23949 and a[17] n24011_not ; n24013
g23950 nor n24012 n24013 ; n24014
g23951 nor n23326 n23330 ; n24015
g23952 and n4694 n22368 ; n24016
g23953 and n4533 n22374 ; n24017
g23954 and n4604 n22371 ; n24018
g23955 nor n24017 n24018 ; n24019
g23956 and n24016_not n24019 ; n24020
g23957 and n4536 n23006 ; n24021
g23958 and n24020 n24021_not ; n24022
g23959 and a[23] n24022_not ; n24023
g23960 nor n24022 n24023 ; n24024
g23961 and a[23] n24023_not ; n24025
g23962 nor n24024 n24025 ; n24026
g23963 nor n23296 n23300 ; n24027
g23964 and n3457 n22387 ; n24028
g23965 and n3542 n22393 ; n24029
g23966 and n3606 n22390 ; n24030
g23967 nor n24029 n24030 ; n24031
g23968 and n24028_not n24031 ; n24032
g23969 and n3368 n22582 ; n24033
g23970 and n24032 n24033_not ; n24034
g23971 and a[29] n24034_not ; n24035
g23972 nor n24034 n24035 ; n24036
g23973 and a[29] n24035_not ; n24037
g23974 nor n24036 n24037 ; n24038
g23975 nor n23270 n23273 ; n24039
g23976 and n116 n511_not ; n24040
g23977 and n514_not n24040 ; n24041
g23978 and n1971 n5002 ; n24042
g23979 and n24041 n24042 ; n24043
g23980 and n4216 n24043 ; n24044
g23981 and n1621 n24044 ; n24045
g23982 and n5296 n24045 ; n24046
g23983 and n916 n24046 ; n24047
g23984 and n3290 n24047 ; n24048
g23985 and n2346 n24048 ; n24049
g23986 and n291 n24049 ; n24050
g23987 and n471 n24050 ; n24051
g23988 and n1531 n24051 ; n24052
g23989 and n520 n24052 ; n24053
g23990 and n118_not n24053 ; n24054
g23991 and n102_not n24054 ; n24055
g23992 and n791_not n24055 ; n24056
g23993 and n225_not n24056 ; n24057
g23994 and n3020 n22396 ; n24058
g23995 and n3028 n22399 ; n24059
g23996 and n3023 n22402 ; n24060
g23997 and n75 n22595 ; n24061
g23998 nor n24060 n24061 ; n24062
g23999 and n24059_not n24062 ; n24063
g24000 and n24058_not n24063 ; n24064
g24001 nor n24057 n24064 ; n24065
g24002 nor n24057 n24065 ; n24066
g24003 nor n24064 n24065 ; n24067
g24004 nor n24066 n24067 ; n24068
g24005 nor n24039 n24068 ; n24069
g24006 nor n24039 n24069 ; n24070
g24007 nor n24068 n24069 ; n24071
g24008 nor n24070 n24071 ; n24072
g24009 nor n24038 n24072 ; n24073
g24010 nor n24038 n24073 ; n24074
g24011 nor n24072 n24073 ; n24075
g24012 nor n24074 n24075 ; n24076
g24013 nor n23277 n23283 ; n24077
g24014 and n24076 n24077 ; n24078
g24015 nor n24076 n24077 ; n24079
g24016 nor n24078 n24079 ; n24080
g24017 and n3884 n22377 ; n24081
g24018 and n3967 n22384 ; n24082
g24019 and n4046 n22380 ; n24083
g24020 nor n24082 n24083 ; n24084
g24021 and n24081_not n24084 ; n24085
g24022 and n4050_not n24085 ; n24086
g24023 and n22834 n24085 ; n24087
g24024 nor n24086 n24087 ; n24088
g24025 and a[26] n24088_not ; n24089
g24026 and a[26]_not n24088 ; n24090
g24027 nor n24089 n24090 ; n24091
g24028 and n24080 n24091_not ; n24092
g24029 and n24080 n24092_not ; n24093
g24030 nor n24091 n24092 ; n24094
g24031 nor n24093 n24094 ; n24095
g24032 nor n24027 n24095 ; n24096
g24033 nor n24027 n24096 ; n24097
g24034 nor n24095 n24096 ; n24098
g24035 nor n24097 n24098 ; n24099
g24036 nor n24026 n24099 ; n24100
g24037 nor n24026 n24100 ; n24101
g24038 nor n24099 n24100 ; n24102
g24039 nor n24101 n24102 ; n24103
g24040 nor n23304 n23310 ; n24104
g24041 and n24103 n24104 ; n24105
g24042 nor n24103 n24104 ; n24106
g24043 nor n24105 n24106 ; n24107
g24044 and n5496 n22359 ; n24108
g24045 and n4935 n22365 ; n24109
g24046 and n5407 n22362 ; n24110
g24047 nor n24109 n24110 ; n24111
g24048 and n24108_not n24111 ; n24112
g24049 and n4938_not n24112 ; n24113
g24050 and n23368_not n24112 ; n24114
g24051 nor n24113 n24114 ; n24115
g24052 and a[20] n24115_not ; n24116
g24053 and a[20]_not n24115 ; n24117
g24054 nor n24116 n24117 ; n24118
g24055 and n24107 n24118_not ; n24119
g24056 and n24107 n24119_not ; n24120
g24057 nor n24118 n24119 ; n24121
g24058 nor n24120 n24121 ; n24122
g24059 nor n24015 n24122 ; n24123
g24060 nor n24015 n24123 ; n24124
g24061 nor n24122 n24123 ; n24125
g24062 nor n24124 n24125 ; n24126
g24063 nor n24014 n24126 ; n24127
g24064 nor n24014 n24127 ; n24128
g24065 nor n24126 n24127 ; n24129
g24066 nor n24128 n24129 ; n24130
g24067 nor n23334 n23632 ; n24131
g24068 and n24130 n24131 ; n24132
g24069 nor n24130 n24131 ; n24133
g24070 nor n24132 n24133 ; n24134
g24071 and n7101 n22341 ; n24135
g24072 and n6402 n22347 ; n24136
g24073 and n6951 n22344 ; n24137
g24074 nor n24136 n24137 ; n24138
g24075 and n24135_not n24138 ; n24139
g24076 and n6397_not n24139 ; n24140
g24077 and n22480 n22482_not ; n24141
g24078 nor n22483 n24141 ; n24142
g24079 and n24139 n24142_not ; n24143
g24080 nor n24140 n24143 ; n24144
g24081 and a[14] n24144_not ; n24145
g24082 and a[14]_not n24144 ; n24146
g24083 nor n24145 n24146 ; n24147
g24084 and n24134 n24147_not ; n24148
g24085 and n24134 n24148_not ; n24149
g24086 nor n24147 n24148 ; n24150
g24087 nor n24149 n24150 ; n24151
g24088 nor n24003 n24151 ; n24152
g24089 nor n24003 n24152 ; n24153
g24090 nor n24151 n24152 ; n24154
g24091 nor n24153 n24154 ; n24155
g24092 nor n22548 n24155 ; n24156
g24093 nor n22548 n24156 ; n24157
g24094 nor n24155 n24156 ; n24158
g24095 nor n24157 n24158 ; n24159
g24096 and n7983 n22335 ; n24160
g24097 and n7291 n22341 ; n24161
g24098 and n7632 n22338 ; n24162
g24099 nor n24161 n24162 ; n24163
g24100 and n24160_not n24163 ; n24164
g24101 nor n22488 n22491 ; n24165
g24102 and n22489_not n22492 ; n24166
g24103 nor n24165 n24166 ; n24167
g24104 and n7294 n24167_not ; n24168
g24105 and n24164 n24168_not ; n24169
g24106 and a[11] n24169_not ; n24170
g24107 nor n24169 n24170 ; n24171
g24108 and a[11] n24170_not ; n24172
g24109 nor n24171 n24172 ; n24173
g24110 nor n23998 n24002 ; n24174
g24111 nor n24001 n24002 ; n24175
g24112 nor n24174 n24175 ; n24176
g24113 nor n24173 n24176 ; n24177
g24114 nor n24173 n24177 ; n24178
g24115 nor n24176 n24177 ; n24179
g24116 nor n24178 n24179 ; n24180
g24117 and n7983 n22338 ; n24181
g24118 and n7291 n22344 ; n24182
g24119 and n7632 n22341 ; n24183
g24120 nor n24182 n24183 ; n24184
g24121 and n24181_not n24184 ; n24185
g24122 nor n22484 n22487 ; n24186
g24123 and n22485_not n22488 ; n24187
g24124 nor n24186 n24187 ; n24188
g24125 and n7294 n24188_not ; n24189
g24126 and n24185 n24189_not ; n24190
g24127 and a[11] n24190_not ; n24191
g24128 nor n24190 n24191 ; n24192
g24129 and a[11] n24191_not ; n24193
g24130 nor n24192 n24193 ; n24194
g24131 nor n23993 n23997 ; n24195
g24132 nor n23996 n23997 ; n24196
g24133 nor n24195 n24196 ; n24197
g24134 nor n24194 n24197 ; n24198
g24135 nor n24194 n24198 ; n24199
g24136 nor n24197 n24198 ; n24200
g24137 nor n24199 n24200 ; n24201
g24138 and n23684 n23991 ; n24202
g24139 nor n23992 n24202 ; n24203
g24140 and n7983 n22341 ; n24204
g24141 and n7291 n22347 ; n24205
g24142 and n7632 n22344 ; n24206
g24143 nor n24205 n24206 ; n24207
g24144 and n24204_not n24207 ; n24208
g24145 and n7294_not n24208 ; n24209
g24146 and n24142_not n24208 ; n24210
g24147 nor n24209 n24210 ; n24211
g24148 and a[11] n24211_not ; n24212
g24149 and a[11]_not n24211 ; n24213
g24150 nor n24212 n24213 ; n24214
g24151 and n24203 n24214_not ; n24215
g24152 and n23702 n23989 ; n24216
g24153 nor n23990 n24216 ; n24217
g24154 and n7983 n22344 ; n24218
g24155 and n7291 n22350 ; n24219
g24156 and n7632 n22347 ; n24220
g24157 nor n24219 n24220 ; n24221
g24158 and n24218_not n24221 ; n24222
g24159 and n7294_not n24222 ; n24223
g24160 and n23642 n24222 ; n24224
g24161 nor n24223 n24224 ; n24225
g24162 and a[11] n24225_not ; n24226
g24163 and a[11]_not n24225 ; n24227
g24164 nor n24226 n24227 ; n24228
g24165 and n24217 n24228_not ; n24229
g24166 and n7983 n22347 ; n24230
g24167 and n7291 n22353 ; n24231
g24168 and n7632 n22350 ; n24232
g24169 nor n24231 n24232 ; n24233
g24170 and n24230_not n24233 ; n24234
g24171 and n7294 n23659_not ; n24235
g24172 and n24234 n24235_not ; n24236
g24173 and a[11] n24236_not ; n24237
g24174 nor n24236 n24237 ; n24238
g24175 and a[11] n24237_not ; n24239
g24176 nor n24238 n24239 ; n24240
g24177 and n23985 n23987_not ; n24241
g24178 nor n23988 n24241 ; n24242
g24179 and n24240_not n24242 ; n24243
g24180 nor n24240 n24243 ; n24244
g24181 and n24242 n24243_not ; n24245
g24182 nor n24244 n24245 ; n24246
g24183 and n7983 n22350 ; n24247
g24184 and n7291 n22356 ; n24248
g24185 and n7632 n22353 ; n24249
g24186 nor n24248 n24249 ; n24250
g24187 and n24247_not n24250 ; n24251
g24188 and n7294 n23672 ; n24252
g24189 and n24251 n24252_not ; n24253
g24190 and a[11] n24253_not ; n24254
g24191 nor n24253 n24254 ; n24255
g24192 and a[11] n24254_not ; n24256
g24193 nor n24255 n24256 ; n24257
g24194 nor n23980 n23984 ; n24258
g24195 nor n23983 n23984 ; n24259
g24196 nor n24258 n24259 ; n24260
g24197 nor n24257 n24260 ; n24261
g24198 nor n24257 n24261 ; n24262
g24199 nor n24260 n24261 ; n24263
g24200 nor n24262 n24263 ; n24264
g24201 and n7983 n22353 ; n24265
g24202 and n7291 n22359 ; n24266
g24203 and n7632 n22356 ; n24267
g24204 nor n24266 n24267 ; n24268
g24205 and n24265_not n24268 ; n24269
g24206 and n7294 n22556_not ; n24270
g24207 and n24269 n24270_not ; n24271
g24208 and a[11] n24271_not ; n24272
g24209 nor n24271 n24272 ; n24273
g24210 and a[11] n24272_not ; n24274
g24211 nor n24273 n24274 ; n24275
g24212 nor n23975 n23979 ; n24276
g24213 nor n23978 n23979 ; n24277
g24214 nor n24276 n24277 ; n24278
g24215 nor n24275 n24278 ; n24279
g24216 nor n24275 n24279 ; n24280
g24217 nor n24278 n24279 ; n24281
g24218 nor n24280 n24281 ; n24282
g24219 and n23761 n23973 ; n24283
g24220 nor n23974 n24283 ; n24284
g24221 and n7983 n22356 ; n24285
g24222 and n7291 n22362 ; n24286
g24223 and n7632 n22359 ; n24287
g24224 nor n24286 n24287 ; n24288
g24225 and n24285_not n24288 ; n24289
g24226 and n7294_not n24289 ; n24290
g24227 and n23345 n24289 ; n24291
g24228 nor n24290 n24291 ; n24292
g24229 and a[11] n24292_not ; n24293
g24230 and a[11]_not n24292 ; n24294
g24231 nor n24293 n24294 ; n24295
g24232 and n24284 n24295_not ; n24296
g24233 and n23779 n23971 ; n24297
g24234 nor n23972 n24297 ; n24298
g24235 and n7983 n22359 ; n24299
g24236 and n7291 n22365 ; n24300
g24237 and n7632 n22362 ; n24301
g24238 nor n24300 n24301 ; n24302
g24239 and n24299_not n24302 ; n24303
g24240 and n7294_not n24303 ; n24304
g24241 and n23368_not n24303 ; n24305
g24242 nor n24304 n24305 ; n24306
g24243 and a[11] n24306_not ; n24307
g24244 and a[11]_not n24306 ; n24308
g24245 nor n24307 n24308 ; n24309
g24246 and n24298 n24309_not ; n24310
g24247 and n23797 n23969 ; n24311
g24248 nor n23970 n24311 ; n24312
g24249 and n7983 n22362 ; n24313
g24250 and n7291 n22368 ; n24314
g24251 and n7632 n22365 ; n24315
g24252 nor n24314 n24315 ; n24316
g24253 and n24313_not n24316 ; n24317
g24254 and n7294_not n24317 ; n24318
g24255 and n23320 n24317 ; n24319
g24256 nor n24318 n24319 ; n24320
g24257 and a[11] n24320_not ; n24321
g24258 and a[11]_not n24320 ; n24322
g24259 nor n24321 n24322 ; n24323
g24260 and n24312 n24323_not ; n24324
g24261 and n7983 n22365 ; n24325
g24262 and n7291 n22371 ; n24326
g24263 and n7632 n22368 ; n24327
g24264 nor n24326 n24327 ; n24328
g24265 and n24325_not n24328 ; n24329
g24266 and n7294 n22993_not ; n24330
g24267 and n24329 n24330_not ; n24331
g24268 and a[11] n24331_not ; n24332
g24269 nor n24331 n24332 ; n24333
g24270 and a[11] n24332_not ; n24334
g24271 nor n24333 n24334 ; n24335
g24272 and n23965 n23967_not ; n24336
g24273 nor n23968 n24336 ; n24337
g24274 and n24335_not n24337 ; n24338
g24275 nor n24335 n24338 ; n24339
g24276 and n24337 n24338_not ; n24340
g24277 nor n24339 n24340 ; n24341
g24278 and n7983 n22368 ; n24342
g24279 and n7291 n22374 ; n24343
g24280 and n7632 n22371 ; n24344
g24281 nor n24343 n24344 ; n24345
g24282 and n24342_not n24345 ; n24346
g24283 and n7294 n23006 ; n24347
g24284 and n24346 n24347_not ; n24348
g24285 and a[11] n24348_not ; n24349
g24286 nor n24348 n24349 ; n24350
g24287 and a[11] n24349_not ; n24351
g24288 nor n24350 n24351 ; n24352
g24289 nor n23960 n23964 ; n24353
g24290 nor n23963 n23964 ; n24354
g24291 nor n24353 n24354 ; n24355
g24292 nor n24352 n24355 ; n24356
g24293 nor n24352 n24356 ; n24357
g24294 nor n24355 n24356 ; n24358
g24295 nor n24357 n24358 ; n24359
g24296 and n7983 n22371 ; n24360
g24297 and n7291 n22377 ; n24361
g24298 and n7632 n22374 ; n24362
g24299 nor n24361 n24362 ; n24363
g24300 and n24360_not n24363 ; n24364
g24301 and n7294 n23025 ; n24365
g24302 and n24364 n24365_not ; n24366
g24303 and a[11] n24366_not ; n24367
g24304 nor n24366 n24367 ; n24368
g24305 and a[11] n24367_not ; n24369
g24306 nor n24368 n24369 ; n24370
g24307 nor n23955 n23959 ; n24371
g24308 nor n23958 n23959 ; n24372
g24309 nor n24371 n24372 ; n24373
g24310 nor n24370 n24373 ; n24374
g24311 nor n24370 n24374 ; n24375
g24312 nor n24373 n24374 ; n24376
g24313 nor n24375 n24376 ; n24377
g24314 and n23856 n23953 ; n24378
g24315 nor n23954 n24378 ; n24379
g24316 and n7983 n22374 ; n24380
g24317 and n7291 n22380 ; n24381
g24318 and n7632 n22377 ; n24382
g24319 nor n24381 n24382 ; n24383
g24320 and n24380_not n24383 ; n24384
g24321 and n7294_not n24384 ; n24385
g24322 and n22569_not n24384 ; n24386
g24323 nor n24385 n24386 ; n24387
g24324 and a[11] n24387_not ; n24388
g24325 and a[11]_not n24387 ; n24389
g24326 nor n24388 n24389 ; n24390
g24327 and n24379 n24390_not ; n24391
g24328 and n23949 n23951_not ; n24392
g24329 nor n23952 n24392 ; n24393
g24330 and n7983 n22377 ; n24394
g24331 and n7291 n22384 ; n24395
g24332 and n7632 n22380 ; n24396
g24333 nor n24395 n24396 ; n24397
g24334 and n24394_not n24397 ; n24398
g24335 and n7294_not n24398 ; n24399
g24336 and n22834 n24398 ; n24400
g24337 nor n24399 n24400 ; n24401
g24338 and a[11] n24401_not ; n24402
g24339 and a[11]_not n24401 ; n24403
g24340 nor n24402 n24403 ; n24404
g24341 and n24393 n24404_not ; n24405
g24342 and n23888 n23947 ; n24406
g24343 nor n23948 n24406 ; n24407
g24344 and n7983 n22380 ; n24408
g24345 and n7291 n22387 ; n24409
g24346 and n7632 n22384 ; n24410
g24347 nor n24409 n24410 ; n24411
g24348 and n24408_not n24411 ; n24412
g24349 and n7294_not n24412 ; n24413
g24350 and n22850_not n24412 ; n24414
g24351 nor n24413 n24414 ; n24415
g24352 and a[11] n24415_not ; n24416
g24353 and a[11]_not n24415 ; n24417
g24354 nor n24416 n24417 ; n24418
g24355 and n24407 n24418_not ; n24419
g24356 and n7983 n22384 ; n24420
g24357 and n7291 n22390 ; n24421
g24358 and n7632 n22387 ; n24422
g24359 nor n24421 n24422 ; n24423
g24360 and n24420_not n24423 ; n24424
g24361 and n7294 n22806 ; n24425
g24362 and n24424 n24425_not ; n24426
g24363 and a[11] n24426_not ; n24427
g24364 nor n24426 n24427 ; n24428
g24365 and a[11] n24427_not ; n24429
g24366 nor n24428 n24429 ; n24430
g24367 and n23943 n23945_not ; n24431
g24368 nor n23946 n24431 ; n24432
g24369 and n24430_not n24432 ; n24433
g24370 nor n24430 n24433 ; n24434
g24371 and n24432 n24433_not ; n24435
g24372 nor n24434 n24435 ; n24436
g24373 nor n23930 n23942 ; n24437
g24374 nor n23941 n23942 ; n24438
g24375 nor n24437 n24438 ; n24439
g24376 and n7983 n22387 ; n24440
g24377 and n7291 n22393 ; n24441
g24378 and n7632 n22390 ; n24442
g24379 nor n24441 n24442 ; n24443
g24380 and n24440_not n24443 ; n24444
g24381 and n7294_not n24444 ; n24445
g24382 and n22582_not n24444 ; n24446
g24383 nor n24445 n24446 ; n24447
g24384 and a[11] n24447_not ; n24448
g24385 and a[11]_not n24447 ; n24449
g24386 nor n24448 n24449 ; n24450
g24387 nor n24439 n24450 ; n24451
g24388 and n7983 n22390 ; n24452
g24389 and n7291 n22396 ; n24453
g24390 and n7632 n22393 ; n24454
g24391 nor n24453 n24454 ; n24455
g24392 and n24452_not n24455 ; n24456
g24393 and n7294 n22649 ; n24457
g24394 and n24456 n24457_not ; n24458
g24395 and a[11] n24458_not ; n24459
g24396 nor n24458 n24459 ; n24460
g24397 and a[11] n24459_not ; n24461
g24398 nor n24460 n24461 ; n24462
g24399 and n23914_not n23925 ; n24463
g24400 nor n23926 n24463 ; n24464
g24401 and n24462_not n24464 ; n24465
g24402 nor n24462 n24465 ; n24466
g24403 and n24464 n24465_not ; n24467
g24404 nor n24466 n24467 ; n24468
g24405 and n23911 n23913_not ; n24469
g24406 nor n23914 n24469 ; n24470
g24407 and n7983 n22393 ; n24471
g24408 and n7291 n22399 ; n24472
g24409 and n7632 n22396 ; n24473
g24410 nor n24472 n24473 ; n24474
g24411 and n24471_not n24474 ; n24475
g24412 and n7294_not n24475 ; n24476
g24413 and n22671_not n24475 ; n24477
g24414 nor n24476 n24477 ; n24478
g24415 and a[11] n24478_not ; n24479
g24416 and a[11]_not n24478 ; n24480
g24417 nor n24479 n24480 ; n24481
g24418 and n24470 n24481_not ; n24482
g24419 and n7632 n22406_not ; n24483
g24420 and n7983 n22402 ; n24484
g24421 nor n24483 n24484 ; n24485
g24422 and n7294 n22609_not ; n24486
g24423 and n24485 n24486_not ; n24487
g24424 and a[11] n24487_not ; n24488
g24425 and a[11] n24488_not ; n24489
g24426 nor n24487 n24488 ; n24490
g24427 nor n24489 n24490 ; n24491
g24428 nor n7289 n22406 ; n24492
g24429 and a[11] n24492_not ; n24493
g24430 and n24491_not n24493 ; n24494
g24431 and n7983 n22399 ; n24495
g24432 and n7291 n22406_not ; n24496
g24433 and n7632 n22402 ; n24497
g24434 nor n24496 n24497 ; n24498
g24435 and n24495_not n24498 ; n24499
g24436 and n7294_not n24499 ; n24500
g24437 and n22625 n24499 ; n24501
g24438 nor n24500 n24501 ; n24502
g24439 and a[11] n24502_not ; n24503
g24440 and a[11]_not n24502 ; n24504
g24441 nor n24503 n24504 ; n24505
g24442 and n24494 n24505_not ; n24506
g24443 and n23912 n24506 ; n24507
g24444 and n24506 n24507_not ; n24508
g24445 and n23912 n24507_not ; n24509
g24446 nor n24508 n24509 ; n24510
g24447 and n7983 n22396 ; n24511
g24448 and n7291 n22402 ; n24512
g24449 and n7632 n22399 ; n24513
g24450 nor n24512 n24513 ; n24514
g24451 and n24511_not n24514 ; n24515
g24452 and n7294 n22595 ; n24516
g24453 and n24515 n24516_not ; n24517
g24454 and a[11] n24517_not ; n24518
g24455 and a[11] n24518_not ; n24519
g24456 nor n24517 n24518 ; n24520
g24457 nor n24519 n24520 ; n24521
g24458 nor n24510 n24521 ; n24522
g24459 nor n24507 n24522 ; n24523
g24460 and n24470_not n24481 ; n24524
g24461 nor n24482 n24524 ; n24525
g24462 and n24523_not n24525 ; n24526
g24463 nor n24482 n24526 ; n24527
g24464 nor n24468 n24527 ; n24528
g24465 nor n24465 n24528 ; n24529
g24466 and n24439 n24450 ; n24530
g24467 nor n24451 n24530 ; n24531
g24468 and n24529_not n24531 ; n24532
g24469 nor n24451 n24532 ; n24533
g24470 nor n24436 n24533 ; n24534
g24471 nor n24433 n24534 ; n24535
g24472 and n24407 n24419_not ; n24536
g24473 nor n24418 n24419 ; n24537
g24474 nor n24536 n24537 ; n24538
g24475 nor n24535 n24538 ; n24539
g24476 nor n24419 n24539 ; n24540
g24477 and n24393 n24405_not ; n24541
g24478 nor n24404 n24405 ; n24542
g24479 nor n24541 n24542 ; n24543
g24480 nor n24540 n24543 ; n24544
g24481 nor n24405 n24544 ; n24545
g24482 and n24379_not n24390 ; n24546
g24483 nor n24391 n24546 ; n24547
g24484 and n24545_not n24547 ; n24548
g24485 nor n24391 n24548 ; n24549
g24486 nor n24377 n24549 ; n24550
g24487 nor n24374 n24550 ; n24551
g24488 nor n24359 n24551 ; n24552
g24489 nor n24356 n24552 ; n24553
g24490 nor n24341 n24553 ; n24554
g24491 nor n24338 n24554 ; n24555
g24492 and n24312 n24324_not ; n24556
g24493 nor n24323 n24324 ; n24557
g24494 nor n24556 n24557 ; n24558
g24495 nor n24555 n24558 ; n24559
g24496 nor n24324 n24559 ; n24560
g24497 and n24298 n24310_not ; n24561
g24498 nor n24309 n24310 ; n24562
g24499 nor n24561 n24562 ; n24563
g24500 nor n24560 n24563 ; n24564
g24501 nor n24310 n24564 ; n24565
g24502 and n24284_not n24295 ; n24566
g24503 nor n24296 n24566 ; n24567
g24504 and n24565_not n24567 ; n24568
g24505 nor n24296 n24568 ; n24569
g24506 nor n24282 n24569 ; n24570
g24507 nor n24279 n24570 ; n24571
g24508 nor n24264 n24571 ; n24572
g24509 nor n24261 n24572 ; n24573
g24510 nor n24246 n24573 ; n24574
g24511 nor n24243 n24574 ; n24575
g24512 and n24217 n24229_not ; n24576
g24513 nor n24228 n24229 ; n24577
g24514 nor n24576 n24577 ; n24578
g24515 nor n24575 n24578 ; n24579
g24516 nor n24229 n24579 ; n24580
g24517 and n24203_not n24214 ; n24581
g24518 nor n24215 n24581 ; n24582
g24519 and n24580_not n24582 ; n24583
g24520 nor n24215 n24583 ; n24584
g24521 nor n24201 n24584 ; n24585
g24522 nor n24198 n24585 ; n24586
g24523 nor n24180 n24586 ; n24587
g24524 nor n24177 n24587 ; n24588
g24525 and n24159 n24588 ; n24589
g24526 nor n24159 n24588 ; n24590
g24527 nor n24589 n24590 ; n24591
g24528 and n9331 n22323 ; n24592
g24529 and n8418 n22329 ; n24593
g24530 and n8860 n22326 ; n24594
g24531 nor n24593 n24594 ; n24595
g24532 and n24592_not n24595 ; n24596
g24533 and n8421_not n24596 ; n24597
g24534 and n22504 n22506_not ; n24598
g24535 nor n22507 n24598 ; n24599
g24536 and n24596 n24599_not ; n24600
g24537 nor n24597 n24600 ; n24601
g24538 and a[8] n24601_not ; n24602
g24539 and a[8]_not n24601 ; n24603
g24540 nor n24602 n24603 ; n24604
g24541 and n24591 n24604_not ; n24605
g24542 and n24180 n24586 ; n24606
g24543 nor n24587 n24606 ; n24607
g24544 and n9331 n22326 ; n24608
g24545 and n8418 n22332 ; n24609
g24546 and n8860 n22329 ; n24610
g24547 nor n24609 n24610 ; n24611
g24548 and n24608_not n24611 ; n24612
g24549 and n8421_not n24612 ; n24613
g24550 nor n22500 n22503 ; n24614
g24551 and n22501_not n22504 ; n24615
g24552 nor n24614 n24615 ; n24616
g24553 and n24612 n24616 ; n24617
g24554 nor n24613 n24617 ; n24618
g24555 and a[8] n24618_not ; n24619
g24556 and a[8]_not n24618 ; n24620
g24557 nor n24619 n24620 ; n24621
g24558 and n24607 n24621_not ; n24622
g24559 and n24201 n24584 ; n24623
g24560 nor n24585 n24623 ; n24624
g24561 and n9331 n22329 ; n24625
g24562 and n8418 n22335 ; n24626
g24563 and n8860 n22332 ; n24627
g24564 nor n24626 n24627 ; n24628
g24565 and n24625_not n24628 ; n24629
g24566 and n8421_not n24629 ; n24630
g24567 nor n22496 n22499 ; n24631
g24568 and n22497_not n22500 ; n24632
g24569 nor n24631 n24632 ; n24633
g24570 and n24629 n24633 ; n24634
g24571 nor n24630 n24634 ; n24635
g24572 and a[8] n24635_not ; n24636
g24573 and a[8]_not n24635 ; n24637
g24574 nor n24636 n24637 ; n24638
g24575 and n24624 n24638_not ; n24639
g24576 and n9331 n22332 ; n24640
g24577 and n8418 n22338 ; n24641
g24578 and n8860 n22335 ; n24642
g24579 nor n24641 n24642 ; n24643
g24580 and n24640_not n24643 ; n24644
g24581 and n8421 n22542 ; n24645
g24582 and n24644 n24645_not ; n24646
g24583 and a[8] n24646_not ; n24647
g24584 nor n24646 n24647 ; n24648
g24585 and a[8] n24647_not ; n24649
g24586 nor n24648 n24649 ; n24650
g24587 and n24580 n24582_not ; n24651
g24588 nor n24583 n24651 ; n24652
g24589 and n24650_not n24652 ; n24653
g24590 nor n24650 n24653 ; n24654
g24591 and n24652 n24653_not ; n24655
g24592 nor n24654 n24655 ; n24656
g24593 and n9331 n22335 ; n24657
g24594 and n8418 n22341 ; n24658
g24595 and n8860 n22338 ; n24659
g24596 nor n24658 n24659 ; n24660
g24597 and n24657_not n24660 ; n24661
g24598 and n8421 n24167_not ; n24662
g24599 and n24661 n24662_not ; n24663
g24600 and a[8] n24663_not ; n24664
g24601 nor n24663 n24664 ; n24665
g24602 and a[8] n24664_not ; n24666
g24603 nor n24665 n24666 ; n24667
g24604 nor n24575 n24579 ; n24668
g24605 nor n24578 n24579 ; n24669
g24606 nor n24668 n24669 ; n24670
g24607 nor n24667 n24670 ; n24671
g24608 nor n24667 n24671 ; n24672
g24609 nor n24670 n24671 ; n24673
g24610 nor n24672 n24673 ; n24674
g24611 and n24246 n24573 ; n24675
g24612 nor n24574 n24675 ; n24676
g24613 and n9331 n22338 ; n24677
g24614 and n8418 n22344 ; n24678
g24615 and n8860 n22341 ; n24679
g24616 nor n24678 n24679 ; n24680
g24617 and n24677_not n24680 ; n24681
g24618 and n8421_not n24681 ; n24682
g24619 and n24188 n24681 ; n24683
g24620 nor n24682 n24683 ; n24684
g24621 and a[8] n24684_not ; n24685
g24622 and a[8]_not n24684 ; n24686
g24623 nor n24685 n24686 ; n24687
g24624 and n24676 n24687_not ; n24688
g24625 and n24264 n24571 ; n24689
g24626 nor n24572 n24689 ; n24690
g24627 and n9331 n22341 ; n24691
g24628 and n8418 n22347 ; n24692
g24629 and n8860 n22344 ; n24693
g24630 nor n24692 n24693 ; n24694
g24631 and n24691_not n24694 ; n24695
g24632 and n8421_not n24695 ; n24696
g24633 and n24142_not n24695 ; n24697
g24634 nor n24696 n24697 ; n24698
g24635 and a[8] n24698_not ; n24699
g24636 and a[8]_not n24698 ; n24700
g24637 nor n24699 n24700 ; n24701
g24638 and n24690 n24701_not ; n24702
g24639 and n24282 n24569 ; n24703
g24640 nor n24570 n24703 ; n24704
g24641 and n9331 n22344 ; n24705
g24642 and n8418 n22350 ; n24706
g24643 and n8860 n22347 ; n24707
g24644 nor n24706 n24707 ; n24708
g24645 and n24705_not n24708 ; n24709
g24646 and n8421_not n24709 ; n24710
g24647 and n23642 n24709 ; n24711
g24648 nor n24710 n24711 ; n24712
g24649 and a[8] n24712_not ; n24713
g24650 and a[8]_not n24712 ; n24714
g24651 nor n24713 n24714 ; n24715
g24652 and n24704 n24715_not ; n24716
g24653 and n9331 n22347 ; n24717
g24654 and n8418 n22353 ; n24718
g24655 and n8860 n22350 ; n24719
g24656 nor n24718 n24719 ; n24720
g24657 and n24717_not n24720 ; n24721
g24658 and n8421 n23659_not ; n24722
g24659 and n24721 n24722_not ; n24723
g24660 and a[8] n24723_not ; n24724
g24661 nor n24723 n24724 ; n24725
g24662 and a[8] n24724_not ; n24726
g24663 nor n24725 n24726 ; n24727
g24664 and n24565 n24567_not ; n24728
g24665 nor n24568 n24728 ; n24729
g24666 and n24727_not n24729 ; n24730
g24667 nor n24727 n24730 ; n24731
g24668 and n24729 n24730_not ; n24732
g24669 nor n24731 n24732 ; n24733
g24670 and n9331 n22350 ; n24734
g24671 and n8418 n22356 ; n24735
g24672 and n8860 n22353 ; n24736
g24673 nor n24735 n24736 ; n24737
g24674 and n24734_not n24737 ; n24738
g24675 and n8421 n23672 ; n24739
g24676 and n24738 n24739_not ; n24740
g24677 and a[8] n24740_not ; n24741
g24678 nor n24740 n24741 ; n24742
g24679 and a[8] n24741_not ; n24743
g24680 nor n24742 n24743 ; n24744
g24681 nor n24560 n24564 ; n24745
g24682 nor n24563 n24564 ; n24746
g24683 nor n24745 n24746 ; n24747
g24684 nor n24744 n24747 ; n24748
g24685 nor n24744 n24748 ; n24749
g24686 nor n24747 n24748 ; n24750
g24687 nor n24749 n24750 ; n24751
g24688 and n9331 n22353 ; n24752
g24689 and n8418 n22359 ; n24753
g24690 and n8860 n22356 ; n24754
g24691 nor n24753 n24754 ; n24755
g24692 and n24752_not n24755 ; n24756
g24693 and n8421 n22556_not ; n24757
g24694 and n24756 n24757_not ; n24758
g24695 and a[8] n24758_not ; n24759
g24696 nor n24758 n24759 ; n24760
g24697 and a[8] n24759_not ; n24761
g24698 nor n24760 n24761 ; n24762
g24699 nor n24555 n24559 ; n24763
g24700 nor n24558 n24559 ; n24764
g24701 nor n24763 n24764 ; n24765
g24702 nor n24762 n24765 ; n24766
g24703 nor n24762 n24766 ; n24767
g24704 nor n24765 n24766 ; n24768
g24705 nor n24767 n24768 ; n24769
g24706 and n24341 n24553 ; n24770
g24707 nor n24554 n24770 ; n24771
g24708 and n9331 n22356 ; n24772
g24709 and n8418 n22362 ; n24773
g24710 and n8860 n22359 ; n24774
g24711 nor n24773 n24774 ; n24775
g24712 and n24772_not n24775 ; n24776
g24713 and n8421_not n24776 ; n24777
g24714 and n23345 n24776 ; n24778
g24715 nor n24777 n24778 ; n24779
g24716 and a[8] n24779_not ; n24780
g24717 and a[8]_not n24779 ; n24781
g24718 nor n24780 n24781 ; n24782
g24719 and n24771 n24782_not ; n24783
g24720 and n24359 n24551 ; n24784
g24721 nor n24552 n24784 ; n24785
g24722 and n9331 n22359 ; n24786
g24723 and n8418 n22365 ; n24787
g24724 and n8860 n22362 ; n24788
g24725 nor n24787 n24788 ; n24789
g24726 and n24786_not n24789 ; n24790
g24727 and n8421_not n24790 ; n24791
g24728 and n23368_not n24790 ; n24792
g24729 nor n24791 n24792 ; n24793
g24730 and a[8] n24793_not ; n24794
g24731 and a[8]_not n24793 ; n24795
g24732 nor n24794 n24795 ; n24796
g24733 and n24785 n24796_not ; n24797
g24734 and n24377 n24549 ; n24798
g24735 nor n24550 n24798 ; n24799
g24736 and n9331 n22362 ; n24800
g24737 and n8418 n22368 ; n24801
g24738 and n8860 n22365 ; n24802
g24739 nor n24801 n24802 ; n24803
g24740 and n24800_not n24803 ; n24804
g24741 and n8421_not n24804 ; n24805
g24742 and n23320 n24804 ; n24806
g24743 nor n24805 n24806 ; n24807
g24744 and a[8] n24807_not ; n24808
g24745 and a[8]_not n24807 ; n24809
g24746 nor n24808 n24809 ; n24810
g24747 and n24799 n24810_not ; n24811
g24748 and n9331 n22365 ; n24812
g24749 and n8418 n22371 ; n24813
g24750 and n8860 n22368 ; n24814
g24751 nor n24813 n24814 ; n24815
g24752 and n24812_not n24815 ; n24816
g24753 and n8421 n22993_not ; n24817
g24754 and n24816 n24817_not ; n24818
g24755 and a[8] n24818_not ; n24819
g24756 nor n24818 n24819 ; n24820
g24757 and a[8] n24819_not ; n24821
g24758 nor n24820 n24821 ; n24822
g24759 and n24545 n24547_not ; n24823
g24760 nor n24548 n24823 ; n24824
g24761 and n24822_not n24824 ; n24825
g24762 nor n24822 n24825 ; n24826
g24763 and n24824 n24825_not ; n24827
g24764 nor n24826 n24827 ; n24828
g24765 and n9331 n22368 ; n24829
g24766 and n8418 n22374 ; n24830
g24767 and n8860 n22371 ; n24831
g24768 nor n24830 n24831 ; n24832
g24769 and n24829_not n24832 ; n24833
g24770 and n8421 n23006 ; n24834
g24771 and n24833 n24834_not ; n24835
g24772 and a[8] n24835_not ; n24836
g24773 nor n24835 n24836 ; n24837
g24774 and a[8] n24836_not ; n24838
g24775 nor n24837 n24838 ; n24839
g24776 nor n24540 n24544 ; n24840
g24777 nor n24543 n24544 ; n24841
g24778 nor n24840 n24841 ; n24842
g24779 nor n24839 n24842 ; n24843
g24780 nor n24839 n24843 ; n24844
g24781 nor n24842 n24843 ; n24845
g24782 nor n24844 n24845 ; n24846
g24783 and n9331 n22371 ; n24847
g24784 and n8418 n22377 ; n24848
g24785 and n8860 n22374 ; n24849
g24786 nor n24848 n24849 ; n24850
g24787 and n24847_not n24850 ; n24851
g24788 and n8421 n23025 ; n24852
g24789 and n24851 n24852_not ; n24853
g24790 and a[8] n24853_not ; n24854
g24791 nor n24853 n24854 ; n24855
g24792 and a[8] n24854_not ; n24856
g24793 nor n24855 n24856 ; n24857
g24794 nor n24535 n24539 ; n24858
g24795 nor n24538 n24539 ; n24859
g24796 nor n24858 n24859 ; n24860
g24797 nor n24857 n24860 ; n24861
g24798 nor n24857 n24861 ; n24862
g24799 nor n24860 n24861 ; n24863
g24800 nor n24862 n24863 ; n24864
g24801 and n24436 n24533 ; n24865
g24802 nor n24534 n24865 ; n24866
g24803 and n9331 n22374 ; n24867
g24804 and n8418 n22380 ; n24868
g24805 and n8860 n22377 ; n24869
g24806 nor n24868 n24869 ; n24870
g24807 and n24867_not n24870 ; n24871
g24808 and n8421_not n24871 ; n24872
g24809 and n22569_not n24871 ; n24873
g24810 nor n24872 n24873 ; n24874
g24811 and a[8] n24874_not ; n24875
g24812 and a[8]_not n24874 ; n24876
g24813 nor n24875 n24876 ; n24877
g24814 and n24866 n24877_not ; n24878
g24815 and n24529 n24531_not ; n24879
g24816 nor n24532 n24879 ; n24880
g24817 and n9331 n22377 ; n24881
g24818 and n8418 n22384 ; n24882
g24819 and n8860 n22380 ; n24883
g24820 nor n24882 n24883 ; n24884
g24821 and n24881_not n24884 ; n24885
g24822 and n8421_not n24885 ; n24886
g24823 and n22834 n24885 ; n24887
g24824 nor n24886 n24887 ; n24888
g24825 and a[8] n24888_not ; n24889
g24826 and a[8]_not n24888 ; n24890
g24827 nor n24889 n24890 ; n24891
g24828 and n24880 n24891_not ; n24892
g24829 and n24468 n24527 ; n24893
g24830 nor n24528 n24893 ; n24894
g24831 and n9331 n22380 ; n24895
g24832 and n8418 n22387 ; n24896
g24833 and n8860 n22384 ; n24897
g24834 nor n24896 n24897 ; n24898
g24835 and n24895_not n24898 ; n24899
g24836 and n8421_not n24899 ; n24900
g24837 and n22850_not n24899 ; n24901
g24838 nor n24900 n24901 ; n24902
g24839 and a[8] n24902_not ; n24903
g24840 and a[8]_not n24902 ; n24904
g24841 nor n24903 n24904 ; n24905
g24842 and n24894 n24905_not ; n24906
g24843 and n9331 n22384 ; n24907
g24844 and n8418 n22390 ; n24908
g24845 and n8860 n22387 ; n24909
g24846 nor n24908 n24909 ; n24910
g24847 and n24907_not n24910 ; n24911
g24848 and n8421 n22806 ; n24912
g24849 and n24911 n24912_not ; n24913
g24850 and a[8] n24913_not ; n24914
g24851 nor n24913 n24914 ; n24915
g24852 and a[8] n24914_not ; n24916
g24853 nor n24915 n24916 ; n24917
g24854 and n24523 n24525_not ; n24918
g24855 nor n24526 n24918 ; n24919
g24856 and n24917_not n24919 ; n24920
g24857 nor n24917 n24920 ; n24921
g24858 and n24919 n24920_not ; n24922
g24859 nor n24921 n24922 ; n24923
g24860 nor n24510 n24522 ; n24924
g24861 nor n24521 n24522 ; n24925
g24862 nor n24924 n24925 ; n24926
g24863 and n9331 n22387 ; n24927
g24864 and n8418 n22393 ; n24928
g24865 and n8860 n22390 ; n24929
g24866 nor n24928 n24929 ; n24930
g24867 and n24927_not n24930 ; n24931
g24868 and n8421_not n24931 ; n24932
g24869 and n22582_not n24931 ; n24933
g24870 nor n24932 n24933 ; n24934
g24871 and a[8] n24934_not ; n24935
g24872 and a[8]_not n24934 ; n24936
g24873 nor n24935 n24936 ; n24937
g24874 nor n24926 n24937 ; n24938
g24875 and n9331 n22390 ; n24939
g24876 and n8418 n22396 ; n24940
g24877 and n8860 n22393 ; n24941
g24878 nor n24940 n24941 ; n24942
g24879 and n24939_not n24942 ; n24943
g24880 and n8421 n22649 ; n24944
g24881 and n24943 n24944_not ; n24945
g24882 and a[8] n24945_not ; n24946
g24883 nor n24945 n24946 ; n24947
g24884 and a[8] n24946_not ; n24948
g24885 nor n24947 n24948 ; n24949
g24886 and n24494_not n24505 ; n24950
g24887 nor n24506 n24950 ; n24951
g24888 and n24949_not n24951 ; n24952
g24889 nor n24949 n24952 ; n24953
g24890 and n24951 n24952_not ; n24954
g24891 nor n24953 n24954 ; n24955
g24892 and n24491 n24493_not ; n24956
g24893 nor n24494 n24956 ; n24957
g24894 and n9331 n22393 ; n24958
g24895 and n8418 n22399 ; n24959
g24896 and n8860 n22396 ; n24960
g24897 nor n24959 n24960 ; n24961
g24898 and n24958_not n24961 ; n24962
g24899 and n8421_not n24962 ; n24963
g24900 and n22671_not n24962 ; n24964
g24901 nor n24963 n24964 ; n24965
g24902 and a[8] n24965_not ; n24966
g24903 and a[8]_not n24965 ; n24967
g24904 nor n24966 n24967 ; n24968
g24905 and n24957 n24968_not ; n24969
g24906 and n8860 n22406_not ; n24970
g24907 and n9331 n22402 ; n24971
g24908 nor n24970 n24971 ; n24972
g24909 and n8421 n22609_not ; n24973
g24910 and n24972 n24973_not ; n24974
g24911 and a[8] n24974_not ; n24975
g24912 and a[8] n24975_not ; n24976
g24913 nor n24974 n24975 ; n24977
g24914 nor n24976 n24977 ; n24978
g24915 nor n8416 n22406 ; n24979
g24916 and a[8] n24979_not ; n24980
g24917 and n24978_not n24980 ; n24981
g24918 and n9331 n22399 ; n24982
g24919 and n8418 n22406_not ; n24983
g24920 and n8860 n22402 ; n24984
g24921 nor n24983 n24984 ; n24985
g24922 and n24982_not n24985 ; n24986
g24923 and n8421_not n24986 ; n24987
g24924 and n22625 n24986 ; n24988
g24925 nor n24987 n24988 ; n24989
g24926 and a[8] n24989_not ; n24990
g24927 and a[8]_not n24989 ; n24991
g24928 nor n24990 n24991 ; n24992
g24929 and n24981 n24992_not ; n24993
g24930 and n24492 n24993 ; n24994
g24931 and n24993 n24994_not ; n24995
g24932 and n24492 n24994_not ; n24996
g24933 nor n24995 n24996 ; n24997
g24934 and n9331 n22396 ; n24998
g24935 and n8418 n22402 ; n24999
g24936 and n8860 n22399 ; n25000
g24937 nor n24999 n25000 ; n25001
g24938 and n24998_not n25001 ; n25002
g24939 and n8421 n22595 ; n25003
g24940 and n25002 n25003_not ; n25004
g24941 and a[8] n25004_not ; n25005
g24942 and a[8] n25005_not ; n25006
g24943 nor n25004 n25005 ; n25007
g24944 nor n25006 n25007 ; n25008
g24945 nor n24997 n25008 ; n25009
g24946 nor n24994 n25009 ; n25010
g24947 and n24957_not n24968 ; n25011
g24948 nor n24969 n25011 ; n25012
g24949 and n25010_not n25012 ; n25013
g24950 nor n24969 n25013 ; n25014
g24951 nor n24955 n25014 ; n25015
g24952 nor n24952 n25015 ; n25016
g24953 and n24926 n24937 ; n25017
g24954 nor n24938 n25017 ; n25018
g24955 and n25016_not n25018 ; n25019
g24956 nor n24938 n25019 ; n25020
g24957 nor n24923 n25020 ; n25021
g24958 nor n24920 n25021 ; n25022
g24959 and n24894 n24906_not ; n25023
g24960 nor n24905 n24906 ; n25024
g24961 nor n25023 n25024 ; n25025
g24962 nor n25022 n25025 ; n25026
g24963 nor n24906 n25026 ; n25027
g24964 and n24880 n24892_not ; n25028
g24965 nor n24891 n24892 ; n25029
g24966 nor n25028 n25029 ; n25030
g24967 nor n25027 n25030 ; n25031
g24968 nor n24892 n25031 ; n25032
g24969 and n24866_not n24877 ; n25033
g24970 nor n24878 n25033 ; n25034
g24971 and n25032_not n25034 ; n25035
g24972 nor n24878 n25035 ; n25036
g24973 nor n24864 n25036 ; n25037
g24974 nor n24861 n25037 ; n25038
g24975 nor n24846 n25038 ; n25039
g24976 nor n24843 n25039 ; n25040
g24977 nor n24828 n25040 ; n25041
g24978 nor n24825 n25041 ; n25042
g24979 and n24799 n24811_not ; n25043
g24980 nor n24810 n24811 ; n25044
g24981 nor n25043 n25044 ; n25045
g24982 nor n25042 n25045 ; n25046
g24983 nor n24811 n25046 ; n25047
g24984 and n24785 n24797_not ; n25048
g24985 nor n24796 n24797 ; n25049
g24986 nor n25048 n25049 ; n25050
g24987 nor n25047 n25050 ; n25051
g24988 nor n24797 n25051 ; n25052
g24989 and n24771_not n24782 ; n25053
g24990 nor n24783 n25053 ; n25054
g24991 and n25052_not n25054 ; n25055
g24992 nor n24783 n25055 ; n25056
g24993 nor n24769 n25056 ; n25057
g24994 nor n24766 n25057 ; n25058
g24995 nor n24751 n25058 ; n25059
g24996 nor n24748 n25059 ; n25060
g24997 nor n24733 n25060 ; n25061
g24998 nor n24730 n25061 ; n25062
g24999 and n24704 n24716_not ; n25063
g25000 nor n24715 n24716 ; n25064
g25001 nor n25063 n25064 ; n25065
g25002 nor n25062 n25065 ; n25066
g25003 nor n24716 n25066 ; n25067
g25004 and n24690 n24702_not ; n25068
g25005 nor n24701 n24702 ; n25069
g25006 nor n25068 n25069 ; n25070
g25007 nor n25067 n25070 ; n25071
g25008 nor n24702 n25071 ; n25072
g25009 and n24676_not n24687 ; n25073
g25010 nor n24688 n25073 ; n25074
g25011 and n25072_not n25074 ; n25075
g25012 nor n24688 n25075 ; n25076
g25013 nor n24674 n25076 ; n25077
g25014 nor n24671 n25077 ; n25078
g25015 nor n24656 n25078 ; n25079
g25016 nor n24653 n25079 ; n25080
g25017 and n24624 n24639_not ; n25081
g25018 nor n24638 n24639 ; n25082
g25019 nor n25081 n25082 ; n25083
g25020 nor n25080 n25083 ; n25084
g25021 nor n24639 n25084 ; n25085
g25022 and n24607 n24622_not ; n25086
g25023 nor n24621 n24622 ; n25087
g25024 nor n25086 n25087 ; n25088
g25025 nor n25085 n25088 ; n25089
g25026 nor n24622 n25089 ; n25090
g25027 and n24591 n24605_not ; n25091
g25028 nor n24604 n24605 ; n25092
g25029 nor n25091 n25092 ; n25093
g25030 nor n25090 n25093 ; n25094
g25031 nor n24605 n25094 ; n25095
g25032 and n7983 n22329 ; n25096
g25033 and n7291 n22335 ; n25097
g25034 and n7632 n22332 ; n25098
g25035 nor n25097 n25098 ; n25099
g25036 and n25096_not n25099 ; n25100
g25037 and n7294 n24633_not ; n25101
g25038 and n25100 n25101_not ; n25102
g25039 and a[11] n25102_not ; n25103
g25040 nor n25102 n25103 ; n25104
g25041 and a[11] n25103_not ; n25105
g25042 nor n25104 n25105 ; n25106
g25043 nor n24148 n24152 ; n25107
g25044 and n6233 n22347 ; n25108
g25045 and n5663 n22353 ; n25109
g25046 and n5939 n22350 ; n25110
g25047 nor n25109 n25110 ; n25111
g25048 and n25108_not n25111 ; n25112
g25049 and n5666 n23659_not ; n25113
g25050 and n25112 n25113_not ; n25114
g25051 and a[17] n25114_not ; n25115
g25052 nor n25114 n25115 ; n25116
g25053 and a[17] n25115_not ; n25117
g25054 nor n25116 n25117 ; n25118
g25055 nor n24119 n24123 ; n25119
g25056 and n4694 n22365 ; n25120
g25057 and n4533 n22371 ; n25121
g25058 and n4604 n22368 ; n25122
g25059 nor n25121 n25122 ; n25123
g25060 and n25120_not n25123 ; n25124
g25061 and n4536 n22993_not ; n25125
g25062 and n25124 n25125_not ; n25126
g25063 and a[23] n25126_not ; n25127
g25064 nor n25126 n25127 ; n25128
g25065 and a[23] n25127_not ; n25129
g25066 nor n25128 n25129 ; n25130
g25067 nor n24092 n24096 ; n25131
g25068 and n3457 n22384 ; n25132
g25069 and n3542 n22390 ; n25133
g25070 and n3606 n22387 ; n25134
g25071 nor n25133 n25134 ; n25135
g25072 and n25132_not n25135 ; n25136
g25073 and n3368 n22806 ; n25137
g25074 and n25136 n25137_not ; n25138
g25075 and a[29] n25138_not ; n25139
g25076 nor n25138 n25139 ; n25140
g25077 and a[29] n25139_not ; n25141
g25078 nor n25140 n25141 ; n25142
g25079 nor n24065 n24069 ; n25143
g25080 and n1611 n5748 ; n25144
g25081 and n4269 n25144 ; n25145
g25082 and n691 n25145 ; n25146
g25083 and n204 n25146 ; n25147
g25084 and n13560 n25147 ; n25148
g25085 and n12932 n25148 ; n25149
g25086 and n12909 n25149 ; n25150
g25087 and n15924 n25150 ; n25151
g25088 and n515 n25151 ; n25152
g25089 and n278_not n25152 ; n25153
g25090 and n135_not n25153 ; n25154
g25091 and n568_not n25154 ; n25155
g25092 and n331_not n25155 ; n25156
g25093 and n225_not n25156 ; n25157
g25094 and n3020 n22393 ; n25158
g25095 and n3028 n22396 ; n25159
g25096 and n3023 n22399 ; n25160
g25097 and n75 n22671 ; n25161
g25098 nor n25160 n25161 ; n25162
g25099 and n25159_not n25162 ; n25163
g25100 and n25158_not n25163 ; n25164
g25101 nor n25157 n25164 ; n25165
g25102 nor n25157 n25165 ; n25166
g25103 nor n25164 n25165 ; n25167
g25104 nor n25166 n25167 ; n25168
g25105 nor n25143 n25168 ; n25169
g25106 nor n25143 n25169 ; n25170
g25107 nor n25168 n25169 ; n25171
g25108 nor n25170 n25171 ; n25172
g25109 nor n25142 n25172 ; n25173
g25110 nor n25142 n25173 ; n25174
g25111 nor n25172 n25173 ; n25175
g25112 nor n25174 n25175 ; n25176
g25113 nor n24073 n24079 ; n25177
g25114 and n25176 n25177 ; n25178
g25115 nor n25176 n25177 ; n25179
g25116 nor n25178 n25179 ; n25180
g25117 and n3884 n22374 ; n25181
g25118 and n3967 n22380 ; n25182
g25119 and n4046 n22377 ; n25183
g25120 nor n25182 n25183 ; n25184
g25121 and n25181_not n25184 ; n25185
g25122 and n4050_not n25185 ; n25186
g25123 and n22569_not n25185 ; n25187
g25124 nor n25186 n25187 ; n25188
g25125 and a[26] n25188_not ; n25189
g25126 and a[26]_not n25188 ; n25190
g25127 nor n25189 n25190 ; n25191
g25128 and n25180 n25191_not ; n25192
g25129 and n25180 n25192_not ; n25193
g25130 nor n25191 n25192 ; n25194
g25131 nor n25193 n25194 ; n25195
g25132 nor n25131 n25195 ; n25196
g25133 nor n25131 n25196 ; n25197
g25134 nor n25195 n25196 ; n25198
g25135 nor n25197 n25198 ; n25199
g25136 nor n25130 n25199 ; n25200
g25137 nor n25130 n25200 ; n25201
g25138 nor n25199 n25200 ; n25202
g25139 nor n25201 n25202 ; n25203
g25140 nor n24100 n24106 ; n25204
g25141 and n25203 n25204 ; n25205
g25142 nor n25203 n25204 ; n25206
g25143 nor n25205 n25206 ; n25207
g25144 and n5496 n22356 ; n25208
g25145 and n4935 n22362 ; n25209
g25146 and n5407 n22359 ; n25210
g25147 nor n25209 n25210 ; n25211
g25148 and n25208_not n25211 ; n25212
g25149 and n4938_not n25212 ; n25213
g25150 and n23345 n25212 ; n25214
g25151 nor n25213 n25214 ; n25215
g25152 and a[20] n25215_not ; n25216
g25153 and a[20]_not n25215 ; n25217
g25154 nor n25216 n25217 ; n25218
g25155 and n25207 n25218_not ; n25219
g25156 and n25207 n25219_not ; n25220
g25157 nor n25218 n25219 ; n25221
g25158 nor n25220 n25221 ; n25222
g25159 nor n25119 n25222 ; n25223
g25160 nor n25119 n25223 ; n25224
g25161 nor n25222 n25223 ; n25225
g25162 nor n25224 n25225 ; n25226
g25163 nor n25118 n25226 ; n25227
g25164 nor n25118 n25227 ; n25228
g25165 nor n25226 n25227 ; n25229
g25166 nor n25228 n25229 ; n25230
g25167 nor n24127 n24133 ; n25231
g25168 and n25230 n25231 ; n25232
g25169 nor n25230 n25231 ; n25233
g25170 nor n25232 n25233 ; n25234
g25171 and n7101 n22338 ; n25235
g25172 and n6402 n22344 ; n25236
g25173 and n6951 n22341 ; n25237
g25174 nor n25236 n25237 ; n25238
g25175 and n25235_not n25238 ; n25239
g25176 and n6397_not n25239 ; n25240
g25177 and n24188 n25239 ; n25241
g25178 nor n25240 n25241 ; n25242
g25179 and a[14] n25242_not ; n25243
g25180 and a[14]_not n25242 ; n25244
g25181 nor n25243 n25244 ; n25245
g25182 and n25234 n25245_not ; n25246
g25183 and n25234 n25246_not ; n25247
g25184 nor n25245 n25246 ; n25248
g25185 nor n25247 n25248 ; n25249
g25186 nor n25107 n25249 ; n25250
g25187 nor n25107 n25250 ; n25251
g25188 nor n25249 n25250 ; n25252
g25189 nor n25251 n25252 ; n25253
g25190 nor n25106 n25253 ; n25254
g25191 nor n25106 n25254 ; n25255
g25192 nor n25253 n25254 ; n25256
g25193 nor n25255 n25256 ; n25257
g25194 nor n24156 n24590 ; n25258
g25195 and n25257 n25258 ; n25259
g25196 nor n25257 n25258 ; n25260
g25197 nor n25259 n25260 ; n25261
g25198 and n9331 n22320 ; n25262
g25199 and n8418 n22326 ; n25263
g25200 and n8860 n22323 ; n25264
g25201 nor n25263 n25264 ; n25265
g25202 and n25262_not n25265 ; n25266
g25203 and n8421_not n25266 ; n25267
g25204 nor n22508 n22511 ; n25268
g25205 and n22509_not n22512 ; n25269
g25206 nor n25268 n25269 ; n25270
g25207 and n25266 n25270 ; n25271
g25208 nor n25267 n25271 ; n25272
g25209 and a[8] n25272_not ; n25273
g25210 and a[8]_not n25272 ; n25274
g25211 nor n25273 n25274 ; n25275
g25212 and n25261 n25275_not ; n25276
g25213 and n25261 n25276_not ; n25277
g25214 nor n25275 n25276 ; n25278
g25215 nor n25277 n25278 ; n25279
g25216 nor n25095 n25279 ; n25280
g25217 nor n25095 n25280 ; n25281
g25218 nor n25279 n25280 ; n25282
g25219 nor n25281 n25282 ; n25283
g25220 nor n22535 n25283 ; n25284
g25221 nor n22535 n25284 ; n25285
g25222 nor n25283 n25284 ; n25286
g25223 nor n25285 n25286 ; n25287
g25224 and n71 n22315 ; n25288
g25225 and n9867 n22320 ; n25289
g25226 and n10434 n22312 ; n25290
g25227 nor n25289 n25290 ; n25291
g25228 and n25288_not n25291 ; n25292
g25229 and n22516 n22519_not ; n25293
g25230 nor n22520 n25293 ; n25294
g25231 and n9870 n25294 ; n25295
g25232 and n25292 n25295_not ; n25296
g25233 and a[5] n25296_not ; n25297
g25234 nor n25296 n25297 ; n25298
g25235 and a[5] n25297_not ; n25299
g25236 nor n25298 n25299 ; n25300
g25237 nor n25090 n25094 ; n25301
g25238 nor n25093 n25094 ; n25302
g25239 nor n25301 n25302 ; n25303
g25240 nor n25300 n25303 ; n25304
g25241 nor n25300 n25304 ; n25305
g25242 nor n25303 n25304 ; n25306
g25243 nor n25305 n25306 ; n25307
g25244 and n71 n22312 ; n25308
g25245 and n9867 n22323 ; n25309
g25246 and n10434 n22320 ; n25310
g25247 nor n25309 n25310 ; n25311
g25248 and n25308_not n25311 ; n25312
g25249 nor n22512 n22515 ; n25313
g25250 and n22513_not n22516 ; n25314
g25251 nor n25313 n25314 ; n25315
g25252 and n9870 n25315_not ; n25316
g25253 and n25312 n25316_not ; n25317
g25254 and a[5] n25317_not ; n25318
g25255 nor n25317 n25318 ; n25319
g25256 and a[5] n25318_not ; n25320
g25257 nor n25319 n25320 ; n25321
g25258 nor n25085 n25089 ; n25322
g25259 nor n25088 n25089 ; n25323
g25260 nor n25322 n25323 ; n25324
g25261 nor n25321 n25324 ; n25325
g25262 nor n25321 n25325 ; n25326
g25263 nor n25324 n25325 ; n25327
g25264 nor n25326 n25327 ; n25328
g25265 and n71 n22320 ; n25329
g25266 and n9867 n22326 ; n25330
g25267 and n10434 n22323 ; n25331
g25268 nor n25330 n25331 ; n25332
g25269 and n25329_not n25332 ; n25333
g25270 and n9870 n25270_not ; n25334
g25271 and n25333 n25334_not ; n25335
g25272 and a[5] n25335_not ; n25336
g25273 nor n25335 n25336 ; n25337
g25274 and a[5] n25336_not ; n25338
g25275 nor n25337 n25338 ; n25339
g25276 nor n25080 n25084 ; n25340
g25277 nor n25083 n25084 ; n25341
g25278 nor n25340 n25341 ; n25342
g25279 nor n25339 n25342 ; n25343
g25280 nor n25339 n25343 ; n25344
g25281 nor n25342 n25343 ; n25345
g25282 nor n25344 n25345 ; n25346
g25283 and n24656 n25078 ; n25347
g25284 nor n25079 n25347 ; n25348
g25285 and n71 n22323 ; n25349
g25286 and n9867 n22329 ; n25350
g25287 and n10434 n22326 ; n25351
g25288 nor n25350 n25351 ; n25352
g25289 and n25349_not n25352 ; n25353
g25290 and n9870_not n25353 ; n25354
g25291 and n24599_not n25353 ; n25355
g25292 nor n25354 n25355 ; n25356
g25293 and a[5] n25356_not ; n25357
g25294 and a[5]_not n25356 ; n25358
g25295 nor n25357 n25358 ; n25359
g25296 and n25348 n25359_not ; n25360
g25297 and n24674 n25076 ; n25361
g25298 nor n25077 n25361 ; n25362
g25299 and n71 n22326 ; n25363
g25300 and n9867 n22332 ; n25364
g25301 and n10434 n22329 ; n25365
g25302 nor n25364 n25365 ; n25366
g25303 and n25363_not n25366 ; n25367
g25304 and n9870_not n25367 ; n25368
g25305 and n24616 n25367 ; n25369
g25306 nor n25368 n25369 ; n25370
g25307 and a[5] n25370_not ; n25371
g25308 and a[5]_not n25370 ; n25372
g25309 nor n25371 n25372 ; n25373
g25310 and n25362 n25373_not ; n25374
g25311 and n71 n22329 ; n25375
g25312 and n9867 n22335 ; n25376
g25313 and n10434 n22332 ; n25377
g25314 nor n25376 n25377 ; n25378
g25315 and n25375_not n25378 ; n25379
g25316 and n9870 n24633_not ; n25380
g25317 and n25379 n25380_not ; n25381
g25318 and a[5] n25381_not ; n25382
g25319 nor n25381 n25382 ; n25383
g25320 and a[5] n25382_not ; n25384
g25321 nor n25383 n25384 ; n25385
g25322 and n25072 n25074_not ; n25386
g25323 nor n25075 n25386 ; n25387
g25324 and n25385_not n25387 ; n25388
g25325 nor n25385 n25388 ; n25389
g25326 and n25387 n25388_not ; n25390
g25327 nor n25389 n25390 ; n25391
g25328 and n71 n22332 ; n25392
g25329 and n9867 n22338 ; n25393
g25330 and n10434 n22335 ; n25394
g25331 nor n25393 n25394 ; n25395
g25332 and n25392_not n25395 ; n25396
g25333 and n9870 n22542 ; n25397
g25334 and n25396 n25397_not ; n25398
g25335 and a[5] n25398_not ; n25399
g25336 nor n25398 n25399 ; n25400
g25337 and a[5] n25399_not ; n25401
g25338 nor n25400 n25401 ; n25402
g25339 nor n25067 n25071 ; n25403
g25340 nor n25070 n25071 ; n25404
g25341 nor n25403 n25404 ; n25405
g25342 nor n25402 n25405 ; n25406
g25343 nor n25402 n25406 ; n25407
g25344 nor n25405 n25406 ; n25408
g25345 nor n25407 n25408 ; n25409
g25346 and n71 n22335 ; n25410
g25347 and n9867 n22341 ; n25411
g25348 and n10434 n22338 ; n25412
g25349 nor n25411 n25412 ; n25413
g25350 and n25410_not n25413 ; n25414
g25351 and n9870 n24167_not ; n25415
g25352 and n25414 n25415_not ; n25416
g25353 and a[5] n25416_not ; n25417
g25354 nor n25416 n25417 ; n25418
g25355 and a[5] n25417_not ; n25419
g25356 nor n25418 n25419 ; n25420
g25357 nor n25062 n25066 ; n25421
g25358 nor n25065 n25066 ; n25422
g25359 nor n25421 n25422 ; n25423
g25360 nor n25420 n25423 ; n25424
g25361 nor n25420 n25424 ; n25425
g25362 nor n25423 n25424 ; n25426
g25363 nor n25425 n25426 ; n25427
g25364 and n24733 n25060 ; n25428
g25365 nor n25061 n25428 ; n25429
g25366 and n71 n22338 ; n25430
g25367 and n9867 n22344 ; n25431
g25368 and n10434 n22341 ; n25432
g25369 nor n25431 n25432 ; n25433
g25370 and n25430_not n25433 ; n25434
g25371 and n9870_not n25434 ; n25435
g25372 and n24188 n25434 ; n25436
g25373 nor n25435 n25436 ; n25437
g25374 and a[5] n25437_not ; n25438
g25375 and a[5]_not n25437 ; n25439
g25376 nor n25438 n25439 ; n25440
g25377 and n25429 n25440_not ; n25441
g25378 and n24751 n25058 ; n25442
g25379 nor n25059 n25442 ; n25443
g25380 and n71 n22341 ; n25444
g25381 and n9867 n22347 ; n25445
g25382 and n10434 n22344 ; n25446
g25383 nor n25445 n25446 ; n25447
g25384 and n25444_not n25447 ; n25448
g25385 and n9870_not n25448 ; n25449
g25386 and n24142_not n25448 ; n25450
g25387 nor n25449 n25450 ; n25451
g25388 and a[5] n25451_not ; n25452
g25389 and a[5]_not n25451 ; n25453
g25390 nor n25452 n25453 ; n25454
g25391 and n25443 n25454_not ; n25455
g25392 and n24769 n25056 ; n25456
g25393 nor n25057 n25456 ; n25457
g25394 and n71 n22344 ; n25458
g25395 and n9867 n22350 ; n25459
g25396 and n10434 n22347 ; n25460
g25397 nor n25459 n25460 ; n25461
g25398 and n25458_not n25461 ; n25462
g25399 and n9870_not n25462 ; n25463
g25400 and n23642 n25462 ; n25464
g25401 nor n25463 n25464 ; n25465
g25402 and a[5] n25465_not ; n25466
g25403 and a[5]_not n25465 ; n25467
g25404 nor n25466 n25467 ; n25468
g25405 and n25457 n25468_not ; n25469
g25406 and n71 n22347 ; n25470
g25407 and n9867 n22353 ; n25471
g25408 and n10434 n22350 ; n25472
g25409 nor n25471 n25472 ; n25473
g25410 and n25470_not n25473 ; n25474
g25411 and n9870 n23659_not ; n25475
g25412 and n25474 n25475_not ; n25476
g25413 and a[5] n25476_not ; n25477
g25414 nor n25476 n25477 ; n25478
g25415 and a[5] n25477_not ; n25479
g25416 nor n25478 n25479 ; n25480
g25417 and n25052 n25054_not ; n25481
g25418 nor n25055 n25481 ; n25482
g25419 and n25480_not n25482 ; n25483
g25420 nor n25480 n25483 ; n25484
g25421 and n25482 n25483_not ; n25485
g25422 nor n25484 n25485 ; n25486
g25423 and n71 n22350 ; n25487
g25424 and n9867 n22356 ; n25488
g25425 and n10434 n22353 ; n25489
g25426 nor n25488 n25489 ; n25490
g25427 and n25487_not n25490 ; n25491
g25428 and n9870 n23672 ; n25492
g25429 and n25491 n25492_not ; n25493
g25430 and a[5] n25493_not ; n25494
g25431 nor n25493 n25494 ; n25495
g25432 and a[5] n25494_not ; n25496
g25433 nor n25495 n25496 ; n25497
g25434 nor n25047 n25051 ; n25498
g25435 nor n25050 n25051 ; n25499
g25436 nor n25498 n25499 ; n25500
g25437 nor n25497 n25500 ; n25501
g25438 nor n25497 n25501 ; n25502
g25439 nor n25500 n25501 ; n25503
g25440 nor n25502 n25503 ; n25504
g25441 and n71 n22353 ; n25505
g25442 and n9867 n22359 ; n25506
g25443 and n10434 n22356 ; n25507
g25444 nor n25506 n25507 ; n25508
g25445 and n25505_not n25508 ; n25509
g25446 and n9870 n22556_not ; n25510
g25447 and n25509 n25510_not ; n25511
g25448 and a[5] n25511_not ; n25512
g25449 nor n25511 n25512 ; n25513
g25450 and a[5] n25512_not ; n25514
g25451 nor n25513 n25514 ; n25515
g25452 nor n25042 n25046 ; n25516
g25453 nor n25045 n25046 ; n25517
g25454 nor n25516 n25517 ; n25518
g25455 nor n25515 n25518 ; n25519
g25456 nor n25515 n25519 ; n25520
g25457 nor n25518 n25519 ; n25521
g25458 nor n25520 n25521 ; n25522
g25459 and n24828 n25040 ; n25523
g25460 nor n25041 n25523 ; n25524
g25461 and n71 n22356 ; n25525
g25462 and n9867 n22362 ; n25526
g25463 and n10434 n22359 ; n25527
g25464 nor n25526 n25527 ; n25528
g25465 and n25525_not n25528 ; n25529
g25466 and n9870_not n25529 ; n25530
g25467 and n23345 n25529 ; n25531
g25468 nor n25530 n25531 ; n25532
g25469 and a[5] n25532_not ; n25533
g25470 and a[5]_not n25532 ; n25534
g25471 nor n25533 n25534 ; n25535
g25472 and n25524 n25535_not ; n25536
g25473 and n24846 n25038 ; n25537
g25474 nor n25039 n25537 ; n25538
g25475 and n71 n22359 ; n25539
g25476 and n9867 n22365 ; n25540
g25477 and n10434 n22362 ; n25541
g25478 nor n25540 n25541 ; n25542
g25479 and n25539_not n25542 ; n25543
g25480 and n9870_not n25543 ; n25544
g25481 and n23368_not n25543 ; n25545
g25482 nor n25544 n25545 ; n25546
g25483 and a[5] n25546_not ; n25547
g25484 and a[5]_not n25546 ; n25548
g25485 nor n25547 n25548 ; n25549
g25486 and n25538 n25549_not ; n25550
g25487 and n24864 n25036 ; n25551
g25488 nor n25037 n25551 ; n25552
g25489 and n71 n22362 ; n25553
g25490 and n9867 n22368 ; n25554
g25491 and n10434 n22365 ; n25555
g25492 nor n25554 n25555 ; n25556
g25493 and n25553_not n25556 ; n25557
g25494 and n9870_not n25557 ; n25558
g25495 and n23320 n25557 ; n25559
g25496 nor n25558 n25559 ; n25560
g25497 and a[5] n25560_not ; n25561
g25498 and a[5]_not n25560 ; n25562
g25499 nor n25561 n25562 ; n25563
g25500 and n25552 n25563_not ; n25564
g25501 and n71 n22365 ; n25565
g25502 and n9867 n22371 ; n25566
g25503 and n10434 n22368 ; n25567
g25504 nor n25566 n25567 ; n25568
g25505 and n25565_not n25568 ; n25569
g25506 and n9870 n22993_not ; n25570
g25507 and n25569 n25570_not ; n25571
g25508 and a[5] n25571_not ; n25572
g25509 nor n25571 n25572 ; n25573
g25510 and a[5] n25572_not ; n25574
g25511 nor n25573 n25574 ; n25575
g25512 and n25032 n25034_not ; n25576
g25513 nor n25035 n25576 ; n25577
g25514 and n25575_not n25577 ; n25578
g25515 nor n25575 n25578 ; n25579
g25516 and n25577 n25578_not ; n25580
g25517 nor n25579 n25580 ; n25581
g25518 and n71 n22368 ; n25582
g25519 and n9867 n22374 ; n25583
g25520 and n10434 n22371 ; n25584
g25521 nor n25583 n25584 ; n25585
g25522 and n25582_not n25585 ; n25586
g25523 and n9870 n23006 ; n25587
g25524 and n25586 n25587_not ; n25588
g25525 and a[5] n25588_not ; n25589
g25526 nor n25588 n25589 ; n25590
g25527 and a[5] n25589_not ; n25591
g25528 nor n25590 n25591 ; n25592
g25529 nor n25027 n25031 ; n25593
g25530 nor n25030 n25031 ; n25594
g25531 nor n25593 n25594 ; n25595
g25532 nor n25592 n25595 ; n25596
g25533 nor n25592 n25596 ; n25597
g25534 nor n25595 n25596 ; n25598
g25535 nor n25597 n25598 ; n25599
g25536 and n71 n22371 ; n25600
g25537 and n9867 n22377 ; n25601
g25538 and n10434 n22374 ; n25602
g25539 nor n25601 n25602 ; n25603
g25540 and n25600_not n25603 ; n25604
g25541 and n9870 n23025 ; n25605
g25542 and n25604 n25605_not ; n25606
g25543 and a[5] n25606_not ; n25607
g25544 nor n25606 n25607 ; n25608
g25545 and a[5] n25607_not ; n25609
g25546 nor n25608 n25609 ; n25610
g25547 nor n25022 n25026 ; n25611
g25548 nor n25025 n25026 ; n25612
g25549 nor n25611 n25612 ; n25613
g25550 nor n25610 n25613 ; n25614
g25551 nor n25610 n25614 ; n25615
g25552 nor n25613 n25614 ; n25616
g25553 nor n25615 n25616 ; n25617
g25554 and n24923 n25020 ; n25618
g25555 nor n25021 n25618 ; n25619
g25556 and n71 n22374 ; n25620
g25557 and n9867 n22380 ; n25621
g25558 and n10434 n22377 ; n25622
g25559 nor n25621 n25622 ; n25623
g25560 and n25620_not n25623 ; n25624
g25561 and n9870_not n25624 ; n25625
g25562 and n22569_not n25624 ; n25626
g25563 nor n25625 n25626 ; n25627
g25564 and a[5] n25627_not ; n25628
g25565 and a[5]_not n25627 ; n25629
g25566 nor n25628 n25629 ; n25630
g25567 and n25619 n25630_not ; n25631
g25568 and n25016 n25018_not ; n25632
g25569 nor n25019 n25632 ; n25633
g25570 and n71 n22377 ; n25634
g25571 and n9867 n22384 ; n25635
g25572 and n10434 n22380 ; n25636
g25573 nor n25635 n25636 ; n25637
g25574 and n25634_not n25637 ; n25638
g25575 and n9870_not n25638 ; n25639
g25576 and n22834 n25638 ; n25640
g25577 nor n25639 n25640 ; n25641
g25578 and a[5] n25641_not ; n25642
g25579 and a[5]_not n25641 ; n25643
g25580 nor n25642 n25643 ; n25644
g25581 and n25633 n25644_not ; n25645
g25582 and n24955 n25014 ; n25646
g25583 nor n25015 n25646 ; n25647
g25584 and n71 n22380 ; n25648
g25585 and n9867 n22387 ; n25649
g25586 and n10434 n22384 ; n25650
g25587 nor n25649 n25650 ; n25651
g25588 and n25648_not n25651 ; n25652
g25589 and n9870_not n25652 ; n25653
g25590 and n22850_not n25652 ; n25654
g25591 nor n25653 n25654 ; n25655
g25592 and a[5] n25655_not ; n25656
g25593 and a[5]_not n25655 ; n25657
g25594 nor n25656 n25657 ; n25658
g25595 and n25647 n25658_not ; n25659
g25596 and n71 n22384 ; n25660
g25597 and n9867 n22390 ; n25661
g25598 and n10434 n22387 ; n25662
g25599 nor n25661 n25662 ; n25663
g25600 and n25660_not n25663 ; n25664
g25601 and n9870 n22806 ; n25665
g25602 and n25664 n25665_not ; n25666
g25603 and a[5] n25666_not ; n25667
g25604 nor n25666 n25667 ; n25668
g25605 and a[5] n25667_not ; n25669
g25606 nor n25668 n25669 ; n25670
g25607 and n25010 n25012_not ; n25671
g25608 nor n25013 n25671 ; n25672
g25609 and n25670_not n25672 ; n25673
g25610 nor n25670 n25673 ; n25674
g25611 and n25672 n25673_not ; n25675
g25612 nor n25674 n25675 ; n25676
g25613 nor n24997 n25009 ; n25677
g25614 nor n25008 n25009 ; n25678
g25615 nor n25677 n25678 ; n25679
g25616 and n71 n22387 ; n25680
g25617 and n9867 n22393 ; n25681
g25618 and n10434 n22390 ; n25682
g25619 nor n25681 n25682 ; n25683
g25620 and n25680_not n25683 ; n25684
g25621 and n9870_not n25684 ; n25685
g25622 and n22582_not n25684 ; n25686
g25623 nor n25685 n25686 ; n25687
g25624 and a[5] n25687_not ; n25688
g25625 and a[5]_not n25687 ; n25689
g25626 nor n25688 n25689 ; n25690
g25627 nor n25679 n25690 ; n25691
g25628 and n71 n22390 ; n25692
g25629 and n9867 n22396 ; n25693
g25630 and n10434 n22393 ; n25694
g25631 nor n25693 n25694 ; n25695
g25632 and n25692_not n25695 ; n25696
g25633 and n9870 n22649 ; n25697
g25634 and n25696 n25697_not ; n25698
g25635 and a[5] n25698_not ; n25699
g25636 nor n25698 n25699 ; n25700
g25637 and a[5] n25699_not ; n25701
g25638 nor n25700 n25701 ; n25702
g25639 and n24981_not n24992 ; n25703
g25640 nor n24993 n25703 ; n25704
g25641 and n25702_not n25704 ; n25705
g25642 nor n25702 n25705 ; n25706
g25643 and n25704 n25705_not ; n25707
g25644 nor n25706 n25707 ; n25708
g25645 and n24978 n24980_not ; n25709
g25646 nor n24981 n25709 ; n25710
g25647 and n71 n22393 ; n25711
g25648 and n9867 n22399 ; n25712
g25649 and n10434 n22396 ; n25713
g25650 nor n25712 n25713 ; n25714
g25651 and n25711_not n25714 ; n25715
g25652 and n9870_not n25715 ; n25716
g25653 and n22671_not n25715 ; n25717
g25654 nor n25716 n25717 ; n25718
g25655 and a[5] n25718_not ; n25719
g25656 and a[5]_not n25718 ; n25720
g25657 nor n25719 n25720 ; n25721
g25658 and n25710 n25721_not ; n25722
g25659 and n10434 n22406_not ; n25723
g25660 and n71 n22402 ; n25724
g25661 nor n25723 n25724 ; n25725
g25662 and n9870 n22609_not ; n25726
g25663 and n25725 n25726_not ; n25727
g25664 and a[5] n25727_not ; n25728
g25665 and a[5] n25728_not ; n25729
g25666 nor n25727 n25728 ; n25730
g25667 nor n25729 n25730 ; n25731
g25668 nor n70 n22406 ; n25732
g25669 and a[5] n25732_not ; n25733
g25670 and n25731_not n25733 ; n25734
g25671 and n71 n22399 ; n25735
g25672 and n9867 n22406_not ; n25736
g25673 and n10434 n22402 ; n25737
g25674 nor n25736 n25737 ; n25738
g25675 and n25735_not n25738 ; n25739
g25676 and n9870_not n25739 ; n25740
g25677 and n22625 n25739 ; n25741
g25678 nor n25740 n25741 ; n25742
g25679 and a[5] n25742_not ; n25743
g25680 and a[5]_not n25742 ; n25744
g25681 nor n25743 n25744 ; n25745
g25682 and n25734 n25745_not ; n25746
g25683 and n24979 n25746 ; n25747
g25684 and n25746 n25747_not ; n25748
g25685 and n24979 n25747_not ; n25749
g25686 nor n25748 n25749 ; n25750
g25687 and n71 n22396 ; n25751
g25688 and n9867 n22402 ; n25752
g25689 and n10434 n22399 ; n25753
g25690 nor n25752 n25753 ; n25754
g25691 and n25751_not n25754 ; n25755
g25692 and n9870 n22595 ; n25756
g25693 and n25755 n25756_not ; n25757
g25694 and a[5] n25757_not ; n25758
g25695 and a[5] n25758_not ; n25759
g25696 nor n25757 n25758 ; n25760
g25697 nor n25759 n25760 ; n25761
g25698 nor n25750 n25761 ; n25762
g25699 nor n25747 n25762 ; n25763
g25700 and n25710_not n25721 ; n25764
g25701 nor n25722 n25764 ; n25765
g25702 and n25763_not n25765 ; n25766
g25703 nor n25722 n25766 ; n25767
g25704 nor n25708 n25767 ; n25768
g25705 nor n25705 n25768 ; n25769
g25706 and n25679 n25690 ; n25770
g25707 nor n25691 n25770 ; n25771
g25708 and n25769_not n25771 ; n25772
g25709 nor n25691 n25772 ; n25773
g25710 nor n25676 n25773 ; n25774
g25711 nor n25673 n25774 ; n25775
g25712 and n25647 n25659_not ; n25776
g25713 nor n25658 n25659 ; n25777
g25714 nor n25776 n25777 ; n25778
g25715 nor n25775 n25778 ; n25779
g25716 nor n25659 n25779 ; n25780
g25717 and n25633 n25645_not ; n25781
g25718 nor n25644 n25645 ; n25782
g25719 nor n25781 n25782 ; n25783
g25720 nor n25780 n25783 ; n25784
g25721 nor n25645 n25784 ; n25785
g25722 and n25619_not n25630 ; n25786
g25723 nor n25631 n25786 ; n25787
g25724 and n25785_not n25787 ; n25788
g25725 nor n25631 n25788 ; n25789
g25726 nor n25617 n25789 ; n25790
g25727 nor n25614 n25790 ; n25791
g25728 nor n25599 n25791 ; n25792
g25729 nor n25596 n25792 ; n25793
g25730 nor n25581 n25793 ; n25794
g25731 nor n25578 n25794 ; n25795
g25732 and n25552 n25564_not ; n25796
g25733 nor n25563 n25564 ; n25797
g25734 nor n25796 n25797 ; n25798
g25735 nor n25795 n25798 ; n25799
g25736 nor n25564 n25799 ; n25800
g25737 and n25538 n25550_not ; n25801
g25738 nor n25549 n25550 ; n25802
g25739 nor n25801 n25802 ; n25803
g25740 nor n25800 n25803 ; n25804
g25741 nor n25550 n25804 ; n25805
g25742 and n25524_not n25535 ; n25806
g25743 nor n25536 n25806 ; n25807
g25744 and n25805_not n25807 ; n25808
g25745 nor n25536 n25808 ; n25809
g25746 nor n25522 n25809 ; n25810
g25747 nor n25519 n25810 ; n25811
g25748 nor n25504 n25811 ; n25812
g25749 nor n25501 n25812 ; n25813
g25750 nor n25486 n25813 ; n25814
g25751 nor n25483 n25814 ; n25815
g25752 and n25457 n25469_not ; n25816
g25753 nor n25468 n25469 ; n25817
g25754 nor n25816 n25817 ; n25818
g25755 nor n25815 n25818 ; n25819
g25756 nor n25469 n25819 ; n25820
g25757 and n25443 n25455_not ; n25821
g25758 nor n25454 n25455 ; n25822
g25759 nor n25821 n25822 ; n25823
g25760 nor n25820 n25823 ; n25824
g25761 nor n25455 n25824 ; n25825
g25762 and n25429_not n25440 ; n25826
g25763 nor n25441 n25826 ; n25827
g25764 and n25825_not n25827 ; n25828
g25765 nor n25441 n25828 ; n25829
g25766 nor n25427 n25829 ; n25830
g25767 nor n25424 n25830 ; n25831
g25768 nor n25409 n25831 ; n25832
g25769 nor n25406 n25832 ; n25833
g25770 nor n25391 n25833 ; n25834
g25771 nor n25388 n25834 ; n25835
g25772 and n25362 n25374_not ; n25836
g25773 nor n25373 n25374 ; n25837
g25774 nor n25836 n25837 ; n25838
g25775 nor n25835 n25838 ; n25839
g25776 nor n25374 n25839 ; n25840
g25777 and n25348_not n25359 ; n25841
g25778 nor n25360 n25841 ; n25842
g25779 and n25840_not n25842 ; n25843
g25780 nor n25360 n25843 ; n25844
g25781 nor n25346 n25844 ; n25845
g25782 nor n25343 n25845 ; n25846
g25783 nor n25328 n25846 ; n25847
g25784 nor n25325 n25847 ; n25848
g25785 nor n25307 n25848 ; n25849
g25786 nor n25304 n25849 ; n25850
g25787 and n25287 n25850 ; n25851
g25788 nor n25287 n25850 ; n25852
g25789 nor n25851 n25852 ; n25853
g25790 nor n22284 n22297 ; n25854
g25791 nor n22275 n22278 ; n25855
g25792 nor n22270 n22272 ; n25856
g25793 and n774 n6716 ; n25857
g25794 and n1824 n25857 ; n25858
g25795 and n3886 n25858 ; n25859
g25796 and n619_not n25859 ; n25860
g25797 and n452_not n25860 ; n25861
g25798 and n1203_not n25861 ; n25862
g25799 and n237_not n25862 ; n25863
g25800 and n792 n13063 ; n25864
g25801 and n3432 n25864 ; n25865
g25802 and n3764 n25865 ; n25866
g25803 and n3405 n25866 ; n25867
g25804 and n1601 n25867 ; n25868
g25805 and n25863 n25868 ; n25869
g25806 and n2276 n25869 ; n25870
g25807 and n1367 n25870 ; n25871
g25808 and n364_not n25871 ; n25872
g25809 and n495_not n25872 ; n25873
g25810 and n296_not n25873 ; n25874
g25811 and n25856_not n25874 ; n25875
g25812 and n25856 n25874_not ; n25876
g25813 nor n25875 n25876 ; n25877
g25814 and n3020 n13515 ; n25878
g25815 and n3028 n13521 ; n25879
g25816 and n3023 n13518 ; n25880
g25817 and n75 n13541 ; n25881
g25818 nor n25880 n25881 ; n25882
g25819 and n25879_not n25882 ; n25883
g25820 and n25878_not n25883 ; n25884
g25821 and n25877 n25884_not ; n25885
g25822 and n25877_not n25884 ; n25886
g25823 nor n25885 n25886 ; n25887
g25824 and n25855_not n25887 ; n25888
g25825 and n25855 n25887_not ; n25889
g25826 nor n25888 n25889 ; n25890
g25827 and n3457 n13633 ; n25891
g25828 and n3542 n13597 ; n25892
g25829 and n3606 n13630 ; n25893
g25830 nor n25892 n25893 ; n25894
g25831 and n25891_not n25894 ; n25895
g25832 and n3368_not n25895 ; n25896
g25833 and n13929_not n25895 ; n25897
g25834 nor n25896 n25897 ; n25898
g25835 and a[29] n25898_not ; n25899
g25836 and a[29]_not n25898 ; n25900
g25837 nor n25899 n25900 ; n25901
g25838 and n25890 n25901_not ; n25902
g25839 and n25890_not n25901 ; n25903
g25840 nor n25902 n25903 ; n25904
g25841 and n25854_not n25904 ; n25905
g25842 and n25854 n25904_not ; n25906
g25843 nor n25905 n25906 ; n25907
g25844 and n3884 n13438_not ; n25908
g25845 and n3967 n13627_not ; n25909
g25846 and n4046 n13941 ; n25910
g25847 nor n25909 n25910 ; n25911
g25848 and n25908_not n25911 ; n25912
g25849 and n4050 n14028 ; n25913
g25850 and n25912 n25913_not ; n25914
g25851 and a[26] n25914_not ; n25915
g25852 and a[26] n25915_not ; n25916
g25853 nor n25914 n25915 ; n25917
g25854 nor n25916 n25917 ; n25918
g25855 and n25907 n25918_not ; n25919
g25856 nor n25905 n25919 ; n25920
g25857 and n75 n13612_not ; n25921
g25858 and n3020 n13597 ; n25922
g25859 and n3023 n13521 ; n25923
g25860 and n3028 n13515 ; n25924
g25861 nor n25923 n25924 ; n25925
g25862 and n25922_not n25925 ; n25926
g25863 and n25921_not n25926 ; n25927
g25864 and n473 n1047 ; n25928
g25865 and n3978 n25928 ; n25929
g25866 and n3782 n25929 ; n25930
g25867 and n13063 n25930 ; n25931
g25868 and n1731 n25931 ; n25932
g25869 and n2170 n25932 ; n25933
g25870 and n3757 n25933 ; n25934
g25871 and n746_not n25934 ; n25935
g25872 and n296_not n25935 ; n25936
g25873 and n173_not n25936 ; n25937
g25874 and n601_not n25937 ; n25938
g25875 and n245_not n25938 ; n25939
g25876 and n142_not n25939 ; n25940
g25877 and n25874_not n25940 ; n25941
g25878 and n25874 n25940_not ; n25942
g25879 nor n25927 n25942 ; n25943
g25880 and n25941_not n25943 ; n25944
g25881 nor n25927 n25944 ; n25945
g25882 nor n25942 n25944 ; n25946
g25883 and n25941_not n25946 ; n25947
g25884 nor n25945 n25947 ; n25948
g25885 nor n25875 n25885 ; n25949
g25886 and n25948 n25949 ; n25950
g25887 nor n25948 n25949 ; n25951
g25888 nor n25950 n25951 ; n25952
g25889 nor n25888 n25902 ; n25953
g25890 and n25952_not n25953 ; n25954
g25891 and n25952 n25953_not ; n25955
g25892 nor n25954 n25955 ; n25956
g25893 nor n3884 n4046 ; n25957
g25894 nor n13438 n25957 ; n25958
g25895 and n3967 n13941 ; n25959
g25896 nor n25958 n25959 ; n25960
g25897 and n4050 n13951_not ; n25961
g25898 and n25960 n25961_not ; n25962
g25899 and a[26] n25962_not ; n25963
g25900 nor n25962 n25963 ; n25964
g25901 and a[26] n25963_not ; n25965
g25902 nor n25964 n25965 ; n25966
g25903 and n3457 n13627_not ; n25967
g25904 and n3542 n13630 ; n25968
g25905 and n3606 n13633 ; n25969
g25906 nor n25968 n25969 ; n25970
g25907 and n25967_not n25970 ; n25971
g25908 and n3368 n13654_not ; n25972
g25909 and n25971 n25972_not ; n25973
g25910 and a[29] n25973_not ; n25974
g25911 and a[29] n25974_not ; n25975
g25912 nor n25973 n25974 ; n25976
g25913 nor n25975 n25976 ; n25977
g25914 nor n25966 n25977 ; n25978
g25915 nor n25966 n25978 ; n25979
g25916 nor n25977 n25978 ; n25980
g25917 nor n25979 n25980 ; n25981
g25918 and n25956_not n25981 ; n25982
g25919 and n25956 n25981_not ; n25983
g25920 nor n25982 n25983 ; n25984
g25921 and n25920_not n25984 ; n25985
g25922 and n25907 n25919_not ; n25986
g25923 nor n25918 n25919 ; n25987
g25924 nor n25986 n25987 ; n25988
g25925 nor n22239 n22300 ; n25989
g25926 nor n22236 n25989 ; n25990
g25927 nor n25988 n25990 ; n25991
g25928 nor n25988 n25991 ; n25992
g25929 nor n25990 n25991 ; n25993
g25930 nor n25992 n25993 ; n25994
g25931 nor n22304 n22307 ; n25995
g25932 nor n25994 n25995 ; n25996
g25933 nor n25991 n25996 ; n25997
g25934 and n25920 n25984_not ; n25998
g25935 nor n25985 n25998 ; n25999
g25936 and n25997_not n25999 ; n26000
g25937 nor n25985 n26000 ; n26001
g25938 and n75 n13976 ; n26002
g25939 and n3020 n13630 ; n26003
g25940 and n3023 n13515 ; n26004
g25941 and n3028 n13597 ; n26005
g25942 nor n26004 n26005 ; n26006
g25943 and n26003_not n26006 ; n26007
g25944 and n26002_not n26007 ; n26008
g25945 and n3967_not n25957 ; n26009
g25946 and n4050_not n26009 ; n26010
g25947 nor n13438 n26010 ; n26011
g25948 and a[26] n26011_not ; n26012
g25949 and a[26]_not n26011 ; n26013
g25950 nor n26012 n26013 ; n26014
g25951 and n3873 n3972 ; n26015
g25952 and n296_not n26015 ; n26016
g25953 and n4017 n4040 ; n26017
g25954 and n2740 n26017 ; n26018
g25955 and n26016 n26018 ; n26019
g25956 and n328_not n26019 ; n26020
g25957 and n601_not n26020 ; n26021
g25958 and n25874 n26021 ; n26022
g25959 nor n25874 n26021 ; n26023
g25960 nor n26022 n26023 ; n26024
g25961 and n26014 n26024 ; n26025
g25962 nor n26014 n26024 ; n26026
g25963 nor n26025 n26026 ; n26027
g25964 and n25946_not n26027 ; n26028
g25965 and n25946 n26027_not ; n26029
g25966 nor n26028 n26029 ; n26030
g25967 and n26008_not n26030 ; n26031
g25968 and n26030 n26031_not ; n26032
g25969 nor n26008 n26031 ; n26033
g25970 nor n26032 n26033 ; n26034
g25971 and n3457 n13941 ; n26035
g25972 and n3542 n13633 ; n26036
g25973 and n3606 n13627_not ; n26037
g25974 nor n26036 n26037 ; n26038
g25975 and n26035_not n26038 ; n26039
g25976 and n3368 n14136 ; n26040
g25977 and n26039 n26040_not ; n26041
g25978 and a[29] n26041_not ; n26042
g25979 and a[29] n26042_not ; n26043
g25980 nor n26041 n26042 ; n26044
g25981 nor n26043 n26044 ; n26045
g25982 nor n26034 n26045 ; n26046
g25983 nor n26034 n26046 ; n26047
g25984 nor n26045 n26046 ; n26048
g25985 nor n26047 n26048 ; n26049
g25986 nor n25951 n25955 ; n26050
g25987 and n26049 n26050 ; n26051
g25988 nor n26049 n26050 ; n26052
g25989 nor n26051 n26052 ; n26053
g25990 nor n25978 n25983 ; n26054
g25991 and n26053 n26054_not ; n26055
g25992 and n26053_not n26054 ; n26056
g25993 nor n26055 n26056 ; n26057
g25994 and n26001 n26057_not ; n26058
g25995 and n26001_not n26057 ; n26059
g25996 nor n26058 n26059 ; n26060
g25997 and n11727 n26060 ; n26061
g25998 and n25994 n25995 ; n26062
g25999 nor n25996 n26062 ; n26063
g26000 and n11055 n26063 ; n26064
g26001 and n25997 n25999_not ; n26065
g26002 nor n26000 n26065 ; n26066
g26003 and n11715 n26066 ; n26067
g26004 nor n26064 n26067 ; n26068
g26005 and n26061_not n26068 ; n26069
g26006 and n11057_not n26069 ; n26070
g26007 and n26063 n26066 ; n26071
g26008 and n22309 n26063 ; n26072
g26009 nor n22309 n26063 ; n26073
g26010 nor n22527 n26073 ; n26074
g26011 and n26072_not n26074 ; n26075
g26012 nor n26072 n26075 ; n26076
g26013 nor n26063 n26066 ; n26077
g26014 nor n26076 n26077 ; n26078
g26015 and n26071_not n26078 ; n26079
g26016 nor n26071 n26079 ; n26080
g26017 and n26060 n26066 ; n26081
g26018 nor n26060 n26066 ; n26082
g26019 nor n26080 n26082 ; n26083
g26020 and n26081_not n26083 ; n26084
g26021 nor n26080 n26084 ; n26085
g26022 nor n26081 n26084 ; n26086
g26023 and n26082_not n26086 ; n26087
g26024 nor n26085 n26087 ; n26088
g26025 and n26069 n26088 ; n26089
g26026 nor n26070 n26089 ; n26090
g26027 and a[2] n26090_not ; n26091
g26028 and a[2]_not n26090 ; n26092
g26029 nor n26091 n26092 ; n26093
g26030 and n25853 n26093_not ; n26094
g26031 and n25840 n25842_not ; n26095
g26032 nor n25843 n26095 ; n26096
g26033 and n25825 n25827_not ; n26097
g26034 nor n25828 n26097 ; n26098
g26035 and n25805 n25807_not ; n26099
g26036 nor n25808 n26099 ; n26100
g26037 and n25785 n25787_not ; n26101
g26038 nor n25788 n26101 ; n26102
g26039 and n25763 n25765_not ; n26103
g26040 nor n25766 n26103 ; n26104
g26041 and n25734_not n25745 ; n26105
g26042 nor n25746 n26105 ; n26106
g26043 nor n11794 n22406 ; n26107
g26044 and n11796 n22625_not ; n26108
g26045 and n11727 n22399 ; n26109
g26046 and n11055 n22406_not ; n26110
g26047 and n11715 n22402 ; n26111
g26048 nor n26110 n26111 ; n26112
g26049 and n26109_not n26112 ; n26113
g26050 and a[2] n26113_not ; n26114
g26051 and n11796 n22609_not ; n26115
g26052 and n11805 n22406_not ; n26116
g26053 and n11807 n22402 ; n26117
g26054 and a[2] n26117_not ; n26118
g26055 and n26116_not n26118 ; n26119
g26056 and n26115_not n26119 ; n26120
g26057 and n26114_not n26120 ; n26121
g26058 and n26108_not n26121 ; n26122
g26059 and n26107_not n26122 ; n26123
g26060 and n25732 n26123 ; n26124
g26061 nor n25732 n26123 ; n26125
g26062 and n11727 n22396 ; n26126
g26063 and n11055 n22402 ; n26127
g26064 and n11715 n22399 ; n26128
g26065 nor n26127 n26128 ; n26129
g26066 and n26126_not n26129 ; n26130
g26067 and n11057 n22595 ; n26131
g26068 and n26130 n26131_not ; n26132
g26069 nor a[2] n26132 ; n26133
g26070 and a[2] n26132 ; n26134
g26071 nor n26133 n26134 ; n26135
g26072 nor n26125 n26135 ; n26136
g26073 nor n26124 n26136 ; n26137
g26074 and n11727 n22393 ; n26138
g26075 and n11055 n22399 ; n26139
g26076 and n11715 n22396 ; n26140
g26077 nor n26139 n26140 ; n26141
g26078 and n26138_not n26141 ; n26142
g26079 and n11057_not n26142 ; n26143
g26080 and n22671_not n26142 ; n26144
g26081 nor n26143 n26144 ; n26145
g26082 and a[2] n26145_not ; n26146
g26083 and a[2]_not n26145 ; n26147
g26084 nor n26146 n26147 ; n26148
g26085 and n26137 n26148 ; n26149
g26086 and n25731 n25733_not ; n26150
g26087 nor n25734 n26150 ; n26151
g26088 and n26149_not n26151 ; n26152
g26089 nor n26137 n26148 ; n26153
g26090 nor n26152 n26153 ; n26154
g26091 and n26106 n26154_not ; n26155
g26092 and n26106_not n26154 ; n26156
g26093 and n11727 n22390 ; n26157
g26094 and n11055 n22396 ; n26158
g26095 and n11715 n22393 ; n26159
g26096 nor n26158 n26159 ; n26160
g26097 and n26157_not n26160 ; n26161
g26098 and n11057 n22649 ; n26162
g26099 and n26161 n26162_not ; n26163
g26100 nor a[2] n26163 ; n26164
g26101 and a[2] n26163 ; n26165
g26102 nor n26164 n26165 ; n26166
g26103 nor n26156 n26166 ; n26167
g26104 nor n26155 n26167 ; n26168
g26105 and n11727 n22387 ; n26169
g26106 and n11055 n22393 ; n26170
g26107 and n11715 n22390 ; n26171
g26108 nor n26170 n26171 ; n26172
g26109 and n26169_not n26172 ; n26173
g26110 and n11057_not n26173 ; n26174
g26111 and n22582_not n26173 ; n26175
g26112 nor n26174 n26175 ; n26176
g26113 and a[2] n26176_not ; n26177
g26114 and a[2]_not n26176 ; n26178
g26115 nor n26177 n26178 ; n26179
g26116 nor n26168 n26179 ; n26180
g26117 and n26168 n26179 ; n26181
g26118 and n25750 n25761 ; n26182
g26119 nor n25762 n26182 ; n26183
g26120 and n26181_not n26183 ; n26184
g26121 nor n26180 n26184 ; n26185
g26122 and n26104 n26185_not ; n26186
g26123 and n26104_not n26185 ; n26187
g26124 and n11727 n22384 ; n26188
g26125 and n11055 n22390 ; n26189
g26126 and n11715 n22387 ; n26190
g26127 nor n26189 n26190 ; n26191
g26128 and n26188_not n26191 ; n26192
g26129 and n11057 n22806 ; n26193
g26130 and n26192 n26193_not ; n26194
g26131 nor a[2] n26194 ; n26195
g26132 and a[2] n26194 ; n26196
g26133 nor n26195 n26196 ; n26197
g26134 nor n26187 n26197 ; n26198
g26135 nor n26186 n26198 ; n26199
g26136 and n11727 n22380 ; n26200
g26137 and n11055 n22387 ; n26201
g26138 and n11715 n22384 ; n26202
g26139 nor n26201 n26202 ; n26203
g26140 and n26200_not n26203 ; n26204
g26141 and n11057_not n26204 ; n26205
g26142 and n22850_not n26204 ; n26206
g26143 nor n26205 n26206 ; n26207
g26144 and a[2] n26207_not ; n26208
g26145 and a[2]_not n26207 ; n26209
g26146 nor n26208 n26209 ; n26210
g26147 and n26199 n26210 ; n26211
g26148 and n25708 n25767 ; n26212
g26149 nor n25768 n26212 ; n26213
g26150 and n26211_not n26213 ; n26214
g26151 nor n26199 n26210 ; n26215
g26152 nor n26214 n26215 ; n26216
g26153 and n11727 n22377 ; n26217
g26154 and n11055 n22384 ; n26218
g26155 and n11715 n22380 ; n26219
g26156 nor n26218 n26219 ; n26220
g26157 and n26217_not n26220 ; n26221
g26158 and n11057_not n26221 ; n26222
g26159 and n22834 n26221 ; n26223
g26160 nor n26222 n26223 ; n26224
g26161 and a[2] n26224_not ; n26225
g26162 and a[2]_not n26224 ; n26226
g26163 nor n26225 n26226 ; n26227
g26164 and n26216 n26227 ; n26228
g26165 and n25769 n25771_not ; n26229
g26166 nor n25772 n26229 ; n26230
g26167 and n26228_not n26230 ; n26231
g26168 nor n26216 n26227 ; n26232
g26169 nor n26231 n26232 ; n26233
g26170 and n11727 n22374 ; n26234
g26171 and n11055 n22380 ; n26235
g26172 and n11715 n22377 ; n26236
g26173 nor n26235 n26236 ; n26237
g26174 and n26234_not n26237 ; n26238
g26175 and n11057_not n26238 ; n26239
g26176 and n22569_not n26238 ; n26240
g26177 nor n26239 n26240 ; n26241
g26178 and a[2] n26241_not ; n26242
g26179 and a[2]_not n26241 ; n26243
g26180 nor n26242 n26243 ; n26244
g26181 and n26233 n26244 ; n26245
g26182 and n25676 n25773 ; n26246
g26183 nor n25774 n26246 ; n26247
g26184 and n26245_not n26247 ; n26248
g26185 nor n26233 n26244 ; n26249
g26186 nor n26248 n26249 ; n26250
g26187 and n25775 n25777_not ; n26251
g26188 and n25776_not n26251 ; n26252
g26189 nor n25779 n26252 ; n26253
g26190 and n26250_not n26253 ; n26254
g26191 and n26250 n26253_not ; n26255
g26192 and n11727 n22371 ; n26256
g26193 and n11055 n22377 ; n26257
g26194 and n11715 n22374 ; n26258
g26195 nor n26257 n26258 ; n26259
g26196 and n26256_not n26259 ; n26260
g26197 and n11057 n23025 ; n26261
g26198 and n26260 n26261_not ; n26262
g26199 nor a[2] n26262 ; n26263
g26200 and a[2] n26262 ; n26264
g26201 nor n26263 n26264 ; n26265
g26202 nor n26255 n26265 ; n26266
g26203 nor n26254 n26266 ; n26267
g26204 and n25780 n25782_not ; n26268
g26205 and n25781_not n26268 ; n26269
g26206 nor n25784 n26269 ; n26270
g26207 and n26267_not n26270 ; n26271
g26208 and n26267 n26270_not ; n26272
g26209 and n11727 n22368 ; n26273
g26210 and n11055 n22374 ; n26274
g26211 and n11715 n22371 ; n26275
g26212 nor n26274 n26275 ; n26276
g26213 and n26273_not n26276 ; n26277
g26214 and n11057 n23006 ; n26278
g26215 and n26277 n26278_not ; n26279
g26216 nor a[2] n26279 ; n26280
g26217 and a[2] n26279 ; n26281
g26218 nor n26280 n26281 ; n26282
g26219 nor n26272 n26282 ; n26283
g26220 nor n26271 n26283 ; n26284
g26221 and n26102 n26284_not ; n26285
g26222 and n26102_not n26284 ; n26286
g26223 and n11727 n22365 ; n26287
g26224 and n11055 n22371 ; n26288
g26225 and n11715 n22368 ; n26289
g26226 nor n26288 n26289 ; n26290
g26227 and n26287_not n26290 ; n26291
g26228 and n11057 n22993_not ; n26292
g26229 and n26291 n26292_not ; n26293
g26230 nor a[2] n26293 ; n26294
g26231 and a[2] n26293 ; n26295
g26232 nor n26294 n26295 ; n26296
g26233 nor n26286 n26296 ; n26297
g26234 nor n26285 n26297 ; n26298
g26235 and n11727 n22362 ; n26299
g26236 and n11055 n22368 ; n26300
g26237 and n11715 n22365 ; n26301
g26238 nor n26300 n26301 ; n26302
g26239 and n26299_not n26302 ; n26303
g26240 and n11057_not n26303 ; n26304
g26241 and n23320 n26303 ; n26305
g26242 nor n26304 n26305 ; n26306
g26243 and a[2] n26306_not ; n26307
g26244 and a[2]_not n26306 ; n26308
g26245 nor n26307 n26308 ; n26309
g26246 and n26298 n26309 ; n26310
g26247 and n25617 n25789 ; n26311
g26248 nor n25790 n26311 ; n26312
g26249 and n26310_not n26312 ; n26313
g26250 nor n26298 n26309 ; n26314
g26251 nor n26313 n26314 ; n26315
g26252 and n11727 n22359 ; n26316
g26253 and n11055 n22365 ; n26317
g26254 and n11715 n22362 ; n26318
g26255 nor n26317 n26318 ; n26319
g26256 and n26316_not n26319 ; n26320
g26257 and n11057_not n26320 ; n26321
g26258 and n23368_not n26320 ; n26322
g26259 nor n26321 n26322 ; n26323
g26260 and a[2] n26323_not ; n26324
g26261 and a[2]_not n26323 ; n26325
g26262 nor n26324 n26325 ; n26326
g26263 and n26315 n26326 ; n26327
g26264 and n25599 n25791 ; n26328
g26265 nor n25792 n26328 ; n26329
g26266 and n26327_not n26329 ; n26330
g26267 nor n26315 n26326 ; n26331
g26268 nor n26330 n26331 ; n26332
g26269 and n11727 n22356 ; n26333
g26270 and n11055 n22362 ; n26334
g26271 and n11715 n22359 ; n26335
g26272 nor n26334 n26335 ; n26336
g26273 and n26333_not n26336 ; n26337
g26274 and n11057_not n26337 ; n26338
g26275 and n23345 n26337 ; n26339
g26276 nor n26338 n26339 ; n26340
g26277 and a[2] n26340_not ; n26341
g26278 and a[2]_not n26340 ; n26342
g26279 nor n26341 n26342 ; n26343
g26280 and n26332 n26343 ; n26344
g26281 and n25581 n25793 ; n26345
g26282 nor n25794 n26345 ; n26346
g26283 and n26344_not n26346 ; n26347
g26284 nor n26332 n26343 ; n26348
g26285 nor n26347 n26348 ; n26349
g26286 and n25795 n25797_not ; n26350
g26287 and n25796_not n26350 ; n26351
g26288 nor n25799 n26351 ; n26352
g26289 and n26349_not n26352 ; n26353
g26290 and n26349 n26352_not ; n26354
g26291 and n11727 n22353 ; n26355
g26292 and n11055 n22359 ; n26356
g26293 and n11715 n22356 ; n26357
g26294 nor n26356 n26357 ; n26358
g26295 and n26355_not n26358 ; n26359
g26296 and n11057 n22556_not ; n26360
g26297 and n26359 n26360_not ; n26361
g26298 nor a[2] n26361 ; n26362
g26299 and a[2] n26361 ; n26363
g26300 nor n26362 n26363 ; n26364
g26301 nor n26354 n26364 ; n26365
g26302 nor n26353 n26365 ; n26366
g26303 and n25800 n25802_not ; n26367
g26304 and n25801_not n26367 ; n26368
g26305 nor n25804 n26368 ; n26369
g26306 and n26366_not n26369 ; n26370
g26307 and n26366 n26369_not ; n26371
g26308 and n11727 n22350 ; n26372
g26309 and n11055 n22356 ; n26373
g26310 and n11715 n22353 ; n26374
g26311 nor n26373 n26374 ; n26375
g26312 and n26372_not n26375 ; n26376
g26313 and n11057 n23672 ; n26377
g26314 and n26376 n26377_not ; n26378
g26315 nor a[2] n26378 ; n26379
g26316 and a[2] n26378 ; n26380
g26317 nor n26379 n26380 ; n26381
g26318 nor n26371 n26381 ; n26382
g26319 nor n26370 n26382 ; n26383
g26320 and n26100 n26383_not ; n26384
g26321 and n26100_not n26383 ; n26385
g26322 and n11727 n22347 ; n26386
g26323 and n11055 n22353 ; n26387
g26324 and n11715 n22350 ; n26388
g26325 nor n26387 n26388 ; n26389
g26326 and n26386_not n26389 ; n26390
g26327 and n11057 n23659_not ; n26391
g26328 and n26390 n26391_not ; n26392
g26329 nor a[2] n26392 ; n26393
g26330 and a[2] n26392 ; n26394
g26331 nor n26393 n26394 ; n26395
g26332 nor n26385 n26395 ; n26396
g26333 nor n26384 n26396 ; n26397
g26334 and n11727 n22344 ; n26398
g26335 and n11055 n22350 ; n26399
g26336 and n11715 n22347 ; n26400
g26337 nor n26399 n26400 ; n26401
g26338 and n26398_not n26401 ; n26402
g26339 and n11057_not n26402 ; n26403
g26340 and n23642 n26402 ; n26404
g26341 nor n26403 n26404 ; n26405
g26342 and a[2] n26405_not ; n26406
g26343 and a[2]_not n26405 ; n26407
g26344 nor n26406 n26407 ; n26408
g26345 and n26397 n26408 ; n26409
g26346 and n25522 n25809 ; n26410
g26347 nor n25810 n26410 ; n26411
g26348 and n26409_not n26411 ; n26412
g26349 nor n26397 n26408 ; n26413
g26350 nor n26412 n26413 ; n26414
g26351 and n11727 n22341 ; n26415
g26352 and n11055 n22347 ; n26416
g26353 and n11715 n22344 ; n26417
g26354 nor n26416 n26417 ; n26418
g26355 and n26415_not n26418 ; n26419
g26356 and n11057_not n26419 ; n26420
g26357 and n24142_not n26419 ; n26421
g26358 nor n26420 n26421 ; n26422
g26359 and a[2] n26422_not ; n26423
g26360 and a[2]_not n26422 ; n26424
g26361 nor n26423 n26424 ; n26425
g26362 and n26414 n26425 ; n26426
g26363 and n25504 n25811 ; n26427
g26364 nor n25812 n26427 ; n26428
g26365 and n26426_not n26428 ; n26429
g26366 nor n26414 n26425 ; n26430
g26367 nor n26429 n26430 ; n26431
g26368 and n11727 n22338 ; n26432
g26369 and n11055 n22344 ; n26433
g26370 and n11715 n22341 ; n26434
g26371 nor n26433 n26434 ; n26435
g26372 and n26432_not n26435 ; n26436
g26373 and n11057_not n26436 ; n26437
g26374 and n24188 n26436 ; n26438
g26375 nor n26437 n26438 ; n26439
g26376 and a[2] n26439_not ; n26440
g26377 and a[2]_not n26439 ; n26441
g26378 nor n26440 n26441 ; n26442
g26379 and n26431 n26442 ; n26443
g26380 and n25486 n25813 ; n26444
g26381 nor n25814 n26444 ; n26445
g26382 and n26443_not n26445 ; n26446
g26383 nor n26431 n26442 ; n26447
g26384 nor n26446 n26447 ; n26448
g26385 and n25815 n25817_not ; n26449
g26386 and n25816_not n26449 ; n26450
g26387 nor n25819 n26450 ; n26451
g26388 and n26448_not n26451 ; n26452
g26389 and n26448 n26451_not ; n26453
g26390 and n11727 n22335 ; n26454
g26391 and n11055 n22341 ; n26455
g26392 and n11715 n22338 ; n26456
g26393 nor n26455 n26456 ; n26457
g26394 and n26454_not n26457 ; n26458
g26395 and n11057 n24167_not ; n26459
g26396 and n26458 n26459_not ; n26460
g26397 nor a[2] n26460 ; n26461
g26398 and a[2] n26460 ; n26462
g26399 nor n26461 n26462 ; n26463
g26400 nor n26453 n26463 ; n26464
g26401 nor n26452 n26464 ; n26465
g26402 and n25820 n25822_not ; n26466
g26403 and n25821_not n26466 ; n26467
g26404 nor n25824 n26467 ; n26468
g26405 and n26465_not n26468 ; n26469
g26406 and n26465 n26468_not ; n26470
g26407 and n11727 n22332 ; n26471
g26408 and n11055 n22338 ; n26472
g26409 and n11715 n22335 ; n26473
g26410 nor n26472 n26473 ; n26474
g26411 and n26471_not n26474 ; n26475
g26412 and n11057 n22542 ; n26476
g26413 and n26475 n26476_not ; n26477
g26414 nor a[2] n26477 ; n26478
g26415 and a[2] n26477 ; n26479
g26416 nor n26478 n26479 ; n26480
g26417 nor n26470 n26480 ; n26481
g26418 nor n26469 n26481 ; n26482
g26419 and n26098 n26482_not ; n26483
g26420 and n26098_not n26482 ; n26484
g26421 and n11727 n22329 ; n26485
g26422 and n11055 n22335 ; n26486
g26423 and n11715 n22332 ; n26487
g26424 nor n26486 n26487 ; n26488
g26425 and n26485_not n26488 ; n26489
g26426 and n11057 n24633_not ; n26490
g26427 and n26489 n26490_not ; n26491
g26428 nor a[2] n26491 ; n26492
g26429 and a[2] n26491 ; n26493
g26430 nor n26492 n26493 ; n26494
g26431 nor n26484 n26494 ; n26495
g26432 nor n26483 n26495 ; n26496
g26433 and n11727 n22326 ; n26497
g26434 and n11055 n22332 ; n26498
g26435 and n11715 n22329 ; n26499
g26436 nor n26498 n26499 ; n26500
g26437 and n26497_not n26500 ; n26501
g26438 and n11057_not n26501 ; n26502
g26439 and n24616 n26501 ; n26503
g26440 nor n26502 n26503 ; n26504
g26441 and a[2] n26504_not ; n26505
g26442 and a[2]_not n26504 ; n26506
g26443 nor n26505 n26506 ; n26507
g26444 and n26496 n26507 ; n26508
g26445 and n25427 n25829 ; n26509
g26446 nor n25830 n26509 ; n26510
g26447 and n26508_not n26510 ; n26511
g26448 nor n26496 n26507 ; n26512
g26449 nor n26511 n26512 ; n26513
g26450 and n11727 n22323 ; n26514
g26451 and n11055 n22329 ; n26515
g26452 and n11715 n22326 ; n26516
g26453 nor n26515 n26516 ; n26517
g26454 and n26514_not n26517 ; n26518
g26455 and n11057_not n26518 ; n26519
g26456 and n24599_not n26518 ; n26520
g26457 nor n26519 n26520 ; n26521
g26458 and a[2] n26521_not ; n26522
g26459 and a[2]_not n26521 ; n26523
g26460 nor n26522 n26523 ; n26524
g26461 and n26513 n26524 ; n26525
g26462 and n25409 n25831 ; n26526
g26463 nor n25832 n26526 ; n26527
g26464 and n26525_not n26527 ; n26528
g26465 nor n26513 n26524 ; n26529
g26466 nor n26528 n26529 ; n26530
g26467 and n11727 n22320 ; n26531
g26468 and n11055 n22326 ; n26532
g26469 and n11715 n22323 ; n26533
g26470 nor n26532 n26533 ; n26534
g26471 and n26531_not n26534 ; n26535
g26472 and n11057_not n26535 ; n26536
g26473 and n25270 n26535 ; n26537
g26474 nor n26536 n26537 ; n26538
g26475 and a[2] n26538_not ; n26539
g26476 and a[2]_not n26538 ; n26540
g26477 nor n26539 n26540 ; n26541
g26478 and n26530 n26541 ; n26542
g26479 and n25391 n25833 ; n26543
g26480 nor n25834 n26543 ; n26544
g26481 and n26542_not n26544 ; n26545
g26482 nor n26530 n26541 ; n26546
g26483 nor n26545 n26546 ; n26547
g26484 and n25835 n25837_not ; n26548
g26485 and n25836_not n26548 ; n26549
g26486 nor n25839 n26549 ; n26550
g26487 and n26547_not n26550 ; n26551
g26488 and n26547 n26550_not ; n26552
g26489 and n11727 n22312 ; n26553
g26490 and n11055 n22323 ; n26554
g26491 and n11715 n22320 ; n26555
g26492 nor n26554 n26555 ; n26556
g26493 and n26553_not n26556 ; n26557
g26494 and n11057 n25315_not ; n26558
g26495 and n26557 n26558_not ; n26559
g26496 nor a[2] n26559 ; n26560
g26497 and a[2] n26559 ; n26561
g26498 nor n26560 n26561 ; n26562
g26499 nor n26552 n26562 ; n26563
g26500 nor n26551 n26563 ; n26564
g26501 and n26096 n26564_not ; n26565
g26502 and n26096_not n26564 ; n26566
g26503 and n11727 n22315 ; n26567
g26504 and n11055 n22320 ; n26568
g26505 and n11715 n22312 ; n26569
g26506 nor n26568 n26569 ; n26570
g26507 and n26567_not n26570 ; n26571
g26508 and n11057 n25294 ; n26572
g26509 and n26571 n26572_not ; n26573
g26510 nor a[2] n26573 ; n26574
g26511 and a[2] n26573 ; n26575
g26512 nor n26574 n26575 ; n26576
g26513 nor n26566 n26576 ; n26577
g26514 nor n26565 n26577 ; n26578
g26515 and n11727 n22309 ; n26579
g26516 and n11055 n22312 ; n26580
g26517 and n11715 n22315 ; n26581
g26518 nor n26580 n26581 ; n26582
g26519 and n26579_not n26582 ; n26583
g26520 and n11057_not n26583 ; n26584
g26521 and n22529 n26583 ; n26585
g26522 nor n26584 n26585 ; n26586
g26523 and a[2] n26586_not ; n26587
g26524 and a[2]_not n26586 ; n26588
g26525 nor n26587 n26588 ; n26589
g26526 and n26578 n26589 ; n26590
g26527 and n25346 n25844 ; n26591
g26528 nor n25845 n26591 ; n26592
g26529 and n26590_not n26592 ; n26593
g26530 nor n26578 n26589 ; n26594
g26531 nor n26593 n26594 ; n26595
g26532 and n11727 n26063 ; n26596
g26533 and n11055 n22315 ; n26597
g26534 and n11715 n22309 ; n26598
g26535 nor n26597 n26598 ; n26599
g26536 and n26596_not n26599 ; n26600
g26537 and n11057_not n26600 ; n26601
g26538 nor n22527 n26075 ; n26602
g26539 and n26073_not n26076 ; n26603
g26540 nor n26602 n26603 ; n26604
g26541 and n26600 n26604 ; n26605
g26542 nor n26601 n26605 ; n26606
g26543 and a[2] n26606_not ; n26607
g26544 and a[2]_not n26606 ; n26608
g26545 nor n26607 n26608 ; n26609
g26546 and n26595 n26609 ; n26610
g26547 and n25328 n25846 ; n26611
g26548 nor n25847 n26611 ; n26612
g26549 and n26610_not n26612 ; n26613
g26550 nor n26595 n26609 ; n26614
g26551 nor n26613 n26614 ; n26615
g26552 and n11727 n26066 ; n26616
g26553 and n11055 n22309 ; n26617
g26554 and n11715 n26063 ; n26618
g26555 nor n26617 n26618 ; n26619
g26556 and n26616_not n26619 ; n26620
g26557 and n11057_not n26620 ; n26621
g26558 nor n26076 n26079 ; n26622
g26559 and n26077_not n26080 ; n26623
g26560 nor n26622 n26623 ; n26624
g26561 and n26620 n26624 ; n26625
g26562 nor n26621 n26625 ; n26626
g26563 and a[2] n26626_not ; n26627
g26564 and a[2]_not n26626 ; n26628
g26565 nor n26627 n26628 ; n26629
g26566 and n26615 n26629 ; n26630
g26567 and n25307 n25848 ; n26631
g26568 nor n25849 n26631 ; n26632
g26569 and n26630_not n26632 ; n26633
g26570 nor n26615 n26629 ; n26634
g26571 nor n26633 n26634 ; n26635
g26572 and n25853 n26094_not ; n26636
g26573 nor n26093 n26094 ; n26637
g26574 nor n26636 n26637 ; n26638
g26575 nor n26635 n26638 ; n26639
g26576 nor n26094 n26639 ; n26640
g26577 and n71 n26063 ; n26641
g26578 and n9867 n22315 ; n26642
g26579 and n10434 n22309 ; n26643
g26580 nor n26642 n26643 ; n26644
g26581 and n26641_not n26644 ; n26645
g26582 and n9870 n26604_not ; n26646
g26583 and n26645 n26646_not ; n26647
g26584 and a[5] n26647_not ; n26648
g26585 nor n26647 n26648 ; n26649
g26586 and a[5] n26648_not ; n26650
g26587 nor n26649 n26650 ; n26651
g26588 nor n25276 n25280 ; n26652
g26589 and n7983 n22326 ; n26653
g26590 and n7291 n22332 ; n26654
g26591 and n7632 n22329 ; n26655
g26592 nor n26654 n26655 ; n26656
g26593 and n26653_not n26656 ; n26657
g26594 and n7294 n24616_not ; n26658
g26595 and n26657 n26658_not ; n26659
g26596 and a[11] n26659_not ; n26660
g26597 nor n26659 n26660 ; n26661
g26598 and a[11] n26660_not ; n26662
g26599 nor n26661 n26662 ; n26663
g26600 nor n25246 n25250 ; n26664
g26601 and n6233 n22344 ; n26665
g26602 and n5663 n22350 ; n26666
g26603 and n5939 n22347 ; n26667
g26604 nor n26666 n26667 ; n26668
g26605 and n26665_not n26668 ; n26669
g26606 and n5666 n23642_not ; n26670
g26607 and n26669 n26670_not ; n26671
g26608 and a[17] n26671_not ; n26672
g26609 nor n26671 n26672 ; n26673
g26610 and a[17] n26672_not ; n26674
g26611 nor n26673 n26674 ; n26675
g26612 nor n25219 n25223 ; n26676
g26613 and n4694 n22362 ; n26677
g26614 and n4533 n22368 ; n26678
g26615 and n4604 n22365 ; n26679
g26616 nor n26678 n26679 ; n26680
g26617 and n26677_not n26680 ; n26681
g26618 and n4536 n23320_not ; n26682
g26619 and n26681 n26682_not ; n26683
g26620 and a[23] n26683_not ; n26684
g26621 nor n26683 n26684 ; n26685
g26622 and a[23] n26684_not ; n26686
g26623 nor n26685 n26686 ; n26687
g26624 nor n25192 n25196 ; n26688
g26625 and n3457 n22380 ; n26689
g26626 and n3542 n22387 ; n26690
g26627 and n3606 n22384 ; n26691
g26628 nor n26690 n26691 ; n26692
g26629 and n26689_not n26692 ; n26693
g26630 and n3368 n22850 ; n26694
g26631 and n26693 n26694_not ; n26695
g26632 and a[29] n26695_not ; n26696
g26633 nor n26695 n26696 ; n26697
g26634 and a[29] n26696_not ; n26698
g26635 nor n26697 n26698 ; n26699
g26636 nor n25165 n25169 ; n26700
g26637 and n12397 n13789 ; n26701
g26638 and n4771 n26701 ; n26702
g26639 and n1887 n26702 ; n26703
g26640 and n790 n26703 ; n26704
g26641 and n13677 n26704 ; n26705
g26642 and n4311 n26705 ; n26706
g26643 and n3155 n26706 ; n26707
g26644 and n244 n26707 ; n26708
g26645 and n933 n26708 ; n26709
g26646 and n1237 n26709 ; n26710
g26647 and n116 n26710 ; n26711
g26648 and n1101_not n26711 ; n26712
g26649 and n422_not n26712 ; n26713
g26650 and n493_not n26713 ; n26714
g26651 and n428_not n26714 ; n26715
g26652 and n3020 n22390 ; n26716
g26653 and n3028 n22393 ; n26717
g26654 and n3023 n22396 ; n26718
g26655 and n75 n22649 ; n26719
g26656 nor n26718 n26719 ; n26720
g26657 and n26717_not n26720 ; n26721
g26658 and n26716_not n26721 ; n26722
g26659 nor n26715 n26722 ; n26723
g26660 nor n26715 n26723 ; n26724
g26661 nor n26722 n26723 ; n26725
g26662 nor n26724 n26725 ; n26726
g26663 nor n26700 n26726 ; n26727
g26664 nor n26700 n26727 ; n26728
g26665 nor n26726 n26727 ; n26729
g26666 nor n26728 n26729 ; n26730
g26667 nor n26699 n26730 ; n26731
g26668 nor n26699 n26731 ; n26732
g26669 nor n26730 n26731 ; n26733
g26670 nor n26732 n26733 ; n26734
g26671 nor n25173 n25179 ; n26735
g26672 and n26734 n26735 ; n26736
g26673 nor n26734 n26735 ; n26737
g26674 nor n26736 n26737 ; n26738
g26675 and n3884 n22371 ; n26739
g26676 and n3967 n22377 ; n26740
g26677 and n4046 n22374 ; n26741
g26678 nor n26740 n26741 ; n26742
g26679 and n26739_not n26742 ; n26743
g26680 and n4050_not n26743 ; n26744
g26681 and n23025_not n26743 ; n26745
g26682 nor n26744 n26745 ; n26746
g26683 and a[26] n26746_not ; n26747
g26684 and a[26]_not n26746 ; n26748
g26685 nor n26747 n26748 ; n26749
g26686 and n26738 n26749_not ; n26750
g26687 and n26738 n26750_not ; n26751
g26688 nor n26749 n26750 ; n26752
g26689 nor n26751 n26752 ; n26753
g26690 nor n26688 n26753 ; n26754
g26691 nor n26688 n26754 ; n26755
g26692 nor n26753 n26754 ; n26756
g26693 nor n26755 n26756 ; n26757
g26694 nor n26687 n26757 ; n26758
g26695 nor n26687 n26758 ; n26759
g26696 nor n26757 n26758 ; n26760
g26697 nor n26759 n26760 ; n26761
g26698 nor n25200 n25206 ; n26762
g26699 and n26761 n26762 ; n26763
g26700 nor n26761 n26762 ; n26764
g26701 nor n26763 n26764 ; n26765
g26702 and n5496 n22353 ; n26766
g26703 and n4935 n22359 ; n26767
g26704 and n5407 n22356 ; n26768
g26705 nor n26767 n26768 ; n26769
g26706 and n26766_not n26769 ; n26770
g26707 and n4938_not n26770 ; n26771
g26708 and n22556 n26770 ; n26772
g26709 nor n26771 n26772 ; n26773
g26710 and a[20] n26773_not ; n26774
g26711 and a[20]_not n26773 ; n26775
g26712 nor n26774 n26775 ; n26776
g26713 and n26765 n26776_not ; n26777
g26714 and n26765 n26777_not ; n26778
g26715 nor n26776 n26777 ; n26779
g26716 nor n26778 n26779 ; n26780
g26717 nor n26676 n26780 ; n26781
g26718 nor n26676 n26781 ; n26782
g26719 nor n26780 n26781 ; n26783
g26720 nor n26782 n26783 ; n26784
g26721 nor n26675 n26784 ; n26785
g26722 nor n26675 n26785 ; n26786
g26723 nor n26784 n26785 ; n26787
g26724 nor n26786 n26787 ; n26788
g26725 nor n25227 n25233 ; n26789
g26726 and n26788 n26789 ; n26790
g26727 nor n26788 n26789 ; n26791
g26728 nor n26790 n26791 ; n26792
g26729 and n7101 n22335 ; n26793
g26730 and n6402 n22341 ; n26794
g26731 and n6951 n22338 ; n26795
g26732 nor n26794 n26795 ; n26796
g26733 and n26793_not n26796 ; n26797
g26734 and n6397_not n26797 ; n26798
g26735 and n24167 n26797 ; n26799
g26736 nor n26798 n26799 ; n26800
g26737 and a[14] n26800_not ; n26801
g26738 and a[14]_not n26800 ; n26802
g26739 nor n26801 n26802 ; n26803
g26740 and n26792 n26803_not ; n26804
g26741 and n26792 n26804_not ; n26805
g26742 nor n26803 n26804 ; n26806
g26743 nor n26805 n26806 ; n26807
g26744 nor n26664 n26807 ; n26808
g26745 nor n26664 n26808 ; n26809
g26746 nor n26807 n26808 ; n26810
g26747 nor n26809 n26810 ; n26811
g26748 nor n26663 n26811 ; n26812
g26749 nor n26663 n26812 ; n26813
g26750 nor n26811 n26812 ; n26814
g26751 nor n26813 n26814 ; n26815
g26752 nor n25254 n25260 ; n26816
g26753 and n26815 n26816 ; n26817
g26754 nor n26815 n26816 ; n26818
g26755 nor n26817 n26818 ; n26819
g26756 and n9331 n22312 ; n26820
g26757 and n8418 n22323 ; n26821
g26758 and n8860 n22320 ; n26822
g26759 nor n26821 n26822 ; n26823
g26760 and n26820_not n26823 ; n26824
g26761 and n8421_not n26824 ; n26825
g26762 and n25315 n26824 ; n26826
g26763 nor n26825 n26826 ; n26827
g26764 and a[8] n26827_not ; n26828
g26765 and a[8]_not n26827 ; n26829
g26766 nor n26828 n26829 ; n26830
g26767 and n26819 n26830_not ; n26831
g26768 and n26819 n26831_not ; n26832
g26769 nor n26830 n26831 ; n26833
g26770 nor n26832 n26833 ; n26834
g26771 nor n26652 n26834 ; n26835
g26772 nor n26652 n26835 ; n26836
g26773 nor n26834 n26835 ; n26837
g26774 nor n26836 n26837 ; n26838
g26775 nor n26651 n26838 ; n26839
g26776 nor n26651 n26839 ; n26840
g26777 nor n26838 n26839 ; n26841
g26778 nor n26840 n26841 ; n26842
g26779 nor n25284 n25852 ; n26843
g26780 and n26842 n26843 ; n26844
g26781 nor n26842 n26843 ; n26845
g26782 nor n26844 n26845 ; n26846
g26783 nor n26055 n26059 ; n26847
g26784 nor n26046 n26052 ; n26848
g26785 and n75 n13929 ; n26849
g26786 and n3020 n13633 ; n26850
g26787 and n3023 n13597 ; n26851
g26788 and n3028 n13630 ; n26852
g26789 nor n26851 n26852 ; n26853
g26790 and n26850_not n26853 ; n26854
g26791 and n26849_not n26854 ; n26855
g26792 nor n26023 n26025 ; n26856
g26793 and n4030 n4511 ; n26857
g26794 and n26016 n26857 ; n26858
g26795 and n328_not n26858 ; n26859
g26796 and n26856_not n26859 ; n26860
g26797 and n26856 n26859_not ; n26861
g26798 nor n26860 n26861 ; n26862
g26799 and n26855_not n26862 ; n26863
g26800 nor n26855 n26863 ; n26864
g26801 and n26862 n26863_not ; n26865
g26802 nor n26864 n26865 ; n26866
g26803 nor n26028 n26031 ; n26867
g26804 and n26866 n26867 ; n26868
g26805 nor n26866 n26867 ; n26869
g26806 nor n26868 n26869 ; n26870
g26807 and n3457 n13438_not ; n26871
g26808 and n3542 n13627_not ; n26872
g26809 and n3606 n13941 ; n26873
g26810 nor n26872 n26873 ; n26874
g26811 and n26871_not n26874 ; n26875
g26812 and n3368_not n26875 ; n26876
g26813 and n14028_not n26875 ; n26877
g26814 nor n26876 n26877 ; n26878
g26815 and a[29] n26878_not ; n26879
g26816 and a[29]_not n26878 ; n26880
g26817 nor n26879 n26880 ; n26881
g26818 and n26870 n26881_not ; n26882
g26819 and n26870_not n26881 ; n26883
g26820 nor n26882 n26883 ; n26884
g26821 and n26848_not n26884 ; n26885
g26822 and n26848 n26884_not ; n26886
g26823 nor n26885 n26886 ; n26887
g26824 and n26847_not n26887 ; n26888
g26825 and n26847 n26887_not ; n26889
g26826 nor n26888 n26889 ; n26890
g26827 and n11727 n26890 ; n26891
g26828 and n11055 n26066 ; n26892
g26829 and n11715 n26060 ; n26893
g26830 nor n26892 n26893 ; n26894
g26831 and n26891_not n26894 ; n26895
g26832 and n11057_not n26895 ; n26896
g26833 and n26060 n26890 ; n26897
g26834 nor n26060 n26890 ; n26898
g26835 nor n26086 n26898 ; n26899
g26836 and n26897_not n26899 ; n26900
g26837 nor n26086 n26900 ; n26901
g26838 nor n26897 n26900 ; n26902
g26839 and n26898_not n26902 ; n26903
g26840 nor n26901 n26903 ; n26904
g26841 and n26895 n26904 ; n26905
g26842 nor n26896 n26905 ; n26906
g26843 and a[2] n26906_not ; n26907
g26844 and a[2]_not n26906 ; n26908
g26845 nor n26907 n26908 ; n26909
g26846 and n26846 n26909_not ; n26910
g26847 and n26846_not n26909 ; n26911
g26848 nor n26910 n26911 ; n26912
g26849 and n26640_not n26912 ; n26913
g26850 and n26640 n26912_not ; n26914
g26851 nor n26913 n26914 ; n26915
g26852 nor n26635 n26639 ; n26916
g26853 nor n26638 n26639 ; n26917
g26854 nor n26916 n26917 ; n26918
g26855 and n26915 n26918 ; n26919
g26856 nor n26915 n26918 ; n26920
g26857 or n26919 n26920 ; result[0]
g26858 and n26915 n26918_not ; n26922
g26859 nor n26910 n26913 ; n26923
g26860 and n71 n26066 ; n26924
g26861 and n9867 n22309 ; n26925
g26862 and n10434 n26063 ; n26926
g26863 nor n26925 n26926 ; n26927
g26864 and n26924_not n26927 ; n26928
g26865 and n9870 n26624_not ; n26929
g26866 and n26928 n26929_not ; n26930
g26867 and a[5] n26930_not ; n26931
g26868 nor n26930 n26931 ; n26932
g26869 and a[5] n26931_not ; n26933
g26870 nor n26932 n26933 ; n26934
g26871 nor n26831 n26835 ; n26935
g26872 and n7983 n22323 ; n26936
g26873 and n7291 n22329 ; n26937
g26874 and n7632 n22326 ; n26938
g26875 nor n26937 n26938 ; n26939
g26876 and n26936_not n26939 ; n26940
g26877 and n7294 n24599 ; n26941
g26878 and n26940 n26941_not ; n26942
g26879 and a[11] n26942_not ; n26943
g26880 nor n26942 n26943 ; n26944
g26881 and a[11] n26943_not ; n26945
g26882 nor n26944 n26945 ; n26946
g26883 nor n26804 n26808 ; n26947
g26884 and n6233 n22341 ; n26948
g26885 and n5663 n22347 ; n26949
g26886 and n5939 n22344 ; n26950
g26887 nor n26949 n26950 ; n26951
g26888 and n26948_not n26951 ; n26952
g26889 and n5666 n24142 ; n26953
g26890 and n26952 n26953_not ; n26954
g26891 and a[17] n26954_not ; n26955
g26892 nor n26954 n26955 ; n26956
g26893 and a[17] n26955_not ; n26957
g26894 nor n26956 n26957 ; n26958
g26895 nor n26777 n26781 ; n26959
g26896 and n4694 n22359 ; n26960
g26897 and n4533 n22365 ; n26961
g26898 and n4604 n22362 ; n26962
g26899 nor n26961 n26962 ; n26963
g26900 and n26960_not n26963 ; n26964
g26901 and n4536 n23368 ; n26965
g26902 and n26964 n26965_not ; n26966
g26903 and a[23] n26966_not ; n26967
g26904 nor n26966 n26967 ; n26968
g26905 and a[23] n26967_not ; n26969
g26906 nor n26968 n26969 ; n26970
g26907 nor n26750 n26754 ; n26971
g26908 nor n26731 n26737 ; n26972
g26909 nor n26723 n26727 ; n26973
g26910 and n1603 n3514 ; n26974
g26911 and n2025 n26974 ; n26975
g26912 and n6628 n26975 ; n26976
g26913 and n14544 n26976 ; n26977
g26914 and n6755 n26977 ; n26978
g26915 and n2979 n26978 ; n26979
g26916 and n3544 n26979 ; n26980
g26917 and n1575 n26980 ; n26981
g26918 and n2583 n26981 ; n26982
g26919 and n1237 n26982 ; n26983
g26920 and n2405 n26983 ; n26984
g26921 and n1522 n26984 ; n26985
g26922 and n1246_not n26985 ; n26986
g26923 and n330_not n26986 ; n26987
g26924 and n296_not n26987 ; n26988
g26925 and n372_not n26988 ; n26989
g26926 and n932_not n26989 ; n26990
g26927 and n771_not n26990 ; n26991
g26928 and n3020 n22387 ; n26992
g26929 and n3028 n22390 ; n26993
g26930 and n3023 n22393 ; n26994
g26931 and n75 n22582 ; n26995
g26932 nor n26994 n26995 ; n26996
g26933 and n26993_not n26996 ; n26997
g26934 and n26992_not n26997 ; n26998
g26935 nor n26991 n26998 ; n26999
g26936 nor n26991 n26999 ; n27000
g26937 nor n26998 n26999 ; n27001
g26938 nor n27000 n27001 ; n27002
g26939 nor n26973 n27002 ; n27003
g26940 nor n26973 n27003 ; n27004
g26941 nor n27002 n27003 ; n27005
g26942 nor n27004 n27005 ; n27006
g26943 and n3457 n22377 ; n27007
g26944 and n3542 n22384 ; n27008
g26945 and n3606 n22380 ; n27009
g26946 nor n27008 n27009 ; n27010
g26947 and n27007_not n27010 ; n27011
g26948 and n3368_not n27011 ; n27012
g26949 and n22834 n27011 ; n27013
g26950 nor n27012 n27013 ; n27014
g26951 and a[29] n27014_not ; n27015
g26952 and a[29]_not n27014 ; n27016
g26953 nor n27015 n27016 ; n27017
g26954 nor n27006 n27017 ; n27018
g26955 and n27006 n27017 ; n27019
g26956 nor n27018 n27019 ; n27020
g26957 and n26972_not n27020 ; n27021
g26958 and n26972 n27020_not ; n27022
g26959 nor n27021 n27022 ; n27023
g26960 and n3884 n22368 ; n27024
g26961 and n3967 n22374 ; n27025
g26962 and n4046 n22371 ; n27026
g26963 nor n27025 n27026 ; n27027
g26964 and n27024_not n27027 ; n27028
g26965 and n4050_not n27028 ; n27029
g26966 and n23006_not n27028 ; n27030
g26967 nor n27029 n27030 ; n27031
g26968 and a[26] n27031_not ; n27032
g26969 and a[26]_not n27031 ; n27033
g26970 nor n27032 n27033 ; n27034
g26971 and n27023 n27034_not ; n27035
g26972 and n27023 n27035_not ; n27036
g26973 nor n27034 n27035 ; n27037
g26974 nor n27036 n27037 ; n27038
g26975 nor n26971 n27038 ; n27039
g26976 nor n26971 n27039 ; n27040
g26977 nor n27038 n27039 ; n27041
g26978 nor n27040 n27041 ; n27042
g26979 nor n26970 n27042 ; n27043
g26980 nor n26970 n27043 ; n27044
g26981 nor n27042 n27043 ; n27045
g26982 nor n27044 n27045 ; n27046
g26983 nor n26758 n26764 ; n27047
g26984 and n27046 n27047 ; n27048
g26985 nor n27046 n27047 ; n27049
g26986 nor n27048 n27049 ; n27050
g26987 and n5496 n22350 ; n27051
g26988 and n4935 n22356 ; n27052
g26989 and n5407 n22353 ; n27053
g26990 nor n27052 n27053 ; n27054
g26991 and n27051_not n27054 ; n27055
g26992 and n4938_not n27055 ; n27056
g26993 and n23672_not n27055 ; n27057
g26994 nor n27056 n27057 ; n27058
g26995 and a[20] n27058_not ; n27059
g26996 and a[20]_not n27058 ; n27060
g26997 nor n27059 n27060 ; n27061
g26998 and n27050 n27061_not ; n27062
g26999 and n27050 n27062_not ; n27063
g27000 nor n27061 n27062 ; n27064
g27001 nor n27063 n27064 ; n27065
g27002 nor n26959 n27065 ; n27066
g27003 nor n26959 n27066 ; n27067
g27004 nor n27065 n27066 ; n27068
g27005 nor n27067 n27068 ; n27069
g27006 nor n26958 n27069 ; n27070
g27007 nor n26958 n27070 ; n27071
g27008 nor n27069 n27070 ; n27072
g27009 nor n27071 n27072 ; n27073
g27010 nor n26785 n26791 ; n27074
g27011 and n27073 n27074 ; n27075
g27012 nor n27073 n27074 ; n27076
g27013 nor n27075 n27076 ; n27077
g27014 and n7101 n22332 ; n27078
g27015 and n6402 n22338 ; n27079
g27016 and n6951 n22335 ; n27080
g27017 nor n27079 n27080 ; n27081
g27018 and n27078_not n27081 ; n27082
g27019 and n6397_not n27082 ; n27083
g27020 and n22542_not n27082 ; n27084
g27021 nor n27083 n27084 ; n27085
g27022 and a[14] n27085_not ; n27086
g27023 and a[14]_not n27085 ; n27087
g27024 nor n27086 n27087 ; n27088
g27025 and n27077 n27088_not ; n27089
g27026 and n27077 n27089_not ; n27090
g27027 nor n27088 n27089 ; n27091
g27028 nor n27090 n27091 ; n27092
g27029 nor n26947 n27092 ; n27093
g27030 nor n26947 n27093 ; n27094
g27031 nor n27092 n27093 ; n27095
g27032 nor n27094 n27095 ; n27096
g27033 nor n26946 n27096 ; n27097
g27034 nor n26946 n27097 ; n27098
g27035 nor n27096 n27097 ; n27099
g27036 nor n27098 n27099 ; n27100
g27037 nor n26812 n26818 ; n27101
g27038 and n27100 n27101 ; n27102
g27039 nor n27100 n27101 ; n27103
g27040 nor n27102 n27103 ; n27104
g27041 and n9331 n22315 ; n27105
g27042 and n8418 n22320 ; n27106
g27043 and n8860 n22312 ; n27107
g27044 nor n27106 n27107 ; n27108
g27045 and n27105_not n27108 ; n27109
g27046 and n8421_not n27109 ; n27110
g27047 and n25294_not n27109 ; n27111
g27048 nor n27110 n27111 ; n27112
g27049 and a[8] n27112_not ; n27113
g27050 and a[8]_not n27112 ; n27114
g27051 nor n27113 n27114 ; n27115
g27052 and n27104 n27115_not ; n27116
g27053 and n27104 n27116_not ; n27117
g27054 nor n27115 n27116 ; n27118
g27055 nor n27117 n27118 ; n27119
g27056 nor n26935 n27119 ; n27120
g27057 nor n26935 n27120 ; n27121
g27058 nor n27119 n27120 ; n27122
g27059 nor n27121 n27122 ; n27123
g27060 nor n26934 n27123 ; n27124
g27061 nor n26934 n27124 ; n27125
g27062 nor n27123 n27124 ; n27126
g27063 nor n27125 n27126 ; n27127
g27064 nor n26839 n26845 ; n27128
g27065 and n27127 n27128 ; n27129
g27066 nor n27127 n27128 ; n27130
g27067 nor n27129 n27130 ; n27131
g27068 nor n26885 n26888 ; n27132
g27069 nor n26869 n26882 ; n27133
g27070 nor n26860 n26863 ; n27134
g27071 and n3856 n4514 ; n27135
g27072 and n26859 n27135_not ; n27136
g27073 and n26859_not n27135 ; n27137
g27074 nor n27134 n27137 ; n27138
g27075 and n27136_not n27138 ; n27139
g27076 nor n27134 n27139 ; n27140
g27077 nor n27137 n27139 ; n27141
g27078 and n27136_not n27141 ; n27142
g27079 nor n27140 n27142 ; n27143
g27080 nor n3457 n3606 ; n27144
g27081 nor n13438 n27144 ; n27145
g27082 and n3542 n13941 ; n27146
g27083 nor n27145 n27146 ; n27147
g27084 and n3368 n13951_not ; n27148
g27085 and n27147 n27148_not ; n27149
g27086 and a[29] n27149_not ; n27150
g27087 nor n27149 n27150 ; n27151
g27088 and a[29] n27150_not ; n27152
g27089 nor n27151 n27152 ; n27153
g27090 and n75 n13654_not ; n27154
g27091 and n3020 n13627_not ; n27155
g27092 and n3023 n13630 ; n27156
g27093 and n3028 n13633 ; n27157
g27094 nor n27156 n27157 ; n27158
g27095 and n27155_not n27158 ; n27159
g27096 and n27154_not n27159 ; n27160
g27097 nor n27153 n27160 ; n27161
g27098 nor n27153 n27161 ; n27162
g27099 nor n27160 n27161 ; n27163
g27100 nor n27162 n27163 ; n27164
g27101 and n27143_not n27164 ; n27165
g27102 and n27143 n27164_not ; n27166
g27103 nor n27165 n27166 ; n27167
g27104 nor n27133 n27167 ; n27168
g27105 and n27133 n27167 ; n27169
g27106 nor n27168 n27169 ; n27170
g27107 and n27132_not n27170 ; n27171
g27108 and n27132 n27170_not ; n27172
g27109 nor n27171 n27172 ; n27173
g27110 and n11727 n27173 ; n27174
g27111 and n11055 n26060 ; n27175
g27112 and n11715 n26890 ; n27176
g27113 nor n27175 n27176 ; n27177
g27114 and n27174_not n27177 ; n27178
g27115 and n11057_not n27178 ; n27179
g27116 nor n26890 n27173 ; n27180
g27117 and n26890 n27173 ; n27181
g27118 nor n27180 n27181 ; n27182
g27119 and n26902_not n27182 ; n27183
g27120 and n26902 n27182_not ; n27184
g27121 nor n27183 n27184 ; n27185
g27122 and n27178 n27185_not ; n27186
g27123 nor n27179 n27186 ; n27187
g27124 and a[2] n27187_not ; n27188
g27125 and a[2]_not n27187 ; n27189
g27126 nor n27188 n27189 ; n27190
g27127 and n27131 n27190_not ; n27191
g27128 and n27131_not n27190 ; n27192
g27129 nor n27191 n27192 ; n27193
g27130 and n26923_not n27193 ; n27194
g27131 and n26923 n27193_not ; n27195
g27132 nor n27194 n27195 ; n27196
g27133 and n26922 n27196 ; n27197
g27134 nor n26922 n27196 ; n27198
g27135 nor n27197 n27198 ; result[1]
g27136 nor n27191 n27194 ; n27200
g27137 and n71 n26060 ; n27201
g27138 and n9867 n26063 ; n27202
g27139 and n10434 n26066 ; n27203
g27140 nor n27202 n27203 ; n27204
g27141 and n27201_not n27204 ; n27205
g27142 and n9870 n26088_not ; n27206
g27143 and n27205 n27206_not ; n27207
g27144 and a[5] n27207_not ; n27208
g27145 nor n27207 n27208 ; n27209
g27146 and a[5] n27208_not ; n27210
g27147 nor n27209 n27210 ; n27211
g27148 nor n27116 n27120 ; n27212
g27149 and n7983 n22320 ; n27213
g27150 and n7291 n22326 ; n27214
g27151 and n7632 n22323 ; n27215
g27152 nor n27214 n27215 ; n27216
g27153 and n27213_not n27216 ; n27217
g27154 and n7294 n25270_not ; n27218
g27155 and n27217 n27218_not ; n27219
g27156 and a[11] n27219_not ; n27220
g27157 nor n27219 n27220 ; n27221
g27158 and a[11] n27220_not ; n27222
g27159 nor n27221 n27222 ; n27223
g27160 nor n27089 n27093 ; n27224
g27161 and n6233 n22338 ; n27225
g27162 and n5663 n22344 ; n27226
g27163 and n5939 n22341 ; n27227
g27164 nor n27226 n27227 ; n27228
g27165 and n27225_not n27228 ; n27229
g27166 and n5666 n24188_not ; n27230
g27167 and n27229 n27230_not ; n27231
g27168 and a[17] n27231_not ; n27232
g27169 nor n27231 n27232 ; n27233
g27170 and a[17] n27232_not ; n27234
g27171 nor n27233 n27234 ; n27235
g27172 nor n27062 n27066 ; n27236
g27173 and n4694 n22356 ; n27237
g27174 and n4533 n22362 ; n27238
g27175 and n4604 n22359 ; n27239
g27176 nor n27238 n27239 ; n27240
g27177 and n27237_not n27240 ; n27241
g27178 and n4536 n23345_not ; n27242
g27179 and n27241 n27242_not ; n27243
g27180 and a[23] n27243_not ; n27244
g27181 nor n27243 n27244 ; n27245
g27182 and a[23] n27244_not ; n27246
g27183 nor n27245 n27246 ; n27247
g27184 nor n27035 n27039 ; n27248
g27185 nor n27018 n27021 ; n27249
g27186 nor n26999 n27003 ; n27250
g27187 and n13827 n14561 ; n27251
g27188 and n6717 n27251 ; n27252
g27189 and n2410 n27252 ; n27253
g27190 and n616 n27253 ; n27254
g27191 and n3180 n27254 ; n27255
g27192 and n3191 n27255 ; n27256
g27193 and n1600 n27256 ; n27257
g27194 and n1479 n27257 ; n27258
g27195 and n1844 n27258 ; n27259
g27196 and n515 n27259 ; n27260
g27197 and n1726 n27260 ; n27261
g27198 and n1269 n27261 ; n27262
g27199 and n107_not n27262 ; n27263
g27200 and n490_not n27263 ; n27264
g27201 and n286_not n27264 ; n27265
g27202 and n245_not n27265 ; n27266
g27203 and n470_not n27266 ; n27267
g27204 and n3020 n22384 ; n27268
g27205 and n3028 n22387 ; n27269
g27206 and n3023 n22390 ; n27270
g27207 and n75 n22806 ; n27271
g27208 nor n27270 n27271 ; n27272
g27209 and n27269_not n27272 ; n27273
g27210 and n27268_not n27273 ; n27274
g27211 nor n27267 n27274 ; n27275
g27212 nor n27267 n27275 ; n27276
g27213 nor n27274 n27275 ; n27277
g27214 nor n27276 n27277 ; n27278
g27215 nor n27250 n27278 ; n27279
g27216 nor n27250 n27279 ; n27280
g27217 nor n27278 n27279 ; n27281
g27218 nor n27280 n27281 ; n27282
g27219 and n3457 n22374 ; n27283
g27220 and n3542 n22380 ; n27284
g27221 and n3606 n22377 ; n27285
g27222 nor n27284 n27285 ; n27286
g27223 and n27283_not n27286 ; n27287
g27224 and n3368_not n27287 ; n27288
g27225 and n22569_not n27287 ; n27289
g27226 nor n27288 n27289 ; n27290
g27227 and a[29] n27290_not ; n27291
g27228 and a[29]_not n27290 ; n27292
g27229 nor n27291 n27292 ; n27293
g27230 nor n27282 n27293 ; n27294
g27231 and n27282 n27293 ; n27295
g27232 nor n27294 n27295 ; n27296
g27233 and n27249_not n27296 ; n27297
g27234 and n27249 n27296_not ; n27298
g27235 nor n27297 n27298 ; n27299
g27236 and n3884 n22365 ; n27300
g27237 and n3967 n22371 ; n27301
g27238 and n4046 n22368 ; n27302
g27239 nor n27301 n27302 ; n27303
g27240 and n27300_not n27303 ; n27304
g27241 and n4050_not n27304 ; n27305
g27242 and n22993 n27304 ; n27306
g27243 nor n27305 n27306 ; n27307
g27244 and a[26] n27307_not ; n27308
g27245 and a[26]_not n27307 ; n27309
g27246 nor n27308 n27309 ; n27310
g27247 and n27299 n27310_not ; n27311
g27248 and n27299 n27311_not ; n27312
g27249 nor n27310 n27311 ; n27313
g27250 nor n27312 n27313 ; n27314
g27251 nor n27248 n27314 ; n27315
g27252 nor n27248 n27315 ; n27316
g27253 nor n27314 n27315 ; n27317
g27254 nor n27316 n27317 ; n27318
g27255 nor n27247 n27318 ; n27319
g27256 nor n27247 n27319 ; n27320
g27257 nor n27318 n27319 ; n27321
g27258 nor n27320 n27321 ; n27322
g27259 nor n27043 n27049 ; n27323
g27260 and n27322 n27323 ; n27324
g27261 nor n27322 n27323 ; n27325
g27262 nor n27324 n27325 ; n27326
g27263 and n5496 n22347 ; n27327
g27264 and n4935 n22353 ; n27328
g27265 and n5407 n22350 ; n27329
g27266 nor n27328 n27329 ; n27330
g27267 and n27327_not n27330 ; n27331
g27268 and n4938_not n27331 ; n27332
g27269 and n23659 n27331 ; n27333
g27270 nor n27332 n27333 ; n27334
g27271 and a[20] n27334_not ; n27335
g27272 and a[20]_not n27334 ; n27336
g27273 nor n27335 n27336 ; n27337
g27274 and n27326 n27337_not ; n27338
g27275 and n27326 n27338_not ; n27339
g27276 nor n27337 n27338 ; n27340
g27277 nor n27339 n27340 ; n27341
g27278 nor n27236 n27341 ; n27342
g27279 nor n27236 n27342 ; n27343
g27280 nor n27341 n27342 ; n27344
g27281 nor n27343 n27344 ; n27345
g27282 nor n27235 n27345 ; n27346
g27283 nor n27235 n27346 ; n27347
g27284 nor n27345 n27346 ; n27348
g27285 nor n27347 n27348 ; n27349
g27286 nor n27070 n27076 ; n27350
g27287 and n27349 n27350 ; n27351
g27288 nor n27349 n27350 ; n27352
g27289 nor n27351 n27352 ; n27353
g27290 and n7101 n22329 ; n27354
g27291 and n6402 n22335 ; n27355
g27292 and n6951 n22332 ; n27356
g27293 nor n27355 n27356 ; n27357
g27294 and n27354_not n27357 ; n27358
g27295 and n6397_not n27358 ; n27359
g27296 and n24633 n27358 ; n27360
g27297 nor n27359 n27360 ; n27361
g27298 and a[14] n27361_not ; n27362
g27299 and a[14]_not n27361 ; n27363
g27300 nor n27362 n27363 ; n27364
g27301 and n27353 n27364_not ; n27365
g27302 and n27353 n27365_not ; n27366
g27303 nor n27364 n27365 ; n27367
g27304 nor n27366 n27367 ; n27368
g27305 nor n27224 n27368 ; n27369
g27306 nor n27224 n27369 ; n27370
g27307 nor n27368 n27369 ; n27371
g27308 nor n27370 n27371 ; n27372
g27309 nor n27223 n27372 ; n27373
g27310 nor n27223 n27373 ; n27374
g27311 nor n27372 n27373 ; n27375
g27312 nor n27374 n27375 ; n27376
g27313 nor n27097 n27103 ; n27377
g27314 and n27376 n27377 ; n27378
g27315 nor n27376 n27377 ; n27379
g27316 nor n27378 n27379 ; n27380
g27317 and n9331 n22309 ; n27381
g27318 and n8418 n22312 ; n27382
g27319 and n8860 n22315 ; n27383
g27320 nor n27382 n27383 ; n27384
g27321 and n27381_not n27384 ; n27385
g27322 and n8421_not n27385 ; n27386
g27323 and n22529 n27385 ; n27387
g27324 nor n27386 n27387 ; n27388
g27325 and a[8] n27388_not ; n27389
g27326 and a[8]_not n27388 ; n27390
g27327 nor n27389 n27390 ; n27391
g27328 and n27380 n27391_not ; n27392
g27329 and n27380 n27392_not ; n27393
g27330 nor n27391 n27392 ; n27394
g27331 nor n27393 n27394 ; n27395
g27332 nor n27212 n27395 ; n27396
g27333 nor n27212 n27396 ; n27397
g27334 nor n27395 n27396 ; n27398
g27335 nor n27397 n27398 ; n27399
g27336 nor n27211 n27399 ; n27400
g27337 nor n27211 n27400 ; n27401
g27338 nor n27399 n27400 ; n27402
g27339 nor n27401 n27402 ; n27403
g27340 nor n27124 n27130 ; n27404
g27341 and n27403 n27404 ; n27405
g27342 nor n27403 n27404 ; n27406
g27343 nor n27405 n27406 ; n27407
g27344 nor n27168 n27171 ; n27408
g27345 nor n27143 n27164 ; n27409
g27346 nor n27161 n27409 ; n27410
g27347 and n75 n14136 ; n27411
g27348 and n3020 n13941 ; n27412
g27349 and n3023 n13633 ; n27413
g27350 and n3028 n13627_not ; n27414
g27351 nor n27413 n27414 ; n27415
g27352 and n27412_not n27415 ; n27416
g27353 and n27411_not n27416 ; n27417
g27354 nor n3542 n3606 ; n27418
g27355 and n3367 n27418 ; n27419
g27356 nor n13438 n27419 ; n27420
g27357 and a[29] n27420_not ; n27421
g27358 and a[29]_not n27420 ; n27422
g27359 nor n27421 n27422 ; n27423
g27360 and n13056 n27135 ; n27424
g27361 nor n13056 n27135 ; n27425
g27362 nor n27424 n27425 ; n27426
g27363 and n27423 n27426 ; n27427
g27364 nor n27423 n27426 ; n27428
g27365 nor n27427 n27428 ; n27429
g27366 and n27417_not n27429 ; n27430
g27367 and n27429 n27430_not ; n27431
g27368 nor n27417 n27430 ; n27432
g27369 nor n27431 n27432 ; n27433
g27370 nor n27141 n27433 ; n27434
g27371 and n27141 n27433 ; n27435
g27372 nor n27434 n27435 ; n27436
g27373 and n27410_not n27436 ; n27437
g27374 and n27410 n27436_not ; n27438
g27375 nor n27437 n27438 ; n27439
g27376 and n27408_not n27439 ; n27440
g27377 and n27408 n27439_not ; n27441
g27378 nor n27440 n27441 ; n27442
g27379 and n11727 n27442 ; n27443
g27380 and n11055 n26890 ; n27444
g27381 and n11715 n27173 ; n27445
g27382 nor n27444 n27445 ; n27446
g27383 and n27443_not n27446 ; n27447
g27384 and n11057_not n27447 ; n27448
g27385 nor n27181 n27183 ; n27449
g27386 nor n27173 n27442 ; n27450
g27387 and n27173 n27442 ; n27451
g27388 nor n27450 n27451 ; n27452
g27389 and n27449_not n27452 ; n27453
g27390 and n27449 n27452_not ; n27454
g27391 nor n27453 n27454 ; n27455
g27392 and n27447 n27455_not ; n27456
g27393 nor n27448 n27456 ; n27457
g27394 and a[2] n27457_not ; n27458
g27395 and a[2]_not n27457 ; n27459
g27396 nor n27458 n27459 ; n27460
g27397 and n27407 n27460_not ; n27461
g27398 and n27407_not n27460 ; n27462
g27399 nor n27461 n27462 ; n27463
g27400 and n27200_not n27463 ; n27464
g27401 and n27200 n27463_not ; n27465
g27402 nor n27464 n27465 ; n27466
g27403 and n27197 n27466 ; n27467
g27404 nor n27197 n27466 ; n27468
g27405 nor n27467 n27468 ; result[2]
g27406 nor n27461 n27464 ; n27470
g27407 and n71 n26890 ; n27471
g27408 and n9867 n26066 ; n27472
g27409 and n10434 n26060 ; n27473
g27410 nor n27472 n27473 ; n27474
g27411 and n27471_not n27474 ; n27475
g27412 and n9870 n26904_not ; n27476
g27413 and n27475 n27476_not ; n27477
g27414 and a[5] n27477_not ; n27478
g27415 nor n27477 n27478 ; n27479
g27416 and a[5] n27478_not ; n27480
g27417 nor n27479 n27480 ; n27481
g27418 nor n27392 n27396 ; n27482
g27419 and n7983 n22312 ; n27483
g27420 and n7291 n22323 ; n27484
g27421 and n7632 n22320 ; n27485
g27422 nor n27484 n27485 ; n27486
g27423 and n27483_not n27486 ; n27487
g27424 and n7294 n25315_not ; n27488
g27425 and n27487 n27488_not ; n27489
g27426 and a[11] n27489_not ; n27490
g27427 nor n27489 n27490 ; n27491
g27428 and a[11] n27490_not ; n27492
g27429 nor n27491 n27492 ; n27493
g27430 nor n27365 n27369 ; n27494
g27431 and n6233 n22335 ; n27495
g27432 and n5663 n22341 ; n27496
g27433 and n5939 n22338 ; n27497
g27434 nor n27496 n27497 ; n27498
g27435 and n27495_not n27498 ; n27499
g27436 and n5666 n24167_not ; n27500
g27437 and n27499 n27500_not ; n27501
g27438 and a[17] n27501_not ; n27502
g27439 nor n27501 n27502 ; n27503
g27440 and a[17] n27502_not ; n27504
g27441 nor n27503 n27504 ; n27505
g27442 nor n27338 n27342 ; n27506
g27443 and n4694 n22353 ; n27507
g27444 and n4533 n22359 ; n27508
g27445 and n4604 n22356 ; n27509
g27446 nor n27508 n27509 ; n27510
g27447 and n27507_not n27510 ; n27511
g27448 and n4536 n22556_not ; n27512
g27449 and n27511 n27512_not ; n27513
g27450 and a[23] n27513_not ; n27514
g27451 nor n27513 n27514 ; n27515
g27452 and a[23] n27514_not ; n27516
g27453 nor n27515 n27516 ; n27517
g27454 nor n27311 n27315 ; n27518
g27455 nor n27294 n27297 ; n27519
g27456 nor n27275 n27279 ; n27520
g27457 and n156 n2466 ; n27521
g27458 and n2993 n27521 ; n27522
g27459 and n1721 n1737 ; n27523
g27460 and n27522 n27523 ; n27524
g27461 and n2410 n27524 ; n27525
g27462 and n4769 n27525 ; n27526
g27463 and n15743 n27526 ; n27527
g27464 and n6732 n27527 ; n27528
g27465 and n6769 n27528 ; n27529
g27466 and n2229 n27529 ; n27530
g27467 and n510 n27530 ; n27531
g27468 and n1826 n27531 ; n27532
g27469 and n1182 n27532 ; n27533
g27470 and n191_not n27533 ; n27534
g27471 and n340_not n27534 ; n27535
g27472 and n3020 n22380 ; n27536
g27473 and n3028 n22384 ; n27537
g27474 and n3023 n22387 ; n27538
g27475 and n75 n22850 ; n27539
g27476 nor n27538 n27539 ; n27540
g27477 and n27537_not n27540 ; n27541
g27478 and n27536_not n27541 ; n27542
g27479 nor n27535 n27542 ; n27543
g27480 nor n27535 n27543 ; n27544
g27481 nor n27542 n27543 ; n27545
g27482 nor n27544 n27545 ; n27546
g27483 nor n27520 n27546 ; n27547
g27484 nor n27520 n27547 ; n27548
g27485 nor n27546 n27547 ; n27549
g27486 nor n27548 n27549 ; n27550
g27487 and n3457 n22371 ; n27551
g27488 and n3542 n22377 ; n27552
g27489 and n3606 n22374 ; n27553
g27490 nor n27552 n27553 ; n27554
g27491 and n27551_not n27554 ; n27555
g27492 and n3368_not n27555 ; n27556
g27493 and n23025_not n27555 ; n27557
g27494 nor n27556 n27557 ; n27558
g27495 and a[29] n27558_not ; n27559
g27496 and a[29]_not n27558 ; n27560
g27497 nor n27559 n27560 ; n27561
g27498 nor n27550 n27561 ; n27562
g27499 and n27550 n27561 ; n27563
g27500 nor n27562 n27563 ; n27564
g27501 and n27519_not n27564 ; n27565
g27502 and n27519 n27564_not ; n27566
g27503 nor n27565 n27566 ; n27567
g27504 and n3884 n22362 ; n27568
g27505 and n3967 n22368 ; n27569
g27506 and n4046 n22365 ; n27570
g27507 nor n27569 n27570 ; n27571
g27508 and n27568_not n27571 ; n27572
g27509 and n4050_not n27572 ; n27573
g27510 and n23320 n27572 ; n27574
g27511 nor n27573 n27574 ; n27575
g27512 and a[26] n27575_not ; n27576
g27513 and a[26]_not n27575 ; n27577
g27514 nor n27576 n27577 ; n27578
g27515 and n27567 n27578_not ; n27579
g27516 and n27567 n27579_not ; n27580
g27517 nor n27578 n27579 ; n27581
g27518 nor n27580 n27581 ; n27582
g27519 nor n27518 n27582 ; n27583
g27520 nor n27518 n27583 ; n27584
g27521 nor n27582 n27583 ; n27585
g27522 nor n27584 n27585 ; n27586
g27523 nor n27517 n27586 ; n27587
g27524 nor n27517 n27587 ; n27588
g27525 nor n27586 n27587 ; n27589
g27526 nor n27588 n27589 ; n27590
g27527 nor n27319 n27325 ; n27591
g27528 and n27590 n27591 ; n27592
g27529 nor n27590 n27591 ; n27593
g27530 nor n27592 n27593 ; n27594
g27531 and n5496 n22344 ; n27595
g27532 and n4935 n22350 ; n27596
g27533 and n5407 n22347 ; n27597
g27534 nor n27596 n27597 ; n27598
g27535 and n27595_not n27598 ; n27599
g27536 and n4938_not n27599 ; n27600
g27537 and n23642 n27599 ; n27601
g27538 nor n27600 n27601 ; n27602
g27539 and a[20] n27602_not ; n27603
g27540 and a[20]_not n27602 ; n27604
g27541 nor n27603 n27604 ; n27605
g27542 and n27594 n27605_not ; n27606
g27543 and n27594 n27606_not ; n27607
g27544 nor n27605 n27606 ; n27608
g27545 nor n27607 n27608 ; n27609
g27546 nor n27506 n27609 ; n27610
g27547 nor n27506 n27610 ; n27611
g27548 nor n27609 n27610 ; n27612
g27549 nor n27611 n27612 ; n27613
g27550 nor n27505 n27613 ; n27614
g27551 nor n27505 n27614 ; n27615
g27552 nor n27613 n27614 ; n27616
g27553 nor n27615 n27616 ; n27617
g27554 nor n27346 n27352 ; n27618
g27555 and n27617 n27618 ; n27619
g27556 nor n27617 n27618 ; n27620
g27557 nor n27619 n27620 ; n27621
g27558 and n7101 n22326 ; n27622
g27559 and n6402 n22332 ; n27623
g27560 and n6951 n22329 ; n27624
g27561 nor n27623 n27624 ; n27625
g27562 and n27622_not n27625 ; n27626
g27563 and n6397_not n27626 ; n27627
g27564 and n24616 n27626 ; n27628
g27565 nor n27627 n27628 ; n27629
g27566 and a[14] n27629_not ; n27630
g27567 and a[14]_not n27629 ; n27631
g27568 nor n27630 n27631 ; n27632
g27569 and n27621 n27632_not ; n27633
g27570 and n27621 n27633_not ; n27634
g27571 nor n27632 n27633 ; n27635
g27572 nor n27634 n27635 ; n27636
g27573 nor n27494 n27636 ; n27637
g27574 nor n27494 n27637 ; n27638
g27575 nor n27636 n27637 ; n27639
g27576 nor n27638 n27639 ; n27640
g27577 nor n27493 n27640 ; n27641
g27578 nor n27493 n27641 ; n27642
g27579 nor n27640 n27641 ; n27643
g27580 nor n27642 n27643 ; n27644
g27581 nor n27373 n27379 ; n27645
g27582 and n27644 n27645 ; n27646
g27583 nor n27644 n27645 ; n27647
g27584 nor n27646 n27647 ; n27648
g27585 and n9331 n26063 ; n27649
g27586 and n8418 n22315 ; n27650
g27587 and n8860 n22309 ; n27651
g27588 nor n27650 n27651 ; n27652
g27589 and n27649_not n27652 ; n27653
g27590 and n8421_not n27653 ; n27654
g27591 and n26604 n27653 ; n27655
g27592 nor n27654 n27655 ; n27656
g27593 and a[8] n27656_not ; n27657
g27594 and a[8]_not n27656 ; n27658
g27595 nor n27657 n27658 ; n27659
g27596 and n27648 n27659_not ; n27660
g27597 and n27648 n27660_not ; n27661
g27598 nor n27659 n27660 ; n27662
g27599 nor n27661 n27662 ; n27663
g27600 nor n27482 n27663 ; n27664
g27601 nor n27482 n27664 ; n27665
g27602 nor n27663 n27664 ; n27666
g27603 nor n27665 n27666 ; n27667
g27604 nor n27481 n27667 ; n27668
g27605 nor n27481 n27668 ; n27669
g27606 nor n27667 n27668 ; n27670
g27607 nor n27669 n27670 ; n27671
g27608 nor n27400 n27406 ; n27672
g27609 and n27671 n27672 ; n27673
g27610 nor n27671 n27672 ; n27674
g27611 nor n27673 n27674 ; n27675
g27612 and n75 n14028 ; n27676
g27613 and n3020 n13438_not ; n27677
g27614 and n3023 n13627_not ; n27678
g27615 and n3028 n13941 ; n27679
g27616 nor n27678 n27679 ; n27680
g27617 and n27677_not n27680 ; n27681
g27618 and n27676_not n27681 ; n27682
g27619 nor n27425 n27427 ; n27683
g27620 and n3839 n27683_not ; n27684
g27621 and n3839_not n27683 ; n27685
g27622 nor n27684 n27685 ; n27686
g27623 and n27682_not n27686 ; n27687
g27624 nor n27682 n27687 ; n27688
g27625 and n27686 n27687_not ; n27689
g27626 nor n27688 n27689 ; n27690
g27627 nor n27430 n27434 ; n27691
g27628 and n27690 n27691 ; n27692
g27629 nor n27690 n27691 ; n27693
g27630 nor n27692 n27693 ; n27694
g27631 nor n27437 n27440 ; n27695
g27632 and n27694_not n27695 ; n27696
g27633 and n27694 n27695_not ; n27697
g27634 nor n27696 n27697 ; n27698
g27635 and n11727 n27698 ; n27699
g27636 and n11055 n27173 ; n27700
g27637 and n11715 n27442 ; n27701
g27638 nor n27700 n27701 ; n27702
g27639 and n27699_not n27702 ; n27703
g27640 and n11057_not n27703 ; n27704
g27641 nor n27451 n27453 ; n27705
g27642 and n27442 n27698 ; n27706
g27643 nor n27442 n27698 ; n27707
g27644 nor n27705 n27707 ; n27708
g27645 and n27706_not n27708 ; n27709
g27646 nor n27705 n27709 ; n27710
g27647 nor n27706 n27709 ; n27711
g27648 and n27707_not n27711 ; n27712
g27649 nor n27710 n27712 ; n27713
g27650 and n27703 n27713 ; n27714
g27651 nor n27704 n27714 ; n27715
g27652 and a[2] n27715_not ; n27716
g27653 and a[2]_not n27715 ; n27717
g27654 nor n27716 n27717 ; n27718
g27655 and n27675 n27718_not ; n27719
g27656 and n27675_not n27718 ; n27720
g27657 nor n27719 n27720 ; n27721
g27658 and n27470_not n27721 ; n27722
g27659 and n27470 n27721_not ; n27723
g27660 nor n27722 n27723 ; n27724
g27661 and n27467 n27724 ; n27725
g27662 nor n27467 n27724 ; n27726
g27663 nor n27725 n27726 ; result[3]
g27664 nor n27719 n27722 ; n27728
g27665 and n71 n27173 ; n27729
g27666 and n9867 n26060 ; n27730
g27667 and n10434 n26890 ; n27731
g27668 nor n27730 n27731 ; n27732
g27669 and n27729_not n27732 ; n27733
g27670 and n9870 n27185 ; n27734
g27671 and n27733 n27734_not ; n27735
g27672 and a[5] n27735_not ; n27736
g27673 nor n27735 n27736 ; n27737
g27674 and a[5] n27736_not ; n27738
g27675 nor n27737 n27738 ; n27739
g27676 nor n27660 n27664 ; n27740
g27677 and n7983 n22315 ; n27741
g27678 and n7291 n22320 ; n27742
g27679 and n7632 n22312 ; n27743
g27680 nor n27742 n27743 ; n27744
g27681 and n27741_not n27744 ; n27745
g27682 and n7294 n25294 ; n27746
g27683 and n27745 n27746_not ; n27747
g27684 and a[11] n27747_not ; n27748
g27685 nor n27747 n27748 ; n27749
g27686 and a[11] n27748_not ; n27750
g27687 nor n27749 n27750 ; n27751
g27688 nor n27633 n27637 ; n27752
g27689 and n6233 n22332 ; n27753
g27690 and n5663 n22338 ; n27754
g27691 and n5939 n22335 ; n27755
g27692 nor n27754 n27755 ; n27756
g27693 and n27753_not n27756 ; n27757
g27694 and n5666 n22542 ; n27758
g27695 and n27757 n27758_not ; n27759
g27696 and a[17] n27759_not ; n27760
g27697 nor n27759 n27760 ; n27761
g27698 and a[17] n27760_not ; n27762
g27699 nor n27761 n27762 ; n27763
g27700 nor n27606 n27610 ; n27764
g27701 and n4694 n22350 ; n27765
g27702 and n4533 n22356 ; n27766
g27703 and n4604 n22353 ; n27767
g27704 nor n27766 n27767 ; n27768
g27705 and n27765_not n27768 ; n27769
g27706 and n4536 n23672 ; n27770
g27707 and n27769 n27770_not ; n27771
g27708 and a[23] n27771_not ; n27772
g27709 nor n27771 n27772 ; n27773
g27710 and a[23] n27772_not ; n27774
g27711 nor n27773 n27774 ; n27775
g27712 nor n27579 n27583 ; n27776
g27713 nor n27562 n27565 ; n27777
g27714 nor n27543 n27547 ; n27778
g27715 and n1423 n2093 ; n27779
g27716 and n3544 n27779 ; n27780
g27717 and n1575 n27780 ; n27781
g27718 and n111_not n27781 ; n27782
g27719 and n400_not n27782 ; n27783
g27720 and n226_not n27783 ; n27784
g27721 and n206_not n27784 ; n27785
g27722 and n490_not n27785 ; n27786
g27723 and n165_not n27786 ; n27787
g27724 and n791_not n27787 ; n27788
g27725 and n886_not n27788 ; n27789
g27726 and n1140 n2092 ; n27790
g27727 and n1681 n27790 ; n27791
g27728 and n1240 n27791 ; n27792
g27729 and n526 n27792 ; n27793
g27730 and n3040 n27793 ; n27794
g27731 and n1709 n27794 ; n27795
g27732 and n3127 n27795 ; n27796
g27733 and n4388 n27796 ; n27797
g27734 and n2012 n27797 ; n27798
g27735 and n27789 n27798 ; n27799
g27736 and n120 n27799 ; n27800
g27737 and n978 n27800 ; n27801
g27738 and n570 n27801 ; n27802
g27739 and n330_not n27802 ; n27803
g27740 and n602_not n27803 ; n27804
g27741 and n107_not n27804 ; n27805
g27742 and n245_not n27805 ; n27806
g27743 and n429_not n27806 ; n27807
g27744 and n3020 n22377 ; n27808
g27745 and n3028 n22380 ; n27809
g27746 and n3023 n22384 ; n27810
g27747 and n75 n22834_not ; n27811
g27748 nor n27810 n27811 ; n27812
g27749 and n27809_not n27812 ; n27813
g27750 and n27808_not n27813 ; n27814
g27751 nor n27807 n27814 ; n27815
g27752 nor n27807 n27815 ; n27816
g27753 nor n27814 n27815 ; n27817
g27754 nor n27816 n27817 ; n27818
g27755 nor n27778 n27818 ; n27819
g27756 nor n27778 n27819 ; n27820
g27757 nor n27818 n27819 ; n27821
g27758 nor n27820 n27821 ; n27822
g27759 and n3457 n22368 ; n27823
g27760 and n3542 n22374 ; n27824
g27761 and n3606 n22371 ; n27825
g27762 nor n27824 n27825 ; n27826
g27763 and n27823_not n27826 ; n27827
g27764 and n3368_not n27827 ; n27828
g27765 and n23006_not n27827 ; n27829
g27766 nor n27828 n27829 ; n27830
g27767 and a[29] n27830_not ; n27831
g27768 and a[29]_not n27830 ; n27832
g27769 nor n27831 n27832 ; n27833
g27770 nor n27822 n27833 ; n27834
g27771 and n27822 n27833 ; n27835
g27772 nor n27834 n27835 ; n27836
g27773 and n27777_not n27836 ; n27837
g27774 and n27777 n27836_not ; n27838
g27775 nor n27837 n27838 ; n27839
g27776 and n3884 n22359 ; n27840
g27777 and n3967 n22365 ; n27841
g27778 and n4046 n22362 ; n27842
g27779 nor n27841 n27842 ; n27843
g27780 and n27840_not n27843 ; n27844
g27781 and n4050_not n27844 ; n27845
g27782 and n23368_not n27844 ; n27846
g27783 nor n27845 n27846 ; n27847
g27784 and a[26] n27847_not ; n27848
g27785 and a[26]_not n27847 ; n27849
g27786 nor n27848 n27849 ; n27850
g27787 and n27839 n27850_not ; n27851
g27788 and n27839 n27851_not ; n27852
g27789 nor n27850 n27851 ; n27853
g27790 nor n27852 n27853 ; n27854
g27791 nor n27776 n27854 ; n27855
g27792 nor n27776 n27855 ; n27856
g27793 nor n27854 n27855 ; n27857
g27794 nor n27856 n27857 ; n27858
g27795 nor n27775 n27858 ; n27859
g27796 nor n27775 n27859 ; n27860
g27797 nor n27858 n27859 ; n27861
g27798 nor n27860 n27861 ; n27862
g27799 nor n27587 n27593 ; n27863
g27800 and n27862 n27863 ; n27864
g27801 nor n27862 n27863 ; n27865
g27802 nor n27864 n27865 ; n27866
g27803 and n5496 n22341 ; n27867
g27804 and n4935 n22347 ; n27868
g27805 and n5407 n22344 ; n27869
g27806 nor n27868 n27869 ; n27870
g27807 and n27867_not n27870 ; n27871
g27808 and n4938_not n27871 ; n27872
g27809 and n24142_not n27871 ; n27873
g27810 nor n27872 n27873 ; n27874
g27811 and a[20] n27874_not ; n27875
g27812 and a[20]_not n27874 ; n27876
g27813 nor n27875 n27876 ; n27877
g27814 and n27866 n27877_not ; n27878
g27815 and n27866 n27878_not ; n27879
g27816 nor n27877 n27878 ; n27880
g27817 nor n27879 n27880 ; n27881
g27818 nor n27764 n27881 ; n27882
g27819 nor n27764 n27882 ; n27883
g27820 nor n27881 n27882 ; n27884
g27821 nor n27883 n27884 ; n27885
g27822 nor n27763 n27885 ; n27886
g27823 nor n27763 n27886 ; n27887
g27824 nor n27885 n27886 ; n27888
g27825 nor n27887 n27888 ; n27889
g27826 nor n27614 n27620 ; n27890
g27827 and n27889 n27890 ; n27891
g27828 nor n27889 n27890 ; n27892
g27829 nor n27891 n27892 ; n27893
g27830 and n7101 n22323 ; n27894
g27831 and n6402 n22329 ; n27895
g27832 and n6951 n22326 ; n27896
g27833 nor n27895 n27896 ; n27897
g27834 and n27894_not n27897 ; n27898
g27835 and n6397_not n27898 ; n27899
g27836 and n24599_not n27898 ; n27900
g27837 nor n27899 n27900 ; n27901
g27838 and a[14] n27901_not ; n27902
g27839 and a[14]_not n27901 ; n27903
g27840 nor n27902 n27903 ; n27904
g27841 and n27893 n27904_not ; n27905
g27842 and n27893 n27905_not ; n27906
g27843 nor n27904 n27905 ; n27907
g27844 nor n27906 n27907 ; n27908
g27845 nor n27752 n27908 ; n27909
g27846 nor n27752 n27909 ; n27910
g27847 nor n27908 n27909 ; n27911
g27848 nor n27910 n27911 ; n27912
g27849 nor n27751 n27912 ; n27913
g27850 nor n27751 n27913 ; n27914
g27851 nor n27912 n27913 ; n27915
g27852 nor n27914 n27915 ; n27916
g27853 nor n27641 n27647 ; n27917
g27854 and n27916 n27917 ; n27918
g27855 nor n27916 n27917 ; n27919
g27856 nor n27918 n27919 ; n27920
g27857 and n9331 n26066 ; n27921
g27858 and n8418 n22309 ; n27922
g27859 and n8860 n26063 ; n27923
g27860 nor n27922 n27923 ; n27924
g27861 and n27921_not n27924 ; n27925
g27862 and n8421_not n27925 ; n27926
g27863 and n26624 n27925 ; n27927
g27864 nor n27926 n27927 ; n27928
g27865 and a[8] n27928_not ; n27929
g27866 and a[8]_not n27928 ; n27930
g27867 nor n27929 n27930 ; n27931
g27868 and n27920 n27931_not ; n27932
g27869 and n27920 n27932_not ; n27933
g27870 nor n27931 n27932 ; n27934
g27871 nor n27933 n27934 ; n27935
g27872 nor n27740 n27935 ; n27936
g27873 nor n27740 n27936 ; n27937
g27874 nor n27935 n27936 ; n27938
g27875 nor n27937 n27938 ; n27939
g27876 nor n27739 n27939 ; n27940
g27877 nor n27739 n27940 ; n27941
g27878 nor n27939 n27940 ; n27942
g27879 nor n27941 n27942 ; n27943
g27880 nor n27668 n27674 ; n27944
g27881 and n27943 n27944 ; n27945
g27882 nor n27943 n27944 ; n27946
g27883 nor n27945 n27946 ; n27947
g27884 and n75 n13951_not ; n27948
g27885 nor n3020 n3028 ; n27949
g27886 nor n13438 n27949 ; n27950
g27887 and n3023 n13941 ; n27951
g27888 nor n27950 n27951 ; n27952
g27889 and n27948_not n27952 ; n27953
g27890 and n3839 n27953 ; n27954
g27891 nor n3839 n27953 ; n27955
g27892 nor n27954 n27955 ; n27956
g27893 nor n27684 n27687 ; n27957
g27894 and n27956 n27957 ; n27958
g27895 nor n27956 n27957 ; n27959
g27896 nor n27958 n27959 ; n27960
g27897 nor n27693 n27697 ; n27961
g27898 and n27960_not n27961 ; n27962
g27899 and n27960 n27961_not ; n27963
g27900 nor n27962 n27963 ; n27964
g27901 and n11727 n27964 ; n27965
g27902 and n11055 n27442 ; n27966
g27903 and n11715 n27698 ; n27967
g27904 nor n27966 n27967 ; n27968
g27905 and n27965_not n27968 ; n27969
g27906 and n11057_not n27969 ; n27970
g27907 nor n27698 n27964 ; n27971
g27908 and n27698 n27964 ; n27972
g27909 nor n27971 n27972 ; n27973
g27910 and n27711_not n27973 ; n27974
g27911 and n27711 n27973_not ; n27975
g27912 nor n27974 n27975 ; n27976
g27913 and n27969 n27976_not ; n27977
g27914 nor n27970 n27977 ; n27978
g27915 and a[2] n27978_not ; n27979
g27916 and a[2]_not n27978 ; n27980
g27917 nor n27979 n27980 ; n27981
g27918 and n27947 n27981_not ; n27982
g27919 and n27947_not n27981 ; n27983
g27920 nor n27982 n27983 ; n27984
g27921 and n27728_not n27984 ; n27985
g27922 and n27728 n27984_not ; n27986
g27923 nor n27985 n27986 ; n27987
g27924 and n27725 n27987 ; n27988
g27925 nor n27725 n27987 ; n27989
g27926 nor n27988 n27989 ; result[4]
g27927 nor n27982 n27985 ; n27991
g27928 and n71 n27442 ; n27992
g27929 and n9867 n26890 ; n27993
g27930 and n10434 n27173 ; n27994
g27931 nor n27993 n27994 ; n27995
g27932 and n27992_not n27995 ; n27996
g27933 and n9870 n27455 ; n27997
g27934 and n27996 n27997_not ; n27998
g27935 and a[5] n27998_not ; n27999
g27936 nor n27998 n27999 ; n28000
g27937 and a[5] n27999_not ; n28001
g27938 nor n28000 n28001 ; n28002
g27939 nor n27932 n27936 ; n28003
g27940 and n7983 n22309 ; n28004
g27941 and n7291 n22312 ; n28005
g27942 and n7632 n22315 ; n28006
g27943 nor n28005 n28006 ; n28007
g27944 and n28004_not n28007 ; n28008
g27945 and n7294 n22529_not ; n28009
g27946 and n28008 n28009_not ; n28010
g27947 and a[11] n28010_not ; n28011
g27948 nor n28010 n28011 ; n28012
g27949 and a[11] n28011_not ; n28013
g27950 nor n28012 n28013 ; n28014
g27951 nor n27905 n27909 ; n28015
g27952 and n6233 n22329 ; n28016
g27953 and n5663 n22335 ; n28017
g27954 and n5939 n22332 ; n28018
g27955 nor n28017 n28018 ; n28019
g27956 and n28016_not n28019 ; n28020
g27957 and n5666 n24633_not ; n28021
g27958 and n28020 n28021_not ; n28022
g27959 and a[17] n28022_not ; n28023
g27960 nor n28022 n28023 ; n28024
g27961 and a[17] n28023_not ; n28025
g27962 nor n28024 n28025 ; n28026
g27963 nor n27878 n27882 ; n28027
g27964 and n4694 n22347 ; n28028
g27965 and n4533 n22353 ; n28029
g27966 and n4604 n22350 ; n28030
g27967 nor n28029 n28030 ; n28031
g27968 and n28028_not n28031 ; n28032
g27969 and n4536 n23659_not ; n28033
g27970 and n28032 n28033_not ; n28034
g27971 and a[23] n28034_not ; n28035
g27972 nor n28034 n28035 ; n28036
g27973 and a[23] n28035_not ; n28037
g27974 nor n28036 n28037 ; n28038
g27975 nor n27851 n27855 ; n28039
g27976 nor n27834 n27837 ; n28040
g27977 nor n27815 n27819 ; n28041
g27978 and n207 n3587 ; n28042
g27979 and n690 n28042 ; n28043
g27980 and n12409 n28043 ; n28044
g27981 and n15970 n28044 ; n28045
g27982 and n3644 n28045 ; n28046
g27983 and n5286 n28046 ; n28047
g27984 and n1046 n28047 ; n28048
g27985 and n469_not n28048 ; n28049
g27986 and n111_not n28049 ; n28050
g27987 and n242_not n28050 ; n28051
g27988 and n171_not n28051 ; n28052
g27989 and n601_not n28052 ; n28053
g27990 and n375_not n28053 ; n28054
g27991 and n493_not n28054 ; n28055
g27992 and n161_not n28055 ; n28056
g27993 and n251_not n28056 ; n28057
g27994 and n158_not n28057 ; n28058
g27995 and n222_not n28058 ; n28059
g27996 and n3020 n22374 ; n28060
g27997 and n3028 n22377 ; n28061
g27998 and n3023 n22380 ; n28062
g27999 and n75 n22569 ; n28063
g28000 nor n28062 n28063 ; n28064
g28001 and n28061_not n28064 ; n28065
g28002 and n28060_not n28065 ; n28066
g28003 nor n28059 n28066 ; n28067
g28004 nor n28059 n28067 ; n28068
g28005 nor n28066 n28067 ; n28069
g28006 nor n28068 n28069 ; n28070
g28007 nor n28041 n28070 ; n28071
g28008 nor n28041 n28071 ; n28072
g28009 nor n28070 n28071 ; n28073
g28010 nor n28072 n28073 ; n28074
g28011 and n3457 n22365 ; n28075
g28012 and n3542 n22371 ; n28076
g28013 and n3606 n22368 ; n28077
g28014 nor n28076 n28077 ; n28078
g28015 and n28075_not n28078 ; n28079
g28016 and n3368_not n28079 ; n28080
g28017 and n22993 n28079 ; n28081
g28018 nor n28080 n28081 ; n28082
g28019 and a[29] n28082_not ; n28083
g28020 and a[29]_not n28082 ; n28084
g28021 nor n28083 n28084 ; n28085
g28022 nor n28074 n28085 ; n28086
g28023 and n28074 n28085 ; n28087
g28024 nor n28086 n28087 ; n28088
g28025 and n28040_not n28088 ; n28089
g28026 and n28040 n28088_not ; n28090
g28027 nor n28089 n28090 ; n28091
g28028 and n3884 n22356 ; n28092
g28029 and n3967 n22362 ; n28093
g28030 and n4046 n22359 ; n28094
g28031 nor n28093 n28094 ; n28095
g28032 and n28092_not n28095 ; n28096
g28033 and n4050_not n28096 ; n28097
g28034 and n23345 n28096 ; n28098
g28035 nor n28097 n28098 ; n28099
g28036 and a[26] n28099_not ; n28100
g28037 and a[26]_not n28099 ; n28101
g28038 nor n28100 n28101 ; n28102
g28039 and n28091 n28102_not ; n28103
g28040 and n28091 n28103_not ; n28104
g28041 nor n28102 n28103 ; n28105
g28042 nor n28104 n28105 ; n28106
g28043 nor n28039 n28106 ; n28107
g28044 nor n28039 n28107 ; n28108
g28045 nor n28106 n28107 ; n28109
g28046 nor n28108 n28109 ; n28110
g28047 nor n28038 n28110 ; n28111
g28048 nor n28038 n28111 ; n28112
g28049 nor n28110 n28111 ; n28113
g28050 nor n28112 n28113 ; n28114
g28051 nor n27859 n27865 ; n28115
g28052 and n28114 n28115 ; n28116
g28053 nor n28114 n28115 ; n28117
g28054 nor n28116 n28117 ; n28118
g28055 and n5496 n22338 ; n28119
g28056 and n4935 n22344 ; n28120
g28057 and n5407 n22341 ; n28121
g28058 nor n28120 n28121 ; n28122
g28059 and n28119_not n28122 ; n28123
g28060 and n4938_not n28123 ; n28124
g28061 and n24188 n28123 ; n28125
g28062 nor n28124 n28125 ; n28126
g28063 and a[20] n28126_not ; n28127
g28064 and a[20]_not n28126 ; n28128
g28065 nor n28127 n28128 ; n28129
g28066 and n28118 n28129_not ; n28130
g28067 and n28118 n28130_not ; n28131
g28068 nor n28129 n28130 ; n28132
g28069 nor n28131 n28132 ; n28133
g28070 nor n28027 n28133 ; n28134
g28071 nor n28027 n28134 ; n28135
g28072 nor n28133 n28134 ; n28136
g28073 nor n28135 n28136 ; n28137
g28074 nor n28026 n28137 ; n28138
g28075 nor n28026 n28138 ; n28139
g28076 nor n28137 n28138 ; n28140
g28077 nor n28139 n28140 ; n28141
g28078 nor n27886 n27892 ; n28142
g28079 and n28141 n28142 ; n28143
g28080 nor n28141 n28142 ; n28144
g28081 nor n28143 n28144 ; n28145
g28082 and n7101 n22320 ; n28146
g28083 and n6402 n22326 ; n28147
g28084 and n6951 n22323 ; n28148
g28085 nor n28147 n28148 ; n28149
g28086 and n28146_not n28149 ; n28150
g28087 and n6397_not n28150 ; n28151
g28088 and n25270 n28150 ; n28152
g28089 nor n28151 n28152 ; n28153
g28090 and a[14] n28153_not ; n28154
g28091 and a[14]_not n28153 ; n28155
g28092 nor n28154 n28155 ; n28156
g28093 and n28145 n28156_not ; n28157
g28094 and n28145 n28157_not ; n28158
g28095 nor n28156 n28157 ; n28159
g28096 nor n28158 n28159 ; n28160
g28097 nor n28015 n28160 ; n28161
g28098 nor n28015 n28161 ; n28162
g28099 nor n28160 n28161 ; n28163
g28100 nor n28162 n28163 ; n28164
g28101 nor n28014 n28164 ; n28165
g28102 nor n28014 n28165 ; n28166
g28103 nor n28164 n28165 ; n28167
g28104 nor n28166 n28167 ; n28168
g28105 nor n27913 n27919 ; n28169
g28106 and n28168 n28169 ; n28170
g28107 nor n28168 n28169 ; n28171
g28108 nor n28170 n28171 ; n28172
g28109 and n9331 n26060 ; n28173
g28110 and n8418 n26063 ; n28174
g28111 and n8860 n26066 ; n28175
g28112 nor n28174 n28175 ; n28176
g28113 and n28173_not n28176 ; n28177
g28114 and n8421_not n28177 ; n28178
g28115 and n26088 n28177 ; n28179
g28116 nor n28178 n28179 ; n28180
g28117 and a[8] n28180_not ; n28181
g28118 and a[8]_not n28180 ; n28182
g28119 nor n28181 n28182 ; n28183
g28120 and n28172 n28183_not ; n28184
g28121 and n28172 n28184_not ; n28185
g28122 nor n28183 n28184 ; n28186
g28123 nor n28185 n28186 ; n28187
g28124 nor n28003 n28187 ; n28188
g28125 nor n28003 n28188 ; n28189
g28126 nor n28187 n28188 ; n28190
g28127 nor n28189 n28190 ; n28191
g28128 nor n28002 n28191 ; n28192
g28129 nor n28002 n28192 ; n28193
g28130 nor n28191 n28192 ; n28194
g28131 nor n28193 n28194 ; n28195
g28132 nor n27940 n27946 ; n28196
g28133 and n28195 n28196 ; n28197
g28134 nor n28195 n28196 ; n28198
g28135 nor n28197 n28198 ; n28199
g28136 nor n27959 n27963 ; n28200
g28137 and a[31]_not n97 ; n28201
g28138 nor n13438 n28201 ; n28202
g28139 and n27954 n28202_not ; n28203
g28140 and n27954_not n28202 ; n28204
g28141 nor n28203 n28204 ; n28205
g28142 and n28200 n28205_not ; n28206
g28143 and n28200_not n28205 ; n28207
g28144 nor n28206 n28207 ; n28208
g28145 and n11727 n28208_not ; n28209
g28146 and n11055 n27698 ; n28210
g28147 and n11715 n27964 ; n28211
g28148 nor n28210 n28211 ; n28212
g28149 and n28209_not n28212 ; n28213
g28150 and n11057_not n28213 ; n28214
g28151 nor n27972 n27974 ; n28215
g28152 and n27964 n28208_not ; n28216
g28153 and n27964_not n28208 ; n28217
g28154 nor n28215 n28217 ; n28218
g28155 and n28216_not n28218 ; n28219
g28156 nor n28215 n28219 ; n28220
g28157 nor n28216 n28219 ; n28221
g28158 and n28217_not n28221 ; n28222
g28159 nor n28220 n28222 ; n28223
g28160 and n28213 n28223 ; n28224
g28161 nor n28214 n28224 ; n28225
g28162 and a[2] n28225_not ; n28226
g28163 and a[2]_not n28225 ; n28227
g28164 nor n28226 n28227 ; n28228
g28165 and n28199 n28228_not ; n28229
g28166 and n28199_not n28228 ; n28230
g28167 nor n28229 n28230 ; n28231
g28168 and n27991_not n28231 ; n28232
g28169 and n27991 n28231_not ; n28233
g28170 nor n28232 n28233 ; n28234
g28171 and n27988 n28234 ; n28235
g28172 nor n27988 n28234 ; n28236
g28173 nor n28235 n28236 ; result[5]
g28174 and n71 n27698 ; n28238
g28175 and n9867 n27173 ; n28239
g28176 and n10434 n27442 ; n28240
g28177 nor n28239 n28240 ; n28241
g28178 and n28238_not n28241 ; n28242
g28179 and n9870 n27713_not ; n28243
g28180 and n28242 n28243_not ; n28244
g28181 and a[5] n28244_not ; n28245
g28182 nor n28244 n28245 ; n28246
g28183 and a[5] n28245_not ; n28247
g28184 nor n28246 n28247 ; n28248
g28185 nor n28184 n28188 ; n28249
g28186 and n7983 n26063 ; n28250
g28187 and n7291 n22315 ; n28251
g28188 and n7632 n22309 ; n28252
g28189 nor n28251 n28252 ; n28253
g28190 and n28250_not n28253 ; n28254
g28191 and n7294 n26604_not ; n28255
g28192 and n28254 n28255_not ; n28256
g28193 and a[11] n28256_not ; n28257
g28194 nor n28256 n28257 ; n28258
g28195 and a[11] n28257_not ; n28259
g28196 nor n28258 n28259 ; n28260
g28197 nor n28157 n28161 ; n28261
g28198 and n6233 n22326 ; n28262
g28199 and n5663 n22332 ; n28263
g28200 and n5939 n22329 ; n28264
g28201 nor n28263 n28264 ; n28265
g28202 and n28262_not n28265 ; n28266
g28203 and n5666 n24616_not ; n28267
g28204 and n28266 n28267_not ; n28268
g28205 and a[17] n28268_not ; n28269
g28206 nor n28268 n28269 ; n28270
g28207 and a[17] n28269_not ; n28271
g28208 nor n28270 n28271 ; n28272
g28209 nor n28130 n28134 ; n28273
g28210 and n4694 n22344 ; n28274
g28211 and n4533 n22350 ; n28275
g28212 and n4604 n22347 ; n28276
g28213 nor n28275 n28276 ; n28277
g28214 and n28274_not n28277 ; n28278
g28215 and n4536 n23642_not ; n28279
g28216 and n28278 n28279_not ; n28280
g28217 and a[23] n28280_not ; n28281
g28218 nor n28280 n28281 ; n28282
g28219 and a[23] n28281_not ; n28283
g28220 nor n28282 n28283 ; n28284
g28221 nor n28103 n28107 ; n28285
g28222 nor n28086 n28089 ; n28286
g28223 nor n28067 n28071 ; n28287
g28224 and n1550 n1693 ; n28288
g28225 and n169_not n28288 ; n28289
g28226 and n228_not n28289 ; n28290
g28227 and n191_not n28290 ; n28291
g28228 and n567_not n28291 ; n28292
g28229 and n325_not n28292 ; n28293
g28230 and n158_not n28293 ; n28294
g28231 and n297 n27522 ; n28295
g28232 and n437 n28295 ; n28296
g28233 and n3040 n28296 ; n28297
g28234 and n28294 n28297 ; n28298
g28235 and n14565 n28298 ; n28299
g28236 and n5013 n28299 ; n28300
g28237 and n15047 n28300 ; n28301
g28238 and n507 n28301 ; n28302
g28239 and n978 n28302 ; n28303
g28240 and n227 n28303 ; n28304
g28241 and n2405 n28304 ; n28305
g28242 and n116 n28305 ; n28306
g28243 and n656_not n28306 ; n28307
g28244 and n246_not n28307 ; n28308
g28245 and n372_not n28308 ; n28309
g28246 and n657_not n28309 ; n28310
g28247 and n712_not n28310 ; n28311
g28248 and n95_not n28311 ; n28312
g28249 and n886_not n28312 ; n28313
g28250 and n428_not n28313 ; n28314
g28251 and n3020 n22371 ; n28315
g28252 and n3028 n22374 ; n28316
g28253 and n3023 n22377 ; n28317
g28254 and n75 n23025 ; n28318
g28255 nor n28317 n28318 ; n28319
g28256 and n28316_not n28319 ; n28320
g28257 and n28315_not n28320 ; n28321
g28258 nor n28314 n28321 ; n28322
g28259 nor n28314 n28322 ; n28323
g28260 nor n28321 n28322 ; n28324
g28261 nor n28323 n28324 ; n28325
g28262 nor n28287 n28325 ; n28326
g28263 nor n28287 n28326 ; n28327
g28264 nor n28325 n28326 ; n28328
g28265 nor n28327 n28328 ; n28329
g28266 and n3457 n22362 ; n28330
g28267 and n3542 n22368 ; n28331
g28268 and n3606 n22365 ; n28332
g28269 nor n28331 n28332 ; n28333
g28270 and n28330_not n28333 ; n28334
g28271 and n3368_not n28334 ; n28335
g28272 and n23320 n28334 ; n28336
g28273 nor n28335 n28336 ; n28337
g28274 and a[29] n28337_not ; n28338
g28275 and a[29]_not n28337 ; n28339
g28276 nor n28338 n28339 ; n28340
g28277 nor n28329 n28340 ; n28341
g28278 and n28329 n28340 ; n28342
g28279 nor n28341 n28342 ; n28343
g28280 and n28286_not n28343 ; n28344
g28281 and n28286 n28343_not ; n28345
g28282 nor n28344 n28345 ; n28346
g28283 and n3884 n22353 ; n28347
g28284 and n3967 n22359 ; n28348
g28285 and n4046 n22356 ; n28349
g28286 nor n28348 n28349 ; n28350
g28287 and n28347_not n28350 ; n28351
g28288 and n4050_not n28351 ; n28352
g28289 and n22556 n28351 ; n28353
g28290 nor n28352 n28353 ; n28354
g28291 and a[26] n28354_not ; n28355
g28292 and a[26]_not n28354 ; n28356
g28293 nor n28355 n28356 ; n28357
g28294 and n28346 n28357_not ; n28358
g28295 and n28346_not n28357 ; n28359
g28296 nor n28358 n28359 ; n28360
g28297 and n28285_not n28360 ; n28361
g28298 and n28285 n28360_not ; n28362
g28299 nor n28361 n28362 ; n28363
g28300 and n28284_not n28363 ; n28364
g28301 nor n28284 n28364 ; n28365
g28302 and n28363 n28364_not ; n28366
g28303 nor n28365 n28366 ; n28367
g28304 nor n28111 n28117 ; n28368
g28305 and n28367 n28368 ; n28369
g28306 nor n28367 n28368 ; n28370
g28307 nor n28369 n28370 ; n28371
g28308 and n5496 n22335 ; n28372
g28309 and n4935 n22341 ; n28373
g28310 and n5407 n22338 ; n28374
g28311 nor n28373 n28374 ; n28375
g28312 and n28372_not n28375 ; n28376
g28313 and n4938_not n28376 ; n28377
g28314 and n24167 n28376 ; n28378
g28315 nor n28377 n28378 ; n28379
g28316 and a[20] n28379_not ; n28380
g28317 and a[20]_not n28379 ; n28381
g28318 nor n28380 n28381 ; n28382
g28319 and n28371 n28382_not ; n28383
g28320 and n28371_not n28382 ; n28384
g28321 nor n28383 n28384 ; n28385
g28322 and n28273_not n28385 ; n28386
g28323 and n28273 n28385_not ; n28387
g28324 nor n28386 n28387 ; n28388
g28325 and n28272_not n28388 ; n28389
g28326 nor n28272 n28389 ; n28390
g28327 and n28388 n28389_not ; n28391
g28328 nor n28390 n28391 ; n28392
g28329 nor n28138 n28144 ; n28393
g28330 and n28392 n28393 ; n28394
g28331 nor n28392 n28393 ; n28395
g28332 nor n28394 n28395 ; n28396
g28333 and n7101 n22312 ; n28397
g28334 and n6402 n22323 ; n28398
g28335 and n6951 n22320 ; n28399
g28336 nor n28398 n28399 ; n28400
g28337 and n28397_not n28400 ; n28401
g28338 and n6397_not n28401 ; n28402
g28339 and n25315 n28401 ; n28403
g28340 nor n28402 n28403 ; n28404
g28341 and a[14] n28404_not ; n28405
g28342 and a[14]_not n28404 ; n28406
g28343 nor n28405 n28406 ; n28407
g28344 and n28396 n28407_not ; n28408
g28345 and n28396_not n28407 ; n28409
g28346 nor n28408 n28409 ; n28410
g28347 and n28261_not n28410 ; n28411
g28348 and n28261 n28410_not ; n28412
g28349 nor n28411 n28412 ; n28413
g28350 and n28260_not n28413 ; n28414
g28351 nor n28260 n28414 ; n28415
g28352 and n28413 n28414_not ; n28416
g28353 nor n28415 n28416 ; n28417
g28354 nor n28165 n28171 ; n28418
g28355 and n28417 n28418 ; n28419
g28356 nor n28417 n28418 ; n28420
g28357 nor n28419 n28420 ; n28421
g28358 and n9331 n26890 ; n28422
g28359 and n8418 n26066 ; n28423
g28360 and n8860 n26060 ; n28424
g28361 nor n28423 n28424 ; n28425
g28362 and n28422_not n28425 ; n28426
g28363 and n8421_not n28426 ; n28427
g28364 and n26904 n28426 ; n28428
g28365 nor n28427 n28428 ; n28429
g28366 and a[8] n28429_not ; n28430
g28367 and a[8]_not n28429 ; n28431
g28368 nor n28430 n28431 ; n28432
g28369 and n28421 n28432_not ; n28433
g28370 and n28421_not n28432 ; n28434
g28371 nor n28433 n28434 ; n28435
g28372 and n28249_not n28435 ; n28436
g28373 and n28249 n28435_not ; n28437
g28374 nor n28436 n28437 ; n28438
g28375 and n28248_not n28438 ; n28439
g28376 nor n28248 n28439 ; n28440
g28377 and n28438 n28439_not ; n28441
g28378 nor n28440 n28441 ; n28442
g28379 nor n20821 n28208 ; n28443
g28380 and n11055 n27964 ; n28444
g28381 nor n28443 n28444 ; n28445
g28382 and n11057 n28221_not ; n28446
g28383 and n28445 n28446_not ; n28447
g28384 and a[2] n28447_not ; n28448
g28385 and a[2] n28448_not ; n28449
g28386 nor n28447 n28448 ; n28450
g28387 nor n28449 n28450 ; n28451
g28388 nor n28442 n28451 ; n28452
g28389 nor n28442 n28452 ; n28453
g28390 nor n28451 n28452 ; n28454
g28391 nor n28453 n28454 ; n28455
g28392 nor n28192 n28198 ; n28456
g28393 and n28455 n28456 ; n28457
g28394 nor n28455 n28456 ; n28458
g28395 nor n28457 n28458 ; n28459
g28396 nor n28229 n28232 ; n28460
g28397 and n28459_not n28460 ; n28461
g28398 and n28459 n28460_not ; n28462
g28399 nor n28461 n28462 ; n28463
g28400 and n28235 n28463 ; n28464
g28401 nor n28235 n28463 ; n28465
g28402 nor n28464 n28465 ; result[6]
g28403 nor n28341 n28344 ; n28467
g28404 and n75 n23006 ; n28468
g28405 and n3020 n22368 ; n28469
g28406 and n3023 n22374 ; n28470
g28407 and n3028 n22371 ; n28471
g28408 nor n28470 n28471 ; n28472
g28409 and n28469_not n28472 ; n28473
g28410 and n28468_not n28473 ; n28474
g28411 and n2115 n2423 ; n28475
g28412 and n6734 n28475 ; n28476
g28413 and n13698 n28476 ; n28477
g28414 and n2022 n28477 ; n28478
g28415 and n12944 n28478 ; n28479
g28416 and n1577 n28479 ; n28480
g28417 and n3757 n28480 ; n28481
g28418 and n1884 n28481 ; n28482
g28419 and n1574 n28482 ; n28483
g28420 and n3984 n28483 ; n28484
g28421 and n2483 n28484 ; n28485
g28422 and n1389 n28485 ; n28486
g28423 and n847_not n28486 ; n28487
g28424 and n619_not n28487 ; n28488
g28425 and n601_not n28488 ; n28489
g28426 and n537_not n28489 ; n28490
g28427 and n157_not n28490 ; n28491
g28428 and n531_not n28491 ; n28492
g28429 nor n15031 n28208 ; n28493
g28430 and a[2] n28493_not ; n28494
g28431 and a[2]_not n28493 ; n28495
g28432 nor n28494 n28495 ; n28496
g28433 nor n28492 n28496 ; n28497
g28434 and n28492 n28496 ; n28498
g28435 nor n28474 n28498 ; n28499
g28436 and n28497_not n28499 ; n28500
g28437 nor n28474 n28500 ; n28501
g28438 nor n28497 n28500 ; n28502
g28439 and n28498_not n28502 ; n28503
g28440 nor n28501 n28503 ; n28504
g28441 nor n28322 n28326 ; n28505
g28442 and n28504 n28505 ; n28506
g28443 nor n28504 n28505 ; n28507
g28444 nor n28506 n28507 ; n28508
g28445 and n3457 n22359 ; n28509
g28446 and n3542 n22365 ; n28510
g28447 and n3606 n22362 ; n28511
g28448 nor n28510 n28511 ; n28512
g28449 and n28509_not n28512 ; n28513
g28450 and n3368_not n28513 ; n28514
g28451 and n23368_not n28513 ; n28515
g28452 nor n28514 n28515 ; n28516
g28453 and a[29] n28516_not ; n28517
g28454 and a[29]_not n28516 ; n28518
g28455 nor n28517 n28518 ; n28519
g28456 and n28508 n28519_not ; n28520
g28457 and n28508_not n28519 ; n28521
g28458 nor n28520 n28521 ; n28522
g28459 and n28467_not n28522 ; n28523
g28460 and n28467 n28522_not ; n28524
g28461 nor n28523 n28524 ; n28525
g28462 and n3884 n22350 ; n28526
g28463 and n3967 n22356 ; n28527
g28464 and n4046 n22353 ; n28528
g28465 nor n28527 n28528 ; n28529
g28466 and n28526_not n28529 ; n28530
g28467 and n4050 n23672 ; n28531
g28468 and n28530 n28531_not ; n28532
g28469 and a[26] n28532_not ; n28533
g28470 and a[26] n28533_not ; n28534
g28471 nor n28532 n28533 ; n28535
g28472 nor n28534 n28535 ; n28536
g28473 and n28525 n28536_not ; n28537
g28474 and n28525 n28537_not ; n28538
g28475 nor n28536 n28537 ; n28539
g28476 nor n28538 n28539 ; n28540
g28477 nor n28358 n28361 ; n28541
g28478 and n28540 n28541 ; n28542
g28479 nor n28540 n28541 ; n28543
g28480 nor n28542 n28543 ; n28544
g28481 and n4694 n22341 ; n28545
g28482 and n4533 n22347 ; n28546
g28483 and n4604 n22344 ; n28547
g28484 nor n28546 n28547 ; n28548
g28485 and n28545_not n28548 ; n28549
g28486 and n4536 n24142 ; n28550
g28487 and n28549 n28550_not ; n28551
g28488 and a[23] n28551_not ; n28552
g28489 and a[23] n28552_not ; n28553
g28490 nor n28551 n28552 ; n28554
g28491 nor n28553 n28554 ; n28555
g28492 and n28544 n28555_not ; n28556
g28493 and n28544 n28556_not ; n28557
g28494 nor n28555 n28556 ; n28558
g28495 nor n28557 n28558 ; n28559
g28496 nor n28364 n28370 ; n28560
g28497 and n28559 n28560 ; n28561
g28498 nor n28559 n28560 ; n28562
g28499 nor n28561 n28562 ; n28563
g28500 and n5496 n22332 ; n28564
g28501 and n4935 n22338 ; n28565
g28502 and n5407 n22335 ; n28566
g28503 nor n28565 n28566 ; n28567
g28504 and n28564_not n28567 ; n28568
g28505 and n4938 n22542 ; n28569
g28506 and n28568 n28569_not ; n28570
g28507 and a[20] n28570_not ; n28571
g28508 and a[20] n28571_not ; n28572
g28509 nor n28570 n28571 ; n28573
g28510 nor n28572 n28573 ; n28574
g28511 and n28563 n28574_not ; n28575
g28512 and n28563 n28575_not ; n28576
g28513 nor n28574 n28575 ; n28577
g28514 nor n28576 n28577 ; n28578
g28515 nor n28383 n28386 ; n28579
g28516 and n28578 n28579 ; n28580
g28517 nor n28578 n28579 ; n28581
g28518 nor n28580 n28581 ; n28582
g28519 and n6233 n22323 ; n28583
g28520 and n5663 n22329 ; n28584
g28521 and n5939 n22326 ; n28585
g28522 nor n28584 n28585 ; n28586
g28523 and n28583_not n28586 ; n28587
g28524 and n5666 n24599 ; n28588
g28525 and n28587 n28588_not ; n28589
g28526 and a[17] n28589_not ; n28590
g28527 and a[17] n28590_not ; n28591
g28528 nor n28589 n28590 ; n28592
g28529 nor n28591 n28592 ; n28593
g28530 and n28582 n28593_not ; n28594
g28531 and n28582 n28594_not ; n28595
g28532 nor n28593 n28594 ; n28596
g28533 nor n28595 n28596 ; n28597
g28534 nor n28389 n28395 ; n28598
g28535 and n28597 n28598 ; n28599
g28536 nor n28597 n28598 ; n28600
g28537 nor n28599 n28600 ; n28601
g28538 and n7101 n22315 ; n28602
g28539 and n6402 n22320 ; n28603
g28540 and n6951 n22312 ; n28604
g28541 nor n28603 n28604 ; n28605
g28542 and n28602_not n28605 ; n28606
g28543 and n6397 n25294 ; n28607
g28544 and n28606 n28607_not ; n28608
g28545 and a[14] n28608_not ; n28609
g28546 and a[14] n28609_not ; n28610
g28547 nor n28608 n28609 ; n28611
g28548 nor n28610 n28611 ; n28612
g28549 and n28601 n28612_not ; n28613
g28550 and n28601 n28613_not ; n28614
g28551 nor n28612 n28613 ; n28615
g28552 nor n28614 n28615 ; n28616
g28553 nor n28408 n28411 ; n28617
g28554 and n28616 n28617 ; n28618
g28555 nor n28616 n28617 ; n28619
g28556 nor n28618 n28619 ; n28620
g28557 and n7983 n26066 ; n28621
g28558 and n7291 n22309 ; n28622
g28559 and n7632 n26063 ; n28623
g28560 nor n28622 n28623 ; n28624
g28561 and n28621_not n28624 ; n28625
g28562 and n7294 n26624_not ; n28626
g28563 and n28625 n28626_not ; n28627
g28564 and a[11] n28627_not ; n28628
g28565 and a[11] n28628_not ; n28629
g28566 nor n28627 n28628 ; n28630
g28567 nor n28629 n28630 ; n28631
g28568 and n28620 n28631_not ; n28632
g28569 and n28620 n28632_not ; n28633
g28570 nor n28631 n28632 ; n28634
g28571 nor n28633 n28634 ; n28635
g28572 nor n28414 n28420 ; n28636
g28573 and n28635 n28636 ; n28637
g28574 nor n28635 n28636 ; n28638
g28575 nor n28637 n28638 ; n28639
g28576 and n9331 n27173 ; n28640
g28577 and n8418 n26060 ; n28641
g28578 and n8860 n26890 ; n28642
g28579 nor n28641 n28642 ; n28643
g28580 and n28640_not n28643 ; n28644
g28581 and n8421 n27185 ; n28645
g28582 and n28644 n28645_not ; n28646
g28583 and a[8] n28646_not ; n28647
g28584 and a[8] n28647_not ; n28648
g28585 nor n28646 n28647 ; n28649
g28586 nor n28648 n28649 ; n28650
g28587 and n28639 n28650_not ; n28651
g28588 and n28639 n28651_not ; n28652
g28589 nor n28650 n28651 ; n28653
g28590 nor n28652 n28653 ; n28654
g28591 nor n28433 n28436 ; n28655
g28592 and n28654 n28655 ; n28656
g28593 nor n28654 n28655 ; n28657
g28594 nor n28656 n28657 ; n28658
g28595 and n71 n27964 ; n28659
g28596 and n9867 n27442 ; n28660
g28597 and n10434 n27698 ; n28661
g28598 nor n28660 n28661 ; n28662
g28599 and n28659_not n28662 ; n28663
g28600 and n9870 n27976 ; n28664
g28601 and n28663 n28664_not ; n28665
g28602 and a[5] n28665_not ; n28666
g28603 and a[5] n28666_not ; n28667
g28604 nor n28665 n28666 ; n28668
g28605 nor n28667 n28668 ; n28669
g28606 and n28658 n28669_not ; n28670
g28607 and n28658 n28670_not ; n28671
g28608 nor n28669 n28670 ; n28672
g28609 nor n28671 n28672 ; n28673
g28610 nor n28439 n28452 ; n28674
g28611 and n28673 n28674 ; n28675
g28612 nor n28673 n28674 ; n28676
g28613 nor n28675 n28676 ; n28677
g28614 nor n28458 n28462 ; n28678
g28615 and n28677_not n28678 ; n28679
g28616 and n28677 n28678_not ; n28680
g28617 nor n28679 n28680 ; n28681
g28618 and n28464 n28681 ; n28682
g28619 nor n28464 n28681 ; n28683
g28620 nor n28682 n28683 ; result[7]
g28621 and n720 n16020 ; n28685
g28622 and n301_not n28685 ; n28686
g28623 and n571_not n28686 ; n28687
g28624 and n886_not n28687 ; n28688
g28625 and n1347 n23251 ; n28689
g28626 and n1424 n28689 ; n28690
g28627 and n2410 n28690 ; n28691
g28628 and n28688 n28691 ; n28692
g28629 and n16067 n28692 ; n28693
g28630 and n1313 n28693 ; n28694
g28631 and n1782 n28694 ; n28695
g28632 and n869 n28695 ; n28696
g28633 and n979 n28696 ; n28697
g28634 and n399 n28697 ; n28698
g28635 and n2583 n28698 ; n28699
g28636 and n2088 n28699 ; n28700
g28637 and n3163 n28700 ; n28701
g28638 and n279 n28701 ; n28702
g28639 and n121_not n28702 ; n28703
g28640 and n283_not n28703 ; n28704
g28641 and n666_not n28704 ; n28705
g28642 and n363_not n28705 ; n28706
g28643 nor n28496 n28706 ; n28707
g28644 and n28496 n28706 ; n28708
g28645 nor n28502 n28708 ; n28709
g28646 and n28707_not n28709 ; n28710
g28647 nor n28502 n28710 ; n28711
g28648 nor n28707 n28710 ; n28712
g28649 and n28708_not n28712 ; n28713
g28650 nor n28711 n28713 ; n28714
g28651 and n75 n22993_not ; n28715
g28652 and n3020 n22365 ; n28716
g28653 and n3023 n22371 ; n28717
g28654 and n3028 n22368 ; n28718
g28655 nor n28717 n28718 ; n28719
g28656 and n28716_not n28719 ; n28720
g28657 and n28715_not n28720 ; n28721
g28658 nor n28714 n28721 ; n28722
g28659 nor n28714 n28722 ; n28723
g28660 nor n28721 n28722 ; n28724
g28661 nor n28723 n28724 ; n28725
g28662 nor n28507 n28520 ; n28726
g28663 and n28725 n28726 ; n28727
g28664 nor n28725 n28726 ; n28728
g28665 nor n28727 n28728 ; n28729
g28666 and n3457 n22356 ; n28730
g28667 and n3542 n22362 ; n28731
g28668 and n3606 n22359 ; n28732
g28669 nor n28731 n28732 ; n28733
g28670 and n28730_not n28733 ; n28734
g28671 and n3368 n23345_not ; n28735
g28672 and n28734 n28735_not ; n28736
g28673 and a[29] n28736_not ; n28737
g28674 and a[29] n28737_not ; n28738
g28675 nor n28736 n28737 ; n28739
g28676 nor n28738 n28739 ; n28740
g28677 and n28729 n28740_not ; n28741
g28678 and n28729 n28741_not ; n28742
g28679 nor n28740 n28741 ; n28743
g28680 nor n28742 n28743 ; n28744
g28681 and n3884 n22347 ; n28745
g28682 and n3967 n22353 ; n28746
g28683 and n4046 n22350 ; n28747
g28684 nor n28746 n28747 ; n28748
g28685 and n28745_not n28748 ; n28749
g28686 and n4050 n23659_not ; n28750
g28687 and n28749 n28750_not ; n28751
g28688 and a[26] n28751_not ; n28752
g28689 and a[26] n28752_not ; n28753
g28690 nor n28751 n28752 ; n28754
g28691 nor n28753 n28754 ; n28755
g28692 nor n28744 n28755 ; n28756
g28693 nor n28744 n28756 ; n28757
g28694 nor n28755 n28756 ; n28758
g28695 nor n28757 n28758 ; n28759
g28696 nor n28523 n28537 ; n28760
g28697 and n28759 n28760 ; n28761
g28698 nor n28759 n28760 ; n28762
g28699 nor n28761 n28762 ; n28763
g28700 and n4694 n22338 ; n28764
g28701 and n4533 n22344 ; n28765
g28702 and n4604 n22341 ; n28766
g28703 nor n28765 n28766 ; n28767
g28704 and n28764_not n28767 ; n28768
g28705 and n4536 n24188_not ; n28769
g28706 and n28768 n28769_not ; n28770
g28707 and a[23] n28770_not ; n28771
g28708 and a[23] n28771_not ; n28772
g28709 nor n28770 n28771 ; n28773
g28710 nor n28772 n28773 ; n28774
g28711 and n28763 n28774_not ; n28775
g28712 and n28763 n28775_not ; n28776
g28713 nor n28774 n28775 ; n28777
g28714 nor n28776 n28777 ; n28778
g28715 nor n28543 n28556 ; n28779
g28716 and n28778 n28779 ; n28780
g28717 nor n28778 n28779 ; n28781
g28718 nor n28780 n28781 ; n28782
g28719 and n5496 n22329 ; n28783
g28720 and n4935 n22335 ; n28784
g28721 and n5407 n22332 ; n28785
g28722 nor n28784 n28785 ; n28786
g28723 and n28783_not n28786 ; n28787
g28724 and n4938 n24633_not ; n28788
g28725 and n28787 n28788_not ; n28789
g28726 and a[20] n28789_not ; n28790
g28727 and a[20] n28790_not ; n28791
g28728 nor n28789 n28790 ; n28792
g28729 nor n28791 n28792 ; n28793
g28730 and n28782 n28793_not ; n28794
g28731 and n28782 n28794_not ; n28795
g28732 nor n28793 n28794 ; n28796
g28733 nor n28795 n28796 ; n28797
g28734 nor n28562 n28575 ; n28798
g28735 and n28797 n28798 ; n28799
g28736 nor n28797 n28798 ; n28800
g28737 nor n28799 n28800 ; n28801
g28738 and n6233 n22320 ; n28802
g28739 and n5663 n22326 ; n28803
g28740 and n5939 n22323 ; n28804
g28741 nor n28803 n28804 ; n28805
g28742 and n28802_not n28805 ; n28806
g28743 and n5666 n25270_not ; n28807
g28744 and n28806 n28807_not ; n28808
g28745 and a[17] n28808_not ; n28809
g28746 and a[17] n28809_not ; n28810
g28747 nor n28808 n28809 ; n28811
g28748 nor n28810 n28811 ; n28812
g28749 and n28801 n28812_not ; n28813
g28750 and n28801 n28813_not ; n28814
g28751 nor n28812 n28813 ; n28815
g28752 nor n28814 n28815 ; n28816
g28753 nor n28581 n28594 ; n28817
g28754 and n28816 n28817 ; n28818
g28755 nor n28816 n28817 ; n28819
g28756 nor n28818 n28819 ; n28820
g28757 and n7101 n22309 ; n28821
g28758 and n6402 n22312 ; n28822
g28759 and n6951 n22315 ; n28823
g28760 nor n28822 n28823 ; n28824
g28761 and n28821_not n28824 ; n28825
g28762 and n6397 n22529_not ; n28826
g28763 and n28825 n28826_not ; n28827
g28764 and a[14] n28827_not ; n28828
g28765 and a[14] n28828_not ; n28829
g28766 nor n28827 n28828 ; n28830
g28767 nor n28829 n28830 ; n28831
g28768 and n28820 n28831_not ; n28832
g28769 and n28820 n28832_not ; n28833
g28770 nor n28831 n28832 ; n28834
g28771 nor n28833 n28834 ; n28835
g28772 nor n28600 n28613 ; n28836
g28773 and n28835 n28836 ; n28837
g28774 nor n28835 n28836 ; n28838
g28775 nor n28837 n28838 ; n28839
g28776 and n7983 n26060 ; n28840
g28777 and n7291 n26063 ; n28841
g28778 and n7632 n26066 ; n28842
g28779 nor n28841 n28842 ; n28843
g28780 and n28840_not n28843 ; n28844
g28781 and n7294 n26088_not ; n28845
g28782 and n28844 n28845_not ; n28846
g28783 and a[11] n28846_not ; n28847
g28784 and a[11] n28847_not ; n28848
g28785 nor n28846 n28847 ; n28849
g28786 nor n28848 n28849 ; n28850
g28787 and n28839 n28850_not ; n28851
g28788 and n28839 n28851_not ; n28852
g28789 nor n28850 n28851 ; n28853
g28790 nor n28852 n28853 ; n28854
g28791 nor n28619 n28632 ; n28855
g28792 and n28854 n28855 ; n28856
g28793 nor n28854 n28855 ; n28857
g28794 nor n28856 n28857 ; n28858
g28795 and n9331 n27442 ; n28859
g28796 and n8418 n26890 ; n28860
g28797 and n8860 n27173 ; n28861
g28798 nor n28860 n28861 ; n28862
g28799 and n28859_not n28862 ; n28863
g28800 and n8421 n27455 ; n28864
g28801 and n28863 n28864_not ; n28865
g28802 and a[8] n28865_not ; n28866
g28803 and a[8] n28866_not ; n28867
g28804 nor n28865 n28866 ; n28868
g28805 nor n28867 n28868 ; n28869
g28806 and n28858 n28869_not ; n28870
g28807 and n28858 n28870_not ; n28871
g28808 nor n28869 n28870 ; n28872
g28809 nor n28871 n28872 ; n28873
g28810 nor n28638 n28651 ; n28874
g28811 and n28873 n28874 ; n28875
g28812 nor n28873 n28874 ; n28876
g28813 nor n28875 n28876 ; n28877
g28814 and n71 n28208_not ; n28878
g28815 and n9867 n27698 ; n28879
g28816 and n10434 n27964 ; n28880
g28817 nor n28879 n28880 ; n28881
g28818 and n28878_not n28881 ; n28882
g28819 and n9870 n28223_not ; n28883
g28820 and n28882 n28883_not ; n28884
g28821 and a[5] n28884_not ; n28885
g28822 and a[5] n28885_not ; n28886
g28823 nor n28884 n28885 ; n28887
g28824 nor n28886 n28887 ; n28888
g28825 and n28877 n28888_not ; n28889
g28826 and n28877 n28889_not ; n28890
g28827 nor n28888 n28889 ; n28891
g28828 nor n28890 n28891 ; n28892
g28829 nor n28657 n28670 ; n28893
g28830 and n28892 n28893 ; n28894
g28831 nor n28892 n28893 ; n28895
g28832 nor n28894 n28895 ; n28896
g28833 nor n28676 n28680 ; n28897
g28834 and n28896_not n28897 ; n28898
g28835 and n28896 n28897_not ; n28899
g28836 nor n28898 n28899 ; n28900
g28837 and n28682 n28900 ; n28901
g28838 nor n28682 n28900 ; n28902
g28839 nor n28901 n28902 ; result[8]
g28840 and n2424 n15286 ; n28904
g28841 and n2704 n28904 ; n28905
g28842 and n1103 n28905 ; n28906
g28843 and n3685 n28906 ; n28907
g28844 and n5199 n28907 ; n28908
g28845 and n770 n28908 ; n28909
g28846 and n415 n28909 ; n28910
g28847 and n1182 n28910 ; n28911
g28848 and n2443 n28911 ; n28912
g28849 and n937 n28912 ; n28913
g28850 and n2167 n28913 ; n28914
g28851 and n276_not n28914 ; n28915
g28852 and n1011_not n28915 ; n28916
g28853 and n255_not n28916 ; n28917
g28854 and n150_not n28917 ; n28918
g28855 and n295_not n28918 ; n28919
g28856 nor n28496 n28919 ; n28920
g28857 and n28496 n28919 ; n28921
g28858 nor n28712 n28921 ; n28922
g28859 and n28920_not n28922 ; n28923
g28860 nor n28712 n28923 ; n28924
g28861 nor n28920 n28923 ; n28925
g28862 and n28921_not n28925 ; n28926
g28863 nor n28924 n28926 ; n28927
g28864 and n75 n23320_not ; n28928
g28865 and n3020 n22362 ; n28929
g28866 and n3023 n22368 ; n28930
g28867 and n3028 n22365 ; n28931
g28868 nor n28930 n28931 ; n28932
g28869 and n28929_not n28932 ; n28933
g28870 and n28928_not n28933 ; n28934
g28871 nor n28927 n28934 ; n28935
g28872 nor n28927 n28935 ; n28936
g28873 nor n28934 n28935 ; n28937
g28874 nor n28936 n28937 ; n28938
g28875 nor n28722 n28728 ; n28939
g28876 and n28938 n28939 ; n28940
g28877 nor n28938 n28939 ; n28941
g28878 nor n28940 n28941 ; n28942
g28879 and n3457 n22353 ; n28943
g28880 and n3542 n22359 ; n28944
g28881 and n3606 n22356 ; n28945
g28882 nor n28944 n28945 ; n28946
g28883 and n28943_not n28946 ; n28947
g28884 and n3368 n22556_not ; n28948
g28885 and n28947 n28948_not ; n28949
g28886 and a[29] n28949_not ; n28950
g28887 and a[29] n28950_not ; n28951
g28888 nor n28949 n28950 ; n28952
g28889 nor n28951 n28952 ; n28953
g28890 and n28942 n28953_not ; n28954
g28891 and n28942 n28954_not ; n28955
g28892 nor n28953 n28954 ; n28956
g28893 nor n28955 n28956 ; n28957
g28894 and n3884 n22344 ; n28958
g28895 and n3967 n22350 ; n28959
g28896 and n4046 n22347 ; n28960
g28897 nor n28959 n28960 ; n28961
g28898 and n28958_not n28961 ; n28962
g28899 and n4050 n23642_not ; n28963
g28900 and n28962 n28963_not ; n28964
g28901 and a[26] n28964_not ; n28965
g28902 and a[26] n28965_not ; n28966
g28903 nor n28964 n28965 ; n28967
g28904 nor n28966 n28967 ; n28968
g28905 nor n28957 n28968 ; n28969
g28906 nor n28957 n28969 ; n28970
g28907 nor n28968 n28969 ; n28971
g28908 nor n28970 n28971 ; n28972
g28909 nor n28741 n28756 ; n28973
g28910 and n28972 n28973 ; n28974
g28911 nor n28972 n28973 ; n28975
g28912 nor n28974 n28975 ; n28976
g28913 and n4694 n22335 ; n28977
g28914 and n4533 n22341 ; n28978
g28915 and n4604 n22338 ; n28979
g28916 nor n28978 n28979 ; n28980
g28917 and n28977_not n28980 ; n28981
g28918 and n4536 n24167_not ; n28982
g28919 and n28981 n28982_not ; n28983
g28920 and a[23] n28983_not ; n28984
g28921 and a[23] n28984_not ; n28985
g28922 nor n28983 n28984 ; n28986
g28923 nor n28985 n28986 ; n28987
g28924 and n28976 n28987_not ; n28988
g28925 and n28976 n28988_not ; n28989
g28926 nor n28987 n28988 ; n28990
g28927 nor n28989 n28990 ; n28991
g28928 nor n28762 n28775 ; n28992
g28929 and n28991 n28992 ; n28993
g28930 nor n28991 n28992 ; n28994
g28931 nor n28993 n28994 ; n28995
g28932 and n5496 n22326 ; n28996
g28933 and n4935 n22332 ; n28997
g28934 and n5407 n22329 ; n28998
g28935 nor n28997 n28998 ; n28999
g28936 and n28996_not n28999 ; n29000
g28937 and n4938 n24616_not ; n29001
g28938 and n29000 n29001_not ; n29002
g28939 and a[20] n29002_not ; n29003
g28940 and a[20] n29003_not ; n29004
g28941 nor n29002 n29003 ; n29005
g28942 nor n29004 n29005 ; n29006
g28943 and n28995 n29006_not ; n29007
g28944 and n28995 n29007_not ; n29008
g28945 nor n29006 n29007 ; n29009
g28946 nor n29008 n29009 ; n29010
g28947 nor n28781 n28794 ; n29011
g28948 and n29010 n29011 ; n29012
g28949 nor n29010 n29011 ; n29013
g28950 nor n29012 n29013 ; n29014
g28951 and n6233 n22312 ; n29015
g28952 and n5663 n22323 ; n29016
g28953 and n5939 n22320 ; n29017
g28954 nor n29016 n29017 ; n29018
g28955 and n29015_not n29018 ; n29019
g28956 and n5666 n25315_not ; n29020
g28957 and n29019 n29020_not ; n29021
g28958 and a[17] n29021_not ; n29022
g28959 and a[17] n29022_not ; n29023
g28960 nor n29021 n29022 ; n29024
g28961 nor n29023 n29024 ; n29025
g28962 and n29014 n29025_not ; n29026
g28963 and n29014 n29026_not ; n29027
g28964 nor n29025 n29026 ; n29028
g28965 nor n29027 n29028 ; n29029
g28966 nor n28800 n28813 ; n29030
g28967 and n29029 n29030 ; n29031
g28968 nor n29029 n29030 ; n29032
g28969 nor n29031 n29032 ; n29033
g28970 and n7101 n26063 ; n29034
g28971 and n6402 n22315 ; n29035
g28972 and n6951 n22309 ; n29036
g28973 nor n29035 n29036 ; n29037
g28974 and n29034_not n29037 ; n29038
g28975 and n6397 n26604_not ; n29039
g28976 and n29038 n29039_not ; n29040
g28977 and a[14] n29040_not ; n29041
g28978 and a[14] n29041_not ; n29042
g28979 nor n29040 n29041 ; n29043
g28980 nor n29042 n29043 ; n29044
g28981 and n29033 n29044_not ; n29045
g28982 and n29033 n29045_not ; n29046
g28983 nor n29044 n29045 ; n29047
g28984 nor n29046 n29047 ; n29048
g28985 nor n28819 n28832 ; n29049
g28986 and n29048 n29049 ; n29050
g28987 nor n29048 n29049 ; n29051
g28988 nor n29050 n29051 ; n29052
g28989 and n7983 n26890 ; n29053
g28990 and n7291 n26066 ; n29054
g28991 and n7632 n26060 ; n29055
g28992 nor n29054 n29055 ; n29056
g28993 and n29053_not n29056 ; n29057
g28994 and n7294 n26904_not ; n29058
g28995 and n29057 n29058_not ; n29059
g28996 and a[11] n29059_not ; n29060
g28997 and a[11] n29060_not ; n29061
g28998 nor n29059 n29060 ; n29062
g28999 nor n29061 n29062 ; n29063
g29000 and n29052 n29063_not ; n29064
g29001 and n29052 n29064_not ; n29065
g29002 nor n29063 n29064 ; n29066
g29003 nor n29065 n29066 ; n29067
g29004 nor n28838 n28851 ; n29068
g29005 and n29067 n29068 ; n29069
g29006 nor n29067 n29068 ; n29070
g29007 nor n29069 n29070 ; n29071
g29008 and n9331 n27698 ; n29072
g29009 and n8418 n27173 ; n29073
g29010 and n8860 n27442 ; n29074
g29011 nor n29073 n29074 ; n29075
g29012 and n29072_not n29075 ; n29076
g29013 and n8421 n27713_not ; n29077
g29014 and n29076 n29077_not ; n29078
g29015 and a[8] n29078_not ; n29079
g29016 and a[8] n29079_not ; n29080
g29017 nor n29078 n29079 ; n29081
g29018 nor n29080 n29081 ; n29082
g29019 and n29071 n29082_not ; n29083
g29020 and n29071 n29083_not ; n29084
g29021 nor n29082 n29083 ; n29085
g29022 nor n29084 n29085 ; n29086
g29023 nor n28857 n28870 ; n29087
g29024 nor n15076 n28208 ; n29088
g29025 and n9867 n27964 ; n29089
g29026 nor n29088 n29089 ; n29090
g29027 and n9870_not n29090 ; n29091
g29028 and n28221 n29090 ; n29092
g29029 nor n29091 n29092 ; n29093
g29030 and a[5] n29093_not ; n29094
g29031 and a[5]_not n29093 ; n29095
g29032 nor n29094 n29095 ; n29096
g29033 nor n29087 n29096 ; n29097
g29034 and n29087 n29096 ; n29098
g29035 nor n29097 n29098 ; n29099
g29036 and n29086_not n29099 ; n29100
g29037 nor n29086 n29100 ; n29101
g29038 and n29099 n29100_not ; n29102
g29039 nor n29101 n29102 ; n29103
g29040 nor n28876 n28889 ; n29104
g29041 and n29103 n29104 ; n29105
g29042 nor n29103 n29104 ; n29106
g29043 nor n29105 n29106 ; n29107
g29044 nor n28895 n28899 ; n29108
g29045 and n29107_not n29108 ; n29109
g29046 and n29107 n29108_not ; n29110
g29047 nor n29109 n29110 ; n29111
g29048 and n28901 n29111 ; n29112
g29049 nor n28901 n29111 ; n29113
g29050 nor n29112 n29113 ; result[9]
g29051 nor n29106 n29110 ; n29115
g29052 nor n29097 n29100 ; n29116
g29053 nor n28935 n28941 ; n29117
g29054 and n1859 n4335 ; n29118
g29055 and n1073 n29118 ; n29119
g29056 and n4357 n29119 ; n29120
g29057 and n960 n29120 ; n29121
g29058 and n526 n29121 ; n29122
g29059 and n13826 n29122 ; n29123
g29060 and n3057 n29123 ; n29124
g29061 and n2467 n29124 ; n29125
g29062 and n3886 n29125 ; n29126
g29063 and n1761 n29126 ; n29127
g29064 and n22748 n29127 ; n29128
g29065 and n746_not n29128 ; n29129
g29066 and n280_not n29129 ; n29130
g29067 and n119_not n29130 ; n29131
g29068 and n358_not n29131 ; n29132
g29069 and n28496 n29132 ; n29133
g29070 nor n28496 n29132 ; n29134
g29071 nor n29133 n29134 ; n29135
g29072 nor n15078 n28208 ; n29136
g29073 and a[5]_not n29136 ; n29137
g29074 and a[5] n29136_not ; n29138
g29075 nor n29135 n29138 ; n29139
g29076 and n29137_not n29139 ; n29140
g29077 nor n29135 n29140 ; n29141
g29078 nor n29138 n29140 ; n29142
g29079 and n29137_not n29142 ; n29143
g29080 nor n29141 n29143 ; n29144
g29081 and n28925_not n29144 ; n29145
g29082 and n28925 n29144_not ; n29146
g29083 nor n29145 n29146 ; n29147
g29084 and n75 n23368 ; n29148
g29085 and n3020 n22359 ; n29149
g29086 and n3023 n22365 ; n29150
g29087 and n3028 n22362 ; n29151
g29088 nor n29150 n29151 ; n29152
g29089 and n29149_not n29152 ; n29153
g29090 and n29148_not n29153 ; n29154
g29091 nor n29147 n29154 ; n29155
g29092 and n29147 n29154 ; n29156
g29093 nor n29155 n29156 ; n29157
g29094 and n29117 n29157_not ; n29158
g29095 and n29117_not n29157 ; n29159
g29096 nor n29158 n29159 ; n29160
g29097 and n3457 n22350 ; n29161
g29098 and n3542 n22356 ; n29162
g29099 and n3606 n22353 ; n29163
g29100 nor n29162 n29163 ; n29164
g29101 and n29161_not n29164 ; n29165
g29102 and n3368 n23672 ; n29166
g29103 and n29165 n29166_not ; n29167
g29104 and a[29] n29167_not ; n29168
g29105 and a[29] n29168_not ; n29169
g29106 nor n29167 n29168 ; n29170
g29107 nor n29169 n29170 ; n29171
g29108 and n29160 n29171_not ; n29172
g29109 and n29160 n29172_not ; n29173
g29110 nor n29171 n29172 ; n29174
g29111 nor n29173 n29174 ; n29175
g29112 and n3884 n22341 ; n29176
g29113 and n3967 n22347 ; n29177
g29114 and n4046 n22344 ; n29178
g29115 nor n29177 n29178 ; n29179
g29116 and n29176_not n29179 ; n29180
g29117 and n4050 n24142 ; n29181
g29118 and n29180 n29181_not ; n29182
g29119 and a[26] n29182_not ; n29183
g29120 and a[26] n29183_not ; n29184
g29121 nor n29182 n29183 ; n29185
g29122 nor n29184 n29185 ; n29186
g29123 nor n29175 n29186 ; n29187
g29124 nor n29175 n29187 ; n29188
g29125 nor n29186 n29187 ; n29189
g29126 nor n29188 n29189 ; n29190
g29127 nor n28954 n28969 ; n29191
g29128 and n29190 n29191 ; n29192
g29129 nor n29190 n29191 ; n29193
g29130 nor n29192 n29193 ; n29194
g29131 and n4694 n22332 ; n29195
g29132 and n4533 n22338 ; n29196
g29133 and n4604 n22335 ; n29197
g29134 nor n29196 n29197 ; n29198
g29135 and n29195_not n29198 ; n29199
g29136 and n4536 n22542 ; n29200
g29137 and n29199 n29200_not ; n29201
g29138 and a[23] n29201_not ; n29202
g29139 and a[23] n29202_not ; n29203
g29140 nor n29201 n29202 ; n29204
g29141 nor n29203 n29204 ; n29205
g29142 and n29194 n29205_not ; n29206
g29143 and n29194 n29206_not ; n29207
g29144 nor n29205 n29206 ; n29208
g29145 nor n29207 n29208 ; n29209
g29146 nor n28975 n28988 ; n29210
g29147 and n29209 n29210 ; n29211
g29148 nor n29209 n29210 ; n29212
g29149 nor n29211 n29212 ; n29213
g29150 and n5496 n22323 ; n29214
g29151 and n4935 n22329 ; n29215
g29152 and n5407 n22326 ; n29216
g29153 nor n29215 n29216 ; n29217
g29154 and n29214_not n29217 ; n29218
g29155 and n4938 n24599 ; n29219
g29156 and n29218 n29219_not ; n29220
g29157 and a[20] n29220_not ; n29221
g29158 and a[20] n29221_not ; n29222
g29159 nor n29220 n29221 ; n29223
g29160 nor n29222 n29223 ; n29224
g29161 and n29213 n29224_not ; n29225
g29162 and n29213 n29225_not ; n29226
g29163 nor n29224 n29225 ; n29227
g29164 nor n29226 n29227 ; n29228
g29165 nor n28994 n29007 ; n29229
g29166 and n29228 n29229 ; n29230
g29167 nor n29228 n29229 ; n29231
g29168 nor n29230 n29231 ; n29232
g29169 and n6233 n22315 ; n29233
g29170 and n5663 n22320 ; n29234
g29171 and n5939 n22312 ; n29235
g29172 nor n29234 n29235 ; n29236
g29173 and n29233_not n29236 ; n29237
g29174 and n5666 n25294 ; n29238
g29175 and n29237 n29238_not ; n29239
g29176 and a[17] n29239_not ; n29240
g29177 and a[17] n29240_not ; n29241
g29178 nor n29239 n29240 ; n29242
g29179 nor n29241 n29242 ; n29243
g29180 and n29232 n29243_not ; n29244
g29181 and n29232 n29244_not ; n29245
g29182 nor n29243 n29244 ; n29246
g29183 nor n29245 n29246 ; n29247
g29184 nor n29013 n29026 ; n29248
g29185 and n29247 n29248 ; n29249
g29186 nor n29247 n29248 ; n29250
g29187 nor n29249 n29250 ; n29251
g29188 nor n29032 n29045 ; n29252
g29189 and n7101 n26066 ; n29253
g29190 and n6402 n22309 ; n29254
g29191 and n6951 n26063 ; n29255
g29192 nor n29254 n29255 ; n29256
g29193 and n29253_not n29256 ; n29257
g29194 and n6397 n26624_not ; n29258
g29195 and n29257 n29258_not ; n29259
g29196 and a[14] n29259_not ; n29260
g29197 and a[14] n29260_not ; n29261
g29198 nor n29259 n29260 ; n29262
g29199 nor n29261 n29262 ; n29263
g29200 nor n29252 n29263 ; n29264
g29201 nor n29252 n29264 ; n29265
g29202 nor n29263 n29264 ; n29266
g29203 nor n29265 n29266 ; n29267
g29204 and n29251_not n29267 ; n29268
g29205 and n29251 n29267_not ; n29269
g29206 nor n29268 n29269 ; n29270
g29207 and n7983 n27173 ; n29271
g29208 and n7291 n26060 ; n29272
g29209 and n7632 n26890 ; n29273
g29210 nor n29272 n29273 ; n29274
g29211 and n29271_not n29274 ; n29275
g29212 and n7294 n27185 ; n29276
g29213 and n29275 n29276_not ; n29277
g29214 and a[11] n29277_not ; n29278
g29215 and a[11] n29278_not ; n29279
g29216 nor n29277 n29278 ; n29280
g29217 nor n29279 n29280 ; n29281
g29218 and n29270 n29281_not ; n29282
g29219 and n29270 n29282_not ; n29283
g29220 nor n29281 n29282 ; n29284
g29221 nor n29283 n29284 ; n29285
g29222 nor n29051 n29064 ; n29286
g29223 and n29285 n29286 ; n29287
g29224 nor n29285 n29286 ; n29288
g29225 nor n29287 n29288 ; n29289
g29226 nor n29070 n29083 ; n29290
g29227 and n9331 n27964 ; n29291
g29228 and n8418 n27442 ; n29292
g29229 and n8860 n27698 ; n29293
g29230 nor n29292 n29293 ; n29294
g29231 and n29291_not n29294 ; n29295
g29232 and n8421 n27976 ; n29296
g29233 and n29295 n29296_not ; n29297
g29234 and a[8] n29297_not ; n29298
g29235 and a[8] n29298_not ; n29299
g29236 nor n29297 n29298 ; n29300
g29237 nor n29299 n29300 ; n29301
g29238 nor n29290 n29301 ; n29302
g29239 nor n29290 n29302 ; n29303
g29240 nor n29301 n29302 ; n29304
g29241 nor n29303 n29304 ; n29305
g29242 and n29289_not n29305 ; n29306
g29243 and n29289 n29305_not ; n29307
g29244 nor n29306 n29307 ; n29308
g29245 and n29116_not n29308 ; n29309
g29246 and n29116 n29308_not ; n29310
g29247 nor n29309 n29310 ; n29311
g29248 and n29115_not n29311 ; n29312
g29249 and n29115 n29311_not ; n29313
g29250 nor n29312 n29313 ; n29314
g29251 nor n29112 n29314 ; n29315
g29252 and n29112 n29314 ; n29316
g29253 nor n29315 n29316 ; result[10]
g29254 nor n29159 n29172 ; n29318
g29255 and n75 n23345_not ; n29319
g29256 and n3020 n22356 ; n29320
g29257 and n3023 n22362 ; n29321
g29258 and n3028 n22359 ; n29322
g29259 nor n29321 n29322 ; n29323
g29260 and n29320_not n29323 ; n29324
g29261 and n29319_not n29324 ; n29325
g29262 and n1324 n6056 ; n29326
g29263 and n1206 n29326 ; n29327
g29264 and n1346 n29327 ; n29328
g29265 and n6705 n29328 ; n29329
g29266 and n654 n29329 ; n29330
g29267 and n3470 n29330 ; n29331
g29268 and n869 n29331 ; n29332
g29269 and n1141 n29332 ; n29333
g29270 and n229_not n29333 ; n29334
g29271 and n121_not n29334 ; n29335
g29272 and n248_not n29335 ; n29336
g29273 and n206_not n29336 ; n29337
g29274 and n1732 n2263 ; n29338
g29275 and n3160 n29338 ; n29339
g29276 and n6771 n29339 ; n29340
g29277 and n29337 n29340 ; n29341
g29278 and n1378 n29341 ; n29342
g29279 and n2678 n29342 ; n29343
g29280 and n600 n29343 ; n29344
g29281 and n488 n29344 ; n29345
g29282 and n1009 n29345 ; n29346
g29283 and n1825 n29346 ; n29347
g29284 and n1522 n29347 ; n29348
g29285 and n1011_not n29348 ; n29349
g29286 and n1246_not n29349 ; n29350
g29287 and n275_not n29350 ; n29351
g29288 and n357_not n29351 ; n29352
g29289 and n165_not n29352 ; n29353
g29290 and n493_not n29353 ; n29354
g29291 and n655_not n29354 ; n29355
g29292 and n28496 n29132_not ; n29356
g29293 nor n29140 n29356 ; n29357
g29294 and n29355 n29357_not ; n29358
g29295 and n29355_not n29357 ; n29359
g29296 nor n29358 n29359 ; n29360
g29297 and n29325_not n29360 ; n29361
g29298 nor n29325 n29361 ; n29362
g29299 and n29360 n29361_not ; n29363
g29300 nor n29362 n29363 ; n29364
g29301 nor n28925 n29144 ; n29365
g29302 nor n29155 n29365 ; n29366
g29303 and n29364 n29366 ; n29367
g29304 nor n29364 n29366 ; n29368
g29305 nor n29367 n29368 ; n29369
g29306 and n3457 n22347 ; n29370
g29307 and n3542 n22353 ; n29371
g29308 and n3606 n22350 ; n29372
g29309 nor n29371 n29372 ; n29373
g29310 and n29370_not n29373 ; n29374
g29311 and n3368_not n29374 ; n29375
g29312 and n23659 n29374 ; n29376
g29313 nor n29375 n29376 ; n29377
g29314 and a[29] n29377_not ; n29378
g29315 and a[29]_not n29377 ; n29379
g29316 nor n29378 n29379 ; n29380
g29317 and n29369 n29380_not ; n29381
g29318 and n29369_not n29380 ; n29382
g29319 nor n29381 n29382 ; n29383
g29320 and n29318_not n29383 ; n29384
g29321 and n29318 n29383_not ; n29385
g29322 nor n29384 n29385 ; n29386
g29323 and n3884 n22338 ; n29387
g29324 and n3967 n22344 ; n29388
g29325 and n4046 n22341 ; n29389
g29326 nor n29388 n29389 ; n29390
g29327 and n29387_not n29390 ; n29391
g29328 and n4050 n24188_not ; n29392
g29329 and n29391 n29392_not ; n29393
g29330 and a[26] n29393_not ; n29394
g29331 and a[26] n29394_not ; n29395
g29332 nor n29393 n29394 ; n29396
g29333 nor n29395 n29396 ; n29397
g29334 and n29386 n29397_not ; n29398
g29335 and n29386 n29398_not ; n29399
g29336 nor n29397 n29398 ; n29400
g29337 nor n29399 n29400 ; n29401
g29338 nor n29187 n29193 ; n29402
g29339 and n29401 n29402 ; n29403
g29340 nor n29401 n29402 ; n29404
g29341 nor n29403 n29404 ; n29405
g29342 and n4694 n22329 ; n29406
g29343 and n4533 n22335 ; n29407
g29344 and n4604 n22332 ; n29408
g29345 nor n29407 n29408 ; n29409
g29346 and n29406_not n29409 ; n29410
g29347 and n4536 n24633_not ; n29411
g29348 and n29410 n29411_not ; n29412
g29349 and a[23] n29412_not ; n29413
g29350 and a[23] n29413_not ; n29414
g29351 nor n29412 n29413 ; n29415
g29352 nor n29414 n29415 ; n29416
g29353 and n29405 n29416_not ; n29417
g29354 and n29405 n29417_not ; n29418
g29355 nor n29416 n29417 ; n29419
g29356 nor n29418 n29419 ; n29420
g29357 nor n29206 n29212 ; n29421
g29358 and n29420 n29421 ; n29422
g29359 nor n29420 n29421 ; n29423
g29360 nor n29422 n29423 ; n29424
g29361 and n5496 n22320 ; n29425
g29362 and n4935 n22326 ; n29426
g29363 and n5407 n22323 ; n29427
g29364 nor n29426 n29427 ; n29428
g29365 and n29425_not n29428 ; n29429
g29366 and n4938 n25270_not ; n29430
g29367 and n29429 n29430_not ; n29431
g29368 and a[20] n29431_not ; n29432
g29369 and a[20] n29432_not ; n29433
g29370 nor n29431 n29432 ; n29434
g29371 nor n29433 n29434 ; n29435
g29372 and n29424 n29435_not ; n29436
g29373 and n29424 n29436_not ; n29437
g29374 nor n29435 n29436 ; n29438
g29375 nor n29437 n29438 ; n29439
g29376 nor n29225 n29231 ; n29440
g29377 and n29439 n29440 ; n29441
g29378 nor n29439 n29440 ; n29442
g29379 nor n29441 n29442 ; n29443
g29380 and n6233 n22309 ; n29444
g29381 and n5663 n22312 ; n29445
g29382 and n5939 n22315 ; n29446
g29383 nor n29445 n29446 ; n29447
g29384 and n29444_not n29447 ; n29448
g29385 and n5666 n22529_not ; n29449
g29386 and n29448 n29449_not ; n29450
g29387 and a[17] n29450_not ; n29451
g29388 and a[17] n29451_not ; n29452
g29389 nor n29450 n29451 ; n29453
g29390 nor n29452 n29453 ; n29454
g29391 and n29443 n29454_not ; n29455
g29392 and n29443 n29455_not ; n29456
g29393 nor n29454 n29455 ; n29457
g29394 nor n29456 n29457 ; n29458
g29395 nor n29244 n29250 ; n29459
g29396 and n29458 n29459 ; n29460
g29397 nor n29458 n29459 ; n29461
g29398 nor n29460 n29461 ; n29462
g29399 and n7101 n26060 ; n29463
g29400 and n6402 n26063 ; n29464
g29401 and n6951 n26066 ; n29465
g29402 nor n29464 n29465 ; n29466
g29403 and n29463_not n29466 ; n29467
g29404 and n6397 n26088_not ; n29468
g29405 and n29467 n29468_not ; n29469
g29406 and a[14] n29469_not ; n29470
g29407 and a[14] n29470_not ; n29471
g29408 nor n29469 n29470 ; n29472
g29409 nor n29471 n29472 ; n29473
g29410 and n29462 n29473_not ; n29474
g29411 and n29462 n29474_not ; n29475
g29412 nor n29473 n29474 ; n29476
g29413 nor n29475 n29476 ; n29477
g29414 nor n29264 n29269 ; n29478
g29415 nor n29477 n29478 ; n29479
g29416 nor n29477 n29479 ; n29480
g29417 nor n29478 n29479 ; n29481
g29418 nor n29480 n29481 ; n29482
g29419 and n7983 n27442 ; n29483
g29420 and n7291 n26890 ; n29484
g29421 and n7632 n27173 ; n29485
g29422 nor n29484 n29485 ; n29486
g29423 and n29483_not n29486 ; n29487
g29424 and n7294 n27455 ; n29488
g29425 and n29487 n29488_not ; n29489
g29426 and a[11] n29489_not ; n29490
g29427 and a[11] n29490_not ; n29491
g29428 nor n29489 n29490 ; n29492
g29429 nor n29491 n29492 ; n29493
g29430 nor n29482 n29493 ; n29494
g29431 nor n29482 n29494 ; n29495
g29432 nor n29493 n29494 ; n29496
g29433 nor n29495 n29496 ; n29497
g29434 nor n29282 n29288 ; n29498
g29435 and n29497 n29498 ; n29499
g29436 nor n29497 n29498 ; n29500
g29437 nor n29499 n29500 ; n29501
g29438 and n9331 n28208_not ; n29502
g29439 and n8418 n27698 ; n29503
g29440 and n8860 n27964 ; n29504
g29441 nor n29503 n29504 ; n29505
g29442 and n29502_not n29505 ; n29506
g29443 and n8421 n28223_not ; n29507
g29444 and n29506 n29507_not ; n29508
g29445 and a[8] n29508_not ; n29509
g29446 and a[8] n29509_not ; n29510
g29447 nor n29508 n29509 ; n29511
g29448 nor n29510 n29511 ; n29512
g29449 and n29501 n29512_not ; n29513
g29450 and n29501 n29513_not ; n29514
g29451 nor n29512 n29513 ; n29515
g29452 nor n29514 n29515 ; n29516
g29453 nor n29302 n29307 ; n29517
g29454 nor n29516 n29517 ; n29518
g29455 nor n29516 n29518 ; n29519
g29456 nor n29517 n29518 ; n29520
g29457 nor n29519 n29520 ; n29521
g29458 nor n29309 n29312 ; n29522
g29459 and n29521 n29522 ; n29523
g29460 nor n29521 n29522 ; n29524
g29461 nor n29523 n29524 ; n29525
g29462 and n29316_not n29525 ; n29526
g29463 and n29316 n29525_not ; n29527
g29464 or n29526 n29527 ; result[11]
g29465 and n29316 n29525 ; n29529
g29466 nor n29358 n29361 ; n29530
g29467 nor n175 n255 ; n29531
g29468 and n299_not n29531 ; n29532
g29469 and n305_not n29532 ; n29533
g29470 and n492_not n29533 ; n29534
g29471 and n165_not n29534 ; n29535
g29472 and n592_not n29535 ; n29536
g29473 and n672_not n29536 ; n29537
g29474 and n270_not n29537 ; n29538
g29475 and n2442 n12712 ; n29539
g29476 and n940 n29539 ; n29540
g29477 and n4295 n29540 ; n29541
g29478 and n2406 n29541 ; n29542
g29479 and n1046 n29542 ; n29543
g29480 and n2417 n29543 ; n29544
g29481 and n885 n29544 ; n29545
g29482 and n289_not n29545 ; n29546
g29483 and n155_not n29546 ; n29547
g29484 and n164_not n29547 ; n29548
g29485 and n191_not n29548 ; n29549
g29486 and n245_not n29549 ; n29550
g29487 and n12911 n13808 ; n29551
g29488 and n6548 n29551 ; n29552
g29489 and n29550 n29552 ; n29553
g29490 and n29538 n29553 ; n29554
g29491 and n3065 n29554 ; n29555
g29492 and n12396 n29555 ; n29556
g29493 and n194_not n29556 ; n29557
g29494 and n254_not n29557 ; n29558
g29495 and n435_not n29558 ; n29559
g29496 and n243_not n29559 ; n29560
g29497 and n466_not n29560 ; n29561
g29498 and n537_not n29561 ; n29562
g29499 and n332_not n29562 ; n29563
g29500 and n325_not n29563 ; n29564
g29501 and n29355_not n29564 ; n29565
g29502 and n29355 n29564_not ; n29566
g29503 nor n29530 n29566 ; n29567
g29504 and n29565_not n29567 ; n29568
g29505 nor n29530 n29568 ; n29569
g29506 nor n29566 n29568 ; n29570
g29507 and n29565_not n29570 ; n29571
g29508 nor n29569 n29571 ; n29572
g29509 and n75 n22556_not ; n29573
g29510 and n3020 n22353 ; n29574
g29511 and n3023 n22359 ; n29575
g29512 and n3028 n22356 ; n29576
g29513 nor n29575 n29576 ; n29577
g29514 and n29574_not n29577 ; n29578
g29515 and n29573_not n29578 ; n29579
g29516 nor n29572 n29579 ; n29580
g29517 nor n29572 n29580 ; n29581
g29518 nor n29579 n29580 ; n29582
g29519 nor n29581 n29582 ; n29583
g29520 nor n29368 n29381 ; n29584
g29521 and n29583 n29584 ; n29585
g29522 nor n29583 n29584 ; n29586
g29523 nor n29585 n29586 ; n29587
g29524 and n3457 n22344 ; n29588
g29525 and n3542 n22350 ; n29589
g29526 and n3606 n22347 ; n29590
g29527 nor n29589 n29590 ; n29591
g29528 and n29588_not n29591 ; n29592
g29529 and n3368 n23642_not ; n29593
g29530 and n29592 n29593_not ; n29594
g29531 and a[29] n29594_not ; n29595
g29532 and a[29] n29595_not ; n29596
g29533 nor n29594 n29595 ; n29597
g29534 nor n29596 n29597 ; n29598
g29535 and n29587 n29598_not ; n29599
g29536 and n29587 n29599_not ; n29600
g29537 nor n29598 n29599 ; n29601
g29538 nor n29600 n29601 ; n29602
g29539 and n3884 n22335 ; n29603
g29540 and n3967 n22341 ; n29604
g29541 and n4046 n22338 ; n29605
g29542 nor n29604 n29605 ; n29606
g29543 and n29603_not n29606 ; n29607
g29544 and n4050 n24167_not ; n29608
g29545 and n29607 n29608_not ; n29609
g29546 and a[26] n29609_not ; n29610
g29547 and a[26] n29610_not ; n29611
g29548 nor n29609 n29610 ; n29612
g29549 nor n29611 n29612 ; n29613
g29550 nor n29602 n29613 ; n29614
g29551 nor n29602 n29614 ; n29615
g29552 nor n29613 n29614 ; n29616
g29553 nor n29615 n29616 ; n29617
g29554 nor n29384 n29398 ; n29618
g29555 and n29617 n29618 ; n29619
g29556 nor n29617 n29618 ; n29620
g29557 nor n29619 n29620 ; n29621
g29558 and n4694 n22326 ; n29622
g29559 and n4533 n22332 ; n29623
g29560 and n4604 n22329 ; n29624
g29561 nor n29623 n29624 ; n29625
g29562 and n29622_not n29625 ; n29626
g29563 and n4536 n24616_not ; n29627
g29564 and n29626 n29627_not ; n29628
g29565 and a[23] n29628_not ; n29629
g29566 and a[23] n29629_not ; n29630
g29567 nor n29628 n29629 ; n29631
g29568 nor n29630 n29631 ; n29632
g29569 and n29621 n29632_not ; n29633
g29570 and n29621 n29633_not ; n29634
g29571 nor n29632 n29633 ; n29635
g29572 nor n29634 n29635 ; n29636
g29573 nor n29404 n29417 ; n29637
g29574 and n29636 n29637 ; n29638
g29575 nor n29636 n29637 ; n29639
g29576 nor n29638 n29639 ; n29640
g29577 and n5496 n22312 ; n29641
g29578 and n4935 n22323 ; n29642
g29579 and n5407 n22320 ; n29643
g29580 nor n29642 n29643 ; n29644
g29581 and n29641_not n29644 ; n29645
g29582 and n4938 n25315_not ; n29646
g29583 and n29645 n29646_not ; n29647
g29584 and a[20] n29647_not ; n29648
g29585 and a[20] n29648_not ; n29649
g29586 nor n29647 n29648 ; n29650
g29587 nor n29649 n29650 ; n29651
g29588 and n29640 n29651_not ; n29652
g29589 and n29640 n29652_not ; n29653
g29590 nor n29651 n29652 ; n29654
g29591 nor n29653 n29654 ; n29655
g29592 nor n29423 n29436 ; n29656
g29593 and n29655 n29656 ; n29657
g29594 nor n29655 n29656 ; n29658
g29595 nor n29657 n29658 ; n29659
g29596 and n6233 n26063 ; n29660
g29597 and n5663 n22315 ; n29661
g29598 and n5939 n22309 ; n29662
g29599 nor n29661 n29662 ; n29663
g29600 and n29660_not n29663 ; n29664
g29601 and n5666 n26604_not ; n29665
g29602 and n29664 n29665_not ; n29666
g29603 and a[17] n29666_not ; n29667
g29604 and a[17] n29667_not ; n29668
g29605 nor n29666 n29667 ; n29669
g29606 nor n29668 n29669 ; n29670
g29607 and n29659 n29670_not ; n29671
g29608 and n29659 n29671_not ; n29672
g29609 nor n29670 n29671 ; n29673
g29610 nor n29672 n29673 ; n29674
g29611 nor n29442 n29455 ; n29675
g29612 and n29674 n29675 ; n29676
g29613 nor n29674 n29675 ; n29677
g29614 nor n29676 n29677 ; n29678
g29615 and n7101 n26890 ; n29679
g29616 and n6402 n26066 ; n29680
g29617 and n6951 n26060 ; n29681
g29618 nor n29680 n29681 ; n29682
g29619 and n29679_not n29682 ; n29683
g29620 and n6397 n26904_not ; n29684
g29621 and n29683 n29684_not ; n29685
g29622 and a[14] n29685_not ; n29686
g29623 and a[14] n29686_not ; n29687
g29624 nor n29685 n29686 ; n29688
g29625 nor n29687 n29688 ; n29689
g29626 and n29678 n29689_not ; n29690
g29627 and n29678 n29690_not ; n29691
g29628 nor n29689 n29690 ; n29692
g29629 nor n29691 n29692 ; n29693
g29630 nor n29461 n29474 ; n29694
g29631 and n29693 n29694 ; n29695
g29632 nor n29693 n29694 ; n29696
g29633 nor n29695 n29696 ; n29697
g29634 and n7983 n27698 ; n29698
g29635 and n7291 n27173 ; n29699
g29636 and n7632 n27442 ; n29700
g29637 nor n29699 n29700 ; n29701
g29638 and n29698_not n29701 ; n29702
g29639 and n7294 n27713_not ; n29703
g29640 and n29702 n29703_not ; n29704
g29641 and a[11] n29704_not ; n29705
g29642 and a[11] n29705_not ; n29706
g29643 nor n29704 n29705 ; n29707
g29644 nor n29706 n29707 ; n29708
g29645 and n29697 n29708_not ; n29709
g29646 and n29697 n29709_not ; n29710
g29647 nor n29708 n29709 ; n29711
g29648 nor n29710 n29711 ; n29712
g29649 nor n29479 n29494 ; n29713
g29650 nor n14590 n28208 ; n29714
g29651 and n8418 n27964 ; n29715
g29652 nor n29714 n29715 ; n29716
g29653 and n8421_not n29716 ; n29717
g29654 and n28221 n29716 ; n29718
g29655 nor n29717 n29718 ; n29719
g29656 and a[8] n29719_not ; n29720
g29657 and a[8]_not n29719 ; n29721
g29658 nor n29720 n29721 ; n29722
g29659 nor n29713 n29722 ; n29723
g29660 and n29713 n29722 ; n29724
g29661 nor n29723 n29724 ; n29725
g29662 and n29712_not n29725 ; n29726
g29663 nor n29712 n29726 ; n29727
g29664 and n29725 n29726_not ; n29728
g29665 nor n29727 n29728 ; n29729
g29666 nor n29500 n29513 ; n29730
g29667 and n29729 n29730 ; n29731
g29668 nor n29729 n29730 ; n29732
g29669 nor n29731 n29732 ; n29733
g29670 nor n29518 n29524 ; n29734
g29671 and n29733_not n29734 ; n29735
g29672 and n29733 n29734_not ; n29736
g29673 nor n29735 n29736 ; n29737
g29674 and n29529 n29737 ; n29738
g29675 nor n29529 n29737 ; n29739
g29676 nor n29738 n29739 ; result[12]
g29677 nor n29732 n29736 ; n29741
g29678 nor n29723 n29726 ; n29742
g29679 and n75 n23672 ; n29743
g29680 and n3020 n22350 ; n29744
g29681 and n3023 n22356 ; n29745
g29682 and n3028 n22353 ; n29746
g29683 nor n29745 n29746 ; n29747
g29684 and n29744_not n29747 ; n29748
g29685 and n29743_not n29748 ; n29749
g29686 nor n14592 n28208 ; n29750
g29687 and a[8] n29750_not ; n29751
g29688 and a[8]_not n29750 ; n29752
g29689 nor n29751 n29752 ; n29753
g29690 and n960 n3474 ; n29754
g29691 and n1422 n29754 ; n29755
g29692 and n300 n29755 ; n29756
g29693 and n13773 n29756 ; n29757
g29694 and n2006 n29757 ; n29758
g29695 and n1575 n29758 ; n29759
g29696 and n2697 n29759 ; n29760
g29697 and n235 n29760 ; n29761
g29698 and n2958 n29761 ; n29762
g29699 and n2484 n29762 ; n29763
g29700 and n2170 n29763 ; n29764
g29701 and n156 n29764 ; n29765
g29702 and n713_not n29765 ; n29766
g29703 and n368_not n29766 ; n29767
g29704 and n29355 n29767 ; n29768
g29705 nor n29355 n29767 ; n29769
g29706 nor n29768 n29769 ; n29770
g29707 and n29753 n29770 ; n29771
g29708 nor n29753 n29770 ; n29772
g29709 nor n29771 n29772 ; n29773
g29710 and n29570_not n29773 ; n29774
g29711 and n29570 n29773_not ; n29775
g29712 nor n29774 n29775 ; n29776
g29713 and n29749_not n29776 ; n29777
g29714 and n29776 n29777_not ; n29778
g29715 nor n29749 n29777 ; n29779
g29716 nor n29778 n29779 ; n29780
g29717 and n3457 n22341 ; n29781
g29718 and n3542 n22347 ; n29782
g29719 and n3606 n22344 ; n29783
g29720 nor n29782 n29783 ; n29784
g29721 and n29781_not n29784 ; n29785
g29722 and n3368 n24142 ; n29786
g29723 and n29785 n29786_not ; n29787
g29724 and a[29] n29787_not ; n29788
g29725 and a[29] n29788_not ; n29789
g29726 nor n29787 n29788 ; n29790
g29727 nor n29789 n29790 ; n29791
g29728 nor n29780 n29791 ; n29792
g29729 nor n29780 n29792 ; n29793
g29730 nor n29791 n29792 ; n29794
g29731 nor n29793 n29794 ; n29795
g29732 nor n29580 n29586 ; n29796
g29733 and n29795 n29796 ; n29797
g29734 nor n29795 n29796 ; n29798
g29735 nor n29797 n29798 ; n29799
g29736 and n3884 n22332 ; n29800
g29737 and n3967 n22338 ; n29801
g29738 and n4046 n22335 ; n29802
g29739 nor n29801 n29802 ; n29803
g29740 and n29800_not n29803 ; n29804
g29741 and n4050 n22542 ; n29805
g29742 and n29804 n29805_not ; n29806
g29743 and a[26] n29806_not ; n29807
g29744 and a[26] n29807_not ; n29808
g29745 nor n29806 n29807 ; n29809
g29746 nor n29808 n29809 ; n29810
g29747 and n29799 n29810_not ; n29811
g29748 and n29799 n29811_not ; n29812
g29749 nor n29810 n29811 ; n29813
g29750 nor n29812 n29813 ; n29814
g29751 nor n29599 n29614 ; n29815
g29752 and n29814 n29815 ; n29816
g29753 nor n29814 n29815 ; n29817
g29754 nor n29816 n29817 ; n29818
g29755 and n4694 n22323 ; n29819
g29756 and n4533 n22329 ; n29820
g29757 and n4604 n22326 ; n29821
g29758 nor n29820 n29821 ; n29822
g29759 and n29819_not n29822 ; n29823
g29760 and n4536 n24599 ; n29824
g29761 and n29823 n29824_not ; n29825
g29762 and a[23] n29825_not ; n29826
g29763 and a[23] n29826_not ; n29827
g29764 nor n29825 n29826 ; n29828
g29765 nor n29827 n29828 ; n29829
g29766 and n29818 n29829_not ; n29830
g29767 and n29818 n29830_not ; n29831
g29768 nor n29829 n29830 ; n29832
g29769 nor n29831 n29832 ; n29833
g29770 nor n29620 n29633 ; n29834
g29771 and n29833 n29834 ; n29835
g29772 nor n29833 n29834 ; n29836
g29773 nor n29835 n29836 ; n29837
g29774 and n5496 n22315 ; n29838
g29775 and n4935 n22320 ; n29839
g29776 and n5407 n22312 ; n29840
g29777 nor n29839 n29840 ; n29841
g29778 and n29838_not n29841 ; n29842
g29779 and n4938 n25294 ; n29843
g29780 and n29842 n29843_not ; n29844
g29781 and a[20] n29844_not ; n29845
g29782 and a[20] n29845_not ; n29846
g29783 nor n29844 n29845 ; n29847
g29784 nor n29846 n29847 ; n29848
g29785 and n29837 n29848_not ; n29849
g29786 and n29837 n29849_not ; n29850
g29787 nor n29848 n29849 ; n29851
g29788 nor n29850 n29851 ; n29852
g29789 nor n29639 n29652 ; n29853
g29790 and n29852 n29853 ; n29854
g29791 nor n29852 n29853 ; n29855
g29792 nor n29854 n29855 ; n29856
g29793 nor n29658 n29671 ; n29857
g29794 and n6233 n26066 ; n29858
g29795 and n5663 n22309 ; n29859
g29796 and n5939 n26063 ; n29860
g29797 nor n29859 n29860 ; n29861
g29798 and n29858_not n29861 ; n29862
g29799 and n5666 n26624_not ; n29863
g29800 and n29862 n29863_not ; n29864
g29801 and a[17] n29864_not ; n29865
g29802 and a[17] n29865_not ; n29866
g29803 nor n29864 n29865 ; n29867
g29804 nor n29866 n29867 ; n29868
g29805 nor n29857 n29868 ; n29869
g29806 nor n29857 n29869 ; n29870
g29807 nor n29868 n29869 ; n29871
g29808 nor n29870 n29871 ; n29872
g29809 and n29856_not n29872 ; n29873
g29810 and n29856 n29872_not ; n29874
g29811 nor n29873 n29874 ; n29875
g29812 and n7101 n27173 ; n29876
g29813 and n6402 n26060 ; n29877
g29814 and n6951 n26890 ; n29878
g29815 nor n29877 n29878 ; n29879
g29816 and n29876_not n29879 ; n29880
g29817 and n6397 n27185 ; n29881
g29818 and n29880 n29881_not ; n29882
g29819 and a[14] n29882_not ; n29883
g29820 and a[14] n29883_not ; n29884
g29821 nor n29882 n29883 ; n29885
g29822 nor n29884 n29885 ; n29886
g29823 and n29875 n29886_not ; n29887
g29824 and n29875 n29887_not ; n29888
g29825 nor n29886 n29887 ; n29889
g29826 nor n29888 n29889 ; n29890
g29827 nor n29677 n29690 ; n29891
g29828 and n29890 n29891 ; n29892
g29829 nor n29890 n29891 ; n29893
g29830 nor n29892 n29893 ; n29894
g29831 nor n29696 n29709 ; n29895
g29832 and n7983 n27964 ; n29896
g29833 and n7291 n27442 ; n29897
g29834 and n7632 n27698 ; n29898
g29835 nor n29897 n29898 ; n29899
g29836 and n29896_not n29899 ; n29900
g29837 and n7294 n27976 ; n29901
g29838 and n29900 n29901_not ; n29902
g29839 and a[11] n29902_not ; n29903
g29840 and a[11] n29903_not ; n29904
g29841 nor n29902 n29903 ; n29905
g29842 nor n29904 n29905 ; n29906
g29843 nor n29895 n29906 ; n29907
g29844 nor n29895 n29907 ; n29908
g29845 nor n29906 n29907 ; n29909
g29846 nor n29908 n29909 ; n29910
g29847 and n29894_not n29910 ; n29911
g29848 and n29894 n29910_not ; n29912
g29849 nor n29911 n29912 ; n29913
g29850 and n29742_not n29913 ; n29914
g29851 and n29742 n29913_not ; n29915
g29852 nor n29914 n29915 ; n29916
g29853 and n29741_not n29916 ; n29917
g29854 and n29741 n29916_not ; n29918
g29855 nor n29917 n29918 ; n29919
g29856 nor n29738 n29919 ; n29920
g29857 and n29738 n29919 ; n29921
g29858 nor n29920 n29921 ; result[13]
g29859 nor n29792 n29798 ; n29923
g29860 and n75 n23659_not ; n29924
g29861 and n3020 n22347 ; n29925
g29862 and n3023 n22353 ; n29926
g29863 and n3028 n22350 ; n29927
g29864 nor n29926 n29927 ; n29928
g29865 and n29925_not n29928 ; n29929
g29866 and n29924_not n29929 ; n29930
g29867 nor n29769 n29771 ; n29931
g29868 and n962 n1490 ; n29932
g29869 and n15854 n29932 ; n29933
g29870 and n14407 n29933 ; n29934
g29871 and n4767 n29934 ; n29935
g29872 and n4786 n29935 ; n29936
g29873 and n1719 n29936 ; n29937
g29874 and n3559 n29937 ; n29938
g29875 and n2635 n29938 ; n29939
g29876 and n242_not n29939 ; n29940
g29877 and n150_not n29940 ; n29941
g29878 and n357_not n29941 ; n29942
g29879 and n286_not n29942 ; n29943
g29880 and n980_not n29943 ; n29944
g29881 and n1010_not n29944 ; n29945
g29882 and n270_not n29945 ; n29946
g29883 and n29931_not n29946 ; n29947
g29884 and n29931 n29946_not ; n29948
g29885 nor n29947 n29948 ; n29949
g29886 and n29930_not n29949 ; n29950
g29887 nor n29930 n29950 ; n29951
g29888 and n29949 n29950_not ; n29952
g29889 nor n29951 n29952 ; n29953
g29890 nor n29774 n29777 ; n29954
g29891 and n29953 n29954 ; n29955
g29892 nor n29953 n29954 ; n29956
g29893 nor n29955 n29956 ; n29957
g29894 and n3457 n22338 ; n29958
g29895 and n3542 n22344 ; n29959
g29896 and n3606 n22341 ; n29960
g29897 nor n29959 n29960 ; n29961
g29898 and n29958_not n29961 ; n29962
g29899 and n3368_not n29962 ; n29963
g29900 and n24188 n29962 ; n29964
g29901 nor n29963 n29964 ; n29965
g29902 and a[29] n29965_not ; n29966
g29903 and a[29]_not n29965 ; n29967
g29904 nor n29966 n29967 ; n29968
g29905 and n29957 n29968_not ; n29969
g29906 and n29957_not n29968 ; n29970
g29907 nor n29969 n29970 ; n29971
g29908 and n29923_not n29971 ; n29972
g29909 and n29923 n29971_not ; n29973
g29910 nor n29972 n29973 ; n29974
g29911 and n3884 n22329 ; n29975
g29912 and n3967 n22335 ; n29976
g29913 and n4046 n22332 ; n29977
g29914 nor n29976 n29977 ; n29978
g29915 and n29975_not n29978 ; n29979
g29916 and n4050 n24633_not ; n29980
g29917 and n29979 n29980_not ; n29981
g29918 and a[26] n29981_not ; n29982
g29919 and a[26] n29982_not ; n29983
g29920 nor n29981 n29982 ; n29984
g29921 nor n29983 n29984 ; n29985
g29922 and n29974 n29985_not ; n29986
g29923 and n29974 n29986_not ; n29987
g29924 nor n29985 n29986 ; n29988
g29925 nor n29987 n29988 ; n29989
g29926 nor n29811 n29817 ; n29990
g29927 and n29989 n29990 ; n29991
g29928 nor n29989 n29990 ; n29992
g29929 nor n29991 n29992 ; n29993
g29930 and n4694 n22320 ; n29994
g29931 and n4533 n22326 ; n29995
g29932 and n4604 n22323 ; n29996
g29933 nor n29995 n29996 ; n29997
g29934 and n29994_not n29997 ; n29998
g29935 and n4536 n25270_not ; n29999
g29936 and n29998 n29999_not ; n30000
g29937 and a[23] n30000_not ; n30001
g29938 and a[23] n30001_not ; n30002
g29939 nor n30000 n30001 ; n30003
g29940 nor n30002 n30003 ; n30004
g29941 and n29993 n30004_not ; n30005
g29942 and n29993 n30005_not ; n30006
g29943 nor n30004 n30005 ; n30007
g29944 nor n30006 n30007 ; n30008
g29945 nor n29830 n29836 ; n30009
g29946 and n30008 n30009 ; n30010
g29947 nor n30008 n30009 ; n30011
g29948 nor n30010 n30011 ; n30012
g29949 and n5496 n22309 ; n30013
g29950 and n4935 n22312 ; n30014
g29951 and n5407 n22315 ; n30015
g29952 nor n30014 n30015 ; n30016
g29953 and n30013_not n30016 ; n30017
g29954 and n4938 n22529_not ; n30018
g29955 and n30017 n30018_not ; n30019
g29956 and a[20] n30019_not ; n30020
g29957 and a[20] n30020_not ; n30021
g29958 nor n30019 n30020 ; n30022
g29959 nor n30021 n30022 ; n30023
g29960 and n30012 n30023_not ; n30024
g29961 and n30012 n30024_not ; n30025
g29962 nor n30023 n30024 ; n30026
g29963 nor n30025 n30026 ; n30027
g29964 nor n29849 n29855 ; n30028
g29965 and n30027 n30028 ; n30029
g29966 nor n30027 n30028 ; n30030
g29967 nor n30029 n30030 ; n30031
g29968 and n6233 n26060 ; n30032
g29969 and n5663 n26063 ; n30033
g29970 and n5939 n26066 ; n30034
g29971 nor n30033 n30034 ; n30035
g29972 and n30032_not n30035 ; n30036
g29973 and n5666 n26088_not ; n30037
g29974 and n30036 n30037_not ; n30038
g29975 and a[17] n30038_not ; n30039
g29976 and a[17] n30039_not ; n30040
g29977 nor n30038 n30039 ; n30041
g29978 nor n30040 n30041 ; n30042
g29979 and n30031 n30042_not ; n30043
g29980 and n30031 n30043_not ; n30044
g29981 nor n30042 n30043 ; n30045
g29982 nor n30044 n30045 ; n30046
g29983 nor n29869 n29874 ; n30047
g29984 nor n30046 n30047 ; n30048
g29985 nor n30046 n30048 ; n30049
g29986 nor n30047 n30048 ; n30050
g29987 nor n30049 n30050 ; n30051
g29988 and n7101 n27442 ; n30052
g29989 and n6402 n26890 ; n30053
g29990 and n6951 n27173 ; n30054
g29991 nor n30053 n30054 ; n30055
g29992 and n30052_not n30055 ; n30056
g29993 and n6397 n27455 ; n30057
g29994 and n30056 n30057_not ; n30058
g29995 and a[14] n30058_not ; n30059
g29996 and a[14] n30059_not ; n30060
g29997 nor n30058 n30059 ; n30061
g29998 nor n30060 n30061 ; n30062
g29999 nor n30051 n30062 ; n30063
g30000 nor n30051 n30063 ; n30064
g30001 nor n30062 n30063 ; n30065
g30002 nor n30064 n30065 ; n30066
g30003 nor n29887 n29893 ; n30067
g30004 and n30066 n30067 ; n30068
g30005 nor n30066 n30067 ; n30069
g30006 nor n30068 n30069 ; n30070
g30007 and n7983 n28208_not ; n30071
g30008 and n7291 n27698 ; n30072
g30009 and n7632 n27964 ; n30073
g30010 nor n30072 n30073 ; n30074
g30011 and n30071_not n30074 ; n30075
g30012 and n7294 n28223_not ; n30076
g30013 and n30075 n30076_not ; n30077
g30014 and a[11] n30077_not ; n30078
g30015 and a[11] n30078_not ; n30079
g30016 nor n30077 n30078 ; n30080
g30017 nor n30079 n30080 ; n30081
g30018 and n30070 n30081_not ; n30082
g30019 and n30070 n30082_not ; n30083
g30020 nor n30081 n30082 ; n30084
g30021 nor n30083 n30084 ; n30085
g30022 nor n29907 n29912 ; n30086
g30023 nor n30085 n30086 ; n30087
g30024 nor n30085 n30087 ; n30088
g30025 nor n30086 n30087 ; n30089
g30026 nor n30088 n30089 ; n30090
g30027 nor n29914 n29917 ; n30091
g30028 and n30090 n30091 ; n30092
g30029 nor n30090 n30091 ; n30093
g30030 nor n30092 n30093 ; n30094
g30031 and n29921 n30094_not ; n30095
g30032 and n29921_not n30094 ; n30096
g30033 or n30095 n30096 ; result[14]
g30034 nor n29956 n29969 ; n30098
g30035 nor n29947 n29950 ; n30099
g30036 and n2705 n2811 ; n30100
g30037 and n2007 n30100 ; n30101
g30038 and n1012 n30101 ; n30102
g30039 and n877 n30102 ; n30103
g30040 and n13768 n30103 ; n30104
g30041 and n15312 n30104 ; n30105
g30042 and n5286 n30105 ; n30106
g30043 and n2651 n30106 ; n30107
g30044 and n291 n30107 ; n30108
g30045 and n1330 n30108 ; n30109
g30046 and n29337 n30109 ; n30110
g30047 and n731 n30110 ; n30111
g30048 and n1247 n30111 ; n30112
g30049 and n426_not n30112 ; n30113
g30050 and n292_not n30113 ; n30114
g30051 and n102_not n30114 ; n30115
g30052 and n422_not n30115 ; n30116
g30053 and n531_not n30116 ; n30117
g30054 and n29946_not n30117 ; n30118
g30055 and n29946 n30117_not ; n30119
g30056 nor n30099 n30119 ; n30120
g30057 and n30118_not n30120 ; n30121
g30058 nor n30099 n30121 ; n30122
g30059 nor n30119 n30121 ; n30123
g30060 and n30118_not n30123 ; n30124
g30061 nor n30122 n30124 ; n30125
g30062 and n75 n23642_not ; n30126
g30063 and n3020 n22344 ; n30127
g30064 and n3023 n22350 ; n30128
g30065 and n3028 n22347 ; n30129
g30066 nor n30128 n30129 ; n30130
g30067 and n30127_not n30130 ; n30131
g30068 and n30126_not n30131 ; n30132
g30069 nor n30125 n30132 ; n30133
g30070 nor n30125 n30133 ; n30134
g30071 nor n30132 n30133 ; n30135
g30072 nor n30134 n30135 ; n30136
g30073 and n3457 n22335 ; n30137
g30074 and n3542 n22341 ; n30138
g30075 and n3606 n22338 ; n30139
g30076 nor n30138 n30139 ; n30140
g30077 and n30137_not n30140 ; n30141
g30078 and n3368_not n30141 ; n30142
g30079 and n24167 n30141 ; n30143
g30080 nor n30142 n30143 ; n30144
g30081 and a[29] n30144_not ; n30145
g30082 and a[29]_not n30144 ; n30146
g30083 nor n30145 n30146 ; n30147
g30084 nor n30136 n30147 ; n30148
g30085 and n30136 n30147 ; n30149
g30086 nor n30148 n30149 ; n30150
g30087 and n30098_not n30150 ; n30151
g30088 and n30098 n30150_not ; n30152
g30089 nor n30151 n30152 ; n30153
g30090 and n3884 n22326 ; n30154
g30091 and n3967 n22332 ; n30155
g30092 and n4046 n22329 ; n30156
g30093 nor n30155 n30156 ; n30157
g30094 and n30154_not n30157 ; n30158
g30095 and n4050 n24616_not ; n30159
g30096 and n30158 n30159_not ; n30160
g30097 and a[26] n30160_not ; n30161
g30098 and a[26] n30161_not ; n30162
g30099 nor n30160 n30161 ; n30163
g30100 nor n30162 n30163 ; n30164
g30101 and n30153 n30164_not ; n30165
g30102 and n30153 n30165_not ; n30166
g30103 nor n30164 n30165 ; n30167
g30104 nor n30166 n30167 ; n30168
g30105 nor n29972 n29986 ; n30169
g30106 and n30168 n30169 ; n30170
g30107 nor n30168 n30169 ; n30171
g30108 nor n30170 n30171 ; n30172
g30109 and n4694 n22312 ; n30173
g30110 and n4533 n22323 ; n30174
g30111 and n4604 n22320 ; n30175
g30112 nor n30174 n30175 ; n30176
g30113 and n30173_not n30176 ; n30177
g30114 and n4536 n25315_not ; n30178
g30115 and n30177 n30178_not ; n30179
g30116 and a[23] n30179_not ; n30180
g30117 and a[23] n30180_not ; n30181
g30118 nor n30179 n30180 ; n30182
g30119 nor n30181 n30182 ; n30183
g30120 and n30172 n30183_not ; n30184
g30121 and n30172 n30184_not ; n30185
g30122 nor n30183 n30184 ; n30186
g30123 nor n30185 n30186 ; n30187
g30124 nor n29992 n30005 ; n30188
g30125 and n30187 n30188 ; n30189
g30126 nor n30187 n30188 ; n30190
g30127 nor n30189 n30190 ; n30191
g30128 and n5496 n26063 ; n30192
g30129 and n4935 n22315 ; n30193
g30130 and n5407 n22309 ; n30194
g30131 nor n30193 n30194 ; n30195
g30132 and n30192_not n30195 ; n30196
g30133 and n4938 n26604_not ; n30197
g30134 and n30196 n30197_not ; n30198
g30135 and a[20] n30198_not ; n30199
g30136 and a[20] n30199_not ; n30200
g30137 nor n30198 n30199 ; n30201
g30138 nor n30200 n30201 ; n30202
g30139 and n30191 n30202_not ; n30203
g30140 and n30191 n30203_not ; n30204
g30141 nor n30202 n30203 ; n30205
g30142 nor n30204 n30205 ; n30206
g30143 nor n30011 n30024 ; n30207
g30144 and n30206 n30207 ; n30208
g30145 nor n30206 n30207 ; n30209
g30146 nor n30208 n30209 ; n30210
g30147 and n6233 n26890 ; n30211
g30148 and n5663 n26066 ; n30212
g30149 and n5939 n26060 ; n30213
g30150 nor n30212 n30213 ; n30214
g30151 and n30211_not n30214 ; n30215
g30152 and n5666 n26904_not ; n30216
g30153 and n30215 n30216_not ; n30217
g30154 and a[17] n30217_not ; n30218
g30155 and a[17] n30218_not ; n30219
g30156 nor n30217 n30218 ; n30220
g30157 nor n30219 n30220 ; n30221
g30158 and n30210 n30221_not ; n30222
g30159 and n30210 n30222_not ; n30223
g30160 nor n30221 n30222 ; n30224
g30161 nor n30223 n30224 ; n30225
g30162 nor n30030 n30043 ; n30226
g30163 and n30225 n30226 ; n30227
g30164 nor n30225 n30226 ; n30228
g30165 nor n30227 n30228 ; n30229
g30166 and n7101 n27698 ; n30230
g30167 and n6402 n27173 ; n30231
g30168 and n6951 n27442 ; n30232
g30169 nor n30231 n30232 ; n30233
g30170 and n30230_not n30233 ; n30234
g30171 and n6397 n27713_not ; n30235
g30172 and n30234 n30235_not ; n30236
g30173 and a[14] n30236_not ; n30237
g30174 and a[14] n30237_not ; n30238
g30175 nor n30236 n30237 ; n30239
g30176 nor n30238 n30239 ; n30240
g30177 and n30229 n30240_not ; n30241
g30178 and n30229 n30241_not ; n30242
g30179 nor n30240 n30241 ; n30243
g30180 nor n30242 n30243 ; n30244
g30181 nor n30048 n30063 ; n30245
g30182 nor n14424 n28208 ; n30246
g30183 and n7291 n27964 ; n30247
g30184 nor n30246 n30247 ; n30248
g30185 and n7294_not n30248 ; n30249
g30186 and n28221 n30248 ; n30250
g30187 nor n30249 n30250 ; n30251
g30188 and a[11] n30251_not ; n30252
g30189 and a[11]_not n30251 ; n30253
g30190 nor n30252 n30253 ; n30254
g30191 nor n30245 n30254 ; n30255
g30192 and n30245 n30254 ; n30256
g30193 nor n30255 n30256 ; n30257
g30194 and n30244_not n30257 ; n30258
g30195 nor n30244 n30258 ; n30259
g30196 and n30257 n30258_not ; n30260
g30197 nor n30259 n30260 ; n30261
g30198 nor n30069 n30082 ; n30262
g30199 and n30261 n30262 ; n30263
g30200 nor n30261 n30262 ; n30264
g30201 nor n30263 n30264 ; n30265
g30202 nor n30087 n30093 ; n30266
g30203 and n30265_not n30266 ; n30267
g30204 and n30265 n30266_not ; n30268
g30205 nor n30267 n30268 ; n30269
g30206 and n29921 n30094 ; n30270
g30207 and n30269 n30270 ; n30271
g30208 nor n30269 n30270 ; n30272
g30209 nor n30271 n30272 ; result[15]
g30210 nor n30264 n30268 ; n30274
g30211 nor n30255 n30258 ; n30275
g30212 nor n30133 n30148 ; n30276
g30213 and n75 n24142 ; n30277
g30214 and n3020 n22341 ; n30278
g30215 and n3023 n22347 ; n30279
g30216 and n3028 n22344 ; n30280
g30217 nor n30279 n30280 ; n30281
g30218 and n30278_not n30281 ; n30282
g30219 and n30277_not n30282 ; n30283
g30220 nor n14426 n28208 ; n30284
g30221 and a[11] n30284_not ; n30285
g30222 and a[11]_not n30284 ; n30286
g30223 nor n30285 n30286 ; n30287
g30224 and n675 n2174 ; n30288
g30225 and n5038 n30288 ; n30289
g30226 and n2808 n30289 ; n30290
g30227 and n5019 n30290 ; n30291
g30228 and n1407 n30291 ; n30292
g30229 and n3510 n30292 ; n30293
g30230 and n241 n30293 ; n30294
g30231 and n1435 n30294 ; n30295
g30232 and n1576 n30295 ; n30296
g30233 and n1252 n30296 ; n30297
g30234 and n3886 n30297 ; n30298
g30235 and n590 n30298 ; n30299
g30236 and n242_not n30299 ; n30300
g30237 and n435_not n30300 ; n30301
g30238 and n532_not n30301 ; n30302
g30239 and n363_not n30302 ; n30303
g30240 and n29946 n30303 ; n30304
g30241 nor n29946 n30303 ; n30305
g30242 nor n30304 n30305 ; n30306
g30243 and n30287 n30306 ; n30307
g30244 nor n30287 n30306 ; n30308
g30245 nor n30307 n30308 ; n30309
g30246 and n30283_not n30309 ; n30310
g30247 and n30309 n30310_not ; n30311
g30248 nor n30283 n30310 ; n30312
g30249 nor n30311 n30312 ; n30313
g30250 nor n30123 n30313 ; n30314
g30251 nor n30313 n30314 ; n30315
g30252 nor n30123 n30314 ; n30316
g30253 nor n30315 n30316 ; n30317
g30254 nor n30276 n30317 ; n30318
g30255 nor n30276 n30318 ; n30319
g30256 nor n30317 n30318 ; n30320
g30257 nor n30319 n30320 ; n30321
g30258 and n3457 n22332 ; n30322
g30259 and n3542 n22338 ; n30323
g30260 and n3606 n22335 ; n30324
g30261 nor n30323 n30324 ; n30325
g30262 and n30322_not n30325 ; n30326
g30263 and n3368 n22542 ; n30327
g30264 and n30326 n30327_not ; n30328
g30265 and a[29] n30328_not ; n30329
g30266 and a[29] n30329_not ; n30330
g30267 nor n30328 n30329 ; n30331
g30268 nor n30330 n30331 ; n30332
g30269 nor n30321 n30332 ; n30333
g30270 nor n30321 n30333 ; n30334
g30271 nor n30332 n30333 ; n30335
g30272 nor n30334 n30335 ; n30336
g30273 and n3884 n22323 ; n30337
g30274 and n3967 n22329 ; n30338
g30275 and n4046 n22326 ; n30339
g30276 nor n30338 n30339 ; n30340
g30277 and n30337_not n30340 ; n30341
g30278 and n4050 n24599 ; n30342
g30279 and n30341 n30342_not ; n30343
g30280 and a[26] n30343_not ; n30344
g30281 and a[26] n30344_not ; n30345
g30282 nor n30343 n30344 ; n30346
g30283 nor n30345 n30346 ; n30347
g30284 nor n30336 n30347 ; n30348
g30285 nor n30336 n30348 ; n30349
g30286 nor n30347 n30348 ; n30350
g30287 nor n30349 n30350 ; n30351
g30288 nor n30151 n30165 ; n30352
g30289 and n30351 n30352 ; n30353
g30290 nor n30351 n30352 ; n30354
g30291 nor n30353 n30354 ; n30355
g30292 and n4694 n22315 ; n30356
g30293 and n4533 n22320 ; n30357
g30294 and n4604 n22312 ; n30358
g30295 nor n30357 n30358 ; n30359
g30296 and n30356_not n30359 ; n30360
g30297 and n4536 n25294 ; n30361
g30298 and n30360 n30361_not ; n30362
g30299 and a[23] n30362_not ; n30363
g30300 and a[23] n30363_not ; n30364
g30301 nor n30362 n30363 ; n30365
g30302 nor n30364 n30365 ; n30366
g30303 and n30355 n30366_not ; n30367
g30304 and n30355 n30367_not ; n30368
g30305 nor n30366 n30367 ; n30369
g30306 nor n30368 n30369 ; n30370
g30307 nor n30171 n30184 ; n30371
g30308 and n30370 n30371 ; n30372
g30309 nor n30370 n30371 ; n30373
g30310 nor n30372 n30373 ; n30374
g30311 nor n30190 n30203 ; n30375
g30312 and n5496 n26066 ; n30376
g30313 and n4935 n22309 ; n30377
g30314 and n5407 n26063 ; n30378
g30315 nor n30377 n30378 ; n30379
g30316 and n30376_not n30379 ; n30380
g30317 and n4938 n26624_not ; n30381
g30318 and n30380 n30381_not ; n30382
g30319 and a[20] n30382_not ; n30383
g30320 and a[20] n30383_not ; n30384
g30321 nor n30382 n30383 ; n30385
g30322 nor n30384 n30385 ; n30386
g30323 nor n30375 n30386 ; n30387
g30324 nor n30375 n30387 ; n30388
g30325 nor n30386 n30387 ; n30389
g30326 nor n30388 n30389 ; n30390
g30327 and n30374_not n30390 ; n30391
g30328 and n30374 n30390_not ; n30392
g30329 nor n30391 n30392 ; n30393
g30330 and n6233 n27173 ; n30394
g30331 and n5663 n26060 ; n30395
g30332 and n5939 n26890 ; n30396
g30333 nor n30395 n30396 ; n30397
g30334 and n30394_not n30397 ; n30398
g30335 and n5666 n27185 ; n30399
g30336 and n30398 n30399_not ; n30400
g30337 and a[17] n30400_not ; n30401
g30338 and a[17] n30401_not ; n30402
g30339 nor n30400 n30401 ; n30403
g30340 nor n30402 n30403 ; n30404
g30341 and n30393 n30404_not ; n30405
g30342 and n30393 n30405_not ; n30406
g30343 nor n30404 n30405 ; n30407
g30344 nor n30406 n30407 ; n30408
g30345 nor n30209 n30222 ; n30409
g30346 and n30408 n30409 ; n30410
g30347 nor n30408 n30409 ; n30411
g30348 nor n30410 n30411 ; n30412
g30349 nor n30228 n30241 ; n30413
g30350 and n7101 n27964 ; n30414
g30351 and n6402 n27442 ; n30415
g30352 and n6951 n27698 ; n30416
g30353 nor n30415 n30416 ; n30417
g30354 and n30414_not n30417 ; n30418
g30355 and n6397 n27976 ; n30419
g30356 and n30418 n30419_not ; n30420
g30357 and a[14] n30420_not ; n30421
g30358 and a[14] n30421_not ; n30422
g30359 nor n30420 n30421 ; n30423
g30360 nor n30422 n30423 ; n30424
g30361 nor n30413 n30424 ; n30425
g30362 nor n30413 n30425 ; n30426
g30363 nor n30424 n30425 ; n30427
g30364 nor n30426 n30427 ; n30428
g30365 and n30412_not n30428 ; n30429
g30366 and n30412 n30428_not ; n30430
g30367 nor n30429 n30430 ; n30431
g30368 and n30275_not n30431 ; n30432
g30369 and n30275 n30431_not ; n30433
g30370 nor n30432 n30433 ; n30434
g30371 and n30274_not n30434 ; n30435
g30372 and n30274 n30434_not ; n30436
g30373 nor n30435 n30436 ; n30437
g30374 nor n30271 n30437 ; n30438
g30375 and n30271 n30437 ; n30439
g30376 nor n30438 n30439 ; result[16]
g30377 nor n30318 n30333 ; n30441
g30378 and n75 n24188_not ; n30442
g30379 and n3020 n22338 ; n30443
g30380 and n3023 n22344 ; n30444
g30381 and n3028 n22341 ; n30445
g30382 nor n30444 n30445 ; n30446
g30383 and n30443_not n30446 ; n30447
g30384 and n30442_not n30447 ; n30448
g30385 nor n30305 n30307 ; n30449
g30386 and n1499 n2059 ; n30450
g30387 and n778 n30450 ; n30451
g30388 and n3128 n30451 ; n30452
g30389 and n12977 n30452 ; n30453
g30390 and n27789 n30453 ; n30454
g30391 and n13458 n30454 ; n30455
g30392 and n15324 n30455 ; n30456
g30393 and n28294 n30456 ; n30457
g30394 and n1380 n30457 ; n30458
g30395 and n810 n30458 ; n30459
g30396 and n469_not n30459 ; n30460
g30397 and n746_not n30460 ; n30461
g30398 and n1102_not n30461 ; n30462
g30399 and n396_not n30462 ; n30463
g30400 and n470_not n30463 ; n30464
g30401 and n30449_not n30464 ; n30465
g30402 and n30449 n30464_not ; n30466
g30403 nor n30465 n30466 ; n30467
g30404 and n30448_not n30467 ; n30468
g30405 nor n30448 n30468 ; n30469
g30406 and n30467 n30468_not ; n30470
g30407 nor n30469 n30470 ; n30471
g30408 nor n30310 n30314 ; n30472
g30409 and n30471 n30472 ; n30473
g30410 nor n30471 n30472 ; n30474
g30411 nor n30473 n30474 ; n30475
g30412 and n3457 n22329 ; n30476
g30413 and n3542 n22335 ; n30477
g30414 and n3606 n22332 ; n30478
g30415 nor n30477 n30478 ; n30479
g30416 and n30476_not n30479 ; n30480
g30417 and n3368_not n30480 ; n30481
g30418 and n24633 n30480 ; n30482
g30419 nor n30481 n30482 ; n30483
g30420 and a[29] n30483_not ; n30484
g30421 and a[29]_not n30483 ; n30485
g30422 nor n30484 n30485 ; n30486
g30423 and n30475 n30486_not ; n30487
g30424 and n30475_not n30486 ; n30488
g30425 nor n30487 n30488 ; n30489
g30426 and n30441_not n30489 ; n30490
g30427 and n30441 n30489_not ; n30491
g30428 nor n30490 n30491 ; n30492
g30429 and n3884 n22320 ; n30493
g30430 and n3967 n22326 ; n30494
g30431 and n4046 n22323 ; n30495
g30432 nor n30494 n30495 ; n30496
g30433 and n30493_not n30496 ; n30497
g30434 and n4050 n25270_not ; n30498
g30435 and n30497 n30498_not ; n30499
g30436 and a[26] n30499_not ; n30500
g30437 and a[26] n30500_not ; n30501
g30438 nor n30499 n30500 ; n30502
g30439 nor n30501 n30502 ; n30503
g30440 and n30492 n30503_not ; n30504
g30441 and n30492 n30504_not ; n30505
g30442 nor n30503 n30504 ; n30506
g30443 nor n30505 n30506 ; n30507
g30444 nor n30348 n30354 ; n30508
g30445 and n30507 n30508 ; n30509
g30446 nor n30507 n30508 ; n30510
g30447 nor n30509 n30510 ; n30511
g30448 and n4694 n22309 ; n30512
g30449 and n4533 n22312 ; n30513
g30450 and n4604 n22315 ; n30514
g30451 nor n30513 n30514 ; n30515
g30452 and n30512_not n30515 ; n30516
g30453 and n4536 n22529_not ; n30517
g30454 and n30516 n30517_not ; n30518
g30455 and a[23] n30518_not ; n30519
g30456 and a[23] n30519_not ; n30520
g30457 nor n30518 n30519 ; n30521
g30458 nor n30520 n30521 ; n30522
g30459 and n30511 n30522_not ; n30523
g30460 and n30511 n30523_not ; n30524
g30461 nor n30522 n30523 ; n30525
g30462 nor n30524 n30525 ; n30526
g30463 nor n30367 n30373 ; n30527
g30464 and n30526 n30527 ; n30528
g30465 nor n30526 n30527 ; n30529
g30466 nor n30528 n30529 ; n30530
g30467 and n5496 n26060 ; n30531
g30468 and n4935 n26063 ; n30532
g30469 and n5407 n26066 ; n30533
g30470 nor n30532 n30533 ; n30534
g30471 and n30531_not n30534 ; n30535
g30472 and n4938 n26088_not ; n30536
g30473 and n30535 n30536_not ; n30537
g30474 and a[20] n30537_not ; n30538
g30475 and a[20] n30538_not ; n30539
g30476 nor n30537 n30538 ; n30540
g30477 nor n30539 n30540 ; n30541
g30478 and n30530 n30541_not ; n30542
g30479 and n30530 n30542_not ; n30543
g30480 nor n30541 n30542 ; n30544
g30481 nor n30543 n30544 ; n30545
g30482 nor n30387 n30392 ; n30546
g30483 nor n30545 n30546 ; n30547
g30484 nor n30545 n30547 ; n30548
g30485 nor n30546 n30547 ; n30549
g30486 nor n30548 n30549 ; n30550
g30487 and n6233 n27442 ; n30551
g30488 and n5663 n26890 ; n30552
g30489 and n5939 n27173 ; n30553
g30490 nor n30552 n30553 ; n30554
g30491 and n30551_not n30554 ; n30555
g30492 and n5666 n27455 ; n30556
g30493 and n30555 n30556_not ; n30557
g30494 and a[17] n30557_not ; n30558
g30495 and a[17] n30558_not ; n30559
g30496 nor n30557 n30558 ; n30560
g30497 nor n30559 n30560 ; n30561
g30498 nor n30550 n30561 ; n30562
g30499 nor n30550 n30562 ; n30563
g30500 nor n30561 n30562 ; n30564
g30501 nor n30563 n30564 ; n30565
g30502 nor n30405 n30411 ; n30566
g30503 and n30565 n30566 ; n30567
g30504 nor n30565 n30566 ; n30568
g30505 nor n30567 n30568 ; n30569
g30506 and n7101 n28208_not ; n30570
g30507 and n6402 n27698 ; n30571
g30508 and n6951 n27964 ; n30572
g30509 nor n30571 n30572 ; n30573
g30510 and n30570_not n30573 ; n30574
g30511 and n6397 n28223_not ; n30575
g30512 and n30574 n30575_not ; n30576
g30513 and a[14] n30576_not ; n30577
g30514 and a[14] n30577_not ; n30578
g30515 nor n30576 n30577 ; n30579
g30516 nor n30578 n30579 ; n30580
g30517 and n30569 n30580_not ; n30581
g30518 and n30569 n30581_not ; n30582
g30519 nor n30580 n30581 ; n30583
g30520 nor n30582 n30583 ; n30584
g30521 nor n30425 n30430 ; n30585
g30522 nor n30584 n30585 ; n30586
g30523 nor n30584 n30586 ; n30587
g30524 nor n30585 n30586 ; n30588
g30525 nor n30587 n30588 ; n30589
g30526 nor n30432 n30435 ; n30590
g30527 and n30589 n30590 ; n30591
g30528 nor n30589 n30590 ; n30592
g30529 nor n30591 n30592 ; n30593
g30530 and n30439_not n30593 ; n30594
g30531 and n30439 n30593_not ; n30595
g30532 or n30594 n30595 ; result[17]
g30533 and n30439 n30593 ; n30597
g30534 and n75 n24167_not ; n30598
g30535 and n3020 n22335 ; n30599
g30536 and n3023 n22341 ; n30600
g30537 and n3028 n22338 ; n30601
g30538 nor n30600 n30601 ; n30602
g30539 and n30599_not n30602 ; n30603
g30540 and n30598_not n30603 ; n30604
g30541 and n694 n2176 ; n30605
g30542 and n6084 n30605 ; n30606
g30543 and n3108 n30606 ; n30607
g30544 and n12710 n30607 ; n30608
g30545 and n13123 n30608 ; n30609
g30546 and n3386 n30609 ; n30610
g30547 and n2500 n30610 ; n30611
g30548 and n5209 n30611 ; n30612
g30549 and n2739 n30612 ; n30613
g30550 and n558_not n30613 ; n30614
g30551 and n1102_not n30614 ; n30615
g30552 and n155_not n30615 ; n30616
g30553 and n248_not n30616 ; n30617
g30554 and n357_not n30617 ; n30618
g30555 and n205_not n30618 ; n30619
g30556 and n436_not n30619 ; n30620
g30557 and n81_not n30620 ; n30621
g30558 and n30464_not n30621 ; n30622
g30559 and n30464 n30621_not ; n30623
g30560 nor n30604 n30623 ; n30624
g30561 and n30622_not n30624 ; n30625
g30562 nor n30604 n30625 ; n30626
g30563 nor n30623 n30625 ; n30627
g30564 and n30622_not n30627 ; n30628
g30565 nor n30626 n30628 ; n30629
g30566 nor n30465 n30468 ; n30630
g30567 and n30629 n30630 ; n30631
g30568 nor n30629 n30630 ; n30632
g30569 nor n30631 n30632 ; n30633
g30570 nor n30474 n30487 ; n30634
g30571 and n30633_not n30634 ; n30635
g30572 and n30633 n30634_not ; n30636
g30573 nor n30635 n30636 ; n30637
g30574 and n3457 n22326 ; n30638
g30575 and n3542 n22332 ; n30639
g30576 and n3606 n22329 ; n30640
g30577 nor n30639 n30640 ; n30641
g30578 and n30638_not n30641 ; n30642
g30579 and n3368 n24616_not ; n30643
g30580 and n30642 n30643_not ; n30644
g30581 and a[29] n30644_not ; n30645
g30582 and a[29] n30645_not ; n30646
g30583 nor n30644 n30645 ; n30647
g30584 nor n30646 n30647 ; n30648
g30585 and n30637 n30648_not ; n30649
g30586 and n30637 n30649_not ; n30650
g30587 nor n30648 n30649 ; n30651
g30588 nor n30650 n30651 ; n30652
g30589 and n3884 n22312 ; n30653
g30590 and n3967 n22323 ; n30654
g30591 and n4046 n22320 ; n30655
g30592 nor n30654 n30655 ; n30656
g30593 and n30653_not n30656 ; n30657
g30594 and n4050 n25315_not ; n30658
g30595 and n30657 n30658_not ; n30659
g30596 and a[26] n30659_not ; n30660
g30597 and a[26] n30660_not ; n30661
g30598 nor n30659 n30660 ; n30662
g30599 nor n30661 n30662 ; n30663
g30600 nor n30652 n30663 ; n30664
g30601 nor n30652 n30664 ; n30665
g30602 nor n30663 n30664 ; n30666
g30603 nor n30665 n30666 ; n30667
g30604 nor n30490 n30504 ; n30668
g30605 and n30667 n30668 ; n30669
g30606 nor n30667 n30668 ; n30670
g30607 nor n30669 n30670 ; n30671
g30608 and n4694 n26063 ; n30672
g30609 and n4533 n22315 ; n30673
g30610 and n4604 n22309 ; n30674
g30611 nor n30673 n30674 ; n30675
g30612 and n30672_not n30675 ; n30676
g30613 and n4536 n26604_not ; n30677
g30614 and n30676 n30677_not ; n30678
g30615 and a[23] n30678_not ; n30679
g30616 and a[23] n30679_not ; n30680
g30617 nor n30678 n30679 ; n30681
g30618 nor n30680 n30681 ; n30682
g30619 and n30671 n30682_not ; n30683
g30620 and n30671 n30683_not ; n30684
g30621 nor n30682 n30683 ; n30685
g30622 nor n30684 n30685 ; n30686
g30623 nor n30510 n30523 ; n30687
g30624 and n30686 n30687 ; n30688
g30625 nor n30686 n30687 ; n30689
g30626 nor n30688 n30689 ; n30690
g30627 and n5496 n26890 ; n30691
g30628 and n4935 n26066 ; n30692
g30629 and n5407 n26060 ; n30693
g30630 nor n30692 n30693 ; n30694
g30631 and n30691_not n30694 ; n30695
g30632 and n4938 n26904_not ; n30696
g30633 and n30695 n30696_not ; n30697
g30634 and a[20] n30697_not ; n30698
g30635 and a[20] n30698_not ; n30699
g30636 nor n30697 n30698 ; n30700
g30637 nor n30699 n30700 ; n30701
g30638 and n30690 n30701_not ; n30702
g30639 and n30690 n30702_not ; n30703
g30640 nor n30701 n30702 ; n30704
g30641 nor n30703 n30704 ; n30705
g30642 nor n30529 n30542 ; n30706
g30643 and n30705 n30706 ; n30707
g30644 nor n30705 n30706 ; n30708
g30645 nor n30707 n30708 ; n30709
g30646 and n6233 n27698 ; n30710
g30647 and n5663 n27173 ; n30711
g30648 and n5939 n27442 ; n30712
g30649 nor n30711 n30712 ; n30713
g30650 and n30710_not n30713 ; n30714
g30651 and n5666 n27713_not ; n30715
g30652 and n30714 n30715_not ; n30716
g30653 and a[17] n30716_not ; n30717
g30654 and a[17] n30717_not ; n30718
g30655 nor n30716 n30717 ; n30719
g30656 nor n30718 n30719 ; n30720
g30657 and n30709 n30720_not ; n30721
g30658 and n30709 n30721_not ; n30722
g30659 nor n30720 n30721 ; n30723
g30660 nor n30722 n30723 ; n30724
g30661 nor n30547 n30562 ; n30725
g30662 nor n13845 n28208 ; n30726
g30663 and n6402 n27964 ; n30727
g30664 nor n30726 n30727 ; n30728
g30665 and n6397_not n30728 ; n30729
g30666 and n28221 n30728 ; n30730
g30667 nor n30729 n30730 ; n30731
g30668 and a[14] n30731_not ; n30732
g30669 and a[14]_not n30731 ; n30733
g30670 nor n30732 n30733 ; n30734
g30671 nor n30725 n30734 ; n30735
g30672 and n30725 n30734 ; n30736
g30673 nor n30735 n30736 ; n30737
g30674 and n30724_not n30737 ; n30738
g30675 nor n30724 n30738 ; n30739
g30676 and n30737 n30738_not ; n30740
g30677 nor n30739 n30740 ; n30741
g30678 nor n30568 n30581 ; n30742
g30679 and n30741 n30742 ; n30743
g30680 nor n30741 n30742 ; n30744
g30681 nor n30743 n30744 ; n30745
g30682 nor n30586 n30592 ; n30746
g30683 and n30745_not n30746 ; n30747
g30684 and n30745 n30746_not ; n30748
g30685 nor n30747 n30748 ; n30749
g30686 and n30597 n30749 ; n30750
g30687 nor n30597 n30749 ; n30751
g30688 nor n30750 n30751 ; result[18]
g30689 nor n30744 n30748 ; n30753
g30690 nor n30735 n30738 ; n30754
g30691 and n75 n22542 ; n30755
g30692 and n3020 n22332 ; n30756
g30693 and n3023 n22338 ; n30757
g30694 and n3028 n22335 ; n30758
g30695 nor n30757 n30758 ; n30759
g30696 and n30756_not n30759 ; n30760
g30697 and n30755_not n30760 ; n30761
g30698 nor n13847 n28208 ; n30762
g30699 and a[14] n30762_not ; n30763
g30700 and a[14]_not n30762 ; n30764
g30701 nor n30763 n30764 ; n30765
g30702 and n2537 n3045 ; n30766
g30703 and n14482 n30766 ; n30767
g30704 and n1894 n30767 ; n30768
g30705 and n14202 n30768 ; n30769
g30706 and n6714 n30769 ; n30770
g30707 and n1291 n30770 ; n30771
g30708 and n976 n30771 ; n30772
g30709 and n1139 n30772 ; n30773
g30710 and n2219 n30773 ; n30774
g30711 and n357_not n30774 ; n30775
g30712 and n326_not n30775 ; n30776
g30713 and n452_not n30776 ; n30777
g30714 and n30464 n30777 ; n30778
g30715 nor n30464 n30777 ; n30779
g30716 nor n30778 n30779 ; n30780
g30717 and n30765 n30780 ; n30781
g30718 nor n30765 n30780 ; n30782
g30719 nor n30781 n30782 ; n30783
g30720 and n30627_not n30783 ; n30784
g30721 and n30627 n30783_not ; n30785
g30722 nor n30784 n30785 ; n30786
g30723 and n30761_not n30786 ; n30787
g30724 and n30786 n30787_not ; n30788
g30725 nor n30761 n30787 ; n30789
g30726 nor n30788 n30789 ; n30790
g30727 and n3457 n22323 ; n30791
g30728 and n3542 n22329 ; n30792
g30729 and n3606 n22326 ; n30793
g30730 nor n30792 n30793 ; n30794
g30731 and n30791_not n30794 ; n30795
g30732 and n3368 n24599 ; n30796
g30733 and n30795 n30796_not ; n30797
g30734 and a[29] n30797_not ; n30798
g30735 and a[29] n30798_not ; n30799
g30736 nor n30797 n30798 ; n30800
g30737 nor n30799 n30800 ; n30801
g30738 nor n30790 n30801 ; n30802
g30739 nor n30790 n30802 ; n30803
g30740 nor n30801 n30802 ; n30804
g30741 nor n30803 n30804 ; n30805
g30742 nor n30632 n30636 ; n30806
g30743 and n30805 n30806 ; n30807
g30744 nor n30805 n30806 ; n30808
g30745 nor n30807 n30808 ; n30809
g30746 and n3884 n22315 ; n30810
g30747 and n3967 n22320 ; n30811
g30748 and n4046 n22312 ; n30812
g30749 nor n30811 n30812 ; n30813
g30750 and n30810_not n30813 ; n30814
g30751 and n4050 n25294 ; n30815
g30752 and n30814 n30815_not ; n30816
g30753 and a[26] n30816_not ; n30817
g30754 and a[26] n30817_not ; n30818
g30755 nor n30816 n30817 ; n30819
g30756 nor n30818 n30819 ; n30820
g30757 and n30809 n30820_not ; n30821
g30758 and n30809 n30821_not ; n30822
g30759 nor n30820 n30821 ; n30823
g30760 nor n30822 n30823 ; n30824
g30761 nor n30649 n30664 ; n30825
g30762 and n30824 n30825 ; n30826
g30763 nor n30824 n30825 ; n30827
g30764 nor n30826 n30827 ; n30828
g30765 nor n30670 n30683 ; n30829
g30766 and n4694 n26066 ; n30830
g30767 and n4533 n22309 ; n30831
g30768 and n4604 n26063 ; n30832
g30769 nor n30831 n30832 ; n30833
g30770 and n30830_not n30833 ; n30834
g30771 and n4536 n26624_not ; n30835
g30772 and n30834 n30835_not ; n30836
g30773 and a[23] n30836_not ; n30837
g30774 and a[23] n30837_not ; n30838
g30775 nor n30836 n30837 ; n30839
g30776 nor n30838 n30839 ; n30840
g30777 nor n30829 n30840 ; n30841
g30778 nor n30829 n30841 ; n30842
g30779 nor n30840 n30841 ; n30843
g30780 nor n30842 n30843 ; n30844
g30781 and n30828_not n30844 ; n30845
g30782 and n30828 n30844_not ; n30846
g30783 nor n30845 n30846 ; n30847
g30784 and n5496 n27173 ; n30848
g30785 and n4935 n26060 ; n30849
g30786 and n5407 n26890 ; n30850
g30787 nor n30849 n30850 ; n30851
g30788 and n30848_not n30851 ; n30852
g30789 and n4938 n27185 ; n30853
g30790 and n30852 n30853_not ; n30854
g30791 and a[20] n30854_not ; n30855
g30792 and a[20] n30855_not ; n30856
g30793 nor n30854 n30855 ; n30857
g30794 nor n30856 n30857 ; n30858
g30795 and n30847 n30858_not ; n30859
g30796 and n30847 n30859_not ; n30860
g30797 nor n30858 n30859 ; n30861
g30798 nor n30860 n30861 ; n30862
g30799 nor n30689 n30702 ; n30863
g30800 and n30862 n30863 ; n30864
g30801 nor n30862 n30863 ; n30865
g30802 nor n30864 n30865 ; n30866
g30803 nor n30708 n30721 ; n30867
g30804 and n6233 n27964 ; n30868
g30805 and n5663 n27442 ; n30869
g30806 and n5939 n27698 ; n30870
g30807 nor n30869 n30870 ; n30871
g30808 and n30868_not n30871 ; n30872
g30809 and n5666 n27976 ; n30873
g30810 and n30872 n30873_not ; n30874
g30811 and a[17] n30874_not ; n30875
g30812 and a[17] n30875_not ; n30876
g30813 nor n30874 n30875 ; n30877
g30814 nor n30876 n30877 ; n30878
g30815 nor n30867 n30878 ; n30879
g30816 nor n30867 n30879 ; n30880
g30817 nor n30878 n30879 ; n30881
g30818 nor n30880 n30881 ; n30882
g30819 and n30866_not n30882 ; n30883
g30820 and n30866 n30882_not ; n30884
g30821 nor n30883 n30884 ; n30885
g30822 and n30754_not n30885 ; n30886
g30823 and n30754 n30885_not ; n30887
g30824 nor n30886 n30887 ; n30888
g30825 and n30753_not n30888 ; n30889
g30826 and n30753 n30888_not ; n30890
g30827 nor n30889 n30890 ; n30891
g30828 nor n30750 n30891 ; n30892
g30829 and n30750 n30891 ; n30893
g30830 nor n30892 n30893 ; result[19]
g30831 nor n30802 n30808 ; n30895
g30832 and n75 n24633_not ; n30896
g30833 and n3020 n22329 ; n30897
g30834 and n3023 n22335 ; n30898
g30835 and n3028 n22332 ; n30899
g30836 nor n30898 n30899 ; n30900
g30837 and n30897_not n30900 ; n30901
g30838 and n30896_not n30901 ; n30902
g30839 nor n30779 n30781 ; n30903
g30840 and n1369 n3393 ; n30904
g30841 and n2361 n30904 ; n30905
g30842 and n14525 n30905 ; n30906
g30843 and n5034 n30906 ; n30907
g30844 and n5773 n30907 ; n30908
g30845 and n977 n30908 ; n30909
g30846 and n491 n30909 ; n30910
g30847 and n1183 n30910 ; n30911
g30848 and n2346 n30911 ; n30912
g30849 and n2697 n30912 ; n30913
g30850 and n471 n30913 ; n30914
g30851 and n1782 n30914 ; n30915
g30852 and n224_not n30915 ; n30916
g30853 and n146_not n30916 ; n30917
g30854 and n161_not n30917 ; n30918
g30855 and n358_not n30918 ; n30919
g30856 and n30903_not n30919 ; n30920
g30857 and n30903 n30919_not ; n30921
g30858 nor n30920 n30921 ; n30922
g30859 and n30902_not n30922 ; n30923
g30860 nor n30902 n30923 ; n30924
g30861 and n30922 n30923_not ; n30925
g30862 nor n30924 n30925 ; n30926
g30863 nor n30784 n30787 ; n30927
g30864 and n30926 n30927 ; n30928
g30865 nor n30926 n30927 ; n30929
g30866 nor n30928 n30929 ; n30930
g30867 and n3457 n22320 ; n30931
g30868 and n3542 n22326 ; n30932
g30869 and n3606 n22323 ; n30933
g30870 nor n30932 n30933 ; n30934
g30871 and n30931_not n30934 ; n30935
g30872 and n3368_not n30935 ; n30936
g30873 and n25270 n30935 ; n30937
g30874 nor n30936 n30937 ; n30938
g30875 and a[29] n30938_not ; n30939
g30876 and a[29]_not n30938 ; n30940
g30877 nor n30939 n30940 ; n30941
g30878 and n30930 n30941_not ; n30942
g30879 and n30930_not n30941 ; n30943
g30880 nor n30942 n30943 ; n30944
g30881 and n30895_not n30944 ; n30945
g30882 and n30895 n30944_not ; n30946
g30883 nor n30945 n30946 ; n30947
g30884 and n3884 n22309 ; n30948
g30885 and n3967 n22312 ; n30949
g30886 and n4046 n22315 ; n30950
g30887 nor n30949 n30950 ; n30951
g30888 and n30948_not n30951 ; n30952
g30889 and n4050 n22529_not ; n30953
g30890 and n30952 n30953_not ; n30954
g30891 and a[26] n30954_not ; n30955
g30892 and a[26] n30955_not ; n30956
g30893 nor n30954 n30955 ; n30957
g30894 nor n30956 n30957 ; n30958
g30895 and n30947 n30958_not ; n30959
g30896 and n30947 n30959_not ; n30960
g30897 nor n30958 n30959 ; n30961
g30898 nor n30960 n30961 ; n30962
g30899 nor n30821 n30827 ; n30963
g30900 and n30962 n30963 ; n30964
g30901 nor n30962 n30963 ; n30965
g30902 nor n30964 n30965 ; n30966
g30903 and n4694 n26060 ; n30967
g30904 and n4533 n26063 ; n30968
g30905 and n4604 n26066 ; n30969
g30906 nor n30968 n30969 ; n30970
g30907 and n30967_not n30970 ; n30971
g30908 and n4536 n26088_not ; n30972
g30909 and n30971 n30972_not ; n30973
g30910 and a[23] n30973_not ; n30974
g30911 and a[23] n30974_not ; n30975
g30912 nor n30973 n30974 ; n30976
g30913 nor n30975 n30976 ; n30977
g30914 and n30966 n30977_not ; n30978
g30915 and n30966 n30978_not ; n30979
g30916 nor n30977 n30978 ; n30980
g30917 nor n30979 n30980 ; n30981
g30918 nor n30841 n30846 ; n30982
g30919 nor n30981 n30982 ; n30983
g30920 nor n30981 n30983 ; n30984
g30921 nor n30982 n30983 ; n30985
g30922 nor n30984 n30985 ; n30986
g30923 and n5496 n27442 ; n30987
g30924 and n4935 n26890 ; n30988
g30925 and n5407 n27173 ; n30989
g30926 nor n30988 n30989 ; n30990
g30927 and n30987_not n30990 ; n30991
g30928 and n4938 n27455 ; n30992
g30929 and n30991 n30992_not ; n30993
g30930 and a[20] n30993_not ; n30994
g30931 and a[20] n30994_not ; n30995
g30932 nor n30993 n30994 ; n30996
g30933 nor n30995 n30996 ; n30997
g30934 nor n30986 n30997 ; n30998
g30935 nor n30986 n30998 ; n30999
g30936 nor n30997 n30998 ; n31000
g30937 nor n30999 n31000 ; n31001
g30938 nor n30859 n30865 ; n31002
g30939 and n31001 n31002 ; n31003
g30940 nor n31001 n31002 ; n31004
g30941 nor n31003 n31004 ; n31005
g30942 and n6233 n28208_not ; n31006
g30943 and n5663 n27698 ; n31007
g30944 and n5939 n27964 ; n31008
g30945 nor n31007 n31008 ; n31009
g30946 and n31006_not n31009 ; n31010
g30947 and n5666 n28223_not ; n31011
g30948 and n31010 n31011_not ; n31012
g30949 and a[17] n31012_not ; n31013
g30950 and a[17] n31013_not ; n31014
g30951 nor n31012 n31013 ; n31015
g30952 nor n31014 n31015 ; n31016
g30953 and n31005 n31016_not ; n31017
g30954 and n31005 n31017_not ; n31018
g30955 nor n31016 n31017 ; n31019
g30956 nor n31018 n31019 ; n31020
g30957 nor n30879 n30884 ; n31021
g30958 nor n31020 n31021 ; n31022
g30959 nor n31020 n31022 ; n31023
g30960 nor n31021 n31022 ; n31024
g30961 nor n31023 n31024 ; n31025
g30962 nor n30886 n30889 ; n31026
g30963 and n31025 n31026 ; n31027
g30964 nor n31025 n31026 ; n31028
g30965 nor n31027 n31028 ; n31029
g30966 and n30893 n31029_not ; n31030
g30967 and n30893_not n31029 ; n31031
g30968 or n31030 n31031 ; result[20]
g30969 nor n30929 n30942 ; n31033
g30970 nor n30920 n30923 ; n31034
g30971 and n242_not n1253 ; n31035
g30972 and n135_not n31035 ; n31036
g30973 and n376 n2026 ; n31037
g30974 and n31036 n31037 ; n31038
g30975 and n2263 n31038 ; n31039
g30976 and n5188 n31039 ; n31040
g30977 and n13247 n31040 ; n31041
g30978 and n1100 n31041 ; n31042
g30979 and n2506 n31042 ; n31043
g30980 and n1781 n31043 ; n31044
g30981 and n3739 n31044 ; n31045
g30982 and n1380 n31045 ; n31046
g30983 and n1306_not n31046 ; n31047
g30984 and n292_not n31047 ; n31048
g30985 and n240_not n31048 ; n31049
g30986 and n225_not n31049 ; n31050
g30987 and n525_not n31050 ; n31051
g30988 and n489_not n31051 ; n31052
g30989 and n30919 n31052_not ; n31053
g30990 and n30919_not n31052 ; n31054
g30991 nor n31034 n31054 ; n31055
g30992 and n31053_not n31055 ; n31056
g30993 nor n31034 n31056 ; n31057
g30994 nor n31054 n31056 ; n31058
g30995 and n31053_not n31058 ; n31059
g30996 nor n31057 n31059 ; n31060
g30997 and n75 n24616_not ; n31061
g30998 and n3020 n22326 ; n31062
g30999 and n3023 n22332 ; n31063
g31000 and n3028 n22329 ; n31064
g31001 nor n31063 n31064 ; n31065
g31002 and n31062_not n31065 ; n31066
g31003 and n31061_not n31066 ; n31067
g31004 nor n31060 n31067 ; n31068
g31005 nor n31060 n31068 ; n31069
g31006 nor n31067 n31068 ; n31070
g31007 nor n31069 n31070 ; n31071
g31008 and n3457 n22312 ; n31072
g31009 and n3542 n22323 ; n31073
g31010 and n3606 n22320 ; n31074
g31011 nor n31073 n31074 ; n31075
g31012 and n31072_not n31075 ; n31076
g31013 and n3368_not n31076 ; n31077
g31014 and n25315 n31076 ; n31078
g31015 nor n31077 n31078 ; n31079
g31016 and a[29] n31079_not ; n31080
g31017 and a[29]_not n31079 ; n31081
g31018 nor n31080 n31081 ; n31082
g31019 nor n31071 n31082 ; n31083
g31020 and n31071 n31082 ; n31084
g31021 nor n31083 n31084 ; n31085
g31022 and n31033_not n31085 ; n31086
g31023 and n31033 n31085_not ; n31087
g31024 nor n31086 n31087 ; n31088
g31025 and n3884 n26063 ; n31089
g31026 and n3967 n22315 ; n31090
g31027 and n4046 n22309 ; n31091
g31028 nor n31090 n31091 ; n31092
g31029 and n31089_not n31092 ; n31093
g31030 and n4050 n26604_not ; n31094
g31031 and n31093 n31094_not ; n31095
g31032 and a[26] n31095_not ; n31096
g31033 and a[26] n31096_not ; n31097
g31034 nor n31095 n31096 ; n31098
g31035 nor n31097 n31098 ; n31099
g31036 and n31088 n31099_not ; n31100
g31037 and n31088 n31100_not ; n31101
g31038 nor n31099 n31100 ; n31102
g31039 nor n31101 n31102 ; n31103
g31040 nor n30945 n30959 ; n31104
g31041 and n31103 n31104 ; n31105
g31042 nor n31103 n31104 ; n31106
g31043 nor n31105 n31106 ; n31107
g31044 and n4694 n26890 ; n31108
g31045 and n4533 n26066 ; n31109
g31046 and n4604 n26060 ; n31110
g31047 nor n31109 n31110 ; n31111
g31048 and n31108_not n31111 ; n31112
g31049 and n4536 n26904_not ; n31113
g31050 and n31112 n31113_not ; n31114
g31051 and a[23] n31114_not ; n31115
g31052 and a[23] n31115_not ; n31116
g31053 nor n31114 n31115 ; n31117
g31054 nor n31116 n31117 ; n31118
g31055 and n31107 n31118_not ; n31119
g31056 and n31107 n31119_not ; n31120
g31057 nor n31118 n31119 ; n31121
g31058 nor n31120 n31121 ; n31122
g31059 nor n30965 n30978 ; n31123
g31060 and n31122 n31123 ; n31124
g31061 nor n31122 n31123 ; n31125
g31062 nor n31124 n31125 ; n31126
g31063 and n5496 n27698 ; n31127
g31064 and n4935 n27173 ; n31128
g31065 and n5407 n27442 ; n31129
g31066 nor n31128 n31129 ; n31130
g31067 and n31127_not n31130 ; n31131
g31068 and n4938 n27713_not ; n31132
g31069 and n31131 n31132_not ; n31133
g31070 and a[20] n31133_not ; n31134
g31071 and a[20] n31134_not ; n31135
g31072 nor n31133 n31134 ; n31136
g31073 nor n31135 n31136 ; n31137
g31074 and n31126 n31137_not ; n31138
g31075 and n31126 n31138_not ; n31139
g31076 nor n31137 n31138 ; n31140
g31077 nor n31139 n31140 ; n31141
g31078 nor n30983 n30998 ; n31142
g31079 nor n13717 n28208 ; n31143
g31080 and n5663 n27964 ; n31144
g31081 nor n31143 n31144 ; n31145
g31082 and n5666_not n31145 ; n31146
g31083 and n28221 n31145 ; n31147
g31084 nor n31146 n31147 ; n31148
g31085 and a[17] n31148_not ; n31149
g31086 and a[17]_not n31148 ; n31150
g31087 nor n31149 n31150 ; n31151
g31088 nor n31142 n31151 ; n31152
g31089 and n31142 n31151 ; n31153
g31090 nor n31152 n31153 ; n31154
g31091 and n31141_not n31154 ; n31155
g31092 nor n31141 n31155 ; n31156
g31093 and n31154 n31155_not ; n31157
g31094 nor n31156 n31157 ; n31158
g31095 nor n31004 n31017 ; n31159
g31096 and n31158 n31159 ; n31160
g31097 nor n31158 n31159 ; n31161
g31098 nor n31160 n31161 ; n31162
g31099 nor n31022 n31028 ; n31163
g31100 and n31162_not n31163 ; n31164
g31101 and n31162 n31163_not ; n31165
g31102 nor n31164 n31165 ; n31166
g31103 and n30893 n31029 ; n31167
g31104 and n31166 n31167 ; n31168
g31105 nor n31166 n31167 ; n31169
g31106 nor n31168 n31169 ; result[21]
g31107 nor n31161 n31165 ; n31171
g31108 nor n31152 n31155 ; n31172
g31109 nor n31106 n31119 ; n31173
g31110 nor n31086 n31100 ; n31174
g31111 and n3884 n26066 ; n31175
g31112 and n3967 n22309 ; n31176
g31113 and n4046 n26063 ; n31177
g31114 nor n31176 n31177 ; n31178
g31115 and n31175_not n31178 ; n31179
g31116 and n4050 n26624_not ; n31180
g31117 and n31179 n31180_not ; n31181
g31118 and a[26] n31181_not ; n31182
g31119 and a[26] n31182_not ; n31183
g31120 nor n31181 n31182 ; n31184
g31121 nor n31183 n31184 ; n31185
g31122 nor n31174 n31185 ; n31186
g31123 nor n31174 n31186 ; n31187
g31124 nor n31185 n31186 ; n31188
g31125 nor n31187 n31188 ; n31189
g31126 nor n31068 n31083 ; n31190
g31127 and n75 n24599 ; n31191
g31128 and n3020 n22323 ; n31192
g31129 and n3023 n22329 ; n31193
g31130 and n3028 n22326 ; n31194
g31131 nor n31193 n31194 ; n31195
g31132 and n31192_not n31195 ; n31196
g31133 and n31191_not n31196 ; n31197
g31134 nor n13719 n28208 ; n31198
g31135 and a[17] n31198_not ; n31199
g31136 and a[17]_not n31198 ; n31200
g31137 nor n31199 n31200 ; n31201
g31138 and n1143 n24041 ; n31202
g31139 and n2719 n31202 ; n31203
g31140 and n4785 n31203 ; n31204
g31141 and n3282 n31204 ; n31205
g31142 and n12924 n31205 ; n31206
g31143 and n882 n31206 ; n31207
g31144 and n448 n31207 ; n31208
g31145 and n279 n31208 ; n31209
g31146 and n229_not n31209 ; n31210
g31147 and n335_not n31210 ; n31211
g31148 and n299_not n31211 ; n31212
g31149 and n525_not n31212 ; n31213
g31150 and n771_not n31213 ; n31214
g31151 and n31052 n31214 ; n31215
g31152 nor n31052 n31214 ; n31216
g31153 nor n31215 n31216 ; n31217
g31154 and n31201 n31217 ; n31218
g31155 nor n31201 n31217 ; n31219
g31156 nor n31218 n31219 ; n31220
g31157 and n31197_not n31220 ; n31221
g31158 and n31220 n31221_not ; n31222
g31159 nor n31197 n31221 ; n31223
g31160 nor n31222 n31223 ; n31224
g31161 nor n31058 n31224 ; n31225
g31162 nor n31224 n31225 ; n31226
g31163 nor n31058 n31225 ; n31227
g31164 nor n31226 n31227 ; n31228
g31165 nor n31190 n31228 ; n31229
g31166 nor n31190 n31229 ; n31230
g31167 nor n31228 n31229 ; n31231
g31168 nor n31230 n31231 ; n31232
g31169 and n3457 n22315 ; n31233
g31170 and n3542 n22320 ; n31234
g31171 and n3606 n22312 ; n31235
g31172 nor n31234 n31235 ; n31236
g31173 and n31233_not n31236 ; n31237
g31174 and n3368 n25294 ; n31238
g31175 and n31237 n31238_not ; n31239
g31176 and a[29] n31239_not ; n31240
g31177 and a[29] n31240_not ; n31241
g31178 nor n31239 n31240 ; n31242
g31179 nor n31241 n31242 ; n31243
g31180 nor n31232 n31243 ; n31244
g31181 nor n31232 n31244 ; n31245
g31182 nor n31243 n31244 ; n31246
g31183 nor n31245 n31246 ; n31247
g31184 and n31189_not n31247 ; n31248
g31185 and n31189 n31247_not ; n31249
g31186 nor n31248 n31249 ; n31250
g31187 and n4694 n27173 ; n31251
g31188 and n4533 n26060 ; n31252
g31189 and n4604 n26890 ; n31253
g31190 nor n31252 n31253 ; n31254
g31191 and n31251_not n31254 ; n31255
g31192 and n4536 n27185 ; n31256
g31193 and n31255 n31256_not ; n31257
g31194 and a[23] n31257_not ; n31258
g31195 and a[23] n31258_not ; n31259
g31196 nor n31257 n31258 ; n31260
g31197 nor n31259 n31260 ; n31261
g31198 nor n31250 n31261 ; n31262
g31199 and n31250 n31261 ; n31263
g31200 nor n31262 n31263 ; n31264
g31201 and n31173 n31264_not ; n31265
g31202 and n31173_not n31264 ; n31266
g31203 nor n31265 n31266 ; n31267
g31204 nor n31125 n31138 ; n31268
g31205 and n5496 n27964 ; n31269
g31206 and n4935 n27442 ; n31270
g31207 and n5407 n27698 ; n31271
g31208 nor n31270 n31271 ; n31272
g31209 and n31269_not n31272 ; n31273
g31210 and n4938 n27976 ; n31274
g31211 and n31273 n31274_not ; n31275
g31212 and a[20] n31275_not ; n31276
g31213 and a[20] n31276_not ; n31277
g31214 nor n31275 n31276 ; n31278
g31215 nor n31277 n31278 ; n31279
g31216 nor n31268 n31279 ; n31280
g31217 nor n31268 n31280 ; n31281
g31218 nor n31279 n31280 ; n31282
g31219 nor n31281 n31282 ; n31283
g31220 and n31267_not n31283 ; n31284
g31221 and n31267 n31283_not ; n31285
g31222 nor n31284 n31285 ; n31286
g31223 and n31172_not n31286 ; n31287
g31224 and n31172 n31286_not ; n31288
g31225 nor n31287 n31288 ; n31289
g31226 and n31171_not n31289 ; n31290
g31227 and n31171 n31289_not ; n31291
g31228 nor n31290 n31291 ; n31292
g31229 nor n31168 n31292 ; n31293
g31230 and n31168 n31292 ; n31294
g31231 nor n31293 n31294 ; result[22]
g31232 nor n31229 n31244 ; n31296
g31233 and n75 n25270_not ; n31297
g31234 and n3020 n22320 ; n31298
g31235 and n3023 n22326 ; n31299
g31236 and n3028 n22323 ; n31300
g31237 nor n31299 n31300 ; n31301
g31238 and n31298_not n31301 ; n31302
g31239 and n31297_not n31302 ; n31303
g31240 nor n31216 n31218 ; n31304
g31241 and n632 n13014 ; n31305
g31242 and n2656 n31305 ; n31306
g31243 and n6514 n31306 ; n31307
g31244 and n2543 n31307 ; n31308
g31245 and n3497 n31308 ; n31309
g31246 and n29550 n31309 ; n31310
g31247 and n423 n31310 ; n31311
g31248 and n418 n31311 ; n31312
g31249 and n4101 n31312 ; n31313
g31250 and n330_not n31313 ; n31314
g31251 and n329_not n31314 ; n31315
g31252 and n280_not n31315 ; n31316
g31253 and n203_not n31316 ; n31317
g31254 and n619_not n31317 ; n31318
g31255 and n536_not n31318 ; n31319
g31256 and n31304_not n31319 ; n31320
g31257 and n31304 n31319_not ; n31321
g31258 nor n31320 n31321 ; n31322
g31259 and n31303_not n31322 ; n31323
g31260 nor n31303 n31323 ; n31324
g31261 and n31322 n31323_not ; n31325
g31262 nor n31324 n31325 ; n31326
g31263 nor n31221 n31225 ; n31327
g31264 and n31326 n31327 ; n31328
g31265 nor n31326 n31327 ; n31329
g31266 nor n31328 n31329 ; n31330
g31267 and n3457 n22309 ; n31331
g31268 and n3542 n22312 ; n31332
g31269 and n3606 n22315 ; n31333
g31270 nor n31332 n31333 ; n31334
g31271 and n31331_not n31334 ; n31335
g31272 and n3368_not n31335 ; n31336
g31273 and n22529 n31335 ; n31337
g31274 nor n31336 n31337 ; n31338
g31275 and a[29] n31338_not ; n31339
g31276 and a[29]_not n31338 ; n31340
g31277 nor n31339 n31340 ; n31341
g31278 and n31330 n31341_not ; n31342
g31279 and n31330_not n31341 ; n31343
g31280 nor n31342 n31343 ; n31344
g31281 and n31296_not n31344 ; n31345
g31282 and n31296 n31344_not ; n31346
g31283 nor n31345 n31346 ; n31347
g31284 and n3884 n26060 ; n31348
g31285 and n3967 n26063 ; n31349
g31286 and n4046 n26066 ; n31350
g31287 nor n31349 n31350 ; n31351
g31288 and n31348_not n31351 ; n31352
g31289 and n4050 n26088_not ; n31353
g31290 and n31352 n31353_not ; n31354
g31291 and a[26] n31354_not ; n31355
g31292 and a[26] n31355_not ; n31356
g31293 nor n31354 n31355 ; n31357
g31294 nor n31356 n31357 ; n31358
g31295 and n31347 n31358_not ; n31359
g31296 and n31347 n31359_not ; n31360
g31297 nor n31358 n31359 ; n31361
g31298 nor n31360 n31361 ; n31362
g31299 nor n31189 n31247 ; n31363
g31300 nor n31186 n31363 ; n31364
g31301 nor n31362 n31364 ; n31365
g31302 nor n31362 n31365 ; n31366
g31303 nor n31364 n31365 ; n31367
g31304 nor n31366 n31367 ; n31368
g31305 and n4694 n27442 ; n31369
g31306 and n4533 n26890 ; n31370
g31307 and n4604 n27173 ; n31371
g31308 nor n31370 n31371 ; n31372
g31309 and n31369_not n31372 ; n31373
g31310 and n4536 n27455 ; n31374
g31311 and n31373 n31374_not ; n31375
g31312 and a[23] n31375_not ; n31376
g31313 and a[23] n31376_not ; n31377
g31314 nor n31375 n31376 ; n31378
g31315 nor n31377 n31378 ; n31379
g31316 nor n31368 n31379 ; n31380
g31317 nor n31368 n31380 ; n31381
g31318 nor n31379 n31380 ; n31382
g31319 nor n31381 n31382 ; n31383
g31320 nor n31262 n31266 ; n31384
g31321 and n31383 n31384 ; n31385
g31322 nor n31383 n31384 ; n31386
g31323 nor n31385 n31386 ; n31387
g31324 and n5496 n28208_not ; n31388
g31325 and n4935 n27698 ; n31389
g31326 and n5407 n27964 ; n31390
g31327 nor n31389 n31390 ; n31391
g31328 and n31388_not n31391 ; n31392
g31329 and n4938 n28223_not ; n31393
g31330 and n31392 n31393_not ; n31394
g31331 and a[20] n31394_not ; n31395
g31332 and a[20] n31395_not ; n31396
g31333 nor n31394 n31395 ; n31397
g31334 nor n31396 n31397 ; n31398
g31335 and n31387 n31398_not ; n31399
g31336 and n31387 n31399_not ; n31400
g31337 nor n31398 n31399 ; n31401
g31338 nor n31400 n31401 ; n31402
g31339 nor n31280 n31285 ; n31403
g31340 nor n31402 n31403 ; n31404
g31341 nor n31402 n31404 ; n31405
g31342 nor n31403 n31404 ; n31406
g31343 nor n31405 n31406 ; n31407
g31344 nor n31287 n31290 ; n31408
g31345 and n31407 n31408 ; n31409
g31346 nor n31407 n31408 ; n31410
g31347 nor n31409 n31410 ; n31411
g31348 and n31294_not n31411 ; n31412
g31349 and n31294 n31411_not ; n31413
g31350 or n31412 n31413 ; result[23]
g31351 and n31294 n31411 ; n31415
g31352 and n75 n25315_not ; n31416
g31353 and n3020 n22312 ; n31417
g31354 and n3023 n22323 ; n31418
g31355 and n3028 n22320 ; n31419
g31356 nor n31418 n31419 ; n31420
g31357 and n31417_not n31420 ; n31421
g31358 and n31416_not n31421 ; n31422
g31359 and n12941 n31036 ; n31423
g31360 and n4366 n31423 ; n31424
g31361 and n6561 n31424 ; n31425
g31362 and n3259 n31425 ; n31426
g31363 and n2651 n31426 ; n31427
g31364 and n2683 n31427 ; n31428
g31365 and n230 n31428 ; n31429
g31366 and n488 n31429 ; n31430
g31367 and n28688 n31430 ; n31431
g31368 and n602_not n31431 ; n31432
g31369 and n1101_not n31432 ; n31433
g31370 and n142_not n31433 ; n31434
g31371 and n125_not n31434 ; n31435
g31372 and n31319_not n31435 ; n31436
g31373 and n31319 n31435_not ; n31437
g31374 nor n31422 n31437 ; n31438
g31375 and n31436_not n31438 ; n31439
g31376 nor n31422 n31439 ; n31440
g31377 nor n31437 n31439 ; n31441
g31378 and n31436_not n31441 ; n31442
g31379 nor n31440 n31442 ; n31443
g31380 nor n31320 n31323 ; n31444
g31381 and n31443 n31444 ; n31445
g31382 nor n31443 n31444 ; n31446
g31383 nor n31445 n31446 ; n31447
g31384 nor n31329 n31342 ; n31448
g31385 and n31447_not n31448 ; n31449
g31386 and n31447 n31448_not ; n31450
g31387 nor n31449 n31450 ; n31451
g31388 and n3457 n26063 ; n31452
g31389 and n3542 n22315 ; n31453
g31390 and n3606 n22309 ; n31454
g31391 nor n31453 n31454 ; n31455
g31392 and n31452_not n31455 ; n31456
g31393 and n3368 n26604_not ; n31457
g31394 and n31456 n31457_not ; n31458
g31395 and a[29] n31458_not ; n31459
g31396 and a[29] n31459_not ; n31460
g31397 nor n31458 n31459 ; n31461
g31398 nor n31460 n31461 ; n31462
g31399 and n31451 n31462_not ; n31463
g31400 and n31451 n31463_not ; n31464
g31401 nor n31462 n31463 ; n31465
g31402 nor n31464 n31465 ; n31466
g31403 and n3884 n26890 ; n31467
g31404 and n3967 n26066 ; n31468
g31405 and n4046 n26060 ; n31469
g31406 nor n31468 n31469 ; n31470
g31407 and n31467_not n31470 ; n31471
g31408 and n4050 n26904_not ; n31472
g31409 and n31471 n31472_not ; n31473
g31410 and a[26] n31473_not ; n31474
g31411 and a[26] n31474_not ; n31475
g31412 nor n31473 n31474 ; n31476
g31413 nor n31475 n31476 ; n31477
g31414 nor n31466 n31477 ; n31478
g31415 nor n31466 n31478 ; n31479
g31416 nor n31477 n31478 ; n31480
g31417 nor n31479 n31480 ; n31481
g31418 nor n31345 n31359 ; n31482
g31419 and n31481 n31482 ; n31483
g31420 nor n31481 n31482 ; n31484
g31421 nor n31483 n31484 ; n31485
g31422 and n4694 n27698 ; n31486
g31423 and n4533 n27173 ; n31487
g31424 and n4604 n27442 ; n31488
g31425 nor n31487 n31488 ; n31489
g31426 and n31486_not n31489 ; n31490
g31427 and n4536 n27713_not ; n31491
g31428 and n31490 n31491_not ; n31492
g31429 and a[23] n31492_not ; n31493
g31430 and a[23] n31493_not ; n31494
g31431 nor n31492 n31493 ; n31495
g31432 nor n31494 n31495 ; n31496
g31433 and n31485 n31496_not ; n31497
g31434 and n31485 n31497_not ; n31498
g31435 nor n31496 n31497 ; n31499
g31436 nor n31498 n31499 ; n31500
g31437 nor n31365 n31380 ; n31501
g31438 nor n13439 n28208 ; n31502
g31439 and n4935 n27964 ; n31503
g31440 nor n31502 n31503 ; n31504
g31441 and n4938_not n31504 ; n31505
g31442 and n28221 n31504 ; n31506
g31443 nor n31505 n31506 ; n31507
g31444 and a[20] n31507_not ; n31508
g31445 and a[20]_not n31507 ; n31509
g31446 nor n31508 n31509 ; n31510
g31447 nor n31501 n31510 ; n31511
g31448 and n31501 n31510 ; n31512
g31449 nor n31511 n31512 ; n31513
g31450 and n31500_not n31513 ; n31514
g31451 nor n31500 n31514 ; n31515
g31452 and n31513 n31514_not ; n31516
g31453 nor n31515 n31516 ; n31517
g31454 nor n31386 n31399 ; n31518
g31455 and n31517 n31518 ; n31519
g31456 nor n31517 n31518 ; n31520
g31457 nor n31519 n31520 ; n31521
g31458 nor n31404 n31410 ; n31522
g31459 and n31521_not n31522 ; n31523
g31460 and n31521 n31522_not ; n31524
g31461 nor n31523 n31524 ; n31525
g31462 and n31415 n31525 ; n31526
g31463 nor n31415 n31525 ; n31527
g31464 nor n31526 n31527 ; result[24]
g31465 nor n31520 n31524 ; n31529
g31466 nor n31511 n31514 ; n31530
g31467 and n75 n25294 ; n31531
g31468 and n3020 n22315 ; n31532
g31469 and n3023 n22320 ; n31533
g31470 and n3028 n22312 ; n31534
g31471 nor n31533 n31534 ; n31535
g31472 and n31532_not n31535 ; n31536
g31473 and n31531_not n31536 ; n31537
g31474 nor n13441 n28208 ; n31538
g31475 and a[20] n31538_not ; n31539
g31476 and a[20]_not n31538 ; n31540
g31477 nor n31539 n31540 ; n31541
g31478 and n2753 n3370 ; n31542
g31479 and n530 n31542 ; n31543
g31480 and n15050 n31543 ; n31544
g31481 and n15953 n31544 ; n31545
g31482 and n4293 n31545 ; n31546
g31483 and n1008 n31546 ; n31547
g31484 and n805 n31547 ; n31548
g31485 and n539 n31548 ; n31549
g31486 and n2506 n31549 ; n31550
g31487 and n615 n31550 ; n31551
g31488 and n1574 n31551 ; n31552
g31489 and n558_not n31552 ; n31553
g31490 and n420_not n31553 ; n31554
g31491 and n189_not n31554 ; n31555
g31492 and n716_not n31555 ; n31556
g31493 and n452_not n31556 ; n31557
g31494 and n201_not n31557 ; n31558
g31495 and n31319 n31558 ; n31559
g31496 nor n31319 n31558 ; n31560
g31497 nor n31559 n31560 ; n31561
g31498 and n31541 n31561 ; n31562
g31499 nor n31541 n31561 ; n31563
g31500 nor n31562 n31563 ; n31564
g31501 and n31441_not n31564 ; n31565
g31502 and n31441 n31564_not ; n31566
g31503 nor n31565 n31566 ; n31567
g31504 and n31537_not n31567 ; n31568
g31505 and n31567 n31568_not ; n31569
g31506 nor n31537 n31568 ; n31570
g31507 nor n31569 n31570 ; n31571
g31508 nor n31446 n31450 ; n31572
g31509 and n31571 n31572 ; n31573
g31510 nor n31571 n31572 ; n31574
g31511 nor n31573 n31574 ; n31575
g31512 and n3457 n26066 ; n31576
g31513 and n3542 n22309 ; n31577
g31514 and n3606 n26063 ; n31578
g31515 nor n31577 n31578 ; n31579
g31516 and n31576_not n31579 ; n31580
g31517 and n3368 n26624_not ; n31581
g31518 and n31580 n31581_not ; n31582
g31519 and a[29] n31582_not ; n31583
g31520 and a[29] n31583_not ; n31584
g31521 nor n31582 n31583 ; n31585
g31522 nor n31584 n31585 ; n31586
g31523 and n31575 n31586_not ; n31587
g31524 and n31575 n31587_not ; n31588
g31525 nor n31586 n31587 ; n31589
g31526 nor n31588 n31589 ; n31590
g31527 and n3884 n27173 ; n31591
g31528 and n3967 n26060 ; n31592
g31529 and n4046 n26890 ; n31593
g31530 nor n31592 n31593 ; n31594
g31531 and n31591_not n31594 ; n31595
g31532 and n4050 n27185 ; n31596
g31533 and n31595 n31596_not ; n31597
g31534 and a[26] n31597_not ; n31598
g31535 and a[26] n31598_not ; n31599
g31536 nor n31597 n31598 ; n31600
g31537 nor n31599 n31600 ; n31601
g31538 nor n31590 n31601 ; n31602
g31539 nor n31590 n31602 ; n31603
g31540 nor n31601 n31602 ; n31604
g31541 nor n31603 n31604 ; n31605
g31542 nor n31463 n31478 ; n31606
g31543 and n31605 n31606 ; n31607
g31544 nor n31605 n31606 ; n31608
g31545 nor n31607 n31608 ; n31609
g31546 nor n31484 n31497 ; n31610
g31547 and n4694 n27964 ; n31611
g31548 and n4533 n27442 ; n31612
g31549 and n4604 n27698 ; n31613
g31550 nor n31612 n31613 ; n31614
g31551 and n31611_not n31614 ; n31615
g31552 and n4536 n27976 ; n31616
g31553 and n31615 n31616_not ; n31617
g31554 and a[23] n31617_not ; n31618
g31555 and a[23] n31618_not ; n31619
g31556 nor n31617 n31618 ; n31620
g31557 nor n31619 n31620 ; n31621
g31558 nor n31610 n31621 ; n31622
g31559 nor n31610 n31622 ; n31623
g31560 nor n31621 n31622 ; n31624
g31561 nor n31623 n31624 ; n31625
g31562 and n31609_not n31625 ; n31626
g31563 and n31609 n31625_not ; n31627
g31564 nor n31626 n31627 ; n31628
g31565 and n31530_not n31628 ; n31629
g31566 and n31530 n31628_not ; n31630
g31567 nor n31629 n31630 ; n31631
g31568 and n31529_not n31631 ; n31632
g31569 and n31529 n31631_not ; n31633
g31570 nor n31632 n31633 ; n31634
g31571 nor n31526 n31634 ; n31635
g31572 and n31526 n31634 ; n31636
g31573 nor n31635 n31636 ; result[25]
g31574 nor n31574 n31587 ; n31638
g31575 and n75 n22529_not ; n31639
g31576 and n3020 n22309 ; n31640
g31577 and n3023 n22312 ; n31641
g31578 and n3028 n22315 ; n31642
g31579 nor n31641 n31642 ; n31643
g31580 and n31640_not n31643 ; n31644
g31581 and n31639_not n31644 ; n31645
g31582 nor n31560 n31562 ; n31646
g31583 and n1740 n4828 ; n31647
g31584 and n1604 n31647 ; n31648
g31585 and n1640 n31648 ; n31649
g31586 and n14534 n31649 ; n31650
g31587 and n1029 n31650 ; n31651
g31588 and n3282 n31651 ; n31652
g31589 and n1679 n31652 ; n31653
g31590 and n3039 n31653 ; n31654
g31591 and n16055 n31654 ; n31655
g31592 and n1252 n31655 ; n31656
g31593 and n1246_not n31656 ; n31657
g31594 and n602_not n31657 ; n31658
g31595 and n145_not n31658 ; n31659
g31596 and n298_not n31659 ; n31660
g31597 and n222_not n31660 ; n31661
g31598 and n31646_not n31661 ; n31662
g31599 and n31646 n31661_not ; n31663
g31600 nor n31662 n31663 ; n31664
g31601 and n31645_not n31664 ; n31665
g31602 nor n31645 n31665 ; n31666
g31603 and n31664 n31665_not ; n31667
g31604 nor n31666 n31667 ; n31668
g31605 nor n31565 n31568 ; n31669
g31606 and n31668 n31669 ; n31670
g31607 nor n31668 n31669 ; n31671
g31608 nor n31670 n31671 ; n31672
g31609 and n3457 n26060 ; n31673
g31610 and n3542 n26063 ; n31674
g31611 and n3606 n26066 ; n31675
g31612 nor n31674 n31675 ; n31676
g31613 and n31673_not n31676 ; n31677
g31614 and n3368_not n31677 ; n31678
g31615 and n26088 n31677 ; n31679
g31616 nor n31678 n31679 ; n31680
g31617 and a[29] n31680_not ; n31681
g31618 and a[29]_not n31680 ; n31682
g31619 nor n31681 n31682 ; n31683
g31620 and n31672 n31683_not ; n31684
g31621 and n31672_not n31683 ; n31685
g31622 nor n31684 n31685 ; n31686
g31623 and n31638_not n31686 ; n31687
g31624 and n31638 n31686_not ; n31688
g31625 nor n31687 n31688 ; n31689
g31626 and n3884 n27442 ; n31690
g31627 and n3967 n26890 ; n31691
g31628 and n4046 n27173 ; n31692
g31629 nor n31691 n31692 ; n31693
g31630 and n31690_not n31693 ; n31694
g31631 and n4050 n27455 ; n31695
g31632 and n31694 n31695_not ; n31696
g31633 and a[26] n31696_not ; n31697
g31634 and a[26] n31697_not ; n31698
g31635 nor n31696 n31697 ; n31699
g31636 nor n31698 n31699 ; n31700
g31637 and n31689 n31700_not ; n31701
g31638 and n31689 n31701_not ; n31702
g31639 nor n31700 n31701 ; n31703
g31640 nor n31702 n31703 ; n31704
g31641 nor n31602 n31608 ; n31705
g31642 and n31704 n31705 ; n31706
g31643 nor n31704 n31705 ; n31707
g31644 nor n31706 n31707 ; n31708
g31645 and n4694 n28208_not ; n31709
g31646 and n4533 n27698 ; n31710
g31647 and n4604 n27964 ; n31711
g31648 nor n31710 n31711 ; n31712
g31649 and n31709_not n31712 ; n31713
g31650 and n4536 n28223_not ; n31714
g31651 and n31713 n31714_not ; n31715
g31652 and a[23] n31715_not ; n31716
g31653 and a[23] n31716_not ; n31717
g31654 nor n31715 n31716 ; n31718
g31655 nor n31717 n31718 ; n31719
g31656 and n31708 n31719_not ; n31720
g31657 and n31708 n31720_not ; n31721
g31658 nor n31719 n31720 ; n31722
g31659 nor n31721 n31722 ; n31723
g31660 nor n31622 n31627 ; n31724
g31661 nor n31723 n31724 ; n31725
g31662 nor n31723 n31725 ; n31726
g31663 nor n31724 n31725 ; n31727
g31664 nor n31726 n31727 ; n31728
g31665 nor n31629 n31632 ; n31729
g31666 and n31728 n31729 ; n31730
g31667 nor n31728 n31729 ; n31731
g31668 nor n31730 n31731 ; n31732
g31669 and n31636 n31732_not ; n31733
g31670 and n31636_not n31732 ; n31734
g31671 or n31733 n31734 ; result[26]
g31672 nor n31662 n31665 ; n31736
g31673 and n3459 n13016 ; n31737
g31674 and n1070 n31737 ; n31738
g31675 and n15882 n31738 ; n31739
g31676 and n25863 n31739 ; n31740
g31677 and n4232 n31740 ; n31741
g31678 and n2651 n31741 ; n31742
g31679 and n29538 n31742 ; n31743
g31680 and n285 n31743 ; n31744
g31681 and n1252 n31744 ; n31745
g31682 and n720 n31745 ; n31746
g31683 and n22762 n31746 ; n31747
g31684 and n334_not n31747 ; n31748
g31685 and n233_not n31748 ; n31749
g31686 and n302_not n31749 ; n31750
g31687 and n714_not n31750 ; n31751
g31688 and n31661 n31751_not ; n31752
g31689 and n31661_not n31751 ; n31753
g31690 nor n31736 n31753 ; n31754
g31691 and n31752_not n31754 ; n31755
g31692 nor n31736 n31755 ; n31756
g31693 nor n31753 n31755 ; n31757
g31694 and n31752_not n31757 ; n31758
g31695 nor n31756 n31758 ; n31759
g31696 and n75 n26604_not ; n31760
g31697 and n3020 n26063 ; n31761
g31698 and n3023 n22315 ; n31762
g31699 and n3028 n22309 ; n31763
g31700 nor n31762 n31763 ; n31764
g31701 and n31761_not n31764 ; n31765
g31702 and n31760_not n31765 ; n31766
g31703 nor n31759 n31766 ; n31767
g31704 nor n31759 n31767 ; n31768
g31705 nor n31766 n31767 ; n31769
g31706 nor n31768 n31769 ; n31770
g31707 nor n31671 n31684 ; n31771
g31708 and n31770 n31771 ; n31772
g31709 nor n31770 n31771 ; n31773
g31710 nor n31772 n31773 ; n31774
g31711 and n3457 n26890 ; n31775
g31712 and n3542 n26066 ; n31776
g31713 and n3606 n26060 ; n31777
g31714 nor n31776 n31777 ; n31778
g31715 and n31775_not n31778 ; n31779
g31716 and n3368 n26904_not ; n31780
g31717 and n31779 n31780_not ; n31781
g31718 and a[29] n31781_not ; n31782
g31719 and a[29] n31782_not ; n31783
g31720 nor n31781 n31782 ; n31784
g31721 nor n31783 n31784 ; n31785
g31722 and n31774 n31785_not ; n31786
g31723 and n31774 n31786_not ; n31787
g31724 nor n31785 n31786 ; n31788
g31725 nor n31787 n31788 ; n31789
g31726 and n3884 n27698 ; n31790
g31727 and n3967 n27173 ; n31791
g31728 and n4046 n27442 ; n31792
g31729 nor n31791 n31792 ; n31793
g31730 and n31790_not n31793 ; n31794
g31731 and n4050 n27713_not ; n31795
g31732 and n31794 n31795_not ; n31796
g31733 and a[26] n31796_not ; n31797
g31734 and a[26] n31797_not ; n31798
g31735 nor n31796 n31797 ; n31799
g31736 nor n31798 n31799 ; n31800
g31737 nor n31789 n31800 ; n31801
g31738 nor n31789 n31801 ; n31802
g31739 nor n31800 n31801 ; n31803
g31740 nor n31802 n31803 ; n31804
g31741 nor n31687 n31701 ; n31805
g31742 nor n13938 n28208 ; n31806
g31743 and n4533 n27964 ; n31807
g31744 nor n31806 n31807 ; n31808
g31745 and n4536_not n31808 ; n31809
g31746 and n28221 n31808 ; n31810
g31747 nor n31809 n31810 ; n31811
g31748 and a[23] n31811_not ; n31812
g31749 and a[23]_not n31811 ; n31813
g31750 nor n31812 n31813 ; n31814
g31751 nor n31805 n31814 ; n31815
g31752 and n31805 n31814 ; n31816
g31753 nor n31815 n31816 ; n31817
g31754 and n31804_not n31817 ; n31818
g31755 nor n31804 n31818 ; n31819
g31756 and n31817 n31818_not ; n31820
g31757 nor n31819 n31820 ; n31821
g31758 nor n31707 n31720 ; n31822
g31759 and n31821 n31822 ; n31823
g31760 nor n31821 n31822 ; n31824
g31761 nor n31823 n31824 ; n31825
g31762 nor n31725 n31731 ; n31826
g31763 and n31825_not n31826 ; n31827
g31764 and n31825 n31826_not ; n31828
g31765 nor n31827 n31828 ; n31829
g31766 and n31636 n31732 ; n31830
g31767 and n31829 n31830 ; n31831
g31768 nor n31829 n31830 ; n31832
g31769 nor n31831 n31832 ; result[27]
g31770 nor n31824 n31828 ; n31834
g31771 nor n31815 n31818 ; n31835
g31772 nor n31786 n31801 ; n31836
g31773 and n3884 n27964 ; n31837
g31774 and n3967 n27442 ; n31838
g31775 and n4046 n27698 ; n31839
g31776 nor n31838 n31839 ; n31840
g31777 and n31837_not n31840 ; n31841
g31778 and n4050 n27976 ; n31842
g31779 and n31841 n31842_not ; n31843
g31780 and a[26] n31843_not ; n31844
g31781 and a[26] n31844_not ; n31845
g31782 nor n31843 n31844 ; n31846
g31783 nor n31845 n31846 ; n31847
g31784 nor n31836 n31847 ; n31848
g31785 nor n31836 n31848 ; n31849
g31786 nor n31847 n31848 ; n31850
g31787 nor n31849 n31850 ; n31851
g31788 and n75 n26624_not ; n31852
g31789 and n3020 n26066 ; n31853
g31790 and n3023 n22309 ; n31854
g31791 and n3028 n26063 ; n31855
g31792 nor n31854 n31855 ; n31856
g31793 and n31853_not n31856 ; n31857
g31794 and n31852_not n31857 ; n31858
g31795 nor n22248 n28208 ; n31859
g31796 and a[23] n31859_not ; n31860
g31797 and a[23]_not n31859 ; n31861
g31798 nor n31860 n31861 ; n31862
g31799 and n4799 n13161 ; n31863
g31800 and n1155 n31863 ; n31864
g31801 and n4003 n31864 ; n31865
g31802 and n3866 n31865 ; n31866
g31803 and n288 n31866 ; n31867
g31804 and n937 n31867 ; n31868
g31805 and n1478 n31868 ; n31869
g31806 and n193 n31869 ; n31870
g31807 and n509_not n31870 ; n31871
g31808 and n1011_not n31871 ; n31872
g31809 and n228_not n31872 ; n31873
g31810 and n825_not n31873 ; n31874
g31811 and n568_not n31874 ; n31875
g31812 and n519_not n31875 ; n31876
g31813 and n31751 n31876 ; n31877
g31814 nor n31751 n31876 ; n31878
g31815 nor n31877 n31878 ; n31879
g31816 and n31862 n31879 ; n31880
g31817 nor n31862 n31879 ; n31881
g31818 nor n31880 n31881 ; n31882
g31819 and n31757_not n31882 ; n31883
g31820 and n31757 n31882_not ; n31884
g31821 nor n31883 n31884 ; n31885
g31822 and n31858_not n31885 ; n31886
g31823 and n31885 n31886_not ; n31887
g31824 nor n31858 n31886 ; n31888
g31825 nor n31887 n31888 ; n31889
g31826 nor n31767 n31773 ; n31890
g31827 and n31889 n31890 ; n31891
g31828 nor n31889 n31890 ; n31892
g31829 nor n31891 n31892 ; n31893
g31830 and n3457 n27173 ; n31894
g31831 and n3542 n26060 ; n31895
g31832 and n3606 n26890 ; n31896
g31833 nor n31895 n31896 ; n31897
g31834 and n31894_not n31897 ; n31898
g31835 and n3368 n27185 ; n31899
g31836 and n31898 n31899_not ; n31900
g31837 and a[29] n31900_not ; n31901
g31838 and a[29] n31901_not ; n31902
g31839 nor n31900 n31901 ; n31903
g31840 nor n31902 n31903 ; n31904
g31841 and n31893 n31904_not ; n31905
g31842 and n31893 n31905_not ; n31906
g31843 nor n31904 n31905 ; n31907
g31844 nor n31906 n31907 ; n31908
g31845 and n31851_not n31908 ; n31909
g31846 and n31851 n31908_not ; n31910
g31847 nor n31909 n31910 ; n31911
g31848 nor n31835 n31911 ; n31912
g31849 and n31835 n31911 ; n31913
g31850 nor n31912 n31913 ; n31914
g31851 and n31834_not n31914 ; n31915
g31852 and n31834 n31914_not ; n31916
g31853 nor n31915 n31916 ; n31917
g31854 nor n31831 n31917 ; n31918
g31855 and n31831 n31917 ; n31919
g31856 nor n31918 n31919 ; result[28]
g31857 nor n31892 n31905 ; n31921
g31858 and n75 n26088_not ; n31922
g31859 and n3020 n26060 ; n31923
g31860 and n3023 n26063 ; n31924
g31861 and n3028 n26066 ; n31925
g31862 nor n31924 n31925 ; n31926
g31863 and n31923_not n31926 ; n31927
g31864 and n31922_not n31927 ; n31928
g31865 nor n31878 n31880 ; n31929
g31866 and n1738 n15012 ; n31930
g31867 and n3438 n31930 ; n31931
g31868 and n6610 n31931 ; n31932
g31869 and n26016 n31932 ; n31933
g31870 and n15880 n31933 ; n31934
g31871 and n3939 n31934 ; n31935
g31872 and n3997 n31935 ; n31936
g31873 and n1183 n31936 ; n31937
g31874 and n1531 n31937 ; n31938
g31875 and n1366 n31938 ; n31939
g31876 and n1783 n31939 ; n31940
g31877 and n100 n31940 ; n31941
g31878 and n420_not n31941 ; n31942
g31879 and n466_not n31942 ; n31943
g31880 and n298_not n31943 ; n31944
g31881 and n251_not n31944 ; n31945
g31882 and n31929_not n31945 ; n31946
g31883 and n31929 n31945_not ; n31947
g31884 nor n31946 n31947 ; n31948
g31885 and n31928_not n31948 ; n31949
g31886 nor n31928 n31949 ; n31950
g31887 and n31948 n31949_not ; n31951
g31888 nor n31950 n31951 ; n31952
g31889 nor n31883 n31886 ; n31953
g31890 and n31952 n31953 ; n31954
g31891 nor n31952 n31953 ; n31955
g31892 nor n31954 n31955 ; n31956
g31893 and n3457 n27442 ; n31957
g31894 and n3542 n26890 ; n31958
g31895 and n3606 n27173 ; n31959
g31896 nor n31958 n31959 ; n31960
g31897 and n31957_not n31960 ; n31961
g31898 and n3368_not n31961 ; n31962
g31899 and n27455_not n31961 ; n31963
g31900 nor n31962 n31963 ; n31964
g31901 and a[29] n31964_not ; n31965
g31902 and a[29]_not n31964 ; n31966
g31903 nor n31965 n31966 ; n31967
g31904 and n31956 n31967_not ; n31968
g31905 and n31956_not n31967 ; n31969
g31906 nor n31968 n31969 ; n31970
g31907 and n31921_not n31970 ; n31971
g31908 and n31921 n31970_not ; n31972
g31909 nor n31971 n31972 ; n31973
g31910 and n3884 n28208_not ; n31974
g31911 and n3967 n27698 ; n31975
g31912 and n4046 n27964 ; n31976
g31913 nor n31975 n31976 ; n31977
g31914 and n31974_not n31977 ; n31978
g31915 and n4050 n28223_not ; n31979
g31916 and n31978 n31979_not ; n31980
g31917 and a[26] n31980_not ; n31981
g31918 and a[26] n31981_not ; n31982
g31919 nor n31980 n31981 ; n31983
g31920 nor n31982 n31983 ; n31984
g31921 and n31973 n31984_not ; n31985
g31922 and n31973 n31985_not ; n31986
g31923 nor n31984 n31985 ; n31987
g31924 nor n31986 n31987 ; n31988
g31925 nor n31851 n31908 ; n31989
g31926 nor n31848 n31989 ; n31990
g31927 nor n31988 n31990 ; n31991
g31928 nor n31988 n31991 ; n31992
g31929 nor n31990 n31991 ; n31993
g31930 nor n31992 n31993 ; n31994
g31931 nor n31912 n31915 ; n31995
g31932 and n31994 n31995 ; n31996
g31933 nor n31994 n31995 ; n31997
g31934 nor n31996 n31997 ; n31998
g31935 and n31919_not n31998 ; n31999
g31936 and n31919 n31998_not ; n32000
g31937 or n31999 n32000 ; result[29]
g31938 and n31919 n31998 ; n32002
g31939 nor n31991 n31997 ; n32003
g31940 nor n31971 n31985 ; n32004
g31941 nor n31946 n31949 ; n32005
g31942 and n4009 n13075 ; n32006
g31943 and n3848 n32006 ; n32007
g31944 and n3839 n32007 ; n32008
g31945 and n2273 n32008 ; n32009
g31946 and n26016 n32009 ; n32010
g31947 and n3984 n32010 ; n32011
g31948 and n825_not n32011 ; n32012
g31949 and n31945_not n32012 ; n32013
g31950 and n31945 n32012_not ; n32014
g31951 nor n32005 n32014 ; n32015
g31952 and n32013_not n32015 ; n32016
g31953 nor n32005 n32016 ; n32017
g31954 nor n32014 n32016 ; n32018
g31955 and n32013_not n32018 ; n32019
g31956 nor n32017 n32019 ; n32020
g31957 and n75 n26904_not ; n32021
g31958 and n3020 n26890 ; n32022
g31959 and n3023 n26066 ; n32023
g31960 and n3028 n26060 ; n32024
g31961 nor n32023 n32024 ; n32025
g31962 and n32022_not n32025 ; n32026
g31963 and n32021_not n32026 ; n32027
g31964 nor n32020 n32027 ; n32028
g31965 nor n32020 n32028 ; n32029
g31966 nor n32027 n32028 ; n32030
g31967 nor n32029 n32030 ; n32031
g31968 nor n31955 n31968 ; n32032
g31969 and n32031 n32032 ; n32033
g31970 nor n32031 n32032 ; n32034
g31971 nor n32033 n32034 ; n32035
g31972 nor n25957 n28208 ; n32036
g31973 and n3967 n27964 ; n32037
g31974 nor n32036 n32037 ; n32038
g31975 and n4050 n28221_not ; n32039
g31976 and n32038 n32039_not ; n32040
g31977 and a[26] n32040_not ; n32041
g31978 nor n32040 n32041 ; n32042
g31979 and a[26] n32041_not ; n32043
g31980 nor n32042 n32043 ; n32044
g31981 and n3457 n27698 ; n32045
g31982 and n3542 n27173 ; n32046
g31983 and n3606 n27442 ; n32047
g31984 nor n32046 n32047 ; n32048
g31985 and n32045_not n32048 ; n32049
g31986 and n3368 n27713_not ; n32050
g31987 and n32049 n32050_not ; n32051
g31988 and a[29] n32051_not ; n32052
g31989 and a[29] n32052_not ; n32053
g31990 nor n32051 n32052 ; n32054
g31991 nor n32053 n32054 ; n32055
g31992 nor n32044 n32055 ; n32056
g31993 nor n32044 n32056 ; n32057
g31994 nor n32055 n32056 ; n32058
g31995 nor n32057 n32058 ; n32059
g31996 and n32035_not n32059 ; n32060
g31997 and n32035 n32059_not ; n32061
g31998 nor n32060 n32061 ; n32062
g31999 and n32004_not n32062 ; n32063
g32000 and n32004 n32062_not ; n32064
g32001 nor n32063 n32064 ; n32065
g32002 and n32003_not n32065 ; n32066
g32003 and n32003 n32065_not ; n32067
g32004 nor n32066 n32067 ; n32068
g32005 nor n32002 n32068 ; n32069
g32006 and n32002 n32068 ; n32070
g32007 nor n32069 n32070 ; result[30]
g32008 nor n32063 n32066 ; n32072
g32009 and n3457 n27964 ; n32073
g32010 and n3542 n27442 ; n32074
g32011 and n3606 n27698 ; n32075
g32012 nor n32074 n32075 ; n32076
g32013 and n32073_not n32076 ; n32077
g32014 and n3368 n27976 ; n32078
g32015 and n32077 n32078_not ; n32079
g32016 nor n32028 n32034 ; n32080
g32017 and a[29] n32080_not ; n32081
g32018 and a[29]_not n32080 ; n32082
g32019 nor n32081 n32082 ; n32083
g32020 and n32079 n32083 ; n32084
g32021 nor n32079 n32083 ; n32085
g32022 nor n32084 n32085 ; n32086
g32023 and n75 n27185 ; n32087
g32024 and n3020 n27173 ; n32088
g32025 and n3023 n26060 ; n32089
g32026 and n3028 n26890 ; n32090
g32027 nor n32089 n32090 ; n32091
g32028 and n32088_not n32091 ; n32092
g32029 and n32087_not n32092 ; n32093
g32030 and n32018 n32093_not ; n32094
g32031 and n32018_not n32093 ; n32095
g32032 nor n32094 n32095 ; n32096
g32033 and n32086 n32096_not ; n32097
g32034 and n32086_not n32096 ; n32098
g32035 nor n32097 n32098 ; n32099
g32036 nor n32056 n32061 ; n32100
g32037 and n3874 n4511 ; n32101
g32038 and n601_not n32101 ; n32102
g32039 and a[26] n32102_not ; n32103
g32040 and a[26]_not n32102 ; n32104
g32041 nor n32103 n32104 ; n32105
g32042 nor n26010 n28208 ; n32106
g32043 and n31945 n32106_not ; n32107
g32044 and n31945_not n32106 ; n32108
g32045 nor n32107 n32108 ; n32109
g32046 and n32105 n32109 ; n32110
g32047 nor n32105 n32109 ; n32111
g32048 nor n32110 n32111 ; n32112
g32049 and n32100 n32112_not ; n32113
g32050 and n32100_not n32112 ; n32114
g32051 nor n32113 n32114 ; n32115
g32052 and n32099 n32115 ; n32116
g32053 nor n32099 n32115 ; n32117
g32054 nor n32116 n32117 ; n32118
g32055 nor n32072 n32118 ; n32119
g32056 and n32072 n32118 ; n32120
g32057 nor n32119 n32120 ; n32121
g32058 and n32070 n32121 ; n32122
g32059 nor n32070 n32121 ; n32123
g32060 or n32122 n32123 ; result[31]
g32061 not n70 ; n70_not
g32062 not n81 ; n81_not
g32063 not n91 ; n91_not
g32064 not n74 ; n74_not
g32065 not n67 ; n67_not
g32066 not n86 ; n86_not
g32067 not n95 ; n95_not
g32068 not n99 ; n99_not
g32069 not n200 ; n200_not
g32070 not n201 ; n201_not
g32071 not n111 ; n111_not
g32072 not n102 ; n102_not
g32073 not n301 ; n301_not
g32074 not n400 ; n400_not
g32075 not n130 ; n130_not
g32076 not n121 ; n121_not
g32077 not n302 ; n302_not
g32078 not n203 ; n203_not
g32079 not n420 ; n420_not
g32080 not n231 ; n231_not
g32081 not n123 ; n123_not
g32082 not n240 ; n240_not
g32083 not n402 ; n402_not
g32084 not n222 ; n222_not
g32085 not n150 ; n150_not
g32086 not n330 ; n330_not
g32087 not n132 ; n132_not
g32088 not n232 ; n232_not
g32089 not n223 ; n223_not
g32090 not n304 ; n304_not
g32091 not n340 ; n340_not
g32092 not n115 ; n115_not
g32093 not n331 ; n331_not
g32094 not n601 ; n601_not
g32095 not n205 ; n205_not
g32096 not n151 ; n151_not
g32097 not n142 ; n142_not
g32098 not n430 ; n430_not
g32099 not n511 ; n511_not
g32100 not n403 ; n403_not
g32101 not n170 ; n170_not
g32102 not n206 ; n206_not
g32103 not n710 ; n710_not
g32104 not n107 ; n107_not
g32105 not n125 ; n125_not
g32106 not n251 ; n251_not
g32107 not n161 ; n161_not
g32108 not n620 ; n620_not
g32109 not n242 ; n242_not
g32110 not n602 ; n602_not
g32111 not n233 ; n233_not
g32112 not n422 ; n422_not
g32113 not n332 ; n332_not
g32114 not n224 ; n224_not
g32115 not n305 ; n305_not
g32116 not n152 ; n152_not
g32117 not n513 ; n513_not
g32118 not n306 ; n306_not
g32119 not n531 ; n531_not
g32120 not n603 ; n603_not
g32121 not n270 ; n270_not
g32122 not n252 ; n252_not
g32123 not n144 ; n144_not
g32124 not n243 ; n243_not
g32125 not n225 ; n225_not
g32126 not n135 ; n135_not
g32127 not n171 ; n171_not
g32128 not n504 ; n504_not
g32129 not n352 ; n352_not
g32130 not n712 ; n712_not
g32131 not n532 ; n532_not
g32132 not n514 ; n514_not
g32133 not n271 ; n271_not
g32134 not n325 ; n325_not
g32135 not n334 ; n334_not
g32136 not n451 ; n451_not
g32137 not n280 ; n280_not
g32138 not n424 ; n424_not
g32139 not n460 ; n460_not
g32140 not n505 ; n505_not
g32141 not n145 ; n145_not
g32142 not n136 ; n136_not
g32143 not n226 ; n226_not
g32144 not n127 ; n127_not
g32145 not n190 ; n190_not
g32146 not n163 ; n163_not
g32147 not n118 ; n118_not
g32148 not n154 ; n154_not
g32149 not n326 ; n326_not
g32150 not n155 ; n155_not
g32151 not n452 ; n452_not
g32152 not n416 ; n416_not
g32153 not n371 ; n371_not
g32154 not n254 ; n254_not
g32155 not n245 ; n245_not
g32156 not n164 ; n164_not
g32157 not n173 ; n173_not
g32158 not n623 ; n623_not
g32159 not n191 ; n191_not
g32160 not n290 ; n290_not
g32161 not n353 ; n353_not
g32162 not n272 ; n272_not
g32163 not n461 ; n461_not
g32164 not n146 ; n146_not
g32165 not n335 ; n335_not
g32166 not n506 ; n506_not
g32167 not n803 ; n803_not
g32168 not n236 ; n236_not
g32169 not n281 ; n281_not
g32170 not n641 ; n641_not
g32171 not n713 ; n713_not
g32172 not n425 ; n425_not
g32173 not n119 ; n119_not
g32174 not n470 ; n470_not
g32175 not n327 ; n327_not
g32176 not n228 ; n228_not
g32177 not n372 ; n372_not
g32178 not n462 ; n462_not
g32179 not n354 ; n354_not
g32180 not n633 ; n633_not
g32181 not n525 ; n525_not
g32182 not n165 ; n165_not
g32183 not n273 ; n273_not
g32184 not n192 ; n192_not
g32185 not n417 ; n417_not
g32186 not n453 ; n453_not
g32187 not n435 ; n435_not
g32188 not n255 ; n255_not
g32189 not n363 ; n363_not
g32190 not n246 ; n246_not
g32191 not n426 ; n426_not
g32192 not n714 ; n714_not
g32193 not n237 ; n237_not
g32194 not n147 ; n147_not
g32195 not n328 ; n328_not
g32196 not n355 ; n355_not
g32197 not n427 ; n427_not
g32198 not n274 ; n274_not
g32199 not n562 ; n562_not
g32200 not n571 ; n571_not
g32201 not n490 ; n490_not
g32202 not n715 ; n715_not
g32203 not n292 ; n292_not
g32204 not n283 ; n283_not
g32205 not n157 ; n157_not
g32206 not n436 ; n436_not
g32207 not n337 ; n337_not
g32208 not n364 ; n364_not
g32209 not n229 ; n229_not
g32210 not n175 ; n175_not
g32211 not n248 ; n248_not
g32212 not n275 ; n275_not
g32213 not n716 ; n716_not
g32214 not n392 ; n392_not
g32215 not n518 ; n518_not
g32216 not n167 ; n167_not
g32217 not n338 ; n338_not
g32218 not n419 ; n419_not
g32219 not n329 ; n329_not
g32220 not n509 ; n509_not
g32221 not n194 ; n194_not
g32222 not n293 ; n293_not
g32223 not n428 ; n428_not
g32224 not n158 ; n158_not
g32225 not n563 ; n563_not
g32226 not n617 ; n617_not
g32227 not n239 ; n239_not
g32228 not n527 ; n527_not
g32229 not n284 ; n284_not
g32230 not n752 ; n752_not
g32231 not n374 ; n374_not
g32232 not n536 ; n536_not
g32233 not n149 ; n149_not
g32234 not n932 ; n932_not
g32235 not n825 ; n825_not
g32236 not n519 ; n519_not
g32237 not n357 ; n357_not
g32238 not n375 ; n375_not
g32239 not n393 ; n393_not
g32240 not n249 ; n249_not
g32241 not n339 ; n339_not
g32242 not n474 ; n474_not
g32243 not n771 ; n771_not
g32244 not n429 ; n429_not
g32245 not n492 ; n492_not
g32246 not n564 ; n564_not
g32247 not n537 ; n537_not
g32248 not n168 ; n168_not
g32249 not n672 ; n672_not
g32250 not n366 ; n366_not
g32251 not n276 ; n276_not
g32252 not n438 ; n438_not
g32253 not n177 ; n177_not
g32254 not n493 ; n493_not
g32255 not n295 ; n295_not
g32256 not n637 ; n637_not
g32257 not n367 ; n367_not
g32258 not n358 ; n358_not
g32259 not n655 ; n655_not
g32260 not n394 ; n394_not
g32261 not n286 ; n286_not
g32262 not n619 ; n619_not
g32263 not n961 ; n961_not
g32264 not n277 ; n277_not
g32265 not n592 ; n592_not
g32266 not n169 ; n169_not
g32267 not n673 ; n673_not
g32268 not n466 ; n466_not
g32269 not n557 ; n557_not
g32270 not n791 ; n791_not
g32271 not n368 ; n368_not
g32272 not n809 ; n809_not
g32273 not n287 ; n287_not
g32274 not n278 ; n278_not
g32275 not n449 ; n449_not
g32276 not n296 ; n296_not
g32277 not n980 ; n980_not
g32278 not n746 ; n746_not
g32279 not n188 ; n188_not
g32280 not n656 ; n656_not
g32281 not n395 ; n395_not
g32282 not n468 ; n468_not
g32283 not n594 ; n594_not
g32284 not n396 ; n396_not
g32285 not n639 ; n639_not
g32286 not n189 ; n189_not
g32287 not n657 ; n657_not
g32288 not n567 ; n567_not
g32289 not n558 ; n558_not
g32290 not n495 ; n495_not
g32291 not n666 ; n666_not
g32292 not n289 ; n289_not
g32293 not n397 ; n397_not
g32294 not n847 ; n847_not
g32295 not n298 ; n298_not
g32296 not n667 ; n667_not
g32297 not n496 ; n496_not
g32298 not n568 ; n568_not
g32299 not n469 ; n469_not
g32300 not n883 ; n883_not
g32301 not n398 ; n398_not
g32302 not n587 ; n587_not
g32303 not n299 ; n299_not
g32304 not n875 ; n875_not
g32305 not n569 ; n569_not
g32306 not n884 ; n884_not
g32307 not n777 ; n777_not
g32308 not n867 ; n867_not
g32309 not n489 ; n489_not
g32310 not n958 ; n958_not
g32311 not n589 ; n589_not
g32312 not n886 ; n886_not
g32313 not n689 ; n689_not
g32314 not n1010 ; n1010_not
g32315 not n1011 ; n1011_not
g32316 not n1101 ; n1101_not
g32317 not n1102 ; n1102_not
g32318 not n3012 ; n3012_not
g32319 not n1203 ; n1203_not
g32320 not n1104 ; n1104_not
g32321 not n4200 ; n4200_not
g32322 not n3021 ; n3021_not
g32323 not n1060 ; n1060_not
g32324 not n4201 ; n4201_not
g32325 not n7000 ; n7000_not
g32326 not n4121 ; n4121_not
g32327 not n5111 ; n5111_not
g32328 not n3032 ; n3032_not
g32329 not n4050 ; n4050_not
g32330 not n5121 ; n5121_not
g32331 not n1062 ; n1062_not
g32332 not n3015 ; n3015_not
g32333 not n6120 ; n6120_not
g32334 not n9000 ; n9000_not
g32335 not n6003 ; n6003_not
g32336 not n7200 ; n7200_not
g32337 not n6210 ; n6210_not
g32338 not n6300 ; n6300_not
g32339 not n1072 ; n1072_not
g32340 not n5410 ; n5410_not
g32341 not n2152 ; n2152_not
g32342 not n6004 ; n6004_not
g32343 not n3241 ; n3241_not
g32344 not n1306 ; n1306_not
g32345 not n9001 ; n9001_not
g32346 not n6400 ; n6400_not
g32347 not n4204 ; n4204_not
g32348 not n3331 ; n3331_not
g32349 not n7102 ; n7102_not
g32350 not n7210 ; n7210_not
g32351 not n1235 ; n1235_not
g32352 not n6122 ; n6122_not
g32353 not n2900 ; n2900_not
g32354 not n1127 ; n1127_not
g32355 not n5510 ; n5510_not
g32356 not n6041 ; n6041_not
g32357 not n5330 ; n5330_not
g32358 not n5114 ; n5114_not
g32359 not n6140 ; n6140_not
g32360 not n5411 ; n5411_not
g32361 not n5600 ; n5600_not
g32362 not n4700 ; n4700_not
g32363 not n4520 ; n4520_not
g32364 not n7022 ; n7022_not
g32365 not n7211 ; n7211_not
g32366 not n3332 ; n3332_not
g32367 not n7310 ; n7310_not
g32368 not n4610 ; n4610_not
g32369 not n7112 ; n7112_not
g32370 not n4430 ; n4430_not
g32371 not n4601 ; n4601_not
g32372 not n4061 ; n4061_not
g32373 not n4070 ; n4070_not
g32374 not n7040 ; n7040_not
g32375 not n5420 ; n5420_not
g32376 not n5124 ; n5124_not
g32377 not n5115 ; n5115_not
g32378 not n9201 ; n9201_not
g32379 not n5502 ; n5502_not
g32380 not n9210 ; n9210_not
g32381 not n3540 ; n3540_not
g32382 not n6222 ; n6222_not
g32383 not n4053 ; n4053_not
g32384 not n3702 ; n3702_not
g32385 not n3018 ; n3018_not
g32386 not n3621 ; n3621_not
g32387 not n9120 ; n9120_not
g32388 not n7131 ; n7131_not
g32389 not n7122 ; n7122_not
g32390 not n9021 ; n9021_not
g32391 not n7410 ; n7410_not
g32392 not n6240 ; n6240_not
g32393 not n6303 ; n6303_not
g32394 not n3333 ; n3333_not
g32395 not n7221 ; n7221_not
g32396 not n2910 ; n2910_not
g32397 not n4701 ; n4701_not
g32398 not n4431 ; n4431_not
g32399 not n8400 ; n8400_not
g32400 not n8013 ; n8013_not
g32401 not n8004 ; n8004_not
g32402 not n4611 ; n4611_not
g32403 not n5322 ; n5322_not
g32404 not n7113 ; n7113_not
g32405 not n6123 ; n6123_not
g32406 not n6150 ; n6150_not
g32407 not n6402 ; n6402_not
g32408 not n9102 ; n9102_not
g32409 not n3027 ; n3027_not
g32410 not n8310 ; n8310_not
g32411 not n7500 ; n7500_not
g32412 not n6204 ; n6204_not
g32413 not n5412 ; n5412_not
g32414 not n7041 ; n7041_not
g32415 not n3711 ; n3711_not
g32416 not n7140 ; n7140_not
g32417 not n7060 ; n7060_not
g32418 not n5116 ; n5116_not
g32419 not n2533 ; n2533_not
g32420 not n7222 ; n7222_not
g32421 not n4045 ; n4045_not
g32422 not n9130 ; n9130_not
g32423 not n6007 ; n6007_not
g32424 not n5170 ; n5170_not
g32425 not n5053 ; n5053_not
g32426 not n4531 ; n4531_not
g32427 not n7150 ; n7150_not
g32428 not n3361 ; n3361_not
g32429 not n4351 ; n4351_not
g32430 not n9202 ; n9202_not
g32431 not n6322 ; n6322_not
g32432 not n1246 ; n1246_not
g32433 not n9013 ; n9013_not
g32434 not n3613 ; n3613_not
g32435 not n9220 ; n9220_not
g32436 not n7015 ; n7015_not
g32437 not n8212 ; n8212_not
g32438 not n9400 ; n9400_not
g32439 not n3820 ; n3820_not
g32440 not n8410 ; n8410_not
g32441 not n4180 ; n4180_not
g32442 not n8401 ; n8401_not
g32443 not n5530 ; n5530_not
g32444 not n8302 ; n8302_not
g32445 not n5503 ; n5503_not
g32446 not n6124 ; n6124_not
g32447 not n5431 ; n5431_not
g32448 not n6043 ; n6043_not
g32449 not n8014 ; n8014_not
g32450 not n6241 ; n6241_not
g32451 not n8050 ; n8050_not
g32452 not n6205 ; n6205_not
g32453 not n3712 ; n3712_not
g32454 not n3703 ; n3703_not
g32455 not n8140 ; n8140_not
g32456 not n8122 ; n8122_not
g32457 not n8104 ; n8104_not
g32458 not n6223 ; n6223_not
g32459 not n5701 ; n5701_not
g32460 not n5350 ; n5350_not
g32461 not n2902 ; n2902_not
g32462 not n4630 ; n4630_not
g32463 not n9040 ; n9040_not
g32464 not n4423 ; n4423_not
g32465 not n3019 ; n3019_not
g32466 not n4702 ; n4702_not
g32467 not n4612 ; n4612_not
g32468 not n7303 ; n7303_not
g32469 not n5602 ; n5602_not
g32470 not n5611 ; n5611_not
g32471 not n3244 ; n3244_not
g32472 not n7240 ; n7240_not
g32473 not n2920 ; n2920_not
g32474 not n4450 ; n4450_not
g32475 not n7511 ; n7511_not
g32476 not n1472 ; n1472_not
g32477 not n5540 ; n5540_not
g32478 not n2057 ; n2057_not
g32479 not n1364 ; n1364_not
g32480 not n2291 ; n2291_not
g32481 not n1913 ; n1913_not
g32482 not n6206 ; n6206_not
g32483 not n8204 ; n8204_not
g32484 not n3605 ; n3605_not
g32485 not n8123 ; n8123_not
g32486 not n8105 ; n8105_not
g32487 not n4730 ; n4730_not
g32488 not n6224 ; n6224_not
g32489 not n5360 ; n5360_not
g32490 not n7034 ; n7034_not
g32491 not n2840 ; n2840_not
g32492 not n3083 ; n3083_not
g32493 not n8141 ; n8141_not
g32494 not n4622 ; n4622_not
g32495 not n4073 ; n4073_not
g32496 not n7421 ; n7421_not
g32497 not n6422 ; n6422_not
g32498 not n8402 ; n8402_not
g32499 not n4064 ; n4064_not
g32500 not n7403 ; n7403_not
g32501 not n3146 ; n3146_not
g32502 not n2912 ; n2912_not
g32503 not n8231 ; n8231_not
g32504 not n7007 ; n7007_not
g32505 not n3812 ; n3812_not
g32506 not n5432 ; n5432_not
g32507 not n9410 ; n9410_not
g32508 not n6143 ; n6143_not
g32509 not n4181 ; n4181_not
g32510 not n5504 ; n5504_not
g32511 not n5450 ; n5450_not
g32512 not n6413 ; n6413_not
g32513 not n5135 ; n5135_not
g32514 not n9140 ; n9140_not
g32515 not n6431 ; n6431_not
g32516 not n9203 ; n9203_not
g32517 not n9050 ; n9050_not
g32518 not n6332 ; n6332_not
g32519 not n8321 ; n8321_not
g32520 not n4055 ; n4055_not
g32521 not n7205 ; n7205_not
g32522 not n7223 ; n7223_not
g32523 not n7250 ; n7250_not
g32524 not n5108 ; n5108_not
g32525 not n7043 ; n7043_not
g32526 not n7241 ; n7241_not
g32527 not n9014 ; n9014_not
g32528 not n8015 ; n8015_not
g32529 not n3632 ; n3632_not
g32530 not n4451 ; n4451_not
g32531 not n7070 ; n7070_not
g32532 not n5342 ; n5342_not
g32533 not n8051 ; n8051_not
g32534 not n8501 ; n8501_not
g32535 not n7133 ; n7133_not
g32536 not n9302 ; n9302_not
g32537 not n7115 ; n7115_not
g32538 not n9320 ; n9320_not
g32539 not n5612 ; n5612_not
g32540 not n9141 ; n9141_not
g32541 not n9222 ; n9222_not
g32542 not n2571 ; n2571_not
g32543 not n9321 ; n9321_not
g32544 not n9105 ; n9105_not
g32545 not n9024 ; n9024_not
g32546 not n9303 ; n9303_not
g32547 not n9231 ; n9231_not
g32548 not n1572 ; n1572_not
g32549 not n5541 ; n5541_not
g32550 not n4515 ; n4515_not
g32551 not n9123 ; n9123_not
g32552 not n8421 ; n8421_not
g32553 not n8502 ; n8502_not
g32554 not n4902 ; n4902_not
g32555 not n4533 ; n4533_not
g32556 not n4173 ; n4173_not
g32557 not n4074 ; n4074_not
g32558 not n3615 ; n3615_not
g32559 not n3624 ; n3624_not
g32560 not n3354 ; n3354_not
g32561 not n2922 ; n2922_not
g32562 not n3327 ; n3327_not
g32563 not n2904 ; n2904_not
g32564 not n2832 ; n2832_not
g32565 not n4560 ; n4560_not
g32566 not n4551 ; n4551_not
g32567 not n4470 ; n4470_not
g32568 not n4461 ; n4461_not
g32569 not n4443 ; n4443_not
g32570 not n5415 ; n5415_not
g32571 not n9600 ; n9600_not
g32572 not n9240 ; n9240_not
g32573 not n9411 ; n9411_not
g32574 not n5451 ; n5451_not
g32575 not n5442 ; n5442_not
g32576 not n5136 ; n5136_not
g32577 not n5325 ; n5325_not
g32578 not n8241 ; n8241_not
g32579 not n8250 ; n8250_not
g32580 not n8070 ; n8070_not
g32581 not n5712 ; n5712_not
g32582 not n7170 ; n7170_not
g32583 not n5640 ; n5640_not
g32584 not n7260 ; n7260_not
g32585 not n8142 ; n8142_not
g32586 not n7107 ; n7107_not
g32587 not n8160 ; n8160_not
g32588 not n8205 ; n8205_not
g32589 not n5622 ; n5622_not
g32590 not n7071 ; n7071_not
g32591 not n8304 ; n8304_not
g32592 not n8124 ; n8124_not
g32593 not n8106 ; n8106_not
g32594 not n7035 ; n7035_not
g32595 not n7503 ; n7503_not
g32596 not n6342 ; n6342_not
g32597 not n6315 ; n6315_not
g32598 not n6234 ; n6234_not
g32599 not n7602 ; n7602_not
g32600 not n5613 ; n5613_not
g32601 not n6144 ; n6144_not
g32602 not n7512 ; n7512_not
g32603 not n8034 ; n8034_not
g32604 not n8610 ; n8610_not
g32605 not n7206 ; n7206_not
g32606 not n2850 ; n2850_not
g32607 not n6153 ; n6153_not
g32608 not n6333 ; n6333_not
g32609 not n7620 ; n7620_not
g32610 not n6432 ; n6432_not
g32611 not n8052 ; n8052_not
g32612 not n8430 ; n8430_not
g32613 not n4633 ; n4633_not
g32614 not n3715 ; n3715_not
g32615 not n2464 ; n2464_not
g32616 not n7810 ; n7810_not
g32617 not n6541 ; n6541_not
g32618 not n3805 ; n3805_not
g32619 not n7711 ; n7711_not
g32620 not n7603 ; n7603_not
g32621 not n7531 ; n7531_not
g32622 not n8341 ; n8341_not
g32623 not n9610 ; n9610_not
g32624 not n8026 ; n8026_not
g32625 not n8413 ; n8413_not
g32626 not n9421 ; n9421_not
g32627 not n9322 ; n9322_not
g32628 not n9304 ; n9304_not
g32629 not n9232 ; n9232_not
g32630 not n8512 ; n8512_not
g32631 not n9142 ; n9142_not
g32632 not n9133 ; n9133_not
g32633 not n4084 ; n4084_not
g32634 not n5335 ; n5335_not
g32635 not n5362 ; n5362_not
g32636 not n8206 ; n8206_not
g32637 not n5416 ; n5416_not
g32638 not n5344 ; n5344_not
g32639 not n5128 ; n5128_not
g32640 not n8260 ; n8260_not
g32641 not n2842 ; n2842_not
g32642 not n3364 ; n3364_not
g32643 not n5254 ; n5254_not
g32644 not n6901 ; n6901_not
g32645 not n4057 ; n4057_not
g32646 not n5650 ; n5650_not
g32647 not n2914 ; n2914_not
g32648 not n7036 ; n7036_not
g32649 not n7054 ; n7054_not
g32650 not n7072 ; n7072_not
g32651 not n4426 ; n4426_not
g32652 not n7135 ; n7135_not
g32653 not n8017 ; n8017_not
g32654 not n7090 ; n7090_not
g32655 not n7108 ; n7108_not
g32656 not n6118 ; n6118_not
g32657 not n6145 ; n6145_not
g32658 not n6190 ; n6190_not
g32659 not n6217 ; n6217_not
g32660 not n6244 ; n6244_not
g32661 not n6280 ; n6280_not
g32662 not n6334 ; n6334_not
g32663 not n6352 ; n6352_not
g32664 not n6370 ; n6370_not
g32665 not n6406 ; n6406_not
g32666 not n6433 ; n6433_not
g32667 not n2860 ; n2860_not
g32668 not n5902 ; n5902_not
g32669 not n7261 ; n7261_not
g32670 not n4705 ; n4705_not
g32671 not n4741 ; n4741_not
g32672 not n4912 ; n4912_not
g32673 not n4930 ; n4930_not
g32674 not n4903 ; n4903_not
g32675 not n7513 ; n7513_not
g32676 not n7504 ; n7504_not
g32677 not n4471 ; n4471_not
g32678 not n4480 ; n4480_not
g32679 not n4516 ; n4516_not
g32680 not n7153 ; n7153_not
g32681 not n4570 ; n4570_not
g32682 not n7207 ; n7207_not
g32683 not n7216 ; n7216_not
g32684 not n7234 ; n7234_not
g32685 not n4525 ; n4525_not
g32686 not n5632 ; n5632_not
g32687 not n4615 ; n4615_not
g32688 not n7306 ; n7306_not
g32689 not n7324 ; n7324_not
g32690 not n8530 ; n8530_not
g32691 not n8620 ; n8620_not
g32692 not n8800 ; n8800_not
g32693 not n3329 ; n3329_not
g32694 not n5507 ; n5507_not
g32695 not n7307 ; n7307_not
g32696 not n1178 ; n1178_not
g32697 not n8405 ; n8405_not
g32698 not n4706 ; n4706_not
g32699 not n4085 ; n4085_not
g32700 not n5471 ; n5471_not
g32701 not n8153 ; n8153_not
g32702 not n8423 ; n8423_not
g32703 not n2852 ; n2852_not
g32704 not n8135 ; n8135_not
g32705 not n4715 ; n4715_not
g32706 not n2924 ; n2924_not
g32707 not n8540 ; n8540_not
g32708 not n9332 ; n9332_not
g32709 not n6272 ; n6272_not
g32710 not n7541 ; n7541_not
g32711 not n7550 ; n7550_not
g32712 not n8180 ; n8180_not
g32713 not n5534 ; n5534_not
g32714 not n6245 ; n6245_not
g32715 not n5561 ; n5561_not
g32716 not n8603 ; n8603_not
g32717 not n6416 ; n6416_not
g32718 not n9530 ; n9530_not
g32719 not n3347 ; n3347_not
g32720 not n6353 ; n6353_not
g32721 not n9512 ; n9512_not
g32722 not n3815 ; n3815_not
g32723 not n9080 ; n9080_not
g32724 not n4067 ; n4067_not
g32725 not n8027 ; n8027_not
g32726 not n2834 ; n2834_not
g32727 not n3806 ; n3806_not
g32728 not n5651 ; n5651_not
g32729 not n2870 ; n2870_not
g32730 not n5831 ; n5831_not
g32731 not n8063 ; n8063_not
g32732 not n8045 ; n8045_not
g32733 not n8720 ; n8720_not
g32734 not n3617 ; n3617_not
g32735 not n8351 ; n8351_not
g32736 not n5633 ; n5633_not
g32737 not n4940 ; n4940_not
g32738 not n9701 ; n9701_not
g32739 not n6911 ; n6911_not
g32740 not n4922 ; n4922_not
g32741 not n4445 ; n4445_not
g32742 not n9035 ; n9035_not
g32743 not n8117 ; n8117_not
g32744 not n5372 ; n5372_not
g32745 not n5930 ; n5930_not
g32746 not n4904 ; n4904_not
g32747 not n8621 ; n8621_not
g32748 not n3248 ; n3248_not
g32749 not n5912 ; n5912_not
g32750 not n4850 ; n4850_not
g32751 not n8081 ; n8081_not
g32752 not n6803 ; n6803_not
g32753 not n6227 ; n6227_not
g32754 not n5606 ; n5606_not
g32755 not n7109 ; n7109_not
g32756 not n6254 ; n6254_not
g32757 not n6074 ; n6074_not
g32758 not n9206 ; n9206_not
g32759 not n4571 ; n4571_not
g32760 not n4436 ; n4436_not
g32761 not n7613 ; n7613_not
g32762 not n7091 ; n7091_not
g32763 not n9233 ; n9233_not
g32764 not n9062 ; n9062_not
g32765 not n7163 ; n7163_not
g32766 not n7802 ; n7802_not
g32767 not n7145 ; n7145_not
g32768 not n5444 ; n5444_not
g32769 not n9116 ; n9116_not
g32770 not n7721 ; n7721_not
g32771 not n9053 ; n9053_not
g32772 not n8270 ; n8270_not
g32773 not n6209 ; n6209_not
g32774 not n4463 ; n4463_not
g32775 not n4193 ; n4193_not
g32776 not n9260 ; n9260_not
g32777 not n7604 ; n7604_not
g32778 not n5480 ; n5480_not
g32779 not n6308 ; n6308_not
g32780 not n7226 ; n7226_not
g32781 not n9134 ; n9134_not
g32782 not n8801 ; n8801_not
g32783 not n2906 ; n2906_not
g32784 not n7055 ; n7055_not
g32785 not n7244 ; n7244_not
g32786 not n3456 ; n3456_not
g32787 not n4059 ; n4059_not
g32788 not n8226 ; n8226_not
g32789 not n7380 ; n7380_not
g32790 not n2736 ; n2736_not
g32791 not n8406 ; n8406_not
g32792 not n9045 ; n9045_not
g32793 not n7173 ; n7173_not
g32794 not n1665 ; n1665_not
g32795 not n4266 ; n4266_not
g32796 not n8271 ; n8271_not
g32797 not n6813 ; n6813_not
g32798 not n8460 ; n8460_not
g32799 not n4077 ; n4077_not
g32800 not n4536 ; n4536_not
g32801 not n4545 ; n4545_not
g32802 not n7056 ; n7056_not
g32803 not n9063 ; n9063_not
g32804 not n8550 ; n8550_not
g32805 not n7146 ; n7146_not
g32806 not n5508 ; n5508_not
g32807 not n9621 ; n9621_not
g32808 not n9081 ; n9081_not
g32809 not n8244 ; n8244_not
g32810 not n5616 ; n5616_not
g32811 not n7065 ; n7065_not
g32812 not n5472 ; n5472_not
g32813 not n9711 ; n9711_not
g32814 not n7317 ; n7317_not
g32815 not n5328 ; n5328_not
g32816 not n4572 ; n4572_not
g32817 not n9504 ; n9504_not
g32818 not n3708 ; n3708_not
g32819 not n4176 ; n4176_not
g32820 not n4086 ; n4086_not
g32821 not n7092 ; n7092_not
g32822 not n6930 ; n6930_not
g32823 not n3357 ; n3357_not
g32824 not n5661 ; n5661_not
g32825 not n5490 ; n5490_not
g32826 not n7029 ; n7029_not
g32827 not n7227 ; n7227_not
g32828 not n8172 ; n8172_not
g32829 not n7344 ; n7344_not
g32830 not n7245 ; n7245_not
g32831 not n5139 ; n5139_not
g32832 not n8622 ; n8622_not
g32833 not n5454 ; n5454_not
g32834 not n4068 ; n4068_not
g32835 not n5382 ; n5382_not
g32836 not n4644 ; n4644_not
g32837 not n4563 ; n4563_not
g32838 not n6912 ; n6912_not
g32839 not n6840 ; n6840_not
g32840 not n9342 ; n9342_not
g32841 not n6363 ; n6363_not
g32842 not n9315 ; n9315_not
g32843 not n6327 ; n6327_not
g32844 not n2844 ; n2844_not
g32845 not n8433 ; n8433_not
g32846 not n7911 ; n7911_not
g32847 not n8370 ; n8370_not
g32848 not n7722 ; n7722_not
g32849 not n2862 ; n2862_not
g32850 not n6462 ; n6462_not
g32851 not n6336 ; n6336_not
g32852 not n7506 ; n7506_not
g32853 not n5544 ; n5544_not
g32854 not n6372 ; n6372_not
g32855 not n6426 ; n6426_not
g32856 not n6417 ; n6417_not
g32857 not n6183 ; n6183_not
g32858 not n9162 ; n9162_not
g32859 not n6165 ; n6165_not
g32860 not n7803 ; n7803_not
g32861 not n9135 ; n9135_not
g32862 not n6138 ; n6138_not
g32863 not n7623 ; n7623_not
g32864 not n6273 ; n6273_not
g32865 not n6228 ; n6228_not
g32866 not n9207 ; n9207_not
g32867 not n8505 ; n8505_not
g32868 not n5517 ; n5517_not
g32869 not n9180 ; n9180_not
g32870 not n7533 ; n7533_not
g32871 not n7704 ; n7704_not
g32872 not n7470 ; n7470_not
g32873 not n3348 ; n3348_not
g32874 not n6642 ; n6642_not
g32875 not n3627 ; n3627_not
g32876 not n4617 ; n4617_not
g32877 not n4671 ; n4671_not
g32878 not n8037 ; n8037_not
g32879 not n5841 ; n5841_not
g32880 not n9540 ; n9540_not
g32881 not n5913 ; n5913_not
g32882 not n4950 ; n4950_not
g32883 not n4923 ; n4923_not
g32884 not n2880 ; n2880_not
g32885 not n2916 ; n2916_not
g32886 not n8910 ; n8910_not
g32887 not n9414 ; n9414_not
g32888 not n7920 ; n7920_not
g32889 not n2674 ; n2674_not
g32890 not n4906 ; n4906_not
g32891 not n4609 ; n4609_not
g32892 not n4708 ; n4708_not
g32893 not n4429 ; n4429_not
g32894 not n7426 ; n7426_not
g32895 not n7750 ; n7750_not
g32896 not n2890 ; n2890_not
g32897 not n7129 ; n7129_not
g32898 not n7444 ; n7444_not
g32899 not n7624 ; n7624_not
g32900 not n7390 ; n7390_not
g32901 not n7408 ; n7408_not
g32902 not n7921 ; n7921_not
g32903 not n8551 ; n8551_not
g32904 not n4726 ; n4726_not
g32905 not n4861 ; n4861_not
g32906 not n7732 ; n7732_not
g32907 not n4717 ; n4717_not
g32908 not n5851 ; n5851_not
g32909 not n7804 ; n7804_not
g32910 not n5329 ; n5329_not
g32911 not n8236 ; n8236_not
g32912 not n4519 ; n4519_not
g32913 not n7840 ; n7840_not
g32914 not n4672 ; n4672_not
g32915 not n7327 ; n7327_not
g32916 not n7273 ; n7273_not
g32917 not n4663 ; n4663_not
g32918 not n7561 ; n7561_not
g32919 not n7255 ; n7255_not
g32920 not n4564 ; n4564_not
g32921 not n4654 ; n4654_not
g32922 not n7543 ; n7543_not
g32923 not n9028 ; n9028_not
g32924 not n7480 ; n7480_not
g32925 not n7462 ; n7462_not
g32926 not n8173 ; n8173_not
g32927 not n8911 ; n8911_not
g32928 not n7831 ; n7831_not
g32929 not n4528 ; n4528_not
g32930 not n8209 ; n8209_not
g32931 not n5383 ; n5383_not
g32932 not n4645 ; n4645_not
g32933 not n7336 ; n7336_not
g32934 not n9046 ; n9046_not
g32935 not n2836 ; n2836_not
g32936 not n7651 ; n7651_not
g32937 not n9208 ; n9208_not
g32938 not n8308 ; n8308_not
g32939 not n6076 ; n6076_not
g32940 not n4069 ; n4069_not
g32941 not n6454 ; n6454_not
g32942 not n6436 ; n6436_not
g32943 not n5491 ; n5491_not
g32944 not n9712 ; n9712_not
g32945 not n6940 ; n6940_not
g32946 not n8470 ; n8470_not
g32947 not n4078 ; n4078_not
g32948 not n3619 ; n3619_not
g32949 not n7039 ; n7039_not
g32950 not n8353 ; n8353_not
g32951 not n9244 ; n9244_not
g32952 not n8290 ; n8290_not
g32953 not n6328 ; n6328_not
g32954 not n8533 ; n8533_not
g32955 not n6292 ; n6292_not
g32956 not n9307 ; n9307_not
g32957 not n9325 ; n9325_not
g32958 not n4186 ; n4186_not
g32959 not n8416 ; n8416_not
g32960 not n6364 ; n6364_not
g32961 not n9352 ; n9352_not
g32962 not n4087 ; n4087_not
g32963 not n9262 ; n9262_not
g32964 not n8713 ; n8713_not
g32965 not n5338 ; n5338_not
g32966 not n5617 ; n5617_not
g32967 not n9550 ; n9550_not
g32968 not n9082 ; n9082_not
g32969 not n3367 ; n3367_not
g32970 not n4933 ; n4933_not
g32971 not n6643 ; n6643_not
g32972 not n8731 ; n8731_not
g32973 not n9640 ; n9640_not
g32974 not n5572 ; n5572_not
g32975 not n2872 ; n2872_not
g32976 not n9424 ; n9424_not
g32977 not n6157 ; n6157_not
g32978 not n2908 ; n2908_not
g32979 not n9442 ; n9442_not
g32980 not n6841 ; n6841_not
g32981 not n3880 ; n3880_not
g32982 not n5923 ; n5923_not
g32983 not n8380 ; n8380_not
g32984 not n8704 ; n8704_not
g32985 not n2926 ; n2926_not
g32986 not n3349 ; n3349_not
g32987 not n9505 ; n9505_not
g32988 not n6283 ; n6283_not
g32989 not n9343 ; n9343_not
g32990 not n6193 ; n6193_not
g32991 not n7075 ; n7075_not
g32992 not n9217 ; n9217_not
g32993 not n8812 ; n8812_not
g32994 not n9145 ; n9145_not
g32995 not n8272 ; n8272_not
g32996 not n9064 ; n9064_not
g32997 not n5464 ; n5464_not
g32998 not n5932 ; n5932_not
g32999 not n6247 ; n6247_not
g33000 not n8281 ; n8281_not
g33001 not n8515 ; n8515_not
g33002 not n9109 ; n9109_not
g33003 not n7291 ; n7291_not
g33004 not n2854 ; n2854_not
g33005 not n9226 ; n9226_not
g33006 not n9172 ; n9172_not
g33007 not n8632 ; n8632_not
g33008 not n7147 ; n7147_not
g33009 not n3368 ; n3368_not
g33010 not n5942 ; n5942_not
g33011 not n9452 ; n9452_not
g33012 not n3539 ; n3539_not
g33013 not n2189 ; n2189_not
g33014 not n5591 ; n5591_not
g33015 not n2882 ; n2882_not
g33016 not n5690 ; n5690_not
g33017 not n5663 ; n5663_not
g33018 not n9155 ; n9155_not
g33019 not n8381 ; n8381_not
g33020 not n4862 ; n4862_not
g33021 not n7490 ; n7490_not
g33022 not n2846 ; n2846_not
g33023 not n5924 ; n5924_not
g33024 not n8660 ; n8660_not
g33025 not n4727 ; n4727_not
g33026 not n7409 ; n7409_not
g33027 not n9551 ; n9551_not
g33028 not n7760 ; n7760_not
g33029 not n7427 ; n7427_not
g33030 not n4439 ; n4439_not
g33031 not n9533 ; n9533_not
g33032 not n7445 ; n7445_not
g33033 not n5852 ; n5852_not
g33034 not n4844 ; n4844_not
g33035 not n7463 ; n7463_not
g33036 not n9119 ; n9119_not
g33037 not n9515 ; n9515_not
g33038 not n6158 ; n6158_not
g33039 not n7283 ; n7283_not
g33040 not n9326 ; n9326_not
g33041 not n5168 ; n5168_not
g33042 not n7832 ; n7832_not
g33043 not n7535 ; n7535_not
g33044 not n7328 ; n7328_not
g33045 not n6383 ; n6383_not
g33046 not n7850 ; n7850_not
g33047 not n8642 ; n8642_not
g33048 not n7553 ; n7553_not
g33049 not n6365 ; n6365_not
g33050 not n7571 ; n7571_not
g33051 not n6347 ; n6347_not
g33052 not n6329 ; n6329_not
g33053 not n6194 ; n6194_not
g33054 not n6293 ; n6293_not
g33055 not n7607 ; n7607_not
g33056 not n7940 ; n7940_not
g33057 not n5861 ; n5861_not
g33058 not n9173 ; n9173_not
g33059 not n5834 ; n5834_not
g33060 not n8543 ; n8543_not
g33061 not n7913 ; n7913_not
g33062 not n7922 ; n7922_not
g33063 not n2864 ; n2864_not
g33064 not n9407 ; n9407_not
g33065 not n4871 ; n4871_not
g33066 not n8606 ; n8606_not
g33067 not n8273 ; n8273_not
g33068 not n6239 ; n6239_not
g33069 not n4961 ; n4961_not
g33070 not n6455 ; n6455_not
g33071 not n7823 ; n7823_not
g33072 not n6419 ; n6419_not
g33073 not n6851 ; n6851_not
g33074 not n9713 ; n9713_not
g33075 not n7337 ; n7337_not
g33076 not n9209 ; n9209_not
g33077 not n7085 ; n7085_not
g33078 not n9047 ; n9047_not
g33079 not n4646 ; n4646_not
g33080 not n5681 ; n5681_not
g33081 not n8804 ; n8804_not
g33082 not n7193 ; n7193_not
g33083 not n5366 ; n5366_not
g33084 not n4565 ; n4565_not
g33085 not n4664 ; n4664_not
g33086 not n4268 ; n4268_not
g33087 not n4484 ; n4484_not
g33088 not n5627 ; n5627_not
g33089 not n4592 ; n4592_not
g33090 not n8183 ; n8183_not
g33091 not n2918 ; n2918_not
g33092 not n8516 ; n8516_not
g33093 not n9425 ; n9425_not
g33094 not n7274 ; n7274_not
g33095 not n7049 ; n7049_not
g33096 not n5474 ; n5474_not
g33097 not n9830 ; n9830_not
g33098 not n9038 ; n9038_not
g33099 not n6941 ; n6941_not
g33100 not n9722 ; n9722_not
g33101 not n9731 ; n9731_not
g33102 not n7256 ; n7256_not
g33103 not n5393 ; n5393_not
g33104 not n5582 ; n5582_not
g33105 not n3818 ; n3818_not
g33106 not n7373 ; n7373_not
g33107 not n7076 ; n7076_not
g33108 not n8822 ; n8822_not
g33109 not n8237 ; n8237_not
g33110 not n9614 ; n9614_not
g33111 not n5357 ; n5357_not
g33112 not n7391 ; n7391_not
g33113 not n8552 ; n8552_not
g33114 not n3458 ; n3458_not
g33115 not n8219 ; n8219_not
g33116 not n5825 ; n5825_not
g33117 not n3629 ; n3629_not
g33118 not n5573 ; n5573_not
g33119 not n9650 ; n9650_not
g33120 not n5645 ; n5645_not
g33121 not n5456 ; n5456_not
g33122 not n4538 ; n4538_not
g33123 not n7257 ; n7257_not
g33124 not n5349 ; n5349_not
g33125 not n2388 ; n2388_not
g33126 not n1992 ; n1992_not
g33127 not n4935 ; n4935_not
g33128 not n2829 ; n2829_not
g33129 not n4485 ; n4485_not
g33130 not n4458 ; n4458_not
g33131 not n4467 ; n4467_not
g33132 not n8661 ; n8661_not
g33133 not n7572 ; n7572_not
g33134 not n7671 ; n7671_not
g33135 not n7707 ; n7707_not
g33136 not n6393 ; n6393_not
g33137 not n7608 ; n7608_not
g33138 not n7095 ; n7095_not
g33139 not n7644 ; n7644_not
g33140 not n6177 ; n6177_not
g33141 not n8418 ; n8418_not
g33142 not n7176 ; n7176_not
g33143 not n6168 ; n6168_not
g33144 not n6591 ; n6591_not
g33145 not n7725 ; n7725_not
g33146 not n7077 ; n7077_not
g33147 not n5646 ; n5646_not
g33148 not n8841 ; n8841_not
g33149 not n7239 ; n7239_not
g33150 not n7059 ; n7059_not
g33151 not n6492 ; n6492_not
g33152 not n4575 ; n4575_not
g33153 not n6807 ; n6807_not
g33154 not n4863 ; n4863_not
g33155 not n4179 ; n4179_not
g33156 not n4683 ; n4683_not
g33157 not n5907 ; n5907_not
g33158 not n7365 ; n7365_not
g33159 not n5925 ; n5925_not
g33160 not n8904 ; n8904_not
g33161 not n4917 ; n4917_not
g33162 not n5655 ; n5655_not
g33163 not n2838 ; n2838_not
g33164 not n4728 ; n4728_not
g33165 not n5835 ; n5835_not
g33166 not n5691 ; n5691_not
g33167 not n7428 ; n7428_not
g33168 not n6816 ; n6816_not
g33169 not n5853 ; n5853_not
g33170 not n7392 ; n7392_not
g33171 not n7446 ; n7446_not
g33172 not n8823 ; n8823_not
g33173 not n7464 ; n7464_not
g33174 not n4971 ; n4971_not
g33175 not n5952 ; n5952_not
g33176 not n6924 ; n6924_not
g33177 not n8544 ; n8544_not
g33178 not n4629 ; n4629_not
g33179 not n6942 ; n6942_not
g33180 not n2874 ; n2874_not
g33181 not n5844 ; n5844_not
g33182 not n6384 ; n6384_not
g33183 not n8940 ; n8940_not
g33184 not n5628 ; n5628_not
g33185 not n6348 ; n6348_not
g33186 not n7275 ; n7275_not
g33187 not n5943 ; n5943_not
g33188 not n6537 ; n6537_not
g33189 not n2928 ; n2928_not
g33190 not n4674 ; n4674_not
g33191 not n4656 ; n4656_not
g33192 not n4665 ; n4665_not
g33193 not n2892 ; n2892_not
g33194 not n7347 ; n7347_not
g33195 not n2856 ; n2856_not
g33196 not n8607 ; n8607_not
g33197 not n6906 ; n6906_not
g33198 not n8922 ; n8922_not
g33199 not n6267 ; n6267_not
g33200 not n6456 ; n6456_not
g33201 not n5394 ; n5394_not
g33202 not n5439 ; n5439_not
g33203 not n8238 ; n8238_not
g33204 not n9057 ; n9057_not
g33205 not n5457 ; n5457_not
g33206 not n8265 ; n8265_not
g33207 not n7491 ; n7491_not
g33208 not n7833 ; n7833_not
g33209 not n7815 ; n7815_not
g33210 not n5592 ; n5592_not
g33211 not n9714 ; n9714_not
g33212 not n8562 ; n8562_not
g33213 not n9543 ; n9543_not
g33214 not n8382 ; n8382_not
g33215 not n9435 ; n9435_not
g33216 not n9372 ; n9372_not
g33217 not n8463 ; n8463_not
g33218 not n9363 ; n9363_not
g33219 not n9345 ; n9345_not
g33220 not n8733 ; n8733_not
g33221 not n9039 ; n9039_not
g33222 not n9174 ; n9174_not
g33223 not n8526 ; n8526_not
g33224 not n8274 ; n8274_not
g33225 not n5574 ; n5574_not
g33226 not n9309 ; n9309_not
g33227 not n9453 ; n9453_not
g33228 not n8319 ; n8319_not
g33229 not n9660 ; n9660_not
g33230 not n9075 ; n9075_not
g33231 not n8337 ; n8337_not
g33232 not n8346 ; n8346_not
g33233 not n9624 ; n9624_not
g33234 not n9246 ; n9246_not
g33235 not n8364 ; n8364_not
g33236 not n9552 ; n9552_not
g33237 not n5547 ; n5547_not
g33238 not n7294 ; n7294_not
g33239 not n8194 ; n8194_not
g33240 not n4558 ; n4558_not
g33241 not n3964 ; n3964_not
g33242 not n5395 ; n5395_not
g33243 not n5629 ; n5629_not
g33244 not n9751 ; n9751_not
g33245 not n8158 ; n8158_not
g33246 not n4639 ; n4639_not
g33247 not n5377 ; n5377_not
g33248 not n5368 ; n5368_not
g33249 not n8266 ; n8266_not
g33250 not n7096 ; n7096_not
g33251 not n7735 ; n7735_not
g33252 not n8257 ; n8257_not
g33253 not n5449 ; n5449_not
g33254 not n7168 ; n7168_not
g33255 not n7186 ; n7186_not
g33256 not n8833 ; n8833_not
g33257 not n7870 ; n7870_not
g33258 not n4585 ; n4585_not
g33259 not n4927 ; n4927_not
g33260 not n7933 ; n7933_not
g33261 not n7915 ; n7915_not
g33262 not n7555 ; n7555_not
g33263 not n7708 ; n7708_not
g33264 not n7861 ; n7861_not
g33265 not n7852 ; n7852_not
g33266 not n8086 ; n8086_not
g33267 not n4684 ; n4684_not
g33268 not n8068 ; n8068_not
g33269 not n8617 ; n8617_not
g33270 not n7960 ; n7960_not
g33271 not n4477 ; n4477_not
g33272 not n4846 ; n4846_not
g33273 not n4918 ; n4918_not
g33274 not n5593 ; n5593_not
g33275 not n7780 ; n7780_not
g33276 not n9382 ; n9382_not
g33277 not n6439 ; n6439_not
g33278 not n6475 ; n6475_not
g33279 not n2848 ; n2848_not
g33280 not n2884 ; n2884_not
g33281 not n5557 ; n5557_not
g33282 not n6538 ; n6538_not
g33283 not n5962 ; n5962_not
g33284 not n5944 ; n5944_not
g33285 not n9463 ; n9463_not
g33286 not n5908 ; n5908_not
g33287 not n9481 ; n9481_not
g33288 not n9490 ; n9490_not
g33289 not n8707 ; n8707_not
g33290 not n9526 ; n9526_not
g33291 not n2866 ; n2866_not
g33292 not n9148 ; n9148_not
g33293 not n9193 ; n9193_not
g33294 not n8491 ; n8491_not
g33295 not n9238 ; n9238_not
g33296 not n9094 ; n9094_not
g33297 not n8806 ; n8806_not
g33298 not n6349 ; n6349_not
g33299 not n8680 ; n8680_not
g33300 not n6358 ; n6358_not
g33301 not n9337 ; n9337_not
g33302 not n8473 ; n8473_not
g33303 not n6385 ; n6385_not
g33304 not n7753 ; n7753_not
g33305 not n8581 ; n8581_not
g33306 not n6925 ; n6925_not
g33307 not n9706 ; n9706_not
g33308 not n9715 ; n9715_not
g33309 not n5485 ; n5485_not
g33310 not n9625 ; n9625_not
g33311 not n9544 ; n9544_not
g33312 not n4189 ; n4189_not
g33313 not n8635 ; n8635_not
g33314 not n5647 ; n5647_not
g33315 not n9832 ; n9832_not
g33316 not n9850 ; n9850_not
g33317 not n8284 ; n8284_not
g33318 not n5539 ; n5539_not
g33319 not n5467 ; n5467_not
g33320 not n5836 ; n5836_not
g33321 not n6691 ; n6691_not
g33322 not n8365 ; n8365_not
g33323 not n9562 ; n9562_not
g33324 not n9580 ; n9580_not
g33325 not n5719 ; n5719_not
g33326 not n9607 ; n9607_not
g33327 not n8347 ; n8347_not
g33328 not n8725 ; n8725_not
g33329 not n6808 ; n6808_not
g33330 not n8545 ; n8545_not
g33331 not n3883 ; n3883_not
g33332 not n8437 ; n8437_not
g33333 not n6970 ; n6970_not
g33334 not n6907 ; n6907_not
g33335 not n4954 ; n4954_not
g33336 not n7582 ; n7582_not
g33337 not n7690 ; n7690_not
g33338 not n4981 ; n4981_not
g33339 not n7537 ; n7537_not
g33340 not n7591 ; n7591_not
g33341 not n7816 ; n7816_not
g33342 not n7663 ; n7663_not
g33343 not n5584 ; n5584_not
g33344 not n7807 ; n7807_not
g33345 not n7492 ; n7492_not
g33346 not n7618 ; n7618_not
g33347 not n1877 ; n1877_not
g33348 not n7646 ; n7646_not
g33349 not n8834 ; n8834_not
g33350 not n7826 ; n7826_not
g33351 not n5675 ; n5675_not
g33352 not n4685 ; n4685_not
g33353 not n7439 ; n7439_not
g33354 not n8672 ; n8672_not
g33355 not n5666 ; n5666_not
g33356 not n8339 ; n8339_not
g33357 not n6449 ; n6449_not
g33358 not n8582 ; n8582_not
g33359 not n4748 ; n4748_not
g33360 not n8456 ; n8456_not
g33361 not n7484 ; n7484_not
g33362 not n9635 ; n9635_not
g33363 not n7169 ; n7169_not
g33364 not n2894 ; n2894_not
g33365 not n8555 ; n8555_not
g33366 not n6368 ; n6368_not
g33367 not n9338 ; n9338_not
g33368 not n5873 ; n5873_not
g33369 not n8348 ; n8348_not
g33370 not n9842 ; n9842_not
g33371 not n8159 ; n8159_not
g33372 not n7457 ; n7457_not
g33373 not n8069 ; n8069_not
g33374 not n7268 ; n7268_not
g33375 not n9095 ; n9095_not
g33376 not n7385 ; n7385_not
g33377 not n2876 ; n2876_not
g33378 not n5558 ; n5558_not
g33379 not n7664 ; n7664_not
g33380 not n9428 ; n9428_not
g33381 not n5972 ; n5972_not
g33382 not n8474 ; n8474_not
g33383 not n9383 ; n9383_not
g33384 not n4577 ; n4577_not
g33385 not n8690 ; n8690_not
g33386 not n5765 ; n5765_not
g33387 not n8366 ; n8366_not
g33388 not n7637 ; n7637_not
g33389 not n6476 ; n6476_not
g33390 not n6692 ; n6692_not
g33391 not n5567 ; n5567_not
g33392 not n3839 ; n3839_not
g33393 not n9545 ; n9545_not
g33394 not n7286 ; n7286_not
g33395 not n2858 ; n2858_not
g33396 not n9365 ; n9365_not
g33397 not n7583 ; n7583_not
g33398 not n5486 ; n5486_not
g33399 not n6188 ; n6188_not
g33400 not n9914 ; n9914_not
g33401 not n7925 ; n7925_not
g33402 not n4658 ; n4658_not
g33403 not n7763 ; n7763_not
g33404 not n6908 ; n6908_not
g33405 not n9932 ; n9932_not
g33406 not n7943 ; n7943_not
g33407 not n5909 ; n5909_not
g33408 not n8627 ; n8627_not
g33409 not n9950 ; n9950_not
g33410 not n4919 ; n4919_not
g33411 not n5918 ; n5918_not
g33412 not n7718 ; n7718_not
g33413 not n9743 ; n9743_not
g33414 not n8519 ; n8519_not
g33415 not n9860 ; n9860_not
g33416 not n8249 ; n8249_not
g33417 not n8654 ; n8654_not
g33418 not n7862 ; n7862_not
g33419 not n9725 ; n9725_not
g33420 not n5378 ; n5378_not
g33421 not n6935 ; n6935_not
g33422 not n9491 ; n9491_not
g33423 not n9707 ; n9707_not
g33424 not n7736 ; n7736_not
g33425 not n6179 ; n6179_not
g33426 not n6926 ; n6926_not
g33427 not n9167 ; n9167_not
g33428 not n8375 ; n8375_not
g33429 not n9185 ; n9185_not
g33430 not n9473 ; n9473_not
g33431 not n6872 ; n6872_not
g33432 not n4892 ; n4892_not
g33433 not n8087 ; n8087_not
g33434 not n4883 ; n4883_not
g33435 not n7079 ; n7079_not
g33436 not n9275 ; n9275_not
g33437 not n9293 ; n9293_not
g33438 not n7619 ; n7619_not
g33439 not n9653 ; n9653_not
g33440 not n7790 ; n7790_not
g33441 not n7358 ; n7358_not
g33442 not n5882 ; n5882_not
g33443 not n3965 ; n3965_not
g33444 not n6890 ; n6890_not
g33445 not n8267 ; n8267_not
g33446 not n4478 ; n4478_not
g33447 not n7493 ; n7493_not
g33448 not n6881 ; n6881_not
g33449 not n1779 ; n1779_not
g33450 not n9870 ; n9870_not
g33451 not n8709 ; n8709_not
g33452 not n4938 ; n4938_not
g33453 not n7278 ; n7278_not
g33454 not n9519 ; n9519_not
g33455 not n7296 ; n7296_not
g33456 not n9492 ; n9492_not
g33457 not n5388 ; n5388_not
g33458 not n9645 ; n9645_not
g33459 not n9672 ; n9672_not
g33460 not n6873 ; n6873_not
g33461 not n4479 ; n4479_not
g33462 not n8817 ; n8817_not
g33463 not n7836 ; n7836_not
g33464 not n6891 ; n6891_not
g33465 not n9951 ; n9951_not
g33466 not n3885 ; n3885_not
g33467 not n9933 ; n9933_not
g33468 not n5487 ; n5487_not
g33469 not n9915 ; n9915_not
g33470 not n8286 ; n8286_not
g33471 not n9708 ; n9708_not
g33472 not n8628 ; n8628_not
g33473 not n9357 ; n9357_not
g33474 not n6945 ; n6945_not
g33475 not n9690 ; n9690_not
g33476 not n8187 ; n8187_not
g33477 not n9555 ; n9555_not
g33478 not n8718 ; n8718_not
g33479 not n8295 ; n8295_not
g33480 not n4578 ; n4578_not
g33481 not n8835 ; n8835_not
g33482 not n6963 ; n6963_not
g33483 not n8790 ; n8790_not
g33484 not n6792 ; n6792_not
g33485 not n7485 ; n7485_not
g33486 not n8484 ; n8484_not
g33487 not n8673 ; n8673_not
g33488 not n6369 ; n6369_not
g33489 not n6396 ; n6396_not
g33490 not n9339 ; n9339_not
g33491 not n5586 ; n5586_not
g33492 not n6378 ; n6378_not
g33493 not n7683 ; n7683_not
g33494 not n4974 ; n4974_not
g33495 not n8727 ; n8727_not
g33496 not n7863 ; n7863_not
g33497 not n7539 ; n7539_not
g33498 not n7566 ; n7566_not
g33499 not n8529 ; n8529_not
g33500 not n7548 ; n7548_not
g33501 not n8664 ; n8664_not
g33502 not n5658 ; n5658_not
g33503 not n9186 ; n9186_not
g33504 not n9177 ; n9177_not
g33505 not n4947 ; n4947_not
g33506 not n6189 ; n6189_not
g33507 not n7584 ; n7584_not
g33508 not n5865 ; n5865_not
g33509 not n7764 ; n7764_not
g33510 not n7665 ; n7665_not
g33511 not n4668 ; n4668_not
g33512 not n8088 ; n8088_not
g33513 not n2868 ; n2868_not
g33514 not n9861 ; n9861_not
g33515 not n5982 ; n5982_not
g33516 not n9474 ; n9474_not
g33517 not n4848 ; n4848_not
g33518 not n5928 ; n5928_not
g33519 not n9438 ; n9438_not
g33520 not n2886 ; n2886_not
g33521 not n8592 ; n8592_not
g33522 not n4695 ; n4695_not
g33523 not n9456 ; n9456_not
g33524 not n5379 ; n5379_not
g33525 not n7746 ; n7746_not
g33526 not n5892 ; n5892_not
g33527 not n7944 ; n7944_not
g33528 not n6459 ; n6459_not
g33529 not n9393 ; n9393_not
g33530 not n8385 ; n8385_not
g33531 not n4875 ; n4875_not
g33532 not n9466 ; n9466_not
g33533 not n3877 ; n3877_not
g33534 not n6397 ; n6397_not
g33535 not n5596 ; n5596_not
g33536 not n5947 ; n5947_not
g33537 not n5929 ; n5929_not
g33538 not n6919 ; n6919_not
g33539 not n6199 ; n6199_not
g33540 not n8296 ; n8296_not
g33541 not n9439 ; n9439_not
g33542 not n6946 ; n6946_not
g33543 not n9277 ; n9277_not
g33544 not n9475 ; n9475_not
g33545 not n9736 ; n9736_not
g33546 not n9727 ; n9727_not
g33547 not n7927 ; n7927_not
g33548 not n8386 ; n8386_not
g33549 not n9646 ; n9646_not
g33550 not n9295 ; n9295_not
g33551 not n9628 ; n9628_not
g33552 not n6748 ; n6748_not
g33553 not n8449 ; n8449_not
g33554 not n6793 ; n6793_not
g33555 not n8683 ; n8683_not
g33556 not n5668 ; n5668_not
g33557 not n8359 ; n8359_not
g33558 not n6388 ; n6388_not
g33559 not n8719 ; n8719_not
g33560 not n8395 ; n8395_not
g33561 not n5497 ; n5497_not
g33562 not n5893 ; n5893_not
g33563 not n9691 ; n9691_not
g33564 not n9682 ; n9682_not
g33565 not n6892 ; n6892_not
g33566 not n7279 ; n7279_not
g33567 not n9196 ; n9196_not
g33568 not n9529 ; n9529_not
g33569 not n5866 ; n5866_not
g33570 not n6874 ; n6874_not
g33571 not n5767 ; n5767_not
g33572 not n2896 ; n2896_not
g33573 not n2878 ; n2878_not
g33574 not n7693 ; n7693_not
g33575 not n4678 ; n4678_not
g33576 not n9745 ; n9745_not
g33577 not n5398 ; n5398_not
g33578 not n4588 ; n4588_not
g33579 not n8197 ; n8197_not
g33580 not n8818 ; n8818_not
g33581 not n9970 ; n9970_not
g33582 not n9952 ; n9952_not
g33583 not n7549 ; n7549_not
g33584 not n7567 ; n7567_not
g33585 not n4966 ; n4966_not
g33586 not n7954 ; n7954_not
g33587 not n7972 ; n7972_not
g33588 not n8872 ; n8872_not
g33589 not n3967 ; n3967_not
g33590 not n9844 ; n9844_not
g33591 not n4849 ; n4849_not
g33592 not n7486 ; n7486_not
g33593 not n4876 ; n4876_not
g33594 not n7990 ; n7990_not
g33595 not n7837 ; n7837_not
g33596 not n9916 ; n9916_not
g33597 not n8629 ; n8629_not
g33598 not n9934 ; n9934_not
g33599 not n6587 ; n6587_not
g33600 not n6479 ; n6479_not
g33601 not n8387 ; n8387_not
g33602 not n5948 ; n5948_not
g33603 not n6695 ; n6695_not
g33604 not n7658 ; n7658_not
g33605 not n4688 ; n4688_not
g33606 not n9449 ; n9449_not
g33607 not n5975 ; n5975_not
g33608 not n2888 ; n2888_not
g33609 not n9872 ; n9872_not
g33610 not n8693 ; n8693_not
g33611 not n9737 ; n9737_not
g33612 not n8567 ; n8567_not
g33613 not n6929 ; n6929_not
g33614 not n8369 ; n8369_not
g33615 not n7739 ; n7739_not
g33616 not n7793 ; n7793_not
g33617 not n4598 ; n4598_not
g33618 not n5858 ; n5858_not
g33619 not n8792 ; n8792_not
g33620 not n8945 ; n8945_not
g33621 not n5876 ; n5876_not
g33622 not n5894 ; n5894_not
g33623 not n9485 ; n9485_not
g33624 not n8099 ; n8099_not
g33625 not n7847 ; n7847_not
g33626 not n7469 ; n7469_not
g33627 not n7991 ; n7991_not
g33628 not n4886 ; n4886_not
g33629 not n7289 ; n7289_not
g33630 not n7973 ; n7973_not
g33631 not n8909 ; n8909_not
g33632 not n8297 ; n8297_not
g33633 not n8927 ; n8927_not
g33634 not n7955 ; n7955_not
g33635 not n7775 ; n7775_not
g33636 not n7694 ; n7694_not
g33637 not n9467 ; n9467_not
g33638 not n4967 ; n4967_not
g33639 not n6488 ; n6488_not
g33640 not n7856 ; n7856_not
g33641 not n9386 ; n9386_not
g33642 not n8891 ; n8891_not
g33643 not n8459 ; n8459_not
g33644 not n7568 ; n7568_not
g33645 not n9359 ; n9359_not
g33646 not n8963 ; n8963_not
g33647 not n6956 ; n6956_not
g33648 not n7577 ; n7577_not
g33649 not n8477 ; n8477_not
g33650 not n6389 ; n6389_not
g33651 not n4868 ; n4868_not
g33652 not n6848 ; n6848_not
g33653 not n8819 ; n8819_not
g33654 not n8981 ; n8981_not
g33655 not n9638 ; n9638_not
g33656 not n7838 ; n7838_not
g33657 not n8747 ; n8747_not
g33658 not n8828 ; n8828_not
g33659 not n5399 ; n5399_not
g33660 not n9647 ; n9647_not
g33661 not n6965 ; n6965_not
g33662 not n5678 ; n5678_not
g33663 not n8558 ; n8558_not
g33664 not n8198 ; n8198_not
g33665 not n7668 ; n7668_not
g33666 not n7749 ; n7749_not
g33667 not n8694 ; n8694_not
g33668 not n9396 ; n9396_not
g33669 not n7785 ; n7785_not
g33670 not n4689 ; n4689_not
g33671 not n8568 ; n8568_not
g33672 not n9738 ; n9738_not
g33673 not n6489 ; n6489_not
g33674 not n7839 ; n7839_not
g33675 not n9927 ; n9927_not
g33676 not n6795 ; n6795_not
g33677 not n5967 ; n5967_not
g33678 not n5679 ; n5679_not
g33679 not n6588 ; n6588_not
g33680 not n9468 ; n9468_not
g33681 not n8838 ; n8838_not
g33682 not n8649 ; n8649_not
g33683 not n9963 ; n9963_not
g33684 not n8928 ; n8928_not
g33685 not n9828 ; n9828_not
g33686 not n4968 ; n4968_not
g33687 not n8964 ; n8964_not
g33688 not n6885 ; n6885_not
g33689 not n9981 ; n9981_not
g33690 not n7938 ; n7938_not
g33691 not n9765 ; n9765_not
g33692 not n7956 ; n7956_not
g33693 not n9945 ; n9945_not
g33694 not n8667 ; n8667_not
g33695 not n6867 ; n6867_not
g33696 not n9837 ; n9837_not
g33697 not n7974 ; n7974_not
g33698 not n8487 ; n8487_not
g33699 not n9297 ; n9297_not
g33700 not n7587 ; n7587_not
g33701 not n9639 ; n9639_not
g33702 not a[0] ; a[0]_not
g33703 not n2898 ; n2898_not
g33704 not n9855 ; n9855_not
g33705 not n8874 ; n8874_not
g33706 not n8892 ; n8892_not
g33707 not n9585 ; n9585_not
g33708 not n9891 ; n9891_not
g33709 not n8982 ; n8982_not
g33710 not n9909 ; n9909_not
g33711 not n9567 ; n9567_not
g33712 not n4986 ; n4986_not
g33713 not n8865 ; n8865_not
g33714 not n8946 ; n8946_not
g33715 not n9882 ; n9882_not
g33716 not n9558 ; n9558_not
g33717 not n8199 ; n8199_not
g33718 not n7597 ; n7597_not
g33719 not n8839 ; n8839_not
g33720 not n9883 ; n9883_not
g33721 not n8848 ; n8848_not
g33722 not n9667 ; n9667_not
g33723 not n7489 ; n7489_not
g33724 not n9838 ; n9838_not
g33725 not n4897 ; n4897_not
g33726 not n7984 ; n7984_not
g33727 not n5896 ; n5896_not
g33728 not n8596 ; n8596_not
g33729 not n9586 ; n9586_not
g33730 not n8929 ; n8929_not
g33731 not n9865 ; n9865_not
g33732 not n8569 ; n8569_not
g33733 not n8983 ; n8983_not
g33734 not n8659 ; n8659_not
g33735 not n7786 ; n7786_not
g33736 not n9685 ; n9685_not
g33737 not n7768 ; n7768_not
g33738 not n5698 ; n5698_not
g33739 not n8893 ; n8893_not
g33740 not n8389 ; n8389_not
g33741 not n7588 ; n7588_not
g33742 not n9379 ; n9379_not
g33743 not n9856 ; n9856_not
g33744 not n8488 ; n8488_not
g33745 not n4987 ; n4987_not
g33746 not n9478 ; n9478_not
g33747 not n9568 ; n9568_not
g33748 not n6895 ; n6895_not
g33749 not n8965 ; n8965_not
g33750 not n7939 ; n7939_not
g33751 not n8794 ; n8794_not
g33752 not n8695 ; n8695_not
g33753 not n8947 ; n8947_not
g33754 not n6877 ; n6877_not
g33755 not n9397 ; n9397_not
g33756 not n5887 ; n5887_not
g33757 not n5968 ; n5968_not
g33758 not a[1] ; a[1]_not
g33759 not n5599 ; n5599_not
g33760 not n8749 ; n8749_not
g33761 not a[2] ; a[2]_not
g33762 not n8696 ; n8696_not
g33763 not n8498 ; n8498_not
g33764 not n9587 ; n9587_not
g33765 not n6986 ; n6986_not
g33766 not n9785 ; n9785_not
g33767 not n9569 ; n9569_not
g33768 not n9767 ; n9767_not
g33769 not n9839 ; n9839_not
g33770 not n7994 ; n7994_not
g33771 not n7967 ; n7967_not
g33772 not n9677 ; n9677_not
g33773 not n7949 ; n7949_not
g33774 not n4898 ; n4898_not
g33775 not n7868 ; n7868_not
g33776 not n9749 ; n9749_not
g33777 not n7697 ; n7697_not
g33778 not n7787 ; n7787_not
g33779 not n4988 ; n4988_not
g33780 not n5987 ; n5987_not
g33781 not n5888 ; n5888_not
g33782 not n5969 ; n5969_not
g33783 not n6896 ; n6896_not
g33784 not n6878 ; n6878_not
g33785 not n9857 ; n9857_not
g33786 not n7589 ; n7589_not
g33787 not n6798 ; n6798_not
g33788 not n9867 ; n9867_not
g33789 not n7797 ; n7797_not
g33790 not n7959 ; n7959_not
g33791 not n6879 ; n6879_not
g33792 not n9678 ; n9678_not
g33793 not n5889 ; n5889_not
g33794 not n8697 ; n8697_not
g33795 not n8994 ; n8994_not
g33796 not n8688 ; n8688_not
g33797 not n8958 ; n8958_not
g33798 not n8886 ; n8886_not
g33799 not n8976 ; n8976_not
g33800 not n7995 ; n7995_not
g33801 not a[3] ; a[3]_not
g33802 not n5988 ; n5988_not
g33803 not n4899 ; n4899_not
g33804 not n6978 ; n6978_not
g33805 not n7977 ; n7977_not
g33806 not n8589 ; n8589_not
g33807 not n9886 ; n9886_not
g33808 not n8689 ; n8689_not
g33809 not n7978 ; n7978_not
g33810 not n9679 ; n9679_not
g33811 not n6979 ; n6979_not
g33812 not n9787 ; n9787_not
g33813 not a[4] ; a[4]_not
g33814 not n5989 ; n5989_not
g33815 not a[5] ; a[5]_not
g33816 not n8879 ; n8879_not
g33817 not n9698 ; n9698_not
g33818 not n9599 ; n9599_not
g33819 not n9896 ; n9896_not
g33820 not n9968 ; n9968_not
g33821 not n9986 ; n9986_not
g33822 not n6989 ; n6989_not
g33823 not n7997 ; n7997_not
g33824 not n9969 ; n9969_not
g33825 not n7989 ; n7989_not
g33826 not a[6] ; a[6]_not
g33827 not n9987 ; n9987_not
g33828 not n9897 ; n9897_not
g33829 not n9879 ; n9879_not
g33830 not n8799 ; n8799_not
g33831 not a[7] ; a[7]_not
g33832 not n9988 ; n9988_not
g33833 not n9898 ; n9898_not
g33834 not a[8] ; a[8]_not
g33835 not n8999 ; n8999_not
g33836 not a[9] ; a[9]_not
g33837 not n9999 ; n9999_not
g33838 not n20000 ; n20000_not
g33839 not n10100 ; n10100_not
g33840 not n30000 ; n30000_not
g33841 not n10110 ; n10110_not
g33842 not n20001 ; n20001_not
g33843 not n11200 ; n11200_not
g33844 not n21010 ; n21010_not
g33845 not n20011 ; n20011_not
g33846 not n12100 ; n12100_not
g33847 not n12001 ; n12001_not
g33848 not n30001 ; n30001_not
g33849 not n13000 ; n13000_not
g33850 not n30020 ; n30020_not
g33851 not n23000 ; n23000_not
g33852 not n20120 ; n20120_not
g33853 not n20210 ; n20210_not
g33854 not n11201 ; n11201_not
g33855 not n10004 ; n10004_not
g33856 not n10040 ; n10040_not
g33857 not n31100 ; n31100_not
g33858 not n10121 ; n10121_not
g33859 not n10202 ; n10202_not
g33860 not n10301 ; n10301_not
g33861 not n22010 ; n22010_not
g33862 not n14000 ; n14000_not
g33863 not n10310 ; n10310_not
g33864 not n21002 ; n21002_not
g33865 not n10220 ; n10220_not
g33866 not n13001 ; n13001_not
g33867 not n21200 ; n21200_not
g33868 not n10140 ; n10140_not
g33869 not n10230 ; n10230_not
g33870 not n10050 ; n10050_not
g33871 not n14010 ; n14010_not
g33872 not n10005 ; n10005_not
g33873 not n10302 ; n10302_not
g33874 not n10320 ; n10320_not
g33875 not n32100 ; n32100_not
g33876 not n11310 ; n11310_not
g33877 not n20013 ; n20013_not
g33878 not n20022 ; n20022_not
g33879 not n20121 ; n20121_not
g33880 not n20130 ; n20130_not
g33881 not n11211 ; n11211_not
g33882 not n20220 ; n20220_not
g33883 not n20031 ; n20031_not
g33884 not n21003 ; n21003_not
g33885 not n11031 ; n11031_not
g33886 not n22002 ; n22002_not
g33887 not n22101 ; n22101_not
g33888 not n22200 ; n22200_not
g33889 not n31011 ; n31011_not
g33890 not n30211 ; n30211_not
g33891 not n20140 ; n20140_not
g33892 not n15010 ; n15010_not
g33893 not n21130 ; n21130_not
g33894 not n20203 ; n20203_not
g33895 not n30202 ; n30202_not
g33896 not n12040 ; n12040_not
g33897 not n11032 ; n11032_not
g33898 not n20302 ; n20302_not
g33899 not n10006 ; n10006_not
g33900 not n10033 ; n10033_not
g33901 not n11401 ; n11401_not
g33902 not n20410 ; n20410_not
g33903 not n10240 ; n10240_not
g33904 not n12031 ; n12031_not
g33905 not n10051 ; n10051_not
g33906 not n20221 ; n20221_not
g33907 not n14101 ; n14101_not
g33908 not n10114 ; n10114_not
g33909 not n30400 ; n30400_not
g33910 not n10150 ; n10150_not
g33911 not n30004 ; n30004_not
g33912 not n24010 ; n24010_not
g33913 not n11320 ; n11320_not
g33914 not n12130 ; n12130_not
g33915 not n22300 ; n22300_not
g33916 not n30013 ; n30013_not
g33917 not n21112 ; n21112_not
g33918 not n10303 ; n10303_not
g33919 not n12301 ; n12301_not
g33920 not n23101 ; n23101_not
g33921 not n15100 ; n15100_not
g33922 not n30310 ; n30310_not
g33923 not n20023 ; n20023_not
g33924 not n31012 ; n31012_not
g33925 not n11500 ; n11500_not
g33926 not n14011 ; n14011_not
g33927 not n21013 ; n21013_not
g33928 not n30203 ; n30203_not
g33929 not n30221 ; n30221_not
g33930 not n30230 ; n30230_not
g33931 not n10340 ; n10340_not
g33932 not n10322 ; n10322_not
g33933 not n10223 ; n10223_not
g33934 not n10241 ; n10241_not
g33935 not n10205 ; n10205_not
g33936 not n11114 ; n11114_not
g33937 not n11132 ; n11132_not
g33938 not n14030 ; n14030_not
g33939 not n30005 ; n30005_not
g33940 not n32102 ; n32102_not
g33941 not n23012 ; n23012_not
g33942 not n11303 ; n11303_not
g33943 not n12311 ; n12311_not
g33944 not n32003 ; n32003_not
g33945 not n11240 ; n11240_not
g33946 not n30023 ; n30023_not
g33947 not n30032 ; n30032_not
g33948 not n23120 ; n23120_not
g33949 not n20024 ; n20024_not
g33950 not n20051 ; n20051_not
g33951 not n20114 ; n20114_not
g33952 not n20141 ; n20141_not
g33953 not n11222 ; n11222_not
g33954 not n31013 ; n31013_not
g33955 not n13031 ; n13031_not
g33956 not n32021 ; n32021_not
g33957 not n20231 ; n20231_not
g33958 not n32012 ; n32012_not
g33959 not n10043 ; n10043_not
g33960 not n20411 ; n20411_not
g33961 not n10052 ; n10052_not
g33962 not n14111 ; n14111_not
g33963 not n12212 ; n12212_not
g33964 not n11150 ; n11150_not
g33965 not n10124 ; n10124_not
g33966 not n22220 ; n22220_not
g33967 not n21131 ; n21131_not
g33968 not n12014 ; n12014_not
g33969 not n22022 ; n22022_not
g33970 not n21203 ; n21203_not
g33971 not n10610 ; n10610_not
g33972 not n11321 ; n11321_not
g33973 not n11402 ; n11402_not
g33974 not n30401 ; n30401_not
g33975 not n21410 ; n21410_not
g33976 not n11060 ; n11060_not
g33977 not n21302 ; n21302_not
g33978 not n21401 ; n21401_not
g33979 not n21122 ; n21122_not
g33980 not n22310 ; n22310_not
g33981 not n16010 ; n16010_not
g33982 not n30500 ; n30500_not
g33983 not n24011 ; n24011_not
g33984 not n11510 ; n11510_not
g33985 not n12113 ; n12113_not
g33986 not n25010 ; n25010_not
g33987 not n10331 ; n10331_not
g33988 not n21320 ; n21320_not
g33989 not n20124 ; n20124_not
g33990 not n23040 ; n23040_not
g33991 not n23220 ; n23220_not
g33992 not n11430 ; n11430_not
g33993 not n21123 ; n21123_not
g33994 not n21204 ; n21204_not
g33995 not n16200 ; n16200_not
g33996 not n21411 ; n21411_not
g33997 not n21321 ; n21321_not
g33998 not n18000 ; n18000_not
g33999 not n22140 ; n22140_not
g34000 not n15003 ; n15003_not
g34001 not n17001 ; n17001_not
g34002 not n11322 ; n11322_not
g34003 not n24021 ; n24021_not
g34004 not n11250 ; n11250_not
g34005 not n22230 ; n22230_not
g34006 not n11610 ; n11610_not
g34007 not n11511 ; n11511_not
g34008 not n12321 ; n12321_not
g34009 not n14310 ; n14310_not
g34010 not n11232 ; n11232_not
g34011 not n22212 ; n22212_not
g34012 not n22104 ; n22104_not
g34013 not n22041 ; n22041_not
g34014 not n22005 ; n22005_not
g34015 not n16101 ; n16101_not
g34016 not n10044 ; n10044_not
g34017 not n10125 ; n10125_not
g34018 not n10233 ; n10233_not
g34019 not n12024 ; n12024_not
g34020 not n26001 ; n26001_not
g34021 not n12051 ; n12051_not
g34022 not n12060 ; n12060_not
g34023 not n15030 ; n15030_not
g34024 not n10242 ; n10242_not
g34025 not n15111 ; n15111_not
g34026 not n10332 ; n10332_not
g34027 not n11115 ; n11115_not
g34028 not n26100 ; n26100_not
g34029 not n21024 ; n21024_not
g34030 not n21042 ; n21042_not
g34031 not n11043 ; n11043_not
g34032 not n21051 ; n21051_not
g34033 not n21105 ; n21105_not
g34034 not n12123 ; n12123_not
g34035 not n12150 ; n12150_not
g34036 not n10026 ; n10026_not
g34037 not n25101 ; n25101_not
g34038 not n12303 ; n12303_not
g34039 not n21312 ; n21312_not
g34040 not n10512 ; n10512_not
g34041 not n12222 ; n12222_not
g34042 not n10062 ; n10062_not
g34043 not n11070 ; n11070_not
g34044 not n11412 ; n11412_not
g34045 not n10080 ; n10080_not
g34046 not n11151 ; n11151_not
g34047 not n10107 ; n10107_not
g34048 not n10800 ; n10800_not
g34049 not n21141 ; n21141_not
g34050 not n11133 ; n11133_not
g34051 not n10422 ; n10422_not
g34052 not n10413 ; n10413_not
g34053 not n20601 ; n20601_not
g34054 not n20610 ; n20610_not
g34055 not n30420 ; n30420_not
g34056 not n30150 ; n30150_not
g34057 not n30222 ; n30222_not
g34058 not n32022 ; n32022_not
g34059 not n32004 ; n32004_not
g34060 not n14004 ; n14004_not
g34061 not n32040 ; n32040_not
g34062 not n31221 ; n31221_not
g34063 not n30024 ; n30024_not
g34064 not n14031 ; n14031_not
g34065 not n31500 ; n31500_not
g34066 not n30240 ; n30240_not
g34067 not n14130 ; n14130_not
g34068 not n32013 ; n32013_not
g34069 not n14022 ; n14022_not
g34070 not n32112 ; n32112_not
g34071 not n13311 ; n13311_not
g34072 not n30042 ; n30042_not
g34073 not n31113 ; n31113_not
g34074 not n14112 ; n14112_not
g34075 not n12313 ; n12313_not
g34076 not n15400 ; n15400_not
g34077 not n20017 ; n20017_not
g34078 not n31132 ; n31132_not
g34079 not n23131 ; n23131_not
g34080 not n31330 ; n31330_not
g34081 not n22204 ; n22204_not
g34082 not n11152 ; n11152_not
g34083 not n25120 ; n25120_not
g34084 not n12007 ; n12007_not
g34085 not n21430 ; n21430_not
g34086 not n30421 ; n30421_not
g34087 not n11170 ; n11170_not
g34088 not n20350 ; n20350_not
g34089 not n12331 ; n12331_not
g34090 not n20008 ; n20008_not
g34091 not n25102 ; n25102_not
g34092 not n15004 ; n15004_not
g34093 not n11215 ; n11215_not
g34094 not n22330 ; n22330_not
g34095 not n21232 ; n21232_not
g34096 not n22150 ; n22150_not
g34097 not n31033 ; n31033_not
g34098 not n21070 ; n21070_not
g34099 not n20053 ; n20053_not
g34100 not n10153 ; n10153_not
g34101 not n20314 ; n20314_not
g34102 not n20404 ; n20404_not
g34103 not n13240 ; n13240_not
g34104 not n31240 ; n31240_not
g34105 not n21124 ; n21124_not
g34106 not n12205 ; n12205_not
g34107 not n10540 ; n10540_not
g34108 not n26011 ; n26011_not
g34109 not n16210 ; n16210_not
g34110 not n30412 ; n30412_not
g34111 not n31303 ; n31303_not
g34112 not n20800 ; n20800_not
g34113 not n11053 ; n11053_not
g34114 not n13501 ; n13501_not
g34115 not n30160 ; n30160_not
g34116 not n20125 ; n20125_not
g34117 not n10522 ; n10522_not
g34118 not n14122 ; n14122_not
g34119 not n20035 ; n20035_not
g34120 not n20431 ; n20431_not
g34121 not n10306 ; n10306_not
g34122 not n23320 ; n23320_not
g34123 not n20071 ; n20071_not
g34124 not n10045 ; n10045_not
g34125 not n24211 ; n24211_not
g34126 not n10135 ; n10135_not
g34127 not n21241 ; n21241_not
g34128 not n31114 ; n31114_not
g34129 not n32050 ; n32050_not
g34130 not n22222 ; n22222_not
g34131 not n12241 ; n12241_not
g34132 not n13321 ; n13321_not
g34133 not n32041 ; n32041_not
g34134 not n20161 ; n20161_not
g34135 not n14320 ; n14320_not
g34136 not n15130 ; n15130_not
g34137 not n20224 ; n20224_not
g34138 not n22240 ; n22240_not
g34139 not n31141 ; n31141_not
g34140 not n13510 ; n13510_not
g34141 not n11116 ; n11116_not
g34142 not n31006 ; n31006_not
g34143 not n22231 ; n22231_not
g34144 not n15112 ; n15112_not
g34145 not n18010 ; n18010_not
g34146 not n20620 ; n20620_not
g34147 not n30322 ; n30322_not
g34148 not n14230 ; n14230_not
g34149 not n12520 ; n12520_not
g34150 not n23041 ; n23041_not
g34151 not n11512 ; n11512_not
g34152 not n24310 ; n24310_not
g34153 not n17200 ; n17200_not
g34154 not n26200 ; n26200_not
g34155 not n22501 ; n22501_not
g34156 not n10234 ; n10234_not
g34157 not n24004 ; n24004_not
g34158 not n11332 ; n11332_not
g34159 not n10216 ; n10216_not
g34160 not n17020 ; n17020_not
g34161 not n11071 ; n11071_not
g34162 not n11422 ; n11422_not
g34163 not n14302 ; n14302_not
g34164 not n31411 ; n31411_not
g34165 not n21214 ; n21214_not
g34166 not n11440 ; n11440_not
g34167 not n15220 ; n15220_not
g34168 not n11044 ; n11044_not
g34169 not n12106 ; n12106_not
g34170 not n30052 ; n30052_not
g34171 not n23113 ; n23113_not
g34172 not n10423 ; n10423_not
g34173 not n25003 ; n25003_not
g34174 not n12601 ; n12601_not
g34175 not n30241 ; n30241_not
g34176 not n21052 ; n21052_not
g34177 not n11233 ; n11233_not
g34178 not n20206 ; n20206_not
g34179 not n24022 ; n24022_not
g34180 not n13420 ; n13420_not
g34181 not n22123 ; n22123_not
g34182 not n10162 ; n10162_not
g34183 not n12142 ; n12142_not
g34184 not n22321 ; n22321_not
g34185 not n10018 ; n10018_not
g34186 not n12043 ; n12043_not
g34187 not n25012 ; n25012_not
g34188 not n10333 ; n10333_not
g34189 not n11134 ; n11134_not
g34190 not n21700 ; n21700_not
g34191 not n10603 ; n10603_not
g34192 not n22033 ; n22033_not
g34193 not n21313 ; n21313_not
g34194 not n26002 ; n26002_not
g34195 not n20305 ; n20305_not
g34196 not n10180 ; n10180_not
g34197 not n11251 ; n11251_not
g34198 not n22411 ; n22411_not
g34199 not n30043 ; n30043_not
g34200 not n21412 ; n21412_not
g34201 not n21034 ; n21034_not
g34202 not n10360 ; n10360_not
g34203 not n26003 ; n26003_not
g34204 not n16211 ; n16211_not
g34205 not n11603 ; n11603_not
g34206 not n31304 ; n31304_not
g34207 not n20315 ; n20315_not
g34208 not n10235 ; n10235_not
g34209 not n11621 ; n11621_not
g34210 not n10424 ; n10424_not
g34211 not n30404 ; n30404_not
g34212 not n22232 ; n22232_not
g34213 not n23411 ; n23411_not
g34214 not n12134 ; n12134_not
g34215 not n30251 ; n30251_not
g34216 not n21035 ; n21035_not
g34217 not n10730 ; n10730_not
g34218 not n22115 ; n22115_not
g34219 not n20540 ; n20540_not
g34220 not n14051 ; n14051_not
g34221 not n30701 ; n30701_not
g34222 not n20630 ; n20630_not
g34223 not n21017 ; n21017_not
g34224 not n31115 ; n31115_not
g34225 not n26102 ; n26102_not
g34226 not n20423 ; n20423_not
g34227 not n15221 ; n15221_not
g34228 not n11522 ; n11522_not
g34229 not n30710 ; n30710_not
g34230 not n20900 ; n20900_not
g34231 not n11423 ; n11423_not
g34232 not n20207 ; n20207_not
g34233 not n20153 ; n20153_not
g34234 not n20810 ; n20810_not
g34235 not n23006 ; n23006_not
g34236 not n27020 ; n27020_not
g34237 not n21134 ; n21134_not
g34238 not n10262 ; n10262_not
g34239 not n22214 ; n22214_not
g34240 not n31331 ; n31331_not
g34241 not n11405 ; n11405_not
g34242 not n13610 ; n13610_not
g34243 not n10280 ; n10280_not
g34244 not n31700 ; n31700_not
g34245 not n31133 ; n31133_not
g34246 not n10712 ; n10712_not
g34247 not n10307 ; n10307_not
g34248 not n22016 ; n22016_not
g34249 not n21071 ; n21071_not
g34250 not n15005 ; n15005_not
g34251 not n21521 ; n21521_not
g34252 not n12035 ; n12035_not
g34253 not n22142 ; n22142_not
g34254 not n20504 ; n20504_not
g34255 not n21053 ; n21053_not
g34256 not n15032 ; n15032_not
g34257 not n24023 ; n24023_not
g34258 not n17120 ; n17120_not
g34259 not n30071 ; n30071_not
g34260 not n18011 ; n18011_not
g34261 not n11234 ; n11234_not
g34262 not n25004 ; n25004_not
g34263 not n24320 ; n24320_not
g34264 not n23123 ; n23123_not
g34265 not n10019 ; n10019_not
g34266 not n23132 ; n23132_not
g34267 not n11027 ; n11027_not
g34268 not n11225 ; n11225_not
g34269 not n17102 ; n17102_not
g34270 not n12341 ; n12341_not
g34271 not n25103 ; n25103_not
g34272 not n12323 ; n12323_not
g34273 not n13430 ; n13430_not
g34274 not n21431 ; n21431_not
g34275 not n24230 ; n24230_not
g34276 not n14123 ; n14123_not
g34277 not n32051 ; n32051_not
g34278 not n21341 ; n21341_not
g34279 not n22421 ; n22421_not
g34280 not n21314 ; n21314_not
g34281 not n10550 ; n10550_not
g34282 not n24203 ; n24203_not
g34283 not n17201 ; n17201_not
g34284 not n31052 ; n31052_not
g34285 not n10523 ; n10523_not
g34286 not n21602 ; n21602_not
g34287 not n21620 ; n21620_not
g34288 not n12503 ; n12503_not
g34289 not n11711 ; n11711_not
g34290 not n12305 ; n12305_not
g34291 not n22700 ; n22700_not
g34292 not n31016 ; n31016_not
g34293 not n14321 ; n14321_not
g34294 not n14303 ; n14303_not
g34295 not n11306 ; n11306_not
g34296 not n11441 ; n11441_not
g34297 not n19100 ; n19100_not
g34298 not n23015 ; n23015_not
g34299 not n24401 ; n24401_not
g34300 not n10613 ; n10613_not
g34301 not n10901 ; n10901_not
g34302 not n23051 ; n23051_not
g34303 not n30512 ; n30512_not
g34304 not n22610 ; n22610_not
g34305 not n30503 ; n30503_not
g34306 not n12611 ; n12611_not
g34307 not n14600 ; n14600_not
g34308 not n13322 ; n13322_not
g34309 not n31061 ; n31061_not
g34310 not n15203 ; n15203_not
g34311 not n28010 ; n28010_not
g34312 not n21260 ; n21260_not
g34313 not n30161 ; n30161_not
g34314 not n30431 ; n30431_not
g34315 not n23312 ; n23312_not
g34316 not n21242 ; n21242_not
g34317 not n10505 ; n10505_not
g34318 not n10145 ; n10145_not
g34319 not n10910 ; n10910_not
g34320 not n10163 ; n10163_not
g34321 not n10181 ; n10181_not
g34322 not n15401 ; n15401_not
g34323 not n21224 ; n21224_not
g34324 not n23402 ; n23402_not
g34325 not n27200 ; n27200_not
g34326 not n20234 ; n20234_not
g34327 not n22241 ; n22241_not
g34328 not n20252 ; n20252_not
g34329 not n10055 ; n10055_not
g34330 not n12233 ; n12233_not
g34331 not n13313 ; n13313_not
g34332 not n11720 ; n11720_not
g34333 not n20135 ; n20135_not
g34334 not n22160 ; n22160_not
g34335 not n31134 ; n31134_not
g34336 not n17400 ; n17400_not
g34337 not n21522 ; n21522_not
g34338 not n10416 ; n10416_not
g34339 not n24420 ; n24420_not
g34340 not n15222 ; n15222_not
g34341 not n31233 ; n31233_not
g34342 not n24204 ; n24204_not
g34343 not n10533 ; n10533_not
g34344 not n21225 ; n21225_not
g34345 not n30531 ; n30531_not
g34346 not n11109 ; n11109_not
g34347 not n17130 ; n17130_not
g34348 not n30342 ; n30342_not
g34349 not n11424 ; n11424_not
g34350 not n21324 ; n21324_not
g34351 not n21027 ; n21027_not
g34352 not n21207 ; n21207_not
g34353 not n17202 ; n17202_not
g34354 not n10470 ; n10470_not
g34355 not n11064 ; n11064_not
g34356 not n20811 ; n20811_not
g34357 not n12621 ; n12621_not
g34358 not n26031 ; n26031_not
g34359 not n30405 ; n30405_not
g34360 not n31341 ; n31341_not
g34361 not n30702 ; n30702_not
g34362 not n13503 ; n13503_not
g34363 not n31323 ; n31323_not
g34364 not n17013 ; n17013_not
g34365 not n10551 ; n10551_not
g34366 not n30414 ; n30414_not
g34367 not n21630 ; n21630_not
g34368 not n26040 ; n26040_not
g34369 not n21108 ; n21108_not
g34370 not n21351 ; n21351_not
g34371 not n21900 ; n21900_not
g34372 not n21261 ; n21261_not
g34373 not n25005 ; n25005_not
g34374 not n24330 ; n24330_not
g34375 not n11091 ; n11091_not
g34376 not n11226 ; n11226_not
g34377 not n25032 ; n25032_not
g34378 not n21405 ; n21405_not
g34379 not n30621 ; n30621_not
g34380 not n24033 ; n24033_not
g34381 not n25113 ; n25113_not
g34382 not n10380 ; n10380_not
g34383 not n12018 ; n12018_not
g34384 not n24240 ; n24240_not
g34385 not n11037 ; n11037_not
g34386 not n25410 ; n25410_not
g34387 not n30522 ; n30522_not
g34388 not n15411 ; n15411_not
g34389 not n21441 ; n21441_not
g34390 not n11307 ; n11307_not
g34391 not n10614 ; n10614_not
g34392 not n30504 ; n30504_not
g34393 not n31251 ; n31251_not
g34394 not n21801 ; n21801_not
g34395 not n21423 ; n21423_not
g34396 not n21720 ; n21720_not
g34397 not n21450 ; n21450_not
g34398 not n21243 ; n21243_not
g34399 not n12063 ; n12063_not
g34400 not n11802 ; n11802_not
g34401 not n21036 ; n21036_not
g34402 not n30441 ; n30441_not
g34403 not n13620 ; n13620_not
g34404 not n10128 ; n10128_not
g34405 not n14070 ; n14070_not
g34406 not n30810 ; n30810_not
g34407 not n13305 ; n13305_not
g34408 not n28011 ; n28011_not
g34409 not n10803 ; n10803_not
g34410 not n20154 ; n20154_not
g34411 not n14403 ; n14403_not
g34412 not n20145 ; n20145_not
g34413 not n23232 ; n23232_not
g34414 not n20136 ; n20136_not
g34415 not n14106 ; n14106_not
g34416 not n22152 ; n22152_not
g34417 not n12216 ; n12216_not
g34418 not n31062 ; n31062_not
g34419 not n13341 ; n13341_not
g34420 not n30144 ; n30144_not
g34421 not n11181 ; n11181_not
g34422 not n20280 ; n20280_not
g34423 not n23412 ; n23412_not
g34424 not n16230 ; n16230_not
g34425 not n27300 ; n27300_not
g34426 not n20262 ; n20262_not
g34427 not n10209 ; n10209_not
g34428 not n14052 ; n14052_not
g34429 not n20217 ; n20217_not
g34430 not n11208 ; n11208_not
g34431 not n10182 ; n10182_not
g34432 not n23025 ; n23025_not
g34433 not n10164 ; n10164_not
g34434 not n16104 ; n16104_not
g34435 not n10146 ; n10146_not
g34436 not n30180 ; n30180_not
g34437 not n23322 ; n23322_not
g34438 not n22602 ; n22602_not
g34439 not n11262 ; n11262_not
g34440 not n22611 ; n22611_not
g34441 not n29100 ; n29100_not
g34442 not n12333 ; n12333_not
g34443 not n31053 ; n31053_not
g34444 not n19110 ; n19110_not
g34445 not n14340 ; n14340_not
g34446 not n23007 ; n23007_not
g34447 not n31017 ; n31017_not
g34448 not n32106 ; n32106_not
g34449 not n30018 ; n30018_not
g34450 not n12315 ; n12315_not
g34451 not n19011 ; n19011_not
g34452 not n22431 ; n22431_not
g34453 not n10308 ; n10308_not
g34454 not n14250 ; n14250_not
g34455 not n22413 ; n22413_not
g34456 not n12270 ; n12270_not
g34457 not n22440 ; n22440_not
g34458 not n14124 ; n14124_not
g34459 not n32052 ; n32052_not
g34460 not n28200 ; n28200_not
g34461 not n12351 ; n12351_not
g34462 not n23142 ; n23142_not
g34463 not n10029 ; n10029_not
g34464 not n30126 ; n30126_not
g34465 not n30117 ; n30117_not
g34466 not n30081 ; n30081_not
g34467 not n22530 ; n22530_not
g34468 not n11244 ; n11244_not
g34469 not n12450 ; n12450_not
g34470 not n29001 ; n29001_not
g34471 not n11163 ; n11163_not
g34472 not n11532 ; n11532_not
g34473 not n30216 ; n30216_not
g34474 not n22206 ; n22206_not
g34475 not n10317 ; n10317_not
g34476 not n22170 ; n22170_not
g34477 not n11415 ; n11415_not
g34478 not n31530 ; n31530_not
g34479 not n15141 ; n15141_not
g34480 not n31611 ; n31611_not
g34481 not n15132 ; n15132_not
g34482 not n12162 ; n12162_not
g34483 not n10722 ; n10722_not
g34484 not n11127 ; n11127_not
g34485 not n10326 ; n10326_not
g34486 not n15114 ; n15114_not
g34487 not n20505 ; n20505_not
g34488 not n22134 ; n22134_not
g34489 not n20631 ; n20631_not
g34490 not n15105 ; n15105_not
g34491 not n10362 ; n10362_not
g34492 not n20604 ; n20604_not
g34493 not n12117 ; n12117_not
g34494 not n26310 ; n26310_not
g34495 not n20037 ; n20037_not
g34496 not n10731 ; n10731_not
g34497 not n31521 ; n31521_not
g34498 not n30720 ; n30720_not
g34499 not n11145 ; n11145_not
g34500 not n27201 ; n27201_not
g34501 not n26211 ; n26211_not
g34502 not n16212 ; n16212_not
g34503 not n20316 ; n20316_not
g34504 not n14034 ; n14034_not
g34505 not n18021 ; n18021_not
g34506 not n13422 ; n13422_not
g34507 not n20343 ; n20343_not
g34508 not n10245 ; n10245_not
g34509 not n23430 ; n23430_not
g34510 not n20235 ; n20235_not
g34511 not n20424 ; n20424_not
g34512 not n31701 ; n31701_not
g34513 not n10344 ; n10344_not
g34514 not n23511 ; n23511_not
g34515 not n20073 ; n20073_not
g34516 not n11550 ; n11550_not
g34517 not n10272 ; n10272_not
g34518 not n24016 ; n24016_not
g34519 not n30721 ; n30721_not
g34520 not n22531 ; n22531_not
g34521 not n10309 ; n10309_not
g34522 not n24502 ; n24502_not
g34523 not n13612 ; n13612_not
g34524 not n22423 ; n22423_not
g34525 not n24430 ; n24430_not
g34526 not n12613 ; n12613_not
g34527 not n22036 ; n22036_not
g34528 not n21613 ; n21613_not
g34529 not n24331 ; n24331_not
g34530 not n12604 ; n12604_not
g34531 not n14233 ; n14233_not
g34532 not n11551 ; n11551_not
g34533 not n24511 ; n24511_not
g34534 not n23026 ; n23026_not
g34535 not n16600 ; n16600_not
g34536 not n22630 ; n22630_not
g34537 not n10651 ; n10651_not
g34538 not n11452 ; n11452_not
g34539 not n22702 ; n22702_not
g34540 not n11803 ; n11803_not
g34541 not n22603 ; n22603_not
g34542 not n22612 ; n22612_not
g34543 not n22711 ; n22711_not
g34544 not n22072 ; n22072_not
g34545 not n23062 ; n23062_not
g34546 not n10642 ; n10642_not
g34547 not n22720 ; n22720_not
g34548 not n23008 ; n23008_not
g34549 not n24034 ; n24034_not
g34550 not n22180 ; n22180_not
g34551 not n23521 ; n23521_not
g34552 not n30820 ; n30820_not
g34553 not n22216 ; n22216_not
g34554 not n22306 ; n22306_not
g34555 not n11281 ; n11281_not
g34556 not n24160 ; n24160_not
g34557 not n24142 ; n24142_not
g34558 not n14323 ; n14323_not
g34559 not n31072 ; n31072_not
g34560 not n30622 ; n30622_not
g34561 not n17023 ; n17023_not
g34562 not n23431 ; n23431_not
g34563 not n10705 ; n10705_not
g34564 not n24115 ; n24115_not
g34565 not n22225 ; n22225_not
g34566 not n12703 ; n12703_not
g34567 not n11416 ; n11416_not
g34568 not n10804 ; n10804_not
g34569 not n23413 ; n23413_not
g34570 not n12730 ; n12730_not
g34571 not n31108 ; n31108_not
g34572 not n22522 ; n22522_not
g34573 not n16402 ; n16402_not
g34574 not n22324 ; n22324_not
g34575 not n23800 ; n23800_not
g34576 not n22504 ; n22504_not
g34577 not n23611 ; n23611_not
g34578 not n24313 ; n24313_not
g34579 not n22333 ; n22333_not
g34580 not n23152 ; n23152_not
g34581 not n22027 ; n22027_not
g34582 not n22342 ; n22342_not
g34583 not n22351 ; n22351_not
g34584 not n22360 ; n22360_not
g34585 not n23080 ; n23080_not
g34586 not n24214 ; n24214_not
g34587 not n23206 ; n23206_not
g34588 not n13720 ; n13720_not
g34589 not n10741 ; n10741_not
g34590 not n16330 ; n16330_not
g34591 not n10930 ; n10930_not
g34592 not n10723 ; n10723_not
g34593 not n21451 ; n21451_not
g34594 not n22162 ; n22162_not
g34595 not n22144 ; n22144_not
g34596 not n26131 ; n26131_not
g34597 not n20911 ; n20911_not
g34598 not n26104 ; n26104_not
g34599 not n20029 ; n20029_not
g34600 not n18220 ; n18220_not
g34601 not n28102 ; n28102_not
g34602 not n20263 ; n20263_not
g34603 not n15160 ; n15160_not
g34604 not n18211 ; n18211_not
g34605 not n20119 ; n20119_not
g34606 not n15142 ; n15142_not
g34607 not n20704 ; n20704_not
g34608 not n20650 ; n20650_not
g34609 not n12244 ; n12244_not
g34610 not n20641 ; n20641_not
g34611 not n14107 ; n14107_not
g34612 not n31522 ; n31522_not
g34613 not n11362 ; n11362_not
g34614 not n12082 ; n12082_not
g34615 not n11227 ; n11227_not
g34616 not n31171 ; n31171_not
g34617 not n12361 ; n12361_not
g34618 not n11623 ; n11623_not
g34619 not n18130 ; n18130_not
g34620 not n10417 ; n10417_not
g34621 not n26041 ; n26041_not
g34622 not n32035 ; n32035_not
g34623 not n11083 ; n11083_not
g34624 not n13513 ; n13513_not
g34625 not n21091 ; n21091_not
g34626 not n21064 ; n21064_not
g34627 not n12307 ; n12307_not
g34628 not n12046 ; n12046_not
g34629 not n11713 ; n11713_not
g34630 not n30361 ; n30361_not
g34631 not n21046 ; n21046_not
g34632 not n26113 ; n26113_not
g34633 not n30343 ; n30343_not
g34634 not n15241 ; n15241_not
g34635 not n10273 ; n10273_not
g34636 not n31720 ; n31720_not
g34637 not n10255 ; n10255_not
g34638 not n20353 ; n20353_not
g34639 not n27031 ; n27031_not
g34640 not n10138 ; n10138_not
g34641 not n27112 ; n27112_not
g34642 not n10147 ; n10147_not
g34643 not n31900 ; n31900_not
g34644 not n20290 ; n20290_not
g34645 not n27220 ; n27220_not
g34646 not n14035 ; n14035_not
g34647 not n12541 ; n12541_not
g34648 not n10219 ; n10219_not
g34649 not n27310 ; n27310_not
g34650 not n14053 ; n14053_not
g34651 not n20245 ; n20245_not
g34652 not n18112 ; n18112_not
g34653 not n13009 ; n13009_not
g34654 not n20137 ; n20137_not
g34655 not n12181 ; n12181_not
g34656 not n20533 ; n20533_not
g34657 not n30244 ; n30244_not
g34658 not n31531 ; n31531_not
g34659 not n31441 ; n31441_not
g34660 not n20506 ; n20506_not
g34661 not n12145 ; n12145_not
g34662 not n30154 ; n30154_not
g34663 not n20164 ; n20164_not
g34664 not n20470 ; n20470_not
g34665 not n28021 ; n28021_not
g34666 not n30235 ; n30235_not
g34667 not n12640 ; n12640_not
g34668 not n20452 ; n20452_not
g34669 not n20182 ; n20182_not
g34670 not n20434 ; n20434_not
g34671 not n30217 ; n30217_not
g34672 not n13306 ; n13306_not
g34673 not n14800 ; n14800_not
g34674 not n21109 ; n21109_not
g34675 not n19021 ; n19021_not
g34676 not n31162 ; n31162_not
g34677 not n11317 ; n11317_not
g34678 not n12532 ; n12532_not
g34679 not n15610 ; n15610_not
g34680 not n31180 ; n31180_not
g34681 not n30442 ; n30442_not
g34682 not n29200 ; n29200_not
g34683 not n32080 ; n32080_not
g34684 not n20632 ; n20632_not
g34685 not n12325 ; n12325_not
g34686 not n19210 ; n19210_not
g34687 not n12343 ; n12343_not
g34688 not n25114 ; n25114_not
g34689 not n21352 ; n21352_not
g34690 not n11038 ; n11038_not
g34691 not n24601 ; n24601_not
g34692 not n10453 ; n10453_not
g34693 not n11902 ; n11902_not
g34694 not n11344 ; n11344_not
g34695 not n11335 ; n11335_not
g34696 not n21550 ; n21550_not
g34697 not n11434 ; n11434_not
g34698 not n17221 ; n17221_not
g34699 not n21532 ; n21532_not
g34700 not n17230 ; n17230_not
g34701 not n30019 ; n30019_not
g34702 not n30541 ; n30541_not
g34703 not n10624 ; n10624_not
g34704 not n21028 ; n21028_not
g34705 not n30523 ; n30523_not
g34706 not n30037 ; n30037_not
g34707 not n22513 ; n22513_not
g34708 not n10552 ; n10552_not
g34709 not n15502 ; n15502_not
g34710 not n11047 ; n11047_not
g34711 not n25510 ; n25510_not
g34712 not n32062 ; n32062_not
g34713 not n25600 ; n25600_not
g34714 not n30082 ; n30082_not
g34715 not n15430 ; n15430_not
g34716 not n14161 ; n14161_not
g34717 not n30118 ; n30118_not
g34718 not n21226 ; n21226_not
g34719 not n10480 ; n10480_not
g34720 not n21217 ; n21217_not
g34721 not n17500 ; n17500_not
g34722 not n30127 ; n30127_not
g34723 not n29020 ; n29020_not
g34724 not n21334 ; n21334_not
g34725 not n15520 ; n15520_not
g34726 not n29002 ; n29002_not
g34727 not n12550 ; n12550_not
g34728 not n25132 ; n25132_not
g34729 not n22406 ; n22406_not
g34730 not n13082 ; n13082_not
g34731 not n20192 ; n20192_not
g34732 not n22136 ; n22136_not
g34733 not n19004 ; n19004_not
g34734 not n13424 ; n13424_not
g34735 not n13343 ; n13343_not
g34736 not n11282 ; n11282_not
g34737 not n11327 ; n11327_not
g34738 not n22712 ; n22712_not
g34739 not n10904 ; n10904_not
g34740 not n13370 ; n13370_not
g34741 not n18212 ; n18212_not
g34742 not n18104 ; n18104_not
g34743 not n13442 ; n13442_not
g34744 not n18140 ; n18140_not
g34745 not n11345 ; n11345_not
g34746 not n19310 ; n19310_not
g34747 not n32045 ; n32045_not
g34748 not n22631 ; n22631_not
g34749 not n16700 ; n16700_not
g34750 not n19130 ; n19130_not
g34751 not n22532 ; n22532_not
g34752 not n19103 ; n19103_not
g34753 not n13352 ; n13352_not
g34754 not n32018 ; n32018_not
g34755 not n13361 ; n13361_not
g34756 not n11363 ; n11363_not
g34757 not n19022 ; n19022_not
g34758 not n22208 ; n22208_not
g34759 not n13541 ; n13541_not
g34760 not n18203 ; n18203_not
g34761 not n11237 ; n11237_not
g34762 not n22415 ; n22415_not
g34763 not n22523 ; n22523_not
g34764 not n18230 ; n18230_not
g34765 not n19211 ; n19211_not
g34766 not n31181 ; n31181_not
g34767 not n21380 ; n21380_not
g34768 not n11057 ; n11057_not
g34769 not n20633 ; n20633_not
g34770 not n21425 ; n21425_not
g34771 not n21353 ; n21353_not
g34772 not n21812 ; n21812_not
g34773 not n21821 ; n21821_not
g34774 not n17060 ; n17060_not
g34775 not n11039 ; n11039_not
g34776 not n17411 ; n17411_not
g34777 not n21281 ; n21281_not
g34778 not n21911 ; n21911_not
g34779 not n21254 ; n21254_not
g34780 not n21920 ; n21920_not
g34781 not n17024 ; n17024_not
g34782 not n21236 ; n21236_not
g34783 not n21560 ; n21560_not
g34784 not n10481 ; n10481_not
g34785 not n17231 ; n17231_not
g34786 not n21641 ; n21641_not
g34787 not n21083 ; n21083_not
g34788 not n21461 ; n21461_not
g34789 not n17123 ; n17123_not
g34790 not n31163 ; n31163_not
g34791 not n21218 ; n21218_not
g34792 not n17213 ; n17213_not
g34793 not n17105 ; n17105_not
g34794 not n21713 ; n21713_not
g34795 not n31118 ; n31118_not
g34796 not n31514 ; n31514_not
g34797 not n20543 ; n20543_not
g34798 not n22109 ; n22109_not
g34799 not n11417 ; n11417_not
g34800 not n31532 ; n31532_not
g34801 not n22118 ; n22118_not
g34802 not n20471 ; n20471_not
g34803 not n21605 ; n21605_not
g34804 not n20462 ; n20462_not
g34805 not n22154 ; n22154_not
g34806 not n22172 ; n22172_not
g34807 not n31631 ; n31631_not
g34808 not n22190 ; n22190_not
g34809 not n31640 ; n31640_not
g34810 not n31811 ; n31811_not
g34811 not n18014 ; n18014_not
g34812 not n20336 ; n20336_not
g34813 not n20309 ; n20309_not
g34814 not n31901 ; n31901_not
g34815 not n20273 ; n20273_not
g34816 not n12902 ; n12902_not
g34817 not n17321 ; n17321_not
g34818 not n31172 ; n31172_not
g34819 not n21164 ; n21164_not
g34820 not n21146 ; n21146_not
g34821 not n21470 ; n21470_not
g34822 not n21137 ; n21137_not
g34823 not n21119 ; n21119_not
g34824 not n13190 ; n13190_not
g34825 not n22019 ; n22019_not
g34826 not n31127 ; n31127_not
g34827 not n21029 ; n21029_not
g34828 not n22055 ; n22055_not
g34829 not n20804 ; n20804_not
g34830 not n10922 ; n10922_not
g34831 not n20291 ; n20291_not
g34832 not n22082 ; n22082_not
g34833 not n20354 ; n20354_not
g34834 not n14009 ; n14009_not
g34835 not n12173 ; n12173_not
g34836 not n24323 ; n24323_not
g34837 not n24332 ; n24332_not
g34838 not n11804 ; n11804_not
g34839 not n30218 ; n30218_not
g34840 not n10652 ; n10652_not
g34841 not n11822 ; n11822_not
g34842 not n24404 ; n24404_not
g34843 not n11840 ; n11840_not
g34844 not n30236 ; n30236_not
g34845 not n24440 ; n24440_not
g34846 not n10382 ; n10382_not
g34847 not n13640 ; n13640_not
g34848 not n30164 ; n30164_not
g34849 not n10724 ; n10724_not
g34850 not n30173 ; n30173_not
g34851 not n11525 ; n11525_not
g34852 not n10157 ; n10157_not
g34853 not n14063 ; n14063_not
g34854 not n10175 ; n10175_not
g34855 not n11570 ; n11570_not
g34856 not n27500 ; n27500_not
g34857 not n27410 ; n27410_not
g34858 not n24035 ; n24035_not
g34859 not n27311 ; n27311_not
g34860 not n27230 ; n27230_not
g34861 not n11615 ; n11615_not
g34862 not n11471 ; n11471_not
g34863 not n27131 ; n27131_not
g34864 not n24170 ; n24170_not
g34865 not n11723 ; n11723_not
g34866 not n27014 ; n27014_not
g34867 not n10670 ; n10670_not
g34868 not n10274 ; n10274_not
g34869 not n15242 ; n15242_not
g34870 not n30443 ; n30443_not
g34871 not n25115 ; n25115_not
g34872 not n12074 ; n12074_not
g34873 not n30344 ; n30344_not
g34874 not n10562 ; n10562_not
g34875 not n30362 ; n30362_not
g34876 not n30434 ; n30434_not
g34877 not n15521 ; n15521_not
g34878 not n25430 ; n25430_not
g34879 not n13730 ; n13730_not
g34880 not n26042 ; n26042_not
g34881 not n25511 ; n25511_not
g34882 not n10139 ; n10139_not
g34883 not n10526 ; n10526_not
g34884 not n11633 ; n11633_not
g34885 not n10508 ; n10508_not
g34886 not n25034 ; n25034_not
g34887 not n13910 ; n13910_not
g34888 not n13532 ; n13532_not
g34889 not n10463 ; n10463_not
g34890 not n15080 ; n15080_not
g34891 not n12632 ; n12632_not
g34892 not n10634 ; n10634_not
g34893 not n30551 ; n30551_not
g34894 not n15107 ; n15107_not
g34895 not n15710 ; n15710_not
g34896 not n14603 ; n14603_not
g34897 not n15125 ; n15125_not
g34898 not n12506 ; n12506_not
g34899 not n24701 ; n24701_not
g34900 not n30542 ; n30542_not
g34901 not n15143 ; n15143_not
g34902 not n24800 ; n24800_not
g34903 not n15161 ; n15161_not
g34904 not n15170 ; n15170_not
g34905 not n25016 ; n25016_not
g34906 not n15215 ; n15215_not
g34907 not n25052 ; n25052_not
g34908 not n26114 ; n26114_not
g34909 not n29003 ; n29003_not
g34910 not n12380 ; n12380_not
g34911 not n16340 ; n16340_not
g34912 not n16331 ; n16331_not
g34913 not n23225 ; n23225_not
g34914 not n16313 ; n16313_not
g34915 not n30137 ; n30137_not
g34916 not n12353 ; n12353_not
g34917 not n30830 ; n30830_not
g34918 not n23243 ; n23243_not
g34919 not n12335 ; n12335_not
g34920 not n28202 ; n28202_not
g34921 not n30821 ; n30821_not
g34922 not n10346 ; n10346_not
g34923 not n12317 ; n12317_not
g34924 not n16250 ; n16250_not
g34925 not n28130 ; n28130_not
g34926 not n11741 ; n11741_not
g34927 not n28103 ; n28103_not
g34928 not n12281 ; n12281_not
g34929 not n12263 ; n12263_not
g34930 not n28040 ; n28040_not
g34931 not n16223 ; n16223_not
g34932 not n16205 ; n16205_not
g34933 not n14252 ; n14252_not
g34934 not n14243 ; n14243_not
g34935 not n14270 ; n14270_not
g34936 not n10832 ; n10832_not
g34937 not n14234 ; n14234_not
g34938 not n16502 ; n16502_not
g34939 not n23009 ; n23009_not
g34940 not n14333 ; n14333_not
g34941 not n22442 ; n22442_not
g34942 not n23027 ; n23027_not
g34943 not n30038 ; n30038_not
g34944 not n29201 ; n29201_not
g34945 not n16403 ; n16403_not
g34946 not n14360 ; n14360_not
g34947 not n23081 ; n23081_not
g34948 not n16421 ; n16421_not
g34949 not n23108 ; n23108_not
g34950 not n12371 ; n12371_not
g34951 not n23126 ; n23126_not
g34952 not n30902 ; n30902_not
g34953 not n23153 ; n23153_not
g34954 not n10814 ; n10814_not
g34955 not n29021 ; n29021_not
g34956 not n23522 ; n23522_not
g34957 not n14108 ; n14108_not
g34958 not n10067 ; n10067_not
g34959 not n10085 ; n10085_not
g34960 not n14612 ; n14612_not
g34961 not n23360 ; n23360_not
g34962 not n14621 ; n14621_not
g34963 not n11507 ; n11507_not
g34964 not n30731 ; n30731_not
g34965 not n28022 ; n28022_not
g34966 not n28004 ; n28004_not
g34967 not n23810 ; n23810_not
g34968 not n14090 ; n14090_not
g34969 not n14117 ; n14117_not
g34970 not n23504 ; n23504_not
g34971 not n10058 ; n10058_not
g34972 not n15243 ; n15243_not
g34973 not n13353 ; n13353_not
g34974 not n27501 ; n27501_not
g34975 not n28221 ; n28221_not
g34976 not n29202 ; n29202_not
g34977 not n29220 ; n29220_not
g34978 not n14343 ; n14343_not
g34979 not n14730 ; n14730_not
g34980 not n21039 ; n21039_not
g34981 not n12057 ; n12057_not
g34982 not n13083 ; n13083_not
g34983 not n20409 ; n20409_not
g34984 not n19032 ; n19032_not
g34985 not n26061 ; n26061_not
g34986 not n10248 ; n10248_not
g34987 not n28023 ; n28023_not
g34988 not n26115 ; n26115_not
g34989 not n31344 ; n31344_not
g34990 not n31353 ; n31353_not
g34991 not n10086 ; n10086_not
g34992 not n13614 ; n13614_not
g34993 not n14028 ; n14028_not
g34994 not n13605 ; n13605_not
g34995 not n15225 ; n15225_not
g34996 not n19140 ; n19140_not
g34997 not n11292 ; n11292_not
g34998 not n14361 ; n14361_not
g34999 not n10194 ; n10194_not
g35000 not n26106 ; n26106_not
g35001 not n30039 ; n30039_not
g35002 not n20814 ; n20814_not
g35003 not n14235 ; n14235_not
g35004 not n11328 ; n11328_not
g35005 not n20175 ; n20175_not
g35006 not n20706 ; n20706_not
g35007 not n11634 ; n11634_not
g35008 not n20382 ; n20382_not
g35009 not n30165 ; n30165_not
g35010 not n13902 ; n13902_not
g35011 not n21147 ; n21147_not
g35012 not n18150 ; n18150_not
g35013 not n10446 ; n10446_not
g35014 not n21165 ; n21165_not
g35015 not n15306 ; n15306_not
g35016 not n18600 ; n18600_not
g35017 not n14910 ; n14910_not
g35018 not n17511 ; n17511_not
g35019 not n11346 ; n11346_not
g35020 not n30363 ; n30363_not
g35021 not n30381 ; n30381_not
g35022 not n21084 ; n21084_not
g35023 not n14145 ; n14145_not
g35024 not n11427 ; n11427_not
g35025 not n12255 ; n12255_not
g35026 not n20364 ; n20364_not
g35027 not n30390 ; n30390_not
g35028 not n13821 ; n13821_not
g35029 not n11364 ; n11364_not
g35030 not n12660 ; n12660_not
g35031 not n17601 ; n17601_not
g35032 not n20391 ; n20391_not
g35033 not n14280 ; n14280_not
g35034 not n21129 ; n21129_not
g35035 not n13911 ; n13911_not
g35036 not n13371 ; n13371_not
g35037 not n27051 ; n27051_not
g35038 not n27132 ; n27132_not
g35039 not n18042 ; n18042_not
g35040 not n30237 ; n30237_not
g35041 not n12345 ; n12345_not
g35042 not n26610 ; n26610_not
g35043 not n27024 ; n27024_not
g35044 not n20526 ; n20526_not
g35045 not n14820 ; n14820_not
g35046 not n10068 ; n10068_not
g35047 not n12363 ; n12363_not
g35048 not n26340 ; n26340_not
g35049 not n13407 ; n13407_not
g35050 not n13326 ; n13326_not
g35051 not n30057 ; n30057_not
g35052 not n28410 ; n28410_not
g35053 not n12291 ; n12291_not
g35054 not n22542 ; n22542_not
g35055 not n20445 ; n20445_not
g35056 not n14127 ; n14127_not
g35057 not n14514 ; n14514_not
g35058 not n12309 ; n12309_not
g35059 not n11049 ; n11049_not
g35060 not n13290 ; n13290_not
g35061 not n30192 ; n30192_not
g35062 not n12156 ; n12156_not
g35063 not n27105 ; n27105_not
g35064 not n18024 ; n18024_not
g35065 not n11391 ; n11391_not
g35066 not n12327 ; n12327_not
g35067 not n20481 ; n20481_not
g35068 not n27150 ; n27150_not
g35069 not n14604 ; n14604_not
g35070 not n26250 ; n26250_not
g35071 not n10338 ; n10338_not
g35072 not n27411 ; n27411_not
g35073 not n20328 ; n20328_not
g35074 not n27420 ; n27420_not
g35075 not n26241 ; n26241_not
g35076 not n20724 ; n20724_not
g35077 not n12372 ; n12372_not
g35078 not n20238 ; n20238_not
g35079 not n29022 ; n29022_not
g35080 not n20193 ; n20193_not
g35081 not n19302 ; n19302_not
g35082 not n18105 ; n18105_not
g35083 not n15180 ; n15180_not
g35084 not n29040 ; n29040_not
g35085 not n19212 ; n19212_not
g35086 not n13074 ; n13074_not
g35087 not n20292 ; n20292_not
g35088 not n30327 ; n30327_not
g35089 not n31452 ; n31452_not
g35090 not n31416 ; n31416_not
g35091 not n27213 ; n27213_not
g35092 not n32073 ; n32073_not
g35093 not n10293 ; n10293_not
g35094 not n20625 ; n20625_not
g35095 not n19050 ; n19050_not
g35096 not n20634 ; n20634_not
g35097 not n19410 ; n19410_not
g35098 not n27231 ; n27231_not
g35099 not n20544 ; n20544_not
g35100 not n20463 ; n20463_not
g35101 not n30183 ; n30183_not
g35102 not n18213 ; n18213_not
g35103 not n11472 ; n11472_not
g35104 not n21435 ; n21435_not
g35105 not n11742 ; n11742_not
g35106 not n10671 ; n10671_not
g35107 not n15900 ; n15900_not
g35108 not n21903 ; n21903_not
g35109 not n31137 ; n31137_not
g35110 not n24144 ; n24144_not
g35111 not n24135 ; n24135_not
g35112 not n24108 ; n24108_not
g35113 not n21651 ; n21651_not
g35114 not n11562 ; n11562_not
g35115 not n30633 ; n30633_not
g35116 not n21471 ; n21471_not
g35117 not n24081 ; n24081_not
g35118 not n30660 ; n30660_not
g35119 not n11580 ; n11580_not
g35120 not n12741 ; n12741_not
g35121 not n24009 ; n24009_not
g35122 not n31119 ; n31119_not
g35123 not n23730 ; n23730_not
g35124 not n22065 ; n22065_not
g35125 not n11544 ; n11544_not
g35126 not n23901 ; n23901_not
g35127 not n17214 ; n17214_not
g35128 not n17205 ; n17205_not
g35129 not n24621 ; n24621_not
g35130 not n30570 ; n30570_not
g35131 not n10635 ; n10635_not
g35132 not n22506 ; n22506_not
g35133 not n10509 ; n10509_not
g35134 not n24324 ; n24324_not
g35135 not n24405 ; n24405_not
g35136 not n21606 ; n21606_not
g35137 not n17151 ; n17151_not
g35138 not n17133 ; n17133_not
g35139 not n24360 ; n24360_not
g35140 not n24342 ; n24342_not
g35141 not n21660 ; n21660_not
g35142 not n21705 ; n21705_not
g35143 not n10653 ; n10653_not
g35144 not n24306 ; n24306_not
g35145 not n24270 ; n24270_not
g35146 not n21732 ; n21732_not
g35147 not n24252 ; n24252_not
g35148 not n24243 ; n24243_not
g35149 not n24225 ; n24225_not
g35150 not n21804 ; n21804_not
g35151 not n16332 ; n16332_not
g35152 not n22425 ; n22425_not
g35153 not n30903 ; n30903_not
g35154 not n23190 ; n23190_not
g35155 not n23172 ; n23172_not
g35156 not n23163 ; n23163_not
g35157 not n23118 ; n23118_not
g35158 not n16413 ; n16413_not
g35159 not n30930 ; n30930_not
g35160 not n23091 ; n23091_not
g35161 not n10824 ; n10824_not
g35162 not n23055 ; n23055_not
g35163 not n23028 ; n23028_not
g35164 not n22632 ; n22632_not
g35165 not n22650 ; n22650_not
g35166 not n23019 ; n23019_not
g35167 not n22920 ; n22920_not
g35168 not n16503 ; n16503_not
g35169 not n22902 ; n22902_not
g35170 not n16512 ; n16512_not
g35171 not n22713 ; n22713_not
g35172 not n31029 ; n31029_not
g35173 not n10851 ; n10851_not
g35174 not n16530 ; n16530_not
g35175 not n11517 ; n11517_not
g35176 not n23712 ; n23712_not
g35177 not n10734 ; n10734_not
g35178 not n22470 ; n22470_not
g35179 not n22146 ; n22146_not
g35180 not n23550 ; n23550_not
g35181 not n22182 ; n22182_not
g35182 not n23154 ; n23154_not
g35183 not n23523 ; n23523_not
g35184 not n23451 ; n23451_not
g35185 not n23424 ; n23424_not
g35186 not n16215 ; n16215_not
g35187 not n16233 ; n16233_not
g35188 not n23406 ; n23406_not
g35189 not n23208 ; n23208_not
g35190 not n23370 ; n23370_not
g35191 not n23361 ; n23361_not
g35192 not n22461 ; n22461_not
g35193 not n23325 ; n23325_not
g35194 not n13731 ; n13731_not
g35195 not n13740 ; n13740_not
g35196 not n23244 ; n23244_not
g35197 not n22164 ; n22164_not
g35198 not n16314 ; n16314_not
g35199 not n23226 ; n23226_not
g35200 not n25125 ; n25125_not
g35201 not n21372 ; n21372_not
g35202 not n24702 ; n24702_not
g35203 not n21381 ; n21381_not
g35204 not n10428 ; n10428_not
g35205 not n31182 ; n31182_not
g35206 not n15603 ; n15603_not
g35207 not n17106 ; n17106_not
g35208 not n15621 ; n15621_not
g35209 not n21417 ; n21417_not
g35210 not n21273 ; n21273_not
g35211 not n24531 ; n24531_not
g35212 not n17250 ; n17250_not
g35213 not n12651 ; n12651_not
g35214 not n24810 ; n24810_not
g35215 not n31155 ; n31155_not
g35216 not n10617 ; n10617_not
g35217 not n25710 ; n25710_not
g35218 not n31173 ; n31173_not
g35219 not n15090 ; n15090_not
g35220 not n21219 ; n21219_not
g35221 not n10491 ; n10491_not
g35222 not n15117 ; n15117_not
g35223 not n15423 ; n15423_not
g35224 not n25620 ; n25620_not
g35225 not n25512 ; n25512_not
g35226 not n20670 ; n20670_not
g35227 not n10536 ; n10536_not
g35228 not n25440 ; n25440_not
g35229 not n17412 ; n17412_not
g35230 not n21309 ; n21309_not
g35231 not n17403 ; n17403_not
g35232 not n31191 ; n31191_not
g35233 not n25242 ; n25242_not
g35234 not n21327 ; n21327_not
g35235 not n15450 ; n15450_not
g35236 not n25215 ; n25215_not
g35237 not n14136 ; n14136_not
g35238 not n12624 ; n12624_not
g35239 not n21543 ; n21543_not
g35240 not n24604 ; n24604_not
g35241 not n10807 ; n10807_not
g35242 not n26053 ; n26053_not
g35243 not n22192 ; n22192_not
g35244 not n20572 ; n20572_not
g35245 not n26323 ; n26323_not
g35246 not n28231 ; n28231_not
g35247 not n22156 ; n22156_not
g35248 not n23227 ; n23227_not
g35249 not n26035 ; n26035_not
g35250 not n30094 ; n30094_not
g35251 not n28330 ; n28330_not
g35252 not n25054 ; n25054_not
g35253 not n30076 ; n30076_not
g35254 not n30058 ; n30058_not
g35255 not n26008 ; n26008_not
g35256 not n32065 ; n32065_not
g35257 not n22417 ; n22417_not
g35258 not n11059 ; n11059_not
g35259 not n21274 ; n21274_not
g35260 not n19600 ; n19600_not
g35261 not n25270 ; n25270_not
g35262 not n26071 ; n26071_not
g35263 not n23542 ; n23542_not
g35264 not n30283 ; n30283_not
g35265 not n23155 ; n23155_not
g35266 not n22174 ; n22174_not
g35267 not n10285 ; n10285_not
g35268 not n21319 ; n21319_not
g35269 not n28060 ; n28060_not
g35270 not n25315 ; n25315_not
g35271 not n21571 ; n21571_not
g35272 not n20554 ; n20554_not
g35273 not n10915 ; n10915_not
g35274 not n20086 ; n20086_not
g35275 not n30274 ; n30274_not
g35276 not n10906 ; n10906_not
g35277 not n21094 ; n21094_not
g35278 not n30382 ; n30382_not
g35279 not n23326 ; n23326_not
g35280 not n22246 ; n22246_not
g35281 not n22291 ; n22291_not
g35282 not n30580 ; n30580_not
g35283 not n22453 ; n22453_not
g35284 not n19060 ; n19060_not
g35285 not n30328 ; n30328_not
g35286 not n29320 ; n29320_not
g35287 not n25702 ; n25702_not
g35288 not n31435 ; n31435_not
g35289 not n22651 ; n22651_not
g35290 not n21166 ; n21166_not
g35291 not n22930 ; n22930_not
g35292 not n10456 ; n10456_not
g35293 not n25711 ; n25711_not
g35294 not n21193 ; n21193_not
g35295 not n31264 ; n31264_not
g35296 not n11329 ; n11329_not
g35297 not n22732 ; n22732_not
g35298 not n18250 ; n18250_not
g35299 not n10870 ; n10870_not
g35300 not n20617 ; n20617_not
g35301 not n10861 ; n10861_not
g35302 not n20626 ; n20626_not
g35303 not n22444 ; n22444_not
g35304 not n10519 ; n10519_not
g35305 not n31507 ; n31507_not
g35306 not n22480 ; n22480_not
g35307 not n22921 ; n22921_not
g35308 not n22516 ; n22516_not
g35309 not n19303 ; n19303_not
g35310 not n30931 ; n30931_not
g35311 not n23119 ; n23119_not
g35312 not n31462 ; n31462_not
g35313 not n25630 ; n25630_not
g35314 not n29041 ; n29041_not
g35315 not n22543 ; n22543_not
g35316 not n22570 ; n22570_not
g35317 not n21229 ; n21229_not
g35318 not n25018 ; n25018_not
g35319 not n23065 ; n23065_not
g35320 not n24640 ; n24640_not
g35321 not n22615 ; n22615_not
g35322 not n21148 ; n21148_not
g35323 not n10825 ; n10825_not
g35324 not n29221 ; n29221_not
g35325 not n29311 ; n29311_not
g35326 not n30517 ; n30517_not
g35327 not n21634 ; n21634_not
g35328 not n31804 ; n31804_not
g35329 not n21850 ; n21850_not
g35330 not n27034 ; n27034_not
g35331 not n27061 ; n27061_not
g35332 not n24433 ; n24433_not
g35333 not n24190 ; n24190_not
g35334 not n31138 ; n31138_not
g35335 not n24181 ; n24181_not
g35336 not n27115 ; n27115_not
g35337 not n30337 ; n30337_not
g35338 not n20329 ; n20329_not
g35339 not n21364 ; n21364_not
g35340 not n20662 ; n20662_not
g35341 not n21616 ; n21616_not
g35342 not n24118 ; n24118_not
g35343 not n26422 ; n26422_not
g35344 not n24811 ; n24811_not
g35345 not n24091 ; n24091_not
g35346 not n26107 ; n26107_not
g35347 not n10537 ; n10537_not
g35348 not n24712 ; n24712_not
g35349 not n24730 ; n24730_not
g35350 not n24325 ; n24325_not
g35351 not n20518 ; n20518_not
g35352 not n24271 ; n24271_not
g35353 not n26521 ; n26521_not
g35354 not n26800 ; n26800_not
g35355 not n21481 ; n21481_not
g35356 not n21751 ; n21751_not
g35357 not n24253 ; n24253_not
g35358 not n10429 ; n10429_not
g35359 not n31714 ; n31714_not
g35360 not n20464 ; n20464_not
g35361 not n24235 ; n24235_not
g35362 not n20392 ; n20392_not
g35363 not n26224 ; n26224_not
g35364 not n24415 ; n24415_not
g35365 not n10267 ; n10267_not
g35366 not n20374 ; n20374_not
g35367 not n31732 ; n31732_not
g35368 not n21436 ; n21436_not
g35369 not n27007 ; n27007_not
g35370 not n26116 ; n26116_not
g35371 not n23911 ; n23911_not
g35372 not n25072 ; n25072_not
g35373 not n24622 ; n24622_not
g35374 not n30715 ; n30715_not
g35375 not n22093 ; n22093_not
g35376 not n21490 ; n21490_not
g35377 not n25108 ; n25108_not
g35378 not n23821 ; n23821_not
g35379 not n23740 ; n23740_not
g35380 not n10087 ; n10087_not
g35381 not n10636 ; n10636_not
g35382 not n21346 ; n21346_not
g35383 not n25126 ; n25126_not
g35384 not n22138 ; n22138_not
g35385 not n30265 ; n30265_not
g35386 not n28033 ; n28033_not
g35387 not n23443 ; n23443_not
g35388 not n21535 ; n21535_not
g35389 not n23551 ; n23551_not
g35390 not n25801 ; n25801_not
g35391 not n10069 ; n10069_not
g35392 not n30724 ; n30724_not
g35393 not n24505 ; n24505_not
g35394 not n24523 ; n24523_not
g35395 not n27232 ; n27232_not
g35396 not n30184 ; n30184_not
g35397 not n30634 ; n30634_not
g35398 not n20266 ; n20266_not
g35399 not n10708 ; n10708_not
g35400 not n31921 ; n31921_not
g35401 not n27412 ; n27412_not
g35402 not n20248 ; n20248_not
g35403 not n30643 ; n30643_not
g35404 not n24028 ; n24028_not
g35405 not n27430 ; n27430_not
g35406 not n31354 ; n31354_not
g35407 not n21382 ; n21382_not
g35408 not n10627 ; n10627_not
g35409 not n20644 ; n20644_not
g35410 not n31192 ; n31192_not
g35411 not n22048 ; n22048_not
g35412 not n23704 ; n23704_not
g35413 not n27502 ; n27502_not
g35414 not n10195 ; n10195_not
g35415 not n31417 ; n31417_not
g35416 not n14443 ; n14443_not
g35417 not n15811 ; n15811_not
g35418 not n13543 ; n13543_not
g35419 not n17053 ; n17053_not
g35420 not n16171 ; n16171_not
g35421 not n18007 ; n18007_not
g35422 not n17116 ; n17116_not
g35423 not n14029 ; n14029_not
g35424 not n11806 ; n11806_not
g35425 not n14083 ; n14083_not
g35426 not n11617 ; n11617_not
g35427 not n13291 ; n13291_not
g35428 not n16090 ; n16090_not
g35429 not n17161 ; n17161_not
g35430 not n14137 ; n14137_not
g35431 not n17404 ; n17404_not
g35432 not n12490 ; n12490_not
g35433 not n17224 ; n17224_not
g35434 not n13633 ; n13633_not
g35435 not n13426 ; n13426_not
g35436 not n11086 ; n11086_not
g35437 not n11482 ; n11482_not
g35438 not n12319 ; n12319_not
g35439 not n13912 ; n13912_not
g35440 not n15181 ; n15181_not
g35441 not n13516 ; n13516_not
g35442 not n12337 ; n12337_not
g35443 not n18151 ; n18151_not
g35444 not n18133 ; n18133_not
g35445 not n18115 ; n18115_not
g35446 not n12373 ; n12373_not
g35447 not n13930 ; n13930_not
g35448 not n14461 ; n14461_not
g35449 not n13660 ; n13660_not
g35450 not n12616 ; n12616_not
g35451 not n14434 ; n14434_not
g35452 not n18052 ; n18052_not
g35453 not n14263 ; n14263_not
g35454 not n10924 ; n10924_not
g35455 not n15901 ; n15901_not
g35456 not n11554 ; n11554_not
g35457 not n15433 ; n15433_not
g35458 not n14344 ; n14344_not
g35459 not n14317 ; n14317_not
g35460 not n15028 ; n15028_not
g35461 not n12139 ; n12139_not
g35462 not n15118 ; n15118_not
g35463 not n11563 ; n11563_not
g35464 not n15091 ; n15091_not
g35465 not n14128 ; n14128_not
g35466 not n16009 ; n16009_not
g35467 not n15613 ; n15613_not
g35468 not n14281 ; n14281_not
g35469 not n17710 ; n17710_not
g35470 not n11608 ; n11608_not
g35471 not n13318 ; n13318_not
g35472 not n15154 ; n15154_not
g35473 not n13642 ; n13642_not
g35474 not n17260 ; n17260_not
g35475 not n11770 ; n11770_not
g35476 not n17134 ; n17134_not
g35477 not n12355 ; n12355_not
g35478 not n17332 ; n17332_not
g35479 not n12544 ; n12544_not
g35480 not n15631 ; n15631_not
g35481 not n15136 ; n15136_not
g35482 not n17350 ; n17350_not
g35483 not n13174 ; n13174_not
g35484 not n11518 ; n11518_not
g35485 not n13606 ; n13606_not
g35486 not n13183 ; n13183_not
g35487 not n17413 ; n17413_not
g35488 not n17422 ; n17422_not
g35489 not n11752 ; n11752_not
g35490 not n17440 ; n17440_not
g35491 not n14245 ; n14245_not
g35492 not n12670 ; n12670_not
g35493 not n15514 ; n15514_not
g35494 not n14605 ; n14605_not
g35495 not n13507 ; n13507_not
g35496 not n16315 ; n16315_not
g35497 not n12643 ; n12643_not
g35498 not n12517 ; n12517_not
g35499 not n14632 ; n14632_not
g35500 not n13732 ; n13732_not
g35501 not n13480 ; n13480_not
g35502 not n13750 ; n13750_not
g35503 not n13327 ; n13327_not
g35504 not n14641 ; n14641_not
g35505 not n11860 ; n11860_not
g35506 not n16621 ; n16621_not
g35507 not n16603 ; n16603_not
g35508 not n18331 ; n18331_not
g35509 not n14803 ; n14803_not
g35510 not n12454 ; n12454_not
g35511 not n12742 ; n12742_not
g35512 not n18025 ; n18025_not
g35513 not n16414 ; n16414_not
g35514 not n11941 ; n11941_not
g35515 not n14713 ; n14713_not
g35516 not n11653 ; n11653_not
g35517 not n14452 ; n14452_not
g35518 not n16513 ; n16513_not
g35519 not n14731 ; n14731_not
g35520 not n13336 ; n13336_not
g35521 not n14740 ; n14740_not
g35522 not n12229 ; n12229_not
g35523 not n18241 ; n18241_not
g35524 not n12238 ; n12238_not
g35525 not n11932 ; n11932_not
g35526 not n16216 ; n16216_not
g35527 not n15226 ; n15226_not
g35528 not n18232 ; n18232_not
g35529 not n16234 ; n16234_not
g35530 not n14821 ; n14821_not
g35531 not n30059 ; n30059_not
g35532 not n12068 ; n12068_not
g35533 not n20609 ; n20609_not
g35534 not n18053 ; n18053_not
g35535 not n24218 ; n24218_not
g35536 not n15128 ; n15128_not
g35537 not n30716 ; n30716_not
g35538 not n12752 ; n12752_not
g35539 not n14228 ; n14228_not
g35540 not n22625 ; n22625_not
g35541 not n30653 ; n30653_not
g35542 not n30644 ; n30644_not
g35543 not n12581 ; n12581_not
g35544 not n20627 ; n20627_not
g35545 not n12293 ; n12293_not
g35546 not n15146 ; n15146_not
g35547 not n30464 ; n30464_not
g35548 not n13805 ; n13805_not
g35549 not n30419 ; n30419_not
g35550 not n30374 ; n30374_not
g35551 not n24236 ; n24236_not
g35552 not n12734 ; n12734_not
g35553 not n11357 ; n11357_not
g35554 not n30275 ; n30275_not
g35555 not n11249 ; n11249_not
g35556 not n26054 ; n26054_not
g35557 not n23642 ; n23642_not
g35558 not n24092 ; n24092_not
g35559 not n10691 ; n10691_not
g35560 not n30428 ; n30428_not
g35561 not n15092 ; n15092_not
g35562 not n24119 ; n24119_not
g35563 not n20825 ; n20825_not
g35564 not n24650 ; n24650_not
g35565 not n12635 ; n12635_not
g35566 not n19412 ; n19412_not
g35567 not n26306 ; n26306_not
g35568 not n20249 ; n20249_not
g35569 not n11654 ; n11654_not
g35570 not n26072 ; n26072_not
g35571 not n26270 ; n26270_not
g35572 not n18206 ; n18206_not
g35573 not n26261 ; n26261_not
g35574 not n24191 ; n24191_not
g35575 not n30815 ; n30815_not
g35576 not n26126 ; n26126_not
g35577 not n26081 ; n26081_not
g35578 not n11735 ; n11735_not
g35579 not n30761 ; n30761_not
g35580 not n26090 ; n26090_not
g35581 not n24335 ; n24335_not
g35582 not n13940 ; n13940_not
g35583 not n20393 ; n20393_not
g35584 not n24380 ; n24380_not
g35585 not n20375 ; n20375_not
g35586 not n11168 ; n11168_not
g35587 not n20357 ; n20357_not
g35588 not n18242 ; n18242_not
g35589 not n26117 ; n26117_not
g35590 not n30266 ; n30266_not
g35591 not n20339 ; n20339_not
g35592 not n12608 ; n12608_not
g35593 not n18035 ; n18035_not
g35594 not n26162 ; n26162_not
g35595 not n13931 ; n13931_not
g35596 not n30284 ; n30284_not
g35597 not n15812 ; n15812_not
g35598 not n13652 ; n13652_not
g35599 not n10646 ; n10646_not
g35600 not n22850 ; n22850_not
g35601 not n20276 ; n20276_not
g35602 not n11186 ; n11186_not
g35603 not n24425 ; n24425_not
g35604 not n11384 ; n11384_not
g35605 not n15236 ; n15236_not
g35606 not n30329 ; n30329_not
g35607 not n30581 ; n30581_not
g35608 not n30383 ; n30383_not
g35609 not n20591 ; n20591_not
g35610 not n28223 ; n28223_not
g35611 not n24470 ; n24470_not
g35612 not n11780 ; n11780_not
g35613 not n24254 ; n24254_not
g35614 not n20168 ; n20168_not
g35615 not n30077 ; n30077_not
g35616 not n20564 ; n20564_not
g35617 not n26234 ; n26234_not
g35618 not n24452 ; n24452_not
g35619 not n14138 ; n14138_not
g35620 not n18152 ; n18152_not
g35621 not n26108 ; n26108_not
g35622 not n12509 ; n12509_not
g35623 not n24272 ; n24272_not
g35624 not n20519 ; n20519_not
g35625 not n18143 ; n18143_not
g35626 not n15164 ; n15164_not
g35627 not n10664 ; n10664_not
g35628 not n20474 ; n20474_not
g35629 not n30536 ; n30536_not
g35630 not n26207 ; n26207_not
g35631 not n20438 ; n20438_not
g35632 not n30518 ; n30518_not
g35633 not n30356 ; n30356_not
g35634 not n16262 ; n16262_not
g35635 not n27170 ; n27170_not
g35636 not n10916 ; n10916_not
g35637 not n11726 ; n11726_not
g35638 not n13580 ; n13580_not
g35639 not n22274 ; n22274_not
g35640 not n14822 ; n14822_not
g35641 not n22292 ; n22292_not
g35642 not n23273 ; n23273_not
g35643 not n14039 ; n14039_not
g35644 not n22184 ; n22184_not
g35645 not n28061 ; n28061_not
g35646 not n27206 ; n27206_not
g35647 not n22148 ; n22148_not
g35648 not n16730 ; n16730_not
g35649 not n22409 ; n22409_not
g35650 not n14624 ; n14624_not
g35651 not n27035 ; n27035_not
g35652 not n27062 ; n27062_not
g35653 not n23192 ; n23192_not
g35654 not n23444 ; n23444_not
g35655 not n27116 ; n27116_not
g35656 not n12653 ; n12653_not
g35657 not n16244 ; n16244_not
g35658 not n22076 ; n22076_not
g35659 not n21491 ; n21491_not
g35660 not n14516 ; n14516_not
g35661 not n28250 ; n28250_not
g35662 not n21563 ; n21563_not
g35663 not n27143 ; n27143_not
g35664 not n12347 ; n12347_not
g35665 not n22166 ; n22166_not
g35666 not n23345 ; n23345_not
g35667 not n12329 ; n12329_not
g35668 not n28205 ; n28205_not
g35669 not n27242 ; n27242_not
g35670 not n22931 ; n22931_not
g35671 not n22706 ; n22706_not
g35672 not n16415 ; n16415_not
g35673 not n10817 ; n10817_not
g35674 not n22733 ; n22733_not
g35675 not n10880 ; n10880_not
g35676 not n16541 ; n16541_not
g35677 not n22427 ; n22427_not
g35678 not n23048 ; n23048_not
g35679 not n22382 ; n22382_not
g35680 not n27602 ; n27602_not
g35681 not n16523 ; n16523_not
g35682 not n14714 ; n14714_not
g35683 not n16460 ; n16460_not
g35684 not n16514 ; n16514_not
g35685 not n27512 ; n27512_not
g35686 not n14732 ; n14732_not
g35687 not n10826 ; n10826_not
g35688 not n23237 ; n23237_not
g35689 not n22436 ; n22436_not
g35690 not n28034 ; n28034_not
g35691 not n16325 ; n16325_not
g35692 not n12176 ; n12176_not
g35693 not n28016 ; n28016_not
g35694 not n22544 ; n22544_not
g35695 not n23066 ; n23066_not
g35696 not n22571 ; n22571_not
g35697 not n14255 ; n14255_not
g35698 not n16622 ; n16622_not
g35699 not n22607 ; n22607_not
g35700 not n23156 ; n23156_not
g35701 not n16604 ; n16604_not
g35702 not n22643 ; n22643_not
g35703 not n23147 ; n23147_not
g35704 not n22652 ; n22652_not
g35705 not n22616 ; n22616_not
g35706 not n11519 ; n11519_not
g35707 not n12167 ; n12167_not
g35708 not n17441 ; n17441_not
g35709 not n21284 ; n21284_not
g35710 not n23840 ; n23840_not
g35711 not n10448 ; n10448_not
g35712 not n14354 ; n14354_not
g35713 not n26531 ; n26531_not
g35714 not n21356 ; n21356_not
g35715 not n21365 ; n21365_not
g35716 not n16082 ; n16082_not
g35717 not n17333 ; n17333_not
g35718 not n26630 ; n26630_not
g35719 not n17162 ; n17162_not
g35720 not n17261 ; n17261_not
g35721 not n23750 ; n23750_not
g35722 not n26333 ; n26333_not
g35723 not n11609 ; n11609_not
g35724 not n12077 ; n12077_not
g35725 not n12590 ; n12590_not
g35726 not n17702 ; n17702_not
g35727 not n26360 ; n26360_not
g35728 not n20726 ; n20726_not
g35729 not n25802 ; n25802_not
g35730 not n11573 ; n11573_not
g35731 not n29411 ; n29411_not
g35732 not n15074 ; n15074_not
g35733 not n11096 ; n11096_not
g35734 not n26405 ; n26405_not
g35735 not n29132 ; n29132_not
g35736 not n26432 ; n26432_not
g35737 not n23912 ; n23912_not
g35738 not n11069 ; n11069_not
g35739 not n29240 ; n29240_not
g35740 not n26504 ; n26504_not
g35741 not n10286 ; n10286_not
g35742 not n23624 ; n23624_not
g35743 not n23534 ; n23534_not
g35744 not n10628 ; n10628_not
g35745 not n10277 ; n10277_not
g35746 not n14921 ; n14921_not
g35747 not n17081 ; n17081_not
g35748 not n23552 ; n23552_not
g35749 not n17063 ; n17063_not
g35750 not n21824 ; n21824_not
g35751 not n21653 ; n21653_not
g35752 not n10709 ; n10709_not
g35753 not n16181 ; n16181_not
g35754 not n23516 ; n23516_not
g35755 not n14903 ; n14903_not
g35756 not n21455 ; n21455_not
g35757 not n28421 ; n28421_not
g35758 not n21923 ; n21923_not
g35759 not n17018 ; n17018_not
g35760 not n29060 ; n29060_not
g35761 not n17234 ; n17234_not
g35762 not n21536 ; n21536_not
g35763 not n12365 ; n12365_not
g35764 not n23705 ; n23705_not
g35765 not n12491 ; n12491_not
g35766 not n29015 ; n29015_not
g35767 not n29006 ; n29006_not
g35768 not n12473 ; n12473_not
g35769 not n17144 ; n17144_not
g35770 not n21644 ; n21644_not
g35771 not n12383 ; n12383_not
g35772 not n21419 ; n21419_not
g35773 not n23651 ; n23651_not
g35774 not n25262 ; n25262_not
g35775 not n15614 ; n15614_not
g35776 not n13238 ; n13238_not
g35777 not n25235 ; n25235_not
g35778 not n24902 ; n24902_not
g35779 not n15434 ; n15434_not
g35780 not n31148 ; n31148_not
g35781 not n31760 ; n31760_not
g35782 not n19331 ; n19331_not
g35783 not n31175 ; n31175_not
g35784 not n15632 ; n15632_not
g35785 not n19025 ; n19025_not
g35786 not n31661 ; n31661_not
g35787 not n31751 ; n31751_not
g35788 not n25334 ; n25334_not
g35789 not n31319 ; n31319_not
g35790 not n11339 ; n11339_not
g35791 not n31463 ; n31463_not
g35792 not n19304 ; n19304_not
g35793 not n25316 ; n25316_not
g35794 not n31922 ; n31922_not
g35795 not n31472 ; n31472_not
g35796 not n24740 ; n24740_not
g35797 not n31085 ; n31085_not
g35798 not n10466 ; n10466_not
g35799 not n11267 ; n11267_not
g35800 not n31094 ; n31094_not
g35801 not n31904 ; n31904_not
g35802 not n25505 ; n25505_not
g35803 not n15524 ; n15524_not
g35804 not n24605 ; n24605_not
g35805 not n25901 ; n25901_not
g35806 not n31247 ; n31247_not
g35807 not n18341 ; n18341_not
g35808 not n25532 ; n25532_not
g35809 not n31616 ; n31616_not
g35810 not n10565 ; n10565_not
g35811 not n25181 ; n25181_not
g35812 not n31625 ; n31625_not
g35813 not n31256 ; n31256_not
g35814 not n25127 ; n25127_not
g35815 not n15542 ; n15542_not
g35816 not n15650 ; n15650_not
g35817 not n10574 ; n10574_not
g35818 not n10439 ; n10439_not
g35819 not n19250 ; n19250_not
g35820 not n15353 ; n15353_not
g35821 not n31274 ; n31274_not
g35822 not n13526 ; n13526_not
g35823 not n24812 ; n24812_not
g35824 not n15560 ; n15560_not
g35825 not n25550 ; n25550_not
g35826 not n13535 ; n13535_not
g35827 not n18710 ; n18710_not
g35828 not n19007 ; n19007_not
g35829 not n19340 ; n19340_not
g35830 not n25208 ; n25208_not
g35831 not n18422 ; n18422_not
g35832 not n31238 ; n31238_not
g35833 not n31715 ; n31715_not
g35834 not n31283 ; n31283_not
g35835 not n13661 ; n13661_not
g35836 not n18431 ; n18431_not
g35837 not n24722 ; n24722_not
g35838 not n25415 ; n25415_not
g35839 not n10547 ; n10547_not
g35840 not n18323 ; n18323_not
g35841 not n30923 ; n30923_not
g35842 not n30941 ; n30941_not
g35843 not n25370 ; n25370_not
g35844 not n25451 ; n25451_not
g35845 not n19232 ; n19232_not
g35846 not n19151 ; n19151_not
g35847 not n32093 ; n32093_not
g35848 not n31355 ; n31355_not
g35849 not n25721 ; n25721_not
g35850 not n26027 ; n26027_not
g35851 not n31436 ; n31436_not
g35852 not n18611 ; n18611_not
g35853 not n13418 ; n13418_not
g35854 not n11915 ; n11915_not
g35855 not n32039 ; n32039_not
g35856 not n18503 ; n18503_not
g35857 not n19205 ; n19205_not
g35858 not n19115 ; n19115_not
g35859 not n24920 ; n24920_not
g35860 not n19106 ; n19106_not
g35861 not n12842 ; n12842_not
g35862 not n18521 ; n18521_not
g35863 not n10484 ; n10484_not
g35864 not n20790 ; n20790_not
g35865 not n21546 ; n21546_not
g35866 not n10467 ; n10467_not
g35867 not n11637 ; n11637_not
g35868 not n31581 ; n31581_not
g35869 not n29610 ; n29610_not
g35870 not n17235 ; n17235_not
g35871 not n19170 ; n19170_not
g35872 not n23733 ; n23733_not
g35873 not n20916 ; n20916_not
g35874 not n14274 ; n14274_not
g35875 not n14931 ; n14931_not
g35876 not n23634 ; n23634_not
g35877 not n11457 ; n11457_not
g35878 not n16083 ; n16083_not
g35879 not n26604 ; n26604_not
g35880 not n24147 ; n24147_not
g35881 not n20934 ; n20934_not
g35882 not n15408 ; n15408_not
g35883 not n15543 ; n15543_not
g35884 not n20817 ; n20817_not
g35885 not n21627 ; n21627_not
g35886 not n20826 ; n20826_not
g35887 not n10296 ; n10296_not
g35888 not n11439 ; n11439_not
g35889 not n18432 ; n18432_not
g35890 not n29007 ; n29007_not
g35891 not n31617 ; n31617_not
g35892 not n26316 ; n26316_not
g35893 not n25137 ; n25137_not
g35894 not n20844 ; n20844_not
g35895 not n23661 ; n23661_not
g35896 not n29025 ; n29025_not
g35897 not n22482 ; n22482_not
g35898 not n29034 ; n29034_not
g35899 not n20862 ; n20862_not
g35900 not n21564 ; n21564_not
g35901 not n22473 ; n22473_not
g35902 not n23715 ; n23715_not
g35903 not n17208 ; n17208_not
g35904 not n11376 ; n11376_not
g35905 not n20880 ; n20880_not
g35906 not n10737 ; n10737_not
g35907 not n26820 ; n26820_not
g35908 not n14454 ; n14454_not
g35909 not n29214 ; n29214_not
g35910 not n29412 ; n29412_not
g35911 not n15255 ; n15255_not
g35912 not n15444 ; n15444_not
g35913 not n24633 ; n24633_not
g35914 not n26514 ; n26514_not
g35915 not n11097 ; n11097_not
g35916 not n15417 ; n15417_not
g35917 not n31491 ; n31491_not
g35918 not n23850 ; n23850_not
g35919 not n17370 ; n17370_not
g35920 not n25605 ; n25605_not
g35921 not n12159 ; n12159_not
g35922 not n25821 ; n25821_not
g35923 not n26451 ; n26451_not
g35924 not n22671 ; n22671_not
g35925 not n31473 ; n31473_not
g35926 not n21186 ; n21186_not
g35927 not n11673 ; n11673_not
g35928 not n12096 ; n12096_not
g35929 not n29115 ; n29115_not
g35930 not n26415 ; n26415_not
g35931 not n19116 ; n19116_not
g35932 not n23931 ; n23931_not
g35933 not n21159 ; n21159_not
g35934 not n10719 ; n10719_not
g35935 not n23922 ; n23922_not
g35936 not n20952 ; n20952_not
g35937 not n23751 ; n23751_not
g35938 not n20970 ; n20970_not
g35939 not n17064 ; n17064_not
g35940 not n14292 ; n14292_not
g35941 not n15561 ; n15561_not
g35942 not n25560 ; n25560_not
g35943 not n17703 ; n17703_not
g35944 not n18414 ; n18414_not
g35945 not n17334 ; n17334_not
g35946 not n10494 ; n10494_not
g35947 not n29502 ; n29502_not
g35948 not n26073 ; n26073_not
g35949 not n26352 ; n26352_not
g35950 not n13158 ; n13158_not
g35951 not n21375 ; n21375_not
g35952 not n17343 ; n17343_not
g35953 not n12339 ; n12339_not
g35954 not n19035 ; n19035_not
g35955 not n11583 ; n11583_not
g35956 not n29430 ; n29430_not
g35957 not n23814 ; n23814_not
g35958 not n26550 ; n26550_not
g35959 not n25641 ; n25641_not
g35960 not n19053 ; n19053_not
g35961 not n18342 ; n18342_not
g35962 not n20664 ; n20664_not
g35963 not n21069 ; n21069_not
g35964 not n29205 ; n29205_not
g35965 not n17406 ; n17406_not
g35966 not n28035 ; n28035_not
g35967 not n25335 ; n25335_not
g35968 not n16182 ; n16182_not
g35969 not n16308 ; n16308_not
g35970 not n14625 ; n14625_not
g35971 not n25470 ; n25470_not
g35972 not n16650 ; n16650_not
g35973 not n16335 ; n16335_not
g35974 not n27207 ; n27207_not
g35975 not n22536 ; n22536_not
g35976 not n10557 ; n10557_not
g35977 not n22545 ; n22545_not
g35978 not n23184 ; n23184_not
g35979 not n22563 ; n22563_not
g35980 not n27711 ; n27711_not
g35981 not n22572 ; n22572_not
g35982 not n23166 ; n23166_not
g35983 not n16623 ; n16623_not
g35984 not n12258 ; n12258_not
g35985 not n31905 ; n31905_not
g35986 not n31851 ; n31851_not
g35987 not n16272 ; n16272_not
g35988 not n16290 ; n16290_not
g35989 not n12249 ; n12249_not
g35990 not n25308 ; n25308_not
g35991 not n18711 ; n18711_not
g35992 not n22176 ; n22176_not
g35993 not n20835 ; n20835_not
g35994 not n21519 ; n21519_not
g35995 not n16740 ; n16740_not
g35996 not n31914 ; n31914_not
g35997 not n31923 ; n31923_not
g35998 not n12195 ; n12195_not
g35999 not n25317 ; n25317_not
g36000 not n23238 ; n23238_not
g36001 not n12645 ; n12645_not
g36002 not n11493 ; n11493_not
g36003 not n10890 ; n10890_not
g36004 not n13392 ; n13392_not
g36005 not n23094 ; n23094_not
g36006 not n16551 ; n16551_not
g36007 not n25074 ; n25074_not
g36008 not n22734 ; n22734_not
g36009 not n23076 ; n23076_not
g36010 not n16533 ; n16533_not
g36011 not n22806 ; n22806_not
g36012 not n18540 ; n18540_not
g36013 not n14715 ; n14715_not
g36014 not n18522 ; n18522_not
g36015 not n25416 ; n25416_not
g36016 not n27513 ; n27513_not
g36017 not n18504 ; n18504_not
g36018 not n22446 ; n22446_not
g36019 not n13374 ; n13374_not
g36020 not n22932 ; n22932_not
g36021 not n14643 ; n14643_not
g36022 not n22617 ; n22617_not
g36023 not n18621 ; n18621_not
g36024 not n15480 ; n15480_not
g36025 not n16434 ; n16434_not
g36026 not n14652 ; n14652_not
g36027 not n13059 ; n13059_not
g36028 not n22419 ; n22419_not
g36029 not n23148 ; n23148_not
g36030 not n16380 ; n16380_not
g36031 not n27225 ; n27225_not
g36032 not n23139 ; n23139_not
g36033 not n14670 ; n14670_not
g36034 not n13428 ; n13428_not
g36035 not n27243 ; n27243_not
g36036 not n25380 ; n25380_not
g36037 not n21843 ; n21843_not
g36038 not n23535 ; n23535_not
g36039 not n23526 ; n23526_not
g36040 not n21861 ; n21861_not
g36041 not n14913 ; n14913_not
g36042 not n10944 ; n10944_not
g36043 not n17046 ; n17046_not
g36044 not n21906 ; n21906_not
g36045 not n25191 ; n25191_not
g36046 not n21456 ; n21456_not
g36047 not n31716 ; n31716_not
g36048 not n17019 ; n17019_not
g36049 not n21942 ; n21942_not
g36050 not n28422 ; n28422_not
g36051 not n28260 ; n28260_not
g36052 not n17109 ; n17109_not
g36053 not n21708 ; n21708_not
g36054 not n12384 ; n12384_not
g36055 not n10575 ; n10575_not
g36056 not n21744 ; n21744_not
g36057 not n17091 ; n17091_not
g36058 not n31680 ; n31680_not
g36059 not n21762 ; n21762_not
g36060 not n23580 ; n23580_not
g36061 not n23571 ; n23571_not
g36062 not n15462 ; n15462_not
g36063 not n26640 ; n26640_not
g36064 not n10746 ; n10746_not
g36065 not n10683 ; n10683_not
g36066 not n21807 ; n21807_not
g36067 not n28602 ; n28602_not
g36068 not n18900 ; n18900_not
g36069 not n16902 ; n16902_not
g36070 not n21591 ; n21591_not
g36071 not n23373 ; n23373_not
g36072 not n22158 ; n22158_not
g36073 not n15525 ; n15525_not
g36074 not n23346 ; n23346_not
g36075 not n25245 ; n25245_not
g36076 not n31842 ; n31842_not
g36077 not n22509 ; n22509_not
g36078 not n16263 ; n16263_not
g36079 not n16830 ; n16830_not
g36080 not n10917 ; n10917_not
g36081 not n25272 ; n25272_not
g36082 not n16812 ; n16812_not
g36083 not n23292 ; n23292_not
g36084 not n22293 ; n22293_not
g36085 not n22239 ; n22239_not
g36086 not n11781 ; n11781_not
g36087 not n18450 ; n18450_not
g36088 not n21960 ; n21960_not
g36089 not n23490 ; n23490_not
g36090 not n28404 ; n28404_not
g36091 not n10818 ; n10818_not
g36092 not n23472 ; n23472_not
g36093 not n14427 ; n14427_not
g36094 not n10764 ; n10764_not
g36095 not n23454 ; n23454_not
g36096 not n31752 ; n31752_not
g36097 not n27135 ; n27135_not
g36098 not n22059 ; n22059_not
g36099 not n31761 ; n31761_not
g36100 not n16245 ; n16245_not
g36101 not n12357 ; n12357_not
g36102 not n25218 ; n25218_not
g36103 not n21645 ; n21645_not
g36104 not n24507 ; n24507_not
g36105 not n11853 ; n11853_not
g36106 not n12690 ; n12690_not
g36107 not n17910 ; n17910_not
g36108 not n26217 ; n26217_not
g36109 not n24309 ; n24309_not
g36110 not n30537 ; n30537_not
g36111 not n19332 ; n19332_not
g36112 not n12663 ; n12663_not
g36113 not n30519 ; n30519_not
g36114 not n18270 ; n18270_not
g36115 not n24741 ; n24741_not
g36116 not n11808 ; n11808_not
g36117 not n20448 ; n20448_not
g36118 not n31095 ; n31095_not
g36119 not n13860 ; n13860_not
g36120 not n18144 ; n18144_not
g36121 not n15147 ; n15147_not
g36122 not n30483 ; n30483_not
g36123 not n12681 ; n12681_not
g36124 not n11961 ; n11961_not
g36125 not n30717 ; n30717_not
g36126 not n11952 ; n11952_not
g36127 not n24705 ; n24705_not
g36128 not n11268 ; n11268_not
g36129 not n31338 ; n31338_not
g36130 not n30078 ; n30078_not
g36131 not n20565 ; n20565_not
g36132 not n24525 ; n24525_not
g36133 not n30672 ; n30672_not
g36134 not n30645 ; n30645_not
g36135 not n14166 ; n14166_not
g36136 not n20547 ; n20547_not
g36137 not n12861 ; n12861_not
g36138 not n14148 ; n14148_not
g36139 not n14139 ; n14139_not
g36140 not n24912 ; n24912_not
g36141 not n20529 ; n20529_not
g36142 not n24723 ; n24723_not
g36143 not n26109 ; n26109_not
g36144 not n19323 ; n19323_not
g36145 not n25920 ; n25920_not
g36146 not n30159 ; n30159_not
g36147 not n24516 ; n24516_not
g36148 not n13095 ; n13095_not
g36149 not n20088 ; n20088_not
g36150 not n19224 ; n19224_not
g36151 not n24408 ; n24408_not
g36152 not n18063 ; n18063_not
g36153 not n13941 ; n13941_not
g36154 not n26145 ; n26145_not
g36155 not n20178 ; n20178_not
g36156 not n31257 ; n31257_not
g36157 not n24822 ; n24822_not
g36158 not n20196 ; n20196_not
g36159 not n20259 ; n20259_not
g36160 not n31239 ; n31239_not
g36161 not n30366 ; n30366_not
g36162 not n11187 ; n11187_not
g36163 not n18081 ; n18081_not
g36164 not n13923 ; n13923_not
g36165 not n18126 ; n18126_not
g36166 not n24426 ; n24426_not
g36167 not n18090 ; n18090_not
g36168 not n13644 ; n13644_not
g36169 not n13932 ; n13932_not
g36170 not n26154 ; n26154_not
g36171 not n19008 ; n19008_not
g36172 not n18243 ; n18243_not
g36173 not n11628 ; n11628_not
g36174 not n26181 ; n26181_not
g36175 not n11817 ; n11817_not
g36176 not n10395 ; n10395_not
g36177 not n20376 ; n20376_not
g36178 not n19350 ; n19350_not
g36179 not n15165 ; n15165_not
g36180 not n19512 ; n19512_not
g36181 not n13806 ; n13806_not
g36182 not n11925 ; n11925_not
g36183 not n20367 ; n20367_not
g36184 not n25524 ; n25524_not
g36185 not n24390 ; n24390_not
g36186 not n18216 ; n18216_not
g36187 not n30258 ; n30258_not
g36188 not n11169 ; n11169_not
g36189 not n24471 ; n24471_not
g36190 not n23913 ; n23913_not
g36191 not n24462 ; n24462_not
g36192 not n31275 ; n31275_not
g36193 not n30762 ; n30762_not
g36194 not n17820 ; n17820_not
g36195 not n30627 ; n30627_not
g36196 not n26082 ; n26082_not
g36197 not n19260 ; n19260_not
g36198 not n24228 ; n24228_not
g36199 not n15372 ; n15372_not
g36200 not n14184 ; n14184_not
g36201 not n30816 ; n30816_not
g36202 not n20646 ; n20646_not
g36203 not n14256 ; n14256_not
g36204 not n20655 ; n20655_not
g36205 not n26253 ; n26253_not
g36206 not n12843 ; n12843_not
g36207 not n31374 ; n31374_not
g36208 not n20277 ; n20277_not
g36209 not n10629 ; n10629_not
g36210 not n30753 ; n30753_not
g36211 not n19710 ; n19710_not
g36212 not n25731 ; n25731_not
g36213 not n24237 ; n24237_not
g36214 not n11763 ; n11763_not
g36215 not n18217 ; n18217_not
g36216 not n18541 ; n18541_not
g36217 not n13654 ; n13654_not
g36218 not n10639 ; n10639_not
g36219 not n12367 ; n12367_not
g36220 not n27136 ; n27136_not
g36221 not n16246 ; n16246_not
g36222 not n10846 ; n10846_not
g36223 not n13951 ; n13951_not
g36224 not n25921 ; n25921_not
g36225 not n30844 ; n30844_not
g36226 not n27307 ; n27307_not
g36227 not n31780 ; n31780_not
g36228 not n14464 ; n14464_not
g36229 not n30853 ; n30853_not
g36230 not n22843 ; n22843_not
g36231 not n12772 ; n12772_not
g36232 not n13339 ; n13339_not
g36233 not n16228 ; n16228_not
g36234 not n14455 ; n14455_not
g36235 not n13438 ; n13438_not
g36236 not n13627 ; n13627_not
g36237 not n13285 ; n13285_not
g36238 not n18802 ; n18802_not
g36239 not n22852 ; n22852_not
g36240 not n18523 ; n18523_not
g36241 not n10765 ; n10765_not
g36242 not n28315 ; n28315_not
g36243 not n30835 ; n30835_not
g36244 not n23347 ; n23347_not
g36245 not n18622 ; n18622_not
g36246 not n12880 ; n12880_not
g36247 not n28216 ; n28216_not
g36248 not n28225 ; n28225_not
g36249 not n22168 ; n22168_not
g36250 not n32086 ; n32086_not
g36251 not n11629 ; n11629_not
g36252 not n30448 ; n30448_not
g36253 not n12349 ; n12349_not
g36254 not n10819 ; n10819_not
g36255 not n27154 ; n27154_not
g36256 not n28243 ; n28243_not
g36257 not n24580 ; n24580_not
g36258 not n24481 ; n24481_not
g36259 not n22627 ; n22627_not
g36260 not n25219 ; n25219_not
g36261 not n22609 ; n22609_not
g36262 not n22780 ; n22780_not
g36263 not n21619 ; n21619_not
g36264 not n27622 ; n27622_not
g36265 not n13375 ; n13375_not
g36266 not n16912 ; n16912_not
g36267 not n24616 ; n24616_not
g36268 not n11791 ; n11791_not
g36269 not n21934 ; n21934_not
g36270 not n10099 ; n10099_not
g36271 not n28432 ; n28432_not
g36272 not n19720 ; n19720_not
g36273 not n18145 ; n18145_not
g36274 not n25192 ; n25192_not
g36275 not n14725 ; n14725_not
g36276 not n30754 ; n30754_not
g36277 not n25417 ; n25417_not
g36278 not n16507 ; n16507_not
g36279 not n12457 ; n12457_not
g36280 not n11845 ; n11845_not
g36281 not n12763 ; n12763_not
g36282 not n22825 ; n22825_not
g36283 not n22960 ; n22960_not
g36284 not n11377 ; n11377_not
g36285 not n22582 ; n22582_not
g36286 not n12466 ; n12466_not
g36287 not n22915 ; n22915_not
g36288 not n22942 ; n22942_not
g36289 not n25525 ; n25525_not
g36290 not n16183 ; n16183_not
g36291 not n28522 ; n28522_not
g36292 not n28531 ; n28531_not
g36293 not n15463 ; n15463_not
g36294 not n27460 ; n27460_not
g36295 not n32059 ; n32059_not
g36296 not n30394 ; n30394_not
g36297 not n21475 ; n21475_not
g36298 not n18190 ; n18190_not
g36299 not n31636 ; n31636_not
g36300 not n28360 ; n28360_not
g36301 not n23914 ; n23914_not
g36302 not n27334 ; n27334_not
g36303 not n27361 ; n27361_not
g36304 not n13915 ; n13915_not
g36305 not n18820 ; n18820_not
g36306 not n22870 ; n22870_not
g36307 not n23149 ; n23149_not
g36308 not n23482 ; n23482_not
g36309 not n28261 ; n28261_not
g36310 not n18172 ; n18172_not
g36311 not n18505 ; n18505_not
g36312 not n30376 ; n30376_not
g36313 not n28414 ; n28414_not
g36314 not n18604 ; n18604_not
g36315 not n27514 ; n27514_not
g36316 not n30367 ; n30367_not
g36317 not n23491 ; n23491_not
g36318 not n15760 ; n15760_not
g36319 not n24625 ; n24625_not
g36320 not n22492 ; n22492_not
g36321 not n22339 ; n22339_not
g36322 not n15724 ; n15724_not
g36323 not n22348 ; n22348_not
g36324 not n14437 ; n14437_not
g36325 not n22357 ; n22357_not
g36326 not n22456 ; n22456_not
g36327 not n22366 ; n22366_not
g36328 not n13492 ; n13492_not
g36329 not n22690 ; n22690_not
g36330 not n24724 ; n24724_not
g36331 not n30439 ; n30439_not
g36332 not n25318 ; n25318_not
g36333 not n22429 ; n22429_not
g36334 not n24517 ; n24517_not
g36335 not n23239 ; n23239_not
g36336 not n16408 ; n16408_not
g36337 not n27901 ; n27901_not
g36338 not n16723 ; n16723_not
g36339 not n12691 ; n12691_not
g36340 not n18451 ; n18451_not
g36341 not n27721 ; n27721_not
g36342 not n16741 ; n16741_not
g36343 not n14815 ; n14815_not
g36344 not n16552 ; n16552_not
g36345 not n27208 ; n27208_not
g36346 not n15364 ; n15364_not
g36347 not n25363 ; n25363_not
g36348 not n22438 ; n22438_not
g36349 not n11872 ; n11872_not
g36350 not n14635 ; n14635_not
g36351 not n18640 ; n18640_not
g36352 not n22465 ; n22465_not
g36353 not n28009 ; n28009_not
g36354 not n19801 ; n19801_not
g36355 not n16345 ; n16345_not
g36356 not n24715 ; n24715_not
g36357 not n16363 ; n16363_not
g36358 not n16336 ; n16336_not
g36359 not n15256 ; n15256_not
g36360 not n11908 ; n11908_not
g36361 not n12862 ; n12862_not
g36362 not n12871 ; n12871_not
g36363 not n16534 ; n16534_not
g36364 not n10558 ; n10558_not
g36365 not n19900 ; n19900_not
g36366 not n25336 ; n25336_not
g36367 not n31852 ; n31852_not
g36368 not n30493 ; n30493_not
g36369 not n25444 ; n25444_not
g36370 not n16813 ; n16813_not
g36371 not n30745 ; n30745_not
g36372 not n30475 ; n30475_not
g36373 not n26902 ; n26902_not
g36374 not n22249 ; n22249_not
g36375 not n31096 ; n31096_not
g36376 not n28153 ; n28153_not
g36377 not n16264 ; n16264_not
g36378 not n24229 ; n24229_not
g36379 not n23086 ; n23086_not
g36380 not n16831 ; n16831_not
g36381 not n14653 ; n14653_not
g36382 not n28180 ; n28180_not
g36383 not n16426 ; n16426_not
g36384 not n31843 ; n31843_not
g36385 not n25246 ; n25246_not
g36386 not n10864 ; n10864_not
g36387 not n31825 ; n31825_not
g36388 not n15652 ; n15652_not
g36389 not n23338 ; n23338_not
g36390 not n16606 ; n16606_not
g36391 not n30556 ; n30556_not
g36392 not n30682 ; n30682_not
g36393 not n16291 ; n16291_not
g36394 not n27244 ; n27244_not
g36395 not n25381 ; n25381_not
g36396 not n31834 ; n31834_not
g36397 not n30538 ; n30538_not
g36398 not n22834 ; n22834_not
g36399 not n22663 ; n22663_not
g36400 not n12637 ; n12637_not
g36401 not n11944 ; n11944_not
g36402 not n27190 ; n27190_not
g36403 not n30817 ; n30817_not
g36404 not n30691 ; n30691_not
g36405 not n12277 ; n12277_not
g36406 not n10891 ; n10891_not
g36407 not n11755 ; n11755_not
g36408 not n16381 ; n16381_not
g36409 not n18721 ; n18721_not
g36410 not n12295 ; n12295_not
g36411 not n25480 ; n25480_not
g36412 not n22519 ; n22519_not
g36413 not n28126 ; n28126_not
g36414 not n29233 ; n29233_not
g36415 not n23860 ; n23860_not
g36416 not n21259 ; n21259_not
g36417 not n24913 ; n24913_not
g36418 not n19081 ; n19081_not
g36419 not n31492 ; n31492_not
g36420 not n29224 ; n29224_not
g36421 not n17434 ; n17434_not
g36422 not n21295 ; n21295_not
g36423 not n29206 ; n29206_not
g36424 not n25570 ; n25570_not
g36425 not n19063 ; n19063_not
g36426 not n24247 ; n24247_not
g36427 not n11674 ; n11674_not
g36428 not n24265 ; n24265_not
g36429 not n20566 ; n20566_not
g36430 not n29116 ; n29116_not
g36431 not n29305 ; n29305_not
g36432 not n11539 ; n11539_not
g36433 not n26443 ; n26443_not
g36434 not n20557 ; n20557_not
g36435 not n29251 ; n29251_not
g36436 not n29260 ; n29260_not
g36437 not n25606 ; n25606_not
g36438 not n14167 ; n14167_not
g36439 not n25822 ; n25822_not
g36440 not n31474 ; n31474_not
g36441 not n19333 ; n19333_not
g36442 not n29107 ; n29107_not
g36443 not n18415 ; n18415_not
g36444 not n26641 ; n26641_not
g36445 not n17038 ; n17038_not
g36446 not n12574 ; n12574_not
g36447 not n17092 ; n17092_not
g36448 not n31564 ; n31564_not
g36449 not n23752 ; n23752_not
g36450 not n19018 ; n19018_not
g36451 not n12673 ; n12673_not
g36452 not n13870 ; n13870_not
g36453 not n18325 ; n18325_not
g36454 not n31537 ; n31537_not
g36455 not n21439 ; n21439_not
g36456 not n17254 ; n17254_not
g36457 not n24292 ; n24292_not
g36458 not n26542 ; n26542_not
g36459 not n23824 ; n23824_not
g36460 not n29161 ; n29161_not
g36461 not n10729 ; n10729_not
g36462 not n14095 ; n14095_not
g36463 not n13186 ; n13186_not
g36464 not n14914 ; n14914_not
g36465 not n17353 ; n17353_not
g36466 not n15445 ; n15445_not
g36467 not n15175 ; n15175_not
g36468 not n17911 ; n17911_not
g36469 not n30178 ; n30178_not
g36470 not n21385 ; n21385_not
g36471 not n19225 ; n19225_not
g36472 not n20827 ; n20827_not
g36473 not n20368 ; n20368_not
g36474 not n20845 ; n20845_not
g36475 not n11728 ; n11728_not
g36476 not n20863 ; n20863_not
g36477 not n14608 ; n14608_not
g36478 not n31375 ; n31375_not
g36479 not n20449 ; n20449_not
g36480 not n20881 ; n20881_not
g36481 not n31294 ; n31294_not
g36482 not n19180 ; n19180_not
g36483 not n17236 ; n17236_not
g36484 not n13177 ; n13177_not
g36485 not n20917 ; n20917_not
g36486 not n25660 ; n25660_not
g36487 not n17731 ; n17731_not
g36488 not n20179 ; n20179_not
g36489 not n18370 ; n18370_not
g36490 not n24148 ; n24148_not
g36491 not n14266 ; n14266_not
g36492 not n20791 ; n20791_not
g36493 not n29800 ; n29800_not
g36494 not n20809 ; n20809_not
g36495 not n15940 ; n15940_not
g36496 not n11692 ; n11692_not
g36497 not n10684 ; n10684_not
g36498 not n17740 ; n17740_not
g36499 not n31393 ; n31393_not
g36500 not n11584 ; n11584_not
g36501 not n19144 ; n19144_not
g36502 not n31348 ; n31348_not
g36503 not n29413 ; n29413_not
g36504 not n19270 ; n19270_not
g36505 not n11098 ; n11098_not
g36506 not n11296 ; n11296_not
g36507 not n12565 ; n12565_not
g36508 not n11557 ; n11557_not
g36509 not n12556 ; n12556_not
g36510 not n19117 ; n19117_not
g36511 not n12619 ; n12619_not
g36512 not n12628 ; n12628_not
g36513 not n14338 ; n14338_not
g36514 not n20935 ; n20935_not
g36515 not n25705 ; n25705_not
g36516 not n20656 ; n20656_not
g36517 not n20953 ; n20953_not
g36518 not n24058 ; n24058_not
g36519 not n20971 ; n20971_not
g36520 not n14284 ; n14284_not
g36521 not n31447 ; n31447_not
g36522 not n26344 ; n26344_not
g36523 not n17704 ; n17704_not
g36524 not n10477 ; n10477_not
g36525 not n29512 ; n29512_not
g36526 not n26245 ; n26245_not
g36527 not n11269 ; n11269_not
g36528 not n25732 ; n25732_not
g36529 not n29431 ; n29431_not
g36530 not n19315 ; n19315_not
g36531 not n26830 ; n26830_not
g36532 not n10576 ; n10576_not
g36533 not n16156 ; n16156_not
g36534 not n21682 ; n21682_not
g36535 not n30277 ; n30277_not
g36536 not n23644 ; n23644_not
g36537 not n31645 ; n31645_not
g36538 not n18028 ; n18028_not
g36539 not n21664 ; n21664_not
g36540 not n25138 ; n25138_not
g36541 not n25840 ; n25840_not
g36542 not n13546 ; n13546_not
g36543 not n17119 ; n17119_not
g36544 not n18433 ; n18433_not
g36545 not n31276 ; n31276_not
g36546 not n26803 ; n26803_not
g36547 not n17137 ; n17137_not
g36548 not n13960 ; n13960_not
g36549 not n31609 ; n31609_not
g36550 not n23626 ; n23626_not
g36551 not n17173 ; n17173_not
g36552 not n14950 ; n14950_not
g36553 not n31618 ; n31618_not
g36554 not n21592 ; n21592_not
g36555 not n14932 ; n14932_not
g36556 not n31690 ; n31690_not
g36557 not n19036 ; n19036_not
g36558 not n18091 ; n18091_not
g36559 not n11188 ; n11188_not
g36560 not n10747 ; n10747_not
g36561 not n31672 ; n31672_not
g36562 not n21835 ; n21835_not
g36563 not n23545 ; n23545_not
g36564 not n18901 ; n18901_not
g36565 not n24427 ; n24427_not
g36566 not n16165 ; n16165_not
g36567 not n17074 ; n17074_not
g36568 not n28612 ; n28612_not
g36569 not n28621 ; n28621_not
g36570 not n12538 ; n12538_not
g36571 not n11836 ; n11836_not
g36572 not n18073 ; n18073_not
g36573 not n24418 ; n24418_not
g36574 not n20287 ; n20287_not
g36575 not n23581 ; n23581_not
g36576 not n21655 ; n21655_not
g36577 not n21736 ; n21736_not
g36578 not n31258 ; n31258_not
g36579 not n21727 ; n21727_not
g36580 not n11458 ; n11458_not
g36581 not n17191 ; n17191_not
g36582 not n31267 ; n31267_not
g36583 not n15193 ; n15193_not
g36584 not n20386 ; n20386_not
g36585 not n29044 ; n29044_not
g36586 not n15544 ; n15544_not
g36587 not n29053 ; n29053_not
g36588 not n31582 ; n31582_not
g36589 not n21529 ; n21529_not
g36590 not n18352 ; n18352_not
g36591 not n17245 ; n17245_not
g36592 not n23743 ; n23743_not
g36593 not n21178 ; n21178_not
g36594 not n29026 ; n29026_not
g36595 not n21574 ; n21574_not
g36596 not n10495 ; n10495_not
g36597 not n31591 ; n31591_not
g36598 not n23069 ; n23069_not
g36599 not n23249 ; n23249_not
g36600 not n10559 ; n10559_not
g36601 not n27155 ; n27155_not
g36602 not n16427 ; n16427_not
g36603 not n26327 ; n26327_not
g36604 not n15356 ; n15356_not
g36605 not n27290 ; n27290_not
g36606 not n15905 ; n15905_not
g36607 not n24338 ; n24338_not
g36608 not n11648 ; n11648_not
g36609 not n14780 ; n14780_not
g36610 not n25904 ; n25904_not
g36611 not n23762 ; n23762_not
g36612 not n24752 ; n24752_not
g36613 not n24167 ; n24167_not
g36614 not n24716 ; n24716_not
g36615 not n16418 ; n16418_not
g36616 not n11639 ; n11639_not
g36617 not n23672 ; n23672_not
g36618 not n24635 ; n24635_not
g36619 not n11990 ; n11990_not
g36620 not n10694 ; n10694_not
g36621 not n26138 ; n26138_not
g36622 not n23087 ; n23087_not
g36623 not n24059 ; n24059_not
g36624 not n26606 ; n26606_not
g36625 not n10766 ; n10766_not
g36626 not n23780 ; n23780_not
g36627 not n10793 ; n10793_not
g36628 not n25553 ; n25553_not
g36629 not n23726 ; n23726_not
g36630 not n23582 ; n23582_not
g36631 not n11738 ; n11738_not
g36632 not n26525 ; n26525_not
g36633 not n26660 ; n26660_not
g36634 not n15446 ; n15446_not
g36635 not n24419 ; n24419_not
g36636 not n15626 ; n15626_not
g36637 not n11585 ; n11585_not
g36638 not n16094 ; n16094_not
g36639 not n26930 ; n26930_not
g36640 not n26273 ; n26273_not
g36641 not n14825 ; n14825_not
g36642 not n25940 ; n25940_not
g36643 not n22556 ; n22556_not
g36644 not n22907 ; n22907_not
g36645 not n27443 ; n27443_not
g36646 not n27452 ; n27452_not
g36647 not n25571 ; n25571_not
g36648 not n24905 ; n24905_not
g36649 not n15491 ; n15491_not
g36650 not n27182 ; n27182_not
g36651 not n27407 ; n27407_not
g36652 not n26912 ; n26912_not
g36653 not n16454 ; n16454_not
g36654 not n23186 ; n23186_not
g36655 not n11657 ; n11657_not
g36656 not n25670 ; n25670_not
g36657 not n26624 ; n26624_not
g36658 not n24653 ; n24653_not
g36659 not n23555 ; n23555_not
g36660 not n13736 ; n13736_not
g36661 not n16472 ; n16472_not
g36662 not n24662 ; n24662_not
g36663 not n25733 ; n25733_not
g36664 not n23285 ; n23285_not
g36665 not n24491 ; n24491_not
g36666 not n15257 ; n15257_not
g36667 not n11936 ; n11936_not
g36668 not n26057 ; n26057_not
g36669 not n10748 ; n10748_not
g36670 not n25454 ; n25454_not
g36671 not n23168 ; n23168_not
g36672 not n15662 ; n15662_not
g36673 not n25607 ; n25607_not
g36674 not n23915 ; n23915_not
g36675 not n25742 ; n25742_not
g36676 not n23384 ; n23384_not
g36677 not n25373 ; n25373_not
g36678 not n27218 ; n27218_not
g36679 not n15428 ; n15428_not
g36680 not n23348 ; n23348_not
g36681 not n26804 ; n26804_not
g36682 not n16364 ; n16364_not
g36683 not n26426 ; n26426_not
g36684 not n24365 ; n24365_not
g36685 not n16229 ; n16229_not
g36686 not n15419 ; n15419_not
g36687 not n23681 ; n23681_not
g36688 not n24545 ; n24545_not
g36689 not n15194 ; n15194_not
g36690 not n26228 ; n26228_not
g36691 not n26471 ; n26471_not
g36692 not n16346 ; n16346_not
g36693 not n15761 ; n15761_not
g36694 not n24914 ; n24914_not
g36695 not n26750 ; n26750_not
g36696 not n24284 ; n24284_not
g36697 not n25805 ; n25805_not
g36698 not n11549 ; n11549_not
g36699 not n15464 ; n15464_not
g36700 not n24518 ; n24518_not
g36701 not n23177 ; n23177_not
g36702 not n25922 ; n25922_not
g36703 not n23906 ; n23906_not
g36704 not n25634 ; n25634_not
g36705 not n23690 ; n23690_not
g36706 not n12089 ; n12089_not
g36707 not n23807 ; n23807_not
g36708 not n25751 ; n25751_not
g36709 not n11756 ; n11756_not
g36710 not n10397 ; n10397_not
g36711 not n16049 ; n16049_not
g36712 not n23609 ; n23609_not
g36713 not n26831 ; n26831_not
g36714 not n23483 ; n23483_not
g36715 not n11594 ; n11594_not
g36716 not n23465 ; n23465_not
g36717 not n15554 ; n15554_not
g36718 not n25382 ; n25382_not
g36719 not n15284 ; n15284_not
g36720 not n15176 ; n15176_not
g36721 not n25913 ; n25913_not
g36722 not n26093 ; n26093_not
g36723 not n15608 ; n15608_not
g36724 not n24734 ; n24734_not
g36725 not n16085 ; n16085_not
g36726 not n15473 ; n15473_not
g36727 not n27164 ; n27164_not
g36728 not n11891 ; n11891_not
g36729 not n25139 ; n25139_not
g36730 not n23825 ; n23825_not
g36731 not n23744 ; n23744_not
g36732 not n25535 ; n25535_not
g36733 not n10892 ; n10892_not
g36734 not n23951 ; n23951_not
g36735 not n23429 ; n23429_not
g36736 not n24608 ; n24608_not
g36737 not n26372 ; n26372_not
g36738 not n24347 ; n24347_not
g36739 not n15725 ; n15725_not
g36740 not n30791 ; n30791_not
g36741 not n21386 ; n21386_not
g36742 not n30836 ; n30836_not
g36743 not n17327 ; n17327_not
g36744 not n30854 ; n30854_not
g36745 not n27713 ; n27713_not
g36746 not n29072 ; n29072_not
g36747 not n29063 ; n29063_not
g36748 not n21494 ; n21494_not
g36749 not n29045 ; n29045_not
g36750 not n30944 ; n30944_not
g36751 not n21557 ; n21557_not
g36752 not n22529 ; n22529_not
g36753 not n30953 ; n30953_not
g36754 not n17183 ; n17183_not
g36755 not n12485 ; n12485_not
g36756 not n28208 ; n28208_not
g36757 not n12854 ; n12854_not
g36758 not n17147 ; n17147_not
g36759 not n12872 ; n12872_not
g36760 not n17471 ; n17471_not
g36761 not n30593 ; n30593_not
g36762 not n19910 ; n19910_not
g36763 not n29243 ; n29243_not
g36764 not n30638 ; n30638_not
g36765 not n29225 ; n29225_not
g36766 not n17354 ; n17354_not
g36767 not n17444 ; n17444_not
g36768 not n30683 ; n30683_not
g36769 not n14285 ; n14285_not
g36770 not n14249 ; n14249_not
g36771 not n29171 ; n29171_not
g36772 not n29117 ; n29117_not
g36773 not n29144 ; n29144_not
g36774 not n30746 ; n30746_not
g36775 not n30755 ; n30755_not
g36776 not n21359 ; n21359_not
g36777 not n29108 ; n29108_not
g36778 not n13097 ; n13097_not
g36779 not n21818 ; n21818_not
g36780 not n13484 ; n13484_not
g36781 not n19064 ; n19064_not
g36782 not n28550 ; n28550_not
g36783 not n28532 ; n28532_not
g36784 not n19361 ; n19361_not
g36785 not n28460 ; n28460_not
g36786 not n17039 ; n17039_not
g36787 not n16913 ; n16913_not
g36788 not n21917 ; n21917_not
g36789 not n12458 ; n12458_not
g36790 not n19352 ; n19352_not
g36791 not n13655 ; n13655_not
g36792 not n31286 ; n31286_not
g36793 not n19316 ; n19316_not
g36794 not n18353 ; n18353_not
g36795 not n19307 ; n19307_not
g36796 not n13628 ; n13628_not
g36797 not n28343 ; n28343_not
g36798 not n31079 ; n31079_not
g36799 not n21665 ; n21665_not
g36800 not n13727 ; n13727_not
g36801 not n28802 ; n28802_not
g36802 not n28730 ; n28730_not
g36803 not n19505 ; n19505_not
g36804 not n10964 ; n10964_not
g36805 not n11459 ; n11459_not
g36806 not n28640 ; n28640_not
g36807 not n28631 ; n28631_not
g36808 not n28613 ; n28613_not
g36809 not n17750 ; n17750_not
g36810 not n13916 ; n13916_not
g36811 not n20369 ; n20369_not
g36812 not n13664 ; n13664_not
g36813 not n29810 ; n29810_not
g36814 not n30278 ; n30278_not
g36815 not n18038 ; n18038_not
g36816 not n17732 ; n17732_not
g36817 not n11387 ; n11387_not
g36818 not n20792 ; n20792_not
g36819 not n20297 ; n20297_not
g36820 not n17723 ; n17723_not
g36821 not n18056 ; n18056_not
g36822 not n20846 ; n20846_not
g36823 not n20864 ; n20864_not
g36824 not n20882 ; n20882_not
g36825 not n18074 ; n18074_not
g36826 not n29603 ; n29603_not
g36827 not n20918 ; n20918_not
g36828 not n20486 ; n20486_not
g36829 not n20477 ; n20477_not
g36830 not n30098 ; n30098_not
g36831 not n17840 ; n17840_not
g36832 not n20459 ; n20459_not
g36833 not n14168 ; n14168_not
g36834 not n12665 ; n12665_not
g36835 not n17930 ; n17930_not
g36836 not n30179 ; n30179_not
g36837 not n30197 ; n30197_not
g36838 not n12584 ; n12584_not
g36839 not n17813 ; n17813_not
g36840 not n13745 ; n13745_not
g36841 not n20657 ; n20657_not
g36842 not n20558 ; n20558_not
g36843 not n13970 ; n13970_not
g36844 not n20684 ; n20684_not
g36845 not n13880 ; n13880_not
g36846 not n30449 ; n30449_not
g36847 not n18227 ; n18227_not
g36848 not n18236 ; n18236_not
g36849 not n17570 ; n17570_not
g36850 not n30476 ; n30476_not
g36851 not n14339 ; n14339_not
g36852 not n18254 ; n18254_not
g36853 not n17552 ; n17552_not
g36854 not n21179 ; n21179_not
g36855 not n17534 ; n17534_not
g36856 not n12647 ; n12647_not
g36857 not n30557 ; n30557_not
g36858 not n17516 ; n17516_not
g36859 not n19370 ; n19370_not
g36860 not n30575 ; n30575_not
g36861 not n17480 ; n17480_not
g36862 not n12692 ; n12692_not
g36863 not n20936 ; n20936_not
g36864 not n20954 ; n20954_not
g36865 not n20972 ; n20972_not
g36866 not n18092 ; n18092_not
g36867 not n20990 ; n20990_not
g36868 not n29513 ; n29513_not
g36869 not n17237 ; n17237_not
g36870 not n18119 ; n18119_not
g36871 not n29450 ; n29450_not
g36872 not n29432 ; n29432_not
g36873 not n20189 ; n20189_not
g36874 not n17660 ; n17660_not
g36875 not n10946 ; n10946_not
g36876 not n18155 ; n18155_not
g36877 not n21098 ; n21098_not
g36878 not n17624 ; n17624_not
g36879 not n18182 ; n18182_not
g36880 not n17606 ; n17606_not
g36881 not n22583 ; n22583_not
g36882 not n31583 ; n31583_not
g36883 not n31628 ; n31628_not
g36884 not n31529 ; n31529_not
g36885 not n31646 ; n31646_not
g36886 not n16616 ; n16616_not
g36887 not n31673 ; n31673_not
g36888 not n18911 ; n18911_not
g36889 not n18902 ; n18902_not
g36890 not n27830 ; n27830_not
g36891 not n22655 ; n22655_not
g36892 not n14654 ; n14654_not
g36893 not n22664 ; n22664_not
g36894 not n22673 ; n22673_not
g36895 not n14663 ; n14663_not
g36896 not n31709 ; n31709_not
g36897 not n16814 ; n16814_not
g36898 not n22286 ; n22286_not
g36899 not n19091 ; n19091_not
g36900 not n28082 ; n28082_not
g36901 not n11783 ; n11783_not
g36902 not n16760 ; n16760_not
g36903 not n31493 ; n31493_not
g36904 not n16742 ; n16742_not
g36905 not n13574 ; n13574_not
g36906 not n12188 ; n12188_not
g36907 not n16715 ; n16715_not
g36908 not n11486 ; n11486_not
g36909 not n28028 ; n28028_not
g36910 not n19046 ; n19046_not
g36911 not n16670 ; n16670_not
g36912 not n31538 ; n31538_not
g36913 not n14177 ; n14177_not
g36914 not n18416 ; n18416_not
g36915 not n27605 ; n27605_not
g36916 not n22826 ; n22826_not
g36917 not n31970 ; n31970_not
g36918 not n22862 ; n22862_not
g36919 not n27551 ; n27551_not
g36920 not n13493 ; n13493_not
g36921 not n18272 ; n18272_not
g36922 not n18623 ; n18623_not
g36923 not n18614 ; n18614_not
g36924 not n32078 ; n32078_not
g36925 not n32087 ; n32087_not
g36926 not n10829 ; n10829_not
g36927 not n13358 ; n13358_not
g36928 not n14735 ; n14735_not
g36929 not n32096 ; n32096_not
g36930 not n22925 ; n22925_not
g36931 not n13538 ; n13538_not
g36932 not n14681 ; n14681_not
g36933 not n16580 ; n16580_not
g36934 not n27470 ; n27470_not
g36935 not n31781 ; n31781_not
g36936 not n16562 ; n16562_not
g36937 not n22718 ; n22718_not
g36938 not n22727 ; n22727_not
g36939 not n31790 ; n31790_not
g36940 not n31826 ; n31826_not
g36941 not n18218 ; n18218_not
g36942 not n27632 ; n27632_not
g36943 not n31844 ; n31844_not
g36944 not n10856 ; n10856_not
g36945 not n14708 ; n14708_not
g36946 not n31853 ; n31853_not
g36947 not n18731 ; n18731_not
g36948 not n22808 ; n22808_not
g36949 not n14447 ; n14447_not
g36950 not n28316 ; n28316_not
g36951 not n13529 ; n13529_not
g36952 not n19271 ; n19271_not
g36953 not n31394 ; n31394_not
g36954 not n14456 ; n14456_not
g36955 not n31457 ; n31457_not
g36956 not n10928 ; n10928_not
g36957 not n19253 ; n19253_not
g36958 not n19154 ; n19154_not
g36959 not n12656 ; n12656_not
g36960 not n16148 ; n16148_not
g36961 not n28217 ; n28217_not
g36962 not n14438 ; n14438_not
g36963 not n31376 ; n31376_not
g36964 not n16940 ; n16940_not
g36965 not n31448 ; n31448_not
g36966 not n21647 ; n21647_not
g36967 not n22196 ; n22196_not
g36968 not n28262 ; n28262_not
g36969 not n19235 ; n19235_not
g36970 not n21476 ; n21476_not
g36971 not n12359 ; n12359_not
g36972 not n31358 ; n31358_not
g36973 not n28280 ; n28280_not
g36974 not n28244 ; n28244_not
g36975 not n19362 ; n19362_not
g36976 not n25275 ; n25275_not
g36977 not n13485 ; n13485_not
g36978 not n18075 ; n18075_not
g36979 not n18363 ; n18363_not
g36980 not n25374 ; n25374_not
g36981 not n18066 ; n18066_not
g36982 not n15195 ; n15195_not
g36983 not n15816 ; n15816_not
g36984 not n13917 ; n13917_not
g36985 not n31197 ; n31197_not
g36986 not n18165 ; n18165_not
g36987 not n31782 ; n31782_not
g36988 not n11289 ; n11289_not
g36989 not n24447 ; n24447_not
g36990 not n24825 ; n24825_not
g36991 not n19092 ; n19092_not
g36992 not n31818 ; n31818_not
g36993 not n13584 ; n13584_not
g36994 not n18129 ; n18129_not
g36995 not n24834 ; n24834_not
g36996 not n19155 ; n19155_not
g36997 not n18219 ; n18219_not
g36998 not n18750 ; n18750_not
g36999 not n24852 ; n24852_not
g37000 not n15357 ; n15357_not
g37001 not n18822 ; n18822_not
g37002 not n13935 ; n13935_not
g37003 not n13656 ; n13656_not
g37004 not n31269 ; n31269_not
g37005 not n15375 ; n15375_not
g37006 not n13647 ; n13647_not
g37007 not n26904 ; n26904_not
g37008 not n18354 ; n18354_not
g37009 not n13548 ; n13548_not
g37010 not n26193 ; n26193_not
g37011 not n30198 ; n30198_not
g37012 not n15483 ; n15483_not
g37013 not n17940 ; n17940_not
g37014 not n18570 ; n18570_not
g37015 not n25392 ; n25392_not
g37016 not n31296 ; n31296_not
g37017 not n18480 ; n18480_not
g37018 not n25437 ; n25437_not
g37019 not n15843 ; n15843_not
g37020 not n15492 ; n15492_not
g37021 not n15177 ; n15177_not
g37022 not n11586 ; n11586_not
g37023 not n15708 ; n15708_not
g37024 not n20469 ; n20469_not
g37025 not n14088 ; n14088_not
g37026 not n18552 ; n18552_not
g37027 not n18534 ; n18534_not
g37028 not n18516 ; n18516_not
g37029 not n31908 ; n31908_not
g37030 not n15519 ; n15519_not
g37031 not n31359 ; n31359_not
g37032 not n25455 ; n25455_not
g37033 not n31980 ; n31980_not
g37034 not n20298 ; n20298_not
g37035 not n13953 ; n13953_not
g37036 not n26157 ; n26157_not
g37037 not n25329 ; n25329_not
g37038 not n18462 ; n18462_not
g37039 not n11829 ; n11829_not
g37040 not n25356 ; n25356_not
g37041 not n18651 ; n18651_not
g37042 not n13296 ; n13296_not
g37043 not n18633 ; n18633_not
g37044 not n20379 ; n20379_not
g37045 not n19263 ; n19263_not
g37046 not n24366 ; n24366_not
g37047 not n19326 ; n19326_not
g37048 not n19272 ; n19272_not
g37049 not n24348 ; n24348_not
g37050 not n32088 ; n32088_not
g37051 not n25572 ; n25572_not
g37052 not n24582 ; n24582_not
g37053 not n30828 ; n30828_not
g37054 not n30837 ; n30837_not
g37055 not n24645 ; n24645_not
g37056 not n15609 ; n15609_not
g37057 not n13575 ; n13575_not
g37058 not n12873 ; n12873_not
g37059 not n25563 ; n25563_not
g37060 not n12684 ; n12684_not
g37061 not n13755 ; n13755_not
g37062 not n13179 ; n13179_not
g37063 not n30783 ; n30783_not
g37064 not n15726 ; n15726_not
g37065 not n10596 ; n10596_not
g37066 not n24618 ; n24618_not
g37067 not n30756 ; n30756_not
g37068 not n25644 ; n25644_not
g37069 not n31089 ; n31089_not
g37070 not n19812 ; n19812_not
g37071 not n19551 ; n19551_not
g37072 not n30738 ; n30738_not
g37073 not n24717 ; n24717_not
g37074 not n31467 ; n31467_not
g37075 not n24906 ; n24906_not
g37076 not n15429 ; n15429_not
g37077 not n19641 ; n19641_not
g37078 not n15690 ; n15690_not
g37079 not n30972 ; n30972_not
g37080 not n30954 ; n30954_not
g37081 not n11964 ; n11964_not
g37082 not n31458 ; n31458_not
g37083 not n19623 ; n19623_not
g37084 not n18381 ; n18381_not
g37085 not n12855 ; n12855_not
g37086 not n24771 ; n24771_not
g37087 not n30882 ; n30882_not
g37088 not n19605 ; n19605_not
g37089 not n24663 ; n24663_not
g37090 not n19137 ; n19137_not
g37091 not n19731 ; n19731_not
g37092 not n30873 ; n30873_not
g37093 not n11649 ; n11649_not
g37094 not n30855 ; n30855_not
g37095 not n19074 ; n19074_not
g37096 not n31395 ; n31395_not
g37097 not n30558 ; n30558_not
g37098 not n25158 ; n25158_not
g37099 not n31683 ; n31683_not
g37100 not n11793 ; n11793_not
g37101 not n11919 ; n11919_not
g37102 not n25914 ; n25914_not
g37103 not n24492 ; n24492_not
g37104 not n30486 ; n30486_not
g37105 not n31638 ; n31638_not
g37106 not n24807 ; n24807_not
g37107 not n30468 ; n30468_not
g37108 not n25680 ; n25680_not
g37109 not n18615 ; n18615_not
g37110 not n31719 ; n31719_not
g37111 not n19911 ; n19911_not
g37112 not n19830 ; n19830_not
g37113 not n15537 ; n15537_not
g37114 not n18444 ; n18444_not
g37115 not n24465 ; n24465_not
g37116 not n18183 ; n18183_not
g37117 not n15627 ; n15627_not
g37118 not n25842 ; n25842_not
g37119 not n12756 ; n12756_not
g37120 not n25734 ; n25734_not
g37121 not n15564 ; n15564_not
g37122 not n19542 ; n19542_not
g37123 not n25941 ; n25941_not
g37124 not n13863 ; n13863_not
g37125 not n18426 ; n18426_not
g37126 not n30648 ; n30648_not
g37127 not n19515 ; n19515_not
g37128 not n18039 ; n18039_not
g37129 not n15672 ; n15672_not
g37130 not n12774 ; n12774_not
g37131 not n18930 ; n18930_not
g37132 not n18921 ; n18921_not
g37133 not n30576 ; n30576_not
g37134 not n31665 ; n31665_not
g37135 not n18336 ; n18336_not
g37136 not n10569 ; n10569_not
g37137 not n28533 ; n28533_not
g37138 not n17049 ; n17049_not
g37139 not n16185 ; n16185_not
g37140 not n21891 ; n21891_not
g37141 not n23484 ; n23484_not
g37142 not n28407 ; n28407_not
g37143 not n12378 ; n12378_not
g37144 not n28272 ; n28272_not
g37145 not n21990 ; n21990_not
g37146 not n28371 ; n28371_not
g37147 not n16194 ; n16194_not
g37148 not n14439 ; n14439_not
g37149 not n16941 ; n16941_not
g37150 not n16239 ; n16239_not
g37151 not n22089 ; n22089_not
g37152 not n28281 ; n28281_not
g37153 not n22098 ; n22098_not
g37154 not n23394 ; n23394_not
g37155 not n16923 ; n16923_not
g37156 not n28245 ; n28245_not
g37157 not n21549 ; n21549_not
g37158 not n22458 ; n22458_not
g37159 not n14826 ; n14826_not
g37160 not n28209 ; n28209_not
g37161 not n22188 ; n22188_not
g37162 not n16851 ; n16851_not
g37163 not n16257 ; n16257_not
g37164 not n14952 ; n14952_not
g37165 not n28173 ; n28173_not
g37166 not n27174 ; n27174_not
g37167 not n28146 ; n28146_not
g37168 not n23295 ; n23295_not
g37169 not n17238 ; n17238_not
g37170 not n17229 ; n17229_not
g37171 not n26670 ; n26670_not
g37172 not n16095 ; n16095_not
g37173 not n21585 ; n21585_not
g37174 not n23691 ; n23691_not
g37175 not n17184 ; n17184_not
g37176 not n17166 ; n17166_not
g37177 not n23673 ; n23673_not
g37178 not n23664 ; n23664_not
g37179 not n28920 ; n28920_not
g37180 not n21666 ; n21666_not
g37181 not n16149 ; n16149_not
g37182 not n28821 ; n28821_not
g37183 not n28812 ; n28812_not
g37184 not n26850 ; n26850_not
g37185 not n21387 ; n21387_not
g37186 not n21657 ; n21657_not
g37187 not n28740 ; n28740_not
g37188 not n28650 ; n28650_not
g37189 not n28632 ; n28632_not
g37190 not n21792 ; n21792_not
g37191 not n23556 ; n23556_not
g37192 not n16167 ; n16167_not
g37193 not n17067 ; n17067_not
g37194 not n16176 ; n16176_not
g37195 not n28551 ; n28551_not
g37196 not n26931 ; n26931_not
g37197 not n23529 ; n23529_not
g37198 not n27660 ; n27660_not
g37199 not n23079 ; n23079_not
g37200 not n27633 ; n27633_not
g37201 not n10857 ; n10857_not
g37202 not n14781 ; n14781_not
g37203 not n16428 ; n16428_not
g37204 not n16437 ; n16437_not
g37205 not n27606 ; n27606_not
g37206 not n22836 ; n22836_not
g37207 not n10839 ; n10839_not
g37208 not n16455 ; n16455_not
g37209 not n27327 ; n27327_not
g37210 not n14718 ; n14718_not
g37211 not n22863 ; n22863_not
g37212 not n27354 ; n27354_not
g37213 not n27381 ; n27381_not
g37214 not n16482 ; n16482_not
g37215 not n27507 ; n27507_not
g37216 not n14763 ; n14763_not
g37217 not n22449 ; n22449_not
g37218 not n27417 ; n27417_not
g37219 not n22908 ; n22908_not
g37220 not n27408 ; n27408_not
g37221 not n14745 ; n14745_not
g37222 not n22953 ; n22953_not
g37223 not n22944 ; n22944_not
g37224 not n27471 ; n27471_not
g37225 not n22926 ; n22926_not
g37226 not n14736 ; n14736_not
g37227 not n15096 ; n15096_not
g37228 not n22278 ; n22278_not
g37229 not n22296 ; n22296_not
g37230 not n28119 ; n28119_not
g37231 not n28092 ; n28092_not
g37232 not n16284 ; n16284_not
g37233 not n14619 ; n14619_not
g37234 not n11496 ; n11496_not
g37235 not n16644 ; n16644_not
g37236 not n22494 ; n22494_not
g37237 not n22557 ; n22557_not
g37238 not n16347 ; n16347_not
g37239 not n14637 ; n14637_not
g37240 not n23178 ; n23178_not
g37241 not n22584 ; n22584_not
g37242 not n23088 ; n23088_not
g37243 not n22962 ; n22962_not
g37244 not n14691 ; n14691_not
g37245 not n16563 ; n16563_not
g37246 not n27741 ; n27741_not
g37247 not n22683 ; n22683_not
g37248 not n16581 ; n16581_not
g37249 not n14673 ; n14673_not
g37250 not n16392 ; n16392_not
g37251 not n27237 ; n27237_not
g37252 not n27840 ; n27840_not
g37253 not n16419 ; n16419_not
g37254 not n16374 ; n16374_not
g37255 not n27219 ; n27219_not
g37256 not n16365 ; n16365_not
g37257 not n16626 ; n16626_not
g37258 not n27921 ; n27921_not
g37259 not n23907 ; n23907_not
g37260 not n17733 ; n17733_not
g37261 not n22485 ; n22485_not
g37262 not n17445 ; n17445_not
g37263 not n29811 ; n29811_not
g37264 not n10893 ; n10893_not
g37265 not n26508 ; n26508_not
g37266 not n21288 ; n21288_not
g37267 not n17535 ; n17535_not
g37268 not n29451 ; n29451_not
g37269 not n17553 ; n17553_not
g37270 not n29901 ; n29901_not
g37271 not n23925 ; n23925_not
g37272 not n26256 ; n26256_not
g37273 not n23835 ; n23835_not
g37274 not n29181 ; n29181_not
g37275 not n29172 ; n29172_not
g37276 not n29910 ; n29910_not
g37277 not n17715 ; n17715_not
g37278 not n12297 ; n12297_not
g37279 not n17571 ; n17571_not
g37280 not n15087 ; n15087_not
g37281 not n26454 ; n26454_not
g37282 not n29316 ; n29316_not
g37283 not n29622 ; n29622_not
g37284 not n17481 ; n17481_not
g37285 not n29271 ; n29271_not
g37286 not n14268 ; n14268_not
g37287 not n29253 ; n29253_not
g37288 not n26355 ; n26355_not
g37289 not n29703 ; n29703_not
g37290 not n17517 ; n17517_not
g37291 not n29244 ; n29244_not
g37292 not n26490 ; n26490_not
g37293 not n17463 ; n17463_not
g37294 not n29712 ; n29712_not
g37295 not n26292 ; n26292_not
g37296 not n24168 ; n24168_not
g37297 not n21189 ; n21189_not
g37298 not n23853 ; n23853_not
g37299 not n20586 ; n20586_not
g37300 not n17607 ; n17607_not
g37301 not n17850 ; n17850_not
g37302 not n26616 ; n26616_not
g37303 not n20559 ; n20559_not
g37304 not n17625 ; n17625_not
g37305 not n21396 ; n21396_not
g37306 not n11694 ; n11694_not
g37307 not n26094 ; n26094_not
g37308 not n17319 ; n17319_not
g37309 not n24285 ; n24285_not
g37310 not n14097 ; n14097_not
g37311 not n17904 ; n17904_not
g37312 not n26391 ; n26391_not
g37313 not n17148 ; n17148_not
g37314 not n15159 ; n15159_not
g37315 not n29370 ; n29370_not
g37316 not n29082 ; n29082_not
g37317 not n23745 ; n23745_not
g37318 not n20487 ; n20487_not
g37319 not n21459 ; n21459_not
g37320 not n29064 ; n29064_not
g37321 not n17382 ; n17382_not
g37322 not n26553 ; n26553_not
g37323 not n17823 ; n17823_not
g37324 not n29325 ; n29325_not
g37325 not n29361 ; n29361_not
g37326 not n17670 ; n17670_not
g37327 not n17364 ; n17364_not
g37328 not n29406 ; n29406_not
g37329 not n14178 ; n14178_not
g37330 not n23943 ; n23943_not
g37331 not n11766 ; n11766_not
g37332 not n26409 ; n26409_not
g37333 not n29136 ; n29136_not
g37334 not n17337 ; n17337_not
g37335 not n27931 ; n27931_not
g37336 not n13909 ; n13909_not
g37337 not n12199 ; n12199_not
g37338 not n23368 ; n23368_not
g37339 not n27850 ; n27850_not
g37340 not n15457 ; n15457_not
g37341 not n25546 ; n25546_not
g37342 not n15079 ; n15079_not
g37343 not n14647 ; n14647_not
g37344 not n26149 ; n26149_not
g37345 not n14593 ; n14593_not
g37346 not n13288 ; n13288_not
g37347 not n26383 ; n26383_not
g37348 not n29425 ; n29425_not
g37349 not n31576 ; n31576_not
g37350 not n29416 ; n29416_not
g37351 not n27904 ; n27904_not
g37352 not n31639 ; n31639_not
g37353 not n29380 ; n29380_not
g37354 not n29470 ; n29470_not
g37355 not n26185 ; n26185_not
g37356 not n31981 ; n31981_not
g37357 not n31945 ; n31945_not
g37358 not n27337 ; n27337_not
g37359 not n14719 ; n14719_not
g37360 not n13486 ; n13486_not
g37361 not n27364 ; n27364_not
g37362 not n12559 ; n12559_not
g37363 not n30199 ; n30199_not
g37364 not n25465 ; n25465_not
g37365 not n27391 ; n27391_not
g37366 not n14764 ; n14764_not
g37367 not n14179 ; n14179_not
g37368 not n14746 ; n14746_not
g37369 not n27436 ; n27436_not
g37370 not n27490 ; n27490_not
g37371 not n25771 ; n25771_not
g37372 not n27463 ; n27463_not
g37373 not n14089 ; n14089_not
g37374 not n13369 ; n13369_not
g37375 not n27823 ; n27823_not
g37376 not n29632 ; n29632_not
g37377 not n29641 ; n29641_not
g37378 not n27760 ; n27760_not
g37379 not n27715 ; n27715_not
g37380 not n29704 ; n29704_not
g37381 not n27706 ; n27706_not
g37382 not n14692 ; n14692_not
g37383 not n26284 ; n26284_not
g37384 not n31837 ; n31837_not
g37385 not n14674 ; n14674_not
g37386 not n13936 ; n13936_not
g37387 not n26176 ; n26176_not
g37388 not n29830 ; n29830_not
g37389 not n31882 ; n31882_not
g37390 not n27283 ; n27283_not
g37391 not n25492 ; n25492_not
g37392 not n25483 ; n25483_not
g37393 not n29902 ; n29902_not
g37394 not n26572 ; n26572_not
g37395 not n12883 ; n12883_not
g37396 not n29137 ; n29137_not
g37397 not n28750 ; n28750_not
g37398 not n12775 ; n12775_not
g37399 not n28741 ; n28741_not
g37400 not n28651 ; n28651_not
g37401 not n14926 ; n14926_not
g37402 not n25915 ; n25915_not
g37403 not n12685 ; n12685_not
g37404 not n12757 ; n12757_not
g37405 not n12892 ; n12892_not
g37406 not n31198 ; n31198_not
g37407 not n28570 ; n28570_not
g37408 not n28552 ; n28552_not
g37409 not n31189 ; n31189_not
g37410 not n25807 ; n25807_not
g37411 not n29182 ; n29182_not
g37412 not n14359 ; n14359_not
g37413 not n13657 ; n13657_not
g37414 not n15358 ; n15358_not
g37415 not n30658 ; n30658_not
g37416 not n26941 ; n26941_not
g37417 not n30649 ; n30649_not
g37418 not n28516 ; n28516_not
g37419 not n26653 ; n26653_not
g37420 not n30874 ; n30874_not
g37421 not n30919 ; n30919_not
g37422 not n11983 ; n11983_not
g37423 not n26671 ; n26671_not
g37424 not n14962 ; n14962_not
g37425 not n12496 ; n12496_not
g37426 not n30955 ; n30955_not
g37427 not n29083 ; n29083_not
g37428 not n30973 ; n30973_not
g37429 not n11947 ; n11947_not
g37430 not n26716 ; n26716_not
g37431 not n12478 ; n12478_not
g37432 not n26626 ; n26626_not
g37433 not n26077 ; n26077_not
g37434 not n28921 ; n28921_not
g37435 not n12766 ; n12766_not
g37436 not n12469 ; n12469_not
g37437 not n28840 ; n28840_not
g37438 not n28831 ; n28831_not
g37439 not n26590 ; n26590_not
g37440 not n28813 ; n28813_not
g37441 not n31099 ; n31099_not
g37442 not n31369 ; n31369_not
g37443 not n29281 ; n29281_not
g37444 not n12667 ; n12667_not
g37445 not n27148 ; n27148_not
g37446 not n28255 ; n28255_not
g37447 not n28228 ; n28228_not
g37448 not n13855 ; n13855_not
g37449 not n13585 ; n13585_not
g37450 not n29308 ; n29308_not
g37451 not n28183 ; n28183_not
g37452 not n10498 ; n10498_not
g37453 not n28156 ; n28156_not
g37454 not n31459 ; n31459_not
g37455 not n13576 ; n13576_not
g37456 not n25627 ; n25627_not
g37457 not n11668 ; n11668_not
g37458 not n28129 ; n28129_not
g37459 not n31486 ; n31486_not
g37460 not n13891 ; n13891_not
g37461 not n15439 ; n15439_not
g37462 not n26923 ; n26923_not
g37463 not n25582 ; n25582_not
g37464 not n27193 ; n27193_not
g37465 not n28075 ; n28075_not
g37466 not n25348 ; n25348_not
g37467 not n14908 ; n14908_not
g37468 not n25825 ; n25825_not
g37469 not n25429 ; n25429_not
g37470 not n28435 ; n28435_not
g37471 not n12379 ; n12379_not
g37472 not n14881 ; n14881_not
g37473 not n25564 ; n25564_not
g37474 not n25645 ; n25645_not
g37475 not n26482 ; n26482_not
g37476 not n13648 ; n13648_not
g37477 not n28273 ; n28273_not
g37478 not n31297 ; n31297_not
g37479 not n27058 ; n27058_not
g37480 not n28372 ; n28372_not
g37481 not n28354 ; n28354_not
g37482 not n27085 ; n27085_not
g37483 not n25735 ; n25735_not
g37484 not n11785 ; n11785_not
g37485 not n15385 ; n15385_not
g37486 not n30577 ; n30577_not
g37487 not n25294 ; n25294_not
g37488 not n25726 ; n25726_not
g37489 not n12649 ; n12649_not
g37490 not n25816 ; n25816_not
g37491 not n23179 ; n23179_not
g37492 not n17572 ; n17572_not
g37493 not n24691 ; n24691_not
g37494 not n16627 ; n16627_not
g37495 not n17554 ; n17554_not
g37496 not n17536 ; n17536_not
g37497 not n22639 ; n22639_not
g37498 not n15691 ; n15691_not
g37499 not n21577 ; n21577_not
g37500 not n19831 ; n19831_not
g37501 not n17518 ; n17518_not
g37502 not n23755 ; n23755_not
g37503 not n16294 ; n16294_not
g37504 not n17482 ; n17482_not
g37505 not n16483 ; n16483_not
g37506 not n20686 ; n20686_not
g37507 not n17671 ; n17671_not
g37508 not n24529 ; n24529_not
g37509 not n16456 ; n16456_not
g37510 not n24565 ; n24565_not
g37511 not n22576 ; n22576_not
g37512 not n24592 ; n24592_not
g37513 not n17653 ; n17653_not
g37514 not n22585 ; n22585_not
g37515 not n11884 ; n11884_not
g37516 not n17626 ; n17626_not
g37517 not n15709 ; n15709_not
g37518 not n24646 ; n24646_not
g37519 not n16825 ; n16825_not
g37520 not n18067 ; n18067_not
g37521 not n24664 ; n24664_not
g37522 not n17608 ; n17608_not
g37523 not n17590 ; n17590_not
g37524 not n19921 ; n19921_not
g37525 not n19624 ; n19624_not
g37526 not n24817 ; n24817_not
g37527 not n23692 ; n23692_not
g37528 not n17383 ; n17383_not
g37529 not n19606 ; n19606_not
g37530 not n24547 ; n24547_not
g37531 not n19570 ; n19570_not
g37532 not n17365 ; n17365_not
g37533 not n19552 ; n19552_not
g37534 not n23674 ; n23674_not
g37535 not n19534 ; n19534_not
g37536 not n24835 ; n24835_not
g37537 not n24853 ; n24853_not
g37538 not n17266 ; n17266_not
g37539 not n19516 ; n19516_not
g37540 not n18940 ; n18940_not
g37541 not n18922 ; n18922_not
g37542 not n18337 ; n18337_not
g37543 not n24727 ; n24727_not
g37544 not n19741 ; n19741_not
g37545 not n10894 ; n10894_not
g37546 not n17464 ; n17464_not
g37547 not n17338 ; n17338_not
g37548 not n23719 ; n23719_not
g37549 not n16582 ; n16582_not
g37550 not n23269 ; n23269_not
g37551 not n16096 ; n16096_not
g37552 not n24772 ; n24772_not
g37553 not n19660 ; n19660_not
g37554 not n15673 ; n15673_not
g37555 not n21298 ; n21298_not
g37556 not n19642 ; n19642_not
g37557 not n22684 ; n22684_not
g37558 not n20857 ; n20857_not
g37559 not n20668 ; n20668_not
g37560 not n23908 ; n23908_not
g37561 not n20875 ; n20875_not
g37562 not n16708 ; n16708_not
g37563 not n22369 ; n22369_not
g37564 not n22468 ; n22468_not
g37565 not n20893 ; n20893_not
g37566 not n24169 ; n24169_not
g37567 not n16663 ; n16663_not
g37568 not n11677 ; n11677_not
g37569 not n23557 ; n23557_not
g37570 not n17716 ; n17716_not
g37571 not n20596 ; n20596_not
g37572 not n11749 ; n11749_not
g37573 not n16807 ; n16807_not
g37574 not n20785 ; n20785_not
g37575 not n22297 ; n22297_not
g37576 not n23665 ; n23665_not
g37577 not n23890 ; n23890_not
g37578 not n11578 ; n11578_not
g37579 not n12586 ; n12586_not
g37580 not n11587 ; n11587_not
g37581 not n16771 ; n16771_not
g37582 not n17752 ; n17752_not
g37583 not n17761 ; n17761_not
g37584 not n16753 ; n16753_not
g37585 not n24088 ; n24088_not
g37586 not n20839 ; n20839_not
g37587 not n16735 ; n16735_not
g37588 not n11497 ; n11497_not
g37589 not n24349 ; n24349_not
g37590 not n17707 ; n17707_not
g37591 not n24367 ; n24367_not
g37592 not n16384 ; n16384_not
g37593 not n11398 ; n11398_not
g37594 not n18049 ; n18049_not
g37595 not n24394 ; n24394_not
g37596 not n20299 ; n20299_not
g37597 not n18085 ; n18085_not
g37598 not n16834 ; n16834_not
g37599 not n23845 ; n23845_not
g37600 not n24457 ; n24457_not
g37601 not n17770 ; n17770_not
g37602 not n22549 ; n22549_not
g37603 not n18184 ; n18184_not
g37604 not n22558 ; n22558_not
g37605 not n22198 ; n22198_not
g37606 not n11848 ; n11848_not
g37607 not n20929 ; n20929_not
g37608 not n17851 ; n17851_not
g37609 not n20569 ; n20569_not
g37610 not n20947 ; n20947_not
g37611 not n20965 ; n20965_not
g37612 not n20983 ; n20983_not
g37613 not n10669 ; n10669_not
g37614 not n16645 ; n16645_not
g37615 not n24295 ; n24295_not
g37616 not n17419 ; n17419_not
g37617 not n11659 ; n11659_not
g37618 not n20488 ; n20488_not
g37619 not n23872 ; n23872_not
g37620 not n15844 ; n15844_not
g37621 not n17914 ; n17914_not
g37622 not n17824 ; n17824_not
g37623 not n19093 ; n19093_not
g37624 not n18391 ; n18391_not
g37625 not n18724 ; n18724_not
g37626 not n18373 ; n18373_not
g37627 not n19165 ; n19165_not
g37628 not n16528 ; n16528_not
g37629 not n21829 ; n21829_not
g37630 not n16492 ; n16492_not
g37631 not n19183 ; n19183_not
g37632 not n15628 ; n15628_not
g37633 not n21838 ; n21838_not
g37634 not n11479 ; n11479_not
g37635 not n25276 ; n25276_not
g37636 not n21658 ; n21658_not
g37637 not n19192 ; n19192_not
g37638 not n23377 ; n23377_not
g37639 not n18706 ; n18706_not
g37640 not n16564 ; n16564_not
g37641 not n23494 ; n23494_not
g37642 not n19246 ; n19246_not
g37643 not n24493 ; n24493_not
g37644 not n16195 ; n16195_not
g37645 not n21667 ; n21667_not
g37646 not n21388 ; n21388_not
g37647 not n24952 ; n24952_not
g37648 not n23575 ; n23575_not
g37649 not n18670 ; n18670_not
g37650 not n23395 ; n23395_not
g37651 not n22918 ; n22918_not
g37652 not n18814 ; n18814_not
g37653 not n15574 ; n15574_not
g37654 not n18931 ; n18931_not
g37655 not n10885 ; n10885_not
g37656 not n15592 ; n15592_not
g37657 not n21775 ; n21775_not
g37658 not n16546 ; n16546_not
g37659 not n25096 ; n25096_not
g37660 not n15565 ; n15565_not
g37661 not n21739 ; n21739_not
g37662 not n16177 ; n16177_not
g37663 not n10966 ; n10966_not
g37664 not n10858 ; n10858_not
g37665 not n19039 ; n19039_not
g37666 not n18409 ; n18409_not
g37667 not n16159 ; n16159_not
g37668 not n17077 ; n17077_not
g37669 not n15547 ; n15547_not
g37670 not n21649 ; n21649_not
g37671 not n23566 ; n23566_not
g37672 not n22927 ; n22927_not
g37673 not n17095 ; n17095_not
g37674 not n25159 ; n25159_not
g37675 not n10588 ; n10588_not
g37676 not n22477 ; n22477_not
g37677 not n19336 ; n19336_not
g37678 not n22864 ; n22864_not
g37679 not n21928 ; n21928_not
g37680 not n19363 ; n19363_not
g37681 not n23647 ; n23647_not
g37682 not n10786 ; n10786_not
g37683 not n19264 ; n19264_not
g37684 not n21937 ; n21937_not
g37685 not n15493 ; n15493_not
g37686 not n25375 ; n25375_not
g37687 not n19390 ; n19390_not
g37688 not n19129 ; n19129_not
g37689 not n16267 ; n16267_not
g37690 not n18616 ; n18616_not
g37691 not n17248 ; n17248_not
g37692 not n23458 ; n23458_not
g37693 not n15484 ; n15484_not
g37694 not n19471 ; n19471_not
g37695 not n15646 ; n15646_not
g37696 not n23296 ; n23296_not
g37697 not n21973 ; n21973_not
g37698 not n21874 ; n21874_not
g37699 not n16249 ; n16249_not
g37700 not n23593 ; n23593_not
g37701 not n21496 ; n21496_not
g37702 not n10984 ; n10984_not
g37703 not n17158 ; n17158_not
g37704 not n22855 ; n22855_not
g37705 not n18256 ; n18256_not
g37706 not n24934 ; n24934_not
g37707 not n22954 ; n22954_not
g37708 not n17185 ; n17185_not
g37709 not n16924 ; n16924_not
g37710 not n24907 ; n24907_not
g37711 not n10759 ; n10759_not
g37712 not n10778 ; n10778_not
g37713 not n28364 ; n28364_not
g37714 not n11669 ; n11669_not
g37715 not n21857 ; n21857_not
g37716 not n14297 ; n14297_not
g37717 not n28346 ; n28346_not
g37718 not n21785 ; n21785_not
g37719 not n23468 ; n23468_not
g37720 not n17726 ; n17726_not
g37721 not n25817 ; n25817_not
g37722 not n23396 ; n23396_not
g37723 not n21983 ; n21983_not
g37724 not n12299 ; n12299_not
g37725 not n28670 ; n28670_not
g37726 not n29525 ; n29525_not
g37727 not n26960 ; n26960_not
g37728 not n29633 ; n29633_not
g37729 not n28526 ; n28526_not
g37730 not n23927 ; n23927_not
g37731 not n21884 ; n21884_not
g37732 not n28571 ; n28571_not
g37733 not n26465 ; n26465_not
g37734 not n28382 ; n28382_not
g37735 not n23936 ; n23936_not
g37736 not n16835 ; n16835_not
g37737 not n28337 ; n28337_not
g37738 not n23891 ; n23891_not
g37739 not n28607 ; n28607_not
g37740 not n29651 ; n29651_not
g37741 not n16196 ; n16196_not
g37742 not n14279 ; n14279_not
g37743 not n28508 ; n28508_not
g37744 not n28157 ; n28157_not
g37745 not n15764 ; n15764_not
g37746 not n23558 ; n23558_not
g37747 not n23882 ; n23882_not
g37748 not n14909 ; n14909_not
g37749 not n29660 ; n29660_not
g37750 not n21956 ; n21956_not
g37751 not n17393 ; n17393_not
g37752 not n13748 ; n13748_not
g37753 not n17195 ; n17195_not
g37754 not n29219 ; n29219_not
g37755 not n21578 ; n21578_not
g37756 not n16925 ; n16925_not
g37757 not n26672 ; n26672_not
g37758 not n17465 ; n17465_not
g37759 not n23729 ; n23729_not
g37760 not n14927 ; n14927_not
g37761 not n16907 ; n16907_not
g37762 not n21668 ; n21668_not
g37763 not n29282 ; n29282_not
g37764 not n29291 ; n29291_not
g37765 not n26870 ; n26870_not
g37766 not n21659 ; n21659_not
g37767 not n21299 ; n21299_not
g37768 not n17078 ; n17078_not
g37769 not n29093 ; n29093_not
g37770 not n28274 ; n28274_not
g37771 not n21389 ; n21389_not
g37772 not n21479 ; n21479_not
g37773 not n17348 ; n17348_not
g37774 not n27185 ; n27185_not
g37775 not n23666 ; n23666_not
g37776 not n15944 ; n15944_not
g37777 not n23675 ; n23675_not
g37778 not n16268 ; n16268_not
g37779 not n26717 ; n26717_not
g37780 not n17366 ; n17366_not
g37781 not n28256 ; n28256_not
g37782 not n17384 ; n17384_not
g37783 not n29039 ; n29039_not
g37784 not n29183 ; n29183_not
g37785 not n24188 ; n24188_not
g37786 not n26924 ; n26924_not
g37787 not n17672 ; n17672_not
g37788 not n29435 ; n29435_not
g37789 not n28751 ; n28751_not
g37790 not n29444 ; n29444_not
g37791 not n28184 ; n28184_not
g37792 not n16178 ; n16178_not
g37793 not n26942 ; n26942_not
g37794 not n21758 ; n21758_not
g37795 not n14792 ; n14792_not
g37796 not n29507 ; n29507_not
g37797 not n23846 ; n23846_not
g37798 not n27149 ; n27149_not
g37799 not n28715 ; n28715_not
g37800 not n16952 ; n16952_not
g37801 not n28850 ; n28850_not
g37802 not n16295 ; n16295_not
g37803 not n28238 ; n28238_not
g37804 not n14972 ; n14972_not
g37805 not n16358 ; n16358_not
g37806 not n16880 ; n16880_not
g37807 not n28832 ; n28832_not
g37808 not n21677 ; n21677_not
g37809 not n16934 ; n16934_not
g37810 not n26906 ; n26906_not
g37811 not n29318 ; n29318_not
g37812 not n26096 ; n26096_not
g37813 not n26564 ; n26564_not
g37814 not n29417 ; n29417_not
g37815 not n17663 ; n17663_not
g37816 not n23387 ; n23387_not
g37817 not n23828 ; n23828_not
g37818 not n25619 ; n25619_not
g37819 not n25763 ; n25763_not
g37820 not n27770 ; n27770_not
g37821 not n22955 ; n22955_not
g37822 not n19337 ; n19337_not
g37823 not n31289 ; n31289_not
g37824 not n25745 ; n25745_not
g37825 not n24917 ; n24917_not
g37826 not n31298 ; n31298_not
g37827 not n24944 ; n24944_not
g37828 not n19292 ; n19292_not
g37829 not n25727 ; n25727_not
g37830 not n27734 ; n27734_not
g37831 not n19265 ; n19265_not
g37832 not n24494 ; n24494_not
g37833 not n27455 ; n27455_not
g37834 not n25718 ; n25718_not
g37835 not n15386 ; n15386_not
g37836 not n15395 ; n15395_not
g37837 not n24980 ; n24980_not
g37838 not n31388 ; n31388_not
g37839 not n19193 ; n19193_not
g37840 not n30974 ; n30974_not
g37841 not n30992 ; n30992_not
g37842 not n19625 ; n19625_not
g37843 not n24818 ; n24818_not
g37844 not n12866 ; n12866_not
g37845 not n19607 ; n19607_not
g37846 not n30893 ; n30893_not
g37847 not n22685 ; n22685_not
g37848 not n19571 ; n19571_not
g37849 not n12677 ; n12677_not
g37850 not n19553 ; n19553_not
g37851 not n14747 ; n14747_not
g37852 not n19535 ; n19535_not
g37853 not n24836 ; n24836_not
g37854 not n22856 ; n22856_not
g37855 not n24854 ; n24854_not
g37856 not n12776 ; n12776_not
g37857 not n19481 ; n19481_not
g37858 not n24881 ; n24881_not
g37859 not n19463 ; n19463_not
g37860 not n18338 ; n18338_not
g37861 not n18347 ; n18347_not
g37862 not n15449 ; n15449_not
g37863 not n15548 ; n15548_not
g37864 not n18743 ; n18743_not
g37865 not n10589 ; n10589_not
g37866 not n31757 ; n31757_not
g37867 not n18716 ; n18716_not
g37868 not n15467 ; n15467_not
g37869 not n25493 ; n25493_not
g37870 not n25295 ; n25295_not
g37871 not n31928 ; n31928_not
g37872 not n31964 ; n31964_not
g37873 not n25475 ; n25475_not
g37874 not n25349 ; n25349_not
g37875 not n31919 ; n31919_not
g37876 not n18671 ; n18671_not
g37877 not n13496 ; n13496_not
g37878 not n18626 ; n18626_not
g37879 not n25385 ; n25385_not
g37880 not n27536 ; n27536_not
g37881 not n13397 ; n13397_not
g37882 not n18590 ; n18590_not
g37883 not n27707 ; n27707_not
g37884 not n25673 ; n25673_not
g37885 not n19175 ; n19175_not
g37886 not n13586 ; n13586_not
g37887 not n14837 ; n14837_not
g37888 not n25655 ; n25655_not
g37889 not n18392 ; n18392_not
g37890 not n31496 ; n31496_not
g37891 not n18374 ; n18374_not
g37892 not n19067 ; n19067_not
g37893 not n19049 ; n19049_not
g37894 not n18419 ; n18419_not
g37895 not n31568 ; n31568_not
g37896 not n31586 ; n31586_not
g37897 not n10886 ; n10886_not
g37898 not n15593 ; n15593_not
g37899 not n10877 ; n10877_not
g37900 not n18905 ; n18905_not
g37901 not n16547 ; n16547_not
g37902 not n18851 ; n18851_not
g37903 not n15575 ; n15575_not
g37904 not n18761 ; n18761_not
g37905 not n31775 ; n31775_not
g37906 not n25565 ; n25565_not
g37907 not n16529 ; n16529_not
g37908 not n20579 ; n20579_not
g37909 not n17852 ; n17852_not
g37910 not n29921 ; n29921_not
g37911 not n11777 ; n11777_not
g37912 not n17870 ; n17870_not
g37913 not n13883 ; n13883_not
g37914 not n17915 ; n17915_not
g37915 not n15188 ; n15188_not
g37916 not n11795 ; n11795_not
g37917 not n17951 ; n17951_not
g37918 not n18068 ; n18068_not
g37919 not n23945 ; n23945_not
g37920 not n13919 ; n13919_not
g37921 not n24458 ; n24458_not
g37922 not n18158 ; n18158_not
g37923 not n15791 ; n15791_not
g37924 not n22559 ; n22559_not
g37925 not n14774 ; n14774_not
g37926 not n20795 ; n20795_not
g37927 not n29705 ; n29705_not
g37928 not n20777 ; n20777_not
g37929 not n29750 ; n29750_not
g37930 not n23648 ; n23648_not
g37931 not n29570 ; n29570_not
g37932 not n26366 ; n26366_not
g37933 not n11579 ; n11579_not
g37934 not n11597 ; n11597_not
g37935 not n29903 ; n29903_not
g37936 not n29741 ; n29741_not
g37937 not n29930 ; n29930_not
g37938 not n17762 ; n17762_not
g37939 not n12569 ; n12569_not
g37940 not n17834 ; n17834_not
g37941 not n26267 ; n26267_not
g37942 not n25781 ; n25781_not
g37943 not n16646 ; n16646_not
g37944 not n20597 ; n20597_not
g37945 not n12596 ; n12596_not
g37946 not n30659 ; n30659_not
g37947 not n30677 ; n30677_not
g37948 not n19841 ; n19841_not
g37949 not n27851 ; n27851_not
g37950 not n15692 ; n15692_not
g37951 not n27365 ; n27365_not
g37952 not n12758 ; n12758_not
g37953 not n12686 ; n12686_not
g37954 not n22658 ; n22658_not
g37955 not n19805 ; n19805_not
g37956 not n19760 ; n19760_not
g37957 not n14765 ; n14765_not
g37958 not n19742 ; n19742_not
g37959 not n30848 ; n30848_not
g37960 not n27392 ; n27392_not
g37961 not n30875 ; n30875_not
g37962 not n25961 ; n25961_not
g37963 not n30866 ; n30866_not
g37964 not n19724 ; n19724_not
g37965 not n25952 ; n25952_not
g37966 not n30938 ; n30938_not
g37967 not n14657 ; n14657_not
g37968 not n19661 ; n19661_not
g37969 not n24782 ; n24782_not
g37970 not n22676 ; n22676_not
g37971 not n19643 ; n19643_not
g37972 not n15368 ; n15368_not
g37973 not n27932 ; n27932_not
g37974 not n24638 ; n24638_not
g37975 not n27338 ; n27338_not
g37976 not n24647 ; n24647_not
g37977 not n16385 ; n16385_not
g37978 not n18248 ; n18248_not
g37979 not n11867 ; n11867_not
g37980 not n11975 ; n11975_not
g37981 not n12749 ; n12749_not
g37982 not n27905 ; n27905_not
g37983 not n19931 ; n19931_not
g37984 not n11876 ; n11876_not
g37985 not n27537 ; n27537_not
g37986 not n27960 ; n27960_not
g37987 not n10869 ; n10869_not
g37988 not n16575 ; n16575_not
g37989 not n22857 ; n22857_not
g37990 not n28284 ; n28284_not
g37991 not n19518 ; n19518_not
g37992 not n16908 ; n16908_not
g37993 not n27519 ; n27519_not
g37994 not n11688 ; n11688_not
g37995 not n28257 ; n28257_not
g37996 not n28347 ; n28347_not
g37997 not n16557 ; n16557_not
g37998 not n27735 ; n27735_not
g37999 not n16845 ; n16845_not
g38000 not n27564 ; n27564_not
g38001 not n22839 ; n22839_not
g38002 not n10887 ; n10887_not
g38003 not n27771 ; n27771_not
g38004 not n16593 ; n16593_not
g38005 not n16962 ; n16962_not
g38006 not n22596 ; n22596_not
g38007 not n16944 ; n16944_not
g38008 not n14658 ; n14658_not
g38009 not n16548 ; n16548_not
g38010 not n27753 ; n27753_not
g38011 not n19482 ; n19482_not
g38012 not n19536 ; n19536_not
g38013 not n13749 ; n13749_not
g38014 not n30993 ; n30993_not
g38015 not n26088 ; n26088_not
g38016 not n30948 ; n30948_not
g38017 not n30885 ; n30885_not
g38018 not n30858 ; n30858_not
g38019 not n19734 ; n19734_not
g38020 not n19743 ; n19743_not
g38021 not n12777 ; n12777_not
g38022 not n19815 ; n19815_not
g38023 not n10986 ; n10986_not
g38024 not n12696 ; n12696_not
g38025 not n30696 ; n30696_not
g38026 not n19392 ; n19392_not
g38027 not n13947 ; n13947_not
g38028 not n20499 ; n20499_not
g38029 not n18078 ; n18078_not
g38030 not n18177 ; n18177_not
g38031 not n30399 ; n30399_not
g38032 not n13884 ; n13884_not
g38033 not n13758 ; n13758_not
g38034 not n13695 ; n13695_not
g38035 not n18195 ; n18195_not
g38036 not n30489 ; n30489_not
g38037 not n30498 ; n30498_not
g38038 not n13848 ; n13848_not
g38039 not n19338 ; n19338_not
g38040 not n19932 ; n19932_not
g38041 not n19914 ; n19914_not
g38042 not n30678 ; n30678_not
g38043 not n18906 ; n18906_not
g38044 not n18924 ; n18924_not
g38045 not n31686 ; n31686_not
g38046 not n31695 ; n31695_not
g38047 not n18807 ; n18807_not
g38048 not n31785 ; n31785_not
g38049 not n18762 ; n18762_not
g38050 not n18753 ; n18753_not
g38051 not n18717 ; n18717_not
g38052 not n31929 ; n31929_not
g38053 not n31956 ; n31956_not
g38054 not n31974 ; n31974_not
g38055 not n18681 ; n18681_not
g38056 not n13497 ; n13497_not
g38057 not n13299 ; n13299_not
g38058 not n13398 ; n13398_not
g38059 not n12858 ; n12858_not
g38060 not n19374 ; n19374_not
g38061 not n19356 ; n19356_not
g38062 not n19347 ; n19347_not
g38063 not n18357 ; n18357_not
g38064 not n19275 ; n19275_not
g38065 not n18816 ; n18816_not
g38066 not n19239 ; n19239_not
g38067 not n19194 ; n19194_not
g38068 not n31398 ; n31398_not
g38069 not n19176 ; n19176_not
g38070 not n19158 ; n19158_not
g38071 not n19077 ; n19077_not
g38072 not n31497 ; n31497_not
g38073 not n31587 ; n31587_not
g38074 not n31596 ; n31596_not
g38075 not n21696 ; n21696_not
g38076 not n28851 ; n28851_not
g38077 not n28950 ; n28950_not
g38078 not n17178 ; n17178_not
g38079 not n21588 ; n21588_not
g38080 not n13929 ; n13929_not
g38081 not n16836 ; n16836_not
g38082 not n29058 ; n29058_not
g38083 not n17259 ; n17259_not
g38084 not n21399 ; n21399_not
g38085 not n17349 ; n17349_not
g38086 not n29148 ; n29148_not
g38087 not n29157 ; n29157_not
g38088 not n29166 ; n29166_not
g38089 not n17439 ; n17439_not
g38090 not n29238 ; n29238_not
g38091 not n21966 ; n21966_not
g38092 not n28248 ; n28248_not
g38093 not n28446 ; n28446_not
g38094 not n28509 ; n28509_not
g38095 not n16890 ; n16890_not
g38096 not n21867 ; n21867_not
g38097 not n28536 ; n28536_not
g38098 not n28545 ; n28545_not
g38099 not n28590 ; n28590_not
g38100 not n28608 ; n28608_not
g38101 not n28626 ; n28626_not
g38102 not n17088 ; n17088_not
g38103 not n28707 ; n28707_not
g38104 not n28716 ; n28716_not
g38105 not n21768 ; n21768_not
g38106 not n28752 ; n28752_not
g38107 not n28770 ; n28770_not
g38108 not n14298 ; n14298_not
g38109 not n29355 ; n29355_not
g38110 not n29652 ; n29652_not
g38111 not n29670 ; n29670_not
g38112 not n20796 ; n20796_not
g38113 not n29733 ; n29733_not
g38114 not n29805 ; n29805_not
g38115 not n17736 ; n17736_not
g38116 not n29742 ; n29742_not
g38117 not n29913 ; n29913_not
g38118 not n29931 ; n29931_not
g38119 not n17763 ; n17763_not
g38120 not n17664 ; n17664_not
g38121 not n12588 ; n12588_not
g38122 not n17835 ; n17835_not
g38123 not n20598 ; n20598_not
g38124 not n17475 ; n17475_not
g38125 not n17493 ; n17493_not
g38126 not n17529 ; n17529_not
g38127 not n17547 ; n17547_not
g38128 not n17565 ; n17565_not
g38129 not n29319 ; n29319_not
g38130 not n17583 ; n17583_not
g38131 not n17619 ; n17619_not
g38132 not n17646 ; n17646_not
g38133 not n29436 ; n29436_not
g38134 not n17268 ; n17268_not
g38135 not n29454 ; n29454_not
g38136 not n29463 ; n29463_not
g38137 not n29490 ; n29490_not
g38138 not n29508 ; n29508_not
g38139 not n15198 ; n15198_not
g38140 not n26871 ; n26871_not
g38141 not n24459 ; n24459_not
g38142 not n27078 ; n27078_not
g38143 not n24486 ; n24486_not
g38144 not n25692 ; n25692_not
g38145 not n24981 ; n24981_not
g38146 not n14856 ; n14856_not
g38147 not n15387 ; n15387_not
g38148 not n24945 ; n24945_not
g38149 not n23847 ; n23847_not
g38150 not n25728 ; n25728_not
g38151 not n22569 ; n22569_not
g38152 not n10599 ; n10599_not
g38153 not n24927 ; n24927_not
g38154 not n15639 ; n15639_not
g38155 not n24495 ; n24495_not
g38156 not n23685 ; n23685_not
g38157 not n25782 ; n25782_not
g38158 not n24189 ; n24189_not
g38159 not n25575 ; n25575_not
g38160 not n14883 ; n14883_not
g38161 not n15576 ; n15576_not
g38162 not n11679 ; n11679_not
g38163 not n14874 ; n14874_not
g38164 not n23559 ; n23559_not
g38165 not n15594 ; n15594_not
g38166 not n24387 ; n24387_not
g38167 not n26682 ; n26682_not
g38168 not n26169 ; n26169_not
g38169 not n25665 ; n25665_not
g38170 not n25854 ; n25854_not
g38171 not n24819 ; n24819_not
g38172 not n25908 ; n25908_not
g38173 not n25836 ; n25836_not
g38174 not n26547 ; n26547_not
g38175 not n10779 ; n10779_not
g38176 not n14973 ; n14973_not
g38177 not n11958 ; n11958_not
g38178 not n14793 ; n14793_not
g38179 not n22785 ; n22785_not
g38180 not n24567 ; n24567_not
g38181 not n25953 ; n25953_not
g38182 not n23595 ; n23595_not
g38183 not n25962 ; n25962_not
g38184 not n16368 ; n16368_not
g38185 not n26646 ; n26646_not
g38186 not n24891 ; n24891_not
g38187 not n27249 ; n27249_not
g38188 not n25827 ; n25827_not
g38189 not n14838 ; n14838_not
g38190 not n22497 ; n22497_not
g38191 not n16449 ; n16449_not
g38192 not n24657 ; n24657_not
g38193 not n24684 ; n24684_not
g38194 not n14991 ; n14991_not
g38195 not n14784 ; n14784_not
g38196 not n23838 ; n23838_not
g38197 not n26538 ; n26538_not
g38198 not n25890 ; n25890_not
g38199 not n14928 ; n14928_not
g38200 not n11787 ; n11787_not
g38201 not n26943 ; n26943_not
g38202 not n14559 ; n14559_not
g38203 not n15468 ; n15468_not
g38204 not n25458 ; n25458_not
g38205 not n26448 ; n26448_not
g38206 not n25359 ; n25359_not
g38207 not n25539 ; n25539_not
g38208 not n25476 ; n25476_not
g38209 not n10698 ; n10698_not
g38210 not n25188 ; n25188_not
g38211 not n23937 ; n23937_not
g38212 not n26349 ; n26349_not
g38213 not n25494 ; n25494_not
g38214 not n25296 ; n25296_not
g38215 not n26439 ; n26439_not
g38216 not n27483 ; n27483_not
g38217 not n22884 ; n22884_not
g38218 not n15486 ; n15486_not
g38219 not n23469 ; n23469_not
g38220 not n24639 ; n24639_not
g38221 not n23388 ; n23388_not
g38222 not n14892 ; n14892_not
g38223 not n14946 ; n14946_not
g38224 not n23938 ; n23938_not
g38225 not n14992 ; n14992_not
g38226 not n30598 ; n30598_not
g38227 not n12697 ; n12697_not
g38228 not n29473 ; n29473_not
g38229 not n17737 ; n17737_not
g38230 not n19924 ; n19924_not
g38231 not n19933 ; n19933_not
g38232 not n29455 ; n29455_not
g38233 not n22993 ; n22993_not
g38234 not n29806 ; n29806_not
g38235 not n29671 ; n29671_not
g38236 not n14839 ; n14839_not
g38237 not n19771 ; n19771_not
g38238 not n25981 ; n25981_not
g38239 not n19339 ; n19339_not
g38240 not n30499 ; n30499_not
g38241 not n28357 ; n28357_not
g38242 not n29824 ; n29824_not
g38243 not n28285 ; n28285_not
g38244 not n12778 ; n12778_not
g38245 not n25765 ; n25765_not
g38246 not n19753 ; n19753_not
g38247 not n16909 ; n16909_not
g38248 not n16918 ; n16918_not
g38249 not n28267 ; n28267_not
g38250 not n23659 ; n23659_not
g38251 not n15685 ; n15685_not
g38252 not n23839 ; n23839_not
g38253 not n23965 ; n23965_not
g38254 not n20779 ; n20779_not
g38255 not n30697 ; n30697_not
g38256 not n17665 ; n17665_not
g38257 not n30679 ; n30679_not
g38258 not n27187 ; n27187_not
g38259 not n26386 ; n26386_not
g38260 not n23569 ; n23569_not
g38261 not n29734 ; n29734_not
g38262 not n10789 ; n10789_not
g38263 not n26953 ; n26953_not
g38264 not n28708 ; n28708_not
g38265 not n30787 ; n30787_not
g38266 not n23389 ; n23389_not
g38267 not n28735 ; n28735_not
g38268 not n25837 ; n25837_not
g38269 not n30796 ; n30796_not
g38270 not n29743 ; n29743_not
g38271 not n26377 ; n26377_not
g38272 not n29923 ; n29923_not
g38273 not n14299 ; n14299_not
g38274 not n28447 ; n28447_not
g38275 not n13858 ; n13858_not
g38276 not n26485 ; n26485_not
g38277 not n21895 ; n21895_not
g38278 not n17638 ; n17638_not
g38279 not n26098 ; n26098_not
g38280 not n26476 ; n26476_not
g38281 not n17818 ; n17818_not
g38282 not n29608 ; n29608_not
g38283 not n22489 ; n22489_not
g38284 not n17944 ; n17944_not
g38285 not n26188 ; n26188_not
g38286 not n11797 ; n11797_not
g38287 not n28771 ; n28771_not
g38288 not n26287 ; n26287_not
g38289 not n17881 ; n17881_not
g38290 not n14875 ; n14875_not
g38291 not n28564 ; n28564_not
g38292 not n28519 ; n28519_not
g38293 not n23479 ; n23479_not
g38294 not n17863 ; n17863_not
g38295 not n17845 ; n17845_not
g38296 not n26278 ; n26278_not
g38297 not n28555 ; n28555_not
g38298 not n14893 ; n14893_not
g38299 not n28537 ; n28537_not
g38300 not n17836 ; n17836_not
g38301 not n28807 ; n28807_not
g38302 not n28645 ; n28645_not
g38303 not n17692 ; n17692_not
g38304 not n13867 ; n13867_not
g38305 not n24379 ; n24379_not
g38306 not n21994 ; n21994_not
g38307 not n11599 ; n11599_not
g38308 not n19816 ; n19816_not
g38309 not n19735 ; n19735_not
g38310 not n16189 ; n16189_not
g38311 not n28627 ; n28627_not
g38312 not n21796 ; n21796_not
g38313 not n29509 ; n29509_not
g38314 not n13894 ; n13894_not
g38315 not n29950 ; n29950_not
g38316 not n12895 ; n12895_not
g38317 not n15199 ; n15199_not
g38318 not n28249 ; n28249_not
g38319 not n16945 ; n16945_not
g38320 not n24478 ; n24478_not
g38321 not n28609 ; n28609_not
g38322 not n28429 ; n28429_not
g38323 not n21949 ; n21949_not
g38324 not n18187 ; n18187_not
g38325 not n23497 ; n23497_not
g38326 not n16963 ; n16963_not
g38327 not n24487 ; n24487_not
g38328 not n16882 ; n16882_not
g38329 not n27088 ; n27088_not
g38330 not n18196 ; n18196_not
g38331 not n29176 ; n29176_not
g38332 not n17377 ; n17377_not
g38333 not n18916 ; n18916_not
g38334 not n14668 ; n14668_not
g38335 not n31696 ; n31696_not
g38336 not n26863 ; n26863_not
g38337 not n14758 ; n14758_not
g38338 not n22678 ; n22678_not
g38339 not n29167 ; n29167_not
g38340 not n14686 ; n14686_not
g38341 not n24676 ; n24676_not
g38342 not n27772 ; n27772_not
g38343 not n22966 ; n22966_not
g38344 not n18808 ; n18808_not
g38345 not n27439 ; n27439_not
g38346 not n31786 ; n31786_not
g38347 not n31795 ; n31795_not
g38348 not n27736 ; n27736_not
g38349 not n31399 ; n31399_not
g38350 not n29239 ; n29239_not
g38351 not n19177 ; n19177_not
g38352 not n24973 ; n24973_not
g38353 not n17458 ; n17458_not
g38354 not n19168 ; n19168_not
g38355 not n25666 ; n25666_not
g38356 not n22399 ; n22399_not
g38357 not n26665 ; n26665_not
g38358 not n18853 ; n18853_not
g38359 not n26683 ; n26683_not
g38360 not n25648 ; n25648_not
g38361 not n24982 ; n24982_not
g38362 not n22588 ; n22588_not
g38363 not n18358 ; n18358_not
g38364 not n24892 ; n24892_not
g38365 not n31597 ; n31597_not
g38366 not n16585 ; n16585_not
g38367 not n27808 ; n27808_not
g38368 not n23587 ; n23587_not
g38369 not n31957 ; n31957_not
g38370 not n25297 ; n25297_not
g38371 not n29086 ; n29086_not
g38372 not n25477 ; n25477_not
g38373 not n13489 ; n13489_not
g38374 not n26773 ; n26773_not
g38375 not n25468 ; n25468_not
g38376 not n31984 ; n31984_not
g38377 not n15478 ; n15478_not
g38378 not n29077 ; n29077_not
g38379 not n15847 ; n15847_not
g38380 not n29059 ; n29059_not
g38381 not n16837 ; n16837_not
g38382 not n12499 ; n12499_not
g38383 not n13399 ; n13399_not
g38384 not n26827 ; n26827_not
g38385 not n22894 ; n22894_not
g38386 not n17188 ; n17188_not
g38387 not n22867 ; n22867_not
g38388 not n18772 ; n18772_not
g38389 not n22948 ; n22948_not
g38390 not n27457 ; n27457_not
g38391 not n16567 ; n16567_not
g38392 not n15559 ; n15559_not
g38393 not n27718 ; n27718_not
g38394 not n25549 ; n25549_not
g38395 not n22939 ; n22939_not
g38396 not n29149 ; n29149_not
g38397 not n31858 ; n31858_not
g38398 not n14785 ; n14785_not
g38399 not n31894 ; n31894_not
g38400 not n27682 ; n27682_not
g38401 not n18718 ; n18718_not
g38402 not n18709 ; n18709_not
g38403 not n25288 ; n25288_not
g38404 not n26746 ; n26746_not
g38405 not n17359 ; n17359_not
g38406 not n26881 ; n26881_not
g38407 not n23785 ; n23785_not
g38408 not n11689 ; n11689_not
g38409 not n30958 ; n30958_not
g38410 not n27268 ; n27268_not
g38411 not n19654 ; n19654_not
g38412 not n19672 ; n19672_not
g38413 not n24847 ; n24847_not
g38414 not n15649 ; n15649_not
g38415 not n16693 ; n16693_not
g38416 not n12886 ; n12886_not
g38417 not n24874 ; n24874_not
g38418 not n23767 ; n23767_not
g38419 not n14794 ; n14794_not
g38420 not n23758 ; n23758_not
g38421 not n25918 ; n25918_not
g38422 not n24793 ; n24793_not
g38423 not n30967 ; n30967_not
g38424 not n30994 ; n30994_not
g38425 not n19636 ; n19636_not
g38426 not n15667 ; n15667_not
g38427 not n19618 ; n19618_not
g38428 not n19582 ; n19582_not
g38429 not n24829 ; n24829_not
g38430 not n25891 ; n25891_not
g38431 not n19564 ; n19564_not
g38432 not n25855 ; n25855_not
g38433 not n19546 ; n19546_not
g38434 not n28870 ; n28870_not
g38435 not n19465 ; n19465_not
g38436 not n12958 ; n12958_not
g38437 not n25747 ; n25747_not
g38438 not n30868 ; n30868_not
g38439 not n30859 ; n30859_not
g38440 not n19285 ; n19285_not
g38441 not n16639 ; n16639_not
g38442 not n16459 ; n16459_not
g38443 not n24946 ; n24946_not
g38444 not n27961 ; n27961_not
g38445 not n19249 ; n19249_not
g38446 not n16369 ; n16369_not
g38447 not n25963 ; n25963_not
g38448 not n16477 ; n16477_not
g38449 not n15397 ; n15397_not
g38450 not n29392 ; n29392_not
g38451 not n22597 ; n22597_not
g38452 not n25972 ; n25972_not
g38453 not n30895 ; n30895_not
g38454 not n19492 ; n19492_not
g38455 not n19690 ; n19690_not
g38456 not n29383 ; n29383_not
g38457 not n19078 ; n19078_not
g38458 not n19717 ; n19717_not
g38459 not n24757 ; n24757_not
g38460 not n15379 ; n15379_not
g38461 not n24739 ; n24739_not
g38462 not n26647 ; n26647_not
g38463 not n25756 ; n25756_not
g38464 not n14939 ; n14939_not
g38465 not n29627 ; n29627_not
g38466 not n29357 ; n29357_not
g38467 not n29078 ; n29078_not
g38468 not n17639 ; n17639_not
g38469 not n29393 ; n29393_not
g38470 not n26567 ; n26567_not
g38471 not n26648 ; n26648_not
g38472 not n17468 ; n17468_not
g38473 not n29258 ; n29258_not
g38474 not n23867 ; n23867_not
g38475 not n14993 ; n14993_not
g38476 not n26684 ; n26684_not
g38477 not n29195 ; n29195_not
g38478 not n29564 ; n29564_not
g38479 not n26468 ; n26468_not
g38480 not n17387 ; n17387_not
g38481 not n29267 ; n29267_not
g38482 not n29276 ; n29276_not
g38483 not n29573 ; n29573_not
g38484 not n29168 ; n29168_not
g38485 not n29483 ; n29483_not
g38486 not n26459 ; n26459_not
g38487 not n29474 ; n29474_not
g38488 not n17369 ; n17369_not
g38489 not n23768 ; n23768_not
g38490 not n23885 ; n23885_not
g38491 not n23678 ; n23678_not
g38492 not n29609 ; n29609_not
g38493 not n17675 ; n17675_not
g38494 not n28925 ; n28925_not
g38495 not n23786 ; n23786_not
g38496 not n26558 ; n26558_not
g38497 not n24866 ; n24866_not
g38498 not n18890 ; n18890_not
g38499 not n18962 ; n18962_not
g38500 not n31598 ; n31598_not
g38501 not n24992 ; n24992_not
g38502 not n19088 ; n19088_not
g38503 not n25658 ; n25658_not
g38504 not n18386 ; n18386_not
g38505 not n25667 ; n25667_not
g38506 not n24974 ; n24974_not
g38507 not n13598 ; n13598_not
g38508 not n24965 ; n24965_not
g38509 not n19187 ; n19187_not
g38510 not n18368 ; n18368_not
g38511 not n25757 ; n25757_not
g38512 not n19169 ; n19169_not
g38513 not n18980 ; n18980_not
g38514 not n25469 ; n25469_not
g38515 not n19493 ; n19493_not
g38516 not n12995 ; n12995_not
g38517 not n12896 ; n12896_not
g38518 not n25856 ; n25856_not
g38519 not n19529 ; n19529_not
g38520 not n25874 ; n25874_not
g38521 not n15668 ; n15668_not
g38522 not n30977 ; n30977_not
g38523 not n18485 ; n18485_not
g38524 not n18539 ; n18539_not
g38525 not n18557 ; n18557_not
g38526 not n18575 ; n18575_not
g38527 not n18467 ; n18467_not
g38528 not n25397 ; n25397_not
g38529 not n25388 ; n25388_not
g38530 not n15479 ; n15479_not
g38531 not n18629 ; n18629_not
g38532 not n18638 ; n18638_not
g38533 not n18656 ; n18656_not
g38534 not n31985 ; n31985_not
g38535 not n18692 ; n18692_not
g38536 not n31967 ; n31967_not
g38537 not n31949 ; n31949_not
g38538 not n25487 ; n25487_not
g38539 not n18449 ; n18449_not
g38540 not n31886 ; n31886_not
g38541 not n31859 ; n31859_not
g38542 not n31796 ; n31796_not
g38543 not n15569 ; n15569_not
g38544 not n18782 ; n18782_not
g38545 not n18809 ; n18809_not
g38546 not n18836 ; n18836_not
g38547 not n31697 ; n31697_not
g38548 not n18917 ; n18917_not
g38549 not n15587 ; n15587_not
g38550 not n24488 ; n24488_not
g38551 not n19709 ; n19709_not
g38552 not n17738 ; n17738_not
g38553 not n13949 ; n13949_not
g38554 not n13994 ; n13994_not
g38555 not n17972 ; n17972_not
g38556 not n17954 ; n17954_not
g38557 not n11798 ; n11798_not
g38558 not n17909 ; n17909_not
g38559 not n17891 ; n17891_not
g38560 not n24299 ; n24299_not
g38561 not n17873 ; n17873_not
g38562 not n17855 ; n17855_not
g38563 not n12599 ; n12599_not
g38564 not n17819 ; n17819_not
g38565 not n17774 ; n17774_not
g38566 not n29924 ; n29924_not
g38567 not n17756 ; n17756_not
g38568 not n29843 ; n29843_not
g38569 not n29825 ; n29825_not
g38570 not n17747 ; n17747_not
g38571 not n29807 ; n29807_not
g38572 not n26369 ; n26369_not
g38573 not n29744 ; n29744_not
g38574 not n29726 ; n29726_not
g38575 not n29708 ; n29708_not
g38576 not n29690 ; n29690_not
g38577 not n30959 ; n30959_not
g38578 not n24758 ; n24758_not
g38579 not n30896 ; n30896_not
g38580 not n19736 ; n19736_not
g38581 not n25973 ; n25973_not
g38582 not n30797 ; n30797_not
g38583 not n25919 ; n25919_not
g38584 not n19826 ; n19826_not
g38585 not n30698 ; n30698_not
g38586 not n15695 ; n15695_not
g38587 not n19844 ; n19844_not
g38588 not n25946 ; n25946_not
g38589 not n19853 ; n19853_not
g38590 not n11969 ; n11969_not
g38591 not n11789 ; n11789_not
g38592 not n19871 ; n19871_not
g38593 not n11978 ; n11978_not
g38594 not n19376 ; n19376_not
g38595 not n12698 ; n12698_not
g38596 not n19907 ; n19907_not
g38597 not n30599 ; n30599_not
g38598 not n24677 ; n24677_not
g38599 not n11879 ; n11879_not
g38600 not n19925 ; n19925_not
g38601 not n13859 ; n13859_not
g38602 not n19790 ; n19790_not
g38603 not n28556 ; n28556_not
g38604 not n26972 ; n26972_not
g38605 not n23489 ; n23489_not
g38606 not n14876 ; n14876_not
g38607 not n21878 ; n21878_not
g38608 not n28493 ; n28493_not
g38609 not n28448 ; n28448_not
g38610 not n28439 ; n28439_not
g38611 not n21977 ; n21977_not
g38612 not n27089 ; n27089_not
g38613 not n28385 ; n28385_not
g38614 not n14849 ; n14849_not
g38615 not n16991 ; n16991_not
g38616 not n28286 ; n28286_not
g38617 not n16199 ; n16199_not
g38618 not n16973 ; n16973_not
g38619 not n23399 ; n23399_not
g38620 not n16928 ; n16928_not
g38621 not n26891 ; n26891_not
g38622 not n28826 ; n28826_not
g38623 not n21689 ; n21689_not
g38624 not n28808 ; n28808_not
g38625 not n26909 ; n26909_not
g38626 not n28790 ; n28790_not
g38627 not n26846 ; n26846_not
g38628 not n26918 ; n26918_not
g38629 not n28745 ; n28745_not
g38630 not n26936 ; n26936_not
g38631 not n28736 ; n28736_not
g38632 not n26954 ; n26954_not
g38633 not n28664 ; n28664_not
g38634 not n28646 ; n28646_not
g38635 not n21779 ; n21779_not
g38636 not n28628 ; n28628_not
g38637 not n28583 ; n28583_not
g38638 not n28574 ; n28574_not
g38639 not n14894 ; n14894_not
g38640 not n16586 ; n16586_not
g38641 not n16478 ; n16478_not
g38642 not n27836 ; n27836_not
g38643 not n27809 ; n27809_not
g38644 not n14669 ; n14669_not
g38645 not n22985 ; n22985_not
g38646 not n22688 ; n22688_not
g38647 not n14687 ; n14687_not
g38648 not n22697 ; n22697_not
g38649 not n27746 ; n27746_not
g38650 not n27449 ; n27449_not
g38651 not n27683 ; n27683_not
g38652 not n27476 ; n27476_not
g38653 not n27656 ; n27656_not
g38654 not n27629 ; n27629_not
g38655 not n22679 ; n22679_not
g38656 not n27575 ; n27575_not
g38657 not n22895 ; n22895_not
g38658 not n22877 ; n22877_not
g38659 not n28268 ; n28268_not
g38660 not n16289 ; n16289_not
g38661 not n16892 ; n16892_not
g38662 not n16856 ; n16856_not
g38663 not n16379 ; n16379_not
g38664 not n16838 ; n16838_not
g38665 not n16397 ; n16397_not
g38666 not n16829 ; n16829_not
g38667 not n28088 ; n28088_not
g38668 not n14696 ; n14696_not
g38669 not n27269 ; n27269_not
g38670 not n16685 ; n16685_not
g38671 not n16649 ; n16649_not
g38672 not n27296 ; n27296_not
g38673 not n27728 ; n27728_not
g38674 not n22589 ; n22589_not
g38675 not n16568 ; n16568_not
g38676 not n14768 ; n14768_not
g38677 not n22598 ; n22598_not
g38678 not n13976 ; n13976_not
g38679 not n21599 ; n21599_not
g38680 not n26855 ; n26855_not
g38681 not n28943 ; n28943_not
g38682 not n17874 ; n17874_not
g38683 not n17892 ; n17892_not
g38684 not n18918 ; n18918_not
g38685 not n28467 ; n28467_not
g38686 not n25587 ; n25587_not
g38687 not n26793 ; n26793_not
g38688 not n26694 ; n26694_not
g38689 not n25776 ; n25776_not
g38690 not n25578 ; n25578_not
g38691 not n17829 ; n17829_not
g38692 not n28575 ; n28575_not
g38693 not n17388 ; n17388_not
g38694 not n22977 ; n22977_not
g38695 not n22995 ; n22995_not
g38696 not n23967 ; n23967_not
g38697 not n17856 ; n17856_not
g38698 not n17937 ; n17937_not
g38699 not n13995 ; n13995_not
g38700 not n13977 ; n13977_not
g38701 not n17982 ; n17982_not
g38702 not n15786 ; n15786_not
g38703 not n28953 ; n28953_not
g38704 not n16929 ; n16929_not
g38705 not n17739 ; n17739_not
g38706 not n13896 ; n13896_not
g38707 not n24957 ; n24957_not
g38708 not n18990 ; n18990_not
g38709 not n14949 ; n14949_not
g38710 not n27495 ; n27495_not
g38711 not n28764 ; n28764_not
g38712 not n20898 ; n20898_not
g38713 not n29628 ; n29628_not
g38714 not n29646 ; n29646_not
g38715 not n28737 ; n28737_not
g38716 not n23949 ; n23949_not
g38717 not n26955 ; n26955_not
g38718 not n27477 ; n27477_not
g38719 not n29709 ; n29709_not
g38720 not n23985 ; n23985_not
g38721 not n18738 ; n18738_not
g38722 not n29781 ; n29781_not
g38723 not n28665 ; n28665_not
g38724 not n28647 ; n28647_not
g38725 not n29826 ; n29826_not
g38726 not n29844 ; n29844_not
g38727 not n16497 ; n16497_not
g38728 not n14688 ; n14688_not
g38729 not n18756 ; n18756_not
g38730 not n27675 ; n27675_not
g38731 not n27729 ; n27729_not
g38732 not n29916 ; n29916_not
g38733 not n29925 ; n29925_not
g38734 not n31797 ; n31797_not
g38735 not n27747 ; n27747_not
g38736 not n18783 ; n18783_not
g38737 not n15939 ; n15939_not
g38738 not n26856 ; n26856_not
g38739 not n27765 ; n27765_not
g38740 not n28593 ; n28593_not
g38741 not n30888 ; n30888_not
g38742 not n30897 ; n30897_not
g38743 not n27954 ; n27954_not
g38744 not n24759 ; n24759_not
g38745 not n16398 ; n16398_not
g38746 not n24786 ; n24786_not
g38747 not n15669 ; n15669_not
g38748 not n30978 ; n30978_not
g38749 not n30987 ; n30987_not
g38750 not n18369 ; n18369_not
g38751 not n14787 ; n14787_not
g38752 not n16794 ; n16794_not
g38753 not n19278 ; n19278_not
g38754 not n16776 ; n16776_not
g38755 not n24939 ; n24939_not
g38756 not n27981 ; n27981_not
g38757 not n25884 ; n25884_not
g38758 not n19539 ; n19539_not
g38759 not n16758 ; n16758_not
g38760 not n18396 ; n18396_not
g38761 not n24867 ; n24867_not
g38762 not n22968 ; n22968_not
g38763 not n12897 ; n12897_not
g38764 not n26766 ; n26766_not
g38765 not n19494 ; n19494_not
g38766 not n19476 ; n19476_not
g38767 not n25758 ; n25758_not
g38768 not n19368 ; n19368_not
g38769 not n25659 ; n25659_not
g38770 not n18954 ; n18954_not
g38771 not n25785 ; n25785_not
g38772 not n13878 ; n13878_not
g38773 not n15597 ; n15597_not
g38774 not n11898 ; n11898_not
g38775 not n19971 ; n19971_not
g38776 not n16992 ; n16992_not
g38777 not n16479 ; n16479_not
g38778 not n19953 ; n19953_not
g38779 not n11997 ; n11997_not
g38780 not n19926 ; n19926_not
g38781 not n24687 ; n24687_not
g38782 not n16974 ; n16974_not
g38783 not n26739 ; n26739_not
g38784 not n19872 ; n19872_not
g38785 not n19854 ; n19854_not
g38786 not n19098 ; n19098_not
g38787 not n15696 ; n15696_not
g38788 not n24975 ; n24975_not
g38789 not n19836 ; n19836_not
g38790 not n28269 ; n28269_not
g38791 not n18387 ; n18387_not
g38792 not n19791 ; n19791_not
g38793 not n30798 ; n30798_not
g38794 not n29079 ; n29079_not
g38795 not n16884 ; n16884_not
g38796 not n25956 ; n25956_not
g38797 not n19746 ; n19746_not
g38798 not n25974 ; n25974_not
g38799 not n14769 ; n14769_not
g38800 not n17955 ; n17955_not
g38801 not n16857 ; n16857_not
g38802 not n16848 ; n16848_not
g38803 not n17685 ; n17685_not
g38804 not n29565 ; n29565_not
g38805 not n18468 ; n18468_not
g38806 not n28809 ; n28809_not
g38807 not n25398 ; n25398_not
g38808 not n29277 ; n29277_not
g38809 not n23787 ; n23787_not
g38810 not n18558 ; n18558_not
g38811 not n29394 ; n29394_not
g38812 not n18639 ; n18639_not
g38813 not n18657 ; n18657_not
g38814 not n23589 ; n23589_not
g38815 not n26847 ; n26847_not
g38816 not n26586 ; n26586_not
g38817 not n18576 ; n18576_not
g38818 not n28845 ; n28845_not
g38819 not n23769 ; n23769_not
g38820 not n23877 ; n23877_not
g38821 not n27558 ; n27558_not
g38822 not n17649 ; n17649_not
g38823 not n20988 ; n20988_not
g38824 not n14967 ; n14967_not
g38825 not n26658 ; n26658_not
g38826 not n22689 ; n22689_not
g38827 not n22896 ; n22896_not
g38828 not n28827 ; n28827_not
g38829 not n29574 ; n29574_not
g38830 not n29259 ; n29259_not
g38831 not n18486 ; n18486_not
g38832 not n24994 ; n24994_not
g38833 not n16849 ; n16849_not
g38834 not n28594 ; n28594_not
g38835 not n13978 ; n13978_not
g38836 not n29971 ; n29971_not
g38837 not n15598 ; n15598_not
g38838 not n17776 ; n17776_not
g38839 not n29980 ; n29980_not
g38840 not n18793 ; n18793_not
g38841 not n27973 ; n27973_not
g38842 not n27964 ; n27964_not
g38843 not n27595 ; n27595_not
g38844 not n20989 ; n20989_not
g38845 not n26992 ; n26992_not
g38846 not n28846 ; n28846_not
g38847 not n15787 ; n15787_not
g38848 not n16894 ; n16894_not
g38849 not n26497 ; n26497_not
g38850 not n18658 ; n18658_not
g38851 not n14986 ; n14986_not
g38852 not n24958 ; n24958_not
g38853 not n19963 ; n19963_not
g38854 not n19297 ; n19297_not
g38855 not n26596 ; n26596_not
g38856 not n18469 ; n18469_not
g38857 not n14968 ; n14968_not
g38858 not a[10] ; a[10]_not
g38859 not n16876 ; n16876_not
g38860 not n27748 ; n27748_not
g38861 not n16777 ; n16777_not
g38862 not n25588 ; n25588_not
g38863 not n14869 ; n14869_not
g38864 not n26695 ; n26695_not
g38865 not n18838 ; n18838_not
g38866 not n26848 ; n26848_not
g38867 not n25399 ; n25399_not
g38868 not n28954 ; n28954_not
g38869 not n17965 ; n17965_not
g38870 not n24796 ; n24796_not
g38871 not n16399 ; n16399_not
g38872 not n17929 ; n17929_not
g38873 not n18955 ; n18955_not
g38874 not n25687 ; n25687_not
g38875 not n26776 ; n26776_not
g38876 not n29449 ; n29449_not
g38877 not n27388 ; n27388_not
g38878 not n28828 ; n28828_not
g38879 not n28396 ; n28396_not
g38880 not n16858 ; n16858_not
g38881 not n26299 ; n26299_not
g38882 not n28963 ; n28963_not
g38883 not n17785 ; n17785_not
g38884 not n28459 ; n28459_not
g38885 not n24949 ; n24949_not
g38886 not n18559 ; n18559_not
g38887 not n27568 ; n27568_not
g38888 not n28099 ; n28099_not
g38889 not n27928 ; n27928_not
g38890 not n17398 ; n17398_not
g38891 not n17839 ; n17839_not
g38892 not n14887 ; n14887_not
g38893 not n16993 ; n16993_not
g38894 not n25777 ; n25777_not
g38895 not n13996 ; n13996_not
g38896 not n28468 ; n28468_not
g38897 not n16795 ; n16795_not
g38898 not n28783 ; n28783_not
g38899 not n19855 ; n19855_not
g38900 not n12997 ; n12997_not
g38901 not n19819 ; n19819_not
g38902 not n26965 ; n26965_not
g38903 not n18388 ; n18388_not
g38904 not n23878 ; n23878_not
g38905 not n27649 ; n27649_not
g38906 not n16678 ; n16678_not
g38907 not n29773 ; n29773_not
g38908 not n19873 ; n19873_not
g38909 not n27694 ; n27694_not
g38910 not n27874 ; n27874_not
g38911 not n29629 ; n29629_not
g38912 not n18685 ; n18685_not
g38913 not n28666 ; n28666_not
g38914 not n15985 ; n15985_not
g38915 not n27478 ; n27478_not
g38916 not n25984 ; n25984_not
g38917 not n19099 ; n19099_not
g38918 not n28864 ; n28864_not
g38919 not n29278 ; n29278_not
g38920 not n19477 ; n19477_not
g38921 not n26398 ; n26398_not
g38922 not n16939 ; n16939_not
g38923 not n15499 ; n15499_not
g38924 not n18577 ; n18577_not
g38925 not n29665 ; n29665_not
g38926 not n16957 ; n16957_not
g38927 not n29719 ; n29719_not
g38928 not n28279 ; n28279_not
g38929 not n28774 ; n28774_not
g38930 not n27676 ; n27676_not
g38931 not n19837 ; n19837_not
g38932 not n29647 ; n29647_not
g38933 not n29872 ; n29872_not
g38934 not n26749 ; n26749_not
g38935 not n29593 ; n29593_not
g38936 not n29863 ; n29863_not
g38937 not n20899 ; n20899_not
g38938 not n16975 ; n16975_not
g38939 not n16498 ; n16498_not
g38940 not n26929 ; n26929_not
g38941 not n29881 ; n29881_not
g38942 not n27847 ; n27847_not
g38943 not n24895 ; n24895_not
g38944 not n29845 ; n29845_not
g38945 not n18784 ; n18784_not
g38946 not n18748 ; n18748_not
g38947 not n26677 ; n26677_not
g38948 not n17983 ; n17983_not
g38949 not n19936 ; n19936_not
g38950 not n27991 ; n27991_not
g38951 not n29377 ; n29377_not
g38952 not n26659 ; n26659_not
g38953 not n18487 ; n18487_not
g38954 not n29296 ; n29296_not
g38955 not n26884 ; n26884_not
g38956 not n14779 ; n14779_not
g38957 not n24877 ; n24877_not
g38958 not n16759 ; n16759_not
g38959 not n18983 ; n18983_not
g38960 not n19838 ; n19838_not
g38961 not a[11] ; a[11]_not
g38962 not a[20] ; a[20]_not
g38963 not n24698 ; n24698_not
g38964 not n26579 ; n26579_not
g38965 not n17678 ; n17678_not
g38966 not n28865 ; n28865_not
g38967 not n19829 ; n19829_not
g38968 not n29387 ; n29387_not
g38969 not n22979 ; n22979_not
g38970 not n28982 ; n28982_not
g38971 not n29369 ; n29369_not
g38972 not n24599 ; n24599_not
g38973 not n25967 ; n25967_not
g38974 not n19964 ; n19964_not
g38975 not n28847 ; n28847_not
g38976 not n28199 ; n28199_not
g38977 not n19946 ; n19946_not
g38978 not n28964 ; n28964_not
g38979 not n28397 ; n28397_not
g38980 not n24968 ; n24968_not
g38981 not n28379 ; n28379_not
g38982 not n16958 ; n16958_not
g38983 not n17894 ; n17894_not
g38984 not n25787 ; n25787_not
g38985 not n17588 ; n17588_not
g38986 not n27947 ; n27947_not
g38987 not n29297 ; n29297_not
g38988 not n18785 ; n18785_not
g38989 not n25796 ; n25796_not
g38990 not n29864 ; n29864_not
g38991 not n29882 ; n29882_not
g38992 not n18749 ; n18749_not
g38993 not n28928 ; n28928_not
g38994 not n15986 ; n15986_not
g38995 not n25877 ; n25877_not
g38996 not n14897 ; n14897_not
g38997 not n26993 ; n26993_not
g38998 not n16886 ; n16886_not
g38999 not n16778 ; n16778_not
g39000 not n27758 ; n27758_not
g39001 not n28883 ; n28883_not
g39002 not n29981 ; n29981_not
g39003 not n17768 ; n17768_not
g39004 not n29594 ; n29594_not
g39005 not n27488 ; n27488_not
g39006 not n17498 ; n17498_not
g39007 not n31979 ; n31979_not
g39008 not n29648 ; n29648_not
g39009 not n26948 ; n26948_not
g39010 not n29666 ; n29666_not
g39011 not n25769 ; n25769_not
g39012 not n27659 ; n27659_not
g39013 not n29684 ; n29684_not
g39014 not n18695 ; n18695_not
g39015 not n28775 ; n28775_not
g39016 not n19478 ; n19478_not
g39017 not n23879 ; n23879_not
g39018 not n27677 ; n27677_not
g39019 not n19487 ; n19487_not
g39020 not n16499 ; n16499_not
g39021 not n27992 ; n27992_not
g39022 not n27695 ; n27695_not
g39023 not n22889 ; n22889_not
g39024 not n22799 ; n22799_not
g39025 not n26966 ; n26966_not
g39026 not n29819 ; n29819_not
g39027 not n24797 ; n24797_not
g39028 not n18929 ; n18929_not
g39029 not n17993 ; n17993_not
g39030 not n13979 ; n13979_not
g39031 not n25697 ; n25697_not
g39032 not n18938 ; n18938_not
g39033 not n29468 ; n29468_not
g39034 not n26777 ; n26777_not
g39035 not n24779 ; n24779_not
g39036 not n28469 ; n28469_not
g39037 not n27965 ; n27965_not
g39038 not n28793 ; n28793_not
g39039 not n17399 ; n17399_not
g39040 not n18884 ; n18884_not
g39041 not n14969 ; n14969_not
g39042 not n27578 ; n27578_not
g39043 not n23987 ; n23987_not
g39044 not n25589 ; n25589_not
g39045 not n18965 ; n18965_not
g39046 not n16796 ; n16796_not
g39047 not n26849 ; n26849_not
g39048 not n26696 ; n26696_not
g39049 not n18498 ; n18498_not
g39050 not n24888 ; n24888_not
g39051 not n14898 ; n14898_not
g39052 not a[12] ; a[12]_not
g39053 not n19677 ; n19677_not
g39054 not n27948 ; n27948_not
g39055 not n19587 ; n19587_not
g39056 not n25887 ; n25887_not
g39057 not n19569 ; n19569_not
g39058 not n28884 ; n28884_not
g39059 not n17589 ; n17589_not
g39060 not n29289 ; n29289_not
g39061 not n28866 ; n28866_not
g39062 not n19749 ; n19749_not
g39063 not n25878 ; n25878_not
g39064 not n29298 ; n29298_not
g39065 not n19758 ; n19758_not
g39066 not n19695 ; n19695_not
g39067 not n19776 ; n19776_not
g39068 not n27894 ; n27894_not
g39069 not n25698 ; n25698_not
g39070 not n16896 ; n16896_not
g39071 not n19497 ; n19497_not
g39072 not n27984 ; n27984_not
g39073 not n17499 ; n17499_not
g39074 not n19659 ; n19659_not
g39075 not n29946 ; n29946_not
g39076 not n18786 ; n18786_not
g39077 not n29982 ; n29982_not
g39078 not n27759 ; n27759_not
g39079 not n27579 ; n27579_not
g39080 not n28794 ; n28794_not
g39081 not n18696 ; n18696_not
g39082 not n28569 ; n28569_not
g39083 not n18885 ; n18885_not
g39084 not n17697 ; n17697_not
g39085 not n17868 ; n17868_not
g39086 not n28497 ; n28497_not
g39087 not n29469 ; n29469_not
g39088 not n12999 ; n12999_not
g39089 not n17958 ; n17958_not
g39090 not n13989 ; n13989_not
g39091 not n22998 ; n22998_not
g39092 not n17787 ; n17787_not
g39093 not n27777 ; n27777_not
g39094 not n28389 ; n28389_not
g39095 not n18993 ; n18993_not
g39096 not a[21] ; a[21]_not
g39097 not n29595 ; n29595_not
g39098 not n16878 ; n16878_not
g39099 not n27489 ; n27489_not
g39100 not n23898 ; n23898_not
g39101 not a[30] ; a[30]_not
g39102 not n29667 ; n29667_not
g39103 not n28929 ; n28929_not
g39104 not n29685 ; n29685_not
g39105 not n23799 ; n23799_not
g39106 not n28677 ; n28677_not
g39107 not n31899 ; n31899_not
g39108 not n27687 ; n27687_not
g39109 not n28659 ; n28659_not
g39110 not n26967 ; n26967_not
g39111 not n29829 ; n29829_not
g39112 not n29838 ; n29838_not
g39113 not n31998 ; n31998_not
g39114 not n18678 ; n18678_not
g39115 not n29865 ; n29865_not
g39116 not n29856 ; n29856_not
g39117 not n29883 ; n29883_not
g39118 not n25797 ; n25797_not
g39119 not n22899 ; n22899_not
g39120 not n18777 ; n18777_not
g39121 not n19893 ; n19893_not
g39122 not n16968 ; n16968_not
g39123 not n26859 ; n26859_not
g39124 not n24978 ; n24978_not
g39125 not n29397 ; n29397_not
g39126 not n16986 ; n16986_not
g39127 not n28965 ; n28965_not
g39128 not n19965 ; n19965_not
g39129 not n18597 ; n18597_not
g39130 not n16959 ; n16959_not
g39131 not n21999 ; n21999_not
g39132 not n19992 ; n19992_not
g39133 not n19866 ; n19866_not
g39134 not n28983 ; n28983_not
g39135 not n19848 ; n19848_not
g39136 not n27867 ; n27867_not
g39137 not n29398 ; n29398_not
g39138 not a[13] ; a[13]_not
g39139 not n18778 ; n18778_not
g39140 not n22999 ; n22999_not
g39141 not n27976 ; n27976_not
g39142 not n29965 ; n29965_not
g39143 not n19885 ; n19885_not
g39144 not n19759 ; n19759_not
g39145 not n19588 ; n19588_not
g39146 not n18796 ; n18796_not
g39147 not n16978 ; n16978_not
g39148 not n28588 ; n28588_not
g39149 not n16996 ; n16996_not
g39150 not n28678 ; n28678_not
g39151 not n28669 ; n28669_not
g39152 not n18769 ; n18769_not
g39153 not n26887 ; n26887_not
g39154 not n28885 ; n28885_not
g39155 not n29749 ; n29749_not
g39156 not n16888 ; n16888_not
g39157 not n25879 ; n25879_not
g39158 not a[31] ; a[31]_not
g39159 not n24979 ; n24979_not
g39160 not n19777 ; n19777_not
g39161 not n18994 ; n18994_not
g39162 not n29848 ; n29848_not
g39163 not n19498 ; n19498_not
g39164 not n27877 ; n27877_not
g39165 not n19678 ; n19678_not
g39166 not a[22] ; a[22]_not
g39167 not n18976 ; n18976_not
g39168 not n17986 ; n17986_not
g39169 not n19993 ; n19993_not
g39170 not n13999 ; n13999_not
g39171 not n17968 ; n17968_not
g39172 not n26878 ; n26878_not
g39173 not n28984 ; n28984_not
g39174 not n19984 ; n19984_not
g39175 not n29686 ; n29686_not
g39176 not n28498 ; n28498_not
g39177 not n29488 ; n29488_not
g39178 not n17869 ; n17869_not
g39179 not n19696 ; n19696_not
g39180 not n18895 ; n18895_not
g39181 not n18886 ; n18886_not
g39182 not n28948 ; n28948_not
g39183 not n19939 ; n19939_not
g39184 not n26689 ; n26689_not
g39185 not n16789 ; n16789_not
g39186 not n25699 ; n25699_not
g39187 not n18589 ; n18589_not
g39188 not a[14] ; a[14]_not
g39189 not n15989 ; n15989_not
g39190 not a[23] ; a[23]_not
g39191 not n24998 ; n24998_not
g39192 not n27878 ; n27878_not
g39193 not n18779 ; n18779_not
g39194 not n24989 ; n24989_not
g39195 not n25997 ; n25997_not
g39196 not n16898 ; n16898_not
g39197 not n19778 ; n19778_not
g39198 not n17969 ; n17969_not
g39199 not n17996 ; n17996_not
g39200 not n19697 ; n19697_not
g39201 not n29588 ; n29588_not
g39202 not n28769 ; n28769_not
g39203 not n19679 ; n19679_not
g39204 not n19976 ; n19976_not
g39205 not n19994 ; n19994_not
g39206 not n19958 ; n19958_not
g39207 not n16997 ; n16997_not
g39208 not n28958 ; n28958_not
g39209 not n29777 ; n29777_not
g39210 not n16979 ; n16979_not
g39211 not n19886 ; n19886_not
g39212 not n29786 ; n29786_not
g39213 not n29858 ; n29858_not
g39214 not n29876 ; n29876_not
g39215 not n29489 ; n29489_not
g39216 not n29894 ; n29894_not
g39217 not n26897 ; n26897_not
g39218 not n28859 ; n28859_not
g39219 not n28589 ; n28589_not
g39220 not n29957 ; n29957_not
g39221 not n29975 ; n29975_not
g39222 not n19589 ; n19589_not
g39223 not n28949 ; n28949_not
g39224 not n29849 ; n29849_not
g39225 not n25898 ; n25898_not
g39226 not n17888 ; n17888_not
g39227 not n18969 ; n18969_not
g39228 not n29985 ; n29985_not
g39229 not n29994 ; n29994_not
g39230 not n18798 ; n18798_not
g39231 not a[24] ; a[24]_not
g39232 not n29958 ; n29958_not
g39233 not n27699 ; n27699_not
g39234 not n29787 ; n29787_not
g39235 not n29886 ; n29886_not
g39236 not n17979 ; n17979_not
g39237 not n18879 ; n18879_not
g39238 not n17997 ; n17997_not
g39239 not n27978 ; n27978_not
g39240 not a[15] ; a[15]_not
g39241 not n29679 ; n29679_not
g39242 not n26898 ; n26898_not
g39243 not n19896 ; n19896_not
g39244 not n18699 ; n18699_not
g39245 not n28977 ; n28977_not
g39246 not n28869 ; n28869_not
g39247 not n28788 ; n28788_not
g39248 not n28878 ; n28878_not
g39249 not n19968 ; n19968_not
g39250 not n19977 ; n19977_not
g39251 not n28896 ; n28896_not
g39252 not n29598 ; n29598_not
g39253 not a[16] ; a[16]_not
g39254 not a[25] ; a[25]_not
g39255 not n28789 ; n28789_not
g39256 not n29788 ; n29788_not
g39257 not n18889 ; n18889_not
g39258 not n29887 ; n29887_not
g39259 not n29896 ; n29896_not
g39260 not n27997 ; n27997_not
g39261 not n29968 ; n29968_not
g39262 not n28888 ; n28888_not
g39263 not n28897 ; n28897_not
g39264 not n28996 ; n28996_not
g39265 not n29986 ; n29986_not
g39266 not n29689 ; n29689_not
g39267 not n18997 ; n18997_not
g39268 not n29599 ; n29599_not
g39269 not n19987 ; n19987_not
g39270 not n29698 ; n29698_not
g39271 not n28987 ; n28987_not
g39272 not n19798 ; n19798_not
g39273 not n18979 ; n18979_not
g39274 not n25999 ; n25999_not
g39275 not a[26] ; a[26]_not
g39276 not a[17] ; a[17]_not
g39277 not n28889 ; n28889_not
g39278 not n28988 ; n28988_not
g39279 not n19997 ; n19997_not
g39280 not n27998 ; n27998_not
g39281 not a[27] ; a[27]_not
g39282 not a[18] ; a[18]_not
g39283 not n27999 ; n27999_not
g39284 not n19998 ; n19998_not
g39285 not a[19] ; a[19]_not
g39286 not a[28] ; a[28]_not
g39287 not n19999 ; n19999_not
g39288 not a[29] ; a[29]_not
g39289 not n29999 ; n29999_not
