name sqrt
i a[0]
i a[1]
i a[2]
i a[3]
i a[4]
i a[5]
i a[6]
i a[7]
i a[8]
i a[9]
i a[10]
i a[11]
i a[12]
i a[13]
i a[14]
i a[15]
i a[16]
i a[17]
i a[18]
i a[19]
i a[20]
i a[21]
i a[22]
i a[23]
i a[24]
i a[25]
i a[26]
i a[27]
i a[28]
i a[29]
i a[30]
i a[31]
i a[32]
i a[33]
i a[34]
i a[35]
i a[36]
i a[37]
i a[38]
i a[39]
i a[40]
i a[41]
i a[42]
i a[43]
i a[44]
i a[45]
i a[46]
i a[47]
i a[48]
i a[49]
i a[50]
i a[51]
i a[52]
i a[53]
i a[54]
i a[55]
i a[56]
i a[57]
i a[58]
i a[59]
i a[60]
i a[61]
i a[62]
i a[63]
i a[64]
i a[65]
i a[66]
i a[67]
i a[68]
i a[69]
i a[70]
i a[71]
i a[72]
i a[73]
i a[74]
i a[75]
i a[76]
i a[77]
i a[78]
i a[79]
i a[80]
i a[81]
i a[82]
i a[83]
i a[84]
i a[85]
i a[86]
i a[87]
i a[88]
i a[89]
i a[90]
i a[91]
i a[92]
i a[93]
i a[94]
i a[95]
i a[96]
i a[97]
i a[98]
i a[99]
i a[100]
i a[101]
i a[102]
i a[103]
i a[104]
i a[105]
i a[106]
i a[107]
i a[108]
i a[109]
i a[110]
i a[111]
i a[112]
i a[113]
i a[114]
i a[115]
i a[116]
i a[117]
i a[118]
i a[119]
i a[120]
i a[121]
i a[122]
i a[123]
i a[124]
i a[125]
i a[126]
i a[127]

o asqrt[0]
o asqrt[1]
o asqrt[2]
o asqrt[3]
o asqrt[4]
o asqrt[5]
o asqrt[6]
o asqrt[7]
o asqrt[8]
o asqrt[9]
o asqrt[10]
o asqrt[11]
o asqrt[12]
o asqrt[13]
o asqrt[14]
o asqrt[15]
o asqrt[16]
o asqrt[17]
o asqrt[18]
o asqrt[19]
o asqrt[20]
o asqrt[21]
o asqrt[22]
o asqrt[23]
o asqrt[24]
o asqrt[25]
o asqrt[26]
o asqrt[27]
o asqrt[28]
o asqrt[29]
o asqrt[30]
o asqrt[31]
o asqrt[32]
o asqrt[33]
o asqrt[34]
o asqrt[35]
o asqrt[36]
o asqrt[37]
o asqrt[38]
o asqrt[39]
o asqrt[40]
o asqrt[41]
o asqrt[42]
o asqrt[43]
o asqrt[44]
o asqrt[45]
o asqrt[46]
o asqrt[47]
o asqrt[48]
o asqrt[49]
o asqrt[50]
o asqrt[51]
o asqrt[52]
o asqrt[53]
o asqrt[54]
o asqrt[55]
o asqrt[56]
o asqrt[57]
o asqrt[58]
o asqrt[59]
o asqrt[60]
o asqrt[61]
o asqrt[62]
o asqrt[63]

g1 or a[126] a[127] ; asqrt[63]
g2 and a[126] a[127] ; n194
g3 and a[126] asqrt[63] ; n195
g4 nor a[124] a[125] ; n196
g5 nor n195 n196 ; n197
g6 or n194 n197 ; asqrt[62]
g7 and a[124] asqrt[62] ; n199
g8 nor a[122] a[123] ; n200
g9 and a[124]_not n200 ; n201
g10 nor n199 n201 ; n202
g11 and a[124]_not asqrt[62] ; n203
g12 and a[125] n203_not ; n204
g13 and n196 asqrt[62] ; n205
g14 nor n204 n205 ; n206
g15 and n202_not n206 ; n207
g16 nor asqrt[63] n207 ; n208
g17 and n202 n206_not ; n209
g18 and a[126] n196 ; n210
g19 nor a[126] n196 ; n211
g20 and a[127] n211_not ; n212
g21 and n210_not n212 ; n213
g22 nor n209 n213 ; n214
g23 nand n208_not n214 ; asqrt[61]
g24 and a[122] asqrt[61] ; n216
g25 nor a[120] a[121] ; n217
g26 and a[122]_not n217 ; n218
g27 nor n216 n218 ; n219
g28 and asqrt[62] n219_not ; n220
g29 nor n194 n218 ; n221
g30 and n197_not n221 ; n222
g31 and n216_not n222 ; n223
g32 and n200 asqrt[61] ; n224
g33 and a[122]_not asqrt[61] ; n225
g34 and a[123] n225_not ; n226
g35 nor n224 n226 ; n227
g36 and n223_not n227 ; n228
g37 nor n220 n228 ; n229
g38 and asqrt[62] n213_not ; n230
g39 and n209_not n230 ; n231
g40 and n208_not n231 ; n232
g41 nor n224 n232 ; n233
g42 and a[124] n233_not ; n234
g43 nor a[124] n232 ; n235
g44 and n224_not n235 ; n236
g45 nor n234 n236 ; n237
g46 and n207 asqrt[61] ; n238
g47 nor n209 n238 ; n239
g48 and n237_not n239 ; n240
g49 and n229_not n240 ; n241
g50 nor asqrt[63] n241 ; n242
g51 and n229 n237 ; n243
g52 and n206 asqrt[61] ; n244
g53 and n202 n244_not ; n245
g54 and asqrt[63] n207_not ; n246
g55 and n245_not n246 ; n247
g56 nor n206 n213 ; n248
g57 and n209_not n248 ; n249
g58 and n208_not n249 ; n250
g59 nor n247 n250 ; n251
g60 and n243_not n251 ; n252
g61 nand n242_not n252 ; asqrt[60]
g62 and a[120] asqrt[60] ; n254
g63 nor a[118] a[119] ; n255
g64 and a[120]_not n255 ; n256
g65 nor n254 n256 ; n257
g66 and asqrt[61] n257_not ; n258
g67 and a[120]_not asqrt[60] ; n259
g68 and a[121] n259_not ; n260
g69 and n217 asqrt[60] ; n261
g70 nor n260 n261 ; n262
g71 nor n213 n256 ; n263
g72 and n209_not n263 ; n264
g73 and n208_not n264 ; n265
g74 and n254_not n265 ; n266
g75 and n262 n266_not ; n267
g76 nor n258 n267 ; n268
g77 and asqrt[62] n268_not ; n269
g78 nor asqrt[62] n258 ; n270
g79 and n267_not n270 ; n271
g80 and asqrt[61] n250_not ; n272
g81 and n247_not n272 ; n273
g82 and n243_not n273 ; n274
g83 and n242_not n274 ; n275
g84 nor n261 n275 ; n276
g85 and a[122] n276_not ; n277
g86 nor a[122] n275 ; n278
g87 and n261_not n278 ; n279
g88 nor n277 n279 ; n280
g89 nor n271 n280 ; n281
g90 nor n269 n281 ; n282
g91 nor n220 n223 ; n283
g92 and n227_not n283 ; n284
g93 and asqrt[60] n284 ; n285
g94 and asqrt[60] n283 ; n286
g95 and n227 n286_not ; n287
g96 nor n285 n287 ; n288
g97 nor n229 n237 ; n289
g98 and asqrt[60] n289 ; n290
g99 nor n243 n290 ; n291
g100 and n288_not n291 ; n292
g101 and n282_not n292 ; n293
g102 nor asqrt[63] n293 ; n294
g103 and n269_not n288 ; n295
g104 and n281_not n295 ; n296
g105 and n229 asqrt[60] ; n297
g106 nor n237 n297 ; n298
g107 and asqrt[63] n243_not ; n299
g108 and n298_not n299 ; n300
g109 nor n236 n250 ; n301
g110 and n234_not n301 ; n302
g111 and n247_not n302 ; n303
g112 and n243_not n303 ; n304
g113 and n242_not n304 ; n305
g114 nor n300 n305 ; n306
g115 and n296_not n306 ; n307
g116 nand n294_not n307 ; asqrt[59]
g117 and a[118] asqrt[59] ; n309
g118 nor a[116] a[117] ; n310
g119 and a[118]_not n310 ; n311
g120 nor n309 n311 ; n312
g121 and asqrt[60] n312_not ; n313
g122 nor n250 n311 ; n314
g123 and n247_not n314 ; n315
g124 and n243_not n315 ; n316
g125 and n242_not n316 ; n317
g126 and n309_not n317 ; n318
g127 and a[118]_not asqrt[59] ; n319
g128 and a[119] n319_not ; n320
g129 and n255 asqrt[59] ; n321
g130 nor n320 n321 ; n322
g131 and n318_not n322 ; n323
g132 nor n313 n323 ; n324
g133 and asqrt[61] n324_not ; n325
g134 nor asqrt[61] n313 ; n326
g135 and n323_not n326 ; n327
g136 and asqrt[60] n305_not ; n328
g137 and n300_not n328 ; n329
g138 and n296_not n329 ; n330
g139 and n294_not n330 ; n331
g140 nor n321 n331 ; n332
g141 and a[120] n332_not ; n333
g142 nor a[120] n331 ; n334
g143 and n321_not n334 ; n335
g144 nor n333 n335 ; n336
g145 nor n327 n336 ; n337
g146 nor n325 n337 ; n338
g147 and asqrt[62] n338_not ; n339
g148 nor asqrt[62] n325 ; n340
g149 and n337_not n340 ; n341
g150 nor n262 n266 ; n342
g151 and n258_not n342 ; n343
g152 and asqrt[59] n343 ; n344
g153 nor n258 n266 ; n345
g154 and asqrt[59] n345 ; n346
g155 and n262 n346_not ; n347
g156 nor n344 n347 ; n348
g157 nor n341 n348 ; n349
g158 nor n339 n349 ; n350
g159 and n271_not n280 ; n351
g160 and n269_not n351 ; n352
g161 and asqrt[59] n352 ; n353
g162 nor n269 n271 ; n354
g163 and asqrt[59] n354 ; n355
g164 nor n280 n355 ; n356
g165 nor n353 n356 ; n357
g166 nor n282 n288 ; n358
g167 and asqrt[59] n358 ; n359
g168 nor n296 n359 ; n360
g169 and n357_not n360 ; n361
g170 and n350_not n361 ; n362
g171 nor asqrt[63] n362 ; n363
g172 and n339_not n357 ; n364
g173 and n349_not n364 ; n365
g174 and n282 asqrt[59] ; n366
g175 nor n288 n366 ; n367
g176 and asqrt[63] n296_not ; n368
g177 and n367_not n368 ; n369
g178 nor n285 n305 ; n370
g179 and n287_not n370 ; n371
g180 and n300_not n371 ; n372
g181 and n296_not n372 ; n373
g182 and n294_not n373 ; n374
g183 nor n369 n374 ; n375
g184 and n365_not n375 ; n376
g185 nand n363_not n376 ; asqrt[58]
g186 and a[116] asqrt[58] ; n378
g187 nor a[114] a[115] ; n379
g188 and a[116]_not n379 ; n380
g189 nor n378 n380 ; n381
g190 and asqrt[59] n381_not ; n382
g191 nor n305 n380 ; n383
g192 and n300_not n383 ; n384
g193 and n296_not n384 ; n385
g194 and n294_not n385 ; n386
g195 and n378_not n386 ; n387
g196 and a[116]_not asqrt[58] ; n388
g197 and a[117] n388_not ; n389
g198 and n310 asqrt[58] ; n390
g199 nor n389 n390 ; n391
g200 and n387_not n391 ; n392
g201 nor n382 n392 ; n393
g202 and asqrt[60] n393_not ; n394
g203 nor asqrt[60] n382 ; n395
g204 and n392_not n395 ; n396
g205 and asqrt[59] n374_not ; n397
g206 and n369_not n397 ; n398
g207 and n365_not n398 ; n399
g208 and n363_not n399 ; n400
g209 nor n390 n400 ; n401
g210 and a[118] n401_not ; n402
g211 nor a[118] n400 ; n403
g212 and n390_not n403 ; n404
g213 nor n402 n404 ; n405
g214 nor n396 n405 ; n406
g215 nor n394 n406 ; n407
g216 and asqrt[61] n407_not ; n408
g217 nor n313 n318 ; n409
g218 and n322_not n409 ; n410
g219 and asqrt[58] n410 ; n411
g220 and asqrt[58] n409 ; n412
g221 and n322 n412_not ; n413
g222 nor n411 n413 ; n414
g223 nor asqrt[61] n394 ; n415
g224 and n406_not n415 ; n416
g225 nor n414 n416 ; n417
g226 nor n408 n417 ; n418
g227 and asqrt[62] n418_not ; n419
g228 and n327_not n336 ; n420
g229 and n325_not n420 ; n421
g230 and asqrt[58] n421 ; n422
g231 nor n325 n327 ; n423
g232 and asqrt[58] n423 ; n424
g233 nor n336 n424 ; n425
g234 nor n422 n425 ; n426
g235 nor asqrt[62] n408 ; n427
g236 and n417_not n427 ; n428
g237 nor n426 n428 ; n429
g238 nor n419 n429 ; n430
g239 and n339_not n348 ; n431
g240 and n341_not n431 ; n432
g241 and asqrt[58] n432 ; n433
g242 nor n339 n341 ; n434
g243 and asqrt[58] n434 ; n435
g244 nor n348 n435 ; n436
g245 nor n433 n436 ; n437
g246 nor n350 n357 ; n438
g247 and asqrt[58] n438 ; n439
g248 nor n365 n439 ; n440
g249 and n437_not n440 ; n441
g250 and n430_not n441 ; n442
g251 nor asqrt[63] n442 ; n443
g252 and n419_not n437 ; n444
g253 and n429_not n444 ; n445
g254 and n357_not asqrt[58] ; n446
g255 and n350 n446_not ; n447
g256 and asqrt[63] n438_not ; n448
g257 and n447_not n448 ; n449
g258 nor n353 n374 ; n450
g259 and n356_not n450 ; n451
g260 and n369_not n451 ; n452
g261 and n365_not n452 ; n453
g262 and n363_not n453 ; n454
g263 nor n449 n454 ; n455
g264 and n445_not n455 ; n456
g265 nand n443_not n456 ; asqrt[57]
g266 and a[114] asqrt[57] ; n458
g267 nor a[112] a[113] ; n459
g268 and a[114]_not n459 ; n460
g269 nor n458 n460 ; n461
g270 and asqrt[58] n461_not ; n462
g271 nor n374 n460 ; n463
g272 and n369_not n463 ; n464
g273 and n365_not n464 ; n465
g274 and n363_not n465 ; n466
g275 and n458_not n466 ; n467
g276 and a[114]_not asqrt[57] ; n468
g277 and a[115] n468_not ; n469
g278 and n379 asqrt[57] ; n470
g279 nor n469 n470 ; n471
g280 and n467_not n471 ; n472
g281 nor n462 n472 ; n473
g282 and asqrt[59] n473_not ; n474
g283 nor asqrt[59] n462 ; n475
g284 and n472_not n475 ; n476
g285 and asqrt[58] n454_not ; n477
g286 and n449_not n477 ; n478
g287 and n445_not n478 ; n479
g288 and n443_not n479 ; n480
g289 nor n470 n480 ; n481
g290 and a[116] n481_not ; n482
g291 nor a[116] n480 ; n483
g292 and n470_not n483 ; n484
g293 nor n482 n484 ; n485
g294 nor n476 n485 ; n486
g295 nor n474 n486 ; n487
g296 and asqrt[60] n487_not ; n488
g297 nor n382 n387 ; n489
g298 and n391_not n489 ; n490
g299 and asqrt[57] n490 ; n491
g300 and asqrt[57] n489 ; n492
g301 and n391 n492_not ; n493
g302 nor n491 n493 ; n494
g303 nor asqrt[60] n474 ; n495
g304 and n486_not n495 ; n496
g305 nor n494 n496 ; n497
g306 nor n488 n497 ; n498
g307 and asqrt[61] n498_not ; n499
g308 and n396_not n405 ; n500
g309 and n394_not n500 ; n501
g310 and asqrt[57] n501 ; n502
g311 nor n394 n396 ; n503
g312 and asqrt[57] n503 ; n504
g313 nor n405 n504 ; n505
g314 nor n502 n505 ; n506
g315 nor asqrt[61] n488 ; n507
g316 and n497_not n507 ; n508
g317 nor n506 n508 ; n509
g318 nor n499 n509 ; n510
g319 and asqrt[62] n510_not ; n511
g320 and n408_not n414 ; n512
g321 and n416_not n512 ; n513
g322 and asqrt[57] n513 ; n514
g323 nor n408 n416 ; n515
g324 and asqrt[57] n515 ; n516
g325 nor n414 n516 ; n517
g326 nor n514 n517 ; n518
g327 nor asqrt[62] n499 ; n519
g328 and n509_not n519 ; n520
g329 nor n518 n520 ; n521
g330 nor n511 n521 ; n522
g331 and n426 n428_not ; n523
g332 and n419_not n523 ; n524
g333 and asqrt[57] n524 ; n525
g334 nor n419 n428 ; n526
g335 and asqrt[57] n526 ; n527
g336 nor n426 n527 ; n528
g337 nor n525 n528 ; n529
g338 nor n430 n437 ; n530
g339 and asqrt[57] n530 ; n531
g340 nor n445 n531 ; n532
g341 and n529_not n532 ; n533
g342 and n522_not n533 ; n534
g343 nor asqrt[63] n534 ; n535
g344 and n511_not n529 ; n536
g345 and n521_not n536 ; n537
g346 and n437_not asqrt[57] ; n538
g347 and n430 n538_not ; n539
g348 and asqrt[63] n530_not ; n540
g349 and n539_not n540 ; n541
g350 nor n433 n454 ; n542
g351 and n436_not n542 ; n543
g352 and n449_not n543 ; n544
g353 and n445_not n544 ; n545
g354 and n443_not n545 ; n546
g355 nor n541 n546 ; n547
g356 and n537_not n547 ; n548
g357 nand n535_not n548 ; asqrt[56]
g358 and a[112] asqrt[56] ; n550
g359 nor a[110] a[111] ; n551
g360 and a[112]_not n551 ; n552
g361 nor n550 n552 ; n553
g362 and asqrt[57] n553_not ; n554
g363 and a[112]_not asqrt[56] ; n555
g364 and a[113] n555_not ; n556
g365 and n459 asqrt[56] ; n557
g366 nor n556 n557 ; n558
g367 nor n454 n552 ; n559
g368 and n449_not n559 ; n560
g369 and n445_not n560 ; n561
g370 and n443_not n561 ; n562
g371 and n550_not n562 ; n563
g372 and n558 n563_not ; n564
g373 nor n554 n564 ; n565
g374 and asqrt[58] n565_not ; n566
g375 nor asqrt[58] n554 ; n567
g376 and n564_not n567 ; n568
g377 and asqrt[57] n546_not ; n569
g378 and n541_not n569 ; n570
g379 and n537_not n570 ; n571
g380 and n535_not n571 ; n572
g381 nor n557 n572 ; n573
g382 and a[114] n573_not ; n574
g383 nor a[114] n572 ; n575
g384 and n557_not n575 ; n576
g385 nor n574 n576 ; n577
g386 nor n568 n577 ; n578
g387 nor n566 n578 ; n579
g388 and asqrt[59] n579_not ; n580
g389 nor n462 n467 ; n581
g390 and n471_not n581 ; n582
g391 and asqrt[56] n582 ; n583
g392 and asqrt[56] n581 ; n584
g393 and n471 n584_not ; n585
g394 nor n583 n585 ; n586
g395 nor asqrt[59] n566 ; n587
g396 and n578_not n587 ; n588
g397 nor n586 n588 ; n589
g398 nor n580 n589 ; n590
g399 and asqrt[60] n590_not ; n591
g400 and n476_not n485 ; n592
g401 and n474_not n592 ; n593
g402 and asqrt[56] n593 ; n594
g403 nor n474 n476 ; n595
g404 and asqrt[56] n595 ; n596
g405 nor n485 n596 ; n597
g406 nor n594 n597 ; n598
g407 nor asqrt[60] n580 ; n599
g408 and n589_not n599 ; n600
g409 nor n598 n600 ; n601
g410 nor n591 n601 ; n602
g411 and asqrt[61] n602_not ; n603
g412 and n488_not n494 ; n604
g413 and n496_not n604 ; n605
g414 and asqrt[56] n605 ; n606
g415 nor n488 n496 ; n607
g416 and asqrt[56] n607 ; n608
g417 nor n494 n608 ; n609
g418 nor n606 n609 ; n610
g419 nor asqrt[61] n591 ; n611
g420 and n601_not n611 ; n612
g421 nor n610 n612 ; n613
g422 nor n603 n613 ; n614
g423 and asqrt[62] n614_not ; n615
g424 and n506 n508_not ; n616
g425 and n499_not n616 ; n617
g426 and asqrt[56] n617 ; n618
g427 nor n499 n508 ; n619
g428 and asqrt[56] n619 ; n620
g429 nor n506 n620 ; n621
g430 nor n618 n621 ; n622
g431 nor asqrt[62] n603 ; n623
g432 and n613_not n623 ; n624
g433 nor n622 n624 ; n625
g434 nor n615 n625 ; n626
g435 and n511_not n518 ; n627
g436 and n520_not n627 ; n628
g437 and asqrt[56] n628 ; n629
g438 nor n511 n520 ; n630
g439 and asqrt[56] n630 ; n631
g440 nor n518 n631 ; n632
g441 nor n629 n632 ; n633
g442 nor n522 n529 ; n634
g443 and asqrt[56] n634 ; n635
g444 nor n537 n635 ; n636
g445 and n633_not n636 ; n637
g446 and n626_not n637 ; n638
g447 nor asqrt[63] n638 ; n639
g448 and n615_not n633 ; n640
g449 and n625_not n640 ; n641
g450 and n529_not asqrt[56] ; n642
g451 and n522 n642_not ; n643
g452 and asqrt[63] n634_not ; n644
g453 and n643_not n644 ; n645
g454 nor n525 n546 ; n646
g455 and n528_not n646 ; n647
g456 and n541_not n647 ; n648
g457 and n537_not n648 ; n649
g458 and n535_not n649 ; n650
g459 nor n645 n650 ; n651
g460 and n641_not n651 ; n652
g461 nand n639_not n652 ; asqrt[55]
g462 and a[110] asqrt[55] ; n654
g463 nor a[108] a[109] ; n655
g464 and a[110]_not n655 ; n656
g465 nor n654 n656 ; n657
g466 and asqrt[56] n657_not ; n658
g467 nor n546 n656 ; n659
g468 and n541_not n659 ; n660
g469 and n537_not n660 ; n661
g470 and n535_not n661 ; n662
g471 and n654_not n662 ; n663
g472 and a[110]_not asqrt[55] ; n664
g473 and a[111] n664_not ; n665
g474 and n551 asqrt[55] ; n666
g475 nor n665 n666 ; n667
g476 and n663_not n667 ; n668
g477 nor n658 n668 ; n669
g478 and asqrt[57] n669_not ; n670
g479 nor asqrt[57] n658 ; n671
g480 and n668_not n671 ; n672
g481 and asqrt[56] n650_not ; n673
g482 and n645_not n673 ; n674
g483 and n641_not n674 ; n675
g484 and n639_not n675 ; n676
g485 nor n666 n676 ; n677
g486 and a[112] n677_not ; n678
g487 nor a[112] n676 ; n679
g488 and n666_not n679 ; n680
g489 nor n678 n680 ; n681
g490 nor n672 n681 ; n682
g491 nor n670 n682 ; n683
g492 and asqrt[58] n683_not ; n684
g493 nor asqrt[58] n670 ; n685
g494 and n682_not n685 ; n686
g495 nor n558 n563 ; n687
g496 and n554_not n687 ; n688
g497 and asqrt[55] n688 ; n689
g498 nor n554 n563 ; n690
g499 and asqrt[55] n690 ; n691
g500 and n558 n691_not ; n692
g501 nor n689 n692 ; n693
g502 nor n686 n693 ; n694
g503 nor n684 n694 ; n695
g504 and asqrt[59] n695_not ; n696
g505 and n568_not n577 ; n697
g506 and n566_not n697 ; n698
g507 and asqrt[55] n698 ; n699
g508 nor n566 n568 ; n700
g509 and asqrt[55] n700 ; n701
g510 nor n577 n701 ; n702
g511 nor n699 n702 ; n703
g512 nor asqrt[59] n684 ; n704
g513 and n694_not n704 ; n705
g514 nor n703 n705 ; n706
g515 nor n696 n706 ; n707
g516 and asqrt[60] n707_not ; n708
g517 and n580_not n586 ; n709
g518 and n588_not n709 ; n710
g519 and asqrt[55] n710 ; n711
g520 nor n580 n588 ; n712
g521 and asqrt[55] n712 ; n713
g522 nor n586 n713 ; n714
g523 nor n711 n714 ; n715
g524 nor asqrt[60] n696 ; n716
g525 and n706_not n716 ; n717
g526 nor n715 n717 ; n718
g527 nor n708 n718 ; n719
g528 and asqrt[61] n719_not ; n720
g529 and n598 n600_not ; n721
g530 and n591_not n721 ; n722
g531 and asqrt[55] n722 ; n723
g532 nor n591 n600 ; n724
g533 and asqrt[55] n724 ; n725
g534 nor n598 n725 ; n726
g535 nor n723 n726 ; n727
g536 nor asqrt[61] n708 ; n728
g537 and n718_not n728 ; n729
g538 nor n727 n729 ; n730
g539 nor n720 n730 ; n731
g540 and asqrt[62] n731_not ; n732
g541 and n603_not n610 ; n733
g542 and n612_not n733 ; n734
g543 and asqrt[55] n734 ; n735
g544 nor n603 n612 ; n736
g545 and asqrt[55] n736 ; n737
g546 nor n610 n737 ; n738
g547 nor n735 n738 ; n739
g548 nor asqrt[62] n720 ; n740
g549 and n730_not n740 ; n741
g550 nor n739 n741 ; n742
g551 nor n732 n742 ; n743
g552 and n622 n624_not ; n744
g553 and n615_not n744 ; n745
g554 and asqrt[55] n745 ; n746
g555 nor n615 n624 ; n747
g556 and asqrt[55] n747 ; n748
g557 nor n622 n748 ; n749
g558 nor n746 n749 ; n750
g559 nor n626 n633 ; n751
g560 and asqrt[55] n751 ; n752
g561 nor n641 n752 ; n753
g562 and n750_not n753 ; n754
g563 and n743_not n754 ; n755
g564 nor asqrt[63] n755 ; n756
g565 and n732_not n750 ; n757
g566 and n742_not n757 ; n758
g567 and n633_not asqrt[55] ; n759
g568 and n626 n759_not ; n760
g569 and asqrt[63] n751_not ; n761
g570 and n760_not n761 ; n762
g571 nor n629 n650 ; n763
g572 and n632_not n763 ; n764
g573 and n645_not n764 ; n765
g574 and n641_not n765 ; n766
g575 and n639_not n766 ; n767
g576 nor n762 n767 ; n768
g577 and n758_not n768 ; n769
g578 nand n756_not n769 ; asqrt[54]
g579 and a[108] asqrt[54] ; n771
g580 nor a[106] a[107] ; n772
g581 and a[108]_not n772 ; n773
g582 nor n771 n773 ; n774
g583 and asqrt[55] n774_not ; n775
g584 nor n650 n773 ; n776
g585 and n645_not n776 ; n777
g586 and n641_not n777 ; n778
g587 and n639_not n778 ; n779
g588 and n771_not n779 ; n780
g589 and a[108]_not asqrt[54] ; n781
g590 and a[109] n781_not ; n782
g591 and n655 asqrt[54] ; n783
g592 nor n782 n783 ; n784
g593 and n780_not n784 ; n785
g594 nor n775 n785 ; n786
g595 and asqrt[56] n786_not ; n787
g596 nor asqrt[56] n775 ; n788
g597 and n785_not n788 ; n789
g598 and asqrt[55] n767_not ; n790
g599 and n762_not n790 ; n791
g600 and n758_not n791 ; n792
g601 and n756_not n792 ; n793
g602 nor n783 n793 ; n794
g603 and a[110] n794_not ; n795
g604 nor a[110] n793 ; n796
g605 and n783_not n796 ; n797
g606 nor n795 n797 ; n798
g607 nor n789 n798 ; n799
g608 nor n787 n799 ; n800
g609 and asqrt[57] n800_not ; n801
g610 nor n658 n663 ; n802
g611 and n667_not n802 ; n803
g612 and asqrt[54] n803 ; n804
g613 and asqrt[54] n802 ; n805
g614 and n667 n805_not ; n806
g615 nor n804 n806 ; n807
g616 nor asqrt[57] n787 ; n808
g617 and n799_not n808 ; n809
g618 nor n807 n809 ; n810
g619 nor n801 n810 ; n811
g620 and asqrt[58] n811_not ; n812
g621 and n672_not n681 ; n813
g622 and n670_not n813 ; n814
g623 and asqrt[54] n814 ; n815
g624 nor n670 n672 ; n816
g625 and asqrt[54] n816 ; n817
g626 nor n681 n817 ; n818
g627 nor n815 n818 ; n819
g628 nor asqrt[58] n801 ; n820
g629 and n810_not n820 ; n821
g630 nor n819 n821 ; n822
g631 nor n812 n822 ; n823
g632 and asqrt[59] n823_not ; n824
g633 nor asqrt[59] n812 ; n825
g634 and n822_not n825 ; n826
g635 and n684_not n693 ; n827
g636 and n686_not n827 ; n828
g637 and asqrt[54] n828 ; n829
g638 nor n684 n686 ; n830
g639 and asqrt[54] n830 ; n831
g640 nor n693 n831 ; n832
g641 nor n829 n832 ; n833
g642 nor n826 n833 ; n834
g643 nor n824 n834 ; n835
g644 and asqrt[60] n835_not ; n836
g645 and n703 n705_not ; n837
g646 and n696_not n837 ; n838
g647 and asqrt[54] n838 ; n839
g648 nor n696 n705 ; n840
g649 and asqrt[54] n840 ; n841
g650 nor n703 n841 ; n842
g651 nor n839 n842 ; n843
g652 nor asqrt[60] n824 ; n844
g653 and n834_not n844 ; n845
g654 nor n843 n845 ; n846
g655 nor n836 n846 ; n847
g656 and asqrt[61] n847_not ; n848
g657 and n708_not n715 ; n849
g658 and n717_not n849 ; n850
g659 and asqrt[54] n850 ; n851
g660 nor n708 n717 ; n852
g661 and asqrt[54] n852 ; n853
g662 nor n715 n853 ; n854
g663 nor n851 n854 ; n855
g664 nor asqrt[61] n836 ; n856
g665 and n846_not n856 ; n857
g666 nor n855 n857 ; n858
g667 nor n848 n858 ; n859
g668 and asqrt[62] n859_not ; n860
g669 and n727 n729_not ; n861
g670 and n720_not n861 ; n862
g671 and asqrt[54] n862 ; n863
g672 nor n720 n729 ; n864
g673 and asqrt[54] n864 ; n865
g674 nor n727 n865 ; n866
g675 nor n863 n866 ; n867
g676 nor asqrt[62] n848 ; n868
g677 and n858_not n868 ; n869
g678 nor n867 n869 ; n870
g679 nor n860 n870 ; n871
g680 and n732_not n739 ; n872
g681 and n741_not n872 ; n873
g682 and asqrt[54] n873 ; n874
g683 nor n732 n741 ; n875
g684 and asqrt[54] n875 ; n876
g685 nor n739 n876 ; n877
g686 nor n874 n877 ; n878
g687 nor n743 n750 ; n879
g688 and asqrt[54] n879 ; n880
g689 nor n758 n880 ; n881
g690 and n878_not n881 ; n882
g691 and n871_not n882 ; n883
g692 nor asqrt[63] n883 ; n884
g693 and n860_not n878 ; n885
g694 and n870_not n885 ; n886
g695 and n750_not asqrt[54] ; n887
g696 and n743 n887_not ; n888
g697 and asqrt[63] n879_not ; n889
g698 and n888_not n889 ; n890
g699 nor n746 n767 ; n891
g700 and n749_not n891 ; n892
g701 and n762_not n892 ; n893
g702 and n758_not n893 ; n894
g703 and n756_not n894 ; n895
g704 nor n890 n895 ; n896
g705 and n886_not n896 ; n897
g706 nand n884_not n897 ; asqrt[53]
g707 and a[106] asqrt[53] ; n899
g708 nor a[104] a[105] ; n900
g709 and a[106]_not n900 ; n901
g710 nor n899 n901 ; n902
g711 and asqrt[54] n902_not ; n903
g712 nor n767 n901 ; n904
g713 and n762_not n904 ; n905
g714 and n758_not n905 ; n906
g715 and n756_not n906 ; n907
g716 and n899_not n907 ; n908
g717 and a[106]_not asqrt[53] ; n909
g718 and a[107] n909_not ; n910
g719 and n772 asqrt[53] ; n911
g720 nor n910 n911 ; n912
g721 and n908_not n912 ; n913
g722 nor n903 n913 ; n914
g723 and asqrt[55] n914_not ; n915
g724 nor asqrt[55] n903 ; n916
g725 and n913_not n916 ; n917
g726 and asqrt[54] n895_not ; n918
g727 and n890_not n918 ; n919
g728 and n886_not n919 ; n920
g729 and n884_not n920 ; n921
g730 nor n911 n921 ; n922
g731 and a[108] n922_not ; n923
g732 nor a[108] n921 ; n924
g733 and n911_not n924 ; n925
g734 nor n923 n925 ; n926
g735 nor n917 n926 ; n927
g736 nor n915 n927 ; n928
g737 and asqrt[56] n928_not ; n929
g738 nor n775 n780 ; n930
g739 and n784_not n930 ; n931
g740 and asqrt[53] n931 ; n932
g741 and asqrt[53] n930 ; n933
g742 and n784 n933_not ; n934
g743 nor n932 n934 ; n935
g744 nor asqrt[56] n915 ; n936
g745 and n927_not n936 ; n937
g746 nor n935 n937 ; n938
g747 nor n929 n938 ; n939
g748 and asqrt[57] n939_not ; n940
g749 and n789_not n798 ; n941
g750 and n787_not n941 ; n942
g751 and asqrt[53] n942 ; n943
g752 nor n787 n789 ; n944
g753 and asqrt[53] n944 ; n945
g754 nor n798 n945 ; n946
g755 nor n943 n946 ; n947
g756 nor asqrt[57] n929 ; n948
g757 and n938_not n948 ; n949
g758 nor n947 n949 ; n950
g759 nor n940 n950 ; n951
g760 and asqrt[58] n951_not ; n952
g761 and n801_not n807 ; n953
g762 and n809_not n953 ; n954
g763 and asqrt[53] n954 ; n955
g764 nor n801 n809 ; n956
g765 and asqrt[53] n956 ; n957
g766 nor n807 n957 ; n958
g767 nor n955 n958 ; n959
g768 nor asqrt[58] n940 ; n960
g769 and n950_not n960 ; n961
g770 nor n959 n961 ; n962
g771 nor n952 n962 ; n963
g772 and asqrt[59] n963_not ; n964
g773 and n819 n821_not ; n965
g774 and n812_not n965 ; n966
g775 and asqrt[53] n966 ; n967
g776 nor n812 n821 ; n968
g777 and asqrt[53] n968 ; n969
g778 nor n819 n969 ; n970
g779 nor n967 n970 ; n971
g780 nor asqrt[59] n952 ; n972
g781 and n962_not n972 ; n973
g782 nor n971 n973 ; n974
g783 nor n964 n974 ; n975
g784 and asqrt[60] n975_not ; n976
g785 nor asqrt[60] n964 ; n977
g786 and n974_not n977 ; n978
g787 and n824_not n833 ; n979
g788 and n826_not n979 ; n980
g789 and asqrt[53] n980 ; n981
g790 nor n824 n826 ; n982
g791 and asqrt[53] n982 ; n983
g792 nor n833 n983 ; n984
g793 nor n981 n984 ; n985
g794 nor n978 n985 ; n986
g795 nor n976 n986 ; n987
g796 and asqrt[61] n987_not ; n988
g797 and n843 n845_not ; n989
g798 and n836_not n989 ; n990
g799 and asqrt[53] n990 ; n991
g800 nor n836 n845 ; n992
g801 and asqrt[53] n992 ; n993
g802 nor n843 n993 ; n994
g803 nor n991 n994 ; n995
g804 nor asqrt[61] n976 ; n996
g805 and n986_not n996 ; n997
g806 nor n995 n997 ; n998
g807 nor n988 n998 ; n999
g808 and asqrt[62] n999_not ; n1000
g809 and n848_not n855 ; n1001
g810 and n857_not n1001 ; n1002
g811 and asqrt[53] n1002 ; n1003
g812 nor n848 n857 ; n1004
g813 and asqrt[53] n1004 ; n1005
g814 nor n855 n1005 ; n1006
g815 nor n1003 n1006 ; n1007
g816 nor asqrt[62] n988 ; n1008
g817 and n998_not n1008 ; n1009
g818 nor n1007 n1009 ; n1010
g819 nor n1000 n1010 ; n1011
g820 and n867 n869_not ; n1012
g821 and n860_not n1012 ; n1013
g822 and asqrt[53] n1013 ; n1014
g823 nor n860 n869 ; n1015
g824 and asqrt[53] n1015 ; n1016
g825 nor n867 n1016 ; n1017
g826 nor n1014 n1017 ; n1018
g827 nor n871 n878 ; n1019
g828 and asqrt[53] n1019 ; n1020
g829 nor n886 n1020 ; n1021
g830 and n1018_not n1021 ; n1022
g831 and n1011_not n1022 ; n1023
g832 nor asqrt[63] n1023 ; n1024
g833 and n1000_not n1018 ; n1025
g834 and n1010_not n1025 ; n1026
g835 and n878_not asqrt[53] ; n1027
g836 and n871 n1027_not ; n1028
g837 and asqrt[63] n1019_not ; n1029
g838 and n1028_not n1029 ; n1030
g839 nor n874 n895 ; n1031
g840 and n877_not n1031 ; n1032
g841 and n890_not n1032 ; n1033
g842 and n886_not n1033 ; n1034
g843 and n884_not n1034 ; n1035
g844 nor n1030 n1035 ; n1036
g845 and n1026_not n1036 ; n1037
g846 nand n1024_not n1037 ; asqrt[52]
g847 and a[104] asqrt[52] ; n1039
g848 nor a[102] a[103] ; n1040
g849 and a[104]_not n1040 ; n1041
g850 nor n1039 n1041 ; n1042
g851 and asqrt[53] n1042_not ; n1043
g852 nor n895 n1041 ; n1044
g853 and n890_not n1044 ; n1045
g854 and n886_not n1045 ; n1046
g855 and n884_not n1046 ; n1047
g856 and n1039_not n1047 ; n1048
g857 and a[104]_not asqrt[52] ; n1049
g858 and a[105] n1049_not ; n1050
g859 and n900 asqrt[52] ; n1051
g860 nor n1050 n1051 ; n1052
g861 and n1048_not n1052 ; n1053
g862 nor n1043 n1053 ; n1054
g863 and asqrt[54] n1054_not ; n1055
g864 nor asqrt[54] n1043 ; n1056
g865 and n1053_not n1056 ; n1057
g866 and asqrt[53] n1035_not ; n1058
g867 and n1030_not n1058 ; n1059
g868 and n1026_not n1059 ; n1060
g869 and n1024_not n1060 ; n1061
g870 nor n1051 n1061 ; n1062
g871 and a[106] n1062_not ; n1063
g872 nor a[106] n1061 ; n1064
g873 and n1051_not n1064 ; n1065
g874 nor n1063 n1065 ; n1066
g875 nor n1057 n1066 ; n1067
g876 nor n1055 n1067 ; n1068
g877 and asqrt[55] n1068_not ; n1069
g878 nor n903 n908 ; n1070
g879 and n912_not n1070 ; n1071
g880 and asqrt[52] n1071 ; n1072
g881 and asqrt[52] n1070 ; n1073
g882 and n912 n1073_not ; n1074
g883 nor n1072 n1074 ; n1075
g884 nor asqrt[55] n1055 ; n1076
g885 and n1067_not n1076 ; n1077
g886 nor n1075 n1077 ; n1078
g887 nor n1069 n1078 ; n1079
g888 and asqrt[56] n1079_not ; n1080
g889 and n917_not n926 ; n1081
g890 and n915_not n1081 ; n1082
g891 and asqrt[52] n1082 ; n1083
g892 nor n915 n917 ; n1084
g893 and asqrt[52] n1084 ; n1085
g894 nor n926 n1085 ; n1086
g895 nor n1083 n1086 ; n1087
g896 nor asqrt[56] n1069 ; n1088
g897 and n1078_not n1088 ; n1089
g898 nor n1087 n1089 ; n1090
g899 nor n1080 n1090 ; n1091
g900 and asqrt[57] n1091_not ; n1092
g901 and n929_not n935 ; n1093
g902 and n937_not n1093 ; n1094
g903 and asqrt[52] n1094 ; n1095
g904 nor n929 n937 ; n1096
g905 and asqrt[52] n1096 ; n1097
g906 nor n935 n1097 ; n1098
g907 nor n1095 n1098 ; n1099
g908 nor asqrt[57] n1080 ; n1100
g909 and n1090_not n1100 ; n1101
g910 nor n1099 n1101 ; n1102
g911 nor n1092 n1102 ; n1103
g912 and asqrt[58] n1103_not ; n1104
g913 and n947 n949_not ; n1105
g914 and n940_not n1105 ; n1106
g915 and asqrt[52] n1106 ; n1107
g916 nor n940 n949 ; n1108
g917 and asqrt[52] n1108 ; n1109
g918 nor n947 n1109 ; n1110
g919 nor n1107 n1110 ; n1111
g920 nor asqrt[58] n1092 ; n1112
g921 and n1102_not n1112 ; n1113
g922 nor n1111 n1113 ; n1114
g923 nor n1104 n1114 ; n1115
g924 and asqrt[59] n1115_not ; n1116
g925 and n952_not n959 ; n1117
g926 and n961_not n1117 ; n1118
g927 and asqrt[52] n1118 ; n1119
g928 nor n952 n961 ; n1120
g929 and asqrt[52] n1120 ; n1121
g930 nor n959 n1121 ; n1122
g931 nor n1119 n1122 ; n1123
g932 nor asqrt[59] n1104 ; n1124
g933 and n1114_not n1124 ; n1125
g934 nor n1123 n1125 ; n1126
g935 nor n1116 n1126 ; n1127
g936 and asqrt[60] n1127_not ; n1128
g937 and n971 n973_not ; n1129
g938 and n964_not n1129 ; n1130
g939 and asqrt[52] n1130 ; n1131
g940 nor n964 n973 ; n1132
g941 and asqrt[52] n1132 ; n1133
g942 nor n971 n1133 ; n1134
g943 nor n1131 n1134 ; n1135
g944 nor asqrt[60] n1116 ; n1136
g945 and n1126_not n1136 ; n1137
g946 nor n1135 n1137 ; n1138
g947 nor n1128 n1138 ; n1139
g948 and asqrt[61] n1139_not ; n1140
g949 nor asqrt[61] n1128 ; n1141
g950 and n1138_not n1141 ; n1142
g951 and n976_not n985 ; n1143
g952 and n978_not n1143 ; n1144
g953 and asqrt[52] n1144 ; n1145
g954 nor n976 n978 ; n1146
g955 and asqrt[52] n1146 ; n1147
g956 nor n985 n1147 ; n1148
g957 nor n1145 n1148 ; n1149
g958 nor n1142 n1149 ; n1150
g959 nor n1140 n1150 ; n1151
g960 and asqrt[62] n1151_not ; n1152
g961 and n995 n997_not ; n1153
g962 and n988_not n1153 ; n1154
g963 and asqrt[52] n1154 ; n1155
g964 nor n988 n997 ; n1156
g965 and asqrt[52] n1156 ; n1157
g966 nor n995 n1157 ; n1158
g967 nor n1155 n1158 ; n1159
g968 nor asqrt[62] n1140 ; n1160
g969 and n1150_not n1160 ; n1161
g970 nor n1159 n1161 ; n1162
g971 nor n1152 n1162 ; n1163
g972 and n1000_not n1007 ; n1164
g973 and n1009_not n1164 ; n1165
g974 and asqrt[52] n1165 ; n1166
g975 nor n1000 n1009 ; n1167
g976 and asqrt[52] n1167 ; n1168
g977 nor n1007 n1168 ; n1169
g978 nor n1166 n1169 ; n1170
g979 nor n1011 n1018 ; n1171
g980 and asqrt[52] n1171 ; n1172
g981 nor n1026 n1172 ; n1173
g982 and n1170_not n1173 ; n1174
g983 and n1163_not n1174 ; n1175
g984 nor asqrt[63] n1175 ; n1176
g985 and n1152_not n1170 ; n1177
g986 and n1162_not n1177 ; n1178
g987 and n1018_not asqrt[52] ; n1179
g988 and n1011 n1179_not ; n1180
g989 and asqrt[63] n1171_not ; n1181
g990 and n1180_not n1181 ; n1182
g991 nor n1014 n1035 ; n1183
g992 and n1017_not n1183 ; n1184
g993 and n1030_not n1184 ; n1185
g994 and n1026_not n1185 ; n1186
g995 and n1024_not n1186 ; n1187
g996 nor n1182 n1187 ; n1188
g997 and n1178_not n1188 ; n1189
g998 nand n1176_not n1189 ; asqrt[51]
g999 and a[102] asqrt[51] ; n1191
g1000 nor a[100] a[101] ; n1192
g1001 and a[102]_not n1192 ; n1193
g1002 nor n1191 n1193 ; n1194
g1003 and asqrt[52] n1194_not ; n1195
g1004 nor n1035 n1193 ; n1196
g1005 and n1030_not n1196 ; n1197
g1006 and n1026_not n1197 ; n1198
g1007 and n1024_not n1198 ; n1199
g1008 and n1191_not n1199 ; n1200
g1009 and a[102]_not asqrt[51] ; n1201
g1010 and a[103] n1201_not ; n1202
g1011 and n1040 asqrt[51] ; n1203
g1012 nor n1202 n1203 ; n1204
g1013 and n1200_not n1204 ; n1205
g1014 nor n1195 n1205 ; n1206
g1015 and asqrt[53] n1206_not ; n1207
g1016 nor asqrt[53] n1195 ; n1208
g1017 and n1205_not n1208 ; n1209
g1018 and asqrt[52] n1187_not ; n1210
g1019 and n1182_not n1210 ; n1211
g1020 and n1178_not n1211 ; n1212
g1021 and n1176_not n1212 ; n1213
g1022 nor n1203 n1213 ; n1214
g1023 and a[104] n1214_not ; n1215
g1024 nor a[104] n1213 ; n1216
g1025 and n1203_not n1216 ; n1217
g1026 nor n1215 n1217 ; n1218
g1027 nor n1209 n1218 ; n1219
g1028 nor n1207 n1219 ; n1220
g1029 and asqrt[54] n1220_not ; n1221
g1030 nor n1043 n1048 ; n1222
g1031 and n1052_not n1222 ; n1223
g1032 and asqrt[51] n1223 ; n1224
g1033 and asqrt[51] n1222 ; n1225
g1034 and n1052 n1225_not ; n1226
g1035 nor n1224 n1226 ; n1227
g1036 nor asqrt[54] n1207 ; n1228
g1037 and n1219_not n1228 ; n1229
g1038 nor n1227 n1229 ; n1230
g1039 nor n1221 n1230 ; n1231
g1040 and asqrt[55] n1231_not ; n1232
g1041 and n1057_not n1066 ; n1233
g1042 and n1055_not n1233 ; n1234
g1043 and asqrt[51] n1234 ; n1235
g1044 nor n1055 n1057 ; n1236
g1045 and asqrt[51] n1236 ; n1237
g1046 nor n1066 n1237 ; n1238
g1047 nor n1235 n1238 ; n1239
g1048 nor asqrt[55] n1221 ; n1240
g1049 and n1230_not n1240 ; n1241
g1050 nor n1239 n1241 ; n1242
g1051 nor n1232 n1242 ; n1243
g1052 and asqrt[56] n1243_not ; n1244
g1053 and n1069_not n1075 ; n1245
g1054 and n1077_not n1245 ; n1246
g1055 and asqrt[51] n1246 ; n1247
g1056 nor n1069 n1077 ; n1248
g1057 and asqrt[51] n1248 ; n1249
g1058 nor n1075 n1249 ; n1250
g1059 nor n1247 n1250 ; n1251
g1060 nor asqrt[56] n1232 ; n1252
g1061 and n1242_not n1252 ; n1253
g1062 nor n1251 n1253 ; n1254
g1063 nor n1244 n1254 ; n1255
g1064 and asqrt[57] n1255_not ; n1256
g1065 and n1087 n1089_not ; n1257
g1066 and n1080_not n1257 ; n1258
g1067 and asqrt[51] n1258 ; n1259
g1068 nor n1080 n1089 ; n1260
g1069 and asqrt[51] n1260 ; n1261
g1070 nor n1087 n1261 ; n1262
g1071 nor n1259 n1262 ; n1263
g1072 nor asqrt[57] n1244 ; n1264
g1073 and n1254_not n1264 ; n1265
g1074 nor n1263 n1265 ; n1266
g1075 nor n1256 n1266 ; n1267
g1076 and asqrt[58] n1267_not ; n1268
g1077 and n1092_not n1099 ; n1269
g1078 and n1101_not n1269 ; n1270
g1079 and asqrt[51] n1270 ; n1271
g1080 nor n1092 n1101 ; n1272
g1081 and asqrt[51] n1272 ; n1273
g1082 nor n1099 n1273 ; n1274
g1083 nor n1271 n1274 ; n1275
g1084 nor asqrt[58] n1256 ; n1276
g1085 and n1266_not n1276 ; n1277
g1086 nor n1275 n1277 ; n1278
g1087 nor n1268 n1278 ; n1279
g1088 and asqrt[59] n1279_not ; n1280
g1089 and n1111 n1113_not ; n1281
g1090 and n1104_not n1281 ; n1282
g1091 and asqrt[51] n1282 ; n1283
g1092 nor n1104 n1113 ; n1284
g1093 and asqrt[51] n1284 ; n1285
g1094 nor n1111 n1285 ; n1286
g1095 nor n1283 n1286 ; n1287
g1096 nor asqrt[59] n1268 ; n1288
g1097 and n1278_not n1288 ; n1289
g1098 nor n1287 n1289 ; n1290
g1099 nor n1280 n1290 ; n1291
g1100 and asqrt[60] n1291_not ; n1292
g1101 and n1116_not n1123 ; n1293
g1102 and n1125_not n1293 ; n1294
g1103 and asqrt[51] n1294 ; n1295
g1104 nor n1116 n1125 ; n1296
g1105 and asqrt[51] n1296 ; n1297
g1106 nor n1123 n1297 ; n1298
g1107 nor n1295 n1298 ; n1299
g1108 nor asqrt[60] n1280 ; n1300
g1109 and n1290_not n1300 ; n1301
g1110 nor n1299 n1301 ; n1302
g1111 nor n1292 n1302 ; n1303
g1112 and asqrt[61] n1303_not ; n1304
g1113 and n1135 n1137_not ; n1305
g1114 and n1128_not n1305 ; n1306
g1115 and asqrt[51] n1306 ; n1307
g1116 nor n1128 n1137 ; n1308
g1117 and asqrt[51] n1308 ; n1309
g1118 nor n1135 n1309 ; n1310
g1119 nor n1307 n1310 ; n1311
g1120 nor asqrt[61] n1292 ; n1312
g1121 and n1302_not n1312 ; n1313
g1122 nor n1311 n1313 ; n1314
g1123 nor n1304 n1314 ; n1315
g1124 and asqrt[62] n1315_not ; n1316
g1125 nor asqrt[62] n1304 ; n1317
g1126 and n1314_not n1317 ; n1318
g1127 and n1140_not n1149 ; n1319
g1128 and n1142_not n1319 ; n1320
g1129 and asqrt[51] n1320 ; n1321
g1130 nor n1140 n1142 ; n1322
g1131 and asqrt[51] n1322 ; n1323
g1132 nor n1149 n1323 ; n1324
g1133 nor n1321 n1324 ; n1325
g1134 nor n1318 n1325 ; n1326
g1135 nor n1316 n1326 ; n1327
g1136 and n1159 n1161_not ; n1328
g1137 and n1152_not n1328 ; n1329
g1138 and asqrt[51] n1329 ; n1330
g1139 nor n1152 n1161 ; n1331
g1140 and asqrt[51] n1331 ; n1332
g1141 nor n1159 n1332 ; n1333
g1142 nor n1330 n1333 ; n1334
g1143 nor n1163 n1170 ; n1335
g1144 and asqrt[51] n1335 ; n1336
g1145 nor n1178 n1336 ; n1337
g1146 and n1334_not n1337 ; n1338
g1147 and n1327_not n1338 ; n1339
g1148 nor asqrt[63] n1339 ; n1340
g1149 and n1316_not n1334 ; n1341
g1150 and n1326_not n1341 ; n1342
g1151 and n1170_not asqrt[51] ; n1343
g1152 and n1163 n1343_not ; n1344
g1153 and asqrt[63] n1335_not ; n1345
g1154 and n1344_not n1345 ; n1346
g1155 nor n1166 n1187 ; n1347
g1156 and n1169_not n1347 ; n1348
g1157 and n1182_not n1348 ; n1349
g1158 and n1178_not n1349 ; n1350
g1159 and n1176_not n1350 ; n1351
g1160 nor n1346 n1351 ; n1352
g1161 and n1342_not n1352 ; n1353
g1162 nand n1340_not n1353 ; asqrt[50]
g1163 and a[100] asqrt[50] ; n1355
g1164 nor a[98] a[99] ; n1356
g1165 and a[100]_not n1356 ; n1357
g1166 nor n1355 n1357 ; n1358
g1167 and asqrt[51] n1358_not ; n1359
g1168 nor n1187 n1357 ; n1360
g1169 and n1182_not n1360 ; n1361
g1170 and n1178_not n1361 ; n1362
g1171 and n1176_not n1362 ; n1363
g1172 and n1355_not n1363 ; n1364
g1173 and a[100]_not asqrt[50] ; n1365
g1174 and a[101] n1365_not ; n1366
g1175 and n1192 asqrt[50] ; n1367
g1176 nor n1366 n1367 ; n1368
g1177 and n1364_not n1368 ; n1369
g1178 nor n1359 n1369 ; n1370
g1179 and asqrt[52] n1370_not ; n1371
g1180 nor asqrt[52] n1359 ; n1372
g1181 and n1369_not n1372 ; n1373
g1182 and asqrt[51] n1351_not ; n1374
g1183 and n1346_not n1374 ; n1375
g1184 and n1342_not n1375 ; n1376
g1185 and n1340_not n1376 ; n1377
g1186 nor n1367 n1377 ; n1378
g1187 and a[102] n1378_not ; n1379
g1188 nor a[102] n1377 ; n1380
g1189 and n1367_not n1380 ; n1381
g1190 nor n1379 n1381 ; n1382
g1191 nor n1373 n1382 ; n1383
g1192 nor n1371 n1383 ; n1384
g1193 and asqrt[53] n1384_not ; n1385
g1194 nor n1195 n1200 ; n1386
g1195 and n1204_not n1386 ; n1387
g1196 and asqrt[50] n1387 ; n1388
g1197 and asqrt[50] n1386 ; n1389
g1198 and n1204 n1389_not ; n1390
g1199 nor n1388 n1390 ; n1391
g1200 nor asqrt[53] n1371 ; n1392
g1201 and n1383_not n1392 ; n1393
g1202 nor n1391 n1393 ; n1394
g1203 nor n1385 n1394 ; n1395
g1204 and asqrt[54] n1395_not ; n1396
g1205 and n1209_not n1218 ; n1397
g1206 and n1207_not n1397 ; n1398
g1207 and asqrt[50] n1398 ; n1399
g1208 nor n1207 n1209 ; n1400
g1209 and asqrt[50] n1400 ; n1401
g1210 nor n1218 n1401 ; n1402
g1211 nor n1399 n1402 ; n1403
g1212 nor asqrt[54] n1385 ; n1404
g1213 and n1394_not n1404 ; n1405
g1214 nor n1403 n1405 ; n1406
g1215 nor n1396 n1406 ; n1407
g1216 and asqrt[55] n1407_not ; n1408
g1217 and n1221_not n1227 ; n1409
g1218 and n1229_not n1409 ; n1410
g1219 and asqrt[50] n1410 ; n1411
g1220 nor n1221 n1229 ; n1412
g1221 and asqrt[50] n1412 ; n1413
g1222 nor n1227 n1413 ; n1414
g1223 nor n1411 n1414 ; n1415
g1224 nor asqrt[55] n1396 ; n1416
g1225 and n1406_not n1416 ; n1417
g1226 nor n1415 n1417 ; n1418
g1227 nor n1408 n1418 ; n1419
g1228 and asqrt[56] n1419_not ; n1420
g1229 and n1239 n1241_not ; n1421
g1230 and n1232_not n1421 ; n1422
g1231 and asqrt[50] n1422 ; n1423
g1232 nor n1232 n1241 ; n1424
g1233 and asqrt[50] n1424 ; n1425
g1234 nor n1239 n1425 ; n1426
g1235 nor n1423 n1426 ; n1427
g1236 nor asqrt[56] n1408 ; n1428
g1237 and n1418_not n1428 ; n1429
g1238 nor n1427 n1429 ; n1430
g1239 nor n1420 n1430 ; n1431
g1240 and asqrt[57] n1431_not ; n1432
g1241 and n1244_not n1251 ; n1433
g1242 and n1253_not n1433 ; n1434
g1243 and asqrt[50] n1434 ; n1435
g1244 nor n1244 n1253 ; n1436
g1245 and asqrt[50] n1436 ; n1437
g1246 nor n1251 n1437 ; n1438
g1247 nor n1435 n1438 ; n1439
g1248 nor asqrt[57] n1420 ; n1440
g1249 and n1430_not n1440 ; n1441
g1250 nor n1439 n1441 ; n1442
g1251 nor n1432 n1442 ; n1443
g1252 and asqrt[58] n1443_not ; n1444
g1253 and n1263 n1265_not ; n1445
g1254 and n1256_not n1445 ; n1446
g1255 and asqrt[50] n1446 ; n1447
g1256 nor n1256 n1265 ; n1448
g1257 and asqrt[50] n1448 ; n1449
g1258 nor n1263 n1449 ; n1450
g1259 nor n1447 n1450 ; n1451
g1260 nor asqrt[58] n1432 ; n1452
g1261 and n1442_not n1452 ; n1453
g1262 nor n1451 n1453 ; n1454
g1263 nor n1444 n1454 ; n1455
g1264 and asqrt[59] n1455_not ; n1456
g1265 and n1268_not n1275 ; n1457
g1266 and n1277_not n1457 ; n1458
g1267 and asqrt[50] n1458 ; n1459
g1268 nor n1268 n1277 ; n1460
g1269 and asqrt[50] n1460 ; n1461
g1270 nor n1275 n1461 ; n1462
g1271 nor n1459 n1462 ; n1463
g1272 nor asqrt[59] n1444 ; n1464
g1273 and n1454_not n1464 ; n1465
g1274 nor n1463 n1465 ; n1466
g1275 nor n1456 n1466 ; n1467
g1276 and asqrt[60] n1467_not ; n1468
g1277 and n1287 n1289_not ; n1469
g1278 and n1280_not n1469 ; n1470
g1279 and asqrt[50] n1470 ; n1471
g1280 nor n1280 n1289 ; n1472
g1281 and asqrt[50] n1472 ; n1473
g1282 nor n1287 n1473 ; n1474
g1283 nor n1471 n1474 ; n1475
g1284 nor asqrt[60] n1456 ; n1476
g1285 and n1466_not n1476 ; n1477
g1286 nor n1475 n1477 ; n1478
g1287 nor n1468 n1478 ; n1479
g1288 and asqrt[61] n1479_not ; n1480
g1289 and n1292_not n1299 ; n1481
g1290 and n1301_not n1481 ; n1482
g1291 and asqrt[50] n1482 ; n1483
g1292 nor n1292 n1301 ; n1484
g1293 and asqrt[50] n1484 ; n1485
g1294 nor n1299 n1485 ; n1486
g1295 nor n1483 n1486 ; n1487
g1296 nor asqrt[61] n1468 ; n1488
g1297 and n1478_not n1488 ; n1489
g1298 nor n1487 n1489 ; n1490
g1299 nor n1480 n1490 ; n1491
g1300 and asqrt[62] n1491_not ; n1492
g1301 and n1311 n1313_not ; n1493
g1302 and n1304_not n1493 ; n1494
g1303 and asqrt[50] n1494 ; n1495
g1304 nor n1304 n1313 ; n1496
g1305 and asqrt[50] n1496 ; n1497
g1306 nor n1311 n1497 ; n1498
g1307 nor n1495 n1498 ; n1499
g1308 nor asqrt[62] n1480 ; n1500
g1309 and n1490_not n1500 ; n1501
g1310 nor n1499 n1501 ; n1502
g1311 nor n1492 n1502 ; n1503
g1312 and n1316_not n1325 ; n1504
g1313 and n1318_not n1504 ; n1505
g1314 and asqrt[50] n1505 ; n1506
g1315 nor n1316 n1318 ; n1507
g1316 and asqrt[50] n1507 ; n1508
g1317 nor n1325 n1508 ; n1509
g1318 nor n1506 n1509 ; n1510
g1319 nor n1327 n1334 ; n1511
g1320 and asqrt[50] n1511 ; n1512
g1321 nor n1342 n1512 ; n1513
g1322 and n1510_not n1513 ; n1514
g1323 and n1503_not n1514 ; n1515
g1324 nor asqrt[63] n1515 ; n1516
g1325 and n1492_not n1510 ; n1517
g1326 and n1502_not n1517 ; n1518
g1327 and n1334_not asqrt[50] ; n1519
g1328 and n1327 n1519_not ; n1520
g1329 and asqrt[63] n1511_not ; n1521
g1330 and n1520_not n1521 ; n1522
g1331 nor n1330 n1351 ; n1523
g1332 and n1333_not n1523 ; n1524
g1333 and n1346_not n1524 ; n1525
g1334 and n1342_not n1525 ; n1526
g1335 and n1340_not n1526 ; n1527
g1336 nor n1522 n1527 ; n1528
g1337 and n1518_not n1528 ; n1529
g1338 nand n1516_not n1529 ; asqrt[49]
g1339 and a[98] asqrt[49] ; n1531
g1340 nor a[96] a[97] ; n1532
g1341 and a[98]_not n1532 ; n1533
g1342 nor n1531 n1533 ; n1534
g1343 and asqrt[50] n1534_not ; n1535
g1344 nor n1351 n1533 ; n1536
g1345 and n1346_not n1536 ; n1537
g1346 and n1342_not n1537 ; n1538
g1347 and n1340_not n1538 ; n1539
g1348 and n1531_not n1539 ; n1540
g1349 and a[98]_not asqrt[49] ; n1541
g1350 and a[99] n1541_not ; n1542
g1351 and n1356 asqrt[49] ; n1543
g1352 nor n1542 n1543 ; n1544
g1353 and n1540_not n1544 ; n1545
g1354 nor n1535 n1545 ; n1546
g1355 and asqrt[51] n1546_not ; n1547
g1356 nor asqrt[51] n1535 ; n1548
g1357 and n1545_not n1548 ; n1549
g1358 and asqrt[50] n1527_not ; n1550
g1359 and n1522_not n1550 ; n1551
g1360 and n1518_not n1551 ; n1552
g1361 and n1516_not n1552 ; n1553
g1362 nor n1543 n1553 ; n1554
g1363 and a[100] n1554_not ; n1555
g1364 nor a[100] n1553 ; n1556
g1365 and n1543_not n1556 ; n1557
g1366 nor n1555 n1557 ; n1558
g1367 nor n1549 n1558 ; n1559
g1368 nor n1547 n1559 ; n1560
g1369 and asqrt[52] n1560_not ; n1561
g1370 nor n1359 n1364 ; n1562
g1371 and n1368_not n1562 ; n1563
g1372 and asqrt[49] n1563 ; n1564
g1373 and asqrt[49] n1562 ; n1565
g1374 and n1368 n1565_not ; n1566
g1375 nor n1564 n1566 ; n1567
g1376 nor asqrt[52] n1547 ; n1568
g1377 and n1559_not n1568 ; n1569
g1378 nor n1567 n1569 ; n1570
g1379 nor n1561 n1570 ; n1571
g1380 and asqrt[53] n1571_not ; n1572
g1381 and n1373_not n1382 ; n1573
g1382 and n1371_not n1573 ; n1574
g1383 and asqrt[49] n1574 ; n1575
g1384 nor n1371 n1373 ; n1576
g1385 and asqrt[49] n1576 ; n1577
g1386 nor n1382 n1577 ; n1578
g1387 nor n1575 n1578 ; n1579
g1388 nor asqrt[53] n1561 ; n1580
g1389 and n1570_not n1580 ; n1581
g1390 nor n1579 n1581 ; n1582
g1391 nor n1572 n1582 ; n1583
g1392 and asqrt[54] n1583_not ; n1584
g1393 and n1385_not n1391 ; n1585
g1394 and n1393_not n1585 ; n1586
g1395 and asqrt[49] n1586 ; n1587
g1396 nor n1385 n1393 ; n1588
g1397 and asqrt[49] n1588 ; n1589
g1398 nor n1391 n1589 ; n1590
g1399 nor n1587 n1590 ; n1591
g1400 nor asqrt[54] n1572 ; n1592
g1401 and n1582_not n1592 ; n1593
g1402 nor n1591 n1593 ; n1594
g1403 nor n1584 n1594 ; n1595
g1404 and asqrt[55] n1595_not ; n1596
g1405 and n1403 n1405_not ; n1597
g1406 and n1396_not n1597 ; n1598
g1407 and asqrt[49] n1598 ; n1599
g1408 nor n1396 n1405 ; n1600
g1409 and asqrt[49] n1600 ; n1601
g1410 nor n1403 n1601 ; n1602
g1411 nor n1599 n1602 ; n1603
g1412 nor asqrt[55] n1584 ; n1604
g1413 and n1594_not n1604 ; n1605
g1414 nor n1603 n1605 ; n1606
g1415 nor n1596 n1606 ; n1607
g1416 and asqrt[56] n1607_not ; n1608
g1417 and n1408_not n1415 ; n1609
g1418 and n1417_not n1609 ; n1610
g1419 and asqrt[49] n1610 ; n1611
g1420 nor n1408 n1417 ; n1612
g1421 and asqrt[49] n1612 ; n1613
g1422 nor n1415 n1613 ; n1614
g1423 nor n1611 n1614 ; n1615
g1424 nor asqrt[56] n1596 ; n1616
g1425 and n1606_not n1616 ; n1617
g1426 nor n1615 n1617 ; n1618
g1427 nor n1608 n1618 ; n1619
g1428 and asqrt[57] n1619_not ; n1620
g1429 and n1427 n1429_not ; n1621
g1430 and n1420_not n1621 ; n1622
g1431 and asqrt[49] n1622 ; n1623
g1432 nor n1420 n1429 ; n1624
g1433 and asqrt[49] n1624 ; n1625
g1434 nor n1427 n1625 ; n1626
g1435 nor n1623 n1626 ; n1627
g1436 nor asqrt[57] n1608 ; n1628
g1437 and n1618_not n1628 ; n1629
g1438 nor n1627 n1629 ; n1630
g1439 nor n1620 n1630 ; n1631
g1440 and asqrt[58] n1631_not ; n1632
g1441 and n1432_not n1439 ; n1633
g1442 and n1441_not n1633 ; n1634
g1443 and asqrt[49] n1634 ; n1635
g1444 nor n1432 n1441 ; n1636
g1445 and asqrt[49] n1636 ; n1637
g1446 nor n1439 n1637 ; n1638
g1447 nor n1635 n1638 ; n1639
g1448 nor asqrt[58] n1620 ; n1640
g1449 and n1630_not n1640 ; n1641
g1450 nor n1639 n1641 ; n1642
g1451 nor n1632 n1642 ; n1643
g1452 and asqrt[59] n1643_not ; n1644
g1453 and n1451 n1453_not ; n1645
g1454 and n1444_not n1645 ; n1646
g1455 and asqrt[49] n1646 ; n1647
g1456 nor n1444 n1453 ; n1648
g1457 and asqrt[49] n1648 ; n1649
g1458 nor n1451 n1649 ; n1650
g1459 nor n1647 n1650 ; n1651
g1460 nor asqrt[59] n1632 ; n1652
g1461 and n1642_not n1652 ; n1653
g1462 nor n1651 n1653 ; n1654
g1463 nor n1644 n1654 ; n1655
g1464 and asqrt[60] n1655_not ; n1656
g1465 and n1456_not n1463 ; n1657
g1466 and n1465_not n1657 ; n1658
g1467 and asqrt[49] n1658 ; n1659
g1468 nor n1456 n1465 ; n1660
g1469 and asqrt[49] n1660 ; n1661
g1470 nor n1463 n1661 ; n1662
g1471 nor n1659 n1662 ; n1663
g1472 nor asqrt[60] n1644 ; n1664
g1473 and n1654_not n1664 ; n1665
g1474 nor n1663 n1665 ; n1666
g1475 nor n1656 n1666 ; n1667
g1476 and asqrt[61] n1667_not ; n1668
g1477 and n1475 n1477_not ; n1669
g1478 and n1468_not n1669 ; n1670
g1479 and asqrt[49] n1670 ; n1671
g1480 nor n1468 n1477 ; n1672
g1481 and asqrt[49] n1672 ; n1673
g1482 nor n1475 n1673 ; n1674
g1483 nor n1671 n1674 ; n1675
g1484 nor asqrt[61] n1656 ; n1676
g1485 and n1666_not n1676 ; n1677
g1486 nor n1675 n1677 ; n1678
g1487 nor n1668 n1678 ; n1679
g1488 and asqrt[62] n1679_not ; n1680
g1489 and n1480_not n1487 ; n1681
g1490 and n1489_not n1681 ; n1682
g1491 and asqrt[49] n1682 ; n1683
g1492 nor n1480 n1489 ; n1684
g1493 and asqrt[49] n1684 ; n1685
g1494 nor n1487 n1685 ; n1686
g1495 nor n1683 n1686 ; n1687
g1496 nor asqrt[62] n1668 ; n1688
g1497 and n1678_not n1688 ; n1689
g1498 nor n1687 n1689 ; n1690
g1499 nor n1680 n1690 ; n1691
g1500 and n1499 n1501_not ; n1692
g1501 and n1492_not n1692 ; n1693
g1502 and asqrt[49] n1693 ; n1694
g1503 nor n1492 n1501 ; n1695
g1504 and asqrt[49] n1695 ; n1696
g1505 nor n1499 n1696 ; n1697
g1506 nor n1694 n1697 ; n1698
g1507 nor n1503 n1510 ; n1699
g1508 and asqrt[49] n1699 ; n1700
g1509 nor n1518 n1700 ; n1701
g1510 and n1698_not n1701 ; n1702
g1511 and n1691_not n1702 ; n1703
g1512 nor asqrt[63] n1703 ; n1704
g1513 and n1680_not n1698 ; n1705
g1514 and n1690_not n1705 ; n1706
g1515 and n1510_not asqrt[49] ; n1707
g1516 and n1503 n1707_not ; n1708
g1517 and asqrt[63] n1699_not ; n1709
g1518 and n1708_not n1709 ; n1710
g1519 nor n1506 n1527 ; n1711
g1520 and n1509_not n1711 ; n1712
g1521 and n1522_not n1712 ; n1713
g1522 and n1518_not n1713 ; n1714
g1523 and n1516_not n1714 ; n1715
g1524 nor n1710 n1715 ; n1716
g1525 and n1706_not n1716 ; n1717
g1526 nand n1704_not n1717 ; asqrt[48]
g1527 and a[96] asqrt[48] ; n1719
g1528 nor a[94] a[95] ; n1720
g1529 and a[96]_not n1720 ; n1721
g1530 nor n1719 n1721 ; n1722
g1531 and asqrt[49] n1722_not ; n1723
g1532 and a[96]_not asqrt[48] ; n1724
g1533 and a[97] n1724_not ; n1725
g1534 and n1532 asqrt[48] ; n1726
g1535 nor n1725 n1726 ; n1727
g1536 nor n1527 n1721 ; n1728
g1537 and n1522_not n1728 ; n1729
g1538 and n1518_not n1729 ; n1730
g1539 and n1516_not n1730 ; n1731
g1540 and n1719_not n1731 ; n1732
g1541 and n1727 n1732_not ; n1733
g1542 nor n1723 n1733 ; n1734
g1543 and asqrt[50] n1734_not ; n1735
g1544 nor asqrt[50] n1723 ; n1736
g1545 and n1733_not n1736 ; n1737
g1546 and asqrt[49] n1715_not ; n1738
g1547 and n1710_not n1738 ; n1739
g1548 and n1706_not n1739 ; n1740
g1549 and n1704_not n1740 ; n1741
g1550 nor n1726 n1741 ; n1742
g1551 and a[98] n1742_not ; n1743
g1552 nor a[98] n1741 ; n1744
g1553 and n1726_not n1744 ; n1745
g1554 nor n1743 n1745 ; n1746
g1555 nor n1737 n1746 ; n1747
g1556 nor n1735 n1747 ; n1748
g1557 and asqrt[51] n1748_not ; n1749
g1558 nor n1535 n1540 ; n1750
g1559 and n1544_not n1750 ; n1751
g1560 and asqrt[48] n1751 ; n1752
g1561 and asqrt[48] n1750 ; n1753
g1562 and n1544 n1753_not ; n1754
g1563 nor n1752 n1754 ; n1755
g1564 nor asqrt[51] n1735 ; n1756
g1565 and n1747_not n1756 ; n1757
g1566 nor n1755 n1757 ; n1758
g1567 nor n1749 n1758 ; n1759
g1568 and asqrt[52] n1759_not ; n1760
g1569 and n1549_not n1558 ; n1761
g1570 and n1547_not n1761 ; n1762
g1571 and asqrt[48] n1762 ; n1763
g1572 nor n1547 n1549 ; n1764
g1573 and asqrt[48] n1764 ; n1765
g1574 nor n1558 n1765 ; n1766
g1575 nor n1763 n1766 ; n1767
g1576 nor asqrt[52] n1749 ; n1768
g1577 and n1758_not n1768 ; n1769
g1578 nor n1767 n1769 ; n1770
g1579 nor n1760 n1770 ; n1771
g1580 and asqrt[53] n1771_not ; n1772
g1581 and n1561_not n1567 ; n1773
g1582 and n1569_not n1773 ; n1774
g1583 and asqrt[48] n1774 ; n1775
g1584 nor n1561 n1569 ; n1776
g1585 and asqrt[48] n1776 ; n1777
g1586 nor n1567 n1777 ; n1778
g1587 nor n1775 n1778 ; n1779
g1588 nor asqrt[53] n1760 ; n1780
g1589 and n1770_not n1780 ; n1781
g1590 nor n1779 n1781 ; n1782
g1591 nor n1772 n1782 ; n1783
g1592 and asqrt[54] n1783_not ; n1784
g1593 and n1579 n1581_not ; n1785
g1594 and n1572_not n1785 ; n1786
g1595 and asqrt[48] n1786 ; n1787
g1596 nor n1572 n1581 ; n1788
g1597 and asqrt[48] n1788 ; n1789
g1598 nor n1579 n1789 ; n1790
g1599 nor n1787 n1790 ; n1791
g1600 nor asqrt[54] n1772 ; n1792
g1601 and n1782_not n1792 ; n1793
g1602 nor n1791 n1793 ; n1794
g1603 nor n1784 n1794 ; n1795
g1604 and asqrt[55] n1795_not ; n1796
g1605 and n1584_not n1591 ; n1797
g1606 and n1593_not n1797 ; n1798
g1607 and asqrt[48] n1798 ; n1799
g1608 nor n1584 n1593 ; n1800
g1609 and asqrt[48] n1800 ; n1801
g1610 nor n1591 n1801 ; n1802
g1611 nor n1799 n1802 ; n1803
g1612 nor asqrt[55] n1784 ; n1804
g1613 and n1794_not n1804 ; n1805
g1614 nor n1803 n1805 ; n1806
g1615 nor n1796 n1806 ; n1807
g1616 and asqrt[56] n1807_not ; n1808
g1617 and n1603 n1605_not ; n1809
g1618 and n1596_not n1809 ; n1810
g1619 and asqrt[48] n1810 ; n1811
g1620 nor n1596 n1605 ; n1812
g1621 and asqrt[48] n1812 ; n1813
g1622 nor n1603 n1813 ; n1814
g1623 nor n1811 n1814 ; n1815
g1624 nor asqrt[56] n1796 ; n1816
g1625 and n1806_not n1816 ; n1817
g1626 nor n1815 n1817 ; n1818
g1627 nor n1808 n1818 ; n1819
g1628 and asqrt[57] n1819_not ; n1820
g1629 and n1608_not n1615 ; n1821
g1630 and n1617_not n1821 ; n1822
g1631 and asqrt[48] n1822 ; n1823
g1632 nor n1608 n1617 ; n1824
g1633 and asqrt[48] n1824 ; n1825
g1634 nor n1615 n1825 ; n1826
g1635 nor n1823 n1826 ; n1827
g1636 nor asqrt[57] n1808 ; n1828
g1637 and n1818_not n1828 ; n1829
g1638 nor n1827 n1829 ; n1830
g1639 nor n1820 n1830 ; n1831
g1640 and asqrt[58] n1831_not ; n1832
g1641 and n1627 n1629_not ; n1833
g1642 and n1620_not n1833 ; n1834
g1643 and asqrt[48] n1834 ; n1835
g1644 nor n1620 n1629 ; n1836
g1645 and asqrt[48] n1836 ; n1837
g1646 nor n1627 n1837 ; n1838
g1647 nor n1835 n1838 ; n1839
g1648 nor asqrt[58] n1820 ; n1840
g1649 and n1830_not n1840 ; n1841
g1650 nor n1839 n1841 ; n1842
g1651 nor n1832 n1842 ; n1843
g1652 and asqrt[59] n1843_not ; n1844
g1653 and n1632_not n1639 ; n1845
g1654 and n1641_not n1845 ; n1846
g1655 and asqrt[48] n1846 ; n1847
g1656 nor n1632 n1641 ; n1848
g1657 and asqrt[48] n1848 ; n1849
g1658 nor n1639 n1849 ; n1850
g1659 nor n1847 n1850 ; n1851
g1660 nor asqrt[59] n1832 ; n1852
g1661 and n1842_not n1852 ; n1853
g1662 nor n1851 n1853 ; n1854
g1663 nor n1844 n1854 ; n1855
g1664 and asqrt[60] n1855_not ; n1856
g1665 and n1651 n1653_not ; n1857
g1666 and n1644_not n1857 ; n1858
g1667 and asqrt[48] n1858 ; n1859
g1668 nor n1644 n1653 ; n1860
g1669 and asqrt[48] n1860 ; n1861
g1670 nor n1651 n1861 ; n1862
g1671 nor n1859 n1862 ; n1863
g1672 nor asqrt[60] n1844 ; n1864
g1673 and n1854_not n1864 ; n1865
g1674 nor n1863 n1865 ; n1866
g1675 nor n1856 n1866 ; n1867
g1676 and asqrt[61] n1867_not ; n1868
g1677 and n1656_not n1663 ; n1869
g1678 and n1665_not n1869 ; n1870
g1679 and asqrt[48] n1870 ; n1871
g1680 nor n1656 n1665 ; n1872
g1681 and asqrt[48] n1872 ; n1873
g1682 nor n1663 n1873 ; n1874
g1683 nor n1871 n1874 ; n1875
g1684 nor asqrt[61] n1856 ; n1876
g1685 and n1866_not n1876 ; n1877
g1686 nor n1875 n1877 ; n1878
g1687 nor n1868 n1878 ; n1879
g1688 and asqrt[62] n1879_not ; n1880
g1689 and n1675 n1677_not ; n1881
g1690 and n1668_not n1881 ; n1882
g1691 and asqrt[48] n1882 ; n1883
g1692 nor n1668 n1677 ; n1884
g1693 and asqrt[48] n1884 ; n1885
g1694 nor n1675 n1885 ; n1886
g1695 nor n1883 n1886 ; n1887
g1696 nor asqrt[62] n1868 ; n1888
g1697 and n1878_not n1888 ; n1889
g1698 nor n1887 n1889 ; n1890
g1699 nor n1880 n1890 ; n1891
g1700 and n1680_not n1687 ; n1892
g1701 and n1689_not n1892 ; n1893
g1702 and asqrt[48] n1893 ; n1894
g1703 nor n1680 n1689 ; n1895
g1704 and asqrt[48] n1895 ; n1896
g1705 nor n1687 n1896 ; n1897
g1706 nor n1894 n1897 ; n1898
g1707 nor n1691 n1698 ; n1899
g1708 and asqrt[48] n1899 ; n1900
g1709 nor n1706 n1900 ; n1901
g1710 and n1898_not n1901 ; n1902
g1711 and n1891_not n1902 ; n1903
g1712 nor asqrt[63] n1903 ; n1904
g1713 and n1880_not n1898 ; n1905
g1714 and n1890_not n1905 ; n1906
g1715 and n1698_not asqrt[48] ; n1907
g1716 and n1691 n1907_not ; n1908
g1717 and asqrt[63] n1899_not ; n1909
g1718 and n1908_not n1909 ; n1910
g1719 nor n1694 n1715 ; n1911
g1720 and n1697_not n1911 ; n1912
g1721 and n1710_not n1912 ; n1913
g1722 and n1706_not n1913 ; n1914
g1723 and n1704_not n1914 ; n1915
g1724 nor n1910 n1915 ; n1916
g1725 and n1906_not n1916 ; n1917
g1726 nand n1904_not n1917 ; asqrt[47]
g1727 and a[94] asqrt[47] ; n1919
g1728 nor a[92] a[93] ; n1920
g1729 and a[94]_not n1920 ; n1921
g1730 nor n1919 n1921 ; n1922
g1731 and asqrt[48] n1922_not ; n1923
g1732 nor n1715 n1921 ; n1924
g1733 and n1710_not n1924 ; n1925
g1734 and n1706_not n1925 ; n1926
g1735 and n1704_not n1926 ; n1927
g1736 and n1919_not n1927 ; n1928
g1737 and a[94]_not asqrt[47] ; n1929
g1738 and a[95] n1929_not ; n1930
g1739 and n1720 asqrt[47] ; n1931
g1740 nor n1930 n1931 ; n1932
g1741 and n1928_not n1932 ; n1933
g1742 nor n1923 n1933 ; n1934
g1743 and asqrt[49] n1934_not ; n1935
g1744 nor asqrt[49] n1923 ; n1936
g1745 and n1933_not n1936 ; n1937
g1746 and asqrt[48] n1915_not ; n1938
g1747 and n1910_not n1938 ; n1939
g1748 and n1906_not n1939 ; n1940
g1749 and n1904_not n1940 ; n1941
g1750 nor n1931 n1941 ; n1942
g1751 and a[96] n1942_not ; n1943
g1752 nor a[96] n1941 ; n1944
g1753 and n1931_not n1944 ; n1945
g1754 nor n1943 n1945 ; n1946
g1755 nor n1937 n1946 ; n1947
g1756 nor n1935 n1947 ; n1948
g1757 and asqrt[50] n1948_not ; n1949
g1758 nor asqrt[50] n1935 ; n1950
g1759 and n1947_not n1950 ; n1951
g1760 nor n1727 n1732 ; n1952
g1761 and n1723_not n1952 ; n1953
g1762 and asqrt[47] n1953 ; n1954
g1763 nor n1723 n1732 ; n1955
g1764 and asqrt[47] n1955 ; n1956
g1765 and n1727 n1956_not ; n1957
g1766 nor n1954 n1957 ; n1958
g1767 nor n1951 n1958 ; n1959
g1768 nor n1949 n1959 ; n1960
g1769 and asqrt[51] n1960_not ; n1961
g1770 and n1737_not n1746 ; n1962
g1771 and n1735_not n1962 ; n1963
g1772 and asqrt[47] n1963 ; n1964
g1773 nor n1735 n1737 ; n1965
g1774 and asqrt[47] n1965 ; n1966
g1775 nor n1746 n1966 ; n1967
g1776 nor n1964 n1967 ; n1968
g1777 nor asqrt[51] n1949 ; n1969
g1778 and n1959_not n1969 ; n1970
g1779 nor n1968 n1970 ; n1971
g1780 nor n1961 n1971 ; n1972
g1781 and asqrt[52] n1972_not ; n1973
g1782 and n1749_not n1755 ; n1974
g1783 and n1757_not n1974 ; n1975
g1784 and asqrt[47] n1975 ; n1976
g1785 nor n1749 n1757 ; n1977
g1786 and asqrt[47] n1977 ; n1978
g1787 nor n1755 n1978 ; n1979
g1788 nor n1976 n1979 ; n1980
g1789 nor asqrt[52] n1961 ; n1981
g1790 and n1971_not n1981 ; n1982
g1791 nor n1980 n1982 ; n1983
g1792 nor n1973 n1983 ; n1984
g1793 and asqrt[53] n1984_not ; n1985
g1794 and n1767 n1769_not ; n1986
g1795 and n1760_not n1986 ; n1987
g1796 and asqrt[47] n1987 ; n1988
g1797 nor n1760 n1769 ; n1989
g1798 and asqrt[47] n1989 ; n1990
g1799 nor n1767 n1990 ; n1991
g1800 nor n1988 n1991 ; n1992
g1801 nor asqrt[53] n1973 ; n1993
g1802 and n1983_not n1993 ; n1994
g1803 nor n1992 n1994 ; n1995
g1804 nor n1985 n1995 ; n1996
g1805 and asqrt[54] n1996_not ; n1997
g1806 and n1772_not n1779 ; n1998
g1807 and n1781_not n1998 ; n1999
g1808 and asqrt[47] n1999 ; n2000
g1809 nor n1772 n1781 ; n2001
g1810 and asqrt[47] n2001 ; n2002
g1811 nor n1779 n2002 ; n2003
g1812 nor n2000 n2003 ; n2004
g1813 nor asqrt[54] n1985 ; n2005
g1814 and n1995_not n2005 ; n2006
g1815 nor n2004 n2006 ; n2007
g1816 nor n1997 n2007 ; n2008
g1817 and asqrt[55] n2008_not ; n2009
g1818 and n1791 n1793_not ; n2010
g1819 and n1784_not n2010 ; n2011
g1820 and asqrt[47] n2011 ; n2012
g1821 nor n1784 n1793 ; n2013
g1822 and asqrt[47] n2013 ; n2014
g1823 nor n1791 n2014 ; n2015
g1824 nor n2012 n2015 ; n2016
g1825 nor asqrt[55] n1997 ; n2017
g1826 and n2007_not n2017 ; n2018
g1827 nor n2016 n2018 ; n2019
g1828 nor n2009 n2019 ; n2020
g1829 and asqrt[56] n2020_not ; n2021
g1830 and n1796_not n1803 ; n2022
g1831 and n1805_not n2022 ; n2023
g1832 and asqrt[47] n2023 ; n2024
g1833 nor n1796 n1805 ; n2025
g1834 and asqrt[47] n2025 ; n2026
g1835 nor n1803 n2026 ; n2027
g1836 nor n2024 n2027 ; n2028
g1837 nor asqrt[56] n2009 ; n2029
g1838 and n2019_not n2029 ; n2030
g1839 nor n2028 n2030 ; n2031
g1840 nor n2021 n2031 ; n2032
g1841 and asqrt[57] n2032_not ; n2033
g1842 and n1815 n1817_not ; n2034
g1843 and n1808_not n2034 ; n2035
g1844 and asqrt[47] n2035 ; n2036
g1845 nor n1808 n1817 ; n2037
g1846 and asqrt[47] n2037 ; n2038
g1847 nor n1815 n2038 ; n2039
g1848 nor n2036 n2039 ; n2040
g1849 nor asqrt[57] n2021 ; n2041
g1850 and n2031_not n2041 ; n2042
g1851 nor n2040 n2042 ; n2043
g1852 nor n2033 n2043 ; n2044
g1853 and asqrt[58] n2044_not ; n2045
g1854 and n1820_not n1827 ; n2046
g1855 and n1829_not n2046 ; n2047
g1856 and asqrt[47] n2047 ; n2048
g1857 nor n1820 n1829 ; n2049
g1858 and asqrt[47] n2049 ; n2050
g1859 nor n1827 n2050 ; n2051
g1860 nor n2048 n2051 ; n2052
g1861 nor asqrt[58] n2033 ; n2053
g1862 and n2043_not n2053 ; n2054
g1863 nor n2052 n2054 ; n2055
g1864 nor n2045 n2055 ; n2056
g1865 and asqrt[59] n2056_not ; n2057
g1866 and n1839 n1841_not ; n2058
g1867 and n1832_not n2058 ; n2059
g1868 and asqrt[47] n2059 ; n2060
g1869 nor n1832 n1841 ; n2061
g1870 and asqrt[47] n2061 ; n2062
g1871 nor n1839 n2062 ; n2063
g1872 nor n2060 n2063 ; n2064
g1873 nor asqrt[59] n2045 ; n2065
g1874 and n2055_not n2065 ; n2066
g1875 nor n2064 n2066 ; n2067
g1876 nor n2057 n2067 ; n2068
g1877 and asqrt[60] n2068_not ; n2069
g1878 and n1844_not n1851 ; n2070
g1879 and n1853_not n2070 ; n2071
g1880 and asqrt[47] n2071 ; n2072
g1881 nor n1844 n1853 ; n2073
g1882 and asqrt[47] n2073 ; n2074
g1883 nor n1851 n2074 ; n2075
g1884 nor n2072 n2075 ; n2076
g1885 nor asqrt[60] n2057 ; n2077
g1886 and n2067_not n2077 ; n2078
g1887 nor n2076 n2078 ; n2079
g1888 nor n2069 n2079 ; n2080
g1889 and asqrt[61] n2080_not ; n2081
g1890 and n1863 n1865_not ; n2082
g1891 and n1856_not n2082 ; n2083
g1892 and asqrt[47] n2083 ; n2084
g1893 nor n1856 n1865 ; n2085
g1894 and asqrt[47] n2085 ; n2086
g1895 nor n1863 n2086 ; n2087
g1896 nor n2084 n2087 ; n2088
g1897 nor asqrt[61] n2069 ; n2089
g1898 and n2079_not n2089 ; n2090
g1899 nor n2088 n2090 ; n2091
g1900 nor n2081 n2091 ; n2092
g1901 and asqrt[62] n2092_not ; n2093
g1902 and n1868_not n1875 ; n2094
g1903 and n1877_not n2094 ; n2095
g1904 and asqrt[47] n2095 ; n2096
g1905 nor n1868 n1877 ; n2097
g1906 and asqrt[47] n2097 ; n2098
g1907 nor n1875 n2098 ; n2099
g1908 nor n2096 n2099 ; n2100
g1909 nor asqrt[62] n2081 ; n2101
g1910 and n2091_not n2101 ; n2102
g1911 nor n2100 n2102 ; n2103
g1912 nor n2093 n2103 ; n2104
g1913 and n1887 n1889_not ; n2105
g1914 and n1880_not n2105 ; n2106
g1915 and asqrt[47] n2106 ; n2107
g1916 nor n1880 n1889 ; n2108
g1917 and asqrt[47] n2108 ; n2109
g1918 nor n1887 n2109 ; n2110
g1919 nor n2107 n2110 ; n2111
g1920 nor n1891 n1898 ; n2112
g1921 and asqrt[47] n2112 ; n2113
g1922 nor n1906 n2113 ; n2114
g1923 and n2111_not n2114 ; n2115
g1924 and n2104_not n2115 ; n2116
g1925 nor asqrt[63] n2116 ; n2117
g1926 and n2093_not n2111 ; n2118
g1927 and n2103_not n2118 ; n2119
g1928 and n1898_not asqrt[47] ; n2120
g1929 and n1891 n2120_not ; n2121
g1930 and asqrt[63] n2112_not ; n2122
g1931 and n2121_not n2122 ; n2123
g1932 nor n1894 n1915 ; n2124
g1933 and n1897_not n2124 ; n2125
g1934 and n1910_not n2125 ; n2126
g1935 and n1906_not n2126 ; n2127
g1936 and n1904_not n2127 ; n2128
g1937 nor n2123 n2128 ; n2129
g1938 and n2119_not n2129 ; n2130
g1939 nand n2117_not n2130 ; asqrt[46]
g1940 and a[92] asqrt[46] ; n2132
g1941 nor a[90] a[91] ; n2133
g1942 and a[92]_not n2133 ; n2134
g1943 nor n2132 n2134 ; n2135
g1944 and asqrt[47] n2135_not ; n2136
g1945 nor n1915 n2134 ; n2137
g1946 and n1910_not n2137 ; n2138
g1947 and n1906_not n2138 ; n2139
g1948 and n1904_not n2139 ; n2140
g1949 and n2132_not n2140 ; n2141
g1950 and a[92]_not asqrt[46] ; n2142
g1951 and a[93] n2142_not ; n2143
g1952 and n1920 asqrt[46] ; n2144
g1953 nor n2143 n2144 ; n2145
g1954 and n2141_not n2145 ; n2146
g1955 nor n2136 n2146 ; n2147
g1956 and asqrt[48] n2147_not ; n2148
g1957 nor asqrt[48] n2136 ; n2149
g1958 and n2146_not n2149 ; n2150
g1959 and asqrt[47] n2128_not ; n2151
g1960 and n2123_not n2151 ; n2152
g1961 and n2119_not n2152 ; n2153
g1962 and n2117_not n2153 ; n2154
g1963 nor n2144 n2154 ; n2155
g1964 and a[94] n2155_not ; n2156
g1965 nor a[94] n2154 ; n2157
g1966 and n2144_not n2157 ; n2158
g1967 nor n2156 n2158 ; n2159
g1968 nor n2150 n2159 ; n2160
g1969 nor n2148 n2160 ; n2161
g1970 and asqrt[49] n2161_not ; n2162
g1971 nor n1923 n1928 ; n2163
g1972 and n1932_not n2163 ; n2164
g1973 and asqrt[46] n2164 ; n2165
g1974 and asqrt[46] n2163 ; n2166
g1975 and n1932 n2166_not ; n2167
g1976 nor n2165 n2167 ; n2168
g1977 nor asqrt[49] n2148 ; n2169
g1978 and n2160_not n2169 ; n2170
g1979 nor n2168 n2170 ; n2171
g1980 nor n2162 n2171 ; n2172
g1981 and asqrt[50] n2172_not ; n2173
g1982 and n1937_not n1946 ; n2174
g1983 and n1935_not n2174 ; n2175
g1984 and asqrt[46] n2175 ; n2176
g1985 nor n1935 n1937 ; n2177
g1986 and asqrt[46] n2177 ; n2178
g1987 nor n1946 n2178 ; n2179
g1988 nor n2176 n2179 ; n2180
g1989 nor asqrt[50] n2162 ; n2181
g1990 and n2171_not n2181 ; n2182
g1991 nor n2180 n2182 ; n2183
g1992 nor n2173 n2183 ; n2184
g1993 and asqrt[51] n2184_not ; n2185
g1994 nor asqrt[51] n2173 ; n2186
g1995 and n2183_not n2186 ; n2187
g1996 and n1949_not n1958 ; n2188
g1997 and n1951_not n2188 ; n2189
g1998 and asqrt[46] n2189 ; n2190
g1999 nor n1949 n1951 ; n2191
g2000 and asqrt[46] n2191 ; n2192
g2001 nor n1958 n2192 ; n2193
g2002 nor n2190 n2193 ; n2194
g2003 nor n2187 n2194 ; n2195
g2004 nor n2185 n2195 ; n2196
g2005 and asqrt[52] n2196_not ; n2197
g2006 and n1968 n1970_not ; n2198
g2007 and n1961_not n2198 ; n2199
g2008 and asqrt[46] n2199 ; n2200
g2009 nor n1961 n1970 ; n2201
g2010 and asqrt[46] n2201 ; n2202
g2011 nor n1968 n2202 ; n2203
g2012 nor n2200 n2203 ; n2204
g2013 nor asqrt[52] n2185 ; n2205
g2014 and n2195_not n2205 ; n2206
g2015 nor n2204 n2206 ; n2207
g2016 nor n2197 n2207 ; n2208
g2017 and asqrt[53] n2208_not ; n2209
g2018 and n1973_not n1980 ; n2210
g2019 and n1982_not n2210 ; n2211
g2020 and asqrt[46] n2211 ; n2212
g2021 nor n1973 n1982 ; n2213
g2022 and asqrt[46] n2213 ; n2214
g2023 nor n1980 n2214 ; n2215
g2024 nor n2212 n2215 ; n2216
g2025 nor asqrt[53] n2197 ; n2217
g2026 and n2207_not n2217 ; n2218
g2027 nor n2216 n2218 ; n2219
g2028 nor n2209 n2219 ; n2220
g2029 and asqrt[54] n2220_not ; n2221
g2030 and n1992 n1994_not ; n2222
g2031 and n1985_not n2222 ; n2223
g2032 and asqrt[46] n2223 ; n2224
g2033 nor n1985 n1994 ; n2225
g2034 and asqrt[46] n2225 ; n2226
g2035 nor n1992 n2226 ; n2227
g2036 nor n2224 n2227 ; n2228
g2037 nor asqrt[54] n2209 ; n2229
g2038 and n2219_not n2229 ; n2230
g2039 nor n2228 n2230 ; n2231
g2040 nor n2221 n2231 ; n2232
g2041 and asqrt[55] n2232_not ; n2233
g2042 and n1997_not n2004 ; n2234
g2043 and n2006_not n2234 ; n2235
g2044 and asqrt[46] n2235 ; n2236
g2045 nor n1997 n2006 ; n2237
g2046 and asqrt[46] n2237 ; n2238
g2047 nor n2004 n2238 ; n2239
g2048 nor n2236 n2239 ; n2240
g2049 nor asqrt[55] n2221 ; n2241
g2050 and n2231_not n2241 ; n2242
g2051 nor n2240 n2242 ; n2243
g2052 nor n2233 n2243 ; n2244
g2053 and asqrt[56] n2244_not ; n2245
g2054 and n2016 n2018_not ; n2246
g2055 and n2009_not n2246 ; n2247
g2056 and asqrt[46] n2247 ; n2248
g2057 nor n2009 n2018 ; n2249
g2058 and asqrt[46] n2249 ; n2250
g2059 nor n2016 n2250 ; n2251
g2060 nor n2248 n2251 ; n2252
g2061 nor asqrt[56] n2233 ; n2253
g2062 and n2243_not n2253 ; n2254
g2063 nor n2252 n2254 ; n2255
g2064 nor n2245 n2255 ; n2256
g2065 and asqrt[57] n2256_not ; n2257
g2066 and n2021_not n2028 ; n2258
g2067 and n2030_not n2258 ; n2259
g2068 and asqrt[46] n2259 ; n2260
g2069 nor n2021 n2030 ; n2261
g2070 and asqrt[46] n2261 ; n2262
g2071 nor n2028 n2262 ; n2263
g2072 nor n2260 n2263 ; n2264
g2073 nor asqrt[57] n2245 ; n2265
g2074 and n2255_not n2265 ; n2266
g2075 nor n2264 n2266 ; n2267
g2076 nor n2257 n2267 ; n2268
g2077 and asqrt[58] n2268_not ; n2269
g2078 and n2040 n2042_not ; n2270
g2079 and n2033_not n2270 ; n2271
g2080 and asqrt[46] n2271 ; n2272
g2081 nor n2033 n2042 ; n2273
g2082 and asqrt[46] n2273 ; n2274
g2083 nor n2040 n2274 ; n2275
g2084 nor n2272 n2275 ; n2276
g2085 nor asqrt[58] n2257 ; n2277
g2086 and n2267_not n2277 ; n2278
g2087 nor n2276 n2278 ; n2279
g2088 nor n2269 n2279 ; n2280
g2089 and asqrt[59] n2280_not ; n2281
g2090 and n2045_not n2052 ; n2282
g2091 and n2054_not n2282 ; n2283
g2092 and asqrt[46] n2283 ; n2284
g2093 nor n2045 n2054 ; n2285
g2094 and asqrt[46] n2285 ; n2286
g2095 nor n2052 n2286 ; n2287
g2096 nor n2284 n2287 ; n2288
g2097 nor asqrt[59] n2269 ; n2289
g2098 and n2279_not n2289 ; n2290
g2099 nor n2288 n2290 ; n2291
g2100 nor n2281 n2291 ; n2292
g2101 and asqrt[60] n2292_not ; n2293
g2102 and n2064 n2066_not ; n2294
g2103 and n2057_not n2294 ; n2295
g2104 and asqrt[46] n2295 ; n2296
g2105 nor n2057 n2066 ; n2297
g2106 and asqrt[46] n2297 ; n2298
g2107 nor n2064 n2298 ; n2299
g2108 nor n2296 n2299 ; n2300
g2109 nor asqrt[60] n2281 ; n2301
g2110 and n2291_not n2301 ; n2302
g2111 nor n2300 n2302 ; n2303
g2112 nor n2293 n2303 ; n2304
g2113 and asqrt[61] n2304_not ; n2305
g2114 and n2069_not n2076 ; n2306
g2115 and n2078_not n2306 ; n2307
g2116 and asqrt[46] n2307 ; n2308
g2117 nor n2069 n2078 ; n2309
g2118 and asqrt[46] n2309 ; n2310
g2119 nor n2076 n2310 ; n2311
g2120 nor n2308 n2311 ; n2312
g2121 nor asqrt[61] n2293 ; n2313
g2122 and n2303_not n2313 ; n2314
g2123 nor n2312 n2314 ; n2315
g2124 nor n2305 n2315 ; n2316
g2125 and asqrt[62] n2316_not ; n2317
g2126 and n2088 n2090_not ; n2318
g2127 and n2081_not n2318 ; n2319
g2128 and asqrt[46] n2319 ; n2320
g2129 nor n2081 n2090 ; n2321
g2130 and asqrt[46] n2321 ; n2322
g2131 nor n2088 n2322 ; n2323
g2132 nor n2320 n2323 ; n2324
g2133 nor asqrt[62] n2305 ; n2325
g2134 and n2315_not n2325 ; n2326
g2135 nor n2324 n2326 ; n2327
g2136 nor n2317 n2327 ; n2328
g2137 and n2093_not n2100 ; n2329
g2138 and n2102_not n2329 ; n2330
g2139 and asqrt[46] n2330 ; n2331
g2140 nor n2093 n2102 ; n2332
g2141 and asqrt[46] n2332 ; n2333
g2142 nor n2100 n2333 ; n2334
g2143 nor n2331 n2334 ; n2335
g2144 nor n2104 n2111 ; n2336
g2145 and asqrt[46] n2336 ; n2337
g2146 nor n2119 n2337 ; n2338
g2147 and n2335_not n2338 ; n2339
g2148 and n2328_not n2339 ; n2340
g2149 nor asqrt[63] n2340 ; n2341
g2150 and n2317_not n2335 ; n2342
g2151 and n2327_not n2342 ; n2343
g2152 and n2111_not asqrt[46] ; n2344
g2153 and n2104 n2344_not ; n2345
g2154 and asqrt[63] n2336_not ; n2346
g2155 and n2345_not n2346 ; n2347
g2156 nor n2107 n2128 ; n2348
g2157 and n2110_not n2348 ; n2349
g2158 and n2123_not n2349 ; n2350
g2159 and n2119_not n2350 ; n2351
g2160 and n2117_not n2351 ; n2352
g2161 nor n2347 n2352 ; n2353
g2162 and n2343_not n2353 ; n2354
g2163 nand n2341_not n2354 ; asqrt[45]
g2164 and a[90] asqrt[45] ; n2356
g2165 nor a[88] a[89] ; n2357
g2166 and a[90]_not n2357 ; n2358
g2167 nor n2356 n2358 ; n2359
g2168 and asqrt[46] n2359_not ; n2360
g2169 nor n2128 n2358 ; n2361
g2170 and n2123_not n2361 ; n2362
g2171 and n2119_not n2362 ; n2363
g2172 and n2117_not n2363 ; n2364
g2173 and n2356_not n2364 ; n2365
g2174 and a[90]_not asqrt[45] ; n2366
g2175 and a[91] n2366_not ; n2367
g2176 and n2133 asqrt[45] ; n2368
g2177 nor n2367 n2368 ; n2369
g2178 and n2365_not n2369 ; n2370
g2179 nor n2360 n2370 ; n2371
g2180 and asqrt[47] n2371_not ; n2372
g2181 nor asqrt[47] n2360 ; n2373
g2182 and n2370_not n2373 ; n2374
g2183 and asqrt[46] n2352_not ; n2375
g2184 and n2347_not n2375 ; n2376
g2185 and n2343_not n2376 ; n2377
g2186 and n2341_not n2377 ; n2378
g2187 nor n2368 n2378 ; n2379
g2188 and a[92] n2379_not ; n2380
g2189 nor a[92] n2378 ; n2381
g2190 and n2368_not n2381 ; n2382
g2191 nor n2380 n2382 ; n2383
g2192 nor n2374 n2383 ; n2384
g2193 nor n2372 n2384 ; n2385
g2194 and asqrt[48] n2385_not ; n2386
g2195 nor n2136 n2141 ; n2387
g2196 and n2145_not n2387 ; n2388
g2197 and asqrt[45] n2388 ; n2389
g2198 and asqrt[45] n2387 ; n2390
g2199 and n2145 n2390_not ; n2391
g2200 nor n2389 n2391 ; n2392
g2201 nor asqrt[48] n2372 ; n2393
g2202 and n2384_not n2393 ; n2394
g2203 nor n2392 n2394 ; n2395
g2204 nor n2386 n2395 ; n2396
g2205 and asqrt[49] n2396_not ; n2397
g2206 and n2150_not n2159 ; n2398
g2207 and n2148_not n2398 ; n2399
g2208 and asqrt[45] n2399 ; n2400
g2209 nor n2148 n2150 ; n2401
g2210 and asqrt[45] n2401 ; n2402
g2211 nor n2159 n2402 ; n2403
g2212 nor n2400 n2403 ; n2404
g2213 nor asqrt[49] n2386 ; n2405
g2214 and n2395_not n2405 ; n2406
g2215 nor n2404 n2406 ; n2407
g2216 nor n2397 n2407 ; n2408
g2217 and asqrt[50] n2408_not ; n2409
g2218 and n2162_not n2168 ; n2410
g2219 and n2170_not n2410 ; n2411
g2220 and asqrt[45] n2411 ; n2412
g2221 nor n2162 n2170 ; n2413
g2222 and asqrt[45] n2413 ; n2414
g2223 nor n2168 n2414 ; n2415
g2224 nor n2412 n2415 ; n2416
g2225 nor asqrt[50] n2397 ; n2417
g2226 and n2407_not n2417 ; n2418
g2227 nor n2416 n2418 ; n2419
g2228 nor n2409 n2419 ; n2420
g2229 and asqrt[51] n2420_not ; n2421
g2230 and n2180 n2182_not ; n2422
g2231 and n2173_not n2422 ; n2423
g2232 and asqrt[45] n2423 ; n2424
g2233 nor n2173 n2182 ; n2425
g2234 and asqrt[45] n2425 ; n2426
g2235 nor n2180 n2426 ; n2427
g2236 nor n2424 n2427 ; n2428
g2237 nor asqrt[51] n2409 ; n2429
g2238 and n2419_not n2429 ; n2430
g2239 nor n2428 n2430 ; n2431
g2240 nor n2421 n2431 ; n2432
g2241 and asqrt[52] n2432_not ; n2433
g2242 nor asqrt[52] n2421 ; n2434
g2243 and n2431_not n2434 ; n2435
g2244 and n2185_not n2194 ; n2436
g2245 and n2187_not n2436 ; n2437
g2246 and asqrt[45] n2437 ; n2438
g2247 nor n2185 n2187 ; n2439
g2248 and asqrt[45] n2439 ; n2440
g2249 nor n2194 n2440 ; n2441
g2250 nor n2438 n2441 ; n2442
g2251 nor n2435 n2442 ; n2443
g2252 nor n2433 n2443 ; n2444
g2253 and asqrt[53] n2444_not ; n2445
g2254 and n2204 n2206_not ; n2446
g2255 and n2197_not n2446 ; n2447
g2256 and asqrt[45] n2447 ; n2448
g2257 nor n2197 n2206 ; n2449
g2258 and asqrt[45] n2449 ; n2450
g2259 nor n2204 n2450 ; n2451
g2260 nor n2448 n2451 ; n2452
g2261 nor asqrt[53] n2433 ; n2453
g2262 and n2443_not n2453 ; n2454
g2263 nor n2452 n2454 ; n2455
g2264 nor n2445 n2455 ; n2456
g2265 and asqrt[54] n2456_not ; n2457
g2266 and n2209_not n2216 ; n2458
g2267 and n2218_not n2458 ; n2459
g2268 and asqrt[45] n2459 ; n2460
g2269 nor n2209 n2218 ; n2461
g2270 and asqrt[45] n2461 ; n2462
g2271 nor n2216 n2462 ; n2463
g2272 nor n2460 n2463 ; n2464
g2273 nor asqrt[54] n2445 ; n2465
g2274 and n2455_not n2465 ; n2466
g2275 nor n2464 n2466 ; n2467
g2276 nor n2457 n2467 ; n2468
g2277 and asqrt[55] n2468_not ; n2469
g2278 and n2228 n2230_not ; n2470
g2279 and n2221_not n2470 ; n2471
g2280 and asqrt[45] n2471 ; n2472
g2281 nor n2221 n2230 ; n2473
g2282 and asqrt[45] n2473 ; n2474
g2283 nor n2228 n2474 ; n2475
g2284 nor n2472 n2475 ; n2476
g2285 nor asqrt[55] n2457 ; n2477
g2286 and n2467_not n2477 ; n2478
g2287 nor n2476 n2478 ; n2479
g2288 nor n2469 n2479 ; n2480
g2289 and asqrt[56] n2480_not ; n2481
g2290 and n2233_not n2240 ; n2482
g2291 and n2242_not n2482 ; n2483
g2292 and asqrt[45] n2483 ; n2484
g2293 nor n2233 n2242 ; n2485
g2294 and asqrt[45] n2485 ; n2486
g2295 nor n2240 n2486 ; n2487
g2296 nor n2484 n2487 ; n2488
g2297 nor asqrt[56] n2469 ; n2489
g2298 and n2479_not n2489 ; n2490
g2299 nor n2488 n2490 ; n2491
g2300 nor n2481 n2491 ; n2492
g2301 and asqrt[57] n2492_not ; n2493
g2302 and n2252 n2254_not ; n2494
g2303 and n2245_not n2494 ; n2495
g2304 and asqrt[45] n2495 ; n2496
g2305 nor n2245 n2254 ; n2497
g2306 and asqrt[45] n2497 ; n2498
g2307 nor n2252 n2498 ; n2499
g2308 nor n2496 n2499 ; n2500
g2309 nor asqrt[57] n2481 ; n2501
g2310 and n2491_not n2501 ; n2502
g2311 nor n2500 n2502 ; n2503
g2312 nor n2493 n2503 ; n2504
g2313 and asqrt[58] n2504_not ; n2505
g2314 and n2257_not n2264 ; n2506
g2315 and n2266_not n2506 ; n2507
g2316 and asqrt[45] n2507 ; n2508
g2317 nor n2257 n2266 ; n2509
g2318 and asqrt[45] n2509 ; n2510
g2319 nor n2264 n2510 ; n2511
g2320 nor n2508 n2511 ; n2512
g2321 nor asqrt[58] n2493 ; n2513
g2322 and n2503_not n2513 ; n2514
g2323 nor n2512 n2514 ; n2515
g2324 nor n2505 n2515 ; n2516
g2325 and asqrt[59] n2516_not ; n2517
g2326 and n2276 n2278_not ; n2518
g2327 and n2269_not n2518 ; n2519
g2328 and asqrt[45] n2519 ; n2520
g2329 nor n2269 n2278 ; n2521
g2330 and asqrt[45] n2521 ; n2522
g2331 nor n2276 n2522 ; n2523
g2332 nor n2520 n2523 ; n2524
g2333 nor asqrt[59] n2505 ; n2525
g2334 and n2515_not n2525 ; n2526
g2335 nor n2524 n2526 ; n2527
g2336 nor n2517 n2527 ; n2528
g2337 and asqrt[60] n2528_not ; n2529
g2338 and n2281_not n2288 ; n2530
g2339 and n2290_not n2530 ; n2531
g2340 and asqrt[45] n2531 ; n2532
g2341 nor n2281 n2290 ; n2533
g2342 and asqrt[45] n2533 ; n2534
g2343 nor n2288 n2534 ; n2535
g2344 nor n2532 n2535 ; n2536
g2345 nor asqrt[60] n2517 ; n2537
g2346 and n2527_not n2537 ; n2538
g2347 nor n2536 n2538 ; n2539
g2348 nor n2529 n2539 ; n2540
g2349 and asqrt[61] n2540_not ; n2541
g2350 and n2300 n2302_not ; n2542
g2351 and n2293_not n2542 ; n2543
g2352 and asqrt[45] n2543 ; n2544
g2353 nor n2293 n2302 ; n2545
g2354 and asqrt[45] n2545 ; n2546
g2355 nor n2300 n2546 ; n2547
g2356 nor n2544 n2547 ; n2548
g2357 nor asqrt[61] n2529 ; n2549
g2358 and n2539_not n2549 ; n2550
g2359 nor n2548 n2550 ; n2551
g2360 nor n2541 n2551 ; n2552
g2361 and asqrt[62] n2552_not ; n2553
g2362 and n2305_not n2312 ; n2554
g2363 and n2314_not n2554 ; n2555
g2364 and asqrt[45] n2555 ; n2556
g2365 nor n2305 n2314 ; n2557
g2366 and asqrt[45] n2557 ; n2558
g2367 nor n2312 n2558 ; n2559
g2368 nor n2556 n2559 ; n2560
g2369 nor asqrt[62] n2541 ; n2561
g2370 and n2551_not n2561 ; n2562
g2371 nor n2560 n2562 ; n2563
g2372 nor n2553 n2563 ; n2564
g2373 and n2324 n2326_not ; n2565
g2374 and n2317_not n2565 ; n2566
g2375 and asqrt[45] n2566 ; n2567
g2376 nor n2317 n2326 ; n2568
g2377 and asqrt[45] n2568 ; n2569
g2378 nor n2324 n2569 ; n2570
g2379 nor n2567 n2570 ; n2571
g2380 nor n2328 n2335 ; n2572
g2381 and asqrt[45] n2572 ; n2573
g2382 nor n2343 n2573 ; n2574
g2383 and n2571_not n2574 ; n2575
g2384 and n2564_not n2575 ; n2576
g2385 nor asqrt[63] n2576 ; n2577
g2386 and n2553_not n2571 ; n2578
g2387 and n2563_not n2578 ; n2579
g2388 and n2335_not asqrt[45] ; n2580
g2389 and n2328 n2580_not ; n2581
g2390 and asqrt[63] n2572_not ; n2582
g2391 and n2581_not n2582 ; n2583
g2392 nor n2331 n2352 ; n2584
g2393 and n2334_not n2584 ; n2585
g2394 and n2347_not n2585 ; n2586
g2395 and n2343_not n2586 ; n2587
g2396 and n2341_not n2587 ; n2588
g2397 nor n2583 n2588 ; n2589
g2398 and n2579_not n2589 ; n2590
g2399 nand n2577_not n2590 ; asqrt[44]
g2400 and a[88] asqrt[44] ; n2592
g2401 nor a[86] a[87] ; n2593
g2402 and a[88]_not n2593 ; n2594
g2403 nor n2592 n2594 ; n2595
g2404 and asqrt[45] n2595_not ; n2596
g2405 nor n2352 n2594 ; n2597
g2406 and n2347_not n2597 ; n2598
g2407 and n2343_not n2598 ; n2599
g2408 and n2341_not n2599 ; n2600
g2409 and n2592_not n2600 ; n2601
g2410 and a[88]_not asqrt[44] ; n2602
g2411 and a[89] n2602_not ; n2603
g2412 and n2357 asqrt[44] ; n2604
g2413 nor n2603 n2604 ; n2605
g2414 and n2601_not n2605 ; n2606
g2415 nor n2596 n2606 ; n2607
g2416 and asqrt[46] n2607_not ; n2608
g2417 nor asqrt[46] n2596 ; n2609
g2418 and n2606_not n2609 ; n2610
g2419 and asqrt[45] n2588_not ; n2611
g2420 and n2583_not n2611 ; n2612
g2421 and n2579_not n2612 ; n2613
g2422 and n2577_not n2613 ; n2614
g2423 nor n2604 n2614 ; n2615
g2424 and a[90] n2615_not ; n2616
g2425 nor a[90] n2614 ; n2617
g2426 and n2604_not n2617 ; n2618
g2427 nor n2616 n2618 ; n2619
g2428 nor n2610 n2619 ; n2620
g2429 nor n2608 n2620 ; n2621
g2430 and asqrt[47] n2621_not ; n2622
g2431 nor n2360 n2365 ; n2623
g2432 and n2369_not n2623 ; n2624
g2433 and asqrt[44] n2624 ; n2625
g2434 and asqrt[44] n2623 ; n2626
g2435 and n2369 n2626_not ; n2627
g2436 nor n2625 n2627 ; n2628
g2437 nor asqrt[47] n2608 ; n2629
g2438 and n2620_not n2629 ; n2630
g2439 nor n2628 n2630 ; n2631
g2440 nor n2622 n2631 ; n2632
g2441 and asqrt[48] n2632_not ; n2633
g2442 and n2374_not n2383 ; n2634
g2443 and n2372_not n2634 ; n2635
g2444 and asqrt[44] n2635 ; n2636
g2445 nor n2372 n2374 ; n2637
g2446 and asqrt[44] n2637 ; n2638
g2447 nor n2383 n2638 ; n2639
g2448 nor n2636 n2639 ; n2640
g2449 nor asqrt[48] n2622 ; n2641
g2450 and n2631_not n2641 ; n2642
g2451 nor n2640 n2642 ; n2643
g2452 nor n2633 n2643 ; n2644
g2453 and asqrt[49] n2644_not ; n2645
g2454 and n2386_not n2392 ; n2646
g2455 and n2394_not n2646 ; n2647
g2456 and asqrt[44] n2647 ; n2648
g2457 nor n2386 n2394 ; n2649
g2458 and asqrt[44] n2649 ; n2650
g2459 nor n2392 n2650 ; n2651
g2460 nor n2648 n2651 ; n2652
g2461 nor asqrt[49] n2633 ; n2653
g2462 and n2643_not n2653 ; n2654
g2463 nor n2652 n2654 ; n2655
g2464 nor n2645 n2655 ; n2656
g2465 and asqrt[50] n2656_not ; n2657
g2466 and n2404 n2406_not ; n2658
g2467 and n2397_not n2658 ; n2659
g2468 and asqrt[44] n2659 ; n2660
g2469 nor n2397 n2406 ; n2661
g2470 and asqrt[44] n2661 ; n2662
g2471 nor n2404 n2662 ; n2663
g2472 nor n2660 n2663 ; n2664
g2473 nor asqrt[50] n2645 ; n2665
g2474 and n2655_not n2665 ; n2666
g2475 nor n2664 n2666 ; n2667
g2476 nor n2657 n2667 ; n2668
g2477 and asqrt[51] n2668_not ; n2669
g2478 and n2409_not n2416 ; n2670
g2479 and n2418_not n2670 ; n2671
g2480 and asqrt[44] n2671 ; n2672
g2481 nor n2409 n2418 ; n2673
g2482 and asqrt[44] n2673 ; n2674
g2483 nor n2416 n2674 ; n2675
g2484 nor n2672 n2675 ; n2676
g2485 nor asqrt[51] n2657 ; n2677
g2486 and n2667_not n2677 ; n2678
g2487 nor n2676 n2678 ; n2679
g2488 nor n2669 n2679 ; n2680
g2489 and asqrt[52] n2680_not ; n2681
g2490 and n2428 n2430_not ; n2682
g2491 and n2421_not n2682 ; n2683
g2492 and asqrt[44] n2683 ; n2684
g2493 nor n2421 n2430 ; n2685
g2494 and asqrt[44] n2685 ; n2686
g2495 nor n2428 n2686 ; n2687
g2496 nor n2684 n2687 ; n2688
g2497 nor asqrt[52] n2669 ; n2689
g2498 and n2679_not n2689 ; n2690
g2499 nor n2688 n2690 ; n2691
g2500 nor n2681 n2691 ; n2692
g2501 and asqrt[53] n2692_not ; n2693
g2502 nor asqrt[53] n2681 ; n2694
g2503 and n2691_not n2694 ; n2695
g2504 and n2433_not n2442 ; n2696
g2505 and n2435_not n2696 ; n2697
g2506 and asqrt[44] n2697 ; n2698
g2507 nor n2433 n2435 ; n2699
g2508 and asqrt[44] n2699 ; n2700
g2509 nor n2442 n2700 ; n2701
g2510 nor n2698 n2701 ; n2702
g2511 nor n2695 n2702 ; n2703
g2512 nor n2693 n2703 ; n2704
g2513 and asqrt[54] n2704_not ; n2705
g2514 and n2452 n2454_not ; n2706
g2515 and n2445_not n2706 ; n2707
g2516 and asqrt[44] n2707 ; n2708
g2517 nor n2445 n2454 ; n2709
g2518 and asqrt[44] n2709 ; n2710
g2519 nor n2452 n2710 ; n2711
g2520 nor n2708 n2711 ; n2712
g2521 nor asqrt[54] n2693 ; n2713
g2522 and n2703_not n2713 ; n2714
g2523 nor n2712 n2714 ; n2715
g2524 nor n2705 n2715 ; n2716
g2525 and asqrt[55] n2716_not ; n2717
g2526 and n2457_not n2464 ; n2718
g2527 and n2466_not n2718 ; n2719
g2528 and asqrt[44] n2719 ; n2720
g2529 nor n2457 n2466 ; n2721
g2530 and asqrt[44] n2721 ; n2722
g2531 nor n2464 n2722 ; n2723
g2532 nor n2720 n2723 ; n2724
g2533 nor asqrt[55] n2705 ; n2725
g2534 and n2715_not n2725 ; n2726
g2535 nor n2724 n2726 ; n2727
g2536 nor n2717 n2727 ; n2728
g2537 and asqrt[56] n2728_not ; n2729
g2538 and n2476 n2478_not ; n2730
g2539 and n2469_not n2730 ; n2731
g2540 and asqrt[44] n2731 ; n2732
g2541 nor n2469 n2478 ; n2733
g2542 and asqrt[44] n2733 ; n2734
g2543 nor n2476 n2734 ; n2735
g2544 nor n2732 n2735 ; n2736
g2545 nor asqrt[56] n2717 ; n2737
g2546 and n2727_not n2737 ; n2738
g2547 nor n2736 n2738 ; n2739
g2548 nor n2729 n2739 ; n2740
g2549 and asqrt[57] n2740_not ; n2741
g2550 and n2481_not n2488 ; n2742
g2551 and n2490_not n2742 ; n2743
g2552 and asqrt[44] n2743 ; n2744
g2553 nor n2481 n2490 ; n2745
g2554 and asqrt[44] n2745 ; n2746
g2555 nor n2488 n2746 ; n2747
g2556 nor n2744 n2747 ; n2748
g2557 nor asqrt[57] n2729 ; n2749
g2558 and n2739_not n2749 ; n2750
g2559 nor n2748 n2750 ; n2751
g2560 nor n2741 n2751 ; n2752
g2561 and asqrt[58] n2752_not ; n2753
g2562 and n2500 n2502_not ; n2754
g2563 and n2493_not n2754 ; n2755
g2564 and asqrt[44] n2755 ; n2756
g2565 nor n2493 n2502 ; n2757
g2566 and asqrt[44] n2757 ; n2758
g2567 nor n2500 n2758 ; n2759
g2568 nor n2756 n2759 ; n2760
g2569 nor asqrt[58] n2741 ; n2761
g2570 and n2751_not n2761 ; n2762
g2571 nor n2760 n2762 ; n2763
g2572 nor n2753 n2763 ; n2764
g2573 and asqrt[59] n2764_not ; n2765
g2574 and n2505_not n2512 ; n2766
g2575 and n2514_not n2766 ; n2767
g2576 and asqrt[44] n2767 ; n2768
g2577 nor n2505 n2514 ; n2769
g2578 and asqrt[44] n2769 ; n2770
g2579 nor n2512 n2770 ; n2771
g2580 nor n2768 n2771 ; n2772
g2581 nor asqrt[59] n2753 ; n2773
g2582 and n2763_not n2773 ; n2774
g2583 nor n2772 n2774 ; n2775
g2584 nor n2765 n2775 ; n2776
g2585 and asqrt[60] n2776_not ; n2777
g2586 and n2524 n2526_not ; n2778
g2587 and n2517_not n2778 ; n2779
g2588 and asqrt[44] n2779 ; n2780
g2589 nor n2517 n2526 ; n2781
g2590 and asqrt[44] n2781 ; n2782
g2591 nor n2524 n2782 ; n2783
g2592 nor n2780 n2783 ; n2784
g2593 nor asqrt[60] n2765 ; n2785
g2594 and n2775_not n2785 ; n2786
g2595 nor n2784 n2786 ; n2787
g2596 nor n2777 n2787 ; n2788
g2597 and asqrt[61] n2788_not ; n2789
g2598 and n2529_not n2536 ; n2790
g2599 and n2538_not n2790 ; n2791
g2600 and asqrt[44] n2791 ; n2792
g2601 nor n2529 n2538 ; n2793
g2602 and asqrt[44] n2793 ; n2794
g2603 nor n2536 n2794 ; n2795
g2604 nor n2792 n2795 ; n2796
g2605 nor asqrt[61] n2777 ; n2797
g2606 and n2787_not n2797 ; n2798
g2607 nor n2796 n2798 ; n2799
g2608 nor n2789 n2799 ; n2800
g2609 and asqrt[62] n2800_not ; n2801
g2610 and n2548 n2550_not ; n2802
g2611 and n2541_not n2802 ; n2803
g2612 and asqrt[44] n2803 ; n2804
g2613 nor n2541 n2550 ; n2805
g2614 and asqrt[44] n2805 ; n2806
g2615 nor n2548 n2806 ; n2807
g2616 nor n2804 n2807 ; n2808
g2617 nor asqrt[62] n2789 ; n2809
g2618 and n2799_not n2809 ; n2810
g2619 nor n2808 n2810 ; n2811
g2620 nor n2801 n2811 ; n2812
g2621 and n2553_not n2560 ; n2813
g2622 and n2562_not n2813 ; n2814
g2623 and asqrt[44] n2814 ; n2815
g2624 nor n2553 n2562 ; n2816
g2625 and asqrt[44] n2816 ; n2817
g2626 nor n2560 n2817 ; n2818
g2627 nor n2815 n2818 ; n2819
g2628 nor n2564 n2571 ; n2820
g2629 and asqrt[44] n2820 ; n2821
g2630 nor n2579 n2821 ; n2822
g2631 and n2819_not n2822 ; n2823
g2632 and n2812_not n2823 ; n2824
g2633 nor asqrt[63] n2824 ; n2825
g2634 and n2801_not n2819 ; n2826
g2635 and n2811_not n2826 ; n2827
g2636 and n2571_not asqrt[44] ; n2828
g2637 and n2564 n2828_not ; n2829
g2638 and asqrt[63] n2820_not ; n2830
g2639 and n2829_not n2830 ; n2831
g2640 nor n2567 n2588 ; n2832
g2641 and n2570_not n2832 ; n2833
g2642 and n2583_not n2833 ; n2834
g2643 and n2579_not n2834 ; n2835
g2644 and n2577_not n2835 ; n2836
g2645 nor n2831 n2836 ; n2837
g2646 and n2827_not n2837 ; n2838
g2647 nand n2825_not n2838 ; asqrt[43]
g2648 and a[86] asqrt[43] ; n2840
g2649 nor a[84] a[85] ; n2841
g2650 and a[86]_not n2841 ; n2842
g2651 nor n2840 n2842 ; n2843
g2652 and asqrt[44] n2843_not ; n2844
g2653 nor n2588 n2842 ; n2845
g2654 and n2583_not n2845 ; n2846
g2655 and n2579_not n2846 ; n2847
g2656 and n2577_not n2847 ; n2848
g2657 and n2840_not n2848 ; n2849
g2658 and a[86]_not asqrt[43] ; n2850
g2659 and a[87] n2850_not ; n2851
g2660 and n2593 asqrt[43] ; n2852
g2661 nor n2851 n2852 ; n2853
g2662 and n2849_not n2853 ; n2854
g2663 nor n2844 n2854 ; n2855
g2664 and asqrt[45] n2855_not ; n2856
g2665 nor asqrt[45] n2844 ; n2857
g2666 and n2854_not n2857 ; n2858
g2667 and asqrt[44] n2836_not ; n2859
g2668 and n2831_not n2859 ; n2860
g2669 and n2827_not n2860 ; n2861
g2670 and n2825_not n2861 ; n2862
g2671 nor n2852 n2862 ; n2863
g2672 and a[88] n2863_not ; n2864
g2673 nor a[88] n2862 ; n2865
g2674 and n2852_not n2865 ; n2866
g2675 nor n2864 n2866 ; n2867
g2676 nor n2858 n2867 ; n2868
g2677 nor n2856 n2868 ; n2869
g2678 and asqrt[46] n2869_not ; n2870
g2679 nor n2596 n2601 ; n2871
g2680 and n2605_not n2871 ; n2872
g2681 and asqrt[43] n2872 ; n2873
g2682 and asqrt[43] n2871 ; n2874
g2683 and n2605 n2874_not ; n2875
g2684 nor n2873 n2875 ; n2876
g2685 nor asqrt[46] n2856 ; n2877
g2686 and n2868_not n2877 ; n2878
g2687 nor n2876 n2878 ; n2879
g2688 nor n2870 n2879 ; n2880
g2689 and asqrt[47] n2880_not ; n2881
g2690 and n2610_not n2619 ; n2882
g2691 and n2608_not n2882 ; n2883
g2692 and asqrt[43] n2883 ; n2884
g2693 nor n2608 n2610 ; n2885
g2694 and asqrt[43] n2885 ; n2886
g2695 nor n2619 n2886 ; n2887
g2696 nor n2884 n2887 ; n2888
g2697 nor asqrt[47] n2870 ; n2889
g2698 and n2879_not n2889 ; n2890
g2699 nor n2888 n2890 ; n2891
g2700 nor n2881 n2891 ; n2892
g2701 and asqrt[48] n2892_not ; n2893
g2702 and n2622_not n2628 ; n2894
g2703 and n2630_not n2894 ; n2895
g2704 and asqrt[43] n2895 ; n2896
g2705 nor n2622 n2630 ; n2897
g2706 and asqrt[43] n2897 ; n2898
g2707 nor n2628 n2898 ; n2899
g2708 nor n2896 n2899 ; n2900
g2709 nor asqrt[48] n2881 ; n2901
g2710 and n2891_not n2901 ; n2902
g2711 nor n2900 n2902 ; n2903
g2712 nor n2893 n2903 ; n2904
g2713 and asqrt[49] n2904_not ; n2905
g2714 and n2640 n2642_not ; n2906
g2715 and n2633_not n2906 ; n2907
g2716 and asqrt[43] n2907 ; n2908
g2717 nor n2633 n2642 ; n2909
g2718 and asqrt[43] n2909 ; n2910
g2719 nor n2640 n2910 ; n2911
g2720 nor n2908 n2911 ; n2912
g2721 nor asqrt[49] n2893 ; n2913
g2722 and n2903_not n2913 ; n2914
g2723 nor n2912 n2914 ; n2915
g2724 nor n2905 n2915 ; n2916
g2725 and asqrt[50] n2916_not ; n2917
g2726 and n2645_not n2652 ; n2918
g2727 and n2654_not n2918 ; n2919
g2728 and asqrt[43] n2919 ; n2920
g2729 nor n2645 n2654 ; n2921
g2730 and asqrt[43] n2921 ; n2922
g2731 nor n2652 n2922 ; n2923
g2732 nor n2920 n2923 ; n2924
g2733 nor asqrt[50] n2905 ; n2925
g2734 and n2915_not n2925 ; n2926
g2735 nor n2924 n2926 ; n2927
g2736 nor n2917 n2927 ; n2928
g2737 and asqrt[51] n2928_not ; n2929
g2738 and n2664 n2666_not ; n2930
g2739 and n2657_not n2930 ; n2931
g2740 and asqrt[43] n2931 ; n2932
g2741 nor n2657 n2666 ; n2933
g2742 and asqrt[43] n2933 ; n2934
g2743 nor n2664 n2934 ; n2935
g2744 nor n2932 n2935 ; n2936
g2745 nor asqrt[51] n2917 ; n2937
g2746 and n2927_not n2937 ; n2938
g2747 nor n2936 n2938 ; n2939
g2748 nor n2929 n2939 ; n2940
g2749 and asqrt[52] n2940_not ; n2941
g2750 and n2669_not n2676 ; n2942
g2751 and n2678_not n2942 ; n2943
g2752 and asqrt[43] n2943 ; n2944
g2753 nor n2669 n2678 ; n2945
g2754 and asqrt[43] n2945 ; n2946
g2755 nor n2676 n2946 ; n2947
g2756 nor n2944 n2947 ; n2948
g2757 nor asqrt[52] n2929 ; n2949
g2758 and n2939_not n2949 ; n2950
g2759 nor n2948 n2950 ; n2951
g2760 nor n2941 n2951 ; n2952
g2761 and asqrt[53] n2952_not ; n2953
g2762 and n2688 n2690_not ; n2954
g2763 and n2681_not n2954 ; n2955
g2764 and asqrt[43] n2955 ; n2956
g2765 nor n2681 n2690 ; n2957
g2766 and asqrt[43] n2957 ; n2958
g2767 nor n2688 n2958 ; n2959
g2768 nor n2956 n2959 ; n2960
g2769 nor asqrt[53] n2941 ; n2961
g2770 and n2951_not n2961 ; n2962
g2771 nor n2960 n2962 ; n2963
g2772 nor n2953 n2963 ; n2964
g2773 and asqrt[54] n2964_not ; n2965
g2774 nor asqrt[54] n2953 ; n2966
g2775 and n2963_not n2966 ; n2967
g2776 and n2693_not n2702 ; n2968
g2777 and n2695_not n2968 ; n2969
g2778 and asqrt[43] n2969 ; n2970
g2779 nor n2693 n2695 ; n2971
g2780 and asqrt[43] n2971 ; n2972
g2781 nor n2702 n2972 ; n2973
g2782 nor n2970 n2973 ; n2974
g2783 nor n2967 n2974 ; n2975
g2784 nor n2965 n2975 ; n2976
g2785 and asqrt[55] n2976_not ; n2977
g2786 and n2712 n2714_not ; n2978
g2787 and n2705_not n2978 ; n2979
g2788 and asqrt[43] n2979 ; n2980
g2789 nor n2705 n2714 ; n2981
g2790 and asqrt[43] n2981 ; n2982
g2791 nor n2712 n2982 ; n2983
g2792 nor n2980 n2983 ; n2984
g2793 nor asqrt[55] n2965 ; n2985
g2794 and n2975_not n2985 ; n2986
g2795 nor n2984 n2986 ; n2987
g2796 nor n2977 n2987 ; n2988
g2797 and asqrt[56] n2988_not ; n2989
g2798 and n2717_not n2724 ; n2990
g2799 and n2726_not n2990 ; n2991
g2800 and asqrt[43] n2991 ; n2992
g2801 nor n2717 n2726 ; n2993
g2802 and asqrt[43] n2993 ; n2994
g2803 nor n2724 n2994 ; n2995
g2804 nor n2992 n2995 ; n2996
g2805 nor asqrt[56] n2977 ; n2997
g2806 and n2987_not n2997 ; n2998
g2807 nor n2996 n2998 ; n2999
g2808 nor n2989 n2999 ; n3000
g2809 and asqrt[57] n3000_not ; n3001
g2810 and n2736 n2738_not ; n3002
g2811 and n2729_not n3002 ; n3003
g2812 and asqrt[43] n3003 ; n3004
g2813 nor n2729 n2738 ; n3005
g2814 and asqrt[43] n3005 ; n3006
g2815 nor n2736 n3006 ; n3007
g2816 nor n3004 n3007 ; n3008
g2817 nor asqrt[57] n2989 ; n3009
g2818 and n2999_not n3009 ; n3010
g2819 nor n3008 n3010 ; n3011
g2820 nor n3001 n3011 ; n3012
g2821 and asqrt[58] n3012_not ; n3013
g2822 and n2741_not n2748 ; n3014
g2823 and n2750_not n3014 ; n3015
g2824 and asqrt[43] n3015 ; n3016
g2825 nor n2741 n2750 ; n3017
g2826 and asqrt[43] n3017 ; n3018
g2827 nor n2748 n3018 ; n3019
g2828 nor n3016 n3019 ; n3020
g2829 nor asqrt[58] n3001 ; n3021
g2830 and n3011_not n3021 ; n3022
g2831 nor n3020 n3022 ; n3023
g2832 nor n3013 n3023 ; n3024
g2833 and asqrt[59] n3024_not ; n3025
g2834 and n2760 n2762_not ; n3026
g2835 and n2753_not n3026 ; n3027
g2836 and asqrt[43] n3027 ; n3028
g2837 nor n2753 n2762 ; n3029
g2838 and asqrt[43] n3029 ; n3030
g2839 nor n2760 n3030 ; n3031
g2840 nor n3028 n3031 ; n3032
g2841 nor asqrt[59] n3013 ; n3033
g2842 and n3023_not n3033 ; n3034
g2843 nor n3032 n3034 ; n3035
g2844 nor n3025 n3035 ; n3036
g2845 and asqrt[60] n3036_not ; n3037
g2846 and n2765_not n2772 ; n3038
g2847 and n2774_not n3038 ; n3039
g2848 and asqrt[43] n3039 ; n3040
g2849 nor n2765 n2774 ; n3041
g2850 and asqrt[43] n3041 ; n3042
g2851 nor n2772 n3042 ; n3043
g2852 nor n3040 n3043 ; n3044
g2853 nor asqrt[60] n3025 ; n3045
g2854 and n3035_not n3045 ; n3046
g2855 nor n3044 n3046 ; n3047
g2856 nor n3037 n3047 ; n3048
g2857 and asqrt[61] n3048_not ; n3049
g2858 and n2784 n2786_not ; n3050
g2859 and n2777_not n3050 ; n3051
g2860 and asqrt[43] n3051 ; n3052
g2861 nor n2777 n2786 ; n3053
g2862 and asqrt[43] n3053 ; n3054
g2863 nor n2784 n3054 ; n3055
g2864 nor n3052 n3055 ; n3056
g2865 nor asqrt[61] n3037 ; n3057
g2866 and n3047_not n3057 ; n3058
g2867 nor n3056 n3058 ; n3059
g2868 nor n3049 n3059 ; n3060
g2869 and asqrt[62] n3060_not ; n3061
g2870 and n2789_not n2796 ; n3062
g2871 and n2798_not n3062 ; n3063
g2872 and asqrt[43] n3063 ; n3064
g2873 nor n2789 n2798 ; n3065
g2874 and asqrt[43] n3065 ; n3066
g2875 nor n2796 n3066 ; n3067
g2876 nor n3064 n3067 ; n3068
g2877 nor asqrt[62] n3049 ; n3069
g2878 and n3059_not n3069 ; n3070
g2879 nor n3068 n3070 ; n3071
g2880 nor n3061 n3071 ; n3072
g2881 and n2808 n2810_not ; n3073
g2882 and n2801_not n3073 ; n3074
g2883 and asqrt[43] n3074 ; n3075
g2884 nor n2801 n2810 ; n3076
g2885 and asqrt[43] n3076 ; n3077
g2886 nor n2808 n3077 ; n3078
g2887 nor n3075 n3078 ; n3079
g2888 nor n2812 n2819 ; n3080
g2889 and asqrt[43] n3080 ; n3081
g2890 nor n2827 n3081 ; n3082
g2891 and n3079_not n3082 ; n3083
g2892 and n3072_not n3083 ; n3084
g2893 nor asqrt[63] n3084 ; n3085
g2894 and n3061_not n3079 ; n3086
g2895 and n3071_not n3086 ; n3087
g2896 and n2819_not asqrt[43] ; n3088
g2897 and n2812 n3088_not ; n3089
g2898 and asqrt[63] n3080_not ; n3090
g2899 and n3089_not n3090 ; n3091
g2900 nor n2815 n2836 ; n3092
g2901 and n2818_not n3092 ; n3093
g2902 and n2831_not n3093 ; n3094
g2903 and n2827_not n3094 ; n3095
g2904 and n2825_not n3095 ; n3096
g2905 nor n3091 n3096 ; n3097
g2906 and n3087_not n3097 ; n3098
g2907 nand n3085_not n3098 ; asqrt[42]
g2908 and a[84] asqrt[42] ; n3100
g2909 nor a[82] a[83] ; n3101
g2910 and a[84]_not n3101 ; n3102
g2911 nor n3100 n3102 ; n3103
g2912 and asqrt[43] n3103_not ; n3104
g2913 nor n2836 n3102 ; n3105
g2914 and n2831_not n3105 ; n3106
g2915 and n2827_not n3106 ; n3107
g2916 and n2825_not n3107 ; n3108
g2917 and n3100_not n3108 ; n3109
g2918 and a[84]_not asqrt[42] ; n3110
g2919 and a[85] n3110_not ; n3111
g2920 and n2841 asqrt[42] ; n3112
g2921 nor n3111 n3112 ; n3113
g2922 and n3109_not n3113 ; n3114
g2923 nor n3104 n3114 ; n3115
g2924 and asqrt[44] n3115_not ; n3116
g2925 nor asqrt[44] n3104 ; n3117
g2926 and n3114_not n3117 ; n3118
g2927 and asqrt[43] n3096_not ; n3119
g2928 and n3091_not n3119 ; n3120
g2929 and n3087_not n3120 ; n3121
g2930 and n3085_not n3121 ; n3122
g2931 nor n3112 n3122 ; n3123
g2932 and a[86] n3123_not ; n3124
g2933 nor a[86] n3122 ; n3125
g2934 and n3112_not n3125 ; n3126
g2935 nor n3124 n3126 ; n3127
g2936 nor n3118 n3127 ; n3128
g2937 nor n3116 n3128 ; n3129
g2938 and asqrt[45] n3129_not ; n3130
g2939 nor n2844 n2849 ; n3131
g2940 and n2853_not n3131 ; n3132
g2941 and asqrt[42] n3132 ; n3133
g2942 and asqrt[42] n3131 ; n3134
g2943 and n2853 n3134_not ; n3135
g2944 nor n3133 n3135 ; n3136
g2945 nor asqrt[45] n3116 ; n3137
g2946 and n3128_not n3137 ; n3138
g2947 nor n3136 n3138 ; n3139
g2948 nor n3130 n3139 ; n3140
g2949 and asqrt[46] n3140_not ; n3141
g2950 and n2858_not n2867 ; n3142
g2951 and n2856_not n3142 ; n3143
g2952 and asqrt[42] n3143 ; n3144
g2953 nor n2856 n2858 ; n3145
g2954 and asqrt[42] n3145 ; n3146
g2955 nor n2867 n3146 ; n3147
g2956 nor n3144 n3147 ; n3148
g2957 nor asqrt[46] n3130 ; n3149
g2958 and n3139_not n3149 ; n3150
g2959 nor n3148 n3150 ; n3151
g2960 nor n3141 n3151 ; n3152
g2961 and asqrt[47] n3152_not ; n3153
g2962 and n2870_not n2876 ; n3154
g2963 and n2878_not n3154 ; n3155
g2964 and asqrt[42] n3155 ; n3156
g2965 nor n2870 n2878 ; n3157
g2966 and asqrt[42] n3157 ; n3158
g2967 nor n2876 n3158 ; n3159
g2968 nor n3156 n3159 ; n3160
g2969 nor asqrt[47] n3141 ; n3161
g2970 and n3151_not n3161 ; n3162
g2971 nor n3160 n3162 ; n3163
g2972 nor n3153 n3163 ; n3164
g2973 and asqrt[48] n3164_not ; n3165
g2974 and n2888 n2890_not ; n3166
g2975 and n2881_not n3166 ; n3167
g2976 and asqrt[42] n3167 ; n3168
g2977 nor n2881 n2890 ; n3169
g2978 and asqrt[42] n3169 ; n3170
g2979 nor n2888 n3170 ; n3171
g2980 nor n3168 n3171 ; n3172
g2981 nor asqrt[48] n3153 ; n3173
g2982 and n3163_not n3173 ; n3174
g2983 nor n3172 n3174 ; n3175
g2984 nor n3165 n3175 ; n3176
g2985 and asqrt[49] n3176_not ; n3177
g2986 and n2893_not n2900 ; n3178
g2987 and n2902_not n3178 ; n3179
g2988 and asqrt[42] n3179 ; n3180
g2989 nor n2893 n2902 ; n3181
g2990 and asqrt[42] n3181 ; n3182
g2991 nor n2900 n3182 ; n3183
g2992 nor n3180 n3183 ; n3184
g2993 nor asqrt[49] n3165 ; n3185
g2994 and n3175_not n3185 ; n3186
g2995 nor n3184 n3186 ; n3187
g2996 nor n3177 n3187 ; n3188
g2997 and asqrt[50] n3188_not ; n3189
g2998 and n2912 n2914_not ; n3190
g2999 and n2905_not n3190 ; n3191
g3000 and asqrt[42] n3191 ; n3192
g3001 nor n2905 n2914 ; n3193
g3002 and asqrt[42] n3193 ; n3194
g3003 nor n2912 n3194 ; n3195
g3004 nor n3192 n3195 ; n3196
g3005 nor asqrt[50] n3177 ; n3197
g3006 and n3187_not n3197 ; n3198
g3007 nor n3196 n3198 ; n3199
g3008 nor n3189 n3199 ; n3200
g3009 and asqrt[51] n3200_not ; n3201
g3010 and n2917_not n2924 ; n3202
g3011 and n2926_not n3202 ; n3203
g3012 and asqrt[42] n3203 ; n3204
g3013 nor n2917 n2926 ; n3205
g3014 and asqrt[42] n3205 ; n3206
g3015 nor n2924 n3206 ; n3207
g3016 nor n3204 n3207 ; n3208
g3017 nor asqrt[51] n3189 ; n3209
g3018 and n3199_not n3209 ; n3210
g3019 nor n3208 n3210 ; n3211
g3020 nor n3201 n3211 ; n3212
g3021 and asqrt[52] n3212_not ; n3213
g3022 and n2936 n2938_not ; n3214
g3023 and n2929_not n3214 ; n3215
g3024 and asqrt[42] n3215 ; n3216
g3025 nor n2929 n2938 ; n3217
g3026 and asqrt[42] n3217 ; n3218
g3027 nor n2936 n3218 ; n3219
g3028 nor n3216 n3219 ; n3220
g3029 nor asqrt[52] n3201 ; n3221
g3030 and n3211_not n3221 ; n3222
g3031 nor n3220 n3222 ; n3223
g3032 nor n3213 n3223 ; n3224
g3033 and asqrt[53] n3224_not ; n3225
g3034 and n2941_not n2948 ; n3226
g3035 and n2950_not n3226 ; n3227
g3036 and asqrt[42] n3227 ; n3228
g3037 nor n2941 n2950 ; n3229
g3038 and asqrt[42] n3229 ; n3230
g3039 nor n2948 n3230 ; n3231
g3040 nor n3228 n3231 ; n3232
g3041 nor asqrt[53] n3213 ; n3233
g3042 and n3223_not n3233 ; n3234
g3043 nor n3232 n3234 ; n3235
g3044 nor n3225 n3235 ; n3236
g3045 and asqrt[54] n3236_not ; n3237
g3046 and n2960 n2962_not ; n3238
g3047 and n2953_not n3238 ; n3239
g3048 and asqrt[42] n3239 ; n3240
g3049 nor n2953 n2962 ; n3241
g3050 and asqrt[42] n3241 ; n3242
g3051 nor n2960 n3242 ; n3243
g3052 nor n3240 n3243 ; n3244
g3053 nor asqrt[54] n3225 ; n3245
g3054 and n3235_not n3245 ; n3246
g3055 nor n3244 n3246 ; n3247
g3056 nor n3237 n3247 ; n3248
g3057 and asqrt[55] n3248_not ; n3249
g3058 nor asqrt[55] n3237 ; n3250
g3059 and n3247_not n3250 ; n3251
g3060 and n2965_not n2974 ; n3252
g3061 and n2967_not n3252 ; n3253
g3062 and asqrt[42] n3253 ; n3254
g3063 nor n2965 n2967 ; n3255
g3064 and asqrt[42] n3255 ; n3256
g3065 nor n2974 n3256 ; n3257
g3066 nor n3254 n3257 ; n3258
g3067 nor n3251 n3258 ; n3259
g3068 nor n3249 n3259 ; n3260
g3069 and asqrt[56] n3260_not ; n3261
g3070 and n2984 n2986_not ; n3262
g3071 and n2977_not n3262 ; n3263
g3072 and asqrt[42] n3263 ; n3264
g3073 nor n2977 n2986 ; n3265
g3074 and asqrt[42] n3265 ; n3266
g3075 nor n2984 n3266 ; n3267
g3076 nor n3264 n3267 ; n3268
g3077 nor asqrt[56] n3249 ; n3269
g3078 and n3259_not n3269 ; n3270
g3079 nor n3268 n3270 ; n3271
g3080 nor n3261 n3271 ; n3272
g3081 and asqrt[57] n3272_not ; n3273
g3082 and n2989_not n2996 ; n3274
g3083 and n2998_not n3274 ; n3275
g3084 and asqrt[42] n3275 ; n3276
g3085 nor n2989 n2998 ; n3277
g3086 and asqrt[42] n3277 ; n3278
g3087 nor n2996 n3278 ; n3279
g3088 nor n3276 n3279 ; n3280
g3089 nor asqrt[57] n3261 ; n3281
g3090 and n3271_not n3281 ; n3282
g3091 nor n3280 n3282 ; n3283
g3092 nor n3273 n3283 ; n3284
g3093 and asqrt[58] n3284_not ; n3285
g3094 and n3008 n3010_not ; n3286
g3095 and n3001_not n3286 ; n3287
g3096 and asqrt[42] n3287 ; n3288
g3097 nor n3001 n3010 ; n3289
g3098 and asqrt[42] n3289 ; n3290
g3099 nor n3008 n3290 ; n3291
g3100 nor n3288 n3291 ; n3292
g3101 nor asqrt[58] n3273 ; n3293
g3102 and n3283_not n3293 ; n3294
g3103 nor n3292 n3294 ; n3295
g3104 nor n3285 n3295 ; n3296
g3105 and asqrt[59] n3296_not ; n3297
g3106 and n3013_not n3020 ; n3298
g3107 and n3022_not n3298 ; n3299
g3108 and asqrt[42] n3299 ; n3300
g3109 nor n3013 n3022 ; n3301
g3110 and asqrt[42] n3301 ; n3302
g3111 nor n3020 n3302 ; n3303
g3112 nor n3300 n3303 ; n3304
g3113 nor asqrt[59] n3285 ; n3305
g3114 and n3295_not n3305 ; n3306
g3115 nor n3304 n3306 ; n3307
g3116 nor n3297 n3307 ; n3308
g3117 and asqrt[60] n3308_not ; n3309
g3118 and n3032 n3034_not ; n3310
g3119 and n3025_not n3310 ; n3311
g3120 and asqrt[42] n3311 ; n3312
g3121 nor n3025 n3034 ; n3313
g3122 and asqrt[42] n3313 ; n3314
g3123 nor n3032 n3314 ; n3315
g3124 nor n3312 n3315 ; n3316
g3125 nor asqrt[60] n3297 ; n3317
g3126 and n3307_not n3317 ; n3318
g3127 nor n3316 n3318 ; n3319
g3128 nor n3309 n3319 ; n3320
g3129 and asqrt[61] n3320_not ; n3321
g3130 and n3037_not n3044 ; n3322
g3131 and n3046_not n3322 ; n3323
g3132 and asqrt[42] n3323 ; n3324
g3133 nor n3037 n3046 ; n3325
g3134 and asqrt[42] n3325 ; n3326
g3135 nor n3044 n3326 ; n3327
g3136 nor n3324 n3327 ; n3328
g3137 nor asqrt[61] n3309 ; n3329
g3138 and n3319_not n3329 ; n3330
g3139 nor n3328 n3330 ; n3331
g3140 nor n3321 n3331 ; n3332
g3141 and asqrt[62] n3332_not ; n3333
g3142 and n3056 n3058_not ; n3334
g3143 and n3049_not n3334 ; n3335
g3144 and asqrt[42] n3335 ; n3336
g3145 nor n3049 n3058 ; n3337
g3146 and asqrt[42] n3337 ; n3338
g3147 nor n3056 n3338 ; n3339
g3148 nor n3336 n3339 ; n3340
g3149 nor asqrt[62] n3321 ; n3341
g3150 and n3331_not n3341 ; n3342
g3151 nor n3340 n3342 ; n3343
g3152 nor n3333 n3343 ; n3344
g3153 and n3061_not n3068 ; n3345
g3154 and n3070_not n3345 ; n3346
g3155 and asqrt[42] n3346 ; n3347
g3156 nor n3061 n3070 ; n3348
g3157 and asqrt[42] n3348 ; n3349
g3158 nor n3068 n3349 ; n3350
g3159 nor n3347 n3350 ; n3351
g3160 nor n3072 n3079 ; n3352
g3161 and asqrt[42] n3352 ; n3353
g3162 nor n3087 n3353 ; n3354
g3163 and n3351_not n3354 ; n3355
g3164 and n3344_not n3355 ; n3356
g3165 nor asqrt[63] n3356 ; n3357
g3166 and n3333_not n3351 ; n3358
g3167 and n3343_not n3358 ; n3359
g3168 and n3079_not asqrt[42] ; n3360
g3169 and n3072 n3360_not ; n3361
g3170 and asqrt[63] n3352_not ; n3362
g3171 and n3361_not n3362 ; n3363
g3172 nor n3075 n3096 ; n3364
g3173 and n3078_not n3364 ; n3365
g3174 and n3091_not n3365 ; n3366
g3175 and n3087_not n3366 ; n3367
g3176 and n3085_not n3367 ; n3368
g3177 nor n3363 n3368 ; n3369
g3178 and n3359_not n3369 ; n3370
g3179 nand n3357_not n3370 ; asqrt[41]
g3180 and a[82] asqrt[41] ; n3372
g3181 nor a[80] a[81] ; n3373
g3182 and a[82]_not n3373 ; n3374
g3183 nor n3372 n3374 ; n3375
g3184 and asqrt[42] n3375_not ; n3376
g3185 nor n3096 n3374 ; n3377
g3186 and n3091_not n3377 ; n3378
g3187 and n3087_not n3378 ; n3379
g3188 and n3085_not n3379 ; n3380
g3189 and n3372_not n3380 ; n3381
g3190 and a[82]_not asqrt[41] ; n3382
g3191 and a[83] n3382_not ; n3383
g3192 and n3101 asqrt[41] ; n3384
g3193 nor n3383 n3384 ; n3385
g3194 and n3381_not n3385 ; n3386
g3195 nor n3376 n3386 ; n3387
g3196 and asqrt[43] n3387_not ; n3388
g3197 nor asqrt[43] n3376 ; n3389
g3198 and n3386_not n3389 ; n3390
g3199 and asqrt[42] n3368_not ; n3391
g3200 and n3363_not n3391 ; n3392
g3201 and n3359_not n3392 ; n3393
g3202 and n3357_not n3393 ; n3394
g3203 nor n3384 n3394 ; n3395
g3204 and a[84] n3395_not ; n3396
g3205 nor a[84] n3394 ; n3397
g3206 and n3384_not n3397 ; n3398
g3207 nor n3396 n3398 ; n3399
g3208 nor n3390 n3399 ; n3400
g3209 nor n3388 n3400 ; n3401
g3210 and asqrt[44] n3401_not ; n3402
g3211 nor n3104 n3109 ; n3403
g3212 and n3113_not n3403 ; n3404
g3213 and asqrt[41] n3404 ; n3405
g3214 and asqrt[41] n3403 ; n3406
g3215 and n3113 n3406_not ; n3407
g3216 nor n3405 n3407 ; n3408
g3217 nor asqrt[44] n3388 ; n3409
g3218 and n3400_not n3409 ; n3410
g3219 nor n3408 n3410 ; n3411
g3220 nor n3402 n3411 ; n3412
g3221 and asqrt[45] n3412_not ; n3413
g3222 and n3118_not n3127 ; n3414
g3223 and n3116_not n3414 ; n3415
g3224 and asqrt[41] n3415 ; n3416
g3225 nor n3116 n3118 ; n3417
g3226 and asqrt[41] n3417 ; n3418
g3227 nor n3127 n3418 ; n3419
g3228 nor n3416 n3419 ; n3420
g3229 nor asqrt[45] n3402 ; n3421
g3230 and n3411_not n3421 ; n3422
g3231 nor n3420 n3422 ; n3423
g3232 nor n3413 n3423 ; n3424
g3233 and asqrt[46] n3424_not ; n3425
g3234 and n3130_not n3136 ; n3426
g3235 and n3138_not n3426 ; n3427
g3236 and asqrt[41] n3427 ; n3428
g3237 nor n3130 n3138 ; n3429
g3238 and asqrt[41] n3429 ; n3430
g3239 nor n3136 n3430 ; n3431
g3240 nor n3428 n3431 ; n3432
g3241 nor asqrt[46] n3413 ; n3433
g3242 and n3423_not n3433 ; n3434
g3243 nor n3432 n3434 ; n3435
g3244 nor n3425 n3435 ; n3436
g3245 and asqrt[47] n3436_not ; n3437
g3246 and n3148 n3150_not ; n3438
g3247 and n3141_not n3438 ; n3439
g3248 and asqrt[41] n3439 ; n3440
g3249 nor n3141 n3150 ; n3441
g3250 and asqrt[41] n3441 ; n3442
g3251 nor n3148 n3442 ; n3443
g3252 nor n3440 n3443 ; n3444
g3253 nor asqrt[47] n3425 ; n3445
g3254 and n3435_not n3445 ; n3446
g3255 nor n3444 n3446 ; n3447
g3256 nor n3437 n3447 ; n3448
g3257 and asqrt[48] n3448_not ; n3449
g3258 and n3153_not n3160 ; n3450
g3259 and n3162_not n3450 ; n3451
g3260 and asqrt[41] n3451 ; n3452
g3261 nor n3153 n3162 ; n3453
g3262 and asqrt[41] n3453 ; n3454
g3263 nor n3160 n3454 ; n3455
g3264 nor n3452 n3455 ; n3456
g3265 nor asqrt[48] n3437 ; n3457
g3266 and n3447_not n3457 ; n3458
g3267 nor n3456 n3458 ; n3459
g3268 nor n3449 n3459 ; n3460
g3269 and asqrt[49] n3460_not ; n3461
g3270 and n3172 n3174_not ; n3462
g3271 and n3165_not n3462 ; n3463
g3272 and asqrt[41] n3463 ; n3464
g3273 nor n3165 n3174 ; n3465
g3274 and asqrt[41] n3465 ; n3466
g3275 nor n3172 n3466 ; n3467
g3276 nor n3464 n3467 ; n3468
g3277 nor asqrt[49] n3449 ; n3469
g3278 and n3459_not n3469 ; n3470
g3279 nor n3468 n3470 ; n3471
g3280 nor n3461 n3471 ; n3472
g3281 and asqrt[50] n3472_not ; n3473
g3282 and n3177_not n3184 ; n3474
g3283 and n3186_not n3474 ; n3475
g3284 and asqrt[41] n3475 ; n3476
g3285 nor n3177 n3186 ; n3477
g3286 and asqrt[41] n3477 ; n3478
g3287 nor n3184 n3478 ; n3479
g3288 nor n3476 n3479 ; n3480
g3289 nor asqrt[50] n3461 ; n3481
g3290 and n3471_not n3481 ; n3482
g3291 nor n3480 n3482 ; n3483
g3292 nor n3473 n3483 ; n3484
g3293 and asqrt[51] n3484_not ; n3485
g3294 and n3196 n3198_not ; n3486
g3295 and n3189_not n3486 ; n3487
g3296 and asqrt[41] n3487 ; n3488
g3297 nor n3189 n3198 ; n3489
g3298 and asqrt[41] n3489 ; n3490
g3299 nor n3196 n3490 ; n3491
g3300 nor n3488 n3491 ; n3492
g3301 nor asqrt[51] n3473 ; n3493
g3302 and n3483_not n3493 ; n3494
g3303 nor n3492 n3494 ; n3495
g3304 nor n3485 n3495 ; n3496
g3305 and asqrt[52] n3496_not ; n3497
g3306 and n3201_not n3208 ; n3498
g3307 and n3210_not n3498 ; n3499
g3308 and asqrt[41] n3499 ; n3500
g3309 nor n3201 n3210 ; n3501
g3310 and asqrt[41] n3501 ; n3502
g3311 nor n3208 n3502 ; n3503
g3312 nor n3500 n3503 ; n3504
g3313 nor asqrt[52] n3485 ; n3505
g3314 and n3495_not n3505 ; n3506
g3315 nor n3504 n3506 ; n3507
g3316 nor n3497 n3507 ; n3508
g3317 and asqrt[53] n3508_not ; n3509
g3318 and n3220 n3222_not ; n3510
g3319 and n3213_not n3510 ; n3511
g3320 and asqrt[41] n3511 ; n3512
g3321 nor n3213 n3222 ; n3513
g3322 and asqrt[41] n3513 ; n3514
g3323 nor n3220 n3514 ; n3515
g3324 nor n3512 n3515 ; n3516
g3325 nor asqrt[53] n3497 ; n3517
g3326 and n3507_not n3517 ; n3518
g3327 nor n3516 n3518 ; n3519
g3328 nor n3509 n3519 ; n3520
g3329 and asqrt[54] n3520_not ; n3521
g3330 and n3225_not n3232 ; n3522
g3331 and n3234_not n3522 ; n3523
g3332 and asqrt[41] n3523 ; n3524
g3333 nor n3225 n3234 ; n3525
g3334 and asqrt[41] n3525 ; n3526
g3335 nor n3232 n3526 ; n3527
g3336 nor n3524 n3527 ; n3528
g3337 nor asqrt[54] n3509 ; n3529
g3338 and n3519_not n3529 ; n3530
g3339 nor n3528 n3530 ; n3531
g3340 nor n3521 n3531 ; n3532
g3341 and asqrt[55] n3532_not ; n3533
g3342 and n3244 n3246_not ; n3534
g3343 and n3237_not n3534 ; n3535
g3344 and asqrt[41] n3535 ; n3536
g3345 nor n3237 n3246 ; n3537
g3346 and asqrt[41] n3537 ; n3538
g3347 nor n3244 n3538 ; n3539
g3348 nor n3536 n3539 ; n3540
g3349 nor asqrt[55] n3521 ; n3541
g3350 and n3531_not n3541 ; n3542
g3351 nor n3540 n3542 ; n3543
g3352 nor n3533 n3543 ; n3544
g3353 and asqrt[56] n3544_not ; n3545
g3354 nor asqrt[56] n3533 ; n3546
g3355 and n3543_not n3546 ; n3547
g3356 and n3249_not n3258 ; n3548
g3357 and n3251_not n3548 ; n3549
g3358 and asqrt[41] n3549 ; n3550
g3359 nor n3249 n3251 ; n3551
g3360 and asqrt[41] n3551 ; n3552
g3361 nor n3258 n3552 ; n3553
g3362 nor n3550 n3553 ; n3554
g3363 nor n3547 n3554 ; n3555
g3364 nor n3545 n3555 ; n3556
g3365 and asqrt[57] n3556_not ; n3557
g3366 and n3268 n3270_not ; n3558
g3367 and n3261_not n3558 ; n3559
g3368 and asqrt[41] n3559 ; n3560
g3369 nor n3261 n3270 ; n3561
g3370 and asqrt[41] n3561 ; n3562
g3371 nor n3268 n3562 ; n3563
g3372 nor n3560 n3563 ; n3564
g3373 nor asqrt[57] n3545 ; n3565
g3374 and n3555_not n3565 ; n3566
g3375 nor n3564 n3566 ; n3567
g3376 nor n3557 n3567 ; n3568
g3377 and asqrt[58] n3568_not ; n3569
g3378 and n3273_not n3280 ; n3570
g3379 and n3282_not n3570 ; n3571
g3380 and asqrt[41] n3571 ; n3572
g3381 nor n3273 n3282 ; n3573
g3382 and asqrt[41] n3573 ; n3574
g3383 nor n3280 n3574 ; n3575
g3384 nor n3572 n3575 ; n3576
g3385 nor asqrt[58] n3557 ; n3577
g3386 and n3567_not n3577 ; n3578
g3387 nor n3576 n3578 ; n3579
g3388 nor n3569 n3579 ; n3580
g3389 and asqrt[59] n3580_not ; n3581
g3390 and n3292 n3294_not ; n3582
g3391 and n3285_not n3582 ; n3583
g3392 and asqrt[41] n3583 ; n3584
g3393 nor n3285 n3294 ; n3585
g3394 and asqrt[41] n3585 ; n3586
g3395 nor n3292 n3586 ; n3587
g3396 nor n3584 n3587 ; n3588
g3397 nor asqrt[59] n3569 ; n3589
g3398 and n3579_not n3589 ; n3590
g3399 nor n3588 n3590 ; n3591
g3400 nor n3581 n3591 ; n3592
g3401 and asqrt[60] n3592_not ; n3593
g3402 and n3297_not n3304 ; n3594
g3403 and n3306_not n3594 ; n3595
g3404 and asqrt[41] n3595 ; n3596
g3405 nor n3297 n3306 ; n3597
g3406 and asqrt[41] n3597 ; n3598
g3407 nor n3304 n3598 ; n3599
g3408 nor n3596 n3599 ; n3600
g3409 nor asqrt[60] n3581 ; n3601
g3410 and n3591_not n3601 ; n3602
g3411 nor n3600 n3602 ; n3603
g3412 nor n3593 n3603 ; n3604
g3413 and asqrt[61] n3604_not ; n3605
g3414 and n3316 n3318_not ; n3606
g3415 and n3309_not n3606 ; n3607
g3416 and asqrt[41] n3607 ; n3608
g3417 nor n3309 n3318 ; n3609
g3418 and asqrt[41] n3609 ; n3610
g3419 nor n3316 n3610 ; n3611
g3420 nor n3608 n3611 ; n3612
g3421 nor asqrt[61] n3593 ; n3613
g3422 and n3603_not n3613 ; n3614
g3423 nor n3612 n3614 ; n3615
g3424 nor n3605 n3615 ; n3616
g3425 and asqrt[62] n3616_not ; n3617
g3426 and n3321_not n3328 ; n3618
g3427 and n3330_not n3618 ; n3619
g3428 and asqrt[41] n3619 ; n3620
g3429 nor n3321 n3330 ; n3621
g3430 and asqrt[41] n3621 ; n3622
g3431 nor n3328 n3622 ; n3623
g3432 nor n3620 n3623 ; n3624
g3433 nor asqrt[62] n3605 ; n3625
g3434 and n3615_not n3625 ; n3626
g3435 nor n3624 n3626 ; n3627
g3436 nor n3617 n3627 ; n3628
g3437 and n3340 n3342_not ; n3629
g3438 and n3333_not n3629 ; n3630
g3439 and asqrt[41] n3630 ; n3631
g3440 nor n3333 n3342 ; n3632
g3441 and asqrt[41] n3632 ; n3633
g3442 nor n3340 n3633 ; n3634
g3443 nor n3631 n3634 ; n3635
g3444 nor n3344 n3351 ; n3636
g3445 and asqrt[41] n3636 ; n3637
g3446 nor n3359 n3637 ; n3638
g3447 and n3635_not n3638 ; n3639
g3448 and n3628_not n3639 ; n3640
g3449 nor asqrt[63] n3640 ; n3641
g3450 and n3617_not n3635 ; n3642
g3451 and n3627_not n3642 ; n3643
g3452 and n3351_not asqrt[41] ; n3644
g3453 and n3344 n3644_not ; n3645
g3454 and asqrt[63] n3636_not ; n3646
g3455 and n3645_not n3646 ; n3647
g3456 nor n3347 n3368 ; n3648
g3457 and n3350_not n3648 ; n3649
g3458 and n3363_not n3649 ; n3650
g3459 and n3359_not n3650 ; n3651
g3460 and n3357_not n3651 ; n3652
g3461 nor n3647 n3652 ; n3653
g3462 and n3643_not n3653 ; n3654
g3463 nand n3641_not n3654 ; asqrt[40]
g3464 and a[80] asqrt[40] ; n3656
g3465 nor a[78] a[79] ; n3657
g3466 and a[80]_not n3657 ; n3658
g3467 nor n3656 n3658 ; n3659
g3468 and asqrt[41] n3659_not ; n3660
g3469 nor n3368 n3658 ; n3661
g3470 and n3363_not n3661 ; n3662
g3471 and n3359_not n3662 ; n3663
g3472 and n3357_not n3663 ; n3664
g3473 and n3656_not n3664 ; n3665
g3474 and a[80]_not asqrt[40] ; n3666
g3475 and a[81] n3666_not ; n3667
g3476 and n3373 asqrt[40] ; n3668
g3477 nor n3667 n3668 ; n3669
g3478 and n3665_not n3669 ; n3670
g3479 nor n3660 n3670 ; n3671
g3480 and asqrt[42] n3671_not ; n3672
g3481 nor asqrt[42] n3660 ; n3673
g3482 and n3670_not n3673 ; n3674
g3483 and asqrt[41] n3652_not ; n3675
g3484 and n3647_not n3675 ; n3676
g3485 and n3643_not n3676 ; n3677
g3486 and n3641_not n3677 ; n3678
g3487 nor n3668 n3678 ; n3679
g3488 and a[82] n3679_not ; n3680
g3489 nor a[82] n3678 ; n3681
g3490 and n3668_not n3681 ; n3682
g3491 nor n3680 n3682 ; n3683
g3492 nor n3674 n3683 ; n3684
g3493 nor n3672 n3684 ; n3685
g3494 and asqrt[43] n3685_not ; n3686
g3495 nor n3376 n3381 ; n3687
g3496 and n3385_not n3687 ; n3688
g3497 and asqrt[40] n3688 ; n3689
g3498 and asqrt[40] n3687 ; n3690
g3499 and n3385 n3690_not ; n3691
g3500 nor n3689 n3691 ; n3692
g3501 nor asqrt[43] n3672 ; n3693
g3502 and n3684_not n3693 ; n3694
g3503 nor n3692 n3694 ; n3695
g3504 nor n3686 n3695 ; n3696
g3505 and asqrt[44] n3696_not ; n3697
g3506 and n3390_not n3399 ; n3698
g3507 and n3388_not n3698 ; n3699
g3508 and asqrt[40] n3699 ; n3700
g3509 nor n3388 n3390 ; n3701
g3510 and asqrt[40] n3701 ; n3702
g3511 nor n3399 n3702 ; n3703
g3512 nor n3700 n3703 ; n3704
g3513 nor asqrt[44] n3686 ; n3705
g3514 and n3695_not n3705 ; n3706
g3515 nor n3704 n3706 ; n3707
g3516 nor n3697 n3707 ; n3708
g3517 and asqrt[45] n3708_not ; n3709
g3518 and n3402_not n3408 ; n3710
g3519 and n3410_not n3710 ; n3711
g3520 and asqrt[40] n3711 ; n3712
g3521 nor n3402 n3410 ; n3713
g3522 and asqrt[40] n3713 ; n3714
g3523 nor n3408 n3714 ; n3715
g3524 nor n3712 n3715 ; n3716
g3525 nor asqrt[45] n3697 ; n3717
g3526 and n3707_not n3717 ; n3718
g3527 nor n3716 n3718 ; n3719
g3528 nor n3709 n3719 ; n3720
g3529 and asqrt[46] n3720_not ; n3721
g3530 and n3420 n3422_not ; n3722
g3531 and n3413_not n3722 ; n3723
g3532 and asqrt[40] n3723 ; n3724
g3533 nor n3413 n3422 ; n3725
g3534 and asqrt[40] n3725 ; n3726
g3535 nor n3420 n3726 ; n3727
g3536 nor n3724 n3727 ; n3728
g3537 nor asqrt[46] n3709 ; n3729
g3538 and n3719_not n3729 ; n3730
g3539 nor n3728 n3730 ; n3731
g3540 nor n3721 n3731 ; n3732
g3541 and asqrt[47] n3732_not ; n3733
g3542 and n3425_not n3432 ; n3734
g3543 and n3434_not n3734 ; n3735
g3544 and asqrt[40] n3735 ; n3736
g3545 nor n3425 n3434 ; n3737
g3546 and asqrt[40] n3737 ; n3738
g3547 nor n3432 n3738 ; n3739
g3548 nor n3736 n3739 ; n3740
g3549 nor asqrt[47] n3721 ; n3741
g3550 and n3731_not n3741 ; n3742
g3551 nor n3740 n3742 ; n3743
g3552 nor n3733 n3743 ; n3744
g3553 and asqrt[48] n3744_not ; n3745
g3554 and n3444 n3446_not ; n3746
g3555 and n3437_not n3746 ; n3747
g3556 and asqrt[40] n3747 ; n3748
g3557 nor n3437 n3446 ; n3749
g3558 and asqrt[40] n3749 ; n3750
g3559 nor n3444 n3750 ; n3751
g3560 nor n3748 n3751 ; n3752
g3561 nor asqrt[48] n3733 ; n3753
g3562 and n3743_not n3753 ; n3754
g3563 nor n3752 n3754 ; n3755
g3564 nor n3745 n3755 ; n3756
g3565 and asqrt[49] n3756_not ; n3757
g3566 and n3449_not n3456 ; n3758
g3567 and n3458_not n3758 ; n3759
g3568 and asqrt[40] n3759 ; n3760
g3569 nor n3449 n3458 ; n3761
g3570 and asqrt[40] n3761 ; n3762
g3571 nor n3456 n3762 ; n3763
g3572 nor n3760 n3763 ; n3764
g3573 nor asqrt[49] n3745 ; n3765
g3574 and n3755_not n3765 ; n3766
g3575 nor n3764 n3766 ; n3767
g3576 nor n3757 n3767 ; n3768
g3577 and asqrt[50] n3768_not ; n3769
g3578 and n3468 n3470_not ; n3770
g3579 and n3461_not n3770 ; n3771
g3580 and asqrt[40] n3771 ; n3772
g3581 nor n3461 n3470 ; n3773
g3582 and asqrt[40] n3773 ; n3774
g3583 nor n3468 n3774 ; n3775
g3584 nor n3772 n3775 ; n3776
g3585 nor asqrt[50] n3757 ; n3777
g3586 and n3767_not n3777 ; n3778
g3587 nor n3776 n3778 ; n3779
g3588 nor n3769 n3779 ; n3780
g3589 and asqrt[51] n3780_not ; n3781
g3590 and n3473_not n3480 ; n3782
g3591 and n3482_not n3782 ; n3783
g3592 and asqrt[40] n3783 ; n3784
g3593 nor n3473 n3482 ; n3785
g3594 and asqrt[40] n3785 ; n3786
g3595 nor n3480 n3786 ; n3787
g3596 nor n3784 n3787 ; n3788
g3597 nor asqrt[51] n3769 ; n3789
g3598 and n3779_not n3789 ; n3790
g3599 nor n3788 n3790 ; n3791
g3600 nor n3781 n3791 ; n3792
g3601 and asqrt[52] n3792_not ; n3793
g3602 and n3492 n3494_not ; n3794
g3603 and n3485_not n3794 ; n3795
g3604 and asqrt[40] n3795 ; n3796
g3605 nor n3485 n3494 ; n3797
g3606 and asqrt[40] n3797 ; n3798
g3607 nor n3492 n3798 ; n3799
g3608 nor n3796 n3799 ; n3800
g3609 nor asqrt[52] n3781 ; n3801
g3610 and n3791_not n3801 ; n3802
g3611 nor n3800 n3802 ; n3803
g3612 nor n3793 n3803 ; n3804
g3613 and asqrt[53] n3804_not ; n3805
g3614 and n3497_not n3504 ; n3806
g3615 and n3506_not n3806 ; n3807
g3616 and asqrt[40] n3807 ; n3808
g3617 nor n3497 n3506 ; n3809
g3618 and asqrt[40] n3809 ; n3810
g3619 nor n3504 n3810 ; n3811
g3620 nor n3808 n3811 ; n3812
g3621 nor asqrt[53] n3793 ; n3813
g3622 and n3803_not n3813 ; n3814
g3623 nor n3812 n3814 ; n3815
g3624 nor n3805 n3815 ; n3816
g3625 and asqrt[54] n3816_not ; n3817
g3626 and n3516 n3518_not ; n3818
g3627 and n3509_not n3818 ; n3819
g3628 and asqrt[40] n3819 ; n3820
g3629 nor n3509 n3518 ; n3821
g3630 and asqrt[40] n3821 ; n3822
g3631 nor n3516 n3822 ; n3823
g3632 nor n3820 n3823 ; n3824
g3633 nor asqrt[54] n3805 ; n3825
g3634 and n3815_not n3825 ; n3826
g3635 nor n3824 n3826 ; n3827
g3636 nor n3817 n3827 ; n3828
g3637 and asqrt[55] n3828_not ; n3829
g3638 and n3521_not n3528 ; n3830
g3639 and n3530_not n3830 ; n3831
g3640 and asqrt[40] n3831 ; n3832
g3641 nor n3521 n3530 ; n3833
g3642 and asqrt[40] n3833 ; n3834
g3643 nor n3528 n3834 ; n3835
g3644 nor n3832 n3835 ; n3836
g3645 nor asqrt[55] n3817 ; n3837
g3646 and n3827_not n3837 ; n3838
g3647 nor n3836 n3838 ; n3839
g3648 nor n3829 n3839 ; n3840
g3649 and asqrt[56] n3840_not ; n3841
g3650 and n3540 n3542_not ; n3842
g3651 and n3533_not n3842 ; n3843
g3652 and asqrt[40] n3843 ; n3844
g3653 nor n3533 n3542 ; n3845
g3654 and asqrt[40] n3845 ; n3846
g3655 nor n3540 n3846 ; n3847
g3656 nor n3844 n3847 ; n3848
g3657 nor asqrt[56] n3829 ; n3849
g3658 and n3839_not n3849 ; n3850
g3659 nor n3848 n3850 ; n3851
g3660 nor n3841 n3851 ; n3852
g3661 and asqrt[57] n3852_not ; n3853
g3662 nor asqrt[57] n3841 ; n3854
g3663 and n3851_not n3854 ; n3855
g3664 and n3545_not n3554 ; n3856
g3665 and n3547_not n3856 ; n3857
g3666 and asqrt[40] n3857 ; n3858
g3667 nor n3545 n3547 ; n3859
g3668 and asqrt[40] n3859 ; n3860
g3669 nor n3554 n3860 ; n3861
g3670 nor n3858 n3861 ; n3862
g3671 nor n3855 n3862 ; n3863
g3672 nor n3853 n3863 ; n3864
g3673 and asqrt[58] n3864_not ; n3865
g3674 and n3564 n3566_not ; n3866
g3675 and n3557_not n3866 ; n3867
g3676 and asqrt[40] n3867 ; n3868
g3677 nor n3557 n3566 ; n3869
g3678 and asqrt[40] n3869 ; n3870
g3679 nor n3564 n3870 ; n3871
g3680 nor n3868 n3871 ; n3872
g3681 nor asqrt[58] n3853 ; n3873
g3682 and n3863_not n3873 ; n3874
g3683 nor n3872 n3874 ; n3875
g3684 nor n3865 n3875 ; n3876
g3685 and asqrt[59] n3876_not ; n3877
g3686 and n3569_not n3576 ; n3878
g3687 and n3578_not n3878 ; n3879
g3688 and asqrt[40] n3879 ; n3880
g3689 nor n3569 n3578 ; n3881
g3690 and asqrt[40] n3881 ; n3882
g3691 nor n3576 n3882 ; n3883
g3692 nor n3880 n3883 ; n3884
g3693 nor asqrt[59] n3865 ; n3885
g3694 and n3875_not n3885 ; n3886
g3695 nor n3884 n3886 ; n3887
g3696 nor n3877 n3887 ; n3888
g3697 and asqrt[60] n3888_not ; n3889
g3698 and n3588 n3590_not ; n3890
g3699 and n3581_not n3890 ; n3891
g3700 and asqrt[40] n3891 ; n3892
g3701 nor n3581 n3590 ; n3893
g3702 and asqrt[40] n3893 ; n3894
g3703 nor n3588 n3894 ; n3895
g3704 nor n3892 n3895 ; n3896
g3705 nor asqrt[60] n3877 ; n3897
g3706 and n3887_not n3897 ; n3898
g3707 nor n3896 n3898 ; n3899
g3708 nor n3889 n3899 ; n3900
g3709 and asqrt[61] n3900_not ; n3901
g3710 and n3593_not n3600 ; n3902
g3711 and n3602_not n3902 ; n3903
g3712 and asqrt[40] n3903 ; n3904
g3713 nor n3593 n3602 ; n3905
g3714 and asqrt[40] n3905 ; n3906
g3715 nor n3600 n3906 ; n3907
g3716 nor n3904 n3907 ; n3908
g3717 nor asqrt[61] n3889 ; n3909
g3718 and n3899_not n3909 ; n3910
g3719 nor n3908 n3910 ; n3911
g3720 nor n3901 n3911 ; n3912
g3721 and asqrt[62] n3912_not ; n3913
g3722 and n3612 n3614_not ; n3914
g3723 and n3605_not n3914 ; n3915
g3724 and asqrt[40] n3915 ; n3916
g3725 nor n3605 n3614 ; n3917
g3726 and asqrt[40] n3917 ; n3918
g3727 nor n3612 n3918 ; n3919
g3728 nor n3916 n3919 ; n3920
g3729 nor asqrt[62] n3901 ; n3921
g3730 and n3911_not n3921 ; n3922
g3731 nor n3920 n3922 ; n3923
g3732 nor n3913 n3923 ; n3924
g3733 and n3617_not n3624 ; n3925
g3734 and n3626_not n3925 ; n3926
g3735 and asqrt[40] n3926 ; n3927
g3736 nor n3617 n3626 ; n3928
g3737 and asqrt[40] n3928 ; n3929
g3738 nor n3624 n3929 ; n3930
g3739 nor n3927 n3930 ; n3931
g3740 nor n3628 n3635 ; n3932
g3741 and asqrt[40] n3932 ; n3933
g3742 nor n3643 n3933 ; n3934
g3743 and n3931_not n3934 ; n3935
g3744 and n3924_not n3935 ; n3936
g3745 nor asqrt[63] n3936 ; n3937
g3746 and n3913_not n3931 ; n3938
g3747 and n3923_not n3938 ; n3939
g3748 and n3635_not asqrt[40] ; n3940
g3749 and n3628 n3940_not ; n3941
g3750 and asqrt[63] n3932_not ; n3942
g3751 and n3941_not n3942 ; n3943
g3752 nor n3631 n3652 ; n3944
g3753 and n3634_not n3944 ; n3945
g3754 and n3647_not n3945 ; n3946
g3755 and n3643_not n3946 ; n3947
g3756 and n3641_not n3947 ; n3948
g3757 nor n3943 n3948 ; n3949
g3758 and n3939_not n3949 ; n3950
g3759 nand n3937_not n3950 ; asqrt[39]
g3760 and a[78] asqrt[39] ; n3952
g3761 nor a[76] a[77] ; n3953
g3762 and a[78]_not n3953 ; n3954
g3763 nor n3952 n3954 ; n3955
g3764 and asqrt[40] n3955_not ; n3956
g3765 nor n3652 n3954 ; n3957
g3766 and n3647_not n3957 ; n3958
g3767 and n3643_not n3958 ; n3959
g3768 and n3641_not n3959 ; n3960
g3769 and n3952_not n3960 ; n3961
g3770 and a[78]_not asqrt[39] ; n3962
g3771 and a[79] n3962_not ; n3963
g3772 and n3657 asqrt[39] ; n3964
g3773 nor n3963 n3964 ; n3965
g3774 and n3961_not n3965 ; n3966
g3775 nor n3956 n3966 ; n3967
g3776 and asqrt[41] n3967_not ; n3968
g3777 nor asqrt[41] n3956 ; n3969
g3778 and n3966_not n3969 ; n3970
g3779 and asqrt[40] n3948_not ; n3971
g3780 and n3943_not n3971 ; n3972
g3781 and n3939_not n3972 ; n3973
g3782 and n3937_not n3973 ; n3974
g3783 nor n3964 n3974 ; n3975
g3784 and a[80] n3975_not ; n3976
g3785 nor a[80] n3974 ; n3977
g3786 and n3964_not n3977 ; n3978
g3787 nor n3976 n3978 ; n3979
g3788 nor n3970 n3979 ; n3980
g3789 nor n3968 n3980 ; n3981
g3790 and asqrt[42] n3981_not ; n3982
g3791 nor n3660 n3665 ; n3983
g3792 and n3669_not n3983 ; n3984
g3793 and asqrt[39] n3984 ; n3985
g3794 and asqrt[39] n3983 ; n3986
g3795 and n3669 n3986_not ; n3987
g3796 nor n3985 n3987 ; n3988
g3797 nor asqrt[42] n3968 ; n3989
g3798 and n3980_not n3989 ; n3990
g3799 nor n3988 n3990 ; n3991
g3800 nor n3982 n3991 ; n3992
g3801 and asqrt[43] n3992_not ; n3993
g3802 and n3674_not n3683 ; n3994
g3803 and n3672_not n3994 ; n3995
g3804 and asqrt[39] n3995 ; n3996
g3805 nor n3672 n3674 ; n3997
g3806 and asqrt[39] n3997 ; n3998
g3807 nor n3683 n3998 ; n3999
g3808 nor n3996 n3999 ; n4000
g3809 nor asqrt[43] n3982 ; n4001
g3810 and n3991_not n4001 ; n4002
g3811 nor n4000 n4002 ; n4003
g3812 nor n3993 n4003 ; n4004
g3813 and asqrt[44] n4004_not ; n4005
g3814 and n3686_not n3692 ; n4006
g3815 and n3694_not n4006 ; n4007
g3816 and asqrt[39] n4007 ; n4008
g3817 nor n3686 n3694 ; n4009
g3818 and asqrt[39] n4009 ; n4010
g3819 nor n3692 n4010 ; n4011
g3820 nor n4008 n4011 ; n4012
g3821 nor asqrt[44] n3993 ; n4013
g3822 and n4003_not n4013 ; n4014
g3823 nor n4012 n4014 ; n4015
g3824 nor n4005 n4015 ; n4016
g3825 and asqrt[45] n4016_not ; n4017
g3826 and n3704 n3706_not ; n4018
g3827 and n3697_not n4018 ; n4019
g3828 and asqrt[39] n4019 ; n4020
g3829 nor n3697 n3706 ; n4021
g3830 and asqrt[39] n4021 ; n4022
g3831 nor n3704 n4022 ; n4023
g3832 nor n4020 n4023 ; n4024
g3833 nor asqrt[45] n4005 ; n4025
g3834 and n4015_not n4025 ; n4026
g3835 nor n4024 n4026 ; n4027
g3836 nor n4017 n4027 ; n4028
g3837 and asqrt[46] n4028_not ; n4029
g3838 and n3709_not n3716 ; n4030
g3839 and n3718_not n4030 ; n4031
g3840 and asqrt[39] n4031 ; n4032
g3841 nor n3709 n3718 ; n4033
g3842 and asqrt[39] n4033 ; n4034
g3843 nor n3716 n4034 ; n4035
g3844 nor n4032 n4035 ; n4036
g3845 nor asqrt[46] n4017 ; n4037
g3846 and n4027_not n4037 ; n4038
g3847 nor n4036 n4038 ; n4039
g3848 nor n4029 n4039 ; n4040
g3849 and asqrt[47] n4040_not ; n4041
g3850 and n3728 n3730_not ; n4042
g3851 and n3721_not n4042 ; n4043
g3852 and asqrt[39] n4043 ; n4044
g3853 nor n3721 n3730 ; n4045
g3854 and asqrt[39] n4045 ; n4046
g3855 nor n3728 n4046 ; n4047
g3856 nor n4044 n4047 ; n4048
g3857 nor asqrt[47] n4029 ; n4049
g3858 and n4039_not n4049 ; n4050
g3859 nor n4048 n4050 ; n4051
g3860 nor n4041 n4051 ; n4052
g3861 and asqrt[48] n4052_not ; n4053
g3862 and n3733_not n3740 ; n4054
g3863 and n3742_not n4054 ; n4055
g3864 and asqrt[39] n4055 ; n4056
g3865 nor n3733 n3742 ; n4057
g3866 and asqrt[39] n4057 ; n4058
g3867 nor n3740 n4058 ; n4059
g3868 nor n4056 n4059 ; n4060
g3869 nor asqrt[48] n4041 ; n4061
g3870 and n4051_not n4061 ; n4062
g3871 nor n4060 n4062 ; n4063
g3872 nor n4053 n4063 ; n4064
g3873 and asqrt[49] n4064_not ; n4065
g3874 and n3752 n3754_not ; n4066
g3875 and n3745_not n4066 ; n4067
g3876 and asqrt[39] n4067 ; n4068
g3877 nor n3745 n3754 ; n4069
g3878 and asqrt[39] n4069 ; n4070
g3879 nor n3752 n4070 ; n4071
g3880 nor n4068 n4071 ; n4072
g3881 nor asqrt[49] n4053 ; n4073
g3882 and n4063_not n4073 ; n4074
g3883 nor n4072 n4074 ; n4075
g3884 nor n4065 n4075 ; n4076
g3885 and asqrt[50] n4076_not ; n4077
g3886 and n3757_not n3764 ; n4078
g3887 and n3766_not n4078 ; n4079
g3888 and asqrt[39] n4079 ; n4080
g3889 nor n3757 n3766 ; n4081
g3890 and asqrt[39] n4081 ; n4082
g3891 nor n3764 n4082 ; n4083
g3892 nor n4080 n4083 ; n4084
g3893 nor asqrt[50] n4065 ; n4085
g3894 and n4075_not n4085 ; n4086
g3895 nor n4084 n4086 ; n4087
g3896 nor n4077 n4087 ; n4088
g3897 and asqrt[51] n4088_not ; n4089
g3898 and n3776 n3778_not ; n4090
g3899 and n3769_not n4090 ; n4091
g3900 and asqrt[39] n4091 ; n4092
g3901 nor n3769 n3778 ; n4093
g3902 and asqrt[39] n4093 ; n4094
g3903 nor n3776 n4094 ; n4095
g3904 nor n4092 n4095 ; n4096
g3905 nor asqrt[51] n4077 ; n4097
g3906 and n4087_not n4097 ; n4098
g3907 nor n4096 n4098 ; n4099
g3908 nor n4089 n4099 ; n4100
g3909 and asqrt[52] n4100_not ; n4101
g3910 and n3781_not n3788 ; n4102
g3911 and n3790_not n4102 ; n4103
g3912 and asqrt[39] n4103 ; n4104
g3913 nor n3781 n3790 ; n4105
g3914 and asqrt[39] n4105 ; n4106
g3915 nor n3788 n4106 ; n4107
g3916 nor n4104 n4107 ; n4108
g3917 nor asqrt[52] n4089 ; n4109
g3918 and n4099_not n4109 ; n4110
g3919 nor n4108 n4110 ; n4111
g3920 nor n4101 n4111 ; n4112
g3921 and asqrt[53] n4112_not ; n4113
g3922 and n3800 n3802_not ; n4114
g3923 and n3793_not n4114 ; n4115
g3924 and asqrt[39] n4115 ; n4116
g3925 nor n3793 n3802 ; n4117
g3926 and asqrt[39] n4117 ; n4118
g3927 nor n3800 n4118 ; n4119
g3928 nor n4116 n4119 ; n4120
g3929 nor asqrt[53] n4101 ; n4121
g3930 and n4111_not n4121 ; n4122
g3931 nor n4120 n4122 ; n4123
g3932 nor n4113 n4123 ; n4124
g3933 and asqrt[54] n4124_not ; n4125
g3934 and n3805_not n3812 ; n4126
g3935 and n3814_not n4126 ; n4127
g3936 and asqrt[39] n4127 ; n4128
g3937 nor n3805 n3814 ; n4129
g3938 and asqrt[39] n4129 ; n4130
g3939 nor n3812 n4130 ; n4131
g3940 nor n4128 n4131 ; n4132
g3941 nor asqrt[54] n4113 ; n4133
g3942 and n4123_not n4133 ; n4134
g3943 nor n4132 n4134 ; n4135
g3944 nor n4125 n4135 ; n4136
g3945 and asqrt[55] n4136_not ; n4137
g3946 and n3824 n3826_not ; n4138
g3947 and n3817_not n4138 ; n4139
g3948 and asqrt[39] n4139 ; n4140
g3949 nor n3817 n3826 ; n4141
g3950 and asqrt[39] n4141 ; n4142
g3951 nor n3824 n4142 ; n4143
g3952 nor n4140 n4143 ; n4144
g3953 nor asqrt[55] n4125 ; n4145
g3954 and n4135_not n4145 ; n4146
g3955 nor n4144 n4146 ; n4147
g3956 nor n4137 n4147 ; n4148
g3957 and asqrt[56] n4148_not ; n4149
g3958 and n3829_not n3836 ; n4150
g3959 and n3838_not n4150 ; n4151
g3960 and asqrt[39] n4151 ; n4152
g3961 nor n3829 n3838 ; n4153
g3962 and asqrt[39] n4153 ; n4154
g3963 nor n3836 n4154 ; n4155
g3964 nor n4152 n4155 ; n4156
g3965 nor asqrt[56] n4137 ; n4157
g3966 and n4147_not n4157 ; n4158
g3967 nor n4156 n4158 ; n4159
g3968 nor n4149 n4159 ; n4160
g3969 and asqrt[57] n4160_not ; n4161
g3970 and n3848 n3850_not ; n4162
g3971 and n3841_not n4162 ; n4163
g3972 and asqrt[39] n4163 ; n4164
g3973 nor n3841 n3850 ; n4165
g3974 and asqrt[39] n4165 ; n4166
g3975 nor n3848 n4166 ; n4167
g3976 nor n4164 n4167 ; n4168
g3977 nor asqrt[57] n4149 ; n4169
g3978 and n4159_not n4169 ; n4170
g3979 nor n4168 n4170 ; n4171
g3980 nor n4161 n4171 ; n4172
g3981 and asqrt[58] n4172_not ; n4173
g3982 nor asqrt[58] n4161 ; n4174
g3983 and n4171_not n4174 ; n4175
g3984 and n3853_not n3862 ; n4176
g3985 and n3855_not n4176 ; n4177
g3986 and asqrt[39] n4177 ; n4178
g3987 nor n3853 n3855 ; n4179
g3988 and asqrt[39] n4179 ; n4180
g3989 nor n3862 n4180 ; n4181
g3990 nor n4178 n4181 ; n4182
g3991 nor n4175 n4182 ; n4183
g3992 nor n4173 n4183 ; n4184
g3993 and asqrt[59] n4184_not ; n4185
g3994 and n3872 n3874_not ; n4186
g3995 and n3865_not n4186 ; n4187
g3996 and asqrt[39] n4187 ; n4188
g3997 nor n3865 n3874 ; n4189
g3998 and asqrt[39] n4189 ; n4190
g3999 nor n3872 n4190 ; n4191
g4000 nor n4188 n4191 ; n4192
g4001 nor asqrt[59] n4173 ; n4193
g4002 and n4183_not n4193 ; n4194
g4003 nor n4192 n4194 ; n4195
g4004 nor n4185 n4195 ; n4196
g4005 and asqrt[60] n4196_not ; n4197
g4006 and n3877_not n3884 ; n4198
g4007 and n3886_not n4198 ; n4199
g4008 and asqrt[39] n4199 ; n4200
g4009 nor n3877 n3886 ; n4201
g4010 and asqrt[39] n4201 ; n4202
g4011 nor n3884 n4202 ; n4203
g4012 nor n4200 n4203 ; n4204
g4013 nor asqrt[60] n4185 ; n4205
g4014 and n4195_not n4205 ; n4206
g4015 nor n4204 n4206 ; n4207
g4016 nor n4197 n4207 ; n4208
g4017 and asqrt[61] n4208_not ; n4209
g4018 and n3896 n3898_not ; n4210
g4019 and n3889_not n4210 ; n4211
g4020 and asqrt[39] n4211 ; n4212
g4021 nor n3889 n3898 ; n4213
g4022 and asqrt[39] n4213 ; n4214
g4023 nor n3896 n4214 ; n4215
g4024 nor n4212 n4215 ; n4216
g4025 nor asqrt[61] n4197 ; n4217
g4026 and n4207_not n4217 ; n4218
g4027 nor n4216 n4218 ; n4219
g4028 nor n4209 n4219 ; n4220
g4029 and asqrt[62] n4220_not ; n4221
g4030 and n3901_not n3908 ; n4222
g4031 and n3910_not n4222 ; n4223
g4032 and asqrt[39] n4223 ; n4224
g4033 nor n3901 n3910 ; n4225
g4034 and asqrt[39] n4225 ; n4226
g4035 nor n3908 n4226 ; n4227
g4036 nor n4224 n4227 ; n4228
g4037 nor asqrt[62] n4209 ; n4229
g4038 and n4219_not n4229 ; n4230
g4039 nor n4228 n4230 ; n4231
g4040 nor n4221 n4231 ; n4232
g4041 and n3920 n3922_not ; n4233
g4042 and n3913_not n4233 ; n4234
g4043 and asqrt[39] n4234 ; n4235
g4044 nor n3913 n3922 ; n4236
g4045 and asqrt[39] n4236 ; n4237
g4046 nor n3920 n4237 ; n4238
g4047 nor n4235 n4238 ; n4239
g4048 nor n3924 n3931 ; n4240
g4049 and asqrt[39] n4240 ; n4241
g4050 nor n3939 n4241 ; n4242
g4051 and n4239_not n4242 ; n4243
g4052 and n4232_not n4243 ; n4244
g4053 nor asqrt[63] n4244 ; n4245
g4054 and n4221_not n4239 ; n4246
g4055 and n4231_not n4246 ; n4247
g4056 and n3931_not asqrt[39] ; n4248
g4057 and n3924 n4248_not ; n4249
g4058 and asqrt[63] n4240_not ; n4250
g4059 and n4249_not n4250 ; n4251
g4060 nor n3927 n3948 ; n4252
g4061 and n3930_not n4252 ; n4253
g4062 and n3943_not n4253 ; n4254
g4063 and n3939_not n4254 ; n4255
g4064 and n3937_not n4255 ; n4256
g4065 nor n4251 n4256 ; n4257
g4066 and n4247_not n4257 ; n4258
g4067 nand n4245_not n4258 ; asqrt[38]
g4068 and a[76] asqrt[38] ; n4260
g4069 nor a[74] a[75] ; n4261
g4070 and a[76]_not n4261 ; n4262
g4071 nor n4260 n4262 ; n4263
g4072 and asqrt[39] n4263_not ; n4264
g4073 nor n3948 n4262 ; n4265
g4074 and n3943_not n4265 ; n4266
g4075 and n3939_not n4266 ; n4267
g4076 and n3937_not n4267 ; n4268
g4077 and n4260_not n4268 ; n4269
g4078 and a[76]_not asqrt[38] ; n4270
g4079 and a[77] n4270_not ; n4271
g4080 and n3953 asqrt[38] ; n4272
g4081 nor n4271 n4272 ; n4273
g4082 and n4269_not n4273 ; n4274
g4083 nor n4264 n4274 ; n4275
g4084 and asqrt[40] n4275_not ; n4276
g4085 nor asqrt[40] n4264 ; n4277
g4086 and n4274_not n4277 ; n4278
g4087 and asqrt[39] n4256_not ; n4279
g4088 and n4251_not n4279 ; n4280
g4089 and n4247_not n4280 ; n4281
g4090 and n4245_not n4281 ; n4282
g4091 nor n4272 n4282 ; n4283
g4092 and a[78] n4283_not ; n4284
g4093 nor a[78] n4282 ; n4285
g4094 and n4272_not n4285 ; n4286
g4095 nor n4284 n4286 ; n4287
g4096 nor n4278 n4287 ; n4288
g4097 nor n4276 n4288 ; n4289
g4098 and asqrt[41] n4289_not ; n4290
g4099 nor n3956 n3961 ; n4291
g4100 and n3965_not n4291 ; n4292
g4101 and asqrt[38] n4292 ; n4293
g4102 and asqrt[38] n4291 ; n4294
g4103 and n3965 n4294_not ; n4295
g4104 nor n4293 n4295 ; n4296
g4105 nor asqrt[41] n4276 ; n4297
g4106 and n4288_not n4297 ; n4298
g4107 nor n4296 n4298 ; n4299
g4108 nor n4290 n4299 ; n4300
g4109 and asqrt[42] n4300_not ; n4301
g4110 and n3970_not n3979 ; n4302
g4111 and n3968_not n4302 ; n4303
g4112 and asqrt[38] n4303 ; n4304
g4113 nor n3968 n3970 ; n4305
g4114 and asqrt[38] n4305 ; n4306
g4115 nor n3979 n4306 ; n4307
g4116 nor n4304 n4307 ; n4308
g4117 nor asqrt[42] n4290 ; n4309
g4118 and n4299_not n4309 ; n4310
g4119 nor n4308 n4310 ; n4311
g4120 nor n4301 n4311 ; n4312
g4121 and asqrt[43] n4312_not ; n4313
g4122 and n3982_not n3988 ; n4314
g4123 and n3990_not n4314 ; n4315
g4124 and asqrt[38] n4315 ; n4316
g4125 nor n3982 n3990 ; n4317
g4126 and asqrt[38] n4317 ; n4318
g4127 nor n3988 n4318 ; n4319
g4128 nor n4316 n4319 ; n4320
g4129 nor asqrt[43] n4301 ; n4321
g4130 and n4311_not n4321 ; n4322
g4131 nor n4320 n4322 ; n4323
g4132 nor n4313 n4323 ; n4324
g4133 and asqrt[44] n4324_not ; n4325
g4134 and n4000 n4002_not ; n4326
g4135 and n3993_not n4326 ; n4327
g4136 and asqrt[38] n4327 ; n4328
g4137 nor n3993 n4002 ; n4329
g4138 and asqrt[38] n4329 ; n4330
g4139 nor n4000 n4330 ; n4331
g4140 nor n4328 n4331 ; n4332
g4141 nor asqrt[44] n4313 ; n4333
g4142 and n4323_not n4333 ; n4334
g4143 nor n4332 n4334 ; n4335
g4144 nor n4325 n4335 ; n4336
g4145 and asqrt[45] n4336_not ; n4337
g4146 and n4005_not n4012 ; n4338
g4147 and n4014_not n4338 ; n4339
g4148 and asqrt[38] n4339 ; n4340
g4149 nor n4005 n4014 ; n4341
g4150 and asqrt[38] n4341 ; n4342
g4151 nor n4012 n4342 ; n4343
g4152 nor n4340 n4343 ; n4344
g4153 nor asqrt[45] n4325 ; n4345
g4154 and n4335_not n4345 ; n4346
g4155 nor n4344 n4346 ; n4347
g4156 nor n4337 n4347 ; n4348
g4157 and asqrt[46] n4348_not ; n4349
g4158 and n4024 n4026_not ; n4350
g4159 and n4017_not n4350 ; n4351
g4160 and asqrt[38] n4351 ; n4352
g4161 nor n4017 n4026 ; n4353
g4162 and asqrt[38] n4353 ; n4354
g4163 nor n4024 n4354 ; n4355
g4164 nor n4352 n4355 ; n4356
g4165 nor asqrt[46] n4337 ; n4357
g4166 and n4347_not n4357 ; n4358
g4167 nor n4356 n4358 ; n4359
g4168 nor n4349 n4359 ; n4360
g4169 and asqrt[47] n4360_not ; n4361
g4170 and n4029_not n4036 ; n4362
g4171 and n4038_not n4362 ; n4363
g4172 and asqrt[38] n4363 ; n4364
g4173 nor n4029 n4038 ; n4365
g4174 and asqrt[38] n4365 ; n4366
g4175 nor n4036 n4366 ; n4367
g4176 nor n4364 n4367 ; n4368
g4177 nor asqrt[47] n4349 ; n4369
g4178 and n4359_not n4369 ; n4370
g4179 nor n4368 n4370 ; n4371
g4180 nor n4361 n4371 ; n4372
g4181 and asqrt[48] n4372_not ; n4373
g4182 and n4048 n4050_not ; n4374
g4183 and n4041_not n4374 ; n4375
g4184 and asqrt[38] n4375 ; n4376
g4185 nor n4041 n4050 ; n4377
g4186 and asqrt[38] n4377 ; n4378
g4187 nor n4048 n4378 ; n4379
g4188 nor n4376 n4379 ; n4380
g4189 nor asqrt[48] n4361 ; n4381
g4190 and n4371_not n4381 ; n4382
g4191 nor n4380 n4382 ; n4383
g4192 nor n4373 n4383 ; n4384
g4193 and asqrt[49] n4384_not ; n4385
g4194 and n4053_not n4060 ; n4386
g4195 and n4062_not n4386 ; n4387
g4196 and asqrt[38] n4387 ; n4388
g4197 nor n4053 n4062 ; n4389
g4198 and asqrt[38] n4389 ; n4390
g4199 nor n4060 n4390 ; n4391
g4200 nor n4388 n4391 ; n4392
g4201 nor asqrt[49] n4373 ; n4393
g4202 and n4383_not n4393 ; n4394
g4203 nor n4392 n4394 ; n4395
g4204 nor n4385 n4395 ; n4396
g4205 and asqrt[50] n4396_not ; n4397
g4206 and n4072 n4074_not ; n4398
g4207 and n4065_not n4398 ; n4399
g4208 and asqrt[38] n4399 ; n4400
g4209 nor n4065 n4074 ; n4401
g4210 and asqrt[38] n4401 ; n4402
g4211 nor n4072 n4402 ; n4403
g4212 nor n4400 n4403 ; n4404
g4213 nor asqrt[50] n4385 ; n4405
g4214 and n4395_not n4405 ; n4406
g4215 nor n4404 n4406 ; n4407
g4216 nor n4397 n4407 ; n4408
g4217 and asqrt[51] n4408_not ; n4409
g4218 and n4077_not n4084 ; n4410
g4219 and n4086_not n4410 ; n4411
g4220 and asqrt[38] n4411 ; n4412
g4221 nor n4077 n4086 ; n4413
g4222 and asqrt[38] n4413 ; n4414
g4223 nor n4084 n4414 ; n4415
g4224 nor n4412 n4415 ; n4416
g4225 nor asqrt[51] n4397 ; n4417
g4226 and n4407_not n4417 ; n4418
g4227 nor n4416 n4418 ; n4419
g4228 nor n4409 n4419 ; n4420
g4229 and asqrt[52] n4420_not ; n4421
g4230 and n4096 n4098_not ; n4422
g4231 and n4089_not n4422 ; n4423
g4232 and asqrt[38] n4423 ; n4424
g4233 nor n4089 n4098 ; n4425
g4234 and asqrt[38] n4425 ; n4426
g4235 nor n4096 n4426 ; n4427
g4236 nor n4424 n4427 ; n4428
g4237 nor asqrt[52] n4409 ; n4429
g4238 and n4419_not n4429 ; n4430
g4239 nor n4428 n4430 ; n4431
g4240 nor n4421 n4431 ; n4432
g4241 and asqrt[53] n4432_not ; n4433
g4242 and n4101_not n4108 ; n4434
g4243 and n4110_not n4434 ; n4435
g4244 and asqrt[38] n4435 ; n4436
g4245 nor n4101 n4110 ; n4437
g4246 and asqrt[38] n4437 ; n4438
g4247 nor n4108 n4438 ; n4439
g4248 nor n4436 n4439 ; n4440
g4249 nor asqrt[53] n4421 ; n4441
g4250 and n4431_not n4441 ; n4442
g4251 nor n4440 n4442 ; n4443
g4252 nor n4433 n4443 ; n4444
g4253 and asqrt[54] n4444_not ; n4445
g4254 and n4120 n4122_not ; n4446
g4255 and n4113_not n4446 ; n4447
g4256 and asqrt[38] n4447 ; n4448
g4257 nor n4113 n4122 ; n4449
g4258 and asqrt[38] n4449 ; n4450
g4259 nor n4120 n4450 ; n4451
g4260 nor n4448 n4451 ; n4452
g4261 nor asqrt[54] n4433 ; n4453
g4262 and n4443_not n4453 ; n4454
g4263 nor n4452 n4454 ; n4455
g4264 nor n4445 n4455 ; n4456
g4265 and asqrt[55] n4456_not ; n4457
g4266 and n4125_not n4132 ; n4458
g4267 and n4134_not n4458 ; n4459
g4268 and asqrt[38] n4459 ; n4460
g4269 nor n4125 n4134 ; n4461
g4270 and asqrt[38] n4461 ; n4462
g4271 nor n4132 n4462 ; n4463
g4272 nor n4460 n4463 ; n4464
g4273 nor asqrt[55] n4445 ; n4465
g4274 and n4455_not n4465 ; n4466
g4275 nor n4464 n4466 ; n4467
g4276 nor n4457 n4467 ; n4468
g4277 and asqrt[56] n4468_not ; n4469
g4278 and n4144 n4146_not ; n4470
g4279 and n4137_not n4470 ; n4471
g4280 and asqrt[38] n4471 ; n4472
g4281 nor n4137 n4146 ; n4473
g4282 and asqrt[38] n4473 ; n4474
g4283 nor n4144 n4474 ; n4475
g4284 nor n4472 n4475 ; n4476
g4285 nor asqrt[56] n4457 ; n4477
g4286 and n4467_not n4477 ; n4478
g4287 nor n4476 n4478 ; n4479
g4288 nor n4469 n4479 ; n4480
g4289 and asqrt[57] n4480_not ; n4481
g4290 and n4149_not n4156 ; n4482
g4291 and n4158_not n4482 ; n4483
g4292 and asqrt[38] n4483 ; n4484
g4293 nor n4149 n4158 ; n4485
g4294 and asqrt[38] n4485 ; n4486
g4295 nor n4156 n4486 ; n4487
g4296 nor n4484 n4487 ; n4488
g4297 nor asqrt[57] n4469 ; n4489
g4298 and n4479_not n4489 ; n4490
g4299 nor n4488 n4490 ; n4491
g4300 nor n4481 n4491 ; n4492
g4301 and asqrt[58] n4492_not ; n4493
g4302 and n4168 n4170_not ; n4494
g4303 and n4161_not n4494 ; n4495
g4304 and asqrt[38] n4495 ; n4496
g4305 nor n4161 n4170 ; n4497
g4306 and asqrt[38] n4497 ; n4498
g4307 nor n4168 n4498 ; n4499
g4308 nor n4496 n4499 ; n4500
g4309 nor asqrt[58] n4481 ; n4501
g4310 and n4491_not n4501 ; n4502
g4311 nor n4500 n4502 ; n4503
g4312 nor n4493 n4503 ; n4504
g4313 and asqrt[59] n4504_not ; n4505
g4314 nor asqrt[59] n4493 ; n4506
g4315 and n4503_not n4506 ; n4507
g4316 and n4173_not n4182 ; n4508
g4317 and n4175_not n4508 ; n4509
g4318 and asqrt[38] n4509 ; n4510
g4319 nor n4173 n4175 ; n4511
g4320 and asqrt[38] n4511 ; n4512
g4321 nor n4182 n4512 ; n4513
g4322 nor n4510 n4513 ; n4514
g4323 nor n4507 n4514 ; n4515
g4324 nor n4505 n4515 ; n4516
g4325 and asqrt[60] n4516_not ; n4517
g4326 and n4192 n4194_not ; n4518
g4327 and n4185_not n4518 ; n4519
g4328 and asqrt[38] n4519 ; n4520
g4329 nor n4185 n4194 ; n4521
g4330 and asqrt[38] n4521 ; n4522
g4331 nor n4192 n4522 ; n4523
g4332 nor n4520 n4523 ; n4524
g4333 nor asqrt[60] n4505 ; n4525
g4334 and n4515_not n4525 ; n4526
g4335 nor n4524 n4526 ; n4527
g4336 nor n4517 n4527 ; n4528
g4337 and asqrt[61] n4528_not ; n4529
g4338 and n4197_not n4204 ; n4530
g4339 and n4206_not n4530 ; n4531
g4340 and asqrt[38] n4531 ; n4532
g4341 nor n4197 n4206 ; n4533
g4342 and asqrt[38] n4533 ; n4534
g4343 nor n4204 n4534 ; n4535
g4344 nor n4532 n4535 ; n4536
g4345 nor asqrt[61] n4517 ; n4537
g4346 and n4527_not n4537 ; n4538
g4347 nor n4536 n4538 ; n4539
g4348 nor n4529 n4539 ; n4540
g4349 and asqrt[62] n4540_not ; n4541
g4350 and n4216 n4218_not ; n4542
g4351 and n4209_not n4542 ; n4543
g4352 and asqrt[38] n4543 ; n4544
g4353 nor n4209 n4218 ; n4545
g4354 and asqrt[38] n4545 ; n4546
g4355 nor n4216 n4546 ; n4547
g4356 nor n4544 n4547 ; n4548
g4357 nor asqrt[62] n4529 ; n4549
g4358 and n4539_not n4549 ; n4550
g4359 nor n4548 n4550 ; n4551
g4360 nor n4541 n4551 ; n4552
g4361 and n4221_not n4228 ; n4553
g4362 and n4230_not n4553 ; n4554
g4363 and asqrt[38] n4554 ; n4555
g4364 nor n4221 n4230 ; n4556
g4365 and asqrt[38] n4556 ; n4557
g4366 nor n4228 n4557 ; n4558
g4367 nor n4555 n4558 ; n4559
g4368 nor n4232 n4239 ; n4560
g4369 and asqrt[38] n4560 ; n4561
g4370 nor n4247 n4561 ; n4562
g4371 and n4559_not n4562 ; n4563
g4372 and n4552_not n4563 ; n4564
g4373 nor asqrt[63] n4564 ; n4565
g4374 and n4541_not n4559 ; n4566
g4375 and n4551_not n4566 ; n4567
g4376 and n4239_not asqrt[38] ; n4568
g4377 and n4232 n4568_not ; n4569
g4378 and asqrt[63] n4560_not ; n4570
g4379 and n4569_not n4570 ; n4571
g4380 nor n4235 n4256 ; n4572
g4381 and n4238_not n4572 ; n4573
g4382 and n4251_not n4573 ; n4574
g4383 and n4247_not n4574 ; n4575
g4384 and n4245_not n4575 ; n4576
g4385 nor n4571 n4576 ; n4577
g4386 and n4567_not n4577 ; n4578
g4387 nand n4565_not n4578 ; asqrt[37]
g4388 and a[74] asqrt[37] ; n4580
g4389 nor a[72] a[73] ; n4581
g4390 and a[74]_not n4581 ; n4582
g4391 nor n4580 n4582 ; n4583
g4392 and asqrt[38] n4583_not ; n4584
g4393 nor n4256 n4582 ; n4585
g4394 and n4251_not n4585 ; n4586
g4395 and n4247_not n4586 ; n4587
g4396 and n4245_not n4587 ; n4588
g4397 and n4580_not n4588 ; n4589
g4398 and a[74]_not asqrt[37] ; n4590
g4399 and a[75] n4590_not ; n4591
g4400 and n4261 asqrt[37] ; n4592
g4401 nor n4591 n4592 ; n4593
g4402 and n4589_not n4593 ; n4594
g4403 nor n4584 n4594 ; n4595
g4404 and asqrt[39] n4595_not ; n4596
g4405 nor asqrt[39] n4584 ; n4597
g4406 and n4594_not n4597 ; n4598
g4407 and asqrt[38] n4576_not ; n4599
g4408 and n4571_not n4599 ; n4600
g4409 and n4567_not n4600 ; n4601
g4410 and n4565_not n4601 ; n4602
g4411 nor n4592 n4602 ; n4603
g4412 and a[76] n4603_not ; n4604
g4413 nor a[76] n4602 ; n4605
g4414 and n4592_not n4605 ; n4606
g4415 nor n4604 n4606 ; n4607
g4416 nor n4598 n4607 ; n4608
g4417 nor n4596 n4608 ; n4609
g4418 and asqrt[40] n4609_not ; n4610
g4419 nor n4264 n4269 ; n4611
g4420 and n4273_not n4611 ; n4612
g4421 and asqrt[37] n4612 ; n4613
g4422 and asqrt[37] n4611 ; n4614
g4423 and n4273 n4614_not ; n4615
g4424 nor n4613 n4615 ; n4616
g4425 nor asqrt[40] n4596 ; n4617
g4426 and n4608_not n4617 ; n4618
g4427 nor n4616 n4618 ; n4619
g4428 nor n4610 n4619 ; n4620
g4429 and asqrt[41] n4620_not ; n4621
g4430 and n4278_not n4287 ; n4622
g4431 and n4276_not n4622 ; n4623
g4432 and asqrt[37] n4623 ; n4624
g4433 nor n4276 n4278 ; n4625
g4434 and asqrt[37] n4625 ; n4626
g4435 nor n4287 n4626 ; n4627
g4436 nor n4624 n4627 ; n4628
g4437 nor asqrt[41] n4610 ; n4629
g4438 and n4619_not n4629 ; n4630
g4439 nor n4628 n4630 ; n4631
g4440 nor n4621 n4631 ; n4632
g4441 and asqrt[42] n4632_not ; n4633
g4442 and n4290_not n4296 ; n4634
g4443 and n4298_not n4634 ; n4635
g4444 and asqrt[37] n4635 ; n4636
g4445 nor n4290 n4298 ; n4637
g4446 and asqrt[37] n4637 ; n4638
g4447 nor n4296 n4638 ; n4639
g4448 nor n4636 n4639 ; n4640
g4449 nor asqrt[42] n4621 ; n4641
g4450 and n4631_not n4641 ; n4642
g4451 nor n4640 n4642 ; n4643
g4452 nor n4633 n4643 ; n4644
g4453 and asqrt[43] n4644_not ; n4645
g4454 and n4308 n4310_not ; n4646
g4455 and n4301_not n4646 ; n4647
g4456 and asqrt[37] n4647 ; n4648
g4457 nor n4301 n4310 ; n4649
g4458 and asqrt[37] n4649 ; n4650
g4459 nor n4308 n4650 ; n4651
g4460 nor n4648 n4651 ; n4652
g4461 nor asqrt[43] n4633 ; n4653
g4462 and n4643_not n4653 ; n4654
g4463 nor n4652 n4654 ; n4655
g4464 nor n4645 n4655 ; n4656
g4465 and asqrt[44] n4656_not ; n4657
g4466 and n4313_not n4320 ; n4658
g4467 and n4322_not n4658 ; n4659
g4468 and asqrt[37] n4659 ; n4660
g4469 nor n4313 n4322 ; n4661
g4470 and asqrt[37] n4661 ; n4662
g4471 nor n4320 n4662 ; n4663
g4472 nor n4660 n4663 ; n4664
g4473 nor asqrt[44] n4645 ; n4665
g4474 and n4655_not n4665 ; n4666
g4475 nor n4664 n4666 ; n4667
g4476 nor n4657 n4667 ; n4668
g4477 and asqrt[45] n4668_not ; n4669
g4478 and n4332 n4334_not ; n4670
g4479 and n4325_not n4670 ; n4671
g4480 and asqrt[37] n4671 ; n4672
g4481 nor n4325 n4334 ; n4673
g4482 and asqrt[37] n4673 ; n4674
g4483 nor n4332 n4674 ; n4675
g4484 nor n4672 n4675 ; n4676
g4485 nor asqrt[45] n4657 ; n4677
g4486 and n4667_not n4677 ; n4678
g4487 nor n4676 n4678 ; n4679
g4488 nor n4669 n4679 ; n4680
g4489 and asqrt[46] n4680_not ; n4681
g4490 and n4337_not n4344 ; n4682
g4491 and n4346_not n4682 ; n4683
g4492 and asqrt[37] n4683 ; n4684
g4493 nor n4337 n4346 ; n4685
g4494 and asqrt[37] n4685 ; n4686
g4495 nor n4344 n4686 ; n4687
g4496 nor n4684 n4687 ; n4688
g4497 nor asqrt[46] n4669 ; n4689
g4498 and n4679_not n4689 ; n4690
g4499 nor n4688 n4690 ; n4691
g4500 nor n4681 n4691 ; n4692
g4501 and asqrt[47] n4692_not ; n4693
g4502 and n4356 n4358_not ; n4694
g4503 and n4349_not n4694 ; n4695
g4504 and asqrt[37] n4695 ; n4696
g4505 nor n4349 n4358 ; n4697
g4506 and asqrt[37] n4697 ; n4698
g4507 nor n4356 n4698 ; n4699
g4508 nor n4696 n4699 ; n4700
g4509 nor asqrt[47] n4681 ; n4701
g4510 and n4691_not n4701 ; n4702
g4511 nor n4700 n4702 ; n4703
g4512 nor n4693 n4703 ; n4704
g4513 and asqrt[48] n4704_not ; n4705
g4514 and n4361_not n4368 ; n4706
g4515 and n4370_not n4706 ; n4707
g4516 and asqrt[37] n4707 ; n4708
g4517 nor n4361 n4370 ; n4709
g4518 and asqrt[37] n4709 ; n4710
g4519 nor n4368 n4710 ; n4711
g4520 nor n4708 n4711 ; n4712
g4521 nor asqrt[48] n4693 ; n4713
g4522 and n4703_not n4713 ; n4714
g4523 nor n4712 n4714 ; n4715
g4524 nor n4705 n4715 ; n4716
g4525 and asqrt[49] n4716_not ; n4717
g4526 and n4380 n4382_not ; n4718
g4527 and n4373_not n4718 ; n4719
g4528 and asqrt[37] n4719 ; n4720
g4529 nor n4373 n4382 ; n4721
g4530 and asqrt[37] n4721 ; n4722
g4531 nor n4380 n4722 ; n4723
g4532 nor n4720 n4723 ; n4724
g4533 nor asqrt[49] n4705 ; n4725
g4534 and n4715_not n4725 ; n4726
g4535 nor n4724 n4726 ; n4727
g4536 nor n4717 n4727 ; n4728
g4537 and asqrt[50] n4728_not ; n4729
g4538 and n4385_not n4392 ; n4730
g4539 and n4394_not n4730 ; n4731
g4540 and asqrt[37] n4731 ; n4732
g4541 nor n4385 n4394 ; n4733
g4542 and asqrt[37] n4733 ; n4734
g4543 nor n4392 n4734 ; n4735
g4544 nor n4732 n4735 ; n4736
g4545 nor asqrt[50] n4717 ; n4737
g4546 and n4727_not n4737 ; n4738
g4547 nor n4736 n4738 ; n4739
g4548 nor n4729 n4739 ; n4740
g4549 and asqrt[51] n4740_not ; n4741
g4550 and n4404 n4406_not ; n4742
g4551 and n4397_not n4742 ; n4743
g4552 and asqrt[37] n4743 ; n4744
g4553 nor n4397 n4406 ; n4745
g4554 and asqrt[37] n4745 ; n4746
g4555 nor n4404 n4746 ; n4747
g4556 nor n4744 n4747 ; n4748
g4557 nor asqrt[51] n4729 ; n4749
g4558 and n4739_not n4749 ; n4750
g4559 nor n4748 n4750 ; n4751
g4560 nor n4741 n4751 ; n4752
g4561 and asqrt[52] n4752_not ; n4753
g4562 and n4409_not n4416 ; n4754
g4563 and n4418_not n4754 ; n4755
g4564 and asqrt[37] n4755 ; n4756
g4565 nor n4409 n4418 ; n4757
g4566 and asqrt[37] n4757 ; n4758
g4567 nor n4416 n4758 ; n4759
g4568 nor n4756 n4759 ; n4760
g4569 nor asqrt[52] n4741 ; n4761
g4570 and n4751_not n4761 ; n4762
g4571 nor n4760 n4762 ; n4763
g4572 nor n4753 n4763 ; n4764
g4573 and asqrt[53] n4764_not ; n4765
g4574 and n4428 n4430_not ; n4766
g4575 and n4421_not n4766 ; n4767
g4576 and asqrt[37] n4767 ; n4768
g4577 nor n4421 n4430 ; n4769
g4578 and asqrt[37] n4769 ; n4770
g4579 nor n4428 n4770 ; n4771
g4580 nor n4768 n4771 ; n4772
g4581 nor asqrt[53] n4753 ; n4773
g4582 and n4763_not n4773 ; n4774
g4583 nor n4772 n4774 ; n4775
g4584 nor n4765 n4775 ; n4776
g4585 and asqrt[54] n4776_not ; n4777
g4586 and n4433_not n4440 ; n4778
g4587 and n4442_not n4778 ; n4779
g4588 and asqrt[37] n4779 ; n4780
g4589 nor n4433 n4442 ; n4781
g4590 and asqrt[37] n4781 ; n4782
g4591 nor n4440 n4782 ; n4783
g4592 nor n4780 n4783 ; n4784
g4593 nor asqrt[54] n4765 ; n4785
g4594 and n4775_not n4785 ; n4786
g4595 nor n4784 n4786 ; n4787
g4596 nor n4777 n4787 ; n4788
g4597 and asqrt[55] n4788_not ; n4789
g4598 and n4452 n4454_not ; n4790
g4599 and n4445_not n4790 ; n4791
g4600 and asqrt[37] n4791 ; n4792
g4601 nor n4445 n4454 ; n4793
g4602 and asqrt[37] n4793 ; n4794
g4603 nor n4452 n4794 ; n4795
g4604 nor n4792 n4795 ; n4796
g4605 nor asqrt[55] n4777 ; n4797
g4606 and n4787_not n4797 ; n4798
g4607 nor n4796 n4798 ; n4799
g4608 nor n4789 n4799 ; n4800
g4609 and asqrt[56] n4800_not ; n4801
g4610 and n4457_not n4464 ; n4802
g4611 and n4466_not n4802 ; n4803
g4612 and asqrt[37] n4803 ; n4804
g4613 nor n4457 n4466 ; n4805
g4614 and asqrt[37] n4805 ; n4806
g4615 nor n4464 n4806 ; n4807
g4616 nor n4804 n4807 ; n4808
g4617 nor asqrt[56] n4789 ; n4809
g4618 and n4799_not n4809 ; n4810
g4619 nor n4808 n4810 ; n4811
g4620 nor n4801 n4811 ; n4812
g4621 and asqrt[57] n4812_not ; n4813
g4622 and n4476 n4478_not ; n4814
g4623 and n4469_not n4814 ; n4815
g4624 and asqrt[37] n4815 ; n4816
g4625 nor n4469 n4478 ; n4817
g4626 and asqrt[37] n4817 ; n4818
g4627 nor n4476 n4818 ; n4819
g4628 nor n4816 n4819 ; n4820
g4629 nor asqrt[57] n4801 ; n4821
g4630 and n4811_not n4821 ; n4822
g4631 nor n4820 n4822 ; n4823
g4632 nor n4813 n4823 ; n4824
g4633 and asqrt[58] n4824_not ; n4825
g4634 and n4481_not n4488 ; n4826
g4635 and n4490_not n4826 ; n4827
g4636 and asqrt[37] n4827 ; n4828
g4637 nor n4481 n4490 ; n4829
g4638 and asqrt[37] n4829 ; n4830
g4639 nor n4488 n4830 ; n4831
g4640 nor n4828 n4831 ; n4832
g4641 nor asqrt[58] n4813 ; n4833
g4642 and n4823_not n4833 ; n4834
g4643 nor n4832 n4834 ; n4835
g4644 nor n4825 n4835 ; n4836
g4645 and asqrt[59] n4836_not ; n4837
g4646 and n4500 n4502_not ; n4838
g4647 and n4493_not n4838 ; n4839
g4648 and asqrt[37] n4839 ; n4840
g4649 nor n4493 n4502 ; n4841
g4650 and asqrt[37] n4841 ; n4842
g4651 nor n4500 n4842 ; n4843
g4652 nor n4840 n4843 ; n4844
g4653 nor asqrt[59] n4825 ; n4845
g4654 and n4835_not n4845 ; n4846
g4655 nor n4844 n4846 ; n4847
g4656 nor n4837 n4847 ; n4848
g4657 and asqrt[60] n4848_not ; n4849
g4658 nor asqrt[60] n4837 ; n4850
g4659 and n4847_not n4850 ; n4851
g4660 and n4505_not n4514 ; n4852
g4661 and n4507_not n4852 ; n4853
g4662 and asqrt[37] n4853 ; n4854
g4663 nor n4505 n4507 ; n4855
g4664 and asqrt[37] n4855 ; n4856
g4665 nor n4514 n4856 ; n4857
g4666 nor n4854 n4857 ; n4858
g4667 nor n4851 n4858 ; n4859
g4668 nor n4849 n4859 ; n4860
g4669 and asqrt[61] n4860_not ; n4861
g4670 and n4524 n4526_not ; n4862
g4671 and n4517_not n4862 ; n4863
g4672 and asqrt[37] n4863 ; n4864
g4673 nor n4517 n4526 ; n4865
g4674 and asqrt[37] n4865 ; n4866
g4675 nor n4524 n4866 ; n4867
g4676 nor n4864 n4867 ; n4868
g4677 nor asqrt[61] n4849 ; n4869
g4678 and n4859_not n4869 ; n4870
g4679 nor n4868 n4870 ; n4871
g4680 nor n4861 n4871 ; n4872
g4681 and asqrt[62] n4872_not ; n4873
g4682 and n4529_not n4536 ; n4874
g4683 and n4538_not n4874 ; n4875
g4684 and asqrt[37] n4875 ; n4876
g4685 nor n4529 n4538 ; n4877
g4686 and asqrt[37] n4877 ; n4878
g4687 nor n4536 n4878 ; n4879
g4688 nor n4876 n4879 ; n4880
g4689 nor asqrt[62] n4861 ; n4881
g4690 and n4871_not n4881 ; n4882
g4691 nor n4880 n4882 ; n4883
g4692 nor n4873 n4883 ; n4884
g4693 and n4548 n4550_not ; n4885
g4694 and n4541_not n4885 ; n4886
g4695 and asqrt[37] n4886 ; n4887
g4696 nor n4541 n4550 ; n4888
g4697 and asqrt[37] n4888 ; n4889
g4698 nor n4548 n4889 ; n4890
g4699 nor n4887 n4890 ; n4891
g4700 nor n4552 n4559 ; n4892
g4701 and asqrt[37] n4892 ; n4893
g4702 nor n4567 n4893 ; n4894
g4703 and n4891_not n4894 ; n4895
g4704 and n4884_not n4895 ; n4896
g4705 nor asqrt[63] n4896 ; n4897
g4706 and n4873_not n4891 ; n4898
g4707 and n4883_not n4898 ; n4899
g4708 and n4559_not asqrt[37] ; n4900
g4709 and n4552 n4900_not ; n4901
g4710 and asqrt[63] n4892_not ; n4902
g4711 and n4901_not n4902 ; n4903
g4712 nor n4555 n4576 ; n4904
g4713 and n4558_not n4904 ; n4905
g4714 and n4571_not n4905 ; n4906
g4715 and n4567_not n4906 ; n4907
g4716 and n4565_not n4907 ; n4908
g4717 nor n4903 n4908 ; n4909
g4718 and n4899_not n4909 ; n4910
g4719 nand n4897_not n4910 ; asqrt[36]
g4720 and a[72] asqrt[36] ; n4912
g4721 nor a[70] a[71] ; n4913
g4722 and a[72]_not n4913 ; n4914
g4723 nor n4912 n4914 ; n4915
g4724 and asqrt[37] n4915_not ; n4916
g4725 nor n4576 n4914 ; n4917
g4726 and n4571_not n4917 ; n4918
g4727 and n4567_not n4918 ; n4919
g4728 and n4565_not n4919 ; n4920
g4729 and n4912_not n4920 ; n4921
g4730 and a[72]_not asqrt[36] ; n4922
g4731 and a[73] n4922_not ; n4923
g4732 and n4581 asqrt[36] ; n4924
g4733 nor n4923 n4924 ; n4925
g4734 and n4921_not n4925 ; n4926
g4735 nor n4916 n4926 ; n4927
g4736 and asqrt[38] n4927_not ; n4928
g4737 nor asqrt[38] n4916 ; n4929
g4738 and n4926_not n4929 ; n4930
g4739 and asqrt[37] n4908_not ; n4931
g4740 and n4903_not n4931 ; n4932
g4741 and n4899_not n4932 ; n4933
g4742 and n4897_not n4933 ; n4934
g4743 nor n4924 n4934 ; n4935
g4744 and a[74] n4935_not ; n4936
g4745 nor a[74] n4934 ; n4937
g4746 and n4924_not n4937 ; n4938
g4747 nor n4936 n4938 ; n4939
g4748 nor n4930 n4939 ; n4940
g4749 nor n4928 n4940 ; n4941
g4750 and asqrt[39] n4941_not ; n4942
g4751 nor n4584 n4589 ; n4943
g4752 and n4593_not n4943 ; n4944
g4753 and asqrt[36] n4944 ; n4945
g4754 and asqrt[36] n4943 ; n4946
g4755 and n4593 n4946_not ; n4947
g4756 nor n4945 n4947 ; n4948
g4757 nor asqrt[39] n4928 ; n4949
g4758 and n4940_not n4949 ; n4950
g4759 nor n4948 n4950 ; n4951
g4760 nor n4942 n4951 ; n4952
g4761 and asqrt[40] n4952_not ; n4953
g4762 and n4598_not n4607 ; n4954
g4763 and n4596_not n4954 ; n4955
g4764 and asqrt[36] n4955 ; n4956
g4765 nor n4596 n4598 ; n4957
g4766 and asqrt[36] n4957 ; n4958
g4767 nor n4607 n4958 ; n4959
g4768 nor n4956 n4959 ; n4960
g4769 nor asqrt[40] n4942 ; n4961
g4770 and n4951_not n4961 ; n4962
g4771 nor n4960 n4962 ; n4963
g4772 nor n4953 n4963 ; n4964
g4773 and asqrt[41] n4964_not ; n4965
g4774 and n4610_not n4616 ; n4966
g4775 and n4618_not n4966 ; n4967
g4776 and asqrt[36] n4967 ; n4968
g4777 nor n4610 n4618 ; n4969
g4778 and asqrt[36] n4969 ; n4970
g4779 nor n4616 n4970 ; n4971
g4780 nor n4968 n4971 ; n4972
g4781 nor asqrt[41] n4953 ; n4973
g4782 and n4963_not n4973 ; n4974
g4783 nor n4972 n4974 ; n4975
g4784 nor n4965 n4975 ; n4976
g4785 and asqrt[42] n4976_not ; n4977
g4786 and n4628 n4630_not ; n4978
g4787 and n4621_not n4978 ; n4979
g4788 and asqrt[36] n4979 ; n4980
g4789 nor n4621 n4630 ; n4981
g4790 and asqrt[36] n4981 ; n4982
g4791 nor n4628 n4982 ; n4983
g4792 nor n4980 n4983 ; n4984
g4793 nor asqrt[42] n4965 ; n4985
g4794 and n4975_not n4985 ; n4986
g4795 nor n4984 n4986 ; n4987
g4796 nor n4977 n4987 ; n4988
g4797 and asqrt[43] n4988_not ; n4989
g4798 and n4633_not n4640 ; n4990
g4799 and n4642_not n4990 ; n4991
g4800 and asqrt[36] n4991 ; n4992
g4801 nor n4633 n4642 ; n4993
g4802 and asqrt[36] n4993 ; n4994
g4803 nor n4640 n4994 ; n4995
g4804 nor n4992 n4995 ; n4996
g4805 nor asqrt[43] n4977 ; n4997
g4806 and n4987_not n4997 ; n4998
g4807 nor n4996 n4998 ; n4999
g4808 nor n4989 n4999 ; n5000
g4809 and asqrt[44] n5000_not ; n5001
g4810 and n4652 n4654_not ; n5002
g4811 and n4645_not n5002 ; n5003
g4812 and asqrt[36] n5003 ; n5004
g4813 nor n4645 n4654 ; n5005
g4814 and asqrt[36] n5005 ; n5006
g4815 nor n4652 n5006 ; n5007
g4816 nor n5004 n5007 ; n5008
g4817 nor asqrt[44] n4989 ; n5009
g4818 and n4999_not n5009 ; n5010
g4819 nor n5008 n5010 ; n5011
g4820 nor n5001 n5011 ; n5012
g4821 and asqrt[45] n5012_not ; n5013
g4822 and n4657_not n4664 ; n5014
g4823 and n4666_not n5014 ; n5015
g4824 and asqrt[36] n5015 ; n5016
g4825 nor n4657 n4666 ; n5017
g4826 and asqrt[36] n5017 ; n5018
g4827 nor n4664 n5018 ; n5019
g4828 nor n5016 n5019 ; n5020
g4829 nor asqrt[45] n5001 ; n5021
g4830 and n5011_not n5021 ; n5022
g4831 nor n5020 n5022 ; n5023
g4832 nor n5013 n5023 ; n5024
g4833 and asqrt[46] n5024_not ; n5025
g4834 and n4676 n4678_not ; n5026
g4835 and n4669_not n5026 ; n5027
g4836 and asqrt[36] n5027 ; n5028
g4837 nor n4669 n4678 ; n5029
g4838 and asqrt[36] n5029 ; n5030
g4839 nor n4676 n5030 ; n5031
g4840 nor n5028 n5031 ; n5032
g4841 nor asqrt[46] n5013 ; n5033
g4842 and n5023_not n5033 ; n5034
g4843 nor n5032 n5034 ; n5035
g4844 nor n5025 n5035 ; n5036
g4845 and asqrt[47] n5036_not ; n5037
g4846 and n4681_not n4688 ; n5038
g4847 and n4690_not n5038 ; n5039
g4848 and asqrt[36] n5039 ; n5040
g4849 nor n4681 n4690 ; n5041
g4850 and asqrt[36] n5041 ; n5042
g4851 nor n4688 n5042 ; n5043
g4852 nor n5040 n5043 ; n5044
g4853 nor asqrt[47] n5025 ; n5045
g4854 and n5035_not n5045 ; n5046
g4855 nor n5044 n5046 ; n5047
g4856 nor n5037 n5047 ; n5048
g4857 and asqrt[48] n5048_not ; n5049
g4858 and n4700 n4702_not ; n5050
g4859 and n4693_not n5050 ; n5051
g4860 and asqrt[36] n5051 ; n5052
g4861 nor n4693 n4702 ; n5053
g4862 and asqrt[36] n5053 ; n5054
g4863 nor n4700 n5054 ; n5055
g4864 nor n5052 n5055 ; n5056
g4865 nor asqrt[48] n5037 ; n5057
g4866 and n5047_not n5057 ; n5058
g4867 nor n5056 n5058 ; n5059
g4868 nor n5049 n5059 ; n5060
g4869 and asqrt[49] n5060_not ; n5061
g4870 and n4705_not n4712 ; n5062
g4871 and n4714_not n5062 ; n5063
g4872 and asqrt[36] n5063 ; n5064
g4873 nor n4705 n4714 ; n5065
g4874 and asqrt[36] n5065 ; n5066
g4875 nor n4712 n5066 ; n5067
g4876 nor n5064 n5067 ; n5068
g4877 nor asqrt[49] n5049 ; n5069
g4878 and n5059_not n5069 ; n5070
g4879 nor n5068 n5070 ; n5071
g4880 nor n5061 n5071 ; n5072
g4881 and asqrt[50] n5072_not ; n5073
g4882 and n4724 n4726_not ; n5074
g4883 and n4717_not n5074 ; n5075
g4884 and asqrt[36] n5075 ; n5076
g4885 nor n4717 n4726 ; n5077
g4886 and asqrt[36] n5077 ; n5078
g4887 nor n4724 n5078 ; n5079
g4888 nor n5076 n5079 ; n5080
g4889 nor asqrt[50] n5061 ; n5081
g4890 and n5071_not n5081 ; n5082
g4891 nor n5080 n5082 ; n5083
g4892 nor n5073 n5083 ; n5084
g4893 and asqrt[51] n5084_not ; n5085
g4894 and n4729_not n4736 ; n5086
g4895 and n4738_not n5086 ; n5087
g4896 and asqrt[36] n5087 ; n5088
g4897 nor n4729 n4738 ; n5089
g4898 and asqrt[36] n5089 ; n5090
g4899 nor n4736 n5090 ; n5091
g4900 nor n5088 n5091 ; n5092
g4901 nor asqrt[51] n5073 ; n5093
g4902 and n5083_not n5093 ; n5094
g4903 nor n5092 n5094 ; n5095
g4904 nor n5085 n5095 ; n5096
g4905 and asqrt[52] n5096_not ; n5097
g4906 and n4748 n4750_not ; n5098
g4907 and n4741_not n5098 ; n5099
g4908 and asqrt[36] n5099 ; n5100
g4909 nor n4741 n4750 ; n5101
g4910 and asqrt[36] n5101 ; n5102
g4911 nor n4748 n5102 ; n5103
g4912 nor n5100 n5103 ; n5104
g4913 nor asqrt[52] n5085 ; n5105
g4914 and n5095_not n5105 ; n5106
g4915 nor n5104 n5106 ; n5107
g4916 nor n5097 n5107 ; n5108
g4917 and asqrt[53] n5108_not ; n5109
g4918 and n4753_not n4760 ; n5110
g4919 and n4762_not n5110 ; n5111
g4920 and asqrt[36] n5111 ; n5112
g4921 nor n4753 n4762 ; n5113
g4922 and asqrt[36] n5113 ; n5114
g4923 nor n4760 n5114 ; n5115
g4924 nor n5112 n5115 ; n5116
g4925 nor asqrt[53] n5097 ; n5117
g4926 and n5107_not n5117 ; n5118
g4927 nor n5116 n5118 ; n5119
g4928 nor n5109 n5119 ; n5120
g4929 and asqrt[54] n5120_not ; n5121
g4930 and n4772 n4774_not ; n5122
g4931 and n4765_not n5122 ; n5123
g4932 and asqrt[36] n5123 ; n5124
g4933 nor n4765 n4774 ; n5125
g4934 and asqrt[36] n5125 ; n5126
g4935 nor n4772 n5126 ; n5127
g4936 nor n5124 n5127 ; n5128
g4937 nor asqrt[54] n5109 ; n5129
g4938 and n5119_not n5129 ; n5130
g4939 nor n5128 n5130 ; n5131
g4940 nor n5121 n5131 ; n5132
g4941 and asqrt[55] n5132_not ; n5133
g4942 and n4777_not n4784 ; n5134
g4943 and n4786_not n5134 ; n5135
g4944 and asqrt[36] n5135 ; n5136
g4945 nor n4777 n4786 ; n5137
g4946 and asqrt[36] n5137 ; n5138
g4947 nor n4784 n5138 ; n5139
g4948 nor n5136 n5139 ; n5140
g4949 nor asqrt[55] n5121 ; n5141
g4950 and n5131_not n5141 ; n5142
g4951 nor n5140 n5142 ; n5143
g4952 nor n5133 n5143 ; n5144
g4953 and asqrt[56] n5144_not ; n5145
g4954 and n4796 n4798_not ; n5146
g4955 and n4789_not n5146 ; n5147
g4956 and asqrt[36] n5147 ; n5148
g4957 nor n4789 n4798 ; n5149
g4958 and asqrt[36] n5149 ; n5150
g4959 nor n4796 n5150 ; n5151
g4960 nor n5148 n5151 ; n5152
g4961 nor asqrt[56] n5133 ; n5153
g4962 and n5143_not n5153 ; n5154
g4963 nor n5152 n5154 ; n5155
g4964 nor n5145 n5155 ; n5156
g4965 and asqrt[57] n5156_not ; n5157
g4966 and n4801_not n4808 ; n5158
g4967 and n4810_not n5158 ; n5159
g4968 and asqrt[36] n5159 ; n5160
g4969 nor n4801 n4810 ; n5161
g4970 and asqrt[36] n5161 ; n5162
g4971 nor n4808 n5162 ; n5163
g4972 nor n5160 n5163 ; n5164
g4973 nor asqrt[57] n5145 ; n5165
g4974 and n5155_not n5165 ; n5166
g4975 nor n5164 n5166 ; n5167
g4976 nor n5157 n5167 ; n5168
g4977 and asqrt[58] n5168_not ; n5169
g4978 and n4820 n4822_not ; n5170
g4979 and n4813_not n5170 ; n5171
g4980 and asqrt[36] n5171 ; n5172
g4981 nor n4813 n4822 ; n5173
g4982 and asqrt[36] n5173 ; n5174
g4983 nor n4820 n5174 ; n5175
g4984 nor n5172 n5175 ; n5176
g4985 nor asqrt[58] n5157 ; n5177
g4986 and n5167_not n5177 ; n5178
g4987 nor n5176 n5178 ; n5179
g4988 nor n5169 n5179 ; n5180
g4989 and asqrt[59] n5180_not ; n5181
g4990 and n4825_not n4832 ; n5182
g4991 and n4834_not n5182 ; n5183
g4992 and asqrt[36] n5183 ; n5184
g4993 nor n4825 n4834 ; n5185
g4994 and asqrt[36] n5185 ; n5186
g4995 nor n4832 n5186 ; n5187
g4996 nor n5184 n5187 ; n5188
g4997 nor asqrt[59] n5169 ; n5189
g4998 and n5179_not n5189 ; n5190
g4999 nor n5188 n5190 ; n5191
g5000 nor n5181 n5191 ; n5192
g5001 and asqrt[60] n5192_not ; n5193
g5002 and n4844 n4846_not ; n5194
g5003 and n4837_not n5194 ; n5195
g5004 and asqrt[36] n5195 ; n5196
g5005 nor n4837 n4846 ; n5197
g5006 and asqrt[36] n5197 ; n5198
g5007 nor n4844 n5198 ; n5199
g5008 nor n5196 n5199 ; n5200
g5009 nor asqrt[60] n5181 ; n5201
g5010 and n5191_not n5201 ; n5202
g5011 nor n5200 n5202 ; n5203
g5012 nor n5193 n5203 ; n5204
g5013 and asqrt[61] n5204_not ; n5205
g5014 nor asqrt[61] n5193 ; n5206
g5015 and n5203_not n5206 ; n5207
g5016 and n4849_not n4858 ; n5208
g5017 and n4851_not n5208 ; n5209
g5018 and asqrt[36] n5209 ; n5210
g5019 nor n4849 n4851 ; n5211
g5020 and asqrt[36] n5211 ; n5212
g5021 nor n4858 n5212 ; n5213
g5022 nor n5210 n5213 ; n5214
g5023 nor n5207 n5214 ; n5215
g5024 nor n5205 n5215 ; n5216
g5025 and asqrt[62] n5216_not ; n5217
g5026 and n4868 n4870_not ; n5218
g5027 and n4861_not n5218 ; n5219
g5028 and asqrt[36] n5219 ; n5220
g5029 nor n4861 n4870 ; n5221
g5030 and asqrt[36] n5221 ; n5222
g5031 nor n4868 n5222 ; n5223
g5032 nor n5220 n5223 ; n5224
g5033 nor asqrt[62] n5205 ; n5225
g5034 and n5215_not n5225 ; n5226
g5035 nor n5224 n5226 ; n5227
g5036 nor n5217 n5227 ; n5228
g5037 and n4873_not n4880 ; n5229
g5038 and n4882_not n5229 ; n5230
g5039 and asqrt[36] n5230 ; n5231
g5040 nor n4873 n4882 ; n5232
g5041 and asqrt[36] n5232 ; n5233
g5042 nor n4880 n5233 ; n5234
g5043 nor n5231 n5234 ; n5235
g5044 nor n4884 n4891 ; n5236
g5045 and asqrt[36] n5236 ; n5237
g5046 nor n4899 n5237 ; n5238
g5047 and n5235_not n5238 ; n5239
g5048 and n5228_not n5239 ; n5240
g5049 nor asqrt[63] n5240 ; n5241
g5050 and n5217_not n5235 ; n5242
g5051 and n5227_not n5242 ; n5243
g5052 and n4891_not asqrt[36] ; n5244
g5053 and n4884 n5244_not ; n5245
g5054 and asqrt[63] n5236_not ; n5246
g5055 and n5245_not n5246 ; n5247
g5056 nor n4887 n4908 ; n5248
g5057 and n4890_not n5248 ; n5249
g5058 and n4903_not n5249 ; n5250
g5059 and n4899_not n5250 ; n5251
g5060 and n4897_not n5251 ; n5252
g5061 nor n5247 n5252 ; n5253
g5062 and n5243_not n5253 ; n5254
g5063 nand n5241_not n5254 ; asqrt[35]
g5064 and a[70] asqrt[35] ; n5256
g5065 nor a[68] a[69] ; n5257
g5066 and a[70]_not n5257 ; n5258
g5067 nor n5256 n5258 ; n5259
g5068 and asqrt[36] n5259_not ; n5260
g5069 nor n4908 n5258 ; n5261
g5070 and n4903_not n5261 ; n5262
g5071 and n4899_not n5262 ; n5263
g5072 and n4897_not n5263 ; n5264
g5073 and n5256_not n5264 ; n5265
g5074 and a[70]_not asqrt[35] ; n5266
g5075 and a[71] n5266_not ; n5267
g5076 and n4913 asqrt[35] ; n5268
g5077 nor n5267 n5268 ; n5269
g5078 and n5265_not n5269 ; n5270
g5079 nor n5260 n5270 ; n5271
g5080 and asqrt[37] n5271_not ; n5272
g5081 nor asqrt[37] n5260 ; n5273
g5082 and n5270_not n5273 ; n5274
g5083 and asqrt[36] n5252_not ; n5275
g5084 and n5247_not n5275 ; n5276
g5085 and n5243_not n5276 ; n5277
g5086 and n5241_not n5277 ; n5278
g5087 nor n5268 n5278 ; n5279
g5088 and a[72] n5279_not ; n5280
g5089 nor a[72] n5278 ; n5281
g5090 and n5268_not n5281 ; n5282
g5091 nor n5280 n5282 ; n5283
g5092 nor n5274 n5283 ; n5284
g5093 nor n5272 n5284 ; n5285
g5094 and asqrt[38] n5285_not ; n5286
g5095 nor n4916 n4921 ; n5287
g5096 and n4925_not n5287 ; n5288
g5097 and asqrt[35] n5288 ; n5289
g5098 and asqrt[35] n5287 ; n5290
g5099 and n4925 n5290_not ; n5291
g5100 nor n5289 n5291 ; n5292
g5101 nor asqrt[38] n5272 ; n5293
g5102 and n5284_not n5293 ; n5294
g5103 nor n5292 n5294 ; n5295
g5104 nor n5286 n5295 ; n5296
g5105 and asqrt[39] n5296_not ; n5297
g5106 and n4930_not n4939 ; n5298
g5107 and n4928_not n5298 ; n5299
g5108 and asqrt[35] n5299 ; n5300
g5109 nor n4928 n4930 ; n5301
g5110 and asqrt[35] n5301 ; n5302
g5111 nor n4939 n5302 ; n5303
g5112 nor n5300 n5303 ; n5304
g5113 nor asqrt[39] n5286 ; n5305
g5114 and n5295_not n5305 ; n5306
g5115 nor n5304 n5306 ; n5307
g5116 nor n5297 n5307 ; n5308
g5117 and asqrt[40] n5308_not ; n5309
g5118 and n4942_not n4948 ; n5310
g5119 and n4950_not n5310 ; n5311
g5120 and asqrt[35] n5311 ; n5312
g5121 nor n4942 n4950 ; n5313
g5122 and asqrt[35] n5313 ; n5314
g5123 nor n4948 n5314 ; n5315
g5124 nor n5312 n5315 ; n5316
g5125 nor asqrt[40] n5297 ; n5317
g5126 and n5307_not n5317 ; n5318
g5127 nor n5316 n5318 ; n5319
g5128 nor n5309 n5319 ; n5320
g5129 and asqrt[41] n5320_not ; n5321
g5130 and n4960 n4962_not ; n5322
g5131 and n4953_not n5322 ; n5323
g5132 and asqrt[35] n5323 ; n5324
g5133 nor n4953 n4962 ; n5325
g5134 and asqrt[35] n5325 ; n5326
g5135 nor n4960 n5326 ; n5327
g5136 nor n5324 n5327 ; n5328
g5137 nor asqrt[41] n5309 ; n5329
g5138 and n5319_not n5329 ; n5330
g5139 nor n5328 n5330 ; n5331
g5140 nor n5321 n5331 ; n5332
g5141 and asqrt[42] n5332_not ; n5333
g5142 and n4965_not n4972 ; n5334
g5143 and n4974_not n5334 ; n5335
g5144 and asqrt[35] n5335 ; n5336
g5145 nor n4965 n4974 ; n5337
g5146 and asqrt[35] n5337 ; n5338
g5147 nor n4972 n5338 ; n5339
g5148 nor n5336 n5339 ; n5340
g5149 nor asqrt[42] n5321 ; n5341
g5150 and n5331_not n5341 ; n5342
g5151 nor n5340 n5342 ; n5343
g5152 nor n5333 n5343 ; n5344
g5153 and asqrt[43] n5344_not ; n5345
g5154 and n4984 n4986_not ; n5346
g5155 and n4977_not n5346 ; n5347
g5156 and asqrt[35] n5347 ; n5348
g5157 nor n4977 n4986 ; n5349
g5158 and asqrt[35] n5349 ; n5350
g5159 nor n4984 n5350 ; n5351
g5160 nor n5348 n5351 ; n5352
g5161 nor asqrt[43] n5333 ; n5353
g5162 and n5343_not n5353 ; n5354
g5163 nor n5352 n5354 ; n5355
g5164 nor n5345 n5355 ; n5356
g5165 and asqrt[44] n5356_not ; n5357
g5166 and n4989_not n4996 ; n5358
g5167 and n4998_not n5358 ; n5359
g5168 and asqrt[35] n5359 ; n5360
g5169 nor n4989 n4998 ; n5361
g5170 and asqrt[35] n5361 ; n5362
g5171 nor n4996 n5362 ; n5363
g5172 nor n5360 n5363 ; n5364
g5173 nor asqrt[44] n5345 ; n5365
g5174 and n5355_not n5365 ; n5366
g5175 nor n5364 n5366 ; n5367
g5176 nor n5357 n5367 ; n5368
g5177 and asqrt[45] n5368_not ; n5369
g5178 and n5008 n5010_not ; n5370
g5179 and n5001_not n5370 ; n5371
g5180 and asqrt[35] n5371 ; n5372
g5181 nor n5001 n5010 ; n5373
g5182 and asqrt[35] n5373 ; n5374
g5183 nor n5008 n5374 ; n5375
g5184 nor n5372 n5375 ; n5376
g5185 nor asqrt[45] n5357 ; n5377
g5186 and n5367_not n5377 ; n5378
g5187 nor n5376 n5378 ; n5379
g5188 nor n5369 n5379 ; n5380
g5189 and asqrt[46] n5380_not ; n5381
g5190 and n5013_not n5020 ; n5382
g5191 and n5022_not n5382 ; n5383
g5192 and asqrt[35] n5383 ; n5384
g5193 nor n5013 n5022 ; n5385
g5194 and asqrt[35] n5385 ; n5386
g5195 nor n5020 n5386 ; n5387
g5196 nor n5384 n5387 ; n5388
g5197 nor asqrt[46] n5369 ; n5389
g5198 and n5379_not n5389 ; n5390
g5199 nor n5388 n5390 ; n5391
g5200 nor n5381 n5391 ; n5392
g5201 and asqrt[47] n5392_not ; n5393
g5202 and n5032 n5034_not ; n5394
g5203 and n5025_not n5394 ; n5395
g5204 and asqrt[35] n5395 ; n5396
g5205 nor n5025 n5034 ; n5397
g5206 and asqrt[35] n5397 ; n5398
g5207 nor n5032 n5398 ; n5399
g5208 nor n5396 n5399 ; n5400
g5209 nor asqrt[47] n5381 ; n5401
g5210 and n5391_not n5401 ; n5402
g5211 nor n5400 n5402 ; n5403
g5212 nor n5393 n5403 ; n5404
g5213 and asqrt[48] n5404_not ; n5405
g5214 and n5037_not n5044 ; n5406
g5215 and n5046_not n5406 ; n5407
g5216 and asqrt[35] n5407 ; n5408
g5217 nor n5037 n5046 ; n5409
g5218 and asqrt[35] n5409 ; n5410
g5219 nor n5044 n5410 ; n5411
g5220 nor n5408 n5411 ; n5412
g5221 nor asqrt[48] n5393 ; n5413
g5222 and n5403_not n5413 ; n5414
g5223 nor n5412 n5414 ; n5415
g5224 nor n5405 n5415 ; n5416
g5225 and asqrt[49] n5416_not ; n5417
g5226 and n5056 n5058_not ; n5418
g5227 and n5049_not n5418 ; n5419
g5228 and asqrt[35] n5419 ; n5420
g5229 nor n5049 n5058 ; n5421
g5230 and asqrt[35] n5421 ; n5422
g5231 nor n5056 n5422 ; n5423
g5232 nor n5420 n5423 ; n5424
g5233 nor asqrt[49] n5405 ; n5425
g5234 and n5415_not n5425 ; n5426
g5235 nor n5424 n5426 ; n5427
g5236 nor n5417 n5427 ; n5428
g5237 and asqrt[50] n5428_not ; n5429
g5238 and n5061_not n5068 ; n5430
g5239 and n5070_not n5430 ; n5431
g5240 and asqrt[35] n5431 ; n5432
g5241 nor n5061 n5070 ; n5433
g5242 and asqrt[35] n5433 ; n5434
g5243 nor n5068 n5434 ; n5435
g5244 nor n5432 n5435 ; n5436
g5245 nor asqrt[50] n5417 ; n5437
g5246 and n5427_not n5437 ; n5438
g5247 nor n5436 n5438 ; n5439
g5248 nor n5429 n5439 ; n5440
g5249 and asqrt[51] n5440_not ; n5441
g5250 and n5080 n5082_not ; n5442
g5251 and n5073_not n5442 ; n5443
g5252 and asqrt[35] n5443 ; n5444
g5253 nor n5073 n5082 ; n5445
g5254 and asqrt[35] n5445 ; n5446
g5255 nor n5080 n5446 ; n5447
g5256 nor n5444 n5447 ; n5448
g5257 nor asqrt[51] n5429 ; n5449
g5258 and n5439_not n5449 ; n5450
g5259 nor n5448 n5450 ; n5451
g5260 nor n5441 n5451 ; n5452
g5261 and asqrt[52] n5452_not ; n5453
g5262 and n5085_not n5092 ; n5454
g5263 and n5094_not n5454 ; n5455
g5264 and asqrt[35] n5455 ; n5456
g5265 nor n5085 n5094 ; n5457
g5266 and asqrt[35] n5457 ; n5458
g5267 nor n5092 n5458 ; n5459
g5268 nor n5456 n5459 ; n5460
g5269 nor asqrt[52] n5441 ; n5461
g5270 and n5451_not n5461 ; n5462
g5271 nor n5460 n5462 ; n5463
g5272 nor n5453 n5463 ; n5464
g5273 and asqrt[53] n5464_not ; n5465
g5274 and n5104 n5106_not ; n5466
g5275 and n5097_not n5466 ; n5467
g5276 and asqrt[35] n5467 ; n5468
g5277 nor n5097 n5106 ; n5469
g5278 and asqrt[35] n5469 ; n5470
g5279 nor n5104 n5470 ; n5471
g5280 nor n5468 n5471 ; n5472
g5281 nor asqrt[53] n5453 ; n5473
g5282 and n5463_not n5473 ; n5474
g5283 nor n5472 n5474 ; n5475
g5284 nor n5465 n5475 ; n5476
g5285 and asqrt[54] n5476_not ; n5477
g5286 and n5109_not n5116 ; n5478
g5287 and n5118_not n5478 ; n5479
g5288 and asqrt[35] n5479 ; n5480
g5289 nor n5109 n5118 ; n5481
g5290 and asqrt[35] n5481 ; n5482
g5291 nor n5116 n5482 ; n5483
g5292 nor n5480 n5483 ; n5484
g5293 nor asqrt[54] n5465 ; n5485
g5294 and n5475_not n5485 ; n5486
g5295 nor n5484 n5486 ; n5487
g5296 nor n5477 n5487 ; n5488
g5297 and asqrt[55] n5488_not ; n5489
g5298 and n5128 n5130_not ; n5490
g5299 and n5121_not n5490 ; n5491
g5300 and asqrt[35] n5491 ; n5492
g5301 nor n5121 n5130 ; n5493
g5302 and asqrt[35] n5493 ; n5494
g5303 nor n5128 n5494 ; n5495
g5304 nor n5492 n5495 ; n5496
g5305 nor asqrt[55] n5477 ; n5497
g5306 and n5487_not n5497 ; n5498
g5307 nor n5496 n5498 ; n5499
g5308 nor n5489 n5499 ; n5500
g5309 and asqrt[56] n5500_not ; n5501
g5310 and n5133_not n5140 ; n5502
g5311 and n5142_not n5502 ; n5503
g5312 and asqrt[35] n5503 ; n5504
g5313 nor n5133 n5142 ; n5505
g5314 and asqrt[35] n5505 ; n5506
g5315 nor n5140 n5506 ; n5507
g5316 nor n5504 n5507 ; n5508
g5317 nor asqrt[56] n5489 ; n5509
g5318 and n5499_not n5509 ; n5510
g5319 nor n5508 n5510 ; n5511
g5320 nor n5501 n5511 ; n5512
g5321 and asqrt[57] n5512_not ; n5513
g5322 and n5152 n5154_not ; n5514
g5323 and n5145_not n5514 ; n5515
g5324 and asqrt[35] n5515 ; n5516
g5325 nor n5145 n5154 ; n5517
g5326 and asqrt[35] n5517 ; n5518
g5327 nor n5152 n5518 ; n5519
g5328 nor n5516 n5519 ; n5520
g5329 nor asqrt[57] n5501 ; n5521
g5330 and n5511_not n5521 ; n5522
g5331 nor n5520 n5522 ; n5523
g5332 nor n5513 n5523 ; n5524
g5333 and asqrt[58] n5524_not ; n5525
g5334 and n5157_not n5164 ; n5526
g5335 and n5166_not n5526 ; n5527
g5336 and asqrt[35] n5527 ; n5528
g5337 nor n5157 n5166 ; n5529
g5338 and asqrt[35] n5529 ; n5530
g5339 nor n5164 n5530 ; n5531
g5340 nor n5528 n5531 ; n5532
g5341 nor asqrt[58] n5513 ; n5533
g5342 and n5523_not n5533 ; n5534
g5343 nor n5532 n5534 ; n5535
g5344 nor n5525 n5535 ; n5536
g5345 and asqrt[59] n5536_not ; n5537
g5346 and n5176 n5178_not ; n5538
g5347 and n5169_not n5538 ; n5539
g5348 and asqrt[35] n5539 ; n5540
g5349 nor n5169 n5178 ; n5541
g5350 and asqrt[35] n5541 ; n5542
g5351 nor n5176 n5542 ; n5543
g5352 nor n5540 n5543 ; n5544
g5353 nor asqrt[59] n5525 ; n5545
g5354 and n5535_not n5545 ; n5546
g5355 nor n5544 n5546 ; n5547
g5356 nor n5537 n5547 ; n5548
g5357 and asqrt[60] n5548_not ; n5549
g5358 and n5181_not n5188 ; n5550
g5359 and n5190_not n5550 ; n5551
g5360 and asqrt[35] n5551 ; n5552
g5361 nor n5181 n5190 ; n5553
g5362 and asqrt[35] n5553 ; n5554
g5363 nor n5188 n5554 ; n5555
g5364 nor n5552 n5555 ; n5556
g5365 nor asqrt[60] n5537 ; n5557
g5366 and n5547_not n5557 ; n5558
g5367 nor n5556 n5558 ; n5559
g5368 nor n5549 n5559 ; n5560
g5369 and asqrt[61] n5560_not ; n5561
g5370 and n5200 n5202_not ; n5562
g5371 and n5193_not n5562 ; n5563
g5372 and asqrt[35] n5563 ; n5564
g5373 nor n5193 n5202 ; n5565
g5374 and asqrt[35] n5565 ; n5566
g5375 nor n5200 n5566 ; n5567
g5376 nor n5564 n5567 ; n5568
g5377 nor asqrt[61] n5549 ; n5569
g5378 and n5559_not n5569 ; n5570
g5379 nor n5568 n5570 ; n5571
g5380 nor n5561 n5571 ; n5572
g5381 and asqrt[62] n5572_not ; n5573
g5382 nor asqrt[62] n5561 ; n5574
g5383 and n5571_not n5574 ; n5575
g5384 and n5205_not n5214 ; n5576
g5385 and n5207_not n5576 ; n5577
g5386 and asqrt[35] n5577 ; n5578
g5387 nor n5205 n5207 ; n5579
g5388 and asqrt[35] n5579 ; n5580
g5389 nor n5214 n5580 ; n5581
g5390 nor n5578 n5581 ; n5582
g5391 nor n5575 n5582 ; n5583
g5392 nor n5573 n5583 ; n5584
g5393 and n5224 n5226_not ; n5585
g5394 and n5217_not n5585 ; n5586
g5395 and asqrt[35] n5586 ; n5587
g5396 nor n5217 n5226 ; n5588
g5397 and asqrt[35] n5588 ; n5589
g5398 nor n5224 n5589 ; n5590
g5399 nor n5587 n5590 ; n5591
g5400 nor n5228 n5235 ; n5592
g5401 and asqrt[35] n5592 ; n5593
g5402 nor n5243 n5593 ; n5594
g5403 and n5591_not n5594 ; n5595
g5404 and n5584_not n5595 ; n5596
g5405 nor asqrt[63] n5596 ; n5597
g5406 and n5573_not n5591 ; n5598
g5407 and n5583_not n5598 ; n5599
g5408 and n5235_not asqrt[35] ; n5600
g5409 and n5228 n5600_not ; n5601
g5410 and asqrt[63] n5592_not ; n5602
g5411 and n5601_not n5602 ; n5603
g5412 nor n5231 n5252 ; n5604
g5413 and n5234_not n5604 ; n5605
g5414 and n5247_not n5605 ; n5606
g5415 and n5243_not n5606 ; n5607
g5416 and n5241_not n5607 ; n5608
g5417 nor n5603 n5608 ; n5609
g5418 and n5599_not n5609 ; n5610
g5419 nand n5597_not n5610 ; asqrt[34]
g5420 and a[68] asqrt[34] ; n5612
g5421 nor a[66] a[67] ; n5613
g5422 and a[68]_not n5613 ; n5614
g5423 nor n5612 n5614 ; n5615
g5424 and asqrt[35] n5615_not ; n5616
g5425 nor n5252 n5614 ; n5617
g5426 and n5247_not n5617 ; n5618
g5427 and n5243_not n5618 ; n5619
g5428 and n5241_not n5619 ; n5620
g5429 and n5612_not n5620 ; n5621
g5430 and a[68]_not asqrt[34] ; n5622
g5431 and a[69] n5622_not ; n5623
g5432 and n5257 asqrt[34] ; n5624
g5433 nor n5623 n5624 ; n5625
g5434 and n5621_not n5625 ; n5626
g5435 nor n5616 n5626 ; n5627
g5436 and asqrt[36] n5627_not ; n5628
g5437 nor asqrt[36] n5616 ; n5629
g5438 and n5626_not n5629 ; n5630
g5439 and asqrt[35] n5608_not ; n5631
g5440 and n5603_not n5631 ; n5632
g5441 and n5599_not n5632 ; n5633
g5442 and n5597_not n5633 ; n5634
g5443 nor n5624 n5634 ; n5635
g5444 and a[70] n5635_not ; n5636
g5445 nor a[70] n5634 ; n5637
g5446 and n5624_not n5637 ; n5638
g5447 nor n5636 n5638 ; n5639
g5448 nor n5630 n5639 ; n5640
g5449 nor n5628 n5640 ; n5641
g5450 and asqrt[37] n5641_not ; n5642
g5451 nor n5260 n5265 ; n5643
g5452 and n5269_not n5643 ; n5644
g5453 and asqrt[34] n5644 ; n5645
g5454 and asqrt[34] n5643 ; n5646
g5455 and n5269 n5646_not ; n5647
g5456 nor n5645 n5647 ; n5648
g5457 nor asqrt[37] n5628 ; n5649
g5458 and n5640_not n5649 ; n5650
g5459 nor n5648 n5650 ; n5651
g5460 nor n5642 n5651 ; n5652
g5461 and asqrt[38] n5652_not ; n5653
g5462 and n5274_not n5283 ; n5654
g5463 and n5272_not n5654 ; n5655
g5464 and asqrt[34] n5655 ; n5656
g5465 nor n5272 n5274 ; n5657
g5466 and asqrt[34] n5657 ; n5658
g5467 nor n5283 n5658 ; n5659
g5468 nor n5656 n5659 ; n5660
g5469 nor asqrt[38] n5642 ; n5661
g5470 and n5651_not n5661 ; n5662
g5471 nor n5660 n5662 ; n5663
g5472 nor n5653 n5663 ; n5664
g5473 and asqrt[39] n5664_not ; n5665
g5474 and n5286_not n5292 ; n5666
g5475 and n5294_not n5666 ; n5667
g5476 and asqrt[34] n5667 ; n5668
g5477 nor n5286 n5294 ; n5669
g5478 and asqrt[34] n5669 ; n5670
g5479 nor n5292 n5670 ; n5671
g5480 nor n5668 n5671 ; n5672
g5481 nor asqrt[39] n5653 ; n5673
g5482 and n5663_not n5673 ; n5674
g5483 nor n5672 n5674 ; n5675
g5484 nor n5665 n5675 ; n5676
g5485 and asqrt[40] n5676_not ; n5677
g5486 and n5304 n5306_not ; n5678
g5487 and n5297_not n5678 ; n5679
g5488 and asqrt[34] n5679 ; n5680
g5489 nor n5297 n5306 ; n5681
g5490 and asqrt[34] n5681 ; n5682
g5491 nor n5304 n5682 ; n5683
g5492 nor n5680 n5683 ; n5684
g5493 nor asqrt[40] n5665 ; n5685
g5494 and n5675_not n5685 ; n5686
g5495 nor n5684 n5686 ; n5687
g5496 nor n5677 n5687 ; n5688
g5497 and asqrt[41] n5688_not ; n5689
g5498 and n5309_not n5316 ; n5690
g5499 and n5318_not n5690 ; n5691
g5500 and asqrt[34] n5691 ; n5692
g5501 nor n5309 n5318 ; n5693
g5502 and asqrt[34] n5693 ; n5694
g5503 nor n5316 n5694 ; n5695
g5504 nor n5692 n5695 ; n5696
g5505 nor asqrt[41] n5677 ; n5697
g5506 and n5687_not n5697 ; n5698
g5507 nor n5696 n5698 ; n5699
g5508 nor n5689 n5699 ; n5700
g5509 and asqrt[42] n5700_not ; n5701
g5510 and n5328 n5330_not ; n5702
g5511 and n5321_not n5702 ; n5703
g5512 and asqrt[34] n5703 ; n5704
g5513 nor n5321 n5330 ; n5705
g5514 and asqrt[34] n5705 ; n5706
g5515 nor n5328 n5706 ; n5707
g5516 nor n5704 n5707 ; n5708
g5517 nor asqrt[42] n5689 ; n5709
g5518 and n5699_not n5709 ; n5710
g5519 nor n5708 n5710 ; n5711
g5520 nor n5701 n5711 ; n5712
g5521 and asqrt[43] n5712_not ; n5713
g5522 and n5333_not n5340 ; n5714
g5523 and n5342_not n5714 ; n5715
g5524 and asqrt[34] n5715 ; n5716
g5525 nor n5333 n5342 ; n5717
g5526 and asqrt[34] n5717 ; n5718
g5527 nor n5340 n5718 ; n5719
g5528 nor n5716 n5719 ; n5720
g5529 nor asqrt[43] n5701 ; n5721
g5530 and n5711_not n5721 ; n5722
g5531 nor n5720 n5722 ; n5723
g5532 nor n5713 n5723 ; n5724
g5533 and asqrt[44] n5724_not ; n5725
g5534 and n5352 n5354_not ; n5726
g5535 and n5345_not n5726 ; n5727
g5536 and asqrt[34] n5727 ; n5728
g5537 nor n5345 n5354 ; n5729
g5538 and asqrt[34] n5729 ; n5730
g5539 nor n5352 n5730 ; n5731
g5540 nor n5728 n5731 ; n5732
g5541 nor asqrt[44] n5713 ; n5733
g5542 and n5723_not n5733 ; n5734
g5543 nor n5732 n5734 ; n5735
g5544 nor n5725 n5735 ; n5736
g5545 and asqrt[45] n5736_not ; n5737
g5546 and n5357_not n5364 ; n5738
g5547 and n5366_not n5738 ; n5739
g5548 and asqrt[34] n5739 ; n5740
g5549 nor n5357 n5366 ; n5741
g5550 and asqrt[34] n5741 ; n5742
g5551 nor n5364 n5742 ; n5743
g5552 nor n5740 n5743 ; n5744
g5553 nor asqrt[45] n5725 ; n5745
g5554 and n5735_not n5745 ; n5746
g5555 nor n5744 n5746 ; n5747
g5556 nor n5737 n5747 ; n5748
g5557 and asqrt[46] n5748_not ; n5749
g5558 and n5376 n5378_not ; n5750
g5559 and n5369_not n5750 ; n5751
g5560 and asqrt[34] n5751 ; n5752
g5561 nor n5369 n5378 ; n5753
g5562 and asqrt[34] n5753 ; n5754
g5563 nor n5376 n5754 ; n5755
g5564 nor n5752 n5755 ; n5756
g5565 nor asqrt[46] n5737 ; n5757
g5566 and n5747_not n5757 ; n5758
g5567 nor n5756 n5758 ; n5759
g5568 nor n5749 n5759 ; n5760
g5569 and asqrt[47] n5760_not ; n5761
g5570 and n5381_not n5388 ; n5762
g5571 and n5390_not n5762 ; n5763
g5572 and asqrt[34] n5763 ; n5764
g5573 nor n5381 n5390 ; n5765
g5574 and asqrt[34] n5765 ; n5766
g5575 nor n5388 n5766 ; n5767
g5576 nor n5764 n5767 ; n5768
g5577 nor asqrt[47] n5749 ; n5769
g5578 and n5759_not n5769 ; n5770
g5579 nor n5768 n5770 ; n5771
g5580 nor n5761 n5771 ; n5772
g5581 and asqrt[48] n5772_not ; n5773
g5582 and n5400 n5402_not ; n5774
g5583 and n5393_not n5774 ; n5775
g5584 and asqrt[34] n5775 ; n5776
g5585 nor n5393 n5402 ; n5777
g5586 and asqrt[34] n5777 ; n5778
g5587 nor n5400 n5778 ; n5779
g5588 nor n5776 n5779 ; n5780
g5589 nor asqrt[48] n5761 ; n5781
g5590 and n5771_not n5781 ; n5782
g5591 nor n5780 n5782 ; n5783
g5592 nor n5773 n5783 ; n5784
g5593 and asqrt[49] n5784_not ; n5785
g5594 and n5405_not n5412 ; n5786
g5595 and n5414_not n5786 ; n5787
g5596 and asqrt[34] n5787 ; n5788
g5597 nor n5405 n5414 ; n5789
g5598 and asqrt[34] n5789 ; n5790
g5599 nor n5412 n5790 ; n5791
g5600 nor n5788 n5791 ; n5792
g5601 nor asqrt[49] n5773 ; n5793
g5602 and n5783_not n5793 ; n5794
g5603 nor n5792 n5794 ; n5795
g5604 nor n5785 n5795 ; n5796
g5605 and asqrt[50] n5796_not ; n5797
g5606 and n5424 n5426_not ; n5798
g5607 and n5417_not n5798 ; n5799
g5608 and asqrt[34] n5799 ; n5800
g5609 nor n5417 n5426 ; n5801
g5610 and asqrt[34] n5801 ; n5802
g5611 nor n5424 n5802 ; n5803
g5612 nor n5800 n5803 ; n5804
g5613 nor asqrt[50] n5785 ; n5805
g5614 and n5795_not n5805 ; n5806
g5615 nor n5804 n5806 ; n5807
g5616 nor n5797 n5807 ; n5808
g5617 and asqrt[51] n5808_not ; n5809
g5618 and n5429_not n5436 ; n5810
g5619 and n5438_not n5810 ; n5811
g5620 and asqrt[34] n5811 ; n5812
g5621 nor n5429 n5438 ; n5813
g5622 and asqrt[34] n5813 ; n5814
g5623 nor n5436 n5814 ; n5815
g5624 nor n5812 n5815 ; n5816
g5625 nor asqrt[51] n5797 ; n5817
g5626 and n5807_not n5817 ; n5818
g5627 nor n5816 n5818 ; n5819
g5628 nor n5809 n5819 ; n5820
g5629 and asqrt[52] n5820_not ; n5821
g5630 and n5448 n5450_not ; n5822
g5631 and n5441_not n5822 ; n5823
g5632 and asqrt[34] n5823 ; n5824
g5633 nor n5441 n5450 ; n5825
g5634 and asqrt[34] n5825 ; n5826
g5635 nor n5448 n5826 ; n5827
g5636 nor n5824 n5827 ; n5828
g5637 nor asqrt[52] n5809 ; n5829
g5638 and n5819_not n5829 ; n5830
g5639 nor n5828 n5830 ; n5831
g5640 nor n5821 n5831 ; n5832
g5641 and asqrt[53] n5832_not ; n5833
g5642 and n5453_not n5460 ; n5834
g5643 and n5462_not n5834 ; n5835
g5644 and asqrt[34] n5835 ; n5836
g5645 nor n5453 n5462 ; n5837
g5646 and asqrt[34] n5837 ; n5838
g5647 nor n5460 n5838 ; n5839
g5648 nor n5836 n5839 ; n5840
g5649 nor asqrt[53] n5821 ; n5841
g5650 and n5831_not n5841 ; n5842
g5651 nor n5840 n5842 ; n5843
g5652 nor n5833 n5843 ; n5844
g5653 and asqrt[54] n5844_not ; n5845
g5654 and n5472 n5474_not ; n5846
g5655 and n5465_not n5846 ; n5847
g5656 and asqrt[34] n5847 ; n5848
g5657 nor n5465 n5474 ; n5849
g5658 and asqrt[34] n5849 ; n5850
g5659 nor n5472 n5850 ; n5851
g5660 nor n5848 n5851 ; n5852
g5661 nor asqrt[54] n5833 ; n5853
g5662 and n5843_not n5853 ; n5854
g5663 nor n5852 n5854 ; n5855
g5664 nor n5845 n5855 ; n5856
g5665 and asqrt[55] n5856_not ; n5857
g5666 and n5477_not n5484 ; n5858
g5667 and n5486_not n5858 ; n5859
g5668 and asqrt[34] n5859 ; n5860
g5669 nor n5477 n5486 ; n5861
g5670 and asqrt[34] n5861 ; n5862
g5671 nor n5484 n5862 ; n5863
g5672 nor n5860 n5863 ; n5864
g5673 nor asqrt[55] n5845 ; n5865
g5674 and n5855_not n5865 ; n5866
g5675 nor n5864 n5866 ; n5867
g5676 nor n5857 n5867 ; n5868
g5677 and asqrt[56] n5868_not ; n5869
g5678 and n5496 n5498_not ; n5870
g5679 and n5489_not n5870 ; n5871
g5680 and asqrt[34] n5871 ; n5872
g5681 nor n5489 n5498 ; n5873
g5682 and asqrt[34] n5873 ; n5874
g5683 nor n5496 n5874 ; n5875
g5684 nor n5872 n5875 ; n5876
g5685 nor asqrt[56] n5857 ; n5877
g5686 and n5867_not n5877 ; n5878
g5687 nor n5876 n5878 ; n5879
g5688 nor n5869 n5879 ; n5880
g5689 and asqrt[57] n5880_not ; n5881
g5690 and n5501_not n5508 ; n5882
g5691 and n5510_not n5882 ; n5883
g5692 and asqrt[34] n5883 ; n5884
g5693 nor n5501 n5510 ; n5885
g5694 and asqrt[34] n5885 ; n5886
g5695 nor n5508 n5886 ; n5887
g5696 nor n5884 n5887 ; n5888
g5697 nor asqrt[57] n5869 ; n5889
g5698 and n5879_not n5889 ; n5890
g5699 nor n5888 n5890 ; n5891
g5700 nor n5881 n5891 ; n5892
g5701 and asqrt[58] n5892_not ; n5893
g5702 and n5520 n5522_not ; n5894
g5703 and n5513_not n5894 ; n5895
g5704 and asqrt[34] n5895 ; n5896
g5705 nor n5513 n5522 ; n5897
g5706 and asqrt[34] n5897 ; n5898
g5707 nor n5520 n5898 ; n5899
g5708 nor n5896 n5899 ; n5900
g5709 nor asqrt[58] n5881 ; n5901
g5710 and n5891_not n5901 ; n5902
g5711 nor n5900 n5902 ; n5903
g5712 nor n5893 n5903 ; n5904
g5713 and asqrt[59] n5904_not ; n5905
g5714 and n5525_not n5532 ; n5906
g5715 and n5534_not n5906 ; n5907
g5716 and asqrt[34] n5907 ; n5908
g5717 nor n5525 n5534 ; n5909
g5718 and asqrt[34] n5909 ; n5910
g5719 nor n5532 n5910 ; n5911
g5720 nor n5908 n5911 ; n5912
g5721 nor asqrt[59] n5893 ; n5913
g5722 and n5903_not n5913 ; n5914
g5723 nor n5912 n5914 ; n5915
g5724 nor n5905 n5915 ; n5916
g5725 and asqrt[60] n5916_not ; n5917
g5726 and n5544 n5546_not ; n5918
g5727 and n5537_not n5918 ; n5919
g5728 and asqrt[34] n5919 ; n5920
g5729 nor n5537 n5546 ; n5921
g5730 and asqrt[34] n5921 ; n5922
g5731 nor n5544 n5922 ; n5923
g5732 nor n5920 n5923 ; n5924
g5733 nor asqrt[60] n5905 ; n5925
g5734 and n5915_not n5925 ; n5926
g5735 nor n5924 n5926 ; n5927
g5736 nor n5917 n5927 ; n5928
g5737 and asqrt[61] n5928_not ; n5929
g5738 and n5549_not n5556 ; n5930
g5739 and n5558_not n5930 ; n5931
g5740 and asqrt[34] n5931 ; n5932
g5741 nor n5549 n5558 ; n5933
g5742 and asqrt[34] n5933 ; n5934
g5743 nor n5556 n5934 ; n5935
g5744 nor n5932 n5935 ; n5936
g5745 nor asqrt[61] n5917 ; n5937
g5746 and n5927_not n5937 ; n5938
g5747 nor n5936 n5938 ; n5939
g5748 nor n5929 n5939 ; n5940
g5749 and asqrt[62] n5940_not ; n5941
g5750 and n5568 n5570_not ; n5942
g5751 and n5561_not n5942 ; n5943
g5752 and asqrt[34] n5943 ; n5944
g5753 nor n5561 n5570 ; n5945
g5754 and asqrt[34] n5945 ; n5946
g5755 nor n5568 n5946 ; n5947
g5756 nor n5944 n5947 ; n5948
g5757 nor asqrt[62] n5929 ; n5949
g5758 and n5939_not n5949 ; n5950
g5759 nor n5948 n5950 ; n5951
g5760 nor n5941 n5951 ; n5952
g5761 and n5573_not n5582 ; n5953
g5762 and n5575_not n5953 ; n5954
g5763 and asqrt[34] n5954 ; n5955
g5764 nor n5573 n5575 ; n5956
g5765 and asqrt[34] n5956 ; n5957
g5766 nor n5582 n5957 ; n5958
g5767 nor n5955 n5958 ; n5959
g5768 nor n5584 n5591 ; n5960
g5769 and asqrt[34] n5960 ; n5961
g5770 nor n5599 n5961 ; n5962
g5771 and n5959_not n5962 ; n5963
g5772 and n5952_not n5963 ; n5964
g5773 nor asqrt[63] n5964 ; n5965
g5774 and n5941_not n5959 ; n5966
g5775 and n5951_not n5966 ; n5967
g5776 and n5591_not asqrt[34] ; n5968
g5777 and n5584 n5968_not ; n5969
g5778 and asqrt[63] n5960_not ; n5970
g5779 and n5969_not n5970 ; n5971
g5780 nor n5587 n5608 ; n5972
g5781 and n5590_not n5972 ; n5973
g5782 and n5603_not n5973 ; n5974
g5783 and n5599_not n5974 ; n5975
g5784 and n5597_not n5975 ; n5976
g5785 nor n5971 n5976 ; n5977
g5786 and n5967_not n5977 ; n5978
g5787 nand n5965_not n5978 ; asqrt[33]
g5788 and a[66] asqrt[33] ; n5980
g5789 nor a[64] a[65] ; n5981
g5790 and a[66]_not n5981 ; n5982
g5791 nor n5980 n5982 ; n5983
g5792 and asqrt[34] n5983_not ; n5984
g5793 nor n5608 n5982 ; n5985
g5794 and n5603_not n5985 ; n5986
g5795 and n5599_not n5986 ; n5987
g5796 and n5597_not n5987 ; n5988
g5797 and n5980_not n5988 ; n5989
g5798 and a[66]_not asqrt[33] ; n5990
g5799 and a[67] n5990_not ; n5991
g5800 and n5613 asqrt[33] ; n5992
g5801 nor n5991 n5992 ; n5993
g5802 and n5989_not n5993 ; n5994
g5803 nor n5984 n5994 ; n5995
g5804 and asqrt[35] n5995_not ; n5996
g5805 nor asqrt[35] n5984 ; n5997
g5806 and n5994_not n5997 ; n5998
g5807 and asqrt[34] n5976_not ; n5999
g5808 and n5971_not n5999 ; n6000
g5809 and n5967_not n6000 ; n6001
g5810 and n5965_not n6001 ; n6002
g5811 nor n5992 n6002 ; n6003
g5812 and a[68] n6003_not ; n6004
g5813 nor a[68] n6002 ; n6005
g5814 and n5992_not n6005 ; n6006
g5815 nor n6004 n6006 ; n6007
g5816 nor n5998 n6007 ; n6008
g5817 nor n5996 n6008 ; n6009
g5818 and asqrt[36] n6009_not ; n6010
g5819 nor n5616 n5621 ; n6011
g5820 and n5625_not n6011 ; n6012
g5821 and asqrt[33] n6012 ; n6013
g5822 and asqrt[33] n6011 ; n6014
g5823 and n5625 n6014_not ; n6015
g5824 nor n6013 n6015 ; n6016
g5825 nor asqrt[36] n5996 ; n6017
g5826 and n6008_not n6017 ; n6018
g5827 nor n6016 n6018 ; n6019
g5828 nor n6010 n6019 ; n6020
g5829 and asqrt[37] n6020_not ; n6021
g5830 and n5630_not n5639 ; n6022
g5831 and n5628_not n6022 ; n6023
g5832 and asqrt[33] n6023 ; n6024
g5833 nor n5628 n5630 ; n6025
g5834 and asqrt[33] n6025 ; n6026
g5835 nor n5639 n6026 ; n6027
g5836 nor n6024 n6027 ; n6028
g5837 nor asqrt[37] n6010 ; n6029
g5838 and n6019_not n6029 ; n6030
g5839 nor n6028 n6030 ; n6031
g5840 nor n6021 n6031 ; n6032
g5841 and asqrt[38] n6032_not ; n6033
g5842 and n5642_not n5648 ; n6034
g5843 and n5650_not n6034 ; n6035
g5844 and asqrt[33] n6035 ; n6036
g5845 nor n5642 n5650 ; n6037
g5846 and asqrt[33] n6037 ; n6038
g5847 nor n5648 n6038 ; n6039
g5848 nor n6036 n6039 ; n6040
g5849 nor asqrt[38] n6021 ; n6041
g5850 and n6031_not n6041 ; n6042
g5851 nor n6040 n6042 ; n6043
g5852 nor n6033 n6043 ; n6044
g5853 and asqrt[39] n6044_not ; n6045
g5854 and n5660 n5662_not ; n6046
g5855 and n5653_not n6046 ; n6047
g5856 and asqrt[33] n6047 ; n6048
g5857 nor n5653 n5662 ; n6049
g5858 and asqrt[33] n6049 ; n6050
g5859 nor n5660 n6050 ; n6051
g5860 nor n6048 n6051 ; n6052
g5861 nor asqrt[39] n6033 ; n6053
g5862 and n6043_not n6053 ; n6054
g5863 nor n6052 n6054 ; n6055
g5864 nor n6045 n6055 ; n6056
g5865 and asqrt[40] n6056_not ; n6057
g5866 and n5665_not n5672 ; n6058
g5867 and n5674_not n6058 ; n6059
g5868 and asqrt[33] n6059 ; n6060
g5869 nor n5665 n5674 ; n6061
g5870 and asqrt[33] n6061 ; n6062
g5871 nor n5672 n6062 ; n6063
g5872 nor n6060 n6063 ; n6064
g5873 nor asqrt[40] n6045 ; n6065
g5874 and n6055_not n6065 ; n6066
g5875 nor n6064 n6066 ; n6067
g5876 nor n6057 n6067 ; n6068
g5877 and asqrt[41] n6068_not ; n6069
g5878 and n5684 n5686_not ; n6070
g5879 and n5677_not n6070 ; n6071
g5880 and asqrt[33] n6071 ; n6072
g5881 nor n5677 n5686 ; n6073
g5882 and asqrt[33] n6073 ; n6074
g5883 nor n5684 n6074 ; n6075
g5884 nor n6072 n6075 ; n6076
g5885 nor asqrt[41] n6057 ; n6077
g5886 and n6067_not n6077 ; n6078
g5887 nor n6076 n6078 ; n6079
g5888 nor n6069 n6079 ; n6080
g5889 and asqrt[42] n6080_not ; n6081
g5890 and n5689_not n5696 ; n6082
g5891 and n5698_not n6082 ; n6083
g5892 and asqrt[33] n6083 ; n6084
g5893 nor n5689 n5698 ; n6085
g5894 and asqrt[33] n6085 ; n6086
g5895 nor n5696 n6086 ; n6087
g5896 nor n6084 n6087 ; n6088
g5897 nor asqrt[42] n6069 ; n6089
g5898 and n6079_not n6089 ; n6090
g5899 nor n6088 n6090 ; n6091
g5900 nor n6081 n6091 ; n6092
g5901 and asqrt[43] n6092_not ; n6093
g5902 and n5708 n5710_not ; n6094
g5903 and n5701_not n6094 ; n6095
g5904 and asqrt[33] n6095 ; n6096
g5905 nor n5701 n5710 ; n6097
g5906 and asqrt[33] n6097 ; n6098
g5907 nor n5708 n6098 ; n6099
g5908 nor n6096 n6099 ; n6100
g5909 nor asqrt[43] n6081 ; n6101
g5910 and n6091_not n6101 ; n6102
g5911 nor n6100 n6102 ; n6103
g5912 nor n6093 n6103 ; n6104
g5913 and asqrt[44] n6104_not ; n6105
g5914 and n5713_not n5720 ; n6106
g5915 and n5722_not n6106 ; n6107
g5916 and asqrt[33] n6107 ; n6108
g5917 nor n5713 n5722 ; n6109
g5918 and asqrt[33] n6109 ; n6110
g5919 nor n5720 n6110 ; n6111
g5920 nor n6108 n6111 ; n6112
g5921 nor asqrt[44] n6093 ; n6113
g5922 and n6103_not n6113 ; n6114
g5923 nor n6112 n6114 ; n6115
g5924 nor n6105 n6115 ; n6116
g5925 and asqrt[45] n6116_not ; n6117
g5926 and n5732 n5734_not ; n6118
g5927 and n5725_not n6118 ; n6119
g5928 and asqrt[33] n6119 ; n6120
g5929 nor n5725 n5734 ; n6121
g5930 and asqrt[33] n6121 ; n6122
g5931 nor n5732 n6122 ; n6123
g5932 nor n6120 n6123 ; n6124
g5933 nor asqrt[45] n6105 ; n6125
g5934 and n6115_not n6125 ; n6126
g5935 nor n6124 n6126 ; n6127
g5936 nor n6117 n6127 ; n6128
g5937 and asqrt[46] n6128_not ; n6129
g5938 and n5737_not n5744 ; n6130
g5939 and n5746_not n6130 ; n6131
g5940 and asqrt[33] n6131 ; n6132
g5941 nor n5737 n5746 ; n6133
g5942 and asqrt[33] n6133 ; n6134
g5943 nor n5744 n6134 ; n6135
g5944 nor n6132 n6135 ; n6136
g5945 nor asqrt[46] n6117 ; n6137
g5946 and n6127_not n6137 ; n6138
g5947 nor n6136 n6138 ; n6139
g5948 nor n6129 n6139 ; n6140
g5949 and asqrt[47] n6140_not ; n6141
g5950 and n5756 n5758_not ; n6142
g5951 and n5749_not n6142 ; n6143
g5952 and asqrt[33] n6143 ; n6144
g5953 nor n5749 n5758 ; n6145
g5954 and asqrt[33] n6145 ; n6146
g5955 nor n5756 n6146 ; n6147
g5956 nor n6144 n6147 ; n6148
g5957 nor asqrt[47] n6129 ; n6149
g5958 and n6139_not n6149 ; n6150
g5959 nor n6148 n6150 ; n6151
g5960 nor n6141 n6151 ; n6152
g5961 and asqrt[48] n6152_not ; n6153
g5962 and n5761_not n5768 ; n6154
g5963 and n5770_not n6154 ; n6155
g5964 and asqrt[33] n6155 ; n6156
g5965 nor n5761 n5770 ; n6157
g5966 and asqrt[33] n6157 ; n6158
g5967 nor n5768 n6158 ; n6159
g5968 nor n6156 n6159 ; n6160
g5969 nor asqrt[48] n6141 ; n6161
g5970 and n6151_not n6161 ; n6162
g5971 nor n6160 n6162 ; n6163
g5972 nor n6153 n6163 ; n6164
g5973 and asqrt[49] n6164_not ; n6165
g5974 and n5780 n5782_not ; n6166
g5975 and n5773_not n6166 ; n6167
g5976 and asqrt[33] n6167 ; n6168
g5977 nor n5773 n5782 ; n6169
g5978 and asqrt[33] n6169 ; n6170
g5979 nor n5780 n6170 ; n6171
g5980 nor n6168 n6171 ; n6172
g5981 nor asqrt[49] n6153 ; n6173
g5982 and n6163_not n6173 ; n6174
g5983 nor n6172 n6174 ; n6175
g5984 nor n6165 n6175 ; n6176
g5985 and asqrt[50] n6176_not ; n6177
g5986 and n5785_not n5792 ; n6178
g5987 and n5794_not n6178 ; n6179
g5988 and asqrt[33] n6179 ; n6180
g5989 nor n5785 n5794 ; n6181
g5990 and asqrt[33] n6181 ; n6182
g5991 nor n5792 n6182 ; n6183
g5992 nor n6180 n6183 ; n6184
g5993 nor asqrt[50] n6165 ; n6185
g5994 and n6175_not n6185 ; n6186
g5995 nor n6184 n6186 ; n6187
g5996 nor n6177 n6187 ; n6188
g5997 and asqrt[51] n6188_not ; n6189
g5998 and n5804 n5806_not ; n6190
g5999 and n5797_not n6190 ; n6191
g6000 and asqrt[33] n6191 ; n6192
g6001 nor n5797 n5806 ; n6193
g6002 and asqrt[33] n6193 ; n6194
g6003 nor n5804 n6194 ; n6195
g6004 nor n6192 n6195 ; n6196
g6005 nor asqrt[51] n6177 ; n6197
g6006 and n6187_not n6197 ; n6198
g6007 nor n6196 n6198 ; n6199
g6008 nor n6189 n6199 ; n6200
g6009 and asqrt[52] n6200_not ; n6201
g6010 and n5809_not n5816 ; n6202
g6011 and n5818_not n6202 ; n6203
g6012 and asqrt[33] n6203 ; n6204
g6013 nor n5809 n5818 ; n6205
g6014 and asqrt[33] n6205 ; n6206
g6015 nor n5816 n6206 ; n6207
g6016 nor n6204 n6207 ; n6208
g6017 nor asqrt[52] n6189 ; n6209
g6018 and n6199_not n6209 ; n6210
g6019 nor n6208 n6210 ; n6211
g6020 nor n6201 n6211 ; n6212
g6021 and asqrt[53] n6212_not ; n6213
g6022 and n5828 n5830_not ; n6214
g6023 and n5821_not n6214 ; n6215
g6024 and asqrt[33] n6215 ; n6216
g6025 nor n5821 n5830 ; n6217
g6026 and asqrt[33] n6217 ; n6218
g6027 nor n5828 n6218 ; n6219
g6028 nor n6216 n6219 ; n6220
g6029 nor asqrt[53] n6201 ; n6221
g6030 and n6211_not n6221 ; n6222
g6031 nor n6220 n6222 ; n6223
g6032 nor n6213 n6223 ; n6224
g6033 and asqrt[54] n6224_not ; n6225
g6034 and n5833_not n5840 ; n6226
g6035 and n5842_not n6226 ; n6227
g6036 and asqrt[33] n6227 ; n6228
g6037 nor n5833 n5842 ; n6229
g6038 and asqrt[33] n6229 ; n6230
g6039 nor n5840 n6230 ; n6231
g6040 nor n6228 n6231 ; n6232
g6041 nor asqrt[54] n6213 ; n6233
g6042 and n6223_not n6233 ; n6234
g6043 nor n6232 n6234 ; n6235
g6044 nor n6225 n6235 ; n6236
g6045 and asqrt[55] n6236_not ; n6237
g6046 and n5852 n5854_not ; n6238
g6047 and n5845_not n6238 ; n6239
g6048 and asqrt[33] n6239 ; n6240
g6049 nor n5845 n5854 ; n6241
g6050 and asqrt[33] n6241 ; n6242
g6051 nor n5852 n6242 ; n6243
g6052 nor n6240 n6243 ; n6244
g6053 nor asqrt[55] n6225 ; n6245
g6054 and n6235_not n6245 ; n6246
g6055 nor n6244 n6246 ; n6247
g6056 nor n6237 n6247 ; n6248
g6057 and asqrt[56] n6248_not ; n6249
g6058 and n5857_not n5864 ; n6250
g6059 and n5866_not n6250 ; n6251
g6060 and asqrt[33] n6251 ; n6252
g6061 nor n5857 n5866 ; n6253
g6062 and asqrt[33] n6253 ; n6254
g6063 nor n5864 n6254 ; n6255
g6064 nor n6252 n6255 ; n6256
g6065 nor asqrt[56] n6237 ; n6257
g6066 and n6247_not n6257 ; n6258
g6067 nor n6256 n6258 ; n6259
g6068 nor n6249 n6259 ; n6260
g6069 and asqrt[57] n6260_not ; n6261
g6070 and n5876 n5878_not ; n6262
g6071 and n5869_not n6262 ; n6263
g6072 and asqrt[33] n6263 ; n6264
g6073 nor n5869 n5878 ; n6265
g6074 and asqrt[33] n6265 ; n6266
g6075 nor n5876 n6266 ; n6267
g6076 nor n6264 n6267 ; n6268
g6077 nor asqrt[57] n6249 ; n6269
g6078 and n6259_not n6269 ; n6270
g6079 nor n6268 n6270 ; n6271
g6080 nor n6261 n6271 ; n6272
g6081 and asqrt[58] n6272_not ; n6273
g6082 and n5881_not n5888 ; n6274
g6083 and n5890_not n6274 ; n6275
g6084 and asqrt[33] n6275 ; n6276
g6085 nor n5881 n5890 ; n6277
g6086 and asqrt[33] n6277 ; n6278
g6087 nor n5888 n6278 ; n6279
g6088 nor n6276 n6279 ; n6280
g6089 nor asqrt[58] n6261 ; n6281
g6090 and n6271_not n6281 ; n6282
g6091 nor n6280 n6282 ; n6283
g6092 nor n6273 n6283 ; n6284
g6093 and asqrt[59] n6284_not ; n6285
g6094 and n5900 n5902_not ; n6286
g6095 and n5893_not n6286 ; n6287
g6096 and asqrt[33] n6287 ; n6288
g6097 nor n5893 n5902 ; n6289
g6098 and asqrt[33] n6289 ; n6290
g6099 nor n5900 n6290 ; n6291
g6100 nor n6288 n6291 ; n6292
g6101 nor asqrt[59] n6273 ; n6293
g6102 and n6283_not n6293 ; n6294
g6103 nor n6292 n6294 ; n6295
g6104 nor n6285 n6295 ; n6296
g6105 and asqrt[60] n6296_not ; n6297
g6106 and n5905_not n5912 ; n6298
g6107 and n5914_not n6298 ; n6299
g6108 and asqrt[33] n6299 ; n6300
g6109 nor n5905 n5914 ; n6301
g6110 and asqrt[33] n6301 ; n6302
g6111 nor n5912 n6302 ; n6303
g6112 nor n6300 n6303 ; n6304
g6113 nor asqrt[60] n6285 ; n6305
g6114 and n6295_not n6305 ; n6306
g6115 nor n6304 n6306 ; n6307
g6116 nor n6297 n6307 ; n6308
g6117 and asqrt[61] n6308_not ; n6309
g6118 and n5924 n5926_not ; n6310
g6119 and n5917_not n6310 ; n6311
g6120 and asqrt[33] n6311 ; n6312
g6121 nor n5917 n5926 ; n6313
g6122 and asqrt[33] n6313 ; n6314
g6123 nor n5924 n6314 ; n6315
g6124 nor n6312 n6315 ; n6316
g6125 nor asqrt[61] n6297 ; n6317
g6126 and n6307_not n6317 ; n6318
g6127 nor n6316 n6318 ; n6319
g6128 nor n6309 n6319 ; n6320
g6129 and asqrt[62] n6320_not ; n6321
g6130 and n5929_not n5936 ; n6322
g6131 and n5938_not n6322 ; n6323
g6132 and asqrt[33] n6323 ; n6324
g6133 nor n5929 n5938 ; n6325
g6134 and asqrt[33] n6325 ; n6326
g6135 nor n5936 n6326 ; n6327
g6136 nor n6324 n6327 ; n6328
g6137 nor asqrt[62] n6309 ; n6329
g6138 and n6319_not n6329 ; n6330
g6139 nor n6328 n6330 ; n6331
g6140 nor n6321 n6331 ; n6332
g6141 and n5948 n5950_not ; n6333
g6142 and n5941_not n6333 ; n6334
g6143 and asqrt[33] n6334 ; n6335
g6144 nor n5941 n5950 ; n6336
g6145 and asqrt[33] n6336 ; n6337
g6146 nor n5948 n6337 ; n6338
g6147 nor n6335 n6338 ; n6339
g6148 nor n5952 n5959 ; n6340
g6149 and asqrt[33] n6340 ; n6341
g6150 nor n5967 n6341 ; n6342
g6151 and n6339_not n6342 ; n6343
g6152 and n6332_not n6343 ; n6344
g6153 nor asqrt[63] n6344 ; n6345
g6154 and n6321_not n6339 ; n6346
g6155 and n6331_not n6346 ; n6347
g6156 and n5959_not asqrt[33] ; n6348
g6157 and n5952 n6348_not ; n6349
g6158 and asqrt[63] n6340_not ; n6350
g6159 and n6349_not n6350 ; n6351
g6160 nor n5955 n5976 ; n6352
g6161 and n5958_not n6352 ; n6353
g6162 and n5971_not n6353 ; n6354
g6163 and n5967_not n6354 ; n6355
g6164 and n5965_not n6355 ; n6356
g6165 nor n6351 n6356 ; n6357
g6166 and n6347_not n6357 ; n6358
g6167 nand n6345_not n6358 ; asqrt[32]
g6168 and a[64] asqrt[32] ; n6360
g6169 nor a[62] a[63] ; n6361
g6170 and a[64]_not n6361 ; n6362
g6171 nor n6360 n6362 ; n6363
g6172 and asqrt[33] n6363_not ; n6364
g6173 and a[64]_not asqrt[32] ; n6365
g6174 and a[65] n6365_not ; n6366
g6175 and n5981 asqrt[32] ; n6367
g6176 nor n6366 n6367 ; n6368
g6177 nor n5976 n6362 ; n6369
g6178 and n5971_not n6369 ; n6370
g6179 and n5967_not n6370 ; n6371
g6180 and n5965_not n6371 ; n6372
g6181 and n6360_not n6372 ; n6373
g6182 and n6368 n6373_not ; n6374
g6183 nor n6364 n6374 ; n6375
g6184 and asqrt[34] n6375_not ; n6376
g6185 nor asqrt[34] n6364 ; n6377
g6186 and n6374_not n6377 ; n6378
g6187 and asqrt[33] n6356_not ; n6379
g6188 and n6351_not n6379 ; n6380
g6189 and n6347_not n6380 ; n6381
g6190 and n6345_not n6381 ; n6382
g6191 nor n6367 n6382 ; n6383
g6192 and a[66] n6383_not ; n6384
g6193 nor a[66] n6382 ; n6385
g6194 and n6367_not n6385 ; n6386
g6195 nor n6384 n6386 ; n6387
g6196 nor n6378 n6387 ; n6388
g6197 nor n6376 n6388 ; n6389
g6198 and asqrt[35] n6389_not ; n6390
g6199 nor n5984 n5989 ; n6391
g6200 and n5993_not n6391 ; n6392
g6201 and asqrt[32] n6392 ; n6393
g6202 and asqrt[32] n6391 ; n6394
g6203 and n5993 n6394_not ; n6395
g6204 nor n6393 n6395 ; n6396
g6205 nor asqrt[35] n6376 ; n6397
g6206 and n6388_not n6397 ; n6398
g6207 nor n6396 n6398 ; n6399
g6208 nor n6390 n6399 ; n6400
g6209 and asqrt[36] n6400_not ; n6401
g6210 and n5998_not n6007 ; n6402
g6211 and n5996_not n6402 ; n6403
g6212 and asqrt[32] n6403 ; n6404
g6213 nor n5996 n5998 ; n6405
g6214 and asqrt[32] n6405 ; n6406
g6215 nor n6007 n6406 ; n6407
g6216 nor n6404 n6407 ; n6408
g6217 nor asqrt[36] n6390 ; n6409
g6218 and n6399_not n6409 ; n6410
g6219 nor n6408 n6410 ; n6411
g6220 nor n6401 n6411 ; n6412
g6221 and asqrt[37] n6412_not ; n6413
g6222 and n6010_not n6016 ; n6414
g6223 and n6018_not n6414 ; n6415
g6224 and asqrt[32] n6415 ; n6416
g6225 nor n6010 n6018 ; n6417
g6226 and asqrt[32] n6417 ; n6418
g6227 nor n6016 n6418 ; n6419
g6228 nor n6416 n6419 ; n6420
g6229 nor asqrt[37] n6401 ; n6421
g6230 and n6411_not n6421 ; n6422
g6231 nor n6420 n6422 ; n6423
g6232 nor n6413 n6423 ; n6424
g6233 and asqrt[38] n6424_not ; n6425
g6234 and n6028 n6030_not ; n6426
g6235 and n6021_not n6426 ; n6427
g6236 and asqrt[32] n6427 ; n6428
g6237 nor n6021 n6030 ; n6429
g6238 and asqrt[32] n6429 ; n6430
g6239 nor n6028 n6430 ; n6431
g6240 nor n6428 n6431 ; n6432
g6241 nor asqrt[38] n6413 ; n6433
g6242 and n6423_not n6433 ; n6434
g6243 nor n6432 n6434 ; n6435
g6244 nor n6425 n6435 ; n6436
g6245 and asqrt[39] n6436_not ; n6437
g6246 and n6033_not n6040 ; n6438
g6247 and n6042_not n6438 ; n6439
g6248 and asqrt[32] n6439 ; n6440
g6249 nor n6033 n6042 ; n6441
g6250 and asqrt[32] n6441 ; n6442
g6251 nor n6040 n6442 ; n6443
g6252 nor n6440 n6443 ; n6444
g6253 nor asqrt[39] n6425 ; n6445
g6254 and n6435_not n6445 ; n6446
g6255 nor n6444 n6446 ; n6447
g6256 nor n6437 n6447 ; n6448
g6257 and asqrt[40] n6448_not ; n6449
g6258 and n6052 n6054_not ; n6450
g6259 and n6045_not n6450 ; n6451
g6260 and asqrt[32] n6451 ; n6452
g6261 nor n6045 n6054 ; n6453
g6262 and asqrt[32] n6453 ; n6454
g6263 nor n6052 n6454 ; n6455
g6264 nor n6452 n6455 ; n6456
g6265 nor asqrt[40] n6437 ; n6457
g6266 and n6447_not n6457 ; n6458
g6267 nor n6456 n6458 ; n6459
g6268 nor n6449 n6459 ; n6460
g6269 and asqrt[41] n6460_not ; n6461
g6270 and n6057_not n6064 ; n6462
g6271 and n6066_not n6462 ; n6463
g6272 and asqrt[32] n6463 ; n6464
g6273 nor n6057 n6066 ; n6465
g6274 and asqrt[32] n6465 ; n6466
g6275 nor n6064 n6466 ; n6467
g6276 nor n6464 n6467 ; n6468
g6277 nor asqrt[41] n6449 ; n6469
g6278 and n6459_not n6469 ; n6470
g6279 nor n6468 n6470 ; n6471
g6280 nor n6461 n6471 ; n6472
g6281 and asqrt[42] n6472_not ; n6473
g6282 and n6076 n6078_not ; n6474
g6283 and n6069_not n6474 ; n6475
g6284 and asqrt[32] n6475 ; n6476
g6285 nor n6069 n6078 ; n6477
g6286 and asqrt[32] n6477 ; n6478
g6287 nor n6076 n6478 ; n6479
g6288 nor n6476 n6479 ; n6480
g6289 nor asqrt[42] n6461 ; n6481
g6290 and n6471_not n6481 ; n6482
g6291 nor n6480 n6482 ; n6483
g6292 nor n6473 n6483 ; n6484
g6293 and asqrt[43] n6484_not ; n6485
g6294 and n6081_not n6088 ; n6486
g6295 and n6090_not n6486 ; n6487
g6296 and asqrt[32] n6487 ; n6488
g6297 nor n6081 n6090 ; n6489
g6298 and asqrt[32] n6489 ; n6490
g6299 nor n6088 n6490 ; n6491
g6300 nor n6488 n6491 ; n6492
g6301 nor asqrt[43] n6473 ; n6493
g6302 and n6483_not n6493 ; n6494
g6303 nor n6492 n6494 ; n6495
g6304 nor n6485 n6495 ; n6496
g6305 and asqrt[44] n6496_not ; n6497
g6306 and n6100 n6102_not ; n6498
g6307 and n6093_not n6498 ; n6499
g6308 and asqrt[32] n6499 ; n6500
g6309 nor n6093 n6102 ; n6501
g6310 and asqrt[32] n6501 ; n6502
g6311 nor n6100 n6502 ; n6503
g6312 nor n6500 n6503 ; n6504
g6313 nor asqrt[44] n6485 ; n6505
g6314 and n6495_not n6505 ; n6506
g6315 nor n6504 n6506 ; n6507
g6316 nor n6497 n6507 ; n6508
g6317 and asqrt[45] n6508_not ; n6509
g6318 and n6105_not n6112 ; n6510
g6319 and n6114_not n6510 ; n6511
g6320 and asqrt[32] n6511 ; n6512
g6321 nor n6105 n6114 ; n6513
g6322 and asqrt[32] n6513 ; n6514
g6323 nor n6112 n6514 ; n6515
g6324 nor n6512 n6515 ; n6516
g6325 nor asqrt[45] n6497 ; n6517
g6326 and n6507_not n6517 ; n6518
g6327 nor n6516 n6518 ; n6519
g6328 nor n6509 n6519 ; n6520
g6329 and asqrt[46] n6520_not ; n6521
g6330 and n6124 n6126_not ; n6522
g6331 and n6117_not n6522 ; n6523
g6332 and asqrt[32] n6523 ; n6524
g6333 nor n6117 n6126 ; n6525
g6334 and asqrt[32] n6525 ; n6526
g6335 nor n6124 n6526 ; n6527
g6336 nor n6524 n6527 ; n6528
g6337 nor asqrt[46] n6509 ; n6529
g6338 and n6519_not n6529 ; n6530
g6339 nor n6528 n6530 ; n6531
g6340 nor n6521 n6531 ; n6532
g6341 and asqrt[47] n6532_not ; n6533
g6342 and n6129_not n6136 ; n6534
g6343 and n6138_not n6534 ; n6535
g6344 and asqrt[32] n6535 ; n6536
g6345 nor n6129 n6138 ; n6537
g6346 and asqrt[32] n6537 ; n6538
g6347 nor n6136 n6538 ; n6539
g6348 nor n6536 n6539 ; n6540
g6349 nor asqrt[47] n6521 ; n6541
g6350 and n6531_not n6541 ; n6542
g6351 nor n6540 n6542 ; n6543
g6352 nor n6533 n6543 ; n6544
g6353 and asqrt[48] n6544_not ; n6545
g6354 and n6148 n6150_not ; n6546
g6355 and n6141_not n6546 ; n6547
g6356 and asqrt[32] n6547 ; n6548
g6357 nor n6141 n6150 ; n6549
g6358 and asqrt[32] n6549 ; n6550
g6359 nor n6148 n6550 ; n6551
g6360 nor n6548 n6551 ; n6552
g6361 nor asqrt[48] n6533 ; n6553
g6362 and n6543_not n6553 ; n6554
g6363 nor n6552 n6554 ; n6555
g6364 nor n6545 n6555 ; n6556
g6365 and asqrt[49] n6556_not ; n6557
g6366 and n6153_not n6160 ; n6558
g6367 and n6162_not n6558 ; n6559
g6368 and asqrt[32] n6559 ; n6560
g6369 nor n6153 n6162 ; n6561
g6370 and asqrt[32] n6561 ; n6562
g6371 nor n6160 n6562 ; n6563
g6372 nor n6560 n6563 ; n6564
g6373 nor asqrt[49] n6545 ; n6565
g6374 and n6555_not n6565 ; n6566
g6375 nor n6564 n6566 ; n6567
g6376 nor n6557 n6567 ; n6568
g6377 and asqrt[50] n6568_not ; n6569
g6378 and n6172 n6174_not ; n6570
g6379 and n6165_not n6570 ; n6571
g6380 and asqrt[32] n6571 ; n6572
g6381 nor n6165 n6174 ; n6573
g6382 and asqrt[32] n6573 ; n6574
g6383 nor n6172 n6574 ; n6575
g6384 nor n6572 n6575 ; n6576
g6385 nor asqrt[50] n6557 ; n6577
g6386 and n6567_not n6577 ; n6578
g6387 nor n6576 n6578 ; n6579
g6388 nor n6569 n6579 ; n6580
g6389 and asqrt[51] n6580_not ; n6581
g6390 and n6177_not n6184 ; n6582
g6391 and n6186_not n6582 ; n6583
g6392 and asqrt[32] n6583 ; n6584
g6393 nor n6177 n6186 ; n6585
g6394 and asqrt[32] n6585 ; n6586
g6395 nor n6184 n6586 ; n6587
g6396 nor n6584 n6587 ; n6588
g6397 nor asqrt[51] n6569 ; n6589
g6398 and n6579_not n6589 ; n6590
g6399 nor n6588 n6590 ; n6591
g6400 nor n6581 n6591 ; n6592
g6401 and asqrt[52] n6592_not ; n6593
g6402 and n6196 n6198_not ; n6594
g6403 and n6189_not n6594 ; n6595
g6404 and asqrt[32] n6595 ; n6596
g6405 nor n6189 n6198 ; n6597
g6406 and asqrt[32] n6597 ; n6598
g6407 nor n6196 n6598 ; n6599
g6408 nor n6596 n6599 ; n6600
g6409 nor asqrt[52] n6581 ; n6601
g6410 and n6591_not n6601 ; n6602
g6411 nor n6600 n6602 ; n6603
g6412 nor n6593 n6603 ; n6604
g6413 and asqrt[53] n6604_not ; n6605
g6414 and n6201_not n6208 ; n6606
g6415 and n6210_not n6606 ; n6607
g6416 and asqrt[32] n6607 ; n6608
g6417 nor n6201 n6210 ; n6609
g6418 and asqrt[32] n6609 ; n6610
g6419 nor n6208 n6610 ; n6611
g6420 nor n6608 n6611 ; n6612
g6421 nor asqrt[53] n6593 ; n6613
g6422 and n6603_not n6613 ; n6614
g6423 nor n6612 n6614 ; n6615
g6424 nor n6605 n6615 ; n6616
g6425 and asqrt[54] n6616_not ; n6617
g6426 and n6220 n6222_not ; n6618
g6427 and n6213_not n6618 ; n6619
g6428 and asqrt[32] n6619 ; n6620
g6429 nor n6213 n6222 ; n6621
g6430 and asqrt[32] n6621 ; n6622
g6431 nor n6220 n6622 ; n6623
g6432 nor n6620 n6623 ; n6624
g6433 nor asqrt[54] n6605 ; n6625
g6434 and n6615_not n6625 ; n6626
g6435 nor n6624 n6626 ; n6627
g6436 nor n6617 n6627 ; n6628
g6437 and asqrt[55] n6628_not ; n6629
g6438 and n6225_not n6232 ; n6630
g6439 and n6234_not n6630 ; n6631
g6440 and asqrt[32] n6631 ; n6632
g6441 nor n6225 n6234 ; n6633
g6442 and asqrt[32] n6633 ; n6634
g6443 nor n6232 n6634 ; n6635
g6444 nor n6632 n6635 ; n6636
g6445 nor asqrt[55] n6617 ; n6637
g6446 and n6627_not n6637 ; n6638
g6447 nor n6636 n6638 ; n6639
g6448 nor n6629 n6639 ; n6640
g6449 and asqrt[56] n6640_not ; n6641
g6450 and n6244 n6246_not ; n6642
g6451 and n6237_not n6642 ; n6643
g6452 and asqrt[32] n6643 ; n6644
g6453 nor n6237 n6246 ; n6645
g6454 and asqrt[32] n6645 ; n6646
g6455 nor n6244 n6646 ; n6647
g6456 nor n6644 n6647 ; n6648
g6457 nor asqrt[56] n6629 ; n6649
g6458 and n6639_not n6649 ; n6650
g6459 nor n6648 n6650 ; n6651
g6460 nor n6641 n6651 ; n6652
g6461 and asqrt[57] n6652_not ; n6653
g6462 and n6249_not n6256 ; n6654
g6463 and n6258_not n6654 ; n6655
g6464 and asqrt[32] n6655 ; n6656
g6465 nor n6249 n6258 ; n6657
g6466 and asqrt[32] n6657 ; n6658
g6467 nor n6256 n6658 ; n6659
g6468 nor n6656 n6659 ; n6660
g6469 nor asqrt[57] n6641 ; n6661
g6470 and n6651_not n6661 ; n6662
g6471 nor n6660 n6662 ; n6663
g6472 nor n6653 n6663 ; n6664
g6473 and asqrt[58] n6664_not ; n6665
g6474 and n6268 n6270_not ; n6666
g6475 and n6261_not n6666 ; n6667
g6476 and asqrt[32] n6667 ; n6668
g6477 nor n6261 n6270 ; n6669
g6478 and asqrt[32] n6669 ; n6670
g6479 nor n6268 n6670 ; n6671
g6480 nor n6668 n6671 ; n6672
g6481 nor asqrt[58] n6653 ; n6673
g6482 and n6663_not n6673 ; n6674
g6483 nor n6672 n6674 ; n6675
g6484 nor n6665 n6675 ; n6676
g6485 and asqrt[59] n6676_not ; n6677
g6486 and n6273_not n6280 ; n6678
g6487 and n6282_not n6678 ; n6679
g6488 and asqrt[32] n6679 ; n6680
g6489 nor n6273 n6282 ; n6681
g6490 and asqrt[32] n6681 ; n6682
g6491 nor n6280 n6682 ; n6683
g6492 nor n6680 n6683 ; n6684
g6493 nor asqrt[59] n6665 ; n6685
g6494 and n6675_not n6685 ; n6686
g6495 nor n6684 n6686 ; n6687
g6496 nor n6677 n6687 ; n6688
g6497 and asqrt[60] n6688_not ; n6689
g6498 and n6292 n6294_not ; n6690
g6499 and n6285_not n6690 ; n6691
g6500 and asqrt[32] n6691 ; n6692
g6501 nor n6285 n6294 ; n6693
g6502 and asqrt[32] n6693 ; n6694
g6503 nor n6292 n6694 ; n6695
g6504 nor n6692 n6695 ; n6696
g6505 nor asqrt[60] n6677 ; n6697
g6506 and n6687_not n6697 ; n6698
g6507 nor n6696 n6698 ; n6699
g6508 nor n6689 n6699 ; n6700
g6509 and asqrt[61] n6700_not ; n6701
g6510 and n6297_not n6304 ; n6702
g6511 and n6306_not n6702 ; n6703
g6512 and asqrt[32] n6703 ; n6704
g6513 nor n6297 n6306 ; n6705
g6514 and asqrt[32] n6705 ; n6706
g6515 nor n6304 n6706 ; n6707
g6516 nor n6704 n6707 ; n6708
g6517 nor asqrt[61] n6689 ; n6709
g6518 and n6699_not n6709 ; n6710
g6519 nor n6708 n6710 ; n6711
g6520 nor n6701 n6711 ; n6712
g6521 and asqrt[62] n6712_not ; n6713
g6522 and n6316 n6318_not ; n6714
g6523 and n6309_not n6714 ; n6715
g6524 and asqrt[32] n6715 ; n6716
g6525 nor n6309 n6318 ; n6717
g6526 and asqrt[32] n6717 ; n6718
g6527 nor n6316 n6718 ; n6719
g6528 nor n6716 n6719 ; n6720
g6529 nor asqrt[62] n6701 ; n6721
g6530 and n6711_not n6721 ; n6722
g6531 nor n6720 n6722 ; n6723
g6532 nor n6713 n6723 ; n6724
g6533 and n6321_not n6328 ; n6725
g6534 and n6330_not n6725 ; n6726
g6535 and asqrt[32] n6726 ; n6727
g6536 nor n6321 n6330 ; n6728
g6537 and asqrt[32] n6728 ; n6729
g6538 nor n6328 n6729 ; n6730
g6539 nor n6727 n6730 ; n6731
g6540 nor n6332 n6339 ; n6732
g6541 and asqrt[32] n6732 ; n6733
g6542 nor n6347 n6733 ; n6734
g6543 and n6731_not n6734 ; n6735
g6544 and n6724_not n6735 ; n6736
g6545 nor asqrt[63] n6736 ; n6737
g6546 and n6713_not n6731 ; n6738
g6547 and n6723_not n6738 ; n6739
g6548 and n6339_not asqrt[32] ; n6740
g6549 and n6332 n6740_not ; n6741
g6550 and asqrt[63] n6732_not ; n6742
g6551 and n6741_not n6742 ; n6743
g6552 nor n6335 n6356 ; n6744
g6553 and n6338_not n6744 ; n6745
g6554 and n6351_not n6745 ; n6746
g6555 and n6347_not n6746 ; n6747
g6556 and n6345_not n6747 ; n6748
g6557 nor n6743 n6748 ; n6749
g6558 and n6739_not n6749 ; n6750
g6559 nand n6737_not n6750 ; asqrt[31]
g6560 and a[62] asqrt[31] ; n6752
g6561 nor a[60] a[61] ; n6753
g6562 and a[62]_not n6753 ; n6754
g6563 nor n6752 n6754 ; n6755
g6564 and asqrt[32] n6755_not ; n6756
g6565 nor n6356 n6754 ; n6757
g6566 and n6351_not n6757 ; n6758
g6567 and n6347_not n6758 ; n6759
g6568 and n6345_not n6759 ; n6760
g6569 and n6752_not n6760 ; n6761
g6570 and a[62]_not asqrt[31] ; n6762
g6571 and a[63] n6762_not ; n6763
g6572 and n6361 asqrt[31] ; n6764
g6573 nor n6763 n6764 ; n6765
g6574 and n6761_not n6765 ; n6766
g6575 nor n6756 n6766 ; n6767
g6576 and asqrt[33] n6767_not ; n6768
g6577 nor asqrt[33] n6756 ; n6769
g6578 and n6766_not n6769 ; n6770
g6579 and asqrt[32] n6748_not ; n6771
g6580 and n6743_not n6771 ; n6772
g6581 and n6739_not n6772 ; n6773
g6582 and n6737_not n6773 ; n6774
g6583 nor n6764 n6774 ; n6775
g6584 and a[64] n6775_not ; n6776
g6585 nor a[64] n6774 ; n6777
g6586 and n6764_not n6777 ; n6778
g6587 nor n6776 n6778 ; n6779
g6588 nor n6770 n6779 ; n6780
g6589 nor n6768 n6780 ; n6781
g6590 and asqrt[34] n6781_not ; n6782
g6591 nor asqrt[34] n6768 ; n6783
g6592 and n6780_not n6783 ; n6784
g6593 nor n6368 n6373 ; n6785
g6594 and n6364_not n6785 ; n6786
g6595 and asqrt[31] n6786 ; n6787
g6596 nor n6364 n6373 ; n6788
g6597 and asqrt[31] n6788 ; n6789
g6598 and n6368 n6789_not ; n6790
g6599 nor n6787 n6790 ; n6791
g6600 nor n6784 n6791 ; n6792
g6601 nor n6782 n6792 ; n6793
g6602 and asqrt[35] n6793_not ; n6794
g6603 and n6378_not n6387 ; n6795
g6604 and n6376_not n6795 ; n6796
g6605 and asqrt[31] n6796 ; n6797
g6606 nor n6376 n6378 ; n6798
g6607 and asqrt[31] n6798 ; n6799
g6608 nor n6387 n6799 ; n6800
g6609 nor n6797 n6800 ; n6801
g6610 nor asqrt[35] n6782 ; n6802
g6611 and n6792_not n6802 ; n6803
g6612 nor n6801 n6803 ; n6804
g6613 nor n6794 n6804 ; n6805
g6614 and asqrt[36] n6805_not ; n6806
g6615 and n6390_not n6396 ; n6807
g6616 and n6398_not n6807 ; n6808
g6617 and asqrt[31] n6808 ; n6809
g6618 nor n6390 n6398 ; n6810
g6619 and asqrt[31] n6810 ; n6811
g6620 nor n6396 n6811 ; n6812
g6621 nor n6809 n6812 ; n6813
g6622 nor asqrt[36] n6794 ; n6814
g6623 and n6804_not n6814 ; n6815
g6624 nor n6813 n6815 ; n6816
g6625 nor n6806 n6816 ; n6817
g6626 and asqrt[37] n6817_not ; n6818
g6627 and n6408 n6410_not ; n6819
g6628 and n6401_not n6819 ; n6820
g6629 and asqrt[31] n6820 ; n6821
g6630 nor n6401 n6410 ; n6822
g6631 and asqrt[31] n6822 ; n6823
g6632 nor n6408 n6823 ; n6824
g6633 nor n6821 n6824 ; n6825
g6634 nor asqrt[37] n6806 ; n6826
g6635 and n6816_not n6826 ; n6827
g6636 nor n6825 n6827 ; n6828
g6637 nor n6818 n6828 ; n6829
g6638 and asqrt[38] n6829_not ; n6830
g6639 and n6413_not n6420 ; n6831
g6640 and n6422_not n6831 ; n6832
g6641 and asqrt[31] n6832 ; n6833
g6642 nor n6413 n6422 ; n6834
g6643 and asqrt[31] n6834 ; n6835
g6644 nor n6420 n6835 ; n6836
g6645 nor n6833 n6836 ; n6837
g6646 nor asqrt[38] n6818 ; n6838
g6647 and n6828_not n6838 ; n6839
g6648 nor n6837 n6839 ; n6840
g6649 nor n6830 n6840 ; n6841
g6650 and asqrt[39] n6841_not ; n6842
g6651 and n6432 n6434_not ; n6843
g6652 and n6425_not n6843 ; n6844
g6653 and asqrt[31] n6844 ; n6845
g6654 nor n6425 n6434 ; n6846
g6655 and asqrt[31] n6846 ; n6847
g6656 nor n6432 n6847 ; n6848
g6657 nor n6845 n6848 ; n6849
g6658 nor asqrt[39] n6830 ; n6850
g6659 and n6840_not n6850 ; n6851
g6660 nor n6849 n6851 ; n6852
g6661 nor n6842 n6852 ; n6853
g6662 and asqrt[40] n6853_not ; n6854
g6663 and n6437_not n6444 ; n6855
g6664 and n6446_not n6855 ; n6856
g6665 and asqrt[31] n6856 ; n6857
g6666 nor n6437 n6446 ; n6858
g6667 and asqrt[31] n6858 ; n6859
g6668 nor n6444 n6859 ; n6860
g6669 nor n6857 n6860 ; n6861
g6670 nor asqrt[40] n6842 ; n6862
g6671 and n6852_not n6862 ; n6863
g6672 nor n6861 n6863 ; n6864
g6673 nor n6854 n6864 ; n6865
g6674 and asqrt[41] n6865_not ; n6866
g6675 and n6456 n6458_not ; n6867
g6676 and n6449_not n6867 ; n6868
g6677 and asqrt[31] n6868 ; n6869
g6678 nor n6449 n6458 ; n6870
g6679 and asqrt[31] n6870 ; n6871
g6680 nor n6456 n6871 ; n6872
g6681 nor n6869 n6872 ; n6873
g6682 nor asqrt[41] n6854 ; n6874
g6683 and n6864_not n6874 ; n6875
g6684 nor n6873 n6875 ; n6876
g6685 nor n6866 n6876 ; n6877
g6686 and asqrt[42] n6877_not ; n6878
g6687 and n6461_not n6468 ; n6879
g6688 and n6470_not n6879 ; n6880
g6689 and asqrt[31] n6880 ; n6881
g6690 nor n6461 n6470 ; n6882
g6691 and asqrt[31] n6882 ; n6883
g6692 nor n6468 n6883 ; n6884
g6693 nor n6881 n6884 ; n6885
g6694 nor asqrt[42] n6866 ; n6886
g6695 and n6876_not n6886 ; n6887
g6696 nor n6885 n6887 ; n6888
g6697 nor n6878 n6888 ; n6889
g6698 and asqrt[43] n6889_not ; n6890
g6699 and n6480 n6482_not ; n6891
g6700 and n6473_not n6891 ; n6892
g6701 and asqrt[31] n6892 ; n6893
g6702 nor n6473 n6482 ; n6894
g6703 and asqrt[31] n6894 ; n6895
g6704 nor n6480 n6895 ; n6896
g6705 nor n6893 n6896 ; n6897
g6706 nor asqrt[43] n6878 ; n6898
g6707 and n6888_not n6898 ; n6899
g6708 nor n6897 n6899 ; n6900
g6709 nor n6890 n6900 ; n6901
g6710 and asqrt[44] n6901_not ; n6902
g6711 and n6485_not n6492 ; n6903
g6712 and n6494_not n6903 ; n6904
g6713 and asqrt[31] n6904 ; n6905
g6714 nor n6485 n6494 ; n6906
g6715 and asqrt[31] n6906 ; n6907
g6716 nor n6492 n6907 ; n6908
g6717 nor n6905 n6908 ; n6909
g6718 nor asqrt[44] n6890 ; n6910
g6719 and n6900_not n6910 ; n6911
g6720 nor n6909 n6911 ; n6912
g6721 nor n6902 n6912 ; n6913
g6722 and asqrt[45] n6913_not ; n6914
g6723 and n6504 n6506_not ; n6915
g6724 and n6497_not n6915 ; n6916
g6725 and asqrt[31] n6916 ; n6917
g6726 nor n6497 n6506 ; n6918
g6727 and asqrt[31] n6918 ; n6919
g6728 nor n6504 n6919 ; n6920
g6729 nor n6917 n6920 ; n6921
g6730 nor asqrt[45] n6902 ; n6922
g6731 and n6912_not n6922 ; n6923
g6732 nor n6921 n6923 ; n6924
g6733 nor n6914 n6924 ; n6925
g6734 and asqrt[46] n6925_not ; n6926
g6735 and n6509_not n6516 ; n6927
g6736 and n6518_not n6927 ; n6928
g6737 and asqrt[31] n6928 ; n6929
g6738 nor n6509 n6518 ; n6930
g6739 and asqrt[31] n6930 ; n6931
g6740 nor n6516 n6931 ; n6932
g6741 nor n6929 n6932 ; n6933
g6742 nor asqrt[46] n6914 ; n6934
g6743 and n6924_not n6934 ; n6935
g6744 nor n6933 n6935 ; n6936
g6745 nor n6926 n6936 ; n6937
g6746 and asqrt[47] n6937_not ; n6938
g6747 and n6528 n6530_not ; n6939
g6748 and n6521_not n6939 ; n6940
g6749 and asqrt[31] n6940 ; n6941
g6750 nor n6521 n6530 ; n6942
g6751 and asqrt[31] n6942 ; n6943
g6752 nor n6528 n6943 ; n6944
g6753 nor n6941 n6944 ; n6945
g6754 nor asqrt[47] n6926 ; n6946
g6755 and n6936_not n6946 ; n6947
g6756 nor n6945 n6947 ; n6948
g6757 nor n6938 n6948 ; n6949
g6758 and asqrt[48] n6949_not ; n6950
g6759 and n6533_not n6540 ; n6951
g6760 and n6542_not n6951 ; n6952
g6761 and asqrt[31] n6952 ; n6953
g6762 nor n6533 n6542 ; n6954
g6763 and asqrt[31] n6954 ; n6955
g6764 nor n6540 n6955 ; n6956
g6765 nor n6953 n6956 ; n6957
g6766 nor asqrt[48] n6938 ; n6958
g6767 and n6948_not n6958 ; n6959
g6768 nor n6957 n6959 ; n6960
g6769 nor n6950 n6960 ; n6961
g6770 and asqrt[49] n6961_not ; n6962
g6771 and n6552 n6554_not ; n6963
g6772 and n6545_not n6963 ; n6964
g6773 and asqrt[31] n6964 ; n6965
g6774 nor n6545 n6554 ; n6966
g6775 and asqrt[31] n6966 ; n6967
g6776 nor n6552 n6967 ; n6968
g6777 nor n6965 n6968 ; n6969
g6778 nor asqrt[49] n6950 ; n6970
g6779 and n6960_not n6970 ; n6971
g6780 nor n6969 n6971 ; n6972
g6781 nor n6962 n6972 ; n6973
g6782 and asqrt[50] n6973_not ; n6974
g6783 and n6557_not n6564 ; n6975
g6784 and n6566_not n6975 ; n6976
g6785 and asqrt[31] n6976 ; n6977
g6786 nor n6557 n6566 ; n6978
g6787 and asqrt[31] n6978 ; n6979
g6788 nor n6564 n6979 ; n6980
g6789 nor n6977 n6980 ; n6981
g6790 nor asqrt[50] n6962 ; n6982
g6791 and n6972_not n6982 ; n6983
g6792 nor n6981 n6983 ; n6984
g6793 nor n6974 n6984 ; n6985
g6794 and asqrt[51] n6985_not ; n6986
g6795 and n6576 n6578_not ; n6987
g6796 and n6569_not n6987 ; n6988
g6797 and asqrt[31] n6988 ; n6989
g6798 nor n6569 n6578 ; n6990
g6799 and asqrt[31] n6990 ; n6991
g6800 nor n6576 n6991 ; n6992
g6801 nor n6989 n6992 ; n6993
g6802 nor asqrt[51] n6974 ; n6994
g6803 and n6984_not n6994 ; n6995
g6804 nor n6993 n6995 ; n6996
g6805 nor n6986 n6996 ; n6997
g6806 and asqrt[52] n6997_not ; n6998
g6807 and n6581_not n6588 ; n6999
g6808 and n6590_not n6999 ; n7000
g6809 and asqrt[31] n7000 ; n7001
g6810 nor n6581 n6590 ; n7002
g6811 and asqrt[31] n7002 ; n7003
g6812 nor n6588 n7003 ; n7004
g6813 nor n7001 n7004 ; n7005
g6814 nor asqrt[52] n6986 ; n7006
g6815 and n6996_not n7006 ; n7007
g6816 nor n7005 n7007 ; n7008
g6817 nor n6998 n7008 ; n7009
g6818 and asqrt[53] n7009_not ; n7010
g6819 and n6600 n6602_not ; n7011
g6820 and n6593_not n7011 ; n7012
g6821 and asqrt[31] n7012 ; n7013
g6822 nor n6593 n6602 ; n7014
g6823 and asqrt[31] n7014 ; n7015
g6824 nor n6600 n7015 ; n7016
g6825 nor n7013 n7016 ; n7017
g6826 nor asqrt[53] n6998 ; n7018
g6827 and n7008_not n7018 ; n7019
g6828 nor n7017 n7019 ; n7020
g6829 nor n7010 n7020 ; n7021
g6830 and asqrt[54] n7021_not ; n7022
g6831 and n6605_not n6612 ; n7023
g6832 and n6614_not n7023 ; n7024
g6833 and asqrt[31] n7024 ; n7025
g6834 nor n6605 n6614 ; n7026
g6835 and asqrt[31] n7026 ; n7027
g6836 nor n6612 n7027 ; n7028
g6837 nor n7025 n7028 ; n7029
g6838 nor asqrt[54] n7010 ; n7030
g6839 and n7020_not n7030 ; n7031
g6840 nor n7029 n7031 ; n7032
g6841 nor n7022 n7032 ; n7033
g6842 and asqrt[55] n7033_not ; n7034
g6843 and n6624 n6626_not ; n7035
g6844 and n6617_not n7035 ; n7036
g6845 and asqrt[31] n7036 ; n7037
g6846 nor n6617 n6626 ; n7038
g6847 and asqrt[31] n7038 ; n7039
g6848 nor n6624 n7039 ; n7040
g6849 nor n7037 n7040 ; n7041
g6850 nor asqrt[55] n7022 ; n7042
g6851 and n7032_not n7042 ; n7043
g6852 nor n7041 n7043 ; n7044
g6853 nor n7034 n7044 ; n7045
g6854 and asqrt[56] n7045_not ; n7046
g6855 and n6629_not n6636 ; n7047
g6856 and n6638_not n7047 ; n7048
g6857 and asqrt[31] n7048 ; n7049
g6858 nor n6629 n6638 ; n7050
g6859 and asqrt[31] n7050 ; n7051
g6860 nor n6636 n7051 ; n7052
g6861 nor n7049 n7052 ; n7053
g6862 nor asqrt[56] n7034 ; n7054
g6863 and n7044_not n7054 ; n7055
g6864 nor n7053 n7055 ; n7056
g6865 nor n7046 n7056 ; n7057
g6866 and asqrt[57] n7057_not ; n7058
g6867 and n6648 n6650_not ; n7059
g6868 and n6641_not n7059 ; n7060
g6869 and asqrt[31] n7060 ; n7061
g6870 nor n6641 n6650 ; n7062
g6871 and asqrt[31] n7062 ; n7063
g6872 nor n6648 n7063 ; n7064
g6873 nor n7061 n7064 ; n7065
g6874 nor asqrt[57] n7046 ; n7066
g6875 and n7056_not n7066 ; n7067
g6876 nor n7065 n7067 ; n7068
g6877 nor n7058 n7068 ; n7069
g6878 and asqrt[58] n7069_not ; n7070
g6879 and n6653_not n6660 ; n7071
g6880 and n6662_not n7071 ; n7072
g6881 and asqrt[31] n7072 ; n7073
g6882 nor n6653 n6662 ; n7074
g6883 and asqrt[31] n7074 ; n7075
g6884 nor n6660 n7075 ; n7076
g6885 nor n7073 n7076 ; n7077
g6886 nor asqrt[58] n7058 ; n7078
g6887 and n7068_not n7078 ; n7079
g6888 nor n7077 n7079 ; n7080
g6889 nor n7070 n7080 ; n7081
g6890 and asqrt[59] n7081_not ; n7082
g6891 and n6672 n6674_not ; n7083
g6892 and n6665_not n7083 ; n7084
g6893 and asqrt[31] n7084 ; n7085
g6894 nor n6665 n6674 ; n7086
g6895 and asqrt[31] n7086 ; n7087
g6896 nor n6672 n7087 ; n7088
g6897 nor n7085 n7088 ; n7089
g6898 nor asqrt[59] n7070 ; n7090
g6899 and n7080_not n7090 ; n7091
g6900 nor n7089 n7091 ; n7092
g6901 nor n7082 n7092 ; n7093
g6902 and asqrt[60] n7093_not ; n7094
g6903 and n6677_not n6684 ; n7095
g6904 and n6686_not n7095 ; n7096
g6905 and asqrt[31] n7096 ; n7097
g6906 nor n6677 n6686 ; n7098
g6907 and asqrt[31] n7098 ; n7099
g6908 nor n6684 n7099 ; n7100
g6909 nor n7097 n7100 ; n7101
g6910 nor asqrt[60] n7082 ; n7102
g6911 and n7092_not n7102 ; n7103
g6912 nor n7101 n7103 ; n7104
g6913 nor n7094 n7104 ; n7105
g6914 and asqrt[61] n7105_not ; n7106
g6915 and n6696 n6698_not ; n7107
g6916 and n6689_not n7107 ; n7108
g6917 and asqrt[31] n7108 ; n7109
g6918 nor n6689 n6698 ; n7110
g6919 and asqrt[31] n7110 ; n7111
g6920 nor n6696 n7111 ; n7112
g6921 nor n7109 n7112 ; n7113
g6922 nor asqrt[61] n7094 ; n7114
g6923 and n7104_not n7114 ; n7115
g6924 nor n7113 n7115 ; n7116
g6925 nor n7106 n7116 ; n7117
g6926 and asqrt[62] n7117_not ; n7118
g6927 and n6701_not n6708 ; n7119
g6928 and n6710_not n7119 ; n7120
g6929 and asqrt[31] n7120 ; n7121
g6930 nor n6701 n6710 ; n7122
g6931 and asqrt[31] n7122 ; n7123
g6932 nor n6708 n7123 ; n7124
g6933 nor n7121 n7124 ; n7125
g6934 nor asqrt[62] n7106 ; n7126
g6935 and n7116_not n7126 ; n7127
g6936 nor n7125 n7127 ; n7128
g6937 nor n7118 n7128 ; n7129
g6938 and n6720 n6722_not ; n7130
g6939 and n6713_not n7130 ; n7131
g6940 and asqrt[31] n7131 ; n7132
g6941 nor n6713 n6722 ; n7133
g6942 and asqrt[31] n7133 ; n7134
g6943 nor n6720 n7134 ; n7135
g6944 nor n7132 n7135 ; n7136
g6945 nor n6724 n6731 ; n7137
g6946 and asqrt[31] n7137 ; n7138
g6947 nor n6739 n7138 ; n7139
g6948 and n7136_not n7139 ; n7140
g6949 and n7129_not n7140 ; n7141
g6950 nor asqrt[63] n7141 ; n7142
g6951 and n7118_not n7136 ; n7143
g6952 and n7128_not n7143 ; n7144
g6953 and n6731_not asqrt[31] ; n7145
g6954 and n6724 n7145_not ; n7146
g6955 and asqrt[63] n7137_not ; n7147
g6956 and n7146_not n7147 ; n7148
g6957 nor n6727 n6748 ; n7149
g6958 and n6730_not n7149 ; n7150
g6959 and n6743_not n7150 ; n7151
g6960 and n6739_not n7151 ; n7152
g6961 and n6737_not n7152 ; n7153
g6962 nor n7148 n7153 ; n7154
g6963 and n7144_not n7154 ; n7155
g6964 nand n7142_not n7155 ; asqrt[30]
g6965 and a[60] asqrt[30] ; n7157
g6966 nor a[58] a[59] ; n7158
g6967 and a[60]_not n7158 ; n7159
g6968 nor n7157 n7159 ; n7160
g6969 and asqrt[31] n7160_not ; n7161
g6970 nor n6748 n7159 ; n7162
g6971 and n6743_not n7162 ; n7163
g6972 and n6739_not n7163 ; n7164
g6973 and n6737_not n7164 ; n7165
g6974 and n7157_not n7165 ; n7166
g6975 and a[60]_not asqrt[30] ; n7167
g6976 and a[61] n7167_not ; n7168
g6977 and n6753 asqrt[30] ; n7169
g6978 nor n7168 n7169 ; n7170
g6979 and n7166_not n7170 ; n7171
g6980 nor n7161 n7171 ; n7172
g6981 and asqrt[32] n7172_not ; n7173
g6982 nor asqrt[32] n7161 ; n7174
g6983 and n7171_not n7174 ; n7175
g6984 and asqrt[31] n7153_not ; n7176
g6985 and n7148_not n7176 ; n7177
g6986 and n7144_not n7177 ; n7178
g6987 and n7142_not n7178 ; n7179
g6988 nor n7169 n7179 ; n7180
g6989 and a[62] n7180_not ; n7181
g6990 nor a[62] n7179 ; n7182
g6991 and n7169_not n7182 ; n7183
g6992 nor n7181 n7183 ; n7184
g6993 nor n7175 n7184 ; n7185
g6994 nor n7173 n7185 ; n7186
g6995 and asqrt[33] n7186_not ; n7187
g6996 nor n6756 n6761 ; n7188
g6997 and n6765_not n7188 ; n7189
g6998 and asqrt[30] n7189 ; n7190
g6999 and asqrt[30] n7188 ; n7191
g7000 and n6765 n7191_not ; n7192
g7001 nor n7190 n7192 ; n7193
g7002 nor asqrt[33] n7173 ; n7194
g7003 and n7185_not n7194 ; n7195
g7004 nor n7193 n7195 ; n7196
g7005 nor n7187 n7196 ; n7197
g7006 and asqrt[34] n7197_not ; n7198
g7007 and n6770_not n6779 ; n7199
g7008 and n6768_not n7199 ; n7200
g7009 and asqrt[30] n7200 ; n7201
g7010 nor n6768 n6770 ; n7202
g7011 and asqrt[30] n7202 ; n7203
g7012 nor n6779 n7203 ; n7204
g7013 nor n7201 n7204 ; n7205
g7014 nor asqrt[34] n7187 ; n7206
g7015 and n7196_not n7206 ; n7207
g7016 nor n7205 n7207 ; n7208
g7017 nor n7198 n7208 ; n7209
g7018 and asqrt[35] n7209_not ; n7210
g7019 nor asqrt[35] n7198 ; n7211
g7020 and n7208_not n7211 ; n7212
g7021 and n6782_not n6791 ; n7213
g7022 and n6784_not n7213 ; n7214
g7023 and asqrt[30] n7214 ; n7215
g7024 nor n6782 n6784 ; n7216
g7025 and asqrt[30] n7216 ; n7217
g7026 nor n6791 n7217 ; n7218
g7027 nor n7215 n7218 ; n7219
g7028 nor n7212 n7219 ; n7220
g7029 nor n7210 n7220 ; n7221
g7030 and asqrt[36] n7221_not ; n7222
g7031 and n6801 n6803_not ; n7223
g7032 and n6794_not n7223 ; n7224
g7033 and asqrt[30] n7224 ; n7225
g7034 nor n6794 n6803 ; n7226
g7035 and asqrt[30] n7226 ; n7227
g7036 nor n6801 n7227 ; n7228
g7037 nor n7225 n7228 ; n7229
g7038 nor asqrt[36] n7210 ; n7230
g7039 and n7220_not n7230 ; n7231
g7040 nor n7229 n7231 ; n7232
g7041 nor n7222 n7232 ; n7233
g7042 and asqrt[37] n7233_not ; n7234
g7043 and n6806_not n6813 ; n7235
g7044 and n6815_not n7235 ; n7236
g7045 and asqrt[30] n7236 ; n7237
g7046 nor n6806 n6815 ; n7238
g7047 and asqrt[30] n7238 ; n7239
g7048 nor n6813 n7239 ; n7240
g7049 nor n7237 n7240 ; n7241
g7050 nor asqrt[37] n7222 ; n7242
g7051 and n7232_not n7242 ; n7243
g7052 nor n7241 n7243 ; n7244
g7053 nor n7234 n7244 ; n7245
g7054 and asqrt[38] n7245_not ; n7246
g7055 and n6825 n6827_not ; n7247
g7056 and n6818_not n7247 ; n7248
g7057 and asqrt[30] n7248 ; n7249
g7058 nor n6818 n6827 ; n7250
g7059 and asqrt[30] n7250 ; n7251
g7060 nor n6825 n7251 ; n7252
g7061 nor n7249 n7252 ; n7253
g7062 nor asqrt[38] n7234 ; n7254
g7063 and n7244_not n7254 ; n7255
g7064 nor n7253 n7255 ; n7256
g7065 nor n7246 n7256 ; n7257
g7066 and asqrt[39] n7257_not ; n7258
g7067 and n6830_not n6837 ; n7259
g7068 and n6839_not n7259 ; n7260
g7069 and asqrt[30] n7260 ; n7261
g7070 nor n6830 n6839 ; n7262
g7071 and asqrt[30] n7262 ; n7263
g7072 nor n6837 n7263 ; n7264
g7073 nor n7261 n7264 ; n7265
g7074 nor asqrt[39] n7246 ; n7266
g7075 and n7256_not n7266 ; n7267
g7076 nor n7265 n7267 ; n7268
g7077 nor n7258 n7268 ; n7269
g7078 and asqrt[40] n7269_not ; n7270
g7079 and n6849 n6851_not ; n7271
g7080 and n6842_not n7271 ; n7272
g7081 and asqrt[30] n7272 ; n7273
g7082 nor n6842 n6851 ; n7274
g7083 and asqrt[30] n7274 ; n7275
g7084 nor n6849 n7275 ; n7276
g7085 nor n7273 n7276 ; n7277
g7086 nor asqrt[40] n7258 ; n7278
g7087 and n7268_not n7278 ; n7279
g7088 nor n7277 n7279 ; n7280
g7089 nor n7270 n7280 ; n7281
g7090 and asqrt[41] n7281_not ; n7282
g7091 and n6854_not n6861 ; n7283
g7092 and n6863_not n7283 ; n7284
g7093 and asqrt[30] n7284 ; n7285
g7094 nor n6854 n6863 ; n7286
g7095 and asqrt[30] n7286 ; n7287
g7096 nor n6861 n7287 ; n7288
g7097 nor n7285 n7288 ; n7289
g7098 nor asqrt[41] n7270 ; n7290
g7099 and n7280_not n7290 ; n7291
g7100 nor n7289 n7291 ; n7292
g7101 nor n7282 n7292 ; n7293
g7102 and asqrt[42] n7293_not ; n7294
g7103 and n6873 n6875_not ; n7295
g7104 and n6866_not n7295 ; n7296
g7105 and asqrt[30] n7296 ; n7297
g7106 nor n6866 n6875 ; n7298
g7107 and asqrt[30] n7298 ; n7299
g7108 nor n6873 n7299 ; n7300
g7109 nor n7297 n7300 ; n7301
g7110 nor asqrt[42] n7282 ; n7302
g7111 and n7292_not n7302 ; n7303
g7112 nor n7301 n7303 ; n7304
g7113 nor n7294 n7304 ; n7305
g7114 and asqrt[43] n7305_not ; n7306
g7115 and n6878_not n6885 ; n7307
g7116 and n6887_not n7307 ; n7308
g7117 and asqrt[30] n7308 ; n7309
g7118 nor n6878 n6887 ; n7310
g7119 and asqrt[30] n7310 ; n7311
g7120 nor n6885 n7311 ; n7312
g7121 nor n7309 n7312 ; n7313
g7122 nor asqrt[43] n7294 ; n7314
g7123 and n7304_not n7314 ; n7315
g7124 nor n7313 n7315 ; n7316
g7125 nor n7306 n7316 ; n7317
g7126 and asqrt[44] n7317_not ; n7318
g7127 and n6897 n6899_not ; n7319
g7128 and n6890_not n7319 ; n7320
g7129 and asqrt[30] n7320 ; n7321
g7130 nor n6890 n6899 ; n7322
g7131 and asqrt[30] n7322 ; n7323
g7132 nor n6897 n7323 ; n7324
g7133 nor n7321 n7324 ; n7325
g7134 nor asqrt[44] n7306 ; n7326
g7135 and n7316_not n7326 ; n7327
g7136 nor n7325 n7327 ; n7328
g7137 nor n7318 n7328 ; n7329
g7138 and asqrt[45] n7329_not ; n7330
g7139 and n6902_not n6909 ; n7331
g7140 and n6911_not n7331 ; n7332
g7141 and asqrt[30] n7332 ; n7333
g7142 nor n6902 n6911 ; n7334
g7143 and asqrt[30] n7334 ; n7335
g7144 nor n6909 n7335 ; n7336
g7145 nor n7333 n7336 ; n7337
g7146 nor asqrt[45] n7318 ; n7338
g7147 and n7328_not n7338 ; n7339
g7148 nor n7337 n7339 ; n7340
g7149 nor n7330 n7340 ; n7341
g7150 and asqrt[46] n7341_not ; n7342
g7151 and n6921 n6923_not ; n7343
g7152 and n6914_not n7343 ; n7344
g7153 and asqrt[30] n7344 ; n7345
g7154 nor n6914 n6923 ; n7346
g7155 and asqrt[30] n7346 ; n7347
g7156 nor n6921 n7347 ; n7348
g7157 nor n7345 n7348 ; n7349
g7158 nor asqrt[46] n7330 ; n7350
g7159 and n7340_not n7350 ; n7351
g7160 nor n7349 n7351 ; n7352
g7161 nor n7342 n7352 ; n7353
g7162 and asqrt[47] n7353_not ; n7354
g7163 and n6926_not n6933 ; n7355
g7164 and n6935_not n7355 ; n7356
g7165 and asqrt[30] n7356 ; n7357
g7166 nor n6926 n6935 ; n7358
g7167 and asqrt[30] n7358 ; n7359
g7168 nor n6933 n7359 ; n7360
g7169 nor n7357 n7360 ; n7361
g7170 nor asqrt[47] n7342 ; n7362
g7171 and n7352_not n7362 ; n7363
g7172 nor n7361 n7363 ; n7364
g7173 nor n7354 n7364 ; n7365
g7174 and asqrt[48] n7365_not ; n7366
g7175 and n6945 n6947_not ; n7367
g7176 and n6938_not n7367 ; n7368
g7177 and asqrt[30] n7368 ; n7369
g7178 nor n6938 n6947 ; n7370
g7179 and asqrt[30] n7370 ; n7371
g7180 nor n6945 n7371 ; n7372
g7181 nor n7369 n7372 ; n7373
g7182 nor asqrt[48] n7354 ; n7374
g7183 and n7364_not n7374 ; n7375
g7184 nor n7373 n7375 ; n7376
g7185 nor n7366 n7376 ; n7377
g7186 and asqrt[49] n7377_not ; n7378
g7187 and n6950_not n6957 ; n7379
g7188 and n6959_not n7379 ; n7380
g7189 and asqrt[30] n7380 ; n7381
g7190 nor n6950 n6959 ; n7382
g7191 and asqrt[30] n7382 ; n7383
g7192 nor n6957 n7383 ; n7384
g7193 nor n7381 n7384 ; n7385
g7194 nor asqrt[49] n7366 ; n7386
g7195 and n7376_not n7386 ; n7387
g7196 nor n7385 n7387 ; n7388
g7197 nor n7378 n7388 ; n7389
g7198 and asqrt[50] n7389_not ; n7390
g7199 and n6969 n6971_not ; n7391
g7200 and n6962_not n7391 ; n7392
g7201 and asqrt[30] n7392 ; n7393
g7202 nor n6962 n6971 ; n7394
g7203 and asqrt[30] n7394 ; n7395
g7204 nor n6969 n7395 ; n7396
g7205 nor n7393 n7396 ; n7397
g7206 nor asqrt[50] n7378 ; n7398
g7207 and n7388_not n7398 ; n7399
g7208 nor n7397 n7399 ; n7400
g7209 nor n7390 n7400 ; n7401
g7210 and asqrt[51] n7401_not ; n7402
g7211 and n6974_not n6981 ; n7403
g7212 and n6983_not n7403 ; n7404
g7213 and asqrt[30] n7404 ; n7405
g7214 nor n6974 n6983 ; n7406
g7215 and asqrt[30] n7406 ; n7407
g7216 nor n6981 n7407 ; n7408
g7217 nor n7405 n7408 ; n7409
g7218 nor asqrt[51] n7390 ; n7410
g7219 and n7400_not n7410 ; n7411
g7220 nor n7409 n7411 ; n7412
g7221 nor n7402 n7412 ; n7413
g7222 and asqrt[52] n7413_not ; n7414
g7223 and n6993 n6995_not ; n7415
g7224 and n6986_not n7415 ; n7416
g7225 and asqrt[30] n7416 ; n7417
g7226 nor n6986 n6995 ; n7418
g7227 and asqrt[30] n7418 ; n7419
g7228 nor n6993 n7419 ; n7420
g7229 nor n7417 n7420 ; n7421
g7230 nor asqrt[52] n7402 ; n7422
g7231 and n7412_not n7422 ; n7423
g7232 nor n7421 n7423 ; n7424
g7233 nor n7414 n7424 ; n7425
g7234 and asqrt[53] n7425_not ; n7426
g7235 and n6998_not n7005 ; n7427
g7236 and n7007_not n7427 ; n7428
g7237 and asqrt[30] n7428 ; n7429
g7238 nor n6998 n7007 ; n7430
g7239 and asqrt[30] n7430 ; n7431
g7240 nor n7005 n7431 ; n7432
g7241 nor n7429 n7432 ; n7433
g7242 nor asqrt[53] n7414 ; n7434
g7243 and n7424_not n7434 ; n7435
g7244 nor n7433 n7435 ; n7436
g7245 nor n7426 n7436 ; n7437
g7246 and asqrt[54] n7437_not ; n7438
g7247 and n7017 n7019_not ; n7439
g7248 and n7010_not n7439 ; n7440
g7249 and asqrt[30] n7440 ; n7441
g7250 nor n7010 n7019 ; n7442
g7251 and asqrt[30] n7442 ; n7443
g7252 nor n7017 n7443 ; n7444
g7253 nor n7441 n7444 ; n7445
g7254 nor asqrt[54] n7426 ; n7446
g7255 and n7436_not n7446 ; n7447
g7256 nor n7445 n7447 ; n7448
g7257 nor n7438 n7448 ; n7449
g7258 and asqrt[55] n7449_not ; n7450
g7259 and n7022_not n7029 ; n7451
g7260 and n7031_not n7451 ; n7452
g7261 and asqrt[30] n7452 ; n7453
g7262 nor n7022 n7031 ; n7454
g7263 and asqrt[30] n7454 ; n7455
g7264 nor n7029 n7455 ; n7456
g7265 nor n7453 n7456 ; n7457
g7266 nor asqrt[55] n7438 ; n7458
g7267 and n7448_not n7458 ; n7459
g7268 nor n7457 n7459 ; n7460
g7269 nor n7450 n7460 ; n7461
g7270 and asqrt[56] n7461_not ; n7462
g7271 and n7041 n7043_not ; n7463
g7272 and n7034_not n7463 ; n7464
g7273 and asqrt[30] n7464 ; n7465
g7274 nor n7034 n7043 ; n7466
g7275 and asqrt[30] n7466 ; n7467
g7276 nor n7041 n7467 ; n7468
g7277 nor n7465 n7468 ; n7469
g7278 nor asqrt[56] n7450 ; n7470
g7279 and n7460_not n7470 ; n7471
g7280 nor n7469 n7471 ; n7472
g7281 nor n7462 n7472 ; n7473
g7282 and asqrt[57] n7473_not ; n7474
g7283 and n7046_not n7053 ; n7475
g7284 and n7055_not n7475 ; n7476
g7285 and asqrt[30] n7476 ; n7477
g7286 nor n7046 n7055 ; n7478
g7287 and asqrt[30] n7478 ; n7479
g7288 nor n7053 n7479 ; n7480
g7289 nor n7477 n7480 ; n7481
g7290 nor asqrt[57] n7462 ; n7482
g7291 and n7472_not n7482 ; n7483
g7292 nor n7481 n7483 ; n7484
g7293 nor n7474 n7484 ; n7485
g7294 and asqrt[58] n7485_not ; n7486
g7295 and n7065 n7067_not ; n7487
g7296 and n7058_not n7487 ; n7488
g7297 and asqrt[30] n7488 ; n7489
g7298 nor n7058 n7067 ; n7490
g7299 and asqrt[30] n7490 ; n7491
g7300 nor n7065 n7491 ; n7492
g7301 nor n7489 n7492 ; n7493
g7302 nor asqrt[58] n7474 ; n7494
g7303 and n7484_not n7494 ; n7495
g7304 nor n7493 n7495 ; n7496
g7305 nor n7486 n7496 ; n7497
g7306 and asqrt[59] n7497_not ; n7498
g7307 and n7070_not n7077 ; n7499
g7308 and n7079_not n7499 ; n7500
g7309 and asqrt[30] n7500 ; n7501
g7310 nor n7070 n7079 ; n7502
g7311 and asqrt[30] n7502 ; n7503
g7312 nor n7077 n7503 ; n7504
g7313 nor n7501 n7504 ; n7505
g7314 nor asqrt[59] n7486 ; n7506
g7315 and n7496_not n7506 ; n7507
g7316 nor n7505 n7507 ; n7508
g7317 nor n7498 n7508 ; n7509
g7318 and asqrt[60] n7509_not ; n7510
g7319 and n7089 n7091_not ; n7511
g7320 and n7082_not n7511 ; n7512
g7321 and asqrt[30] n7512 ; n7513
g7322 nor n7082 n7091 ; n7514
g7323 and asqrt[30] n7514 ; n7515
g7324 nor n7089 n7515 ; n7516
g7325 nor n7513 n7516 ; n7517
g7326 nor asqrt[60] n7498 ; n7518
g7327 and n7508_not n7518 ; n7519
g7328 nor n7517 n7519 ; n7520
g7329 nor n7510 n7520 ; n7521
g7330 and asqrt[61] n7521_not ; n7522
g7331 and n7094_not n7101 ; n7523
g7332 and n7103_not n7523 ; n7524
g7333 and asqrt[30] n7524 ; n7525
g7334 nor n7094 n7103 ; n7526
g7335 and asqrt[30] n7526 ; n7527
g7336 nor n7101 n7527 ; n7528
g7337 nor n7525 n7528 ; n7529
g7338 nor asqrt[61] n7510 ; n7530
g7339 and n7520_not n7530 ; n7531
g7340 nor n7529 n7531 ; n7532
g7341 nor n7522 n7532 ; n7533
g7342 and asqrt[62] n7533_not ; n7534
g7343 and n7113 n7115_not ; n7535
g7344 and n7106_not n7535 ; n7536
g7345 and asqrt[30] n7536 ; n7537
g7346 nor n7106 n7115 ; n7538
g7347 and asqrt[30] n7538 ; n7539
g7348 nor n7113 n7539 ; n7540
g7349 nor n7537 n7540 ; n7541
g7350 nor asqrt[62] n7522 ; n7542
g7351 and n7532_not n7542 ; n7543
g7352 nor n7541 n7543 ; n7544
g7353 nor n7534 n7544 ; n7545
g7354 and n7118_not n7125 ; n7546
g7355 and n7127_not n7546 ; n7547
g7356 and asqrt[30] n7547 ; n7548
g7357 nor n7118 n7127 ; n7549
g7358 and asqrt[30] n7549 ; n7550
g7359 nor n7125 n7550 ; n7551
g7360 nor n7548 n7551 ; n7552
g7361 nor n7129 n7136 ; n7553
g7362 and asqrt[30] n7553 ; n7554
g7363 nor n7144 n7554 ; n7555
g7364 and n7552_not n7555 ; n7556
g7365 and n7545_not n7556 ; n7557
g7366 nor asqrt[63] n7557 ; n7558
g7367 and n7534_not n7552 ; n7559
g7368 and n7544_not n7559 ; n7560
g7369 and n7136_not asqrt[30] ; n7561
g7370 and n7129 n7561_not ; n7562
g7371 and asqrt[63] n7553_not ; n7563
g7372 and n7562_not n7563 ; n7564
g7373 nor n7132 n7153 ; n7565
g7374 and n7135_not n7565 ; n7566
g7375 and n7148_not n7566 ; n7567
g7376 and n7144_not n7567 ; n7568
g7377 and n7142_not n7568 ; n7569
g7378 nor n7564 n7569 ; n7570
g7379 and n7560_not n7570 ; n7571
g7380 nand n7558_not n7571 ; asqrt[29]
g7381 and a[58] asqrt[29] ; n7573
g7382 nor a[56] a[57] ; n7574
g7383 and a[58]_not n7574 ; n7575
g7384 nor n7573 n7575 ; n7576
g7385 and asqrt[30] n7576_not ; n7577
g7386 nor n7153 n7575 ; n7578
g7387 and n7148_not n7578 ; n7579
g7388 and n7144_not n7579 ; n7580
g7389 and n7142_not n7580 ; n7581
g7390 and n7573_not n7581 ; n7582
g7391 and a[58]_not asqrt[29] ; n7583
g7392 and a[59] n7583_not ; n7584
g7393 and n7158 asqrt[29] ; n7585
g7394 nor n7584 n7585 ; n7586
g7395 and n7582_not n7586 ; n7587
g7396 nor n7577 n7587 ; n7588
g7397 and asqrt[31] n7588_not ; n7589
g7398 nor asqrt[31] n7577 ; n7590
g7399 and n7587_not n7590 ; n7591
g7400 and asqrt[30] n7569_not ; n7592
g7401 and n7564_not n7592 ; n7593
g7402 and n7560_not n7593 ; n7594
g7403 and n7558_not n7594 ; n7595
g7404 nor n7585 n7595 ; n7596
g7405 and a[60] n7596_not ; n7597
g7406 nor a[60] n7595 ; n7598
g7407 and n7585_not n7598 ; n7599
g7408 nor n7597 n7599 ; n7600
g7409 nor n7591 n7600 ; n7601
g7410 nor n7589 n7601 ; n7602
g7411 and asqrt[32] n7602_not ; n7603
g7412 nor n7161 n7166 ; n7604
g7413 and n7170_not n7604 ; n7605
g7414 and asqrt[29] n7605 ; n7606
g7415 and asqrt[29] n7604 ; n7607
g7416 and n7170 n7607_not ; n7608
g7417 nor n7606 n7608 ; n7609
g7418 nor asqrt[32] n7589 ; n7610
g7419 and n7601_not n7610 ; n7611
g7420 nor n7609 n7611 ; n7612
g7421 nor n7603 n7612 ; n7613
g7422 and asqrt[33] n7613_not ; n7614
g7423 and n7175_not n7184 ; n7615
g7424 and n7173_not n7615 ; n7616
g7425 and asqrt[29] n7616 ; n7617
g7426 nor n7173 n7175 ; n7618
g7427 and asqrt[29] n7618 ; n7619
g7428 nor n7184 n7619 ; n7620
g7429 nor n7617 n7620 ; n7621
g7430 nor asqrt[33] n7603 ; n7622
g7431 and n7612_not n7622 ; n7623
g7432 nor n7621 n7623 ; n7624
g7433 nor n7614 n7624 ; n7625
g7434 and asqrt[34] n7625_not ; n7626
g7435 and n7187_not n7193 ; n7627
g7436 and n7195_not n7627 ; n7628
g7437 and asqrt[29] n7628 ; n7629
g7438 nor n7187 n7195 ; n7630
g7439 and asqrt[29] n7630 ; n7631
g7440 nor n7193 n7631 ; n7632
g7441 nor n7629 n7632 ; n7633
g7442 nor asqrt[34] n7614 ; n7634
g7443 and n7624_not n7634 ; n7635
g7444 nor n7633 n7635 ; n7636
g7445 nor n7626 n7636 ; n7637
g7446 and asqrt[35] n7637_not ; n7638
g7447 and n7205 n7207_not ; n7639
g7448 and n7198_not n7639 ; n7640
g7449 and asqrt[29] n7640 ; n7641
g7450 nor n7198 n7207 ; n7642
g7451 and asqrt[29] n7642 ; n7643
g7452 nor n7205 n7643 ; n7644
g7453 nor n7641 n7644 ; n7645
g7454 nor asqrt[35] n7626 ; n7646
g7455 and n7636_not n7646 ; n7647
g7456 nor n7645 n7647 ; n7648
g7457 nor n7638 n7648 ; n7649
g7458 and asqrt[36] n7649_not ; n7650
g7459 nor asqrt[36] n7638 ; n7651
g7460 and n7648_not n7651 ; n7652
g7461 and n7210_not n7219 ; n7653
g7462 and n7212_not n7653 ; n7654
g7463 and asqrt[29] n7654 ; n7655
g7464 nor n7210 n7212 ; n7656
g7465 and asqrt[29] n7656 ; n7657
g7466 nor n7219 n7657 ; n7658
g7467 nor n7655 n7658 ; n7659
g7468 nor n7652 n7659 ; n7660
g7469 nor n7650 n7660 ; n7661
g7470 and asqrt[37] n7661_not ; n7662
g7471 and n7229 n7231_not ; n7663
g7472 and n7222_not n7663 ; n7664
g7473 and asqrt[29] n7664 ; n7665
g7474 nor n7222 n7231 ; n7666
g7475 and asqrt[29] n7666 ; n7667
g7476 nor n7229 n7667 ; n7668
g7477 nor n7665 n7668 ; n7669
g7478 nor asqrt[37] n7650 ; n7670
g7479 and n7660_not n7670 ; n7671
g7480 nor n7669 n7671 ; n7672
g7481 nor n7662 n7672 ; n7673
g7482 and asqrt[38] n7673_not ; n7674
g7483 and n7234_not n7241 ; n7675
g7484 and n7243_not n7675 ; n7676
g7485 and asqrt[29] n7676 ; n7677
g7486 nor n7234 n7243 ; n7678
g7487 and asqrt[29] n7678 ; n7679
g7488 nor n7241 n7679 ; n7680
g7489 nor n7677 n7680 ; n7681
g7490 nor asqrt[38] n7662 ; n7682
g7491 and n7672_not n7682 ; n7683
g7492 nor n7681 n7683 ; n7684
g7493 nor n7674 n7684 ; n7685
g7494 and asqrt[39] n7685_not ; n7686
g7495 and n7253 n7255_not ; n7687
g7496 and n7246_not n7687 ; n7688
g7497 and asqrt[29] n7688 ; n7689
g7498 nor n7246 n7255 ; n7690
g7499 and asqrt[29] n7690 ; n7691
g7500 nor n7253 n7691 ; n7692
g7501 nor n7689 n7692 ; n7693
g7502 nor asqrt[39] n7674 ; n7694
g7503 and n7684_not n7694 ; n7695
g7504 nor n7693 n7695 ; n7696
g7505 nor n7686 n7696 ; n7697
g7506 and asqrt[40] n7697_not ; n7698
g7507 and n7258_not n7265 ; n7699
g7508 and n7267_not n7699 ; n7700
g7509 and asqrt[29] n7700 ; n7701
g7510 nor n7258 n7267 ; n7702
g7511 and asqrt[29] n7702 ; n7703
g7512 nor n7265 n7703 ; n7704
g7513 nor n7701 n7704 ; n7705
g7514 nor asqrt[40] n7686 ; n7706
g7515 and n7696_not n7706 ; n7707
g7516 nor n7705 n7707 ; n7708
g7517 nor n7698 n7708 ; n7709
g7518 and asqrt[41] n7709_not ; n7710
g7519 and n7277 n7279_not ; n7711
g7520 and n7270_not n7711 ; n7712
g7521 and asqrt[29] n7712 ; n7713
g7522 nor n7270 n7279 ; n7714
g7523 and asqrt[29] n7714 ; n7715
g7524 nor n7277 n7715 ; n7716
g7525 nor n7713 n7716 ; n7717
g7526 nor asqrt[41] n7698 ; n7718
g7527 and n7708_not n7718 ; n7719
g7528 nor n7717 n7719 ; n7720
g7529 nor n7710 n7720 ; n7721
g7530 and asqrt[42] n7721_not ; n7722
g7531 and n7282_not n7289 ; n7723
g7532 and n7291_not n7723 ; n7724
g7533 and asqrt[29] n7724 ; n7725
g7534 nor n7282 n7291 ; n7726
g7535 and asqrt[29] n7726 ; n7727
g7536 nor n7289 n7727 ; n7728
g7537 nor n7725 n7728 ; n7729
g7538 nor asqrt[42] n7710 ; n7730
g7539 and n7720_not n7730 ; n7731
g7540 nor n7729 n7731 ; n7732
g7541 nor n7722 n7732 ; n7733
g7542 and asqrt[43] n7733_not ; n7734
g7543 and n7301 n7303_not ; n7735
g7544 and n7294_not n7735 ; n7736
g7545 and asqrt[29] n7736 ; n7737
g7546 nor n7294 n7303 ; n7738
g7547 and asqrt[29] n7738 ; n7739
g7548 nor n7301 n7739 ; n7740
g7549 nor n7737 n7740 ; n7741
g7550 nor asqrt[43] n7722 ; n7742
g7551 and n7732_not n7742 ; n7743
g7552 nor n7741 n7743 ; n7744
g7553 nor n7734 n7744 ; n7745
g7554 and asqrt[44] n7745_not ; n7746
g7555 and n7306_not n7313 ; n7747
g7556 and n7315_not n7747 ; n7748
g7557 and asqrt[29] n7748 ; n7749
g7558 nor n7306 n7315 ; n7750
g7559 and asqrt[29] n7750 ; n7751
g7560 nor n7313 n7751 ; n7752
g7561 nor n7749 n7752 ; n7753
g7562 nor asqrt[44] n7734 ; n7754
g7563 and n7744_not n7754 ; n7755
g7564 nor n7753 n7755 ; n7756
g7565 nor n7746 n7756 ; n7757
g7566 and asqrt[45] n7757_not ; n7758
g7567 and n7325 n7327_not ; n7759
g7568 and n7318_not n7759 ; n7760
g7569 and asqrt[29] n7760 ; n7761
g7570 nor n7318 n7327 ; n7762
g7571 and asqrt[29] n7762 ; n7763
g7572 nor n7325 n7763 ; n7764
g7573 nor n7761 n7764 ; n7765
g7574 nor asqrt[45] n7746 ; n7766
g7575 and n7756_not n7766 ; n7767
g7576 nor n7765 n7767 ; n7768
g7577 nor n7758 n7768 ; n7769
g7578 and asqrt[46] n7769_not ; n7770
g7579 and n7330_not n7337 ; n7771
g7580 and n7339_not n7771 ; n7772
g7581 and asqrt[29] n7772 ; n7773
g7582 nor n7330 n7339 ; n7774
g7583 and asqrt[29] n7774 ; n7775
g7584 nor n7337 n7775 ; n7776
g7585 nor n7773 n7776 ; n7777
g7586 nor asqrt[46] n7758 ; n7778
g7587 and n7768_not n7778 ; n7779
g7588 nor n7777 n7779 ; n7780
g7589 nor n7770 n7780 ; n7781
g7590 and asqrt[47] n7781_not ; n7782
g7591 and n7349 n7351_not ; n7783
g7592 and n7342_not n7783 ; n7784
g7593 and asqrt[29] n7784 ; n7785
g7594 nor n7342 n7351 ; n7786
g7595 and asqrt[29] n7786 ; n7787
g7596 nor n7349 n7787 ; n7788
g7597 nor n7785 n7788 ; n7789
g7598 nor asqrt[47] n7770 ; n7790
g7599 and n7780_not n7790 ; n7791
g7600 nor n7789 n7791 ; n7792
g7601 nor n7782 n7792 ; n7793
g7602 and asqrt[48] n7793_not ; n7794
g7603 and n7354_not n7361 ; n7795
g7604 and n7363_not n7795 ; n7796
g7605 and asqrt[29] n7796 ; n7797
g7606 nor n7354 n7363 ; n7798
g7607 and asqrt[29] n7798 ; n7799
g7608 nor n7361 n7799 ; n7800
g7609 nor n7797 n7800 ; n7801
g7610 nor asqrt[48] n7782 ; n7802
g7611 and n7792_not n7802 ; n7803
g7612 nor n7801 n7803 ; n7804
g7613 nor n7794 n7804 ; n7805
g7614 and asqrt[49] n7805_not ; n7806
g7615 and n7373 n7375_not ; n7807
g7616 and n7366_not n7807 ; n7808
g7617 and asqrt[29] n7808 ; n7809
g7618 nor n7366 n7375 ; n7810
g7619 and asqrt[29] n7810 ; n7811
g7620 nor n7373 n7811 ; n7812
g7621 nor n7809 n7812 ; n7813
g7622 nor asqrt[49] n7794 ; n7814
g7623 and n7804_not n7814 ; n7815
g7624 nor n7813 n7815 ; n7816
g7625 nor n7806 n7816 ; n7817
g7626 and asqrt[50] n7817_not ; n7818
g7627 and n7378_not n7385 ; n7819
g7628 and n7387_not n7819 ; n7820
g7629 and asqrt[29] n7820 ; n7821
g7630 nor n7378 n7387 ; n7822
g7631 and asqrt[29] n7822 ; n7823
g7632 nor n7385 n7823 ; n7824
g7633 nor n7821 n7824 ; n7825
g7634 nor asqrt[50] n7806 ; n7826
g7635 and n7816_not n7826 ; n7827
g7636 nor n7825 n7827 ; n7828
g7637 nor n7818 n7828 ; n7829
g7638 and asqrt[51] n7829_not ; n7830
g7639 and n7397 n7399_not ; n7831
g7640 and n7390_not n7831 ; n7832
g7641 and asqrt[29] n7832 ; n7833
g7642 nor n7390 n7399 ; n7834
g7643 and asqrt[29] n7834 ; n7835
g7644 nor n7397 n7835 ; n7836
g7645 nor n7833 n7836 ; n7837
g7646 nor asqrt[51] n7818 ; n7838
g7647 and n7828_not n7838 ; n7839
g7648 nor n7837 n7839 ; n7840
g7649 nor n7830 n7840 ; n7841
g7650 and asqrt[52] n7841_not ; n7842
g7651 and n7402_not n7409 ; n7843
g7652 and n7411_not n7843 ; n7844
g7653 and asqrt[29] n7844 ; n7845
g7654 nor n7402 n7411 ; n7846
g7655 and asqrt[29] n7846 ; n7847
g7656 nor n7409 n7847 ; n7848
g7657 nor n7845 n7848 ; n7849
g7658 nor asqrt[52] n7830 ; n7850
g7659 and n7840_not n7850 ; n7851
g7660 nor n7849 n7851 ; n7852
g7661 nor n7842 n7852 ; n7853
g7662 and asqrt[53] n7853_not ; n7854
g7663 and n7421 n7423_not ; n7855
g7664 and n7414_not n7855 ; n7856
g7665 and asqrt[29] n7856 ; n7857
g7666 nor n7414 n7423 ; n7858
g7667 and asqrt[29] n7858 ; n7859
g7668 nor n7421 n7859 ; n7860
g7669 nor n7857 n7860 ; n7861
g7670 nor asqrt[53] n7842 ; n7862
g7671 and n7852_not n7862 ; n7863
g7672 nor n7861 n7863 ; n7864
g7673 nor n7854 n7864 ; n7865
g7674 and asqrt[54] n7865_not ; n7866
g7675 and n7426_not n7433 ; n7867
g7676 and n7435_not n7867 ; n7868
g7677 and asqrt[29] n7868 ; n7869
g7678 nor n7426 n7435 ; n7870
g7679 and asqrt[29] n7870 ; n7871
g7680 nor n7433 n7871 ; n7872
g7681 nor n7869 n7872 ; n7873
g7682 nor asqrt[54] n7854 ; n7874
g7683 and n7864_not n7874 ; n7875
g7684 nor n7873 n7875 ; n7876
g7685 nor n7866 n7876 ; n7877
g7686 and asqrt[55] n7877_not ; n7878
g7687 and n7445 n7447_not ; n7879
g7688 and n7438_not n7879 ; n7880
g7689 and asqrt[29] n7880 ; n7881
g7690 nor n7438 n7447 ; n7882
g7691 and asqrt[29] n7882 ; n7883
g7692 nor n7445 n7883 ; n7884
g7693 nor n7881 n7884 ; n7885
g7694 nor asqrt[55] n7866 ; n7886
g7695 and n7876_not n7886 ; n7887
g7696 nor n7885 n7887 ; n7888
g7697 nor n7878 n7888 ; n7889
g7698 and asqrt[56] n7889_not ; n7890
g7699 and n7450_not n7457 ; n7891
g7700 and n7459_not n7891 ; n7892
g7701 and asqrt[29] n7892 ; n7893
g7702 nor n7450 n7459 ; n7894
g7703 and asqrt[29] n7894 ; n7895
g7704 nor n7457 n7895 ; n7896
g7705 nor n7893 n7896 ; n7897
g7706 nor asqrt[56] n7878 ; n7898
g7707 and n7888_not n7898 ; n7899
g7708 nor n7897 n7899 ; n7900
g7709 nor n7890 n7900 ; n7901
g7710 and asqrt[57] n7901_not ; n7902
g7711 and n7469 n7471_not ; n7903
g7712 and n7462_not n7903 ; n7904
g7713 and asqrt[29] n7904 ; n7905
g7714 nor n7462 n7471 ; n7906
g7715 and asqrt[29] n7906 ; n7907
g7716 nor n7469 n7907 ; n7908
g7717 nor n7905 n7908 ; n7909
g7718 nor asqrt[57] n7890 ; n7910
g7719 and n7900_not n7910 ; n7911
g7720 nor n7909 n7911 ; n7912
g7721 nor n7902 n7912 ; n7913
g7722 and asqrt[58] n7913_not ; n7914
g7723 and n7474_not n7481 ; n7915
g7724 and n7483_not n7915 ; n7916
g7725 and asqrt[29] n7916 ; n7917
g7726 nor n7474 n7483 ; n7918
g7727 and asqrt[29] n7918 ; n7919
g7728 nor n7481 n7919 ; n7920
g7729 nor n7917 n7920 ; n7921
g7730 nor asqrt[58] n7902 ; n7922
g7731 and n7912_not n7922 ; n7923
g7732 nor n7921 n7923 ; n7924
g7733 nor n7914 n7924 ; n7925
g7734 and asqrt[59] n7925_not ; n7926
g7735 and n7493 n7495_not ; n7927
g7736 and n7486_not n7927 ; n7928
g7737 and asqrt[29] n7928 ; n7929
g7738 nor n7486 n7495 ; n7930
g7739 and asqrt[29] n7930 ; n7931
g7740 nor n7493 n7931 ; n7932
g7741 nor n7929 n7932 ; n7933
g7742 nor asqrt[59] n7914 ; n7934
g7743 and n7924_not n7934 ; n7935
g7744 nor n7933 n7935 ; n7936
g7745 nor n7926 n7936 ; n7937
g7746 and asqrt[60] n7937_not ; n7938
g7747 and n7498_not n7505 ; n7939
g7748 and n7507_not n7939 ; n7940
g7749 and asqrt[29] n7940 ; n7941
g7750 nor n7498 n7507 ; n7942
g7751 and asqrt[29] n7942 ; n7943
g7752 nor n7505 n7943 ; n7944
g7753 nor n7941 n7944 ; n7945
g7754 nor asqrt[60] n7926 ; n7946
g7755 and n7936_not n7946 ; n7947
g7756 nor n7945 n7947 ; n7948
g7757 nor n7938 n7948 ; n7949
g7758 and asqrt[61] n7949_not ; n7950
g7759 and n7517 n7519_not ; n7951
g7760 and n7510_not n7951 ; n7952
g7761 and asqrt[29] n7952 ; n7953
g7762 nor n7510 n7519 ; n7954
g7763 and asqrt[29] n7954 ; n7955
g7764 nor n7517 n7955 ; n7956
g7765 nor n7953 n7956 ; n7957
g7766 nor asqrt[61] n7938 ; n7958
g7767 and n7948_not n7958 ; n7959
g7768 nor n7957 n7959 ; n7960
g7769 nor n7950 n7960 ; n7961
g7770 and asqrt[62] n7961_not ; n7962
g7771 and n7522_not n7529 ; n7963
g7772 and n7531_not n7963 ; n7964
g7773 and asqrt[29] n7964 ; n7965
g7774 nor n7522 n7531 ; n7966
g7775 and asqrt[29] n7966 ; n7967
g7776 nor n7529 n7967 ; n7968
g7777 nor n7965 n7968 ; n7969
g7778 nor asqrt[62] n7950 ; n7970
g7779 and n7960_not n7970 ; n7971
g7780 nor n7969 n7971 ; n7972
g7781 nor n7962 n7972 ; n7973
g7782 and n7541 n7543_not ; n7974
g7783 and n7534_not n7974 ; n7975
g7784 and asqrt[29] n7975 ; n7976
g7785 nor n7534 n7543 ; n7977
g7786 and asqrt[29] n7977 ; n7978
g7787 nor n7541 n7978 ; n7979
g7788 nor n7976 n7979 ; n7980
g7789 nor n7545 n7552 ; n7981
g7790 and asqrt[29] n7981 ; n7982
g7791 nor n7560 n7982 ; n7983
g7792 and n7980_not n7983 ; n7984
g7793 and n7973_not n7984 ; n7985
g7794 nor asqrt[63] n7985 ; n7986
g7795 and n7962_not n7980 ; n7987
g7796 and n7972_not n7987 ; n7988
g7797 and n7552_not asqrt[29] ; n7989
g7798 and n7545 n7989_not ; n7990
g7799 and asqrt[63] n7981_not ; n7991
g7800 and n7990_not n7991 ; n7992
g7801 nor n7548 n7569 ; n7993
g7802 and n7551_not n7993 ; n7994
g7803 and n7564_not n7994 ; n7995
g7804 and n7560_not n7995 ; n7996
g7805 and n7558_not n7996 ; n7997
g7806 nor n7992 n7997 ; n7998
g7807 and n7988_not n7998 ; n7999
g7808 nand n7986_not n7999 ; asqrt[28]
g7809 and a[56] asqrt[28] ; n8001
g7810 nor a[54] a[55] ; n8002
g7811 and a[56]_not n8002 ; n8003
g7812 nor n8001 n8003 ; n8004
g7813 and asqrt[29] n8004_not ; n8005
g7814 nor n7569 n8003 ; n8006
g7815 and n7564_not n8006 ; n8007
g7816 and n7560_not n8007 ; n8008
g7817 and n7558_not n8008 ; n8009
g7818 and n8001_not n8009 ; n8010
g7819 and a[56]_not asqrt[28] ; n8011
g7820 and a[57] n8011_not ; n8012
g7821 and n7574 asqrt[28] ; n8013
g7822 nor n8012 n8013 ; n8014
g7823 and n8010_not n8014 ; n8015
g7824 nor n8005 n8015 ; n8016
g7825 and asqrt[30] n8016_not ; n8017
g7826 nor asqrt[30] n8005 ; n8018
g7827 and n8015_not n8018 ; n8019
g7828 and asqrt[29] n7997_not ; n8020
g7829 and n7992_not n8020 ; n8021
g7830 and n7988_not n8021 ; n8022
g7831 and n7986_not n8022 ; n8023
g7832 nor n8013 n8023 ; n8024
g7833 and a[58] n8024_not ; n8025
g7834 nor a[58] n8023 ; n8026
g7835 and n8013_not n8026 ; n8027
g7836 nor n8025 n8027 ; n8028
g7837 nor n8019 n8028 ; n8029
g7838 nor n8017 n8029 ; n8030
g7839 and asqrt[31] n8030_not ; n8031
g7840 nor n7577 n7582 ; n8032
g7841 and n7586_not n8032 ; n8033
g7842 and asqrt[28] n8033 ; n8034
g7843 and asqrt[28] n8032 ; n8035
g7844 and n7586 n8035_not ; n8036
g7845 nor n8034 n8036 ; n8037
g7846 nor asqrt[31] n8017 ; n8038
g7847 and n8029_not n8038 ; n8039
g7848 nor n8037 n8039 ; n8040
g7849 nor n8031 n8040 ; n8041
g7850 and asqrt[32] n8041_not ; n8042
g7851 and n7591_not n7600 ; n8043
g7852 and n7589_not n8043 ; n8044
g7853 and asqrt[28] n8044 ; n8045
g7854 nor n7589 n7591 ; n8046
g7855 and asqrt[28] n8046 ; n8047
g7856 nor n7600 n8047 ; n8048
g7857 nor n8045 n8048 ; n8049
g7858 nor asqrt[32] n8031 ; n8050
g7859 and n8040_not n8050 ; n8051
g7860 nor n8049 n8051 ; n8052
g7861 nor n8042 n8052 ; n8053
g7862 and asqrt[33] n8053_not ; n8054
g7863 and n7603_not n7609 ; n8055
g7864 and n7611_not n8055 ; n8056
g7865 and asqrt[28] n8056 ; n8057
g7866 nor n7603 n7611 ; n8058
g7867 and asqrt[28] n8058 ; n8059
g7868 nor n7609 n8059 ; n8060
g7869 nor n8057 n8060 ; n8061
g7870 nor asqrt[33] n8042 ; n8062
g7871 and n8052_not n8062 ; n8063
g7872 nor n8061 n8063 ; n8064
g7873 nor n8054 n8064 ; n8065
g7874 and asqrt[34] n8065_not ; n8066
g7875 and n7621 n7623_not ; n8067
g7876 and n7614_not n8067 ; n8068
g7877 and asqrt[28] n8068 ; n8069
g7878 nor n7614 n7623 ; n8070
g7879 and asqrt[28] n8070 ; n8071
g7880 nor n7621 n8071 ; n8072
g7881 nor n8069 n8072 ; n8073
g7882 nor asqrt[34] n8054 ; n8074
g7883 and n8064_not n8074 ; n8075
g7884 nor n8073 n8075 ; n8076
g7885 nor n8066 n8076 ; n8077
g7886 and asqrt[35] n8077_not ; n8078
g7887 and n7626_not n7633 ; n8079
g7888 and n7635_not n8079 ; n8080
g7889 and asqrt[28] n8080 ; n8081
g7890 nor n7626 n7635 ; n8082
g7891 and asqrt[28] n8082 ; n8083
g7892 nor n7633 n8083 ; n8084
g7893 nor n8081 n8084 ; n8085
g7894 nor asqrt[35] n8066 ; n8086
g7895 and n8076_not n8086 ; n8087
g7896 nor n8085 n8087 ; n8088
g7897 nor n8078 n8088 ; n8089
g7898 and asqrt[36] n8089_not ; n8090
g7899 and n7645 n7647_not ; n8091
g7900 and n7638_not n8091 ; n8092
g7901 and asqrt[28] n8092 ; n8093
g7902 nor n7638 n7647 ; n8094
g7903 and asqrt[28] n8094 ; n8095
g7904 nor n7645 n8095 ; n8096
g7905 nor n8093 n8096 ; n8097
g7906 nor asqrt[36] n8078 ; n8098
g7907 and n8088_not n8098 ; n8099
g7908 nor n8097 n8099 ; n8100
g7909 nor n8090 n8100 ; n8101
g7910 and asqrt[37] n8101_not ; n8102
g7911 nor asqrt[37] n8090 ; n8103
g7912 and n8100_not n8103 ; n8104
g7913 and n7650_not n7659 ; n8105
g7914 and n7652_not n8105 ; n8106
g7915 and asqrt[28] n8106 ; n8107
g7916 nor n7650 n7652 ; n8108
g7917 and asqrt[28] n8108 ; n8109
g7918 nor n7659 n8109 ; n8110
g7919 nor n8107 n8110 ; n8111
g7920 nor n8104 n8111 ; n8112
g7921 nor n8102 n8112 ; n8113
g7922 and asqrt[38] n8113_not ; n8114
g7923 and n7669 n7671_not ; n8115
g7924 and n7662_not n8115 ; n8116
g7925 and asqrt[28] n8116 ; n8117
g7926 nor n7662 n7671 ; n8118
g7927 and asqrt[28] n8118 ; n8119
g7928 nor n7669 n8119 ; n8120
g7929 nor n8117 n8120 ; n8121
g7930 nor asqrt[38] n8102 ; n8122
g7931 and n8112_not n8122 ; n8123
g7932 nor n8121 n8123 ; n8124
g7933 nor n8114 n8124 ; n8125
g7934 and asqrt[39] n8125_not ; n8126
g7935 and n7674_not n7681 ; n8127
g7936 and n7683_not n8127 ; n8128
g7937 and asqrt[28] n8128 ; n8129
g7938 nor n7674 n7683 ; n8130
g7939 and asqrt[28] n8130 ; n8131
g7940 nor n7681 n8131 ; n8132
g7941 nor n8129 n8132 ; n8133
g7942 nor asqrt[39] n8114 ; n8134
g7943 and n8124_not n8134 ; n8135
g7944 nor n8133 n8135 ; n8136
g7945 nor n8126 n8136 ; n8137
g7946 and asqrt[40] n8137_not ; n8138
g7947 and n7693 n7695_not ; n8139
g7948 and n7686_not n8139 ; n8140
g7949 and asqrt[28] n8140 ; n8141
g7950 nor n7686 n7695 ; n8142
g7951 and asqrt[28] n8142 ; n8143
g7952 nor n7693 n8143 ; n8144
g7953 nor n8141 n8144 ; n8145
g7954 nor asqrt[40] n8126 ; n8146
g7955 and n8136_not n8146 ; n8147
g7956 nor n8145 n8147 ; n8148
g7957 nor n8138 n8148 ; n8149
g7958 and asqrt[41] n8149_not ; n8150
g7959 and n7698_not n7705 ; n8151
g7960 and n7707_not n8151 ; n8152
g7961 and asqrt[28] n8152 ; n8153
g7962 nor n7698 n7707 ; n8154
g7963 and asqrt[28] n8154 ; n8155
g7964 nor n7705 n8155 ; n8156
g7965 nor n8153 n8156 ; n8157
g7966 nor asqrt[41] n8138 ; n8158
g7967 and n8148_not n8158 ; n8159
g7968 nor n8157 n8159 ; n8160
g7969 nor n8150 n8160 ; n8161
g7970 and asqrt[42] n8161_not ; n8162
g7971 and n7717 n7719_not ; n8163
g7972 and n7710_not n8163 ; n8164
g7973 and asqrt[28] n8164 ; n8165
g7974 nor n7710 n7719 ; n8166
g7975 and asqrt[28] n8166 ; n8167
g7976 nor n7717 n8167 ; n8168
g7977 nor n8165 n8168 ; n8169
g7978 nor asqrt[42] n8150 ; n8170
g7979 and n8160_not n8170 ; n8171
g7980 nor n8169 n8171 ; n8172
g7981 nor n8162 n8172 ; n8173
g7982 and asqrt[43] n8173_not ; n8174
g7983 and n7722_not n7729 ; n8175
g7984 and n7731_not n8175 ; n8176
g7985 and asqrt[28] n8176 ; n8177
g7986 nor n7722 n7731 ; n8178
g7987 and asqrt[28] n8178 ; n8179
g7988 nor n7729 n8179 ; n8180
g7989 nor n8177 n8180 ; n8181
g7990 nor asqrt[43] n8162 ; n8182
g7991 and n8172_not n8182 ; n8183
g7992 nor n8181 n8183 ; n8184
g7993 nor n8174 n8184 ; n8185
g7994 and asqrt[44] n8185_not ; n8186
g7995 and n7741 n7743_not ; n8187
g7996 and n7734_not n8187 ; n8188
g7997 and asqrt[28] n8188 ; n8189
g7998 nor n7734 n7743 ; n8190
g7999 and asqrt[28] n8190 ; n8191
g8000 nor n7741 n8191 ; n8192
g8001 nor n8189 n8192 ; n8193
g8002 nor asqrt[44] n8174 ; n8194
g8003 and n8184_not n8194 ; n8195
g8004 nor n8193 n8195 ; n8196
g8005 nor n8186 n8196 ; n8197
g8006 and asqrt[45] n8197_not ; n8198
g8007 and n7746_not n7753 ; n8199
g8008 and n7755_not n8199 ; n8200
g8009 and asqrt[28] n8200 ; n8201
g8010 nor n7746 n7755 ; n8202
g8011 and asqrt[28] n8202 ; n8203
g8012 nor n7753 n8203 ; n8204
g8013 nor n8201 n8204 ; n8205
g8014 nor asqrt[45] n8186 ; n8206
g8015 and n8196_not n8206 ; n8207
g8016 nor n8205 n8207 ; n8208
g8017 nor n8198 n8208 ; n8209
g8018 and asqrt[46] n8209_not ; n8210
g8019 and n7765 n7767_not ; n8211
g8020 and n7758_not n8211 ; n8212
g8021 and asqrt[28] n8212 ; n8213
g8022 nor n7758 n7767 ; n8214
g8023 and asqrt[28] n8214 ; n8215
g8024 nor n7765 n8215 ; n8216
g8025 nor n8213 n8216 ; n8217
g8026 nor asqrt[46] n8198 ; n8218
g8027 and n8208_not n8218 ; n8219
g8028 nor n8217 n8219 ; n8220
g8029 nor n8210 n8220 ; n8221
g8030 and asqrt[47] n8221_not ; n8222
g8031 and n7770_not n7777 ; n8223
g8032 and n7779_not n8223 ; n8224
g8033 and asqrt[28] n8224 ; n8225
g8034 nor n7770 n7779 ; n8226
g8035 and asqrt[28] n8226 ; n8227
g8036 nor n7777 n8227 ; n8228
g8037 nor n8225 n8228 ; n8229
g8038 nor asqrt[47] n8210 ; n8230
g8039 and n8220_not n8230 ; n8231
g8040 nor n8229 n8231 ; n8232
g8041 nor n8222 n8232 ; n8233
g8042 and asqrt[48] n8233_not ; n8234
g8043 and n7789 n7791_not ; n8235
g8044 and n7782_not n8235 ; n8236
g8045 and asqrt[28] n8236 ; n8237
g8046 nor n7782 n7791 ; n8238
g8047 and asqrt[28] n8238 ; n8239
g8048 nor n7789 n8239 ; n8240
g8049 nor n8237 n8240 ; n8241
g8050 nor asqrt[48] n8222 ; n8242
g8051 and n8232_not n8242 ; n8243
g8052 nor n8241 n8243 ; n8244
g8053 nor n8234 n8244 ; n8245
g8054 and asqrt[49] n8245_not ; n8246
g8055 and n7794_not n7801 ; n8247
g8056 and n7803_not n8247 ; n8248
g8057 and asqrt[28] n8248 ; n8249
g8058 nor n7794 n7803 ; n8250
g8059 and asqrt[28] n8250 ; n8251
g8060 nor n7801 n8251 ; n8252
g8061 nor n8249 n8252 ; n8253
g8062 nor asqrt[49] n8234 ; n8254
g8063 and n8244_not n8254 ; n8255
g8064 nor n8253 n8255 ; n8256
g8065 nor n8246 n8256 ; n8257
g8066 and asqrt[50] n8257_not ; n8258
g8067 and n7813 n7815_not ; n8259
g8068 and n7806_not n8259 ; n8260
g8069 and asqrt[28] n8260 ; n8261
g8070 nor n7806 n7815 ; n8262
g8071 and asqrt[28] n8262 ; n8263
g8072 nor n7813 n8263 ; n8264
g8073 nor n8261 n8264 ; n8265
g8074 nor asqrt[50] n8246 ; n8266
g8075 and n8256_not n8266 ; n8267
g8076 nor n8265 n8267 ; n8268
g8077 nor n8258 n8268 ; n8269
g8078 and asqrt[51] n8269_not ; n8270
g8079 and n7818_not n7825 ; n8271
g8080 and n7827_not n8271 ; n8272
g8081 and asqrt[28] n8272 ; n8273
g8082 nor n7818 n7827 ; n8274
g8083 and asqrt[28] n8274 ; n8275
g8084 nor n7825 n8275 ; n8276
g8085 nor n8273 n8276 ; n8277
g8086 nor asqrt[51] n8258 ; n8278
g8087 and n8268_not n8278 ; n8279
g8088 nor n8277 n8279 ; n8280
g8089 nor n8270 n8280 ; n8281
g8090 and asqrt[52] n8281_not ; n8282
g8091 and n7837 n7839_not ; n8283
g8092 and n7830_not n8283 ; n8284
g8093 and asqrt[28] n8284 ; n8285
g8094 nor n7830 n7839 ; n8286
g8095 and asqrt[28] n8286 ; n8287
g8096 nor n7837 n8287 ; n8288
g8097 nor n8285 n8288 ; n8289
g8098 nor asqrt[52] n8270 ; n8290
g8099 and n8280_not n8290 ; n8291
g8100 nor n8289 n8291 ; n8292
g8101 nor n8282 n8292 ; n8293
g8102 and asqrt[53] n8293_not ; n8294
g8103 and n7842_not n7849 ; n8295
g8104 and n7851_not n8295 ; n8296
g8105 and asqrt[28] n8296 ; n8297
g8106 nor n7842 n7851 ; n8298
g8107 and asqrt[28] n8298 ; n8299
g8108 nor n7849 n8299 ; n8300
g8109 nor n8297 n8300 ; n8301
g8110 nor asqrt[53] n8282 ; n8302
g8111 and n8292_not n8302 ; n8303
g8112 nor n8301 n8303 ; n8304
g8113 nor n8294 n8304 ; n8305
g8114 and asqrt[54] n8305_not ; n8306
g8115 and n7861 n7863_not ; n8307
g8116 and n7854_not n8307 ; n8308
g8117 and asqrt[28] n8308 ; n8309
g8118 nor n7854 n7863 ; n8310
g8119 and asqrt[28] n8310 ; n8311
g8120 nor n7861 n8311 ; n8312
g8121 nor n8309 n8312 ; n8313
g8122 nor asqrt[54] n8294 ; n8314
g8123 and n8304_not n8314 ; n8315
g8124 nor n8313 n8315 ; n8316
g8125 nor n8306 n8316 ; n8317
g8126 and asqrt[55] n8317_not ; n8318
g8127 and n7866_not n7873 ; n8319
g8128 and n7875_not n8319 ; n8320
g8129 and asqrt[28] n8320 ; n8321
g8130 nor n7866 n7875 ; n8322
g8131 and asqrt[28] n8322 ; n8323
g8132 nor n7873 n8323 ; n8324
g8133 nor n8321 n8324 ; n8325
g8134 nor asqrt[55] n8306 ; n8326
g8135 and n8316_not n8326 ; n8327
g8136 nor n8325 n8327 ; n8328
g8137 nor n8318 n8328 ; n8329
g8138 and asqrt[56] n8329_not ; n8330
g8139 and n7885 n7887_not ; n8331
g8140 and n7878_not n8331 ; n8332
g8141 and asqrt[28] n8332 ; n8333
g8142 nor n7878 n7887 ; n8334
g8143 and asqrt[28] n8334 ; n8335
g8144 nor n7885 n8335 ; n8336
g8145 nor n8333 n8336 ; n8337
g8146 nor asqrt[56] n8318 ; n8338
g8147 and n8328_not n8338 ; n8339
g8148 nor n8337 n8339 ; n8340
g8149 nor n8330 n8340 ; n8341
g8150 and asqrt[57] n8341_not ; n8342
g8151 and n7890_not n7897 ; n8343
g8152 and n7899_not n8343 ; n8344
g8153 and asqrt[28] n8344 ; n8345
g8154 nor n7890 n7899 ; n8346
g8155 and asqrt[28] n8346 ; n8347
g8156 nor n7897 n8347 ; n8348
g8157 nor n8345 n8348 ; n8349
g8158 nor asqrt[57] n8330 ; n8350
g8159 and n8340_not n8350 ; n8351
g8160 nor n8349 n8351 ; n8352
g8161 nor n8342 n8352 ; n8353
g8162 and asqrt[58] n8353_not ; n8354
g8163 and n7909 n7911_not ; n8355
g8164 and n7902_not n8355 ; n8356
g8165 and asqrt[28] n8356 ; n8357
g8166 nor n7902 n7911 ; n8358
g8167 and asqrt[28] n8358 ; n8359
g8168 nor n7909 n8359 ; n8360
g8169 nor n8357 n8360 ; n8361
g8170 nor asqrt[58] n8342 ; n8362
g8171 and n8352_not n8362 ; n8363
g8172 nor n8361 n8363 ; n8364
g8173 nor n8354 n8364 ; n8365
g8174 and asqrt[59] n8365_not ; n8366
g8175 and n7914_not n7921 ; n8367
g8176 and n7923_not n8367 ; n8368
g8177 and asqrt[28] n8368 ; n8369
g8178 nor n7914 n7923 ; n8370
g8179 and asqrt[28] n8370 ; n8371
g8180 nor n7921 n8371 ; n8372
g8181 nor n8369 n8372 ; n8373
g8182 nor asqrt[59] n8354 ; n8374
g8183 and n8364_not n8374 ; n8375
g8184 nor n8373 n8375 ; n8376
g8185 nor n8366 n8376 ; n8377
g8186 and asqrt[60] n8377_not ; n8378
g8187 and n7933 n7935_not ; n8379
g8188 and n7926_not n8379 ; n8380
g8189 and asqrt[28] n8380 ; n8381
g8190 nor n7926 n7935 ; n8382
g8191 and asqrt[28] n8382 ; n8383
g8192 nor n7933 n8383 ; n8384
g8193 nor n8381 n8384 ; n8385
g8194 nor asqrt[60] n8366 ; n8386
g8195 and n8376_not n8386 ; n8387
g8196 nor n8385 n8387 ; n8388
g8197 nor n8378 n8388 ; n8389
g8198 and asqrt[61] n8389_not ; n8390
g8199 and n7938_not n7945 ; n8391
g8200 and n7947_not n8391 ; n8392
g8201 and asqrt[28] n8392 ; n8393
g8202 nor n7938 n7947 ; n8394
g8203 and asqrt[28] n8394 ; n8395
g8204 nor n7945 n8395 ; n8396
g8205 nor n8393 n8396 ; n8397
g8206 nor asqrt[61] n8378 ; n8398
g8207 and n8388_not n8398 ; n8399
g8208 nor n8397 n8399 ; n8400
g8209 nor n8390 n8400 ; n8401
g8210 and asqrt[62] n8401_not ; n8402
g8211 and n7957 n7959_not ; n8403
g8212 and n7950_not n8403 ; n8404
g8213 and asqrt[28] n8404 ; n8405
g8214 nor n7950 n7959 ; n8406
g8215 and asqrt[28] n8406 ; n8407
g8216 nor n7957 n8407 ; n8408
g8217 nor n8405 n8408 ; n8409
g8218 nor asqrt[62] n8390 ; n8410
g8219 and n8400_not n8410 ; n8411
g8220 nor n8409 n8411 ; n8412
g8221 nor n8402 n8412 ; n8413
g8222 and n7962_not n7969 ; n8414
g8223 and n7971_not n8414 ; n8415
g8224 and asqrt[28] n8415 ; n8416
g8225 nor n7962 n7971 ; n8417
g8226 and asqrt[28] n8417 ; n8418
g8227 nor n7969 n8418 ; n8419
g8228 nor n8416 n8419 ; n8420
g8229 nor n7973 n7980 ; n8421
g8230 and asqrt[28] n8421 ; n8422
g8231 nor n7988 n8422 ; n8423
g8232 and n8420_not n8423 ; n8424
g8233 and n8413_not n8424 ; n8425
g8234 nor asqrt[63] n8425 ; n8426
g8235 and n8402_not n8420 ; n8427
g8236 and n8412_not n8427 ; n8428
g8237 and n7980_not asqrt[28] ; n8429
g8238 and n7973 n8429_not ; n8430
g8239 and asqrt[63] n8421_not ; n8431
g8240 and n8430_not n8431 ; n8432
g8241 nor n7976 n7997 ; n8433
g8242 and n7979_not n8433 ; n8434
g8243 and n7992_not n8434 ; n8435
g8244 and n7988_not n8435 ; n8436
g8245 and n7986_not n8436 ; n8437
g8246 nor n8432 n8437 ; n8438
g8247 and n8428_not n8438 ; n8439
g8248 nand n8426_not n8439 ; asqrt[27]
g8249 and a[54] asqrt[27] ; n8441
g8250 nor a[52] a[53] ; n8442
g8251 and a[54]_not n8442 ; n8443
g8252 nor n8441 n8443 ; n8444
g8253 and asqrt[28] n8444_not ; n8445
g8254 nor n7997 n8443 ; n8446
g8255 and n7992_not n8446 ; n8447
g8256 and n7988_not n8447 ; n8448
g8257 and n7986_not n8448 ; n8449
g8258 and n8441_not n8449 ; n8450
g8259 and a[54]_not asqrt[27] ; n8451
g8260 and a[55] n8451_not ; n8452
g8261 and n8002 asqrt[27] ; n8453
g8262 nor n8452 n8453 ; n8454
g8263 and n8450_not n8454 ; n8455
g8264 nor n8445 n8455 ; n8456
g8265 and asqrt[29] n8456_not ; n8457
g8266 nor asqrt[29] n8445 ; n8458
g8267 and n8455_not n8458 ; n8459
g8268 and asqrt[28] n8437_not ; n8460
g8269 and n8432_not n8460 ; n8461
g8270 and n8428_not n8461 ; n8462
g8271 and n8426_not n8462 ; n8463
g8272 nor n8453 n8463 ; n8464
g8273 and a[56] n8464_not ; n8465
g8274 nor a[56] n8463 ; n8466
g8275 and n8453_not n8466 ; n8467
g8276 nor n8465 n8467 ; n8468
g8277 nor n8459 n8468 ; n8469
g8278 nor n8457 n8469 ; n8470
g8279 and asqrt[30] n8470_not ; n8471
g8280 nor n8005 n8010 ; n8472
g8281 and n8014_not n8472 ; n8473
g8282 and asqrt[27] n8473 ; n8474
g8283 and asqrt[27] n8472 ; n8475
g8284 and n8014 n8475_not ; n8476
g8285 nor n8474 n8476 ; n8477
g8286 nor asqrt[30] n8457 ; n8478
g8287 and n8469_not n8478 ; n8479
g8288 nor n8477 n8479 ; n8480
g8289 nor n8471 n8480 ; n8481
g8290 and asqrt[31] n8481_not ; n8482
g8291 and n8019_not n8028 ; n8483
g8292 and n8017_not n8483 ; n8484
g8293 and asqrt[27] n8484 ; n8485
g8294 nor n8017 n8019 ; n8486
g8295 and asqrt[27] n8486 ; n8487
g8296 nor n8028 n8487 ; n8488
g8297 nor n8485 n8488 ; n8489
g8298 nor asqrt[31] n8471 ; n8490
g8299 and n8480_not n8490 ; n8491
g8300 nor n8489 n8491 ; n8492
g8301 nor n8482 n8492 ; n8493
g8302 and asqrt[32] n8493_not ; n8494
g8303 and n8031_not n8037 ; n8495
g8304 and n8039_not n8495 ; n8496
g8305 and asqrt[27] n8496 ; n8497
g8306 nor n8031 n8039 ; n8498
g8307 and asqrt[27] n8498 ; n8499
g8308 nor n8037 n8499 ; n8500
g8309 nor n8497 n8500 ; n8501
g8310 nor asqrt[32] n8482 ; n8502
g8311 and n8492_not n8502 ; n8503
g8312 nor n8501 n8503 ; n8504
g8313 nor n8494 n8504 ; n8505
g8314 and asqrt[33] n8505_not ; n8506
g8315 and n8049 n8051_not ; n8507
g8316 and n8042_not n8507 ; n8508
g8317 and asqrt[27] n8508 ; n8509
g8318 nor n8042 n8051 ; n8510
g8319 and asqrt[27] n8510 ; n8511
g8320 nor n8049 n8511 ; n8512
g8321 nor n8509 n8512 ; n8513
g8322 nor asqrt[33] n8494 ; n8514
g8323 and n8504_not n8514 ; n8515
g8324 nor n8513 n8515 ; n8516
g8325 nor n8506 n8516 ; n8517
g8326 and asqrt[34] n8517_not ; n8518
g8327 and n8054_not n8061 ; n8519
g8328 and n8063_not n8519 ; n8520
g8329 and asqrt[27] n8520 ; n8521
g8330 nor n8054 n8063 ; n8522
g8331 and asqrt[27] n8522 ; n8523
g8332 nor n8061 n8523 ; n8524
g8333 nor n8521 n8524 ; n8525
g8334 nor asqrt[34] n8506 ; n8526
g8335 and n8516_not n8526 ; n8527
g8336 nor n8525 n8527 ; n8528
g8337 nor n8518 n8528 ; n8529
g8338 and asqrt[35] n8529_not ; n8530
g8339 and n8073 n8075_not ; n8531
g8340 and n8066_not n8531 ; n8532
g8341 and asqrt[27] n8532 ; n8533
g8342 nor n8066 n8075 ; n8534
g8343 and asqrt[27] n8534 ; n8535
g8344 nor n8073 n8535 ; n8536
g8345 nor n8533 n8536 ; n8537
g8346 nor asqrt[35] n8518 ; n8538
g8347 and n8528_not n8538 ; n8539
g8348 nor n8537 n8539 ; n8540
g8349 nor n8530 n8540 ; n8541
g8350 and asqrt[36] n8541_not ; n8542
g8351 and n8078_not n8085 ; n8543
g8352 and n8087_not n8543 ; n8544
g8353 and asqrt[27] n8544 ; n8545
g8354 nor n8078 n8087 ; n8546
g8355 and asqrt[27] n8546 ; n8547
g8356 nor n8085 n8547 ; n8548
g8357 nor n8545 n8548 ; n8549
g8358 nor asqrt[36] n8530 ; n8550
g8359 and n8540_not n8550 ; n8551
g8360 nor n8549 n8551 ; n8552
g8361 nor n8542 n8552 ; n8553
g8362 and asqrt[37] n8553_not ; n8554
g8363 and n8097 n8099_not ; n8555
g8364 and n8090_not n8555 ; n8556
g8365 and asqrt[27] n8556 ; n8557
g8366 nor n8090 n8099 ; n8558
g8367 and asqrt[27] n8558 ; n8559
g8368 nor n8097 n8559 ; n8560
g8369 nor n8557 n8560 ; n8561
g8370 nor asqrt[37] n8542 ; n8562
g8371 and n8552_not n8562 ; n8563
g8372 nor n8561 n8563 ; n8564
g8373 nor n8554 n8564 ; n8565
g8374 and asqrt[38] n8565_not ; n8566
g8375 nor asqrt[38] n8554 ; n8567
g8376 and n8564_not n8567 ; n8568
g8377 and n8102_not n8111 ; n8569
g8378 and n8104_not n8569 ; n8570
g8379 and asqrt[27] n8570 ; n8571
g8380 nor n8102 n8104 ; n8572
g8381 and asqrt[27] n8572 ; n8573
g8382 nor n8111 n8573 ; n8574
g8383 nor n8571 n8574 ; n8575
g8384 nor n8568 n8575 ; n8576
g8385 nor n8566 n8576 ; n8577
g8386 and asqrt[39] n8577_not ; n8578
g8387 and n8121 n8123_not ; n8579
g8388 and n8114_not n8579 ; n8580
g8389 and asqrt[27] n8580 ; n8581
g8390 nor n8114 n8123 ; n8582
g8391 and asqrt[27] n8582 ; n8583
g8392 nor n8121 n8583 ; n8584
g8393 nor n8581 n8584 ; n8585
g8394 nor asqrt[39] n8566 ; n8586
g8395 and n8576_not n8586 ; n8587
g8396 nor n8585 n8587 ; n8588
g8397 nor n8578 n8588 ; n8589
g8398 and asqrt[40] n8589_not ; n8590
g8399 and n8126_not n8133 ; n8591
g8400 and n8135_not n8591 ; n8592
g8401 and asqrt[27] n8592 ; n8593
g8402 nor n8126 n8135 ; n8594
g8403 and asqrt[27] n8594 ; n8595
g8404 nor n8133 n8595 ; n8596
g8405 nor n8593 n8596 ; n8597
g8406 nor asqrt[40] n8578 ; n8598
g8407 and n8588_not n8598 ; n8599
g8408 nor n8597 n8599 ; n8600
g8409 nor n8590 n8600 ; n8601
g8410 and asqrt[41] n8601_not ; n8602
g8411 and n8145 n8147_not ; n8603
g8412 and n8138_not n8603 ; n8604
g8413 and asqrt[27] n8604 ; n8605
g8414 nor n8138 n8147 ; n8606
g8415 and asqrt[27] n8606 ; n8607
g8416 nor n8145 n8607 ; n8608
g8417 nor n8605 n8608 ; n8609
g8418 nor asqrt[41] n8590 ; n8610
g8419 and n8600_not n8610 ; n8611
g8420 nor n8609 n8611 ; n8612
g8421 nor n8602 n8612 ; n8613
g8422 and asqrt[42] n8613_not ; n8614
g8423 and n8150_not n8157 ; n8615
g8424 and n8159_not n8615 ; n8616
g8425 and asqrt[27] n8616 ; n8617
g8426 nor n8150 n8159 ; n8618
g8427 and asqrt[27] n8618 ; n8619
g8428 nor n8157 n8619 ; n8620
g8429 nor n8617 n8620 ; n8621
g8430 nor asqrt[42] n8602 ; n8622
g8431 and n8612_not n8622 ; n8623
g8432 nor n8621 n8623 ; n8624
g8433 nor n8614 n8624 ; n8625
g8434 and asqrt[43] n8625_not ; n8626
g8435 and n8169 n8171_not ; n8627
g8436 and n8162_not n8627 ; n8628
g8437 and asqrt[27] n8628 ; n8629
g8438 nor n8162 n8171 ; n8630
g8439 and asqrt[27] n8630 ; n8631
g8440 nor n8169 n8631 ; n8632
g8441 nor n8629 n8632 ; n8633
g8442 nor asqrt[43] n8614 ; n8634
g8443 and n8624_not n8634 ; n8635
g8444 nor n8633 n8635 ; n8636
g8445 nor n8626 n8636 ; n8637
g8446 and asqrt[44] n8637_not ; n8638
g8447 and n8174_not n8181 ; n8639
g8448 and n8183_not n8639 ; n8640
g8449 and asqrt[27] n8640 ; n8641
g8450 nor n8174 n8183 ; n8642
g8451 and asqrt[27] n8642 ; n8643
g8452 nor n8181 n8643 ; n8644
g8453 nor n8641 n8644 ; n8645
g8454 nor asqrt[44] n8626 ; n8646
g8455 and n8636_not n8646 ; n8647
g8456 nor n8645 n8647 ; n8648
g8457 nor n8638 n8648 ; n8649
g8458 and asqrt[45] n8649_not ; n8650
g8459 and n8193 n8195_not ; n8651
g8460 and n8186_not n8651 ; n8652
g8461 and asqrt[27] n8652 ; n8653
g8462 nor n8186 n8195 ; n8654
g8463 and asqrt[27] n8654 ; n8655
g8464 nor n8193 n8655 ; n8656
g8465 nor n8653 n8656 ; n8657
g8466 nor asqrt[45] n8638 ; n8658
g8467 and n8648_not n8658 ; n8659
g8468 nor n8657 n8659 ; n8660
g8469 nor n8650 n8660 ; n8661
g8470 and asqrt[46] n8661_not ; n8662
g8471 and n8198_not n8205 ; n8663
g8472 and n8207_not n8663 ; n8664
g8473 and asqrt[27] n8664 ; n8665
g8474 nor n8198 n8207 ; n8666
g8475 and asqrt[27] n8666 ; n8667
g8476 nor n8205 n8667 ; n8668
g8477 nor n8665 n8668 ; n8669
g8478 nor asqrt[46] n8650 ; n8670
g8479 and n8660_not n8670 ; n8671
g8480 nor n8669 n8671 ; n8672
g8481 nor n8662 n8672 ; n8673
g8482 and asqrt[47] n8673_not ; n8674
g8483 and n8217 n8219_not ; n8675
g8484 and n8210_not n8675 ; n8676
g8485 and asqrt[27] n8676 ; n8677
g8486 nor n8210 n8219 ; n8678
g8487 and asqrt[27] n8678 ; n8679
g8488 nor n8217 n8679 ; n8680
g8489 nor n8677 n8680 ; n8681
g8490 nor asqrt[47] n8662 ; n8682
g8491 and n8672_not n8682 ; n8683
g8492 nor n8681 n8683 ; n8684
g8493 nor n8674 n8684 ; n8685
g8494 and asqrt[48] n8685_not ; n8686
g8495 and n8222_not n8229 ; n8687
g8496 and n8231_not n8687 ; n8688
g8497 and asqrt[27] n8688 ; n8689
g8498 nor n8222 n8231 ; n8690
g8499 and asqrt[27] n8690 ; n8691
g8500 nor n8229 n8691 ; n8692
g8501 nor n8689 n8692 ; n8693
g8502 nor asqrt[48] n8674 ; n8694
g8503 and n8684_not n8694 ; n8695
g8504 nor n8693 n8695 ; n8696
g8505 nor n8686 n8696 ; n8697
g8506 and asqrt[49] n8697_not ; n8698
g8507 and n8241 n8243_not ; n8699
g8508 and n8234_not n8699 ; n8700
g8509 and asqrt[27] n8700 ; n8701
g8510 nor n8234 n8243 ; n8702
g8511 and asqrt[27] n8702 ; n8703
g8512 nor n8241 n8703 ; n8704
g8513 nor n8701 n8704 ; n8705
g8514 nor asqrt[49] n8686 ; n8706
g8515 and n8696_not n8706 ; n8707
g8516 nor n8705 n8707 ; n8708
g8517 nor n8698 n8708 ; n8709
g8518 and asqrt[50] n8709_not ; n8710
g8519 and n8246_not n8253 ; n8711
g8520 and n8255_not n8711 ; n8712
g8521 and asqrt[27] n8712 ; n8713
g8522 nor n8246 n8255 ; n8714
g8523 and asqrt[27] n8714 ; n8715
g8524 nor n8253 n8715 ; n8716
g8525 nor n8713 n8716 ; n8717
g8526 nor asqrt[50] n8698 ; n8718
g8527 and n8708_not n8718 ; n8719
g8528 nor n8717 n8719 ; n8720
g8529 nor n8710 n8720 ; n8721
g8530 and asqrt[51] n8721_not ; n8722
g8531 and n8265 n8267_not ; n8723
g8532 and n8258_not n8723 ; n8724
g8533 and asqrt[27] n8724 ; n8725
g8534 nor n8258 n8267 ; n8726
g8535 and asqrt[27] n8726 ; n8727
g8536 nor n8265 n8727 ; n8728
g8537 nor n8725 n8728 ; n8729
g8538 nor asqrt[51] n8710 ; n8730
g8539 and n8720_not n8730 ; n8731
g8540 nor n8729 n8731 ; n8732
g8541 nor n8722 n8732 ; n8733
g8542 and asqrt[52] n8733_not ; n8734
g8543 and n8270_not n8277 ; n8735
g8544 and n8279_not n8735 ; n8736
g8545 and asqrt[27] n8736 ; n8737
g8546 nor n8270 n8279 ; n8738
g8547 and asqrt[27] n8738 ; n8739
g8548 nor n8277 n8739 ; n8740
g8549 nor n8737 n8740 ; n8741
g8550 nor asqrt[52] n8722 ; n8742
g8551 and n8732_not n8742 ; n8743
g8552 nor n8741 n8743 ; n8744
g8553 nor n8734 n8744 ; n8745
g8554 and asqrt[53] n8745_not ; n8746
g8555 and n8289 n8291_not ; n8747
g8556 and n8282_not n8747 ; n8748
g8557 and asqrt[27] n8748 ; n8749
g8558 nor n8282 n8291 ; n8750
g8559 and asqrt[27] n8750 ; n8751
g8560 nor n8289 n8751 ; n8752
g8561 nor n8749 n8752 ; n8753
g8562 nor asqrt[53] n8734 ; n8754
g8563 and n8744_not n8754 ; n8755
g8564 nor n8753 n8755 ; n8756
g8565 nor n8746 n8756 ; n8757
g8566 and asqrt[54] n8757_not ; n8758
g8567 and n8294_not n8301 ; n8759
g8568 and n8303_not n8759 ; n8760
g8569 and asqrt[27] n8760 ; n8761
g8570 nor n8294 n8303 ; n8762
g8571 and asqrt[27] n8762 ; n8763
g8572 nor n8301 n8763 ; n8764
g8573 nor n8761 n8764 ; n8765
g8574 nor asqrt[54] n8746 ; n8766
g8575 and n8756_not n8766 ; n8767
g8576 nor n8765 n8767 ; n8768
g8577 nor n8758 n8768 ; n8769
g8578 and asqrt[55] n8769_not ; n8770
g8579 and n8313 n8315_not ; n8771
g8580 and n8306_not n8771 ; n8772
g8581 and asqrt[27] n8772 ; n8773
g8582 nor n8306 n8315 ; n8774
g8583 and asqrt[27] n8774 ; n8775
g8584 nor n8313 n8775 ; n8776
g8585 nor n8773 n8776 ; n8777
g8586 nor asqrt[55] n8758 ; n8778
g8587 and n8768_not n8778 ; n8779
g8588 nor n8777 n8779 ; n8780
g8589 nor n8770 n8780 ; n8781
g8590 and asqrt[56] n8781_not ; n8782
g8591 and n8318_not n8325 ; n8783
g8592 and n8327_not n8783 ; n8784
g8593 and asqrt[27] n8784 ; n8785
g8594 nor n8318 n8327 ; n8786
g8595 and asqrt[27] n8786 ; n8787
g8596 nor n8325 n8787 ; n8788
g8597 nor n8785 n8788 ; n8789
g8598 nor asqrt[56] n8770 ; n8790
g8599 and n8780_not n8790 ; n8791
g8600 nor n8789 n8791 ; n8792
g8601 nor n8782 n8792 ; n8793
g8602 and asqrt[57] n8793_not ; n8794
g8603 and n8337 n8339_not ; n8795
g8604 and n8330_not n8795 ; n8796
g8605 and asqrt[27] n8796 ; n8797
g8606 nor n8330 n8339 ; n8798
g8607 and asqrt[27] n8798 ; n8799
g8608 nor n8337 n8799 ; n8800
g8609 nor n8797 n8800 ; n8801
g8610 nor asqrt[57] n8782 ; n8802
g8611 and n8792_not n8802 ; n8803
g8612 nor n8801 n8803 ; n8804
g8613 nor n8794 n8804 ; n8805
g8614 and asqrt[58] n8805_not ; n8806
g8615 and n8342_not n8349 ; n8807
g8616 and n8351_not n8807 ; n8808
g8617 and asqrt[27] n8808 ; n8809
g8618 nor n8342 n8351 ; n8810
g8619 and asqrt[27] n8810 ; n8811
g8620 nor n8349 n8811 ; n8812
g8621 nor n8809 n8812 ; n8813
g8622 nor asqrt[58] n8794 ; n8814
g8623 and n8804_not n8814 ; n8815
g8624 nor n8813 n8815 ; n8816
g8625 nor n8806 n8816 ; n8817
g8626 and asqrt[59] n8817_not ; n8818
g8627 and n8361 n8363_not ; n8819
g8628 and n8354_not n8819 ; n8820
g8629 and asqrt[27] n8820 ; n8821
g8630 nor n8354 n8363 ; n8822
g8631 and asqrt[27] n8822 ; n8823
g8632 nor n8361 n8823 ; n8824
g8633 nor n8821 n8824 ; n8825
g8634 nor asqrt[59] n8806 ; n8826
g8635 and n8816_not n8826 ; n8827
g8636 nor n8825 n8827 ; n8828
g8637 nor n8818 n8828 ; n8829
g8638 and asqrt[60] n8829_not ; n8830
g8639 and n8366_not n8373 ; n8831
g8640 and n8375_not n8831 ; n8832
g8641 and asqrt[27] n8832 ; n8833
g8642 nor n8366 n8375 ; n8834
g8643 and asqrt[27] n8834 ; n8835
g8644 nor n8373 n8835 ; n8836
g8645 nor n8833 n8836 ; n8837
g8646 nor asqrt[60] n8818 ; n8838
g8647 and n8828_not n8838 ; n8839
g8648 nor n8837 n8839 ; n8840
g8649 nor n8830 n8840 ; n8841
g8650 and asqrt[61] n8841_not ; n8842
g8651 and n8385 n8387_not ; n8843
g8652 and n8378_not n8843 ; n8844
g8653 and asqrt[27] n8844 ; n8845
g8654 nor n8378 n8387 ; n8846
g8655 and asqrt[27] n8846 ; n8847
g8656 nor n8385 n8847 ; n8848
g8657 nor n8845 n8848 ; n8849
g8658 nor asqrt[61] n8830 ; n8850
g8659 and n8840_not n8850 ; n8851
g8660 nor n8849 n8851 ; n8852
g8661 nor n8842 n8852 ; n8853
g8662 and asqrt[62] n8853_not ; n8854
g8663 and n8390_not n8397 ; n8855
g8664 and n8399_not n8855 ; n8856
g8665 and asqrt[27] n8856 ; n8857
g8666 nor n8390 n8399 ; n8858
g8667 and asqrt[27] n8858 ; n8859
g8668 nor n8397 n8859 ; n8860
g8669 nor n8857 n8860 ; n8861
g8670 nor asqrt[62] n8842 ; n8862
g8671 and n8852_not n8862 ; n8863
g8672 nor n8861 n8863 ; n8864
g8673 nor n8854 n8864 ; n8865
g8674 and n8409 n8411_not ; n8866
g8675 and n8402_not n8866 ; n8867
g8676 and asqrt[27] n8867 ; n8868
g8677 nor n8402 n8411 ; n8869
g8678 and asqrt[27] n8869 ; n8870
g8679 nor n8409 n8870 ; n8871
g8680 nor n8868 n8871 ; n8872
g8681 nor n8413 n8420 ; n8873
g8682 and asqrt[27] n8873 ; n8874
g8683 nor n8428 n8874 ; n8875
g8684 and n8872_not n8875 ; n8876
g8685 and n8865_not n8876 ; n8877
g8686 nor asqrt[63] n8877 ; n8878
g8687 and n8854_not n8872 ; n8879
g8688 and n8864_not n8879 ; n8880
g8689 and n8420_not asqrt[27] ; n8881
g8690 and n8413 n8881_not ; n8882
g8691 and asqrt[63] n8873_not ; n8883
g8692 and n8882_not n8883 ; n8884
g8693 nor n8416 n8437 ; n8885
g8694 and n8419_not n8885 ; n8886
g8695 and n8432_not n8886 ; n8887
g8696 and n8428_not n8887 ; n8888
g8697 and n8426_not n8888 ; n8889
g8698 nor n8884 n8889 ; n8890
g8699 and n8880_not n8890 ; n8891
g8700 nand n8878_not n8891 ; asqrt[26]
g8701 and a[52] asqrt[26] ; n8893
g8702 nor a[50] a[51] ; n8894
g8703 and a[52]_not n8894 ; n8895
g8704 nor n8893 n8895 ; n8896
g8705 and asqrt[27] n8896_not ; n8897
g8706 nor n8437 n8895 ; n8898
g8707 and n8432_not n8898 ; n8899
g8708 and n8428_not n8899 ; n8900
g8709 and n8426_not n8900 ; n8901
g8710 and n8893_not n8901 ; n8902
g8711 and a[52]_not asqrt[26] ; n8903
g8712 and a[53] n8903_not ; n8904
g8713 and n8442 asqrt[26] ; n8905
g8714 nor n8904 n8905 ; n8906
g8715 and n8902_not n8906 ; n8907
g8716 nor n8897 n8907 ; n8908
g8717 and asqrt[28] n8908_not ; n8909
g8718 nor asqrt[28] n8897 ; n8910
g8719 and n8907_not n8910 ; n8911
g8720 and asqrt[27] n8889_not ; n8912
g8721 and n8884_not n8912 ; n8913
g8722 and n8880_not n8913 ; n8914
g8723 and n8878_not n8914 ; n8915
g8724 nor n8905 n8915 ; n8916
g8725 and a[54] n8916_not ; n8917
g8726 nor a[54] n8915 ; n8918
g8727 and n8905_not n8918 ; n8919
g8728 nor n8917 n8919 ; n8920
g8729 nor n8911 n8920 ; n8921
g8730 nor n8909 n8921 ; n8922
g8731 and asqrt[29] n8922_not ; n8923
g8732 nor n8445 n8450 ; n8924
g8733 and n8454_not n8924 ; n8925
g8734 and asqrt[26] n8925 ; n8926
g8735 and asqrt[26] n8924 ; n8927
g8736 and n8454 n8927_not ; n8928
g8737 nor n8926 n8928 ; n8929
g8738 nor asqrt[29] n8909 ; n8930
g8739 and n8921_not n8930 ; n8931
g8740 nor n8929 n8931 ; n8932
g8741 nor n8923 n8932 ; n8933
g8742 and asqrt[30] n8933_not ; n8934
g8743 and n8459_not n8468 ; n8935
g8744 and n8457_not n8935 ; n8936
g8745 and asqrt[26] n8936 ; n8937
g8746 nor n8457 n8459 ; n8938
g8747 and asqrt[26] n8938 ; n8939
g8748 nor n8468 n8939 ; n8940
g8749 nor n8937 n8940 ; n8941
g8750 nor asqrt[30] n8923 ; n8942
g8751 and n8932_not n8942 ; n8943
g8752 nor n8941 n8943 ; n8944
g8753 nor n8934 n8944 ; n8945
g8754 and asqrt[31] n8945_not ; n8946
g8755 and n8471_not n8477 ; n8947
g8756 and n8479_not n8947 ; n8948
g8757 and asqrt[26] n8948 ; n8949
g8758 nor n8471 n8479 ; n8950
g8759 and asqrt[26] n8950 ; n8951
g8760 nor n8477 n8951 ; n8952
g8761 nor n8949 n8952 ; n8953
g8762 nor asqrt[31] n8934 ; n8954
g8763 and n8944_not n8954 ; n8955
g8764 nor n8953 n8955 ; n8956
g8765 nor n8946 n8956 ; n8957
g8766 and asqrt[32] n8957_not ; n8958
g8767 and n8489 n8491_not ; n8959
g8768 and n8482_not n8959 ; n8960
g8769 and asqrt[26] n8960 ; n8961
g8770 nor n8482 n8491 ; n8962
g8771 and asqrt[26] n8962 ; n8963
g8772 nor n8489 n8963 ; n8964
g8773 nor n8961 n8964 ; n8965
g8774 nor asqrt[32] n8946 ; n8966
g8775 and n8956_not n8966 ; n8967
g8776 nor n8965 n8967 ; n8968
g8777 nor n8958 n8968 ; n8969
g8778 and asqrt[33] n8969_not ; n8970
g8779 and n8494_not n8501 ; n8971
g8780 and n8503_not n8971 ; n8972
g8781 and asqrt[26] n8972 ; n8973
g8782 nor n8494 n8503 ; n8974
g8783 and asqrt[26] n8974 ; n8975
g8784 nor n8501 n8975 ; n8976
g8785 nor n8973 n8976 ; n8977
g8786 nor asqrt[33] n8958 ; n8978
g8787 and n8968_not n8978 ; n8979
g8788 nor n8977 n8979 ; n8980
g8789 nor n8970 n8980 ; n8981
g8790 and asqrt[34] n8981_not ; n8982
g8791 and n8513 n8515_not ; n8983
g8792 and n8506_not n8983 ; n8984
g8793 and asqrt[26] n8984 ; n8985
g8794 nor n8506 n8515 ; n8986
g8795 and asqrt[26] n8986 ; n8987
g8796 nor n8513 n8987 ; n8988
g8797 nor n8985 n8988 ; n8989
g8798 nor asqrt[34] n8970 ; n8990
g8799 and n8980_not n8990 ; n8991
g8800 nor n8989 n8991 ; n8992
g8801 nor n8982 n8992 ; n8993
g8802 and asqrt[35] n8993_not ; n8994
g8803 and n8518_not n8525 ; n8995
g8804 and n8527_not n8995 ; n8996
g8805 and asqrt[26] n8996 ; n8997
g8806 nor n8518 n8527 ; n8998
g8807 and asqrt[26] n8998 ; n8999
g8808 nor n8525 n8999 ; n9000
g8809 nor n8997 n9000 ; n9001
g8810 nor asqrt[35] n8982 ; n9002
g8811 and n8992_not n9002 ; n9003
g8812 nor n9001 n9003 ; n9004
g8813 nor n8994 n9004 ; n9005
g8814 and asqrt[36] n9005_not ; n9006
g8815 and n8537 n8539_not ; n9007
g8816 and n8530_not n9007 ; n9008
g8817 and asqrt[26] n9008 ; n9009
g8818 nor n8530 n8539 ; n9010
g8819 and asqrt[26] n9010 ; n9011
g8820 nor n8537 n9011 ; n9012
g8821 nor n9009 n9012 ; n9013
g8822 nor asqrt[36] n8994 ; n9014
g8823 and n9004_not n9014 ; n9015
g8824 nor n9013 n9015 ; n9016
g8825 nor n9006 n9016 ; n9017
g8826 and asqrt[37] n9017_not ; n9018
g8827 and n8542_not n8549 ; n9019
g8828 and n8551_not n9019 ; n9020
g8829 and asqrt[26] n9020 ; n9021
g8830 nor n8542 n8551 ; n9022
g8831 and asqrt[26] n9022 ; n9023
g8832 nor n8549 n9023 ; n9024
g8833 nor n9021 n9024 ; n9025
g8834 nor asqrt[37] n9006 ; n9026
g8835 and n9016_not n9026 ; n9027
g8836 nor n9025 n9027 ; n9028
g8837 nor n9018 n9028 ; n9029
g8838 and asqrt[38] n9029_not ; n9030
g8839 and n8561 n8563_not ; n9031
g8840 and n8554_not n9031 ; n9032
g8841 and asqrt[26] n9032 ; n9033
g8842 nor n8554 n8563 ; n9034
g8843 and asqrt[26] n9034 ; n9035
g8844 nor n8561 n9035 ; n9036
g8845 nor n9033 n9036 ; n9037
g8846 nor asqrt[38] n9018 ; n9038
g8847 and n9028_not n9038 ; n9039
g8848 nor n9037 n9039 ; n9040
g8849 nor n9030 n9040 ; n9041
g8850 and asqrt[39] n9041_not ; n9042
g8851 nor asqrt[39] n9030 ; n9043
g8852 and n9040_not n9043 ; n9044
g8853 and n8566_not n8575 ; n9045
g8854 and n8568_not n9045 ; n9046
g8855 and asqrt[26] n9046 ; n9047
g8856 nor n8566 n8568 ; n9048
g8857 and asqrt[26] n9048 ; n9049
g8858 nor n8575 n9049 ; n9050
g8859 nor n9047 n9050 ; n9051
g8860 nor n9044 n9051 ; n9052
g8861 nor n9042 n9052 ; n9053
g8862 and asqrt[40] n9053_not ; n9054
g8863 and n8585 n8587_not ; n9055
g8864 and n8578_not n9055 ; n9056
g8865 and asqrt[26] n9056 ; n9057
g8866 nor n8578 n8587 ; n9058
g8867 and asqrt[26] n9058 ; n9059
g8868 nor n8585 n9059 ; n9060
g8869 nor n9057 n9060 ; n9061
g8870 nor asqrt[40] n9042 ; n9062
g8871 and n9052_not n9062 ; n9063
g8872 nor n9061 n9063 ; n9064
g8873 nor n9054 n9064 ; n9065
g8874 and asqrt[41] n9065_not ; n9066
g8875 and n8590_not n8597 ; n9067
g8876 and n8599_not n9067 ; n9068
g8877 and asqrt[26] n9068 ; n9069
g8878 nor n8590 n8599 ; n9070
g8879 and asqrt[26] n9070 ; n9071
g8880 nor n8597 n9071 ; n9072
g8881 nor n9069 n9072 ; n9073
g8882 nor asqrt[41] n9054 ; n9074
g8883 and n9064_not n9074 ; n9075
g8884 nor n9073 n9075 ; n9076
g8885 nor n9066 n9076 ; n9077
g8886 and asqrt[42] n9077_not ; n9078
g8887 and n8609 n8611_not ; n9079
g8888 and n8602_not n9079 ; n9080
g8889 and asqrt[26] n9080 ; n9081
g8890 nor n8602 n8611 ; n9082
g8891 and asqrt[26] n9082 ; n9083
g8892 nor n8609 n9083 ; n9084
g8893 nor n9081 n9084 ; n9085
g8894 nor asqrt[42] n9066 ; n9086
g8895 and n9076_not n9086 ; n9087
g8896 nor n9085 n9087 ; n9088
g8897 nor n9078 n9088 ; n9089
g8898 and asqrt[43] n9089_not ; n9090
g8899 and n8614_not n8621 ; n9091
g8900 and n8623_not n9091 ; n9092
g8901 and asqrt[26] n9092 ; n9093
g8902 nor n8614 n8623 ; n9094
g8903 and asqrt[26] n9094 ; n9095
g8904 nor n8621 n9095 ; n9096
g8905 nor n9093 n9096 ; n9097
g8906 nor asqrt[43] n9078 ; n9098
g8907 and n9088_not n9098 ; n9099
g8908 nor n9097 n9099 ; n9100
g8909 nor n9090 n9100 ; n9101
g8910 and asqrt[44] n9101_not ; n9102
g8911 and n8633 n8635_not ; n9103
g8912 and n8626_not n9103 ; n9104
g8913 and asqrt[26] n9104 ; n9105
g8914 nor n8626 n8635 ; n9106
g8915 and asqrt[26] n9106 ; n9107
g8916 nor n8633 n9107 ; n9108
g8917 nor n9105 n9108 ; n9109
g8918 nor asqrt[44] n9090 ; n9110
g8919 and n9100_not n9110 ; n9111
g8920 nor n9109 n9111 ; n9112
g8921 nor n9102 n9112 ; n9113
g8922 and asqrt[45] n9113_not ; n9114
g8923 and n8638_not n8645 ; n9115
g8924 and n8647_not n9115 ; n9116
g8925 and asqrt[26] n9116 ; n9117
g8926 nor n8638 n8647 ; n9118
g8927 and asqrt[26] n9118 ; n9119
g8928 nor n8645 n9119 ; n9120
g8929 nor n9117 n9120 ; n9121
g8930 nor asqrt[45] n9102 ; n9122
g8931 and n9112_not n9122 ; n9123
g8932 nor n9121 n9123 ; n9124
g8933 nor n9114 n9124 ; n9125
g8934 and asqrt[46] n9125_not ; n9126
g8935 and n8657 n8659_not ; n9127
g8936 and n8650_not n9127 ; n9128
g8937 and asqrt[26] n9128 ; n9129
g8938 nor n8650 n8659 ; n9130
g8939 and asqrt[26] n9130 ; n9131
g8940 nor n8657 n9131 ; n9132
g8941 nor n9129 n9132 ; n9133
g8942 nor asqrt[46] n9114 ; n9134
g8943 and n9124_not n9134 ; n9135
g8944 nor n9133 n9135 ; n9136
g8945 nor n9126 n9136 ; n9137
g8946 and asqrt[47] n9137_not ; n9138
g8947 and n8662_not n8669 ; n9139
g8948 and n8671_not n9139 ; n9140
g8949 and asqrt[26] n9140 ; n9141
g8950 nor n8662 n8671 ; n9142
g8951 and asqrt[26] n9142 ; n9143
g8952 nor n8669 n9143 ; n9144
g8953 nor n9141 n9144 ; n9145
g8954 nor asqrt[47] n9126 ; n9146
g8955 and n9136_not n9146 ; n9147
g8956 nor n9145 n9147 ; n9148
g8957 nor n9138 n9148 ; n9149
g8958 and asqrt[48] n9149_not ; n9150
g8959 and n8681 n8683_not ; n9151
g8960 and n8674_not n9151 ; n9152
g8961 and asqrt[26] n9152 ; n9153
g8962 nor n8674 n8683 ; n9154
g8963 and asqrt[26] n9154 ; n9155
g8964 nor n8681 n9155 ; n9156
g8965 nor n9153 n9156 ; n9157
g8966 nor asqrt[48] n9138 ; n9158
g8967 and n9148_not n9158 ; n9159
g8968 nor n9157 n9159 ; n9160
g8969 nor n9150 n9160 ; n9161
g8970 and asqrt[49] n9161_not ; n9162
g8971 and n8686_not n8693 ; n9163
g8972 and n8695_not n9163 ; n9164
g8973 and asqrt[26] n9164 ; n9165
g8974 nor n8686 n8695 ; n9166
g8975 and asqrt[26] n9166 ; n9167
g8976 nor n8693 n9167 ; n9168
g8977 nor n9165 n9168 ; n9169
g8978 nor asqrt[49] n9150 ; n9170
g8979 and n9160_not n9170 ; n9171
g8980 nor n9169 n9171 ; n9172
g8981 nor n9162 n9172 ; n9173
g8982 and asqrt[50] n9173_not ; n9174
g8983 and n8705 n8707_not ; n9175
g8984 and n8698_not n9175 ; n9176
g8985 and asqrt[26] n9176 ; n9177
g8986 nor n8698 n8707 ; n9178
g8987 and asqrt[26] n9178 ; n9179
g8988 nor n8705 n9179 ; n9180
g8989 nor n9177 n9180 ; n9181
g8990 nor asqrt[50] n9162 ; n9182
g8991 and n9172_not n9182 ; n9183
g8992 nor n9181 n9183 ; n9184
g8993 nor n9174 n9184 ; n9185
g8994 and asqrt[51] n9185_not ; n9186
g8995 and n8710_not n8717 ; n9187
g8996 and n8719_not n9187 ; n9188
g8997 and asqrt[26] n9188 ; n9189
g8998 nor n8710 n8719 ; n9190
g8999 and asqrt[26] n9190 ; n9191
g9000 nor n8717 n9191 ; n9192
g9001 nor n9189 n9192 ; n9193
g9002 nor asqrt[51] n9174 ; n9194
g9003 and n9184_not n9194 ; n9195
g9004 nor n9193 n9195 ; n9196
g9005 nor n9186 n9196 ; n9197
g9006 and asqrt[52] n9197_not ; n9198
g9007 and n8729 n8731_not ; n9199
g9008 and n8722_not n9199 ; n9200
g9009 and asqrt[26] n9200 ; n9201
g9010 nor n8722 n8731 ; n9202
g9011 and asqrt[26] n9202 ; n9203
g9012 nor n8729 n9203 ; n9204
g9013 nor n9201 n9204 ; n9205
g9014 nor asqrt[52] n9186 ; n9206
g9015 and n9196_not n9206 ; n9207
g9016 nor n9205 n9207 ; n9208
g9017 nor n9198 n9208 ; n9209
g9018 and asqrt[53] n9209_not ; n9210
g9019 and n8734_not n8741 ; n9211
g9020 and n8743_not n9211 ; n9212
g9021 and asqrt[26] n9212 ; n9213
g9022 nor n8734 n8743 ; n9214
g9023 and asqrt[26] n9214 ; n9215
g9024 nor n8741 n9215 ; n9216
g9025 nor n9213 n9216 ; n9217
g9026 nor asqrt[53] n9198 ; n9218
g9027 and n9208_not n9218 ; n9219
g9028 nor n9217 n9219 ; n9220
g9029 nor n9210 n9220 ; n9221
g9030 and asqrt[54] n9221_not ; n9222
g9031 and n8753 n8755_not ; n9223
g9032 and n8746_not n9223 ; n9224
g9033 and asqrt[26] n9224 ; n9225
g9034 nor n8746 n8755 ; n9226
g9035 and asqrt[26] n9226 ; n9227
g9036 nor n8753 n9227 ; n9228
g9037 nor n9225 n9228 ; n9229
g9038 nor asqrt[54] n9210 ; n9230
g9039 and n9220_not n9230 ; n9231
g9040 nor n9229 n9231 ; n9232
g9041 nor n9222 n9232 ; n9233
g9042 and asqrt[55] n9233_not ; n9234
g9043 and n8758_not n8765 ; n9235
g9044 and n8767_not n9235 ; n9236
g9045 and asqrt[26] n9236 ; n9237
g9046 nor n8758 n8767 ; n9238
g9047 and asqrt[26] n9238 ; n9239
g9048 nor n8765 n9239 ; n9240
g9049 nor n9237 n9240 ; n9241
g9050 nor asqrt[55] n9222 ; n9242
g9051 and n9232_not n9242 ; n9243
g9052 nor n9241 n9243 ; n9244
g9053 nor n9234 n9244 ; n9245
g9054 and asqrt[56] n9245_not ; n9246
g9055 and n8777 n8779_not ; n9247
g9056 and n8770_not n9247 ; n9248
g9057 and asqrt[26] n9248 ; n9249
g9058 nor n8770 n8779 ; n9250
g9059 and asqrt[26] n9250 ; n9251
g9060 nor n8777 n9251 ; n9252
g9061 nor n9249 n9252 ; n9253
g9062 nor asqrt[56] n9234 ; n9254
g9063 and n9244_not n9254 ; n9255
g9064 nor n9253 n9255 ; n9256
g9065 nor n9246 n9256 ; n9257
g9066 and asqrt[57] n9257_not ; n9258
g9067 and n8782_not n8789 ; n9259
g9068 and n8791_not n9259 ; n9260
g9069 and asqrt[26] n9260 ; n9261
g9070 nor n8782 n8791 ; n9262
g9071 and asqrt[26] n9262 ; n9263
g9072 nor n8789 n9263 ; n9264
g9073 nor n9261 n9264 ; n9265
g9074 nor asqrt[57] n9246 ; n9266
g9075 and n9256_not n9266 ; n9267
g9076 nor n9265 n9267 ; n9268
g9077 nor n9258 n9268 ; n9269
g9078 and asqrt[58] n9269_not ; n9270
g9079 and n8801 n8803_not ; n9271
g9080 and n8794_not n9271 ; n9272
g9081 and asqrt[26] n9272 ; n9273
g9082 nor n8794 n8803 ; n9274
g9083 and asqrt[26] n9274 ; n9275
g9084 nor n8801 n9275 ; n9276
g9085 nor n9273 n9276 ; n9277
g9086 nor asqrt[58] n9258 ; n9278
g9087 and n9268_not n9278 ; n9279
g9088 nor n9277 n9279 ; n9280
g9089 nor n9270 n9280 ; n9281
g9090 and asqrt[59] n9281_not ; n9282
g9091 and n8806_not n8813 ; n9283
g9092 and n8815_not n9283 ; n9284
g9093 and asqrt[26] n9284 ; n9285
g9094 nor n8806 n8815 ; n9286
g9095 and asqrt[26] n9286 ; n9287
g9096 nor n8813 n9287 ; n9288
g9097 nor n9285 n9288 ; n9289
g9098 nor asqrt[59] n9270 ; n9290
g9099 and n9280_not n9290 ; n9291
g9100 nor n9289 n9291 ; n9292
g9101 nor n9282 n9292 ; n9293
g9102 and asqrt[60] n9293_not ; n9294
g9103 and n8825 n8827_not ; n9295
g9104 and n8818_not n9295 ; n9296
g9105 and asqrt[26] n9296 ; n9297
g9106 nor n8818 n8827 ; n9298
g9107 and asqrt[26] n9298 ; n9299
g9108 nor n8825 n9299 ; n9300
g9109 nor n9297 n9300 ; n9301
g9110 nor asqrt[60] n9282 ; n9302
g9111 and n9292_not n9302 ; n9303
g9112 nor n9301 n9303 ; n9304
g9113 nor n9294 n9304 ; n9305
g9114 and asqrt[61] n9305_not ; n9306
g9115 and n8830_not n8837 ; n9307
g9116 and n8839_not n9307 ; n9308
g9117 and asqrt[26] n9308 ; n9309
g9118 nor n8830 n8839 ; n9310
g9119 and asqrt[26] n9310 ; n9311
g9120 nor n8837 n9311 ; n9312
g9121 nor n9309 n9312 ; n9313
g9122 nor asqrt[61] n9294 ; n9314
g9123 and n9304_not n9314 ; n9315
g9124 nor n9313 n9315 ; n9316
g9125 nor n9306 n9316 ; n9317
g9126 and asqrt[62] n9317_not ; n9318
g9127 and n8849 n8851_not ; n9319
g9128 and n8842_not n9319 ; n9320
g9129 and asqrt[26] n9320 ; n9321
g9130 nor n8842 n8851 ; n9322
g9131 and asqrt[26] n9322 ; n9323
g9132 nor n8849 n9323 ; n9324
g9133 nor n9321 n9324 ; n9325
g9134 nor asqrt[62] n9306 ; n9326
g9135 and n9316_not n9326 ; n9327
g9136 nor n9325 n9327 ; n9328
g9137 nor n9318 n9328 ; n9329
g9138 and n8854_not n8861 ; n9330
g9139 and n8863_not n9330 ; n9331
g9140 and asqrt[26] n9331 ; n9332
g9141 nor n8854 n8863 ; n9333
g9142 and asqrt[26] n9333 ; n9334
g9143 nor n8861 n9334 ; n9335
g9144 nor n9332 n9335 ; n9336
g9145 nor n8865 n8872 ; n9337
g9146 and asqrt[26] n9337 ; n9338
g9147 nor n8880 n9338 ; n9339
g9148 and n9336_not n9339 ; n9340
g9149 and n9329_not n9340 ; n9341
g9150 nor asqrt[63] n9341 ; n9342
g9151 and n9318_not n9336 ; n9343
g9152 and n9328_not n9343 ; n9344
g9153 and n8872_not asqrt[26] ; n9345
g9154 and n8865 n9345_not ; n9346
g9155 and asqrt[63] n9337_not ; n9347
g9156 and n9346_not n9347 ; n9348
g9157 nor n8868 n8889 ; n9349
g9158 and n8871_not n9349 ; n9350
g9159 and n8884_not n9350 ; n9351
g9160 and n8880_not n9351 ; n9352
g9161 and n8878_not n9352 ; n9353
g9162 nor n9348 n9353 ; n9354
g9163 and n9344_not n9354 ; n9355
g9164 nand n9342_not n9355 ; asqrt[25]
g9165 and a[50] asqrt[25] ; n9357
g9166 nor a[48] a[49] ; n9358
g9167 and a[50]_not n9358 ; n9359
g9168 nor n9357 n9359 ; n9360
g9169 and asqrt[26] n9360_not ; n9361
g9170 nor n8889 n9359 ; n9362
g9171 and n8884_not n9362 ; n9363
g9172 and n8880_not n9363 ; n9364
g9173 and n8878_not n9364 ; n9365
g9174 and n9357_not n9365 ; n9366
g9175 and a[50]_not asqrt[25] ; n9367
g9176 and a[51] n9367_not ; n9368
g9177 and n8894 asqrt[25] ; n9369
g9178 nor n9368 n9369 ; n9370
g9179 and n9366_not n9370 ; n9371
g9180 nor n9361 n9371 ; n9372
g9181 and asqrt[27] n9372_not ; n9373
g9182 nor asqrt[27] n9361 ; n9374
g9183 and n9371_not n9374 ; n9375
g9184 and asqrt[26] n9353_not ; n9376
g9185 and n9348_not n9376 ; n9377
g9186 and n9344_not n9377 ; n9378
g9187 and n9342_not n9378 ; n9379
g9188 nor n9369 n9379 ; n9380
g9189 and a[52] n9380_not ; n9381
g9190 nor a[52] n9379 ; n9382
g9191 and n9369_not n9382 ; n9383
g9192 nor n9381 n9383 ; n9384
g9193 nor n9375 n9384 ; n9385
g9194 nor n9373 n9385 ; n9386
g9195 and asqrt[28] n9386_not ; n9387
g9196 nor n8897 n8902 ; n9388
g9197 and n8906_not n9388 ; n9389
g9198 and asqrt[25] n9389 ; n9390
g9199 and asqrt[25] n9388 ; n9391
g9200 and n8906 n9391_not ; n9392
g9201 nor n9390 n9392 ; n9393
g9202 nor asqrt[28] n9373 ; n9394
g9203 and n9385_not n9394 ; n9395
g9204 nor n9393 n9395 ; n9396
g9205 nor n9387 n9396 ; n9397
g9206 and asqrt[29] n9397_not ; n9398
g9207 and n8911_not n8920 ; n9399
g9208 and n8909_not n9399 ; n9400
g9209 and asqrt[25] n9400 ; n9401
g9210 nor n8909 n8911 ; n9402
g9211 and asqrt[25] n9402 ; n9403
g9212 nor n8920 n9403 ; n9404
g9213 nor n9401 n9404 ; n9405
g9214 nor asqrt[29] n9387 ; n9406
g9215 and n9396_not n9406 ; n9407
g9216 nor n9405 n9407 ; n9408
g9217 nor n9398 n9408 ; n9409
g9218 and asqrt[30] n9409_not ; n9410
g9219 and n8923_not n8929 ; n9411
g9220 and n8931_not n9411 ; n9412
g9221 and asqrt[25] n9412 ; n9413
g9222 nor n8923 n8931 ; n9414
g9223 and asqrt[25] n9414 ; n9415
g9224 nor n8929 n9415 ; n9416
g9225 nor n9413 n9416 ; n9417
g9226 nor asqrt[30] n9398 ; n9418
g9227 and n9408_not n9418 ; n9419
g9228 nor n9417 n9419 ; n9420
g9229 nor n9410 n9420 ; n9421
g9230 and asqrt[31] n9421_not ; n9422
g9231 and n8941 n8943_not ; n9423
g9232 and n8934_not n9423 ; n9424
g9233 and asqrt[25] n9424 ; n9425
g9234 nor n8934 n8943 ; n9426
g9235 and asqrt[25] n9426 ; n9427
g9236 nor n8941 n9427 ; n9428
g9237 nor n9425 n9428 ; n9429
g9238 nor asqrt[31] n9410 ; n9430
g9239 and n9420_not n9430 ; n9431
g9240 nor n9429 n9431 ; n9432
g9241 nor n9422 n9432 ; n9433
g9242 and asqrt[32] n9433_not ; n9434
g9243 and n8946_not n8953 ; n9435
g9244 and n8955_not n9435 ; n9436
g9245 and asqrt[25] n9436 ; n9437
g9246 nor n8946 n8955 ; n9438
g9247 and asqrt[25] n9438 ; n9439
g9248 nor n8953 n9439 ; n9440
g9249 nor n9437 n9440 ; n9441
g9250 nor asqrt[32] n9422 ; n9442
g9251 and n9432_not n9442 ; n9443
g9252 nor n9441 n9443 ; n9444
g9253 nor n9434 n9444 ; n9445
g9254 and asqrt[33] n9445_not ; n9446
g9255 and n8965 n8967_not ; n9447
g9256 and n8958_not n9447 ; n9448
g9257 and asqrt[25] n9448 ; n9449
g9258 nor n8958 n8967 ; n9450
g9259 and asqrt[25] n9450 ; n9451
g9260 nor n8965 n9451 ; n9452
g9261 nor n9449 n9452 ; n9453
g9262 nor asqrt[33] n9434 ; n9454
g9263 and n9444_not n9454 ; n9455
g9264 nor n9453 n9455 ; n9456
g9265 nor n9446 n9456 ; n9457
g9266 and asqrt[34] n9457_not ; n9458
g9267 and n8970_not n8977 ; n9459
g9268 and n8979_not n9459 ; n9460
g9269 and asqrt[25] n9460 ; n9461
g9270 nor n8970 n8979 ; n9462
g9271 and asqrt[25] n9462 ; n9463
g9272 nor n8977 n9463 ; n9464
g9273 nor n9461 n9464 ; n9465
g9274 nor asqrt[34] n9446 ; n9466
g9275 and n9456_not n9466 ; n9467
g9276 nor n9465 n9467 ; n9468
g9277 nor n9458 n9468 ; n9469
g9278 and asqrt[35] n9469_not ; n9470
g9279 and n8989 n8991_not ; n9471
g9280 and n8982_not n9471 ; n9472
g9281 and asqrt[25] n9472 ; n9473
g9282 nor n8982 n8991 ; n9474
g9283 and asqrt[25] n9474 ; n9475
g9284 nor n8989 n9475 ; n9476
g9285 nor n9473 n9476 ; n9477
g9286 nor asqrt[35] n9458 ; n9478
g9287 and n9468_not n9478 ; n9479
g9288 nor n9477 n9479 ; n9480
g9289 nor n9470 n9480 ; n9481
g9290 and asqrt[36] n9481_not ; n9482
g9291 and n8994_not n9001 ; n9483
g9292 and n9003_not n9483 ; n9484
g9293 and asqrt[25] n9484 ; n9485
g9294 nor n8994 n9003 ; n9486
g9295 and asqrt[25] n9486 ; n9487
g9296 nor n9001 n9487 ; n9488
g9297 nor n9485 n9488 ; n9489
g9298 nor asqrt[36] n9470 ; n9490
g9299 and n9480_not n9490 ; n9491
g9300 nor n9489 n9491 ; n9492
g9301 nor n9482 n9492 ; n9493
g9302 and asqrt[37] n9493_not ; n9494
g9303 and n9013 n9015_not ; n9495
g9304 and n9006_not n9495 ; n9496
g9305 and asqrt[25] n9496 ; n9497
g9306 nor n9006 n9015 ; n9498
g9307 and asqrt[25] n9498 ; n9499
g9308 nor n9013 n9499 ; n9500
g9309 nor n9497 n9500 ; n9501
g9310 nor asqrt[37] n9482 ; n9502
g9311 and n9492_not n9502 ; n9503
g9312 nor n9501 n9503 ; n9504
g9313 nor n9494 n9504 ; n9505
g9314 and asqrt[38] n9505_not ; n9506
g9315 and n9018_not n9025 ; n9507
g9316 and n9027_not n9507 ; n9508
g9317 and asqrt[25] n9508 ; n9509
g9318 nor n9018 n9027 ; n9510
g9319 and asqrt[25] n9510 ; n9511
g9320 nor n9025 n9511 ; n9512
g9321 nor n9509 n9512 ; n9513
g9322 nor asqrt[38] n9494 ; n9514
g9323 and n9504_not n9514 ; n9515
g9324 nor n9513 n9515 ; n9516
g9325 nor n9506 n9516 ; n9517
g9326 and asqrt[39] n9517_not ; n9518
g9327 and n9037 n9039_not ; n9519
g9328 and n9030_not n9519 ; n9520
g9329 and asqrt[25] n9520 ; n9521
g9330 nor n9030 n9039 ; n9522
g9331 and asqrt[25] n9522 ; n9523
g9332 nor n9037 n9523 ; n9524
g9333 nor n9521 n9524 ; n9525
g9334 nor asqrt[39] n9506 ; n9526
g9335 and n9516_not n9526 ; n9527
g9336 nor n9525 n9527 ; n9528
g9337 nor n9518 n9528 ; n9529
g9338 and asqrt[40] n9529_not ; n9530
g9339 nor asqrt[40] n9518 ; n9531
g9340 and n9528_not n9531 ; n9532
g9341 and n9042_not n9051 ; n9533
g9342 and n9044_not n9533 ; n9534
g9343 and asqrt[25] n9534 ; n9535
g9344 nor n9042 n9044 ; n9536
g9345 and asqrt[25] n9536 ; n9537
g9346 nor n9051 n9537 ; n9538
g9347 nor n9535 n9538 ; n9539
g9348 nor n9532 n9539 ; n9540
g9349 nor n9530 n9540 ; n9541
g9350 and asqrt[41] n9541_not ; n9542
g9351 and n9061 n9063_not ; n9543
g9352 and n9054_not n9543 ; n9544
g9353 and asqrt[25] n9544 ; n9545
g9354 nor n9054 n9063 ; n9546
g9355 and asqrt[25] n9546 ; n9547
g9356 nor n9061 n9547 ; n9548
g9357 nor n9545 n9548 ; n9549
g9358 nor asqrt[41] n9530 ; n9550
g9359 and n9540_not n9550 ; n9551
g9360 nor n9549 n9551 ; n9552
g9361 nor n9542 n9552 ; n9553
g9362 and asqrt[42] n9553_not ; n9554
g9363 and n9066_not n9073 ; n9555
g9364 and n9075_not n9555 ; n9556
g9365 and asqrt[25] n9556 ; n9557
g9366 nor n9066 n9075 ; n9558
g9367 and asqrt[25] n9558 ; n9559
g9368 nor n9073 n9559 ; n9560
g9369 nor n9557 n9560 ; n9561
g9370 nor asqrt[42] n9542 ; n9562
g9371 and n9552_not n9562 ; n9563
g9372 nor n9561 n9563 ; n9564
g9373 nor n9554 n9564 ; n9565
g9374 and asqrt[43] n9565_not ; n9566
g9375 and n9085 n9087_not ; n9567
g9376 and n9078_not n9567 ; n9568
g9377 and asqrt[25] n9568 ; n9569
g9378 nor n9078 n9087 ; n9570
g9379 and asqrt[25] n9570 ; n9571
g9380 nor n9085 n9571 ; n9572
g9381 nor n9569 n9572 ; n9573
g9382 nor asqrt[43] n9554 ; n9574
g9383 and n9564_not n9574 ; n9575
g9384 nor n9573 n9575 ; n9576
g9385 nor n9566 n9576 ; n9577
g9386 and asqrt[44] n9577_not ; n9578
g9387 and n9090_not n9097 ; n9579
g9388 and n9099_not n9579 ; n9580
g9389 and asqrt[25] n9580 ; n9581
g9390 nor n9090 n9099 ; n9582
g9391 and asqrt[25] n9582 ; n9583
g9392 nor n9097 n9583 ; n9584
g9393 nor n9581 n9584 ; n9585
g9394 nor asqrt[44] n9566 ; n9586
g9395 and n9576_not n9586 ; n9587
g9396 nor n9585 n9587 ; n9588
g9397 nor n9578 n9588 ; n9589
g9398 and asqrt[45] n9589_not ; n9590
g9399 and n9109 n9111_not ; n9591
g9400 and n9102_not n9591 ; n9592
g9401 and asqrt[25] n9592 ; n9593
g9402 nor n9102 n9111 ; n9594
g9403 and asqrt[25] n9594 ; n9595
g9404 nor n9109 n9595 ; n9596
g9405 nor n9593 n9596 ; n9597
g9406 nor asqrt[45] n9578 ; n9598
g9407 and n9588_not n9598 ; n9599
g9408 nor n9597 n9599 ; n9600
g9409 nor n9590 n9600 ; n9601
g9410 and asqrt[46] n9601_not ; n9602
g9411 and n9114_not n9121 ; n9603
g9412 and n9123_not n9603 ; n9604
g9413 and asqrt[25] n9604 ; n9605
g9414 nor n9114 n9123 ; n9606
g9415 and asqrt[25] n9606 ; n9607
g9416 nor n9121 n9607 ; n9608
g9417 nor n9605 n9608 ; n9609
g9418 nor asqrt[46] n9590 ; n9610
g9419 and n9600_not n9610 ; n9611
g9420 nor n9609 n9611 ; n9612
g9421 nor n9602 n9612 ; n9613
g9422 and asqrt[47] n9613_not ; n9614
g9423 and n9133 n9135_not ; n9615
g9424 and n9126_not n9615 ; n9616
g9425 and asqrt[25] n9616 ; n9617
g9426 nor n9126 n9135 ; n9618
g9427 and asqrt[25] n9618 ; n9619
g9428 nor n9133 n9619 ; n9620
g9429 nor n9617 n9620 ; n9621
g9430 nor asqrt[47] n9602 ; n9622
g9431 and n9612_not n9622 ; n9623
g9432 nor n9621 n9623 ; n9624
g9433 nor n9614 n9624 ; n9625
g9434 and asqrt[48] n9625_not ; n9626
g9435 and n9138_not n9145 ; n9627
g9436 and n9147_not n9627 ; n9628
g9437 and asqrt[25] n9628 ; n9629
g9438 nor n9138 n9147 ; n9630
g9439 and asqrt[25] n9630 ; n9631
g9440 nor n9145 n9631 ; n9632
g9441 nor n9629 n9632 ; n9633
g9442 nor asqrt[48] n9614 ; n9634
g9443 and n9624_not n9634 ; n9635
g9444 nor n9633 n9635 ; n9636
g9445 nor n9626 n9636 ; n9637
g9446 and asqrt[49] n9637_not ; n9638
g9447 and n9157 n9159_not ; n9639
g9448 and n9150_not n9639 ; n9640
g9449 and asqrt[25] n9640 ; n9641
g9450 nor n9150 n9159 ; n9642
g9451 and asqrt[25] n9642 ; n9643
g9452 nor n9157 n9643 ; n9644
g9453 nor n9641 n9644 ; n9645
g9454 nor asqrt[49] n9626 ; n9646
g9455 and n9636_not n9646 ; n9647
g9456 nor n9645 n9647 ; n9648
g9457 nor n9638 n9648 ; n9649
g9458 and asqrt[50] n9649_not ; n9650
g9459 and n9162_not n9169 ; n9651
g9460 and n9171_not n9651 ; n9652
g9461 and asqrt[25] n9652 ; n9653
g9462 nor n9162 n9171 ; n9654
g9463 and asqrt[25] n9654 ; n9655
g9464 nor n9169 n9655 ; n9656
g9465 nor n9653 n9656 ; n9657
g9466 nor asqrt[50] n9638 ; n9658
g9467 and n9648_not n9658 ; n9659
g9468 nor n9657 n9659 ; n9660
g9469 nor n9650 n9660 ; n9661
g9470 and asqrt[51] n9661_not ; n9662
g9471 and n9181 n9183_not ; n9663
g9472 and n9174_not n9663 ; n9664
g9473 and asqrt[25] n9664 ; n9665
g9474 nor n9174 n9183 ; n9666
g9475 and asqrt[25] n9666 ; n9667
g9476 nor n9181 n9667 ; n9668
g9477 nor n9665 n9668 ; n9669
g9478 nor asqrt[51] n9650 ; n9670
g9479 and n9660_not n9670 ; n9671
g9480 nor n9669 n9671 ; n9672
g9481 nor n9662 n9672 ; n9673
g9482 and asqrt[52] n9673_not ; n9674
g9483 and n9186_not n9193 ; n9675
g9484 and n9195_not n9675 ; n9676
g9485 and asqrt[25] n9676 ; n9677
g9486 nor n9186 n9195 ; n9678
g9487 and asqrt[25] n9678 ; n9679
g9488 nor n9193 n9679 ; n9680
g9489 nor n9677 n9680 ; n9681
g9490 nor asqrt[52] n9662 ; n9682
g9491 and n9672_not n9682 ; n9683
g9492 nor n9681 n9683 ; n9684
g9493 nor n9674 n9684 ; n9685
g9494 and asqrt[53] n9685_not ; n9686
g9495 and n9205 n9207_not ; n9687
g9496 and n9198_not n9687 ; n9688
g9497 and asqrt[25] n9688 ; n9689
g9498 nor n9198 n9207 ; n9690
g9499 and asqrt[25] n9690 ; n9691
g9500 nor n9205 n9691 ; n9692
g9501 nor n9689 n9692 ; n9693
g9502 nor asqrt[53] n9674 ; n9694
g9503 and n9684_not n9694 ; n9695
g9504 nor n9693 n9695 ; n9696
g9505 nor n9686 n9696 ; n9697
g9506 and asqrt[54] n9697_not ; n9698
g9507 and n9210_not n9217 ; n9699
g9508 and n9219_not n9699 ; n9700
g9509 and asqrt[25] n9700 ; n9701
g9510 nor n9210 n9219 ; n9702
g9511 and asqrt[25] n9702 ; n9703
g9512 nor n9217 n9703 ; n9704
g9513 nor n9701 n9704 ; n9705
g9514 nor asqrt[54] n9686 ; n9706
g9515 and n9696_not n9706 ; n9707
g9516 nor n9705 n9707 ; n9708
g9517 nor n9698 n9708 ; n9709
g9518 and asqrt[55] n9709_not ; n9710
g9519 and n9229 n9231_not ; n9711
g9520 and n9222_not n9711 ; n9712
g9521 and asqrt[25] n9712 ; n9713
g9522 nor n9222 n9231 ; n9714
g9523 and asqrt[25] n9714 ; n9715
g9524 nor n9229 n9715 ; n9716
g9525 nor n9713 n9716 ; n9717
g9526 nor asqrt[55] n9698 ; n9718
g9527 and n9708_not n9718 ; n9719
g9528 nor n9717 n9719 ; n9720
g9529 nor n9710 n9720 ; n9721
g9530 and asqrt[56] n9721_not ; n9722
g9531 and n9234_not n9241 ; n9723
g9532 and n9243_not n9723 ; n9724
g9533 and asqrt[25] n9724 ; n9725
g9534 nor n9234 n9243 ; n9726
g9535 and asqrt[25] n9726 ; n9727
g9536 nor n9241 n9727 ; n9728
g9537 nor n9725 n9728 ; n9729
g9538 nor asqrt[56] n9710 ; n9730
g9539 and n9720_not n9730 ; n9731
g9540 nor n9729 n9731 ; n9732
g9541 nor n9722 n9732 ; n9733
g9542 and asqrt[57] n9733_not ; n9734
g9543 and n9253 n9255_not ; n9735
g9544 and n9246_not n9735 ; n9736
g9545 and asqrt[25] n9736 ; n9737
g9546 nor n9246 n9255 ; n9738
g9547 and asqrt[25] n9738 ; n9739
g9548 nor n9253 n9739 ; n9740
g9549 nor n9737 n9740 ; n9741
g9550 nor asqrt[57] n9722 ; n9742
g9551 and n9732_not n9742 ; n9743
g9552 nor n9741 n9743 ; n9744
g9553 nor n9734 n9744 ; n9745
g9554 and asqrt[58] n9745_not ; n9746
g9555 and n9258_not n9265 ; n9747
g9556 and n9267_not n9747 ; n9748
g9557 and asqrt[25] n9748 ; n9749
g9558 nor n9258 n9267 ; n9750
g9559 and asqrt[25] n9750 ; n9751
g9560 nor n9265 n9751 ; n9752
g9561 nor n9749 n9752 ; n9753
g9562 nor asqrt[58] n9734 ; n9754
g9563 and n9744_not n9754 ; n9755
g9564 nor n9753 n9755 ; n9756
g9565 nor n9746 n9756 ; n9757
g9566 and asqrt[59] n9757_not ; n9758
g9567 and n9277 n9279_not ; n9759
g9568 and n9270_not n9759 ; n9760
g9569 and asqrt[25] n9760 ; n9761
g9570 nor n9270 n9279 ; n9762
g9571 and asqrt[25] n9762 ; n9763
g9572 nor n9277 n9763 ; n9764
g9573 nor n9761 n9764 ; n9765
g9574 nor asqrt[59] n9746 ; n9766
g9575 and n9756_not n9766 ; n9767
g9576 nor n9765 n9767 ; n9768
g9577 nor n9758 n9768 ; n9769
g9578 and asqrt[60] n9769_not ; n9770
g9579 and n9282_not n9289 ; n9771
g9580 and n9291_not n9771 ; n9772
g9581 and asqrt[25] n9772 ; n9773
g9582 nor n9282 n9291 ; n9774
g9583 and asqrt[25] n9774 ; n9775
g9584 nor n9289 n9775 ; n9776
g9585 nor n9773 n9776 ; n9777
g9586 nor asqrt[60] n9758 ; n9778
g9587 and n9768_not n9778 ; n9779
g9588 nor n9777 n9779 ; n9780
g9589 nor n9770 n9780 ; n9781
g9590 and asqrt[61] n9781_not ; n9782
g9591 and n9301 n9303_not ; n9783
g9592 and n9294_not n9783 ; n9784
g9593 and asqrt[25] n9784 ; n9785
g9594 nor n9294 n9303 ; n9786
g9595 and asqrt[25] n9786 ; n9787
g9596 nor n9301 n9787 ; n9788
g9597 nor n9785 n9788 ; n9789
g9598 nor asqrt[61] n9770 ; n9790
g9599 and n9780_not n9790 ; n9791
g9600 nor n9789 n9791 ; n9792
g9601 nor n9782 n9792 ; n9793
g9602 and asqrt[62] n9793_not ; n9794
g9603 and n9306_not n9313 ; n9795
g9604 and n9315_not n9795 ; n9796
g9605 and asqrt[25] n9796 ; n9797
g9606 nor n9306 n9315 ; n9798
g9607 and asqrt[25] n9798 ; n9799
g9608 nor n9313 n9799 ; n9800
g9609 nor n9797 n9800 ; n9801
g9610 nor asqrt[62] n9782 ; n9802
g9611 and n9792_not n9802 ; n9803
g9612 nor n9801 n9803 ; n9804
g9613 nor n9794 n9804 ; n9805
g9614 and n9325 n9327_not ; n9806
g9615 and n9318_not n9806 ; n9807
g9616 and asqrt[25] n9807 ; n9808
g9617 nor n9318 n9327 ; n9809
g9618 and asqrt[25] n9809 ; n9810
g9619 nor n9325 n9810 ; n9811
g9620 nor n9808 n9811 ; n9812
g9621 nor n9329 n9336 ; n9813
g9622 and asqrt[25] n9813 ; n9814
g9623 nor n9344 n9814 ; n9815
g9624 and n9812_not n9815 ; n9816
g9625 and n9805_not n9816 ; n9817
g9626 nor asqrt[63] n9817 ; n9818
g9627 and n9794_not n9812 ; n9819
g9628 and n9804_not n9819 ; n9820
g9629 and n9336_not asqrt[25] ; n9821
g9630 and n9329 n9821_not ; n9822
g9631 and asqrt[63] n9813_not ; n9823
g9632 and n9822_not n9823 ; n9824
g9633 nor n9332 n9353 ; n9825
g9634 and n9335_not n9825 ; n9826
g9635 and n9348_not n9826 ; n9827
g9636 and n9344_not n9827 ; n9828
g9637 and n9342_not n9828 ; n9829
g9638 nor n9824 n9829 ; n9830
g9639 and n9820_not n9830 ; n9831
g9640 nand n9818_not n9831 ; asqrt[24]
g9641 and a[48] asqrt[24] ; n9833
g9642 nor a[46] a[47] ; n9834
g9643 and a[48]_not n9834 ; n9835
g9644 nor n9833 n9835 ; n9836
g9645 and asqrt[25] n9836_not ; n9837
g9646 nor n9353 n9835 ; n9838
g9647 and n9348_not n9838 ; n9839
g9648 and n9344_not n9839 ; n9840
g9649 and n9342_not n9840 ; n9841
g9650 and n9833_not n9841 ; n9842
g9651 and a[48]_not asqrt[24] ; n9843
g9652 and a[49] n9843_not ; n9844
g9653 and n9358 asqrt[24] ; n9845
g9654 nor n9844 n9845 ; n9846
g9655 and n9842_not n9846 ; n9847
g9656 nor n9837 n9847 ; n9848
g9657 and asqrt[26] n9848_not ; n9849
g9658 nor asqrt[26] n9837 ; n9850
g9659 and n9847_not n9850 ; n9851
g9660 and asqrt[25] n9829_not ; n9852
g9661 and n9824_not n9852 ; n9853
g9662 and n9820_not n9853 ; n9854
g9663 and n9818_not n9854 ; n9855
g9664 nor n9845 n9855 ; n9856
g9665 and a[50] n9856_not ; n9857
g9666 nor a[50] n9855 ; n9858
g9667 and n9845_not n9858 ; n9859
g9668 nor n9857 n9859 ; n9860
g9669 nor n9851 n9860 ; n9861
g9670 nor n9849 n9861 ; n9862
g9671 and asqrt[27] n9862_not ; n9863
g9672 nor n9361 n9366 ; n9864
g9673 and n9370_not n9864 ; n9865
g9674 and asqrt[24] n9865 ; n9866
g9675 and asqrt[24] n9864 ; n9867
g9676 and n9370 n9867_not ; n9868
g9677 nor n9866 n9868 ; n9869
g9678 nor asqrt[27] n9849 ; n9870
g9679 and n9861_not n9870 ; n9871
g9680 nor n9869 n9871 ; n9872
g9681 nor n9863 n9872 ; n9873
g9682 and asqrt[28] n9873_not ; n9874
g9683 and n9375_not n9384 ; n9875
g9684 and n9373_not n9875 ; n9876
g9685 and asqrt[24] n9876 ; n9877
g9686 nor n9373 n9375 ; n9878
g9687 and asqrt[24] n9878 ; n9879
g9688 nor n9384 n9879 ; n9880
g9689 nor n9877 n9880 ; n9881
g9690 nor asqrt[28] n9863 ; n9882
g9691 and n9872_not n9882 ; n9883
g9692 nor n9881 n9883 ; n9884
g9693 nor n9874 n9884 ; n9885
g9694 and asqrt[29] n9885_not ; n9886
g9695 and n9387_not n9393 ; n9887
g9696 and n9395_not n9887 ; n9888
g9697 and asqrt[24] n9888 ; n9889
g9698 nor n9387 n9395 ; n9890
g9699 and asqrt[24] n9890 ; n9891
g9700 nor n9393 n9891 ; n9892
g9701 nor n9889 n9892 ; n9893
g9702 nor asqrt[29] n9874 ; n9894
g9703 and n9884_not n9894 ; n9895
g9704 nor n9893 n9895 ; n9896
g9705 nor n9886 n9896 ; n9897
g9706 and asqrt[30] n9897_not ; n9898
g9707 and n9405 n9407_not ; n9899
g9708 and n9398_not n9899 ; n9900
g9709 and asqrt[24] n9900 ; n9901
g9710 nor n9398 n9407 ; n9902
g9711 and asqrt[24] n9902 ; n9903
g9712 nor n9405 n9903 ; n9904
g9713 nor n9901 n9904 ; n9905
g9714 nor asqrt[30] n9886 ; n9906
g9715 and n9896_not n9906 ; n9907
g9716 nor n9905 n9907 ; n9908
g9717 nor n9898 n9908 ; n9909
g9718 and asqrt[31] n9909_not ; n9910
g9719 and n9410_not n9417 ; n9911
g9720 and n9419_not n9911 ; n9912
g9721 and asqrt[24] n9912 ; n9913
g9722 nor n9410 n9419 ; n9914
g9723 and asqrt[24] n9914 ; n9915
g9724 nor n9417 n9915 ; n9916
g9725 nor n9913 n9916 ; n9917
g9726 nor asqrt[31] n9898 ; n9918
g9727 and n9908_not n9918 ; n9919
g9728 nor n9917 n9919 ; n9920
g9729 nor n9910 n9920 ; n9921
g9730 and asqrt[32] n9921_not ; n9922
g9731 and n9429 n9431_not ; n9923
g9732 and n9422_not n9923 ; n9924
g9733 and asqrt[24] n9924 ; n9925
g9734 nor n9422 n9431 ; n9926
g9735 and asqrt[24] n9926 ; n9927
g9736 nor n9429 n9927 ; n9928
g9737 nor n9925 n9928 ; n9929
g9738 nor asqrt[32] n9910 ; n9930
g9739 and n9920_not n9930 ; n9931
g9740 nor n9929 n9931 ; n9932
g9741 nor n9922 n9932 ; n9933
g9742 and asqrt[33] n9933_not ; n9934
g9743 and n9434_not n9441 ; n9935
g9744 and n9443_not n9935 ; n9936
g9745 and asqrt[24] n9936 ; n9937
g9746 nor n9434 n9443 ; n9938
g9747 and asqrt[24] n9938 ; n9939
g9748 nor n9441 n9939 ; n9940
g9749 nor n9937 n9940 ; n9941
g9750 nor asqrt[33] n9922 ; n9942
g9751 and n9932_not n9942 ; n9943
g9752 nor n9941 n9943 ; n9944
g9753 nor n9934 n9944 ; n9945
g9754 and asqrt[34] n9945_not ; n9946
g9755 and n9453 n9455_not ; n9947
g9756 and n9446_not n9947 ; n9948
g9757 and asqrt[24] n9948 ; n9949
g9758 nor n9446 n9455 ; n9950
g9759 and asqrt[24] n9950 ; n9951
g9760 nor n9453 n9951 ; n9952
g9761 nor n9949 n9952 ; n9953
g9762 nor asqrt[34] n9934 ; n9954
g9763 and n9944_not n9954 ; n9955
g9764 nor n9953 n9955 ; n9956
g9765 nor n9946 n9956 ; n9957
g9766 and asqrt[35] n9957_not ; n9958
g9767 and n9458_not n9465 ; n9959
g9768 and n9467_not n9959 ; n9960
g9769 and asqrt[24] n9960 ; n9961
g9770 nor n9458 n9467 ; n9962
g9771 and asqrt[24] n9962 ; n9963
g9772 nor n9465 n9963 ; n9964
g9773 nor n9961 n9964 ; n9965
g9774 nor asqrt[35] n9946 ; n9966
g9775 and n9956_not n9966 ; n9967
g9776 nor n9965 n9967 ; n9968
g9777 nor n9958 n9968 ; n9969
g9778 and asqrt[36] n9969_not ; n9970
g9779 and n9477 n9479_not ; n9971
g9780 and n9470_not n9971 ; n9972
g9781 and asqrt[24] n9972 ; n9973
g9782 nor n9470 n9479 ; n9974
g9783 and asqrt[24] n9974 ; n9975
g9784 nor n9477 n9975 ; n9976
g9785 nor n9973 n9976 ; n9977
g9786 nor asqrt[36] n9958 ; n9978
g9787 and n9968_not n9978 ; n9979
g9788 nor n9977 n9979 ; n9980
g9789 nor n9970 n9980 ; n9981
g9790 and asqrt[37] n9981_not ; n9982
g9791 and n9482_not n9489 ; n9983
g9792 and n9491_not n9983 ; n9984
g9793 and asqrt[24] n9984 ; n9985
g9794 nor n9482 n9491 ; n9986
g9795 and asqrt[24] n9986 ; n9987
g9796 nor n9489 n9987 ; n9988
g9797 nor n9985 n9988 ; n9989
g9798 nor asqrt[37] n9970 ; n9990
g9799 and n9980_not n9990 ; n9991
g9800 nor n9989 n9991 ; n9992
g9801 nor n9982 n9992 ; n9993
g9802 and asqrt[38] n9993_not ; n9994
g9803 and n9501 n9503_not ; n9995
g9804 and n9494_not n9995 ; n9996
g9805 and asqrt[24] n9996 ; n9997
g9806 nor n9494 n9503 ; n9998
g9807 and asqrt[24] n9998 ; n9999
g9808 nor n9501 n9999 ; n10000
g9809 nor n9997 n10000 ; n10001
g9810 nor asqrt[38] n9982 ; n10002
g9811 and n9992_not n10002 ; n10003
g9812 nor n10001 n10003 ; n10004
g9813 nor n9994 n10004 ; n10005
g9814 and asqrt[39] n10005_not ; n10006
g9815 and n9506_not n9513 ; n10007
g9816 and n9515_not n10007 ; n10008
g9817 and asqrt[24] n10008 ; n10009
g9818 nor n9506 n9515 ; n10010
g9819 and asqrt[24] n10010 ; n10011
g9820 nor n9513 n10011 ; n10012
g9821 nor n10009 n10012 ; n10013
g9822 nor asqrt[39] n9994 ; n10014
g9823 and n10004_not n10014 ; n10015
g9824 nor n10013 n10015 ; n10016
g9825 nor n10006 n10016 ; n10017
g9826 and asqrt[40] n10017_not ; n10018
g9827 and n9525 n9527_not ; n10019
g9828 and n9518_not n10019 ; n10020
g9829 and asqrt[24] n10020 ; n10021
g9830 nor n9518 n9527 ; n10022
g9831 and asqrt[24] n10022 ; n10023
g9832 nor n9525 n10023 ; n10024
g9833 nor n10021 n10024 ; n10025
g9834 nor asqrt[40] n10006 ; n10026
g9835 and n10016_not n10026 ; n10027
g9836 nor n10025 n10027 ; n10028
g9837 nor n10018 n10028 ; n10029
g9838 and asqrt[41] n10029_not ; n10030
g9839 nor asqrt[41] n10018 ; n10031
g9840 and n10028_not n10031 ; n10032
g9841 and n9530_not n9539 ; n10033
g9842 and n9532_not n10033 ; n10034
g9843 and asqrt[24] n10034 ; n10035
g9844 nor n9530 n9532 ; n10036
g9845 and asqrt[24] n10036 ; n10037
g9846 nor n9539 n10037 ; n10038
g9847 nor n10035 n10038 ; n10039
g9848 nor n10032 n10039 ; n10040
g9849 nor n10030 n10040 ; n10041
g9850 and asqrt[42] n10041_not ; n10042
g9851 and n9549 n9551_not ; n10043
g9852 and n9542_not n10043 ; n10044
g9853 and asqrt[24] n10044 ; n10045
g9854 nor n9542 n9551 ; n10046
g9855 and asqrt[24] n10046 ; n10047
g9856 nor n9549 n10047 ; n10048
g9857 nor n10045 n10048 ; n10049
g9858 nor asqrt[42] n10030 ; n10050
g9859 and n10040_not n10050 ; n10051
g9860 nor n10049 n10051 ; n10052
g9861 nor n10042 n10052 ; n10053
g9862 and asqrt[43] n10053_not ; n10054
g9863 and n9554_not n9561 ; n10055
g9864 and n9563_not n10055 ; n10056
g9865 and asqrt[24] n10056 ; n10057
g9866 nor n9554 n9563 ; n10058
g9867 and asqrt[24] n10058 ; n10059
g9868 nor n9561 n10059 ; n10060
g9869 nor n10057 n10060 ; n10061
g9870 nor asqrt[43] n10042 ; n10062
g9871 and n10052_not n10062 ; n10063
g9872 nor n10061 n10063 ; n10064
g9873 nor n10054 n10064 ; n10065
g9874 and asqrt[44] n10065_not ; n10066
g9875 and n9573 n9575_not ; n10067
g9876 and n9566_not n10067 ; n10068
g9877 and asqrt[24] n10068 ; n10069
g9878 nor n9566 n9575 ; n10070
g9879 and asqrt[24] n10070 ; n10071
g9880 nor n9573 n10071 ; n10072
g9881 nor n10069 n10072 ; n10073
g9882 nor asqrt[44] n10054 ; n10074
g9883 and n10064_not n10074 ; n10075
g9884 nor n10073 n10075 ; n10076
g9885 nor n10066 n10076 ; n10077
g9886 and asqrt[45] n10077_not ; n10078
g9887 and n9578_not n9585 ; n10079
g9888 and n9587_not n10079 ; n10080
g9889 and asqrt[24] n10080 ; n10081
g9890 nor n9578 n9587 ; n10082
g9891 and asqrt[24] n10082 ; n10083
g9892 nor n9585 n10083 ; n10084
g9893 nor n10081 n10084 ; n10085
g9894 nor asqrt[45] n10066 ; n10086
g9895 and n10076_not n10086 ; n10087
g9896 nor n10085 n10087 ; n10088
g9897 nor n10078 n10088 ; n10089
g9898 and asqrt[46] n10089_not ; n10090
g9899 and n9597 n9599_not ; n10091
g9900 and n9590_not n10091 ; n10092
g9901 and asqrt[24] n10092 ; n10093
g9902 nor n9590 n9599 ; n10094
g9903 and asqrt[24] n10094 ; n10095
g9904 nor n9597 n10095 ; n10096
g9905 nor n10093 n10096 ; n10097
g9906 nor asqrt[46] n10078 ; n10098
g9907 and n10088_not n10098 ; n10099
g9908 nor n10097 n10099 ; n10100
g9909 nor n10090 n10100 ; n10101
g9910 and asqrt[47] n10101_not ; n10102
g9911 and n9602_not n9609 ; n10103
g9912 and n9611_not n10103 ; n10104
g9913 and asqrt[24] n10104 ; n10105
g9914 nor n9602 n9611 ; n10106
g9915 and asqrt[24] n10106 ; n10107
g9916 nor n9609 n10107 ; n10108
g9917 nor n10105 n10108 ; n10109
g9918 nor asqrt[47] n10090 ; n10110
g9919 and n10100_not n10110 ; n10111
g9920 nor n10109 n10111 ; n10112
g9921 nor n10102 n10112 ; n10113
g9922 and asqrt[48] n10113_not ; n10114
g9923 and n9621 n9623_not ; n10115
g9924 and n9614_not n10115 ; n10116
g9925 and asqrt[24] n10116 ; n10117
g9926 nor n9614 n9623 ; n10118
g9927 and asqrt[24] n10118 ; n10119
g9928 nor n9621 n10119 ; n10120
g9929 nor n10117 n10120 ; n10121
g9930 nor asqrt[48] n10102 ; n10122
g9931 and n10112_not n10122 ; n10123
g9932 nor n10121 n10123 ; n10124
g9933 nor n10114 n10124 ; n10125
g9934 and asqrt[49] n10125_not ; n10126
g9935 and n9626_not n9633 ; n10127
g9936 and n9635_not n10127 ; n10128
g9937 and asqrt[24] n10128 ; n10129
g9938 nor n9626 n9635 ; n10130
g9939 and asqrt[24] n10130 ; n10131
g9940 nor n9633 n10131 ; n10132
g9941 nor n10129 n10132 ; n10133
g9942 nor asqrt[49] n10114 ; n10134
g9943 and n10124_not n10134 ; n10135
g9944 nor n10133 n10135 ; n10136
g9945 nor n10126 n10136 ; n10137
g9946 and asqrt[50] n10137_not ; n10138
g9947 and n9645 n9647_not ; n10139
g9948 and n9638_not n10139 ; n10140
g9949 and asqrt[24] n10140 ; n10141
g9950 nor n9638 n9647 ; n10142
g9951 and asqrt[24] n10142 ; n10143
g9952 nor n9645 n10143 ; n10144
g9953 nor n10141 n10144 ; n10145
g9954 nor asqrt[50] n10126 ; n10146
g9955 and n10136_not n10146 ; n10147
g9956 nor n10145 n10147 ; n10148
g9957 nor n10138 n10148 ; n10149
g9958 and asqrt[51] n10149_not ; n10150
g9959 and n9650_not n9657 ; n10151
g9960 and n9659_not n10151 ; n10152
g9961 and asqrt[24] n10152 ; n10153
g9962 nor n9650 n9659 ; n10154
g9963 and asqrt[24] n10154 ; n10155
g9964 nor n9657 n10155 ; n10156
g9965 nor n10153 n10156 ; n10157
g9966 nor asqrt[51] n10138 ; n10158
g9967 and n10148_not n10158 ; n10159
g9968 nor n10157 n10159 ; n10160
g9969 nor n10150 n10160 ; n10161
g9970 and asqrt[52] n10161_not ; n10162
g9971 and n9669 n9671_not ; n10163
g9972 and n9662_not n10163 ; n10164
g9973 and asqrt[24] n10164 ; n10165
g9974 nor n9662 n9671 ; n10166
g9975 and asqrt[24] n10166 ; n10167
g9976 nor n9669 n10167 ; n10168
g9977 nor n10165 n10168 ; n10169
g9978 nor asqrt[52] n10150 ; n10170
g9979 and n10160_not n10170 ; n10171
g9980 nor n10169 n10171 ; n10172
g9981 nor n10162 n10172 ; n10173
g9982 and asqrt[53] n10173_not ; n10174
g9983 and n9674_not n9681 ; n10175
g9984 and n9683_not n10175 ; n10176
g9985 and asqrt[24] n10176 ; n10177
g9986 nor n9674 n9683 ; n10178
g9987 and asqrt[24] n10178 ; n10179
g9988 nor n9681 n10179 ; n10180
g9989 nor n10177 n10180 ; n10181
g9990 nor asqrt[53] n10162 ; n10182
g9991 and n10172_not n10182 ; n10183
g9992 nor n10181 n10183 ; n10184
g9993 nor n10174 n10184 ; n10185
g9994 and asqrt[54] n10185_not ; n10186
g9995 and n9693 n9695_not ; n10187
g9996 and n9686_not n10187 ; n10188
g9997 and asqrt[24] n10188 ; n10189
g9998 nor n9686 n9695 ; n10190
g9999 and asqrt[24] n10190 ; n10191
g10000 nor n9693 n10191 ; n10192
g10001 nor n10189 n10192 ; n10193
g10002 nor asqrt[54] n10174 ; n10194
g10003 and n10184_not n10194 ; n10195
g10004 nor n10193 n10195 ; n10196
g10005 nor n10186 n10196 ; n10197
g10006 and asqrt[55] n10197_not ; n10198
g10007 and n9698_not n9705 ; n10199
g10008 and n9707_not n10199 ; n10200
g10009 and asqrt[24] n10200 ; n10201
g10010 nor n9698 n9707 ; n10202
g10011 and asqrt[24] n10202 ; n10203
g10012 nor n9705 n10203 ; n10204
g10013 nor n10201 n10204 ; n10205
g10014 nor asqrt[55] n10186 ; n10206
g10015 and n10196_not n10206 ; n10207
g10016 nor n10205 n10207 ; n10208
g10017 nor n10198 n10208 ; n10209
g10018 and asqrt[56] n10209_not ; n10210
g10019 and n9717 n9719_not ; n10211
g10020 and n9710_not n10211 ; n10212
g10021 and asqrt[24] n10212 ; n10213
g10022 nor n9710 n9719 ; n10214
g10023 and asqrt[24] n10214 ; n10215
g10024 nor n9717 n10215 ; n10216
g10025 nor n10213 n10216 ; n10217
g10026 nor asqrt[56] n10198 ; n10218
g10027 and n10208_not n10218 ; n10219
g10028 nor n10217 n10219 ; n10220
g10029 nor n10210 n10220 ; n10221
g10030 and asqrt[57] n10221_not ; n10222
g10031 and n9722_not n9729 ; n10223
g10032 and n9731_not n10223 ; n10224
g10033 and asqrt[24] n10224 ; n10225
g10034 nor n9722 n9731 ; n10226
g10035 and asqrt[24] n10226 ; n10227
g10036 nor n9729 n10227 ; n10228
g10037 nor n10225 n10228 ; n10229
g10038 nor asqrt[57] n10210 ; n10230
g10039 and n10220_not n10230 ; n10231
g10040 nor n10229 n10231 ; n10232
g10041 nor n10222 n10232 ; n10233
g10042 and asqrt[58] n10233_not ; n10234
g10043 and n9741 n9743_not ; n10235
g10044 and n9734_not n10235 ; n10236
g10045 and asqrt[24] n10236 ; n10237
g10046 nor n9734 n9743 ; n10238
g10047 and asqrt[24] n10238 ; n10239
g10048 nor n9741 n10239 ; n10240
g10049 nor n10237 n10240 ; n10241
g10050 nor asqrt[58] n10222 ; n10242
g10051 and n10232_not n10242 ; n10243
g10052 nor n10241 n10243 ; n10244
g10053 nor n10234 n10244 ; n10245
g10054 and asqrt[59] n10245_not ; n10246
g10055 and n9746_not n9753 ; n10247
g10056 and n9755_not n10247 ; n10248
g10057 and asqrt[24] n10248 ; n10249
g10058 nor n9746 n9755 ; n10250
g10059 and asqrt[24] n10250 ; n10251
g10060 nor n9753 n10251 ; n10252
g10061 nor n10249 n10252 ; n10253
g10062 nor asqrt[59] n10234 ; n10254
g10063 and n10244_not n10254 ; n10255
g10064 nor n10253 n10255 ; n10256
g10065 nor n10246 n10256 ; n10257
g10066 and asqrt[60] n10257_not ; n10258
g10067 and n9765 n9767_not ; n10259
g10068 and n9758_not n10259 ; n10260
g10069 and asqrt[24] n10260 ; n10261
g10070 nor n9758 n9767 ; n10262
g10071 and asqrt[24] n10262 ; n10263
g10072 nor n9765 n10263 ; n10264
g10073 nor n10261 n10264 ; n10265
g10074 nor asqrt[60] n10246 ; n10266
g10075 and n10256_not n10266 ; n10267
g10076 nor n10265 n10267 ; n10268
g10077 nor n10258 n10268 ; n10269
g10078 and asqrt[61] n10269_not ; n10270
g10079 and n9770_not n9777 ; n10271
g10080 and n9779_not n10271 ; n10272
g10081 and asqrt[24] n10272 ; n10273
g10082 nor n9770 n9779 ; n10274
g10083 and asqrt[24] n10274 ; n10275
g10084 nor n9777 n10275 ; n10276
g10085 nor n10273 n10276 ; n10277
g10086 nor asqrt[61] n10258 ; n10278
g10087 and n10268_not n10278 ; n10279
g10088 nor n10277 n10279 ; n10280
g10089 nor n10270 n10280 ; n10281
g10090 and asqrt[62] n10281_not ; n10282
g10091 and n9789 n9791_not ; n10283
g10092 and n9782_not n10283 ; n10284
g10093 and asqrt[24] n10284 ; n10285
g10094 nor n9782 n9791 ; n10286
g10095 and asqrt[24] n10286 ; n10287
g10096 nor n9789 n10287 ; n10288
g10097 nor n10285 n10288 ; n10289
g10098 nor asqrt[62] n10270 ; n10290
g10099 and n10280_not n10290 ; n10291
g10100 nor n10289 n10291 ; n10292
g10101 nor n10282 n10292 ; n10293
g10102 and n9794_not n9801 ; n10294
g10103 and n9803_not n10294 ; n10295
g10104 and asqrt[24] n10295 ; n10296
g10105 nor n9794 n9803 ; n10297
g10106 and asqrt[24] n10297 ; n10298
g10107 nor n9801 n10298 ; n10299
g10108 nor n10296 n10299 ; n10300
g10109 nor n9805 n9812 ; n10301
g10110 and asqrt[24] n10301 ; n10302
g10111 nor n9820 n10302 ; n10303
g10112 and n10300_not n10303 ; n10304
g10113 and n10293_not n10304 ; n10305
g10114 nor asqrt[63] n10305 ; n10306
g10115 and n10282_not n10300 ; n10307
g10116 and n10292_not n10307 ; n10308
g10117 and n9812_not asqrt[24] ; n10309
g10118 and n9805 n10309_not ; n10310
g10119 and asqrt[63] n10301_not ; n10311
g10120 and n10310_not n10311 ; n10312
g10121 nor n9808 n9829 ; n10313
g10122 and n9811_not n10313 ; n10314
g10123 and n9824_not n10314 ; n10315
g10124 and n9820_not n10315 ; n10316
g10125 and n9818_not n10316 ; n10317
g10126 nor n10312 n10317 ; n10318
g10127 and n10308_not n10318 ; n10319
g10128 nand n10306_not n10319 ; asqrt[23]
g10129 and a[46] asqrt[23] ; n10321
g10130 nor a[44] a[45] ; n10322
g10131 and a[46]_not n10322 ; n10323
g10132 nor n10321 n10323 ; n10324
g10133 and asqrt[24] n10324_not ; n10325
g10134 nor n9829 n10323 ; n10326
g10135 and n9824_not n10326 ; n10327
g10136 and n9820_not n10327 ; n10328
g10137 and n9818_not n10328 ; n10329
g10138 and n10321_not n10329 ; n10330
g10139 and a[46]_not asqrt[23] ; n10331
g10140 and a[47] n10331_not ; n10332
g10141 and n9834 asqrt[23] ; n10333
g10142 nor n10332 n10333 ; n10334
g10143 and n10330_not n10334 ; n10335
g10144 nor n10325 n10335 ; n10336
g10145 and asqrt[25] n10336_not ; n10337
g10146 nor asqrt[25] n10325 ; n10338
g10147 and n10335_not n10338 ; n10339
g10148 and asqrt[24] n10317_not ; n10340
g10149 and n10312_not n10340 ; n10341
g10150 and n10308_not n10341 ; n10342
g10151 and n10306_not n10342 ; n10343
g10152 nor n10333 n10343 ; n10344
g10153 and a[48] n10344_not ; n10345
g10154 nor a[48] n10343 ; n10346
g10155 and n10333_not n10346 ; n10347
g10156 nor n10345 n10347 ; n10348
g10157 nor n10339 n10348 ; n10349
g10158 nor n10337 n10349 ; n10350
g10159 and asqrt[26] n10350_not ; n10351
g10160 nor n9837 n9842 ; n10352
g10161 and n9846_not n10352 ; n10353
g10162 and asqrt[23] n10353 ; n10354
g10163 and asqrt[23] n10352 ; n10355
g10164 and n9846 n10355_not ; n10356
g10165 nor n10354 n10356 ; n10357
g10166 nor asqrt[26] n10337 ; n10358
g10167 and n10349_not n10358 ; n10359
g10168 nor n10357 n10359 ; n10360
g10169 nor n10351 n10360 ; n10361
g10170 and asqrt[27] n10361_not ; n10362
g10171 and n9851_not n9860 ; n10363
g10172 and n9849_not n10363 ; n10364
g10173 and asqrt[23] n10364 ; n10365
g10174 nor n9849 n9851 ; n10366
g10175 and asqrt[23] n10366 ; n10367
g10176 nor n9860 n10367 ; n10368
g10177 nor n10365 n10368 ; n10369
g10178 nor asqrt[27] n10351 ; n10370
g10179 and n10360_not n10370 ; n10371
g10180 nor n10369 n10371 ; n10372
g10181 nor n10362 n10372 ; n10373
g10182 and asqrt[28] n10373_not ; n10374
g10183 and n9863_not n9869 ; n10375
g10184 and n9871_not n10375 ; n10376
g10185 and asqrt[23] n10376 ; n10377
g10186 nor n9863 n9871 ; n10378
g10187 and asqrt[23] n10378 ; n10379
g10188 nor n9869 n10379 ; n10380
g10189 nor n10377 n10380 ; n10381
g10190 nor asqrt[28] n10362 ; n10382
g10191 and n10372_not n10382 ; n10383
g10192 nor n10381 n10383 ; n10384
g10193 nor n10374 n10384 ; n10385
g10194 and asqrt[29] n10385_not ; n10386
g10195 and n9881 n9883_not ; n10387
g10196 and n9874_not n10387 ; n10388
g10197 and asqrt[23] n10388 ; n10389
g10198 nor n9874 n9883 ; n10390
g10199 and asqrt[23] n10390 ; n10391
g10200 nor n9881 n10391 ; n10392
g10201 nor n10389 n10392 ; n10393
g10202 nor asqrt[29] n10374 ; n10394
g10203 and n10384_not n10394 ; n10395
g10204 nor n10393 n10395 ; n10396
g10205 nor n10386 n10396 ; n10397
g10206 and asqrt[30] n10397_not ; n10398
g10207 and n9886_not n9893 ; n10399
g10208 and n9895_not n10399 ; n10400
g10209 and asqrt[23] n10400 ; n10401
g10210 nor n9886 n9895 ; n10402
g10211 and asqrt[23] n10402 ; n10403
g10212 nor n9893 n10403 ; n10404
g10213 nor n10401 n10404 ; n10405
g10214 nor asqrt[30] n10386 ; n10406
g10215 and n10396_not n10406 ; n10407
g10216 nor n10405 n10407 ; n10408
g10217 nor n10398 n10408 ; n10409
g10218 and asqrt[31] n10409_not ; n10410
g10219 and n9905 n9907_not ; n10411
g10220 and n9898_not n10411 ; n10412
g10221 and asqrt[23] n10412 ; n10413
g10222 nor n9898 n9907 ; n10414
g10223 and asqrt[23] n10414 ; n10415
g10224 nor n9905 n10415 ; n10416
g10225 nor n10413 n10416 ; n10417
g10226 nor asqrt[31] n10398 ; n10418
g10227 and n10408_not n10418 ; n10419
g10228 nor n10417 n10419 ; n10420
g10229 nor n10410 n10420 ; n10421
g10230 and asqrt[32] n10421_not ; n10422
g10231 and n9910_not n9917 ; n10423
g10232 and n9919_not n10423 ; n10424
g10233 and asqrt[23] n10424 ; n10425
g10234 nor n9910 n9919 ; n10426
g10235 and asqrt[23] n10426 ; n10427
g10236 nor n9917 n10427 ; n10428
g10237 nor n10425 n10428 ; n10429
g10238 nor asqrt[32] n10410 ; n10430
g10239 and n10420_not n10430 ; n10431
g10240 nor n10429 n10431 ; n10432
g10241 nor n10422 n10432 ; n10433
g10242 and asqrt[33] n10433_not ; n10434
g10243 and n9929 n9931_not ; n10435
g10244 and n9922_not n10435 ; n10436
g10245 and asqrt[23] n10436 ; n10437
g10246 nor n9922 n9931 ; n10438
g10247 and asqrt[23] n10438 ; n10439
g10248 nor n9929 n10439 ; n10440
g10249 nor n10437 n10440 ; n10441
g10250 nor asqrt[33] n10422 ; n10442
g10251 and n10432_not n10442 ; n10443
g10252 nor n10441 n10443 ; n10444
g10253 nor n10434 n10444 ; n10445
g10254 and asqrt[34] n10445_not ; n10446
g10255 and n9934_not n9941 ; n10447
g10256 and n9943_not n10447 ; n10448
g10257 and asqrt[23] n10448 ; n10449
g10258 nor n9934 n9943 ; n10450
g10259 and asqrt[23] n10450 ; n10451
g10260 nor n9941 n10451 ; n10452
g10261 nor n10449 n10452 ; n10453
g10262 nor asqrt[34] n10434 ; n10454
g10263 and n10444_not n10454 ; n10455
g10264 nor n10453 n10455 ; n10456
g10265 nor n10446 n10456 ; n10457
g10266 and asqrt[35] n10457_not ; n10458
g10267 and n9953 n9955_not ; n10459
g10268 and n9946_not n10459 ; n10460
g10269 and asqrt[23] n10460 ; n10461
g10270 nor n9946 n9955 ; n10462
g10271 and asqrt[23] n10462 ; n10463
g10272 nor n9953 n10463 ; n10464
g10273 nor n10461 n10464 ; n10465
g10274 nor asqrt[35] n10446 ; n10466
g10275 and n10456_not n10466 ; n10467
g10276 nor n10465 n10467 ; n10468
g10277 nor n10458 n10468 ; n10469
g10278 and asqrt[36] n10469_not ; n10470
g10279 and n9958_not n9965 ; n10471
g10280 and n9967_not n10471 ; n10472
g10281 and asqrt[23] n10472 ; n10473
g10282 nor n9958 n9967 ; n10474
g10283 and asqrt[23] n10474 ; n10475
g10284 nor n9965 n10475 ; n10476
g10285 nor n10473 n10476 ; n10477
g10286 nor asqrt[36] n10458 ; n10478
g10287 and n10468_not n10478 ; n10479
g10288 nor n10477 n10479 ; n10480
g10289 nor n10470 n10480 ; n10481
g10290 and asqrt[37] n10481_not ; n10482
g10291 and n9977 n9979_not ; n10483
g10292 and n9970_not n10483 ; n10484
g10293 and asqrt[23] n10484 ; n10485
g10294 nor n9970 n9979 ; n10486
g10295 and asqrt[23] n10486 ; n10487
g10296 nor n9977 n10487 ; n10488
g10297 nor n10485 n10488 ; n10489
g10298 nor asqrt[37] n10470 ; n10490
g10299 and n10480_not n10490 ; n10491
g10300 nor n10489 n10491 ; n10492
g10301 nor n10482 n10492 ; n10493
g10302 and asqrt[38] n10493_not ; n10494
g10303 and n9982_not n9989 ; n10495
g10304 and n9991_not n10495 ; n10496
g10305 and asqrt[23] n10496 ; n10497
g10306 nor n9982 n9991 ; n10498
g10307 and asqrt[23] n10498 ; n10499
g10308 nor n9989 n10499 ; n10500
g10309 nor n10497 n10500 ; n10501
g10310 nor asqrt[38] n10482 ; n10502
g10311 and n10492_not n10502 ; n10503
g10312 nor n10501 n10503 ; n10504
g10313 nor n10494 n10504 ; n10505
g10314 and asqrt[39] n10505_not ; n10506
g10315 and n10001 n10003_not ; n10507
g10316 and n9994_not n10507 ; n10508
g10317 and asqrt[23] n10508 ; n10509
g10318 nor n9994 n10003 ; n10510
g10319 and asqrt[23] n10510 ; n10511
g10320 nor n10001 n10511 ; n10512
g10321 nor n10509 n10512 ; n10513
g10322 nor asqrt[39] n10494 ; n10514
g10323 and n10504_not n10514 ; n10515
g10324 nor n10513 n10515 ; n10516
g10325 nor n10506 n10516 ; n10517
g10326 and asqrt[40] n10517_not ; n10518
g10327 and n10006_not n10013 ; n10519
g10328 and n10015_not n10519 ; n10520
g10329 and asqrt[23] n10520 ; n10521
g10330 nor n10006 n10015 ; n10522
g10331 and asqrt[23] n10522 ; n10523
g10332 nor n10013 n10523 ; n10524
g10333 nor n10521 n10524 ; n10525
g10334 nor asqrt[40] n10506 ; n10526
g10335 and n10516_not n10526 ; n10527
g10336 nor n10525 n10527 ; n10528
g10337 nor n10518 n10528 ; n10529
g10338 and asqrt[41] n10529_not ; n10530
g10339 and n10025 n10027_not ; n10531
g10340 and n10018_not n10531 ; n10532
g10341 and asqrt[23] n10532 ; n10533
g10342 nor n10018 n10027 ; n10534
g10343 and asqrt[23] n10534 ; n10535
g10344 nor n10025 n10535 ; n10536
g10345 nor n10533 n10536 ; n10537
g10346 nor asqrt[41] n10518 ; n10538
g10347 and n10528_not n10538 ; n10539
g10348 nor n10537 n10539 ; n10540
g10349 nor n10530 n10540 ; n10541
g10350 and asqrt[42] n10541_not ; n10542
g10351 nor asqrt[42] n10530 ; n10543
g10352 and n10540_not n10543 ; n10544
g10353 and n10030_not n10039 ; n10545
g10354 and n10032_not n10545 ; n10546
g10355 and asqrt[23] n10546 ; n10547
g10356 nor n10030 n10032 ; n10548
g10357 and asqrt[23] n10548 ; n10549
g10358 nor n10039 n10549 ; n10550
g10359 nor n10547 n10550 ; n10551
g10360 nor n10544 n10551 ; n10552
g10361 nor n10542 n10552 ; n10553
g10362 and asqrt[43] n10553_not ; n10554
g10363 and n10049 n10051_not ; n10555
g10364 and n10042_not n10555 ; n10556
g10365 and asqrt[23] n10556 ; n10557
g10366 nor n10042 n10051 ; n10558
g10367 and asqrt[23] n10558 ; n10559
g10368 nor n10049 n10559 ; n10560
g10369 nor n10557 n10560 ; n10561
g10370 nor asqrt[43] n10542 ; n10562
g10371 and n10552_not n10562 ; n10563
g10372 nor n10561 n10563 ; n10564
g10373 nor n10554 n10564 ; n10565
g10374 and asqrt[44] n10565_not ; n10566
g10375 and n10054_not n10061 ; n10567
g10376 and n10063_not n10567 ; n10568
g10377 and asqrt[23] n10568 ; n10569
g10378 nor n10054 n10063 ; n10570
g10379 and asqrt[23] n10570 ; n10571
g10380 nor n10061 n10571 ; n10572
g10381 nor n10569 n10572 ; n10573
g10382 nor asqrt[44] n10554 ; n10574
g10383 and n10564_not n10574 ; n10575
g10384 nor n10573 n10575 ; n10576
g10385 nor n10566 n10576 ; n10577
g10386 and asqrt[45] n10577_not ; n10578
g10387 and n10073 n10075_not ; n10579
g10388 and n10066_not n10579 ; n10580
g10389 and asqrt[23] n10580 ; n10581
g10390 nor n10066 n10075 ; n10582
g10391 and asqrt[23] n10582 ; n10583
g10392 nor n10073 n10583 ; n10584
g10393 nor n10581 n10584 ; n10585
g10394 nor asqrt[45] n10566 ; n10586
g10395 and n10576_not n10586 ; n10587
g10396 nor n10585 n10587 ; n10588
g10397 nor n10578 n10588 ; n10589
g10398 and asqrt[46] n10589_not ; n10590
g10399 and n10078_not n10085 ; n10591
g10400 and n10087_not n10591 ; n10592
g10401 and asqrt[23] n10592 ; n10593
g10402 nor n10078 n10087 ; n10594
g10403 and asqrt[23] n10594 ; n10595
g10404 nor n10085 n10595 ; n10596
g10405 nor n10593 n10596 ; n10597
g10406 nor asqrt[46] n10578 ; n10598
g10407 and n10588_not n10598 ; n10599
g10408 nor n10597 n10599 ; n10600
g10409 nor n10590 n10600 ; n10601
g10410 and asqrt[47] n10601_not ; n10602
g10411 and n10097 n10099_not ; n10603
g10412 and n10090_not n10603 ; n10604
g10413 and asqrt[23] n10604 ; n10605
g10414 nor n10090 n10099 ; n10606
g10415 and asqrt[23] n10606 ; n10607
g10416 nor n10097 n10607 ; n10608
g10417 nor n10605 n10608 ; n10609
g10418 nor asqrt[47] n10590 ; n10610
g10419 and n10600_not n10610 ; n10611
g10420 nor n10609 n10611 ; n10612
g10421 nor n10602 n10612 ; n10613
g10422 and asqrt[48] n10613_not ; n10614
g10423 and n10102_not n10109 ; n10615
g10424 and n10111_not n10615 ; n10616
g10425 and asqrt[23] n10616 ; n10617
g10426 nor n10102 n10111 ; n10618
g10427 and asqrt[23] n10618 ; n10619
g10428 nor n10109 n10619 ; n10620
g10429 nor n10617 n10620 ; n10621
g10430 nor asqrt[48] n10602 ; n10622
g10431 and n10612_not n10622 ; n10623
g10432 nor n10621 n10623 ; n10624
g10433 nor n10614 n10624 ; n10625
g10434 and asqrt[49] n10625_not ; n10626
g10435 and n10121 n10123_not ; n10627
g10436 and n10114_not n10627 ; n10628
g10437 and asqrt[23] n10628 ; n10629
g10438 nor n10114 n10123 ; n10630
g10439 and asqrt[23] n10630 ; n10631
g10440 nor n10121 n10631 ; n10632
g10441 nor n10629 n10632 ; n10633
g10442 nor asqrt[49] n10614 ; n10634
g10443 and n10624_not n10634 ; n10635
g10444 nor n10633 n10635 ; n10636
g10445 nor n10626 n10636 ; n10637
g10446 and asqrt[50] n10637_not ; n10638
g10447 and n10126_not n10133 ; n10639
g10448 and n10135_not n10639 ; n10640
g10449 and asqrt[23] n10640 ; n10641
g10450 nor n10126 n10135 ; n10642
g10451 and asqrt[23] n10642 ; n10643
g10452 nor n10133 n10643 ; n10644
g10453 nor n10641 n10644 ; n10645
g10454 nor asqrt[50] n10626 ; n10646
g10455 and n10636_not n10646 ; n10647
g10456 nor n10645 n10647 ; n10648
g10457 nor n10638 n10648 ; n10649
g10458 and asqrt[51] n10649_not ; n10650
g10459 and n10145 n10147_not ; n10651
g10460 and n10138_not n10651 ; n10652
g10461 and asqrt[23] n10652 ; n10653
g10462 nor n10138 n10147 ; n10654
g10463 and asqrt[23] n10654 ; n10655
g10464 nor n10145 n10655 ; n10656
g10465 nor n10653 n10656 ; n10657
g10466 nor asqrt[51] n10638 ; n10658
g10467 and n10648_not n10658 ; n10659
g10468 nor n10657 n10659 ; n10660
g10469 nor n10650 n10660 ; n10661
g10470 and asqrt[52] n10661_not ; n10662
g10471 and n10150_not n10157 ; n10663
g10472 and n10159_not n10663 ; n10664
g10473 and asqrt[23] n10664 ; n10665
g10474 nor n10150 n10159 ; n10666
g10475 and asqrt[23] n10666 ; n10667
g10476 nor n10157 n10667 ; n10668
g10477 nor n10665 n10668 ; n10669
g10478 nor asqrt[52] n10650 ; n10670
g10479 and n10660_not n10670 ; n10671
g10480 nor n10669 n10671 ; n10672
g10481 nor n10662 n10672 ; n10673
g10482 and asqrt[53] n10673_not ; n10674
g10483 and n10169 n10171_not ; n10675
g10484 and n10162_not n10675 ; n10676
g10485 and asqrt[23] n10676 ; n10677
g10486 nor n10162 n10171 ; n10678
g10487 and asqrt[23] n10678 ; n10679
g10488 nor n10169 n10679 ; n10680
g10489 nor n10677 n10680 ; n10681
g10490 nor asqrt[53] n10662 ; n10682
g10491 and n10672_not n10682 ; n10683
g10492 nor n10681 n10683 ; n10684
g10493 nor n10674 n10684 ; n10685
g10494 and asqrt[54] n10685_not ; n10686
g10495 and n10174_not n10181 ; n10687
g10496 and n10183_not n10687 ; n10688
g10497 and asqrt[23] n10688 ; n10689
g10498 nor n10174 n10183 ; n10690
g10499 and asqrt[23] n10690 ; n10691
g10500 nor n10181 n10691 ; n10692
g10501 nor n10689 n10692 ; n10693
g10502 nor asqrt[54] n10674 ; n10694
g10503 and n10684_not n10694 ; n10695
g10504 nor n10693 n10695 ; n10696
g10505 nor n10686 n10696 ; n10697
g10506 and asqrt[55] n10697_not ; n10698
g10507 and n10193 n10195_not ; n10699
g10508 and n10186_not n10699 ; n10700
g10509 and asqrt[23] n10700 ; n10701
g10510 nor n10186 n10195 ; n10702
g10511 and asqrt[23] n10702 ; n10703
g10512 nor n10193 n10703 ; n10704
g10513 nor n10701 n10704 ; n10705
g10514 nor asqrt[55] n10686 ; n10706
g10515 and n10696_not n10706 ; n10707
g10516 nor n10705 n10707 ; n10708
g10517 nor n10698 n10708 ; n10709
g10518 and asqrt[56] n10709_not ; n10710
g10519 and n10198_not n10205 ; n10711
g10520 and n10207_not n10711 ; n10712
g10521 and asqrt[23] n10712 ; n10713
g10522 nor n10198 n10207 ; n10714
g10523 and asqrt[23] n10714 ; n10715
g10524 nor n10205 n10715 ; n10716
g10525 nor n10713 n10716 ; n10717
g10526 nor asqrt[56] n10698 ; n10718
g10527 and n10708_not n10718 ; n10719
g10528 nor n10717 n10719 ; n10720
g10529 nor n10710 n10720 ; n10721
g10530 and asqrt[57] n10721_not ; n10722
g10531 and n10217 n10219_not ; n10723
g10532 and n10210_not n10723 ; n10724
g10533 and asqrt[23] n10724 ; n10725
g10534 nor n10210 n10219 ; n10726
g10535 and asqrt[23] n10726 ; n10727
g10536 nor n10217 n10727 ; n10728
g10537 nor n10725 n10728 ; n10729
g10538 nor asqrt[57] n10710 ; n10730
g10539 and n10720_not n10730 ; n10731
g10540 nor n10729 n10731 ; n10732
g10541 nor n10722 n10732 ; n10733
g10542 and asqrt[58] n10733_not ; n10734
g10543 and n10222_not n10229 ; n10735
g10544 and n10231_not n10735 ; n10736
g10545 and asqrt[23] n10736 ; n10737
g10546 nor n10222 n10231 ; n10738
g10547 and asqrt[23] n10738 ; n10739
g10548 nor n10229 n10739 ; n10740
g10549 nor n10737 n10740 ; n10741
g10550 nor asqrt[58] n10722 ; n10742
g10551 and n10732_not n10742 ; n10743
g10552 nor n10741 n10743 ; n10744
g10553 nor n10734 n10744 ; n10745
g10554 and asqrt[59] n10745_not ; n10746
g10555 and n10241 n10243_not ; n10747
g10556 and n10234_not n10747 ; n10748
g10557 and asqrt[23] n10748 ; n10749
g10558 nor n10234 n10243 ; n10750
g10559 and asqrt[23] n10750 ; n10751
g10560 nor n10241 n10751 ; n10752
g10561 nor n10749 n10752 ; n10753
g10562 nor asqrt[59] n10734 ; n10754
g10563 and n10744_not n10754 ; n10755
g10564 nor n10753 n10755 ; n10756
g10565 nor n10746 n10756 ; n10757
g10566 and asqrt[60] n10757_not ; n10758
g10567 and n10246_not n10253 ; n10759
g10568 and n10255_not n10759 ; n10760
g10569 and asqrt[23] n10760 ; n10761
g10570 nor n10246 n10255 ; n10762
g10571 and asqrt[23] n10762 ; n10763
g10572 nor n10253 n10763 ; n10764
g10573 nor n10761 n10764 ; n10765
g10574 nor asqrt[60] n10746 ; n10766
g10575 and n10756_not n10766 ; n10767
g10576 nor n10765 n10767 ; n10768
g10577 nor n10758 n10768 ; n10769
g10578 and asqrt[61] n10769_not ; n10770
g10579 and n10265 n10267_not ; n10771
g10580 and n10258_not n10771 ; n10772
g10581 and asqrt[23] n10772 ; n10773
g10582 nor n10258 n10267 ; n10774
g10583 and asqrt[23] n10774 ; n10775
g10584 nor n10265 n10775 ; n10776
g10585 nor n10773 n10776 ; n10777
g10586 nor asqrt[61] n10758 ; n10778
g10587 and n10768_not n10778 ; n10779
g10588 nor n10777 n10779 ; n10780
g10589 nor n10770 n10780 ; n10781
g10590 and asqrt[62] n10781_not ; n10782
g10591 and n10270_not n10277 ; n10783
g10592 and n10279_not n10783 ; n10784
g10593 and asqrt[23] n10784 ; n10785
g10594 nor n10270 n10279 ; n10786
g10595 and asqrt[23] n10786 ; n10787
g10596 nor n10277 n10787 ; n10788
g10597 nor n10785 n10788 ; n10789
g10598 nor asqrt[62] n10770 ; n10790
g10599 and n10780_not n10790 ; n10791
g10600 nor n10789 n10791 ; n10792
g10601 nor n10782 n10792 ; n10793
g10602 and n10289 n10291_not ; n10794
g10603 and n10282_not n10794 ; n10795
g10604 and asqrt[23] n10795 ; n10796
g10605 nor n10282 n10291 ; n10797
g10606 and asqrt[23] n10797 ; n10798
g10607 nor n10289 n10798 ; n10799
g10608 nor n10796 n10799 ; n10800
g10609 nor n10293 n10300 ; n10801
g10610 and asqrt[23] n10801 ; n10802
g10611 nor n10308 n10802 ; n10803
g10612 and n10800_not n10803 ; n10804
g10613 and n10793_not n10804 ; n10805
g10614 nor asqrt[63] n10805 ; n10806
g10615 and n10782_not n10800 ; n10807
g10616 and n10792_not n10807 ; n10808
g10617 and n10300_not asqrt[23] ; n10809
g10618 and n10293 n10809_not ; n10810
g10619 and asqrt[63] n10801_not ; n10811
g10620 and n10810_not n10811 ; n10812
g10621 nor n10296 n10317 ; n10813
g10622 and n10299_not n10813 ; n10814
g10623 and n10312_not n10814 ; n10815
g10624 and n10308_not n10815 ; n10816
g10625 and n10306_not n10816 ; n10817
g10626 nor n10812 n10817 ; n10818
g10627 and n10808_not n10818 ; n10819
g10628 nand n10806_not n10819 ; asqrt[22]
g10629 and a[44] asqrt[22] ; n10821
g10630 nor a[42] a[43] ; n10822
g10631 and a[44]_not n10822 ; n10823
g10632 nor n10821 n10823 ; n10824
g10633 and asqrt[23] n10824_not ; n10825
g10634 nor n10317 n10823 ; n10826
g10635 and n10312_not n10826 ; n10827
g10636 and n10308_not n10827 ; n10828
g10637 and n10306_not n10828 ; n10829
g10638 and n10821_not n10829 ; n10830
g10639 and a[44]_not asqrt[22] ; n10831
g10640 and a[45] n10831_not ; n10832
g10641 and n10322 asqrt[22] ; n10833
g10642 nor n10832 n10833 ; n10834
g10643 and n10830_not n10834 ; n10835
g10644 nor n10825 n10835 ; n10836
g10645 and asqrt[24] n10836_not ; n10837
g10646 nor asqrt[24] n10825 ; n10838
g10647 and n10835_not n10838 ; n10839
g10648 and asqrt[23] n10817_not ; n10840
g10649 and n10812_not n10840 ; n10841
g10650 and n10808_not n10841 ; n10842
g10651 and n10806_not n10842 ; n10843
g10652 nor n10833 n10843 ; n10844
g10653 and a[46] n10844_not ; n10845
g10654 nor a[46] n10843 ; n10846
g10655 and n10833_not n10846 ; n10847
g10656 nor n10845 n10847 ; n10848
g10657 nor n10839 n10848 ; n10849
g10658 nor n10837 n10849 ; n10850
g10659 and asqrt[25] n10850_not ; n10851
g10660 nor n10325 n10330 ; n10852
g10661 and n10334_not n10852 ; n10853
g10662 and asqrt[22] n10853 ; n10854
g10663 and asqrt[22] n10852 ; n10855
g10664 and n10334 n10855_not ; n10856
g10665 nor n10854 n10856 ; n10857
g10666 nor asqrt[25] n10837 ; n10858
g10667 and n10849_not n10858 ; n10859
g10668 nor n10857 n10859 ; n10860
g10669 nor n10851 n10860 ; n10861
g10670 and asqrt[26] n10861_not ; n10862
g10671 and n10339_not n10348 ; n10863
g10672 and n10337_not n10863 ; n10864
g10673 and asqrt[22] n10864 ; n10865
g10674 nor n10337 n10339 ; n10866
g10675 and asqrt[22] n10866 ; n10867
g10676 nor n10348 n10867 ; n10868
g10677 nor n10865 n10868 ; n10869
g10678 nor asqrt[26] n10851 ; n10870
g10679 and n10860_not n10870 ; n10871
g10680 nor n10869 n10871 ; n10872
g10681 nor n10862 n10872 ; n10873
g10682 and asqrt[27] n10873_not ; n10874
g10683 and n10351_not n10357 ; n10875
g10684 and n10359_not n10875 ; n10876
g10685 and asqrt[22] n10876 ; n10877
g10686 nor n10351 n10359 ; n10878
g10687 and asqrt[22] n10878 ; n10879
g10688 nor n10357 n10879 ; n10880
g10689 nor n10877 n10880 ; n10881
g10690 nor asqrt[27] n10862 ; n10882
g10691 and n10872_not n10882 ; n10883
g10692 nor n10881 n10883 ; n10884
g10693 nor n10874 n10884 ; n10885
g10694 and asqrt[28] n10885_not ; n10886
g10695 and n10369 n10371_not ; n10887
g10696 and n10362_not n10887 ; n10888
g10697 and asqrt[22] n10888 ; n10889
g10698 nor n10362 n10371 ; n10890
g10699 and asqrt[22] n10890 ; n10891
g10700 nor n10369 n10891 ; n10892
g10701 nor n10889 n10892 ; n10893
g10702 nor asqrt[28] n10874 ; n10894
g10703 and n10884_not n10894 ; n10895
g10704 nor n10893 n10895 ; n10896
g10705 nor n10886 n10896 ; n10897
g10706 and asqrt[29] n10897_not ; n10898
g10707 and n10374_not n10381 ; n10899
g10708 and n10383_not n10899 ; n10900
g10709 and asqrt[22] n10900 ; n10901
g10710 nor n10374 n10383 ; n10902
g10711 and asqrt[22] n10902 ; n10903
g10712 nor n10381 n10903 ; n10904
g10713 nor n10901 n10904 ; n10905
g10714 nor asqrt[29] n10886 ; n10906
g10715 and n10896_not n10906 ; n10907
g10716 nor n10905 n10907 ; n10908
g10717 nor n10898 n10908 ; n10909
g10718 and asqrt[30] n10909_not ; n10910
g10719 and n10393 n10395_not ; n10911
g10720 and n10386_not n10911 ; n10912
g10721 and asqrt[22] n10912 ; n10913
g10722 nor n10386 n10395 ; n10914
g10723 and asqrt[22] n10914 ; n10915
g10724 nor n10393 n10915 ; n10916
g10725 nor n10913 n10916 ; n10917
g10726 nor asqrt[30] n10898 ; n10918
g10727 and n10908_not n10918 ; n10919
g10728 nor n10917 n10919 ; n10920
g10729 nor n10910 n10920 ; n10921
g10730 and asqrt[31] n10921_not ; n10922
g10731 and n10398_not n10405 ; n10923
g10732 and n10407_not n10923 ; n10924
g10733 and asqrt[22] n10924 ; n10925
g10734 nor n10398 n10407 ; n10926
g10735 and asqrt[22] n10926 ; n10927
g10736 nor n10405 n10927 ; n10928
g10737 nor n10925 n10928 ; n10929
g10738 nor asqrt[31] n10910 ; n10930
g10739 and n10920_not n10930 ; n10931
g10740 nor n10929 n10931 ; n10932
g10741 nor n10922 n10932 ; n10933
g10742 and asqrt[32] n10933_not ; n10934
g10743 and n10417 n10419_not ; n10935
g10744 and n10410_not n10935 ; n10936
g10745 and asqrt[22] n10936 ; n10937
g10746 nor n10410 n10419 ; n10938
g10747 and asqrt[22] n10938 ; n10939
g10748 nor n10417 n10939 ; n10940
g10749 nor n10937 n10940 ; n10941
g10750 nor asqrt[32] n10922 ; n10942
g10751 and n10932_not n10942 ; n10943
g10752 nor n10941 n10943 ; n10944
g10753 nor n10934 n10944 ; n10945
g10754 and asqrt[33] n10945_not ; n10946
g10755 and n10422_not n10429 ; n10947
g10756 and n10431_not n10947 ; n10948
g10757 and asqrt[22] n10948 ; n10949
g10758 nor n10422 n10431 ; n10950
g10759 and asqrt[22] n10950 ; n10951
g10760 nor n10429 n10951 ; n10952
g10761 nor n10949 n10952 ; n10953
g10762 nor asqrt[33] n10934 ; n10954
g10763 and n10944_not n10954 ; n10955
g10764 nor n10953 n10955 ; n10956
g10765 nor n10946 n10956 ; n10957
g10766 and asqrt[34] n10957_not ; n10958
g10767 and n10441 n10443_not ; n10959
g10768 and n10434_not n10959 ; n10960
g10769 and asqrt[22] n10960 ; n10961
g10770 nor n10434 n10443 ; n10962
g10771 and asqrt[22] n10962 ; n10963
g10772 nor n10441 n10963 ; n10964
g10773 nor n10961 n10964 ; n10965
g10774 nor asqrt[34] n10946 ; n10966
g10775 and n10956_not n10966 ; n10967
g10776 nor n10965 n10967 ; n10968
g10777 nor n10958 n10968 ; n10969
g10778 and asqrt[35] n10969_not ; n10970
g10779 and n10446_not n10453 ; n10971
g10780 and n10455_not n10971 ; n10972
g10781 and asqrt[22] n10972 ; n10973
g10782 nor n10446 n10455 ; n10974
g10783 and asqrt[22] n10974 ; n10975
g10784 nor n10453 n10975 ; n10976
g10785 nor n10973 n10976 ; n10977
g10786 nor asqrt[35] n10958 ; n10978
g10787 and n10968_not n10978 ; n10979
g10788 nor n10977 n10979 ; n10980
g10789 nor n10970 n10980 ; n10981
g10790 and asqrt[36] n10981_not ; n10982
g10791 and n10465 n10467_not ; n10983
g10792 and n10458_not n10983 ; n10984
g10793 and asqrt[22] n10984 ; n10985
g10794 nor n10458 n10467 ; n10986
g10795 and asqrt[22] n10986 ; n10987
g10796 nor n10465 n10987 ; n10988
g10797 nor n10985 n10988 ; n10989
g10798 nor asqrt[36] n10970 ; n10990
g10799 and n10980_not n10990 ; n10991
g10800 nor n10989 n10991 ; n10992
g10801 nor n10982 n10992 ; n10993
g10802 and asqrt[37] n10993_not ; n10994
g10803 and n10470_not n10477 ; n10995
g10804 and n10479_not n10995 ; n10996
g10805 and asqrt[22] n10996 ; n10997
g10806 nor n10470 n10479 ; n10998
g10807 and asqrt[22] n10998 ; n10999
g10808 nor n10477 n10999 ; n11000
g10809 nor n10997 n11000 ; n11001
g10810 nor asqrt[37] n10982 ; n11002
g10811 and n10992_not n11002 ; n11003
g10812 nor n11001 n11003 ; n11004
g10813 nor n10994 n11004 ; n11005
g10814 and asqrt[38] n11005_not ; n11006
g10815 and n10489 n10491_not ; n11007
g10816 and n10482_not n11007 ; n11008
g10817 and asqrt[22] n11008 ; n11009
g10818 nor n10482 n10491 ; n11010
g10819 and asqrt[22] n11010 ; n11011
g10820 nor n10489 n11011 ; n11012
g10821 nor n11009 n11012 ; n11013
g10822 nor asqrt[38] n10994 ; n11014
g10823 and n11004_not n11014 ; n11015
g10824 nor n11013 n11015 ; n11016
g10825 nor n11006 n11016 ; n11017
g10826 and asqrt[39] n11017_not ; n11018
g10827 and n10494_not n10501 ; n11019
g10828 and n10503_not n11019 ; n11020
g10829 and asqrt[22] n11020 ; n11021
g10830 nor n10494 n10503 ; n11022
g10831 and asqrt[22] n11022 ; n11023
g10832 nor n10501 n11023 ; n11024
g10833 nor n11021 n11024 ; n11025
g10834 nor asqrt[39] n11006 ; n11026
g10835 and n11016_not n11026 ; n11027
g10836 nor n11025 n11027 ; n11028
g10837 nor n11018 n11028 ; n11029
g10838 and asqrt[40] n11029_not ; n11030
g10839 and n10513 n10515_not ; n11031
g10840 and n10506_not n11031 ; n11032
g10841 and asqrt[22] n11032 ; n11033
g10842 nor n10506 n10515 ; n11034
g10843 and asqrt[22] n11034 ; n11035
g10844 nor n10513 n11035 ; n11036
g10845 nor n11033 n11036 ; n11037
g10846 nor asqrt[40] n11018 ; n11038
g10847 and n11028_not n11038 ; n11039
g10848 nor n11037 n11039 ; n11040
g10849 nor n11030 n11040 ; n11041
g10850 and asqrt[41] n11041_not ; n11042
g10851 and n10518_not n10525 ; n11043
g10852 and n10527_not n11043 ; n11044
g10853 and asqrt[22] n11044 ; n11045
g10854 nor n10518 n10527 ; n11046
g10855 and asqrt[22] n11046 ; n11047
g10856 nor n10525 n11047 ; n11048
g10857 nor n11045 n11048 ; n11049
g10858 nor asqrt[41] n11030 ; n11050
g10859 and n11040_not n11050 ; n11051
g10860 nor n11049 n11051 ; n11052
g10861 nor n11042 n11052 ; n11053
g10862 and asqrt[42] n11053_not ; n11054
g10863 and n10537 n10539_not ; n11055
g10864 and n10530_not n11055 ; n11056
g10865 and asqrt[22] n11056 ; n11057
g10866 nor n10530 n10539 ; n11058
g10867 and asqrt[22] n11058 ; n11059
g10868 nor n10537 n11059 ; n11060
g10869 nor n11057 n11060 ; n11061
g10870 nor asqrt[42] n11042 ; n11062
g10871 and n11052_not n11062 ; n11063
g10872 nor n11061 n11063 ; n11064
g10873 nor n11054 n11064 ; n11065
g10874 and asqrt[43] n11065_not ; n11066
g10875 nor asqrt[43] n11054 ; n11067
g10876 and n11064_not n11067 ; n11068
g10877 and n10542_not n10551 ; n11069
g10878 and n10544_not n11069 ; n11070
g10879 and asqrt[22] n11070 ; n11071
g10880 nor n10542 n10544 ; n11072
g10881 and asqrt[22] n11072 ; n11073
g10882 nor n10551 n11073 ; n11074
g10883 nor n11071 n11074 ; n11075
g10884 nor n11068 n11075 ; n11076
g10885 nor n11066 n11076 ; n11077
g10886 and asqrt[44] n11077_not ; n11078
g10887 and n10561 n10563_not ; n11079
g10888 and n10554_not n11079 ; n11080
g10889 and asqrt[22] n11080 ; n11081
g10890 nor n10554 n10563 ; n11082
g10891 and asqrt[22] n11082 ; n11083
g10892 nor n10561 n11083 ; n11084
g10893 nor n11081 n11084 ; n11085
g10894 nor asqrt[44] n11066 ; n11086
g10895 and n11076_not n11086 ; n11087
g10896 nor n11085 n11087 ; n11088
g10897 nor n11078 n11088 ; n11089
g10898 and asqrt[45] n11089_not ; n11090
g10899 and n10566_not n10573 ; n11091
g10900 and n10575_not n11091 ; n11092
g10901 and asqrt[22] n11092 ; n11093
g10902 nor n10566 n10575 ; n11094
g10903 and asqrt[22] n11094 ; n11095
g10904 nor n10573 n11095 ; n11096
g10905 nor n11093 n11096 ; n11097
g10906 nor asqrt[45] n11078 ; n11098
g10907 and n11088_not n11098 ; n11099
g10908 nor n11097 n11099 ; n11100
g10909 nor n11090 n11100 ; n11101
g10910 and asqrt[46] n11101_not ; n11102
g10911 and n10585 n10587_not ; n11103
g10912 and n10578_not n11103 ; n11104
g10913 and asqrt[22] n11104 ; n11105
g10914 nor n10578 n10587 ; n11106
g10915 and asqrt[22] n11106 ; n11107
g10916 nor n10585 n11107 ; n11108
g10917 nor n11105 n11108 ; n11109
g10918 nor asqrt[46] n11090 ; n11110
g10919 and n11100_not n11110 ; n11111
g10920 nor n11109 n11111 ; n11112
g10921 nor n11102 n11112 ; n11113
g10922 and asqrt[47] n11113_not ; n11114
g10923 and n10590_not n10597 ; n11115
g10924 and n10599_not n11115 ; n11116
g10925 and asqrt[22] n11116 ; n11117
g10926 nor n10590 n10599 ; n11118
g10927 and asqrt[22] n11118 ; n11119
g10928 nor n10597 n11119 ; n11120
g10929 nor n11117 n11120 ; n11121
g10930 nor asqrt[47] n11102 ; n11122
g10931 and n11112_not n11122 ; n11123
g10932 nor n11121 n11123 ; n11124
g10933 nor n11114 n11124 ; n11125
g10934 and asqrt[48] n11125_not ; n11126
g10935 and n10609 n10611_not ; n11127
g10936 and n10602_not n11127 ; n11128
g10937 and asqrt[22] n11128 ; n11129
g10938 nor n10602 n10611 ; n11130
g10939 and asqrt[22] n11130 ; n11131
g10940 nor n10609 n11131 ; n11132
g10941 nor n11129 n11132 ; n11133
g10942 nor asqrt[48] n11114 ; n11134
g10943 and n11124_not n11134 ; n11135
g10944 nor n11133 n11135 ; n11136
g10945 nor n11126 n11136 ; n11137
g10946 and asqrt[49] n11137_not ; n11138
g10947 and n10614_not n10621 ; n11139
g10948 and n10623_not n11139 ; n11140
g10949 and asqrt[22] n11140 ; n11141
g10950 nor n10614 n10623 ; n11142
g10951 and asqrt[22] n11142 ; n11143
g10952 nor n10621 n11143 ; n11144
g10953 nor n11141 n11144 ; n11145
g10954 nor asqrt[49] n11126 ; n11146
g10955 and n11136_not n11146 ; n11147
g10956 nor n11145 n11147 ; n11148
g10957 nor n11138 n11148 ; n11149
g10958 and asqrt[50] n11149_not ; n11150
g10959 and n10633 n10635_not ; n11151
g10960 and n10626_not n11151 ; n11152
g10961 and asqrt[22] n11152 ; n11153
g10962 nor n10626 n10635 ; n11154
g10963 and asqrt[22] n11154 ; n11155
g10964 nor n10633 n11155 ; n11156
g10965 nor n11153 n11156 ; n11157
g10966 nor asqrt[50] n11138 ; n11158
g10967 and n11148_not n11158 ; n11159
g10968 nor n11157 n11159 ; n11160
g10969 nor n11150 n11160 ; n11161
g10970 and asqrt[51] n11161_not ; n11162
g10971 and n10638_not n10645 ; n11163
g10972 and n10647_not n11163 ; n11164
g10973 and asqrt[22] n11164 ; n11165
g10974 nor n10638 n10647 ; n11166
g10975 and asqrt[22] n11166 ; n11167
g10976 nor n10645 n11167 ; n11168
g10977 nor n11165 n11168 ; n11169
g10978 nor asqrt[51] n11150 ; n11170
g10979 and n11160_not n11170 ; n11171
g10980 nor n11169 n11171 ; n11172
g10981 nor n11162 n11172 ; n11173
g10982 and asqrt[52] n11173_not ; n11174
g10983 and n10657 n10659_not ; n11175
g10984 and n10650_not n11175 ; n11176
g10985 and asqrt[22] n11176 ; n11177
g10986 nor n10650 n10659 ; n11178
g10987 and asqrt[22] n11178 ; n11179
g10988 nor n10657 n11179 ; n11180
g10989 nor n11177 n11180 ; n11181
g10990 nor asqrt[52] n11162 ; n11182
g10991 and n11172_not n11182 ; n11183
g10992 nor n11181 n11183 ; n11184
g10993 nor n11174 n11184 ; n11185
g10994 and asqrt[53] n11185_not ; n11186
g10995 and n10662_not n10669 ; n11187
g10996 and n10671_not n11187 ; n11188
g10997 and asqrt[22] n11188 ; n11189
g10998 nor n10662 n10671 ; n11190
g10999 and asqrt[22] n11190 ; n11191
g11000 nor n10669 n11191 ; n11192
g11001 nor n11189 n11192 ; n11193
g11002 nor asqrt[53] n11174 ; n11194
g11003 and n11184_not n11194 ; n11195
g11004 nor n11193 n11195 ; n11196
g11005 nor n11186 n11196 ; n11197
g11006 and asqrt[54] n11197_not ; n11198
g11007 and n10681 n10683_not ; n11199
g11008 and n10674_not n11199 ; n11200
g11009 and asqrt[22] n11200 ; n11201
g11010 nor n10674 n10683 ; n11202
g11011 and asqrt[22] n11202 ; n11203
g11012 nor n10681 n11203 ; n11204
g11013 nor n11201 n11204 ; n11205
g11014 nor asqrt[54] n11186 ; n11206
g11015 and n11196_not n11206 ; n11207
g11016 nor n11205 n11207 ; n11208
g11017 nor n11198 n11208 ; n11209
g11018 and asqrt[55] n11209_not ; n11210
g11019 and n10686_not n10693 ; n11211
g11020 and n10695_not n11211 ; n11212
g11021 and asqrt[22] n11212 ; n11213
g11022 nor n10686 n10695 ; n11214
g11023 and asqrt[22] n11214 ; n11215
g11024 nor n10693 n11215 ; n11216
g11025 nor n11213 n11216 ; n11217
g11026 nor asqrt[55] n11198 ; n11218
g11027 and n11208_not n11218 ; n11219
g11028 nor n11217 n11219 ; n11220
g11029 nor n11210 n11220 ; n11221
g11030 and asqrt[56] n11221_not ; n11222
g11031 and n10705 n10707_not ; n11223
g11032 and n10698_not n11223 ; n11224
g11033 and asqrt[22] n11224 ; n11225
g11034 nor n10698 n10707 ; n11226
g11035 and asqrt[22] n11226 ; n11227
g11036 nor n10705 n11227 ; n11228
g11037 nor n11225 n11228 ; n11229
g11038 nor asqrt[56] n11210 ; n11230
g11039 and n11220_not n11230 ; n11231
g11040 nor n11229 n11231 ; n11232
g11041 nor n11222 n11232 ; n11233
g11042 and asqrt[57] n11233_not ; n11234
g11043 and n10710_not n10717 ; n11235
g11044 and n10719_not n11235 ; n11236
g11045 and asqrt[22] n11236 ; n11237
g11046 nor n10710 n10719 ; n11238
g11047 and asqrt[22] n11238 ; n11239
g11048 nor n10717 n11239 ; n11240
g11049 nor n11237 n11240 ; n11241
g11050 nor asqrt[57] n11222 ; n11242
g11051 and n11232_not n11242 ; n11243
g11052 nor n11241 n11243 ; n11244
g11053 nor n11234 n11244 ; n11245
g11054 and asqrt[58] n11245_not ; n11246
g11055 and n10729 n10731_not ; n11247
g11056 and n10722_not n11247 ; n11248
g11057 and asqrt[22] n11248 ; n11249
g11058 nor n10722 n10731 ; n11250
g11059 and asqrt[22] n11250 ; n11251
g11060 nor n10729 n11251 ; n11252
g11061 nor n11249 n11252 ; n11253
g11062 nor asqrt[58] n11234 ; n11254
g11063 and n11244_not n11254 ; n11255
g11064 nor n11253 n11255 ; n11256
g11065 nor n11246 n11256 ; n11257
g11066 and asqrt[59] n11257_not ; n11258
g11067 and n10734_not n10741 ; n11259
g11068 and n10743_not n11259 ; n11260
g11069 and asqrt[22] n11260 ; n11261
g11070 nor n10734 n10743 ; n11262
g11071 and asqrt[22] n11262 ; n11263
g11072 nor n10741 n11263 ; n11264
g11073 nor n11261 n11264 ; n11265
g11074 nor asqrt[59] n11246 ; n11266
g11075 and n11256_not n11266 ; n11267
g11076 nor n11265 n11267 ; n11268
g11077 nor n11258 n11268 ; n11269
g11078 and asqrt[60] n11269_not ; n11270
g11079 and n10753 n10755_not ; n11271
g11080 and n10746_not n11271 ; n11272
g11081 and asqrt[22] n11272 ; n11273
g11082 nor n10746 n10755 ; n11274
g11083 and asqrt[22] n11274 ; n11275
g11084 nor n10753 n11275 ; n11276
g11085 nor n11273 n11276 ; n11277
g11086 nor asqrt[60] n11258 ; n11278
g11087 and n11268_not n11278 ; n11279
g11088 nor n11277 n11279 ; n11280
g11089 nor n11270 n11280 ; n11281
g11090 and asqrt[61] n11281_not ; n11282
g11091 and n10758_not n10765 ; n11283
g11092 and n10767_not n11283 ; n11284
g11093 and asqrt[22] n11284 ; n11285
g11094 nor n10758 n10767 ; n11286
g11095 and asqrt[22] n11286 ; n11287
g11096 nor n10765 n11287 ; n11288
g11097 nor n11285 n11288 ; n11289
g11098 nor asqrt[61] n11270 ; n11290
g11099 and n11280_not n11290 ; n11291
g11100 nor n11289 n11291 ; n11292
g11101 nor n11282 n11292 ; n11293
g11102 and asqrt[62] n11293_not ; n11294
g11103 and n10777 n10779_not ; n11295
g11104 and n10770_not n11295 ; n11296
g11105 and asqrt[22] n11296 ; n11297
g11106 nor n10770 n10779 ; n11298
g11107 and asqrt[22] n11298 ; n11299
g11108 nor n10777 n11299 ; n11300
g11109 nor n11297 n11300 ; n11301
g11110 nor asqrt[62] n11282 ; n11302
g11111 and n11292_not n11302 ; n11303
g11112 nor n11301 n11303 ; n11304
g11113 nor n11294 n11304 ; n11305
g11114 and n10782_not n10789 ; n11306
g11115 and n10791_not n11306 ; n11307
g11116 and asqrt[22] n11307 ; n11308
g11117 nor n10782 n10791 ; n11309
g11118 and asqrt[22] n11309 ; n11310
g11119 nor n10789 n11310 ; n11311
g11120 nor n11308 n11311 ; n11312
g11121 nor n10793 n10800 ; n11313
g11122 and asqrt[22] n11313 ; n11314
g11123 nor n10808 n11314 ; n11315
g11124 and n11312_not n11315 ; n11316
g11125 and n11305_not n11316 ; n11317
g11126 nor asqrt[63] n11317 ; n11318
g11127 and n11294_not n11312 ; n11319
g11128 and n11304_not n11319 ; n11320
g11129 and n10800_not asqrt[22] ; n11321
g11130 and n10793 n11321_not ; n11322
g11131 and asqrt[63] n11313_not ; n11323
g11132 and n11322_not n11323 ; n11324
g11133 nor n10796 n10817 ; n11325
g11134 and n10799_not n11325 ; n11326
g11135 and n10812_not n11326 ; n11327
g11136 and n10808_not n11327 ; n11328
g11137 and n10806_not n11328 ; n11329
g11138 nor n11324 n11329 ; n11330
g11139 and n11320_not n11330 ; n11331
g11140 nand n11318_not n11331 ; asqrt[21]
g11141 and a[42] asqrt[21] ; n11333
g11142 nor a[40] a[41] ; n11334
g11143 and a[42]_not n11334 ; n11335
g11144 nor n11333 n11335 ; n11336
g11145 and asqrt[22] n11336_not ; n11337
g11146 nor n10817 n11335 ; n11338
g11147 and n10812_not n11338 ; n11339
g11148 and n10808_not n11339 ; n11340
g11149 and n10806_not n11340 ; n11341
g11150 and n11333_not n11341 ; n11342
g11151 and a[42]_not asqrt[21] ; n11343
g11152 and a[43] n11343_not ; n11344
g11153 and n10822 asqrt[21] ; n11345
g11154 nor n11344 n11345 ; n11346
g11155 and n11342_not n11346 ; n11347
g11156 nor n11337 n11347 ; n11348
g11157 and asqrt[23] n11348_not ; n11349
g11158 nor asqrt[23] n11337 ; n11350
g11159 and n11347_not n11350 ; n11351
g11160 and asqrt[22] n11329_not ; n11352
g11161 and n11324_not n11352 ; n11353
g11162 and n11320_not n11353 ; n11354
g11163 and n11318_not n11354 ; n11355
g11164 nor n11345 n11355 ; n11356
g11165 and a[44] n11356_not ; n11357
g11166 nor a[44] n11355 ; n11358
g11167 and n11345_not n11358 ; n11359
g11168 nor n11357 n11359 ; n11360
g11169 nor n11351 n11360 ; n11361
g11170 nor n11349 n11361 ; n11362
g11171 and asqrt[24] n11362_not ; n11363
g11172 nor n10825 n10830 ; n11364
g11173 and n10834_not n11364 ; n11365
g11174 and asqrt[21] n11365 ; n11366
g11175 and asqrt[21] n11364 ; n11367
g11176 and n10834 n11367_not ; n11368
g11177 nor n11366 n11368 ; n11369
g11178 nor asqrt[24] n11349 ; n11370
g11179 and n11361_not n11370 ; n11371
g11180 nor n11369 n11371 ; n11372
g11181 nor n11363 n11372 ; n11373
g11182 and asqrt[25] n11373_not ; n11374
g11183 and n10839_not n10848 ; n11375
g11184 and n10837_not n11375 ; n11376
g11185 and asqrt[21] n11376 ; n11377
g11186 nor n10837 n10839 ; n11378
g11187 and asqrt[21] n11378 ; n11379
g11188 nor n10848 n11379 ; n11380
g11189 nor n11377 n11380 ; n11381
g11190 nor asqrt[25] n11363 ; n11382
g11191 and n11372_not n11382 ; n11383
g11192 nor n11381 n11383 ; n11384
g11193 nor n11374 n11384 ; n11385
g11194 and asqrt[26] n11385_not ; n11386
g11195 and n10851_not n10857 ; n11387
g11196 and n10859_not n11387 ; n11388
g11197 and asqrt[21] n11388 ; n11389
g11198 nor n10851 n10859 ; n11390
g11199 and asqrt[21] n11390 ; n11391
g11200 nor n10857 n11391 ; n11392
g11201 nor n11389 n11392 ; n11393
g11202 nor asqrt[26] n11374 ; n11394
g11203 and n11384_not n11394 ; n11395
g11204 nor n11393 n11395 ; n11396
g11205 nor n11386 n11396 ; n11397
g11206 and asqrt[27] n11397_not ; n11398
g11207 and n10869 n10871_not ; n11399
g11208 and n10862_not n11399 ; n11400
g11209 and asqrt[21] n11400 ; n11401
g11210 nor n10862 n10871 ; n11402
g11211 and asqrt[21] n11402 ; n11403
g11212 nor n10869 n11403 ; n11404
g11213 nor n11401 n11404 ; n11405
g11214 nor asqrt[27] n11386 ; n11406
g11215 and n11396_not n11406 ; n11407
g11216 nor n11405 n11407 ; n11408
g11217 nor n11398 n11408 ; n11409
g11218 and asqrt[28] n11409_not ; n11410
g11219 and n10874_not n10881 ; n11411
g11220 and n10883_not n11411 ; n11412
g11221 and asqrt[21] n11412 ; n11413
g11222 nor n10874 n10883 ; n11414
g11223 and asqrt[21] n11414 ; n11415
g11224 nor n10881 n11415 ; n11416
g11225 nor n11413 n11416 ; n11417
g11226 nor asqrt[28] n11398 ; n11418
g11227 and n11408_not n11418 ; n11419
g11228 nor n11417 n11419 ; n11420
g11229 nor n11410 n11420 ; n11421
g11230 and asqrt[29] n11421_not ; n11422
g11231 and n10893 n10895_not ; n11423
g11232 and n10886_not n11423 ; n11424
g11233 and asqrt[21] n11424 ; n11425
g11234 nor n10886 n10895 ; n11426
g11235 and asqrt[21] n11426 ; n11427
g11236 nor n10893 n11427 ; n11428
g11237 nor n11425 n11428 ; n11429
g11238 nor asqrt[29] n11410 ; n11430
g11239 and n11420_not n11430 ; n11431
g11240 nor n11429 n11431 ; n11432
g11241 nor n11422 n11432 ; n11433
g11242 and asqrt[30] n11433_not ; n11434
g11243 and n10898_not n10905 ; n11435
g11244 and n10907_not n11435 ; n11436
g11245 and asqrt[21] n11436 ; n11437
g11246 nor n10898 n10907 ; n11438
g11247 and asqrt[21] n11438 ; n11439
g11248 nor n10905 n11439 ; n11440
g11249 nor n11437 n11440 ; n11441
g11250 nor asqrt[30] n11422 ; n11442
g11251 and n11432_not n11442 ; n11443
g11252 nor n11441 n11443 ; n11444
g11253 nor n11434 n11444 ; n11445
g11254 and asqrt[31] n11445_not ; n11446
g11255 and n10917 n10919_not ; n11447
g11256 and n10910_not n11447 ; n11448
g11257 and asqrt[21] n11448 ; n11449
g11258 nor n10910 n10919 ; n11450
g11259 and asqrt[21] n11450 ; n11451
g11260 nor n10917 n11451 ; n11452
g11261 nor n11449 n11452 ; n11453
g11262 nor asqrt[31] n11434 ; n11454
g11263 and n11444_not n11454 ; n11455
g11264 nor n11453 n11455 ; n11456
g11265 nor n11446 n11456 ; n11457
g11266 and asqrt[32] n11457_not ; n11458
g11267 and n10922_not n10929 ; n11459
g11268 and n10931_not n11459 ; n11460
g11269 and asqrt[21] n11460 ; n11461
g11270 nor n10922 n10931 ; n11462
g11271 and asqrt[21] n11462 ; n11463
g11272 nor n10929 n11463 ; n11464
g11273 nor n11461 n11464 ; n11465
g11274 nor asqrt[32] n11446 ; n11466
g11275 and n11456_not n11466 ; n11467
g11276 nor n11465 n11467 ; n11468
g11277 nor n11458 n11468 ; n11469
g11278 and asqrt[33] n11469_not ; n11470
g11279 and n10941 n10943_not ; n11471
g11280 and n10934_not n11471 ; n11472
g11281 and asqrt[21] n11472 ; n11473
g11282 nor n10934 n10943 ; n11474
g11283 and asqrt[21] n11474 ; n11475
g11284 nor n10941 n11475 ; n11476
g11285 nor n11473 n11476 ; n11477
g11286 nor asqrt[33] n11458 ; n11478
g11287 and n11468_not n11478 ; n11479
g11288 nor n11477 n11479 ; n11480
g11289 nor n11470 n11480 ; n11481
g11290 and asqrt[34] n11481_not ; n11482
g11291 and n10946_not n10953 ; n11483
g11292 and n10955_not n11483 ; n11484
g11293 and asqrt[21] n11484 ; n11485
g11294 nor n10946 n10955 ; n11486
g11295 and asqrt[21] n11486 ; n11487
g11296 nor n10953 n11487 ; n11488
g11297 nor n11485 n11488 ; n11489
g11298 nor asqrt[34] n11470 ; n11490
g11299 and n11480_not n11490 ; n11491
g11300 nor n11489 n11491 ; n11492
g11301 nor n11482 n11492 ; n11493
g11302 and asqrt[35] n11493_not ; n11494
g11303 and n10965 n10967_not ; n11495
g11304 and n10958_not n11495 ; n11496
g11305 and asqrt[21] n11496 ; n11497
g11306 nor n10958 n10967 ; n11498
g11307 and asqrt[21] n11498 ; n11499
g11308 nor n10965 n11499 ; n11500
g11309 nor n11497 n11500 ; n11501
g11310 nor asqrt[35] n11482 ; n11502
g11311 and n11492_not n11502 ; n11503
g11312 nor n11501 n11503 ; n11504
g11313 nor n11494 n11504 ; n11505
g11314 and asqrt[36] n11505_not ; n11506
g11315 and n10970_not n10977 ; n11507
g11316 and n10979_not n11507 ; n11508
g11317 and asqrt[21] n11508 ; n11509
g11318 nor n10970 n10979 ; n11510
g11319 and asqrt[21] n11510 ; n11511
g11320 nor n10977 n11511 ; n11512
g11321 nor n11509 n11512 ; n11513
g11322 nor asqrt[36] n11494 ; n11514
g11323 and n11504_not n11514 ; n11515
g11324 nor n11513 n11515 ; n11516
g11325 nor n11506 n11516 ; n11517
g11326 and asqrt[37] n11517_not ; n11518
g11327 and n10989 n10991_not ; n11519
g11328 and n10982_not n11519 ; n11520
g11329 and asqrt[21] n11520 ; n11521
g11330 nor n10982 n10991 ; n11522
g11331 and asqrt[21] n11522 ; n11523
g11332 nor n10989 n11523 ; n11524
g11333 nor n11521 n11524 ; n11525
g11334 nor asqrt[37] n11506 ; n11526
g11335 and n11516_not n11526 ; n11527
g11336 nor n11525 n11527 ; n11528
g11337 nor n11518 n11528 ; n11529
g11338 and asqrt[38] n11529_not ; n11530
g11339 and n10994_not n11001 ; n11531
g11340 and n11003_not n11531 ; n11532
g11341 and asqrt[21] n11532 ; n11533
g11342 nor n10994 n11003 ; n11534
g11343 and asqrt[21] n11534 ; n11535
g11344 nor n11001 n11535 ; n11536
g11345 nor n11533 n11536 ; n11537
g11346 nor asqrt[38] n11518 ; n11538
g11347 and n11528_not n11538 ; n11539
g11348 nor n11537 n11539 ; n11540
g11349 nor n11530 n11540 ; n11541
g11350 and asqrt[39] n11541_not ; n11542
g11351 and n11013 n11015_not ; n11543
g11352 and n11006_not n11543 ; n11544
g11353 and asqrt[21] n11544 ; n11545
g11354 nor n11006 n11015 ; n11546
g11355 and asqrt[21] n11546 ; n11547
g11356 nor n11013 n11547 ; n11548
g11357 nor n11545 n11548 ; n11549
g11358 nor asqrt[39] n11530 ; n11550
g11359 and n11540_not n11550 ; n11551
g11360 nor n11549 n11551 ; n11552
g11361 nor n11542 n11552 ; n11553
g11362 and asqrt[40] n11553_not ; n11554
g11363 and n11018_not n11025 ; n11555
g11364 and n11027_not n11555 ; n11556
g11365 and asqrt[21] n11556 ; n11557
g11366 nor n11018 n11027 ; n11558
g11367 and asqrt[21] n11558 ; n11559
g11368 nor n11025 n11559 ; n11560
g11369 nor n11557 n11560 ; n11561
g11370 nor asqrt[40] n11542 ; n11562
g11371 and n11552_not n11562 ; n11563
g11372 nor n11561 n11563 ; n11564
g11373 nor n11554 n11564 ; n11565
g11374 and asqrt[41] n11565_not ; n11566
g11375 and n11037 n11039_not ; n11567
g11376 and n11030_not n11567 ; n11568
g11377 and asqrt[21] n11568 ; n11569
g11378 nor n11030 n11039 ; n11570
g11379 and asqrt[21] n11570 ; n11571
g11380 nor n11037 n11571 ; n11572
g11381 nor n11569 n11572 ; n11573
g11382 nor asqrt[41] n11554 ; n11574
g11383 and n11564_not n11574 ; n11575
g11384 nor n11573 n11575 ; n11576
g11385 nor n11566 n11576 ; n11577
g11386 and asqrt[42] n11577_not ; n11578
g11387 and n11042_not n11049 ; n11579
g11388 and n11051_not n11579 ; n11580
g11389 and asqrt[21] n11580 ; n11581
g11390 nor n11042 n11051 ; n11582
g11391 and asqrt[21] n11582 ; n11583
g11392 nor n11049 n11583 ; n11584
g11393 nor n11581 n11584 ; n11585
g11394 nor asqrt[42] n11566 ; n11586
g11395 and n11576_not n11586 ; n11587
g11396 nor n11585 n11587 ; n11588
g11397 nor n11578 n11588 ; n11589
g11398 and asqrt[43] n11589_not ; n11590
g11399 and n11061 n11063_not ; n11591
g11400 and n11054_not n11591 ; n11592
g11401 and asqrt[21] n11592 ; n11593
g11402 nor n11054 n11063 ; n11594
g11403 and asqrt[21] n11594 ; n11595
g11404 nor n11061 n11595 ; n11596
g11405 nor n11593 n11596 ; n11597
g11406 nor asqrt[43] n11578 ; n11598
g11407 and n11588_not n11598 ; n11599
g11408 nor n11597 n11599 ; n11600
g11409 nor n11590 n11600 ; n11601
g11410 and asqrt[44] n11601_not ; n11602
g11411 nor asqrt[44] n11590 ; n11603
g11412 and n11600_not n11603 ; n11604
g11413 and n11066_not n11075 ; n11605
g11414 and n11068_not n11605 ; n11606
g11415 and asqrt[21] n11606 ; n11607
g11416 nor n11066 n11068 ; n11608
g11417 and asqrt[21] n11608 ; n11609
g11418 nor n11075 n11609 ; n11610
g11419 nor n11607 n11610 ; n11611
g11420 nor n11604 n11611 ; n11612
g11421 nor n11602 n11612 ; n11613
g11422 and asqrt[45] n11613_not ; n11614
g11423 and n11085 n11087_not ; n11615
g11424 and n11078_not n11615 ; n11616
g11425 and asqrt[21] n11616 ; n11617
g11426 nor n11078 n11087 ; n11618
g11427 and asqrt[21] n11618 ; n11619
g11428 nor n11085 n11619 ; n11620
g11429 nor n11617 n11620 ; n11621
g11430 nor asqrt[45] n11602 ; n11622
g11431 and n11612_not n11622 ; n11623
g11432 nor n11621 n11623 ; n11624
g11433 nor n11614 n11624 ; n11625
g11434 and asqrt[46] n11625_not ; n11626
g11435 and n11090_not n11097 ; n11627
g11436 and n11099_not n11627 ; n11628
g11437 and asqrt[21] n11628 ; n11629
g11438 nor n11090 n11099 ; n11630
g11439 and asqrt[21] n11630 ; n11631
g11440 nor n11097 n11631 ; n11632
g11441 nor n11629 n11632 ; n11633
g11442 nor asqrt[46] n11614 ; n11634
g11443 and n11624_not n11634 ; n11635
g11444 nor n11633 n11635 ; n11636
g11445 nor n11626 n11636 ; n11637
g11446 and asqrt[47] n11637_not ; n11638
g11447 and n11109 n11111_not ; n11639
g11448 and n11102_not n11639 ; n11640
g11449 and asqrt[21] n11640 ; n11641
g11450 nor n11102 n11111 ; n11642
g11451 and asqrt[21] n11642 ; n11643
g11452 nor n11109 n11643 ; n11644
g11453 nor n11641 n11644 ; n11645
g11454 nor asqrt[47] n11626 ; n11646
g11455 and n11636_not n11646 ; n11647
g11456 nor n11645 n11647 ; n11648
g11457 nor n11638 n11648 ; n11649
g11458 and asqrt[48] n11649_not ; n11650
g11459 and n11114_not n11121 ; n11651
g11460 and n11123_not n11651 ; n11652
g11461 and asqrt[21] n11652 ; n11653
g11462 nor n11114 n11123 ; n11654
g11463 and asqrt[21] n11654 ; n11655
g11464 nor n11121 n11655 ; n11656
g11465 nor n11653 n11656 ; n11657
g11466 nor asqrt[48] n11638 ; n11658
g11467 and n11648_not n11658 ; n11659
g11468 nor n11657 n11659 ; n11660
g11469 nor n11650 n11660 ; n11661
g11470 and asqrt[49] n11661_not ; n11662
g11471 and n11133 n11135_not ; n11663
g11472 and n11126_not n11663 ; n11664
g11473 and asqrt[21] n11664 ; n11665
g11474 nor n11126 n11135 ; n11666
g11475 and asqrt[21] n11666 ; n11667
g11476 nor n11133 n11667 ; n11668
g11477 nor n11665 n11668 ; n11669
g11478 nor asqrt[49] n11650 ; n11670
g11479 and n11660_not n11670 ; n11671
g11480 nor n11669 n11671 ; n11672
g11481 nor n11662 n11672 ; n11673
g11482 and asqrt[50] n11673_not ; n11674
g11483 and n11138_not n11145 ; n11675
g11484 and n11147_not n11675 ; n11676
g11485 and asqrt[21] n11676 ; n11677
g11486 nor n11138 n11147 ; n11678
g11487 and asqrt[21] n11678 ; n11679
g11488 nor n11145 n11679 ; n11680
g11489 nor n11677 n11680 ; n11681
g11490 nor asqrt[50] n11662 ; n11682
g11491 and n11672_not n11682 ; n11683
g11492 nor n11681 n11683 ; n11684
g11493 nor n11674 n11684 ; n11685
g11494 and asqrt[51] n11685_not ; n11686
g11495 and n11157 n11159_not ; n11687
g11496 and n11150_not n11687 ; n11688
g11497 and asqrt[21] n11688 ; n11689
g11498 nor n11150 n11159 ; n11690
g11499 and asqrt[21] n11690 ; n11691
g11500 nor n11157 n11691 ; n11692
g11501 nor n11689 n11692 ; n11693
g11502 nor asqrt[51] n11674 ; n11694
g11503 and n11684_not n11694 ; n11695
g11504 nor n11693 n11695 ; n11696
g11505 nor n11686 n11696 ; n11697
g11506 and asqrt[52] n11697_not ; n11698
g11507 and n11162_not n11169 ; n11699
g11508 and n11171_not n11699 ; n11700
g11509 and asqrt[21] n11700 ; n11701
g11510 nor n11162 n11171 ; n11702
g11511 and asqrt[21] n11702 ; n11703
g11512 nor n11169 n11703 ; n11704
g11513 nor n11701 n11704 ; n11705
g11514 nor asqrt[52] n11686 ; n11706
g11515 and n11696_not n11706 ; n11707
g11516 nor n11705 n11707 ; n11708
g11517 nor n11698 n11708 ; n11709
g11518 and asqrt[53] n11709_not ; n11710
g11519 and n11181 n11183_not ; n11711
g11520 and n11174_not n11711 ; n11712
g11521 and asqrt[21] n11712 ; n11713
g11522 nor n11174 n11183 ; n11714
g11523 and asqrt[21] n11714 ; n11715
g11524 nor n11181 n11715 ; n11716
g11525 nor n11713 n11716 ; n11717
g11526 nor asqrt[53] n11698 ; n11718
g11527 and n11708_not n11718 ; n11719
g11528 nor n11717 n11719 ; n11720
g11529 nor n11710 n11720 ; n11721
g11530 and asqrt[54] n11721_not ; n11722
g11531 and n11186_not n11193 ; n11723
g11532 and n11195_not n11723 ; n11724
g11533 and asqrt[21] n11724 ; n11725
g11534 nor n11186 n11195 ; n11726
g11535 and asqrt[21] n11726 ; n11727
g11536 nor n11193 n11727 ; n11728
g11537 nor n11725 n11728 ; n11729
g11538 nor asqrt[54] n11710 ; n11730
g11539 and n11720_not n11730 ; n11731
g11540 nor n11729 n11731 ; n11732
g11541 nor n11722 n11732 ; n11733
g11542 and asqrt[55] n11733_not ; n11734
g11543 and n11205 n11207_not ; n11735
g11544 and n11198_not n11735 ; n11736
g11545 and asqrt[21] n11736 ; n11737
g11546 nor n11198 n11207 ; n11738
g11547 and asqrt[21] n11738 ; n11739
g11548 nor n11205 n11739 ; n11740
g11549 nor n11737 n11740 ; n11741
g11550 nor asqrt[55] n11722 ; n11742
g11551 and n11732_not n11742 ; n11743
g11552 nor n11741 n11743 ; n11744
g11553 nor n11734 n11744 ; n11745
g11554 and asqrt[56] n11745_not ; n11746
g11555 and n11210_not n11217 ; n11747
g11556 and n11219_not n11747 ; n11748
g11557 and asqrt[21] n11748 ; n11749
g11558 nor n11210 n11219 ; n11750
g11559 and asqrt[21] n11750 ; n11751
g11560 nor n11217 n11751 ; n11752
g11561 nor n11749 n11752 ; n11753
g11562 nor asqrt[56] n11734 ; n11754
g11563 and n11744_not n11754 ; n11755
g11564 nor n11753 n11755 ; n11756
g11565 nor n11746 n11756 ; n11757
g11566 and asqrt[57] n11757_not ; n11758
g11567 and n11229 n11231_not ; n11759
g11568 and n11222_not n11759 ; n11760
g11569 and asqrt[21] n11760 ; n11761
g11570 nor n11222 n11231 ; n11762
g11571 and asqrt[21] n11762 ; n11763
g11572 nor n11229 n11763 ; n11764
g11573 nor n11761 n11764 ; n11765
g11574 nor asqrt[57] n11746 ; n11766
g11575 and n11756_not n11766 ; n11767
g11576 nor n11765 n11767 ; n11768
g11577 nor n11758 n11768 ; n11769
g11578 and asqrt[58] n11769_not ; n11770
g11579 and n11234_not n11241 ; n11771
g11580 and n11243_not n11771 ; n11772
g11581 and asqrt[21] n11772 ; n11773
g11582 nor n11234 n11243 ; n11774
g11583 and asqrt[21] n11774 ; n11775
g11584 nor n11241 n11775 ; n11776
g11585 nor n11773 n11776 ; n11777
g11586 nor asqrt[58] n11758 ; n11778
g11587 and n11768_not n11778 ; n11779
g11588 nor n11777 n11779 ; n11780
g11589 nor n11770 n11780 ; n11781
g11590 and asqrt[59] n11781_not ; n11782
g11591 and n11253 n11255_not ; n11783
g11592 and n11246_not n11783 ; n11784
g11593 and asqrt[21] n11784 ; n11785
g11594 nor n11246 n11255 ; n11786
g11595 and asqrt[21] n11786 ; n11787
g11596 nor n11253 n11787 ; n11788
g11597 nor n11785 n11788 ; n11789
g11598 nor asqrt[59] n11770 ; n11790
g11599 and n11780_not n11790 ; n11791
g11600 nor n11789 n11791 ; n11792
g11601 nor n11782 n11792 ; n11793
g11602 and asqrt[60] n11793_not ; n11794
g11603 and n11258_not n11265 ; n11795
g11604 and n11267_not n11795 ; n11796
g11605 and asqrt[21] n11796 ; n11797
g11606 nor n11258 n11267 ; n11798
g11607 and asqrt[21] n11798 ; n11799
g11608 nor n11265 n11799 ; n11800
g11609 nor n11797 n11800 ; n11801
g11610 nor asqrt[60] n11782 ; n11802
g11611 and n11792_not n11802 ; n11803
g11612 nor n11801 n11803 ; n11804
g11613 nor n11794 n11804 ; n11805
g11614 and asqrt[61] n11805_not ; n11806
g11615 and n11277 n11279_not ; n11807
g11616 and n11270_not n11807 ; n11808
g11617 and asqrt[21] n11808 ; n11809
g11618 nor n11270 n11279 ; n11810
g11619 and asqrt[21] n11810 ; n11811
g11620 nor n11277 n11811 ; n11812
g11621 nor n11809 n11812 ; n11813
g11622 nor asqrt[61] n11794 ; n11814
g11623 and n11804_not n11814 ; n11815
g11624 nor n11813 n11815 ; n11816
g11625 nor n11806 n11816 ; n11817
g11626 and asqrt[62] n11817_not ; n11818
g11627 and n11282_not n11289 ; n11819
g11628 and n11291_not n11819 ; n11820
g11629 and asqrt[21] n11820 ; n11821
g11630 nor n11282 n11291 ; n11822
g11631 and asqrt[21] n11822 ; n11823
g11632 nor n11289 n11823 ; n11824
g11633 nor n11821 n11824 ; n11825
g11634 nor asqrt[62] n11806 ; n11826
g11635 and n11816_not n11826 ; n11827
g11636 nor n11825 n11827 ; n11828
g11637 nor n11818 n11828 ; n11829
g11638 and n11301 n11303_not ; n11830
g11639 and n11294_not n11830 ; n11831
g11640 and asqrt[21] n11831 ; n11832
g11641 nor n11294 n11303 ; n11833
g11642 and asqrt[21] n11833 ; n11834
g11643 nor n11301 n11834 ; n11835
g11644 nor n11832 n11835 ; n11836
g11645 nor n11305 n11312 ; n11837
g11646 and asqrt[21] n11837 ; n11838
g11647 nor n11320 n11838 ; n11839
g11648 and n11836_not n11839 ; n11840
g11649 and n11829_not n11840 ; n11841
g11650 nor asqrt[63] n11841 ; n11842
g11651 and n11818_not n11836 ; n11843
g11652 and n11828_not n11843 ; n11844
g11653 and n11312_not asqrt[21] ; n11845
g11654 and n11305 n11845_not ; n11846
g11655 and asqrt[63] n11837_not ; n11847
g11656 and n11846_not n11847 ; n11848
g11657 nor n11308 n11329 ; n11849
g11658 and n11311_not n11849 ; n11850
g11659 and n11324_not n11850 ; n11851
g11660 and n11320_not n11851 ; n11852
g11661 and n11318_not n11852 ; n11853
g11662 nor n11848 n11853 ; n11854
g11663 and n11844_not n11854 ; n11855
g11664 nand n11842_not n11855 ; asqrt[20]
g11665 and a[40] asqrt[20] ; n11857
g11666 nor a[38] a[39] ; n11858
g11667 and a[40]_not n11858 ; n11859
g11668 nor n11857 n11859 ; n11860
g11669 and asqrt[21] n11860_not ; n11861
g11670 nor n11329 n11859 ; n11862
g11671 and n11324_not n11862 ; n11863
g11672 and n11320_not n11863 ; n11864
g11673 and n11318_not n11864 ; n11865
g11674 and n11857_not n11865 ; n11866
g11675 and a[40]_not asqrt[20] ; n11867
g11676 and a[41] n11867_not ; n11868
g11677 and n11334 asqrt[20] ; n11869
g11678 nor n11868 n11869 ; n11870
g11679 and n11866_not n11870 ; n11871
g11680 nor n11861 n11871 ; n11872
g11681 and asqrt[22] n11872_not ; n11873
g11682 nor asqrt[22] n11861 ; n11874
g11683 and n11871_not n11874 ; n11875
g11684 and asqrt[21] n11853_not ; n11876
g11685 and n11848_not n11876 ; n11877
g11686 and n11844_not n11877 ; n11878
g11687 and n11842_not n11878 ; n11879
g11688 nor n11869 n11879 ; n11880
g11689 and a[42] n11880_not ; n11881
g11690 nor a[42] n11879 ; n11882
g11691 and n11869_not n11882 ; n11883
g11692 nor n11881 n11883 ; n11884
g11693 nor n11875 n11884 ; n11885
g11694 nor n11873 n11885 ; n11886
g11695 and asqrt[23] n11886_not ; n11887
g11696 nor n11337 n11342 ; n11888
g11697 and n11346_not n11888 ; n11889
g11698 and asqrt[20] n11889 ; n11890
g11699 and asqrt[20] n11888 ; n11891
g11700 and n11346 n11891_not ; n11892
g11701 nor n11890 n11892 ; n11893
g11702 nor asqrt[23] n11873 ; n11894
g11703 and n11885_not n11894 ; n11895
g11704 nor n11893 n11895 ; n11896
g11705 nor n11887 n11896 ; n11897
g11706 and asqrt[24] n11897_not ; n11898
g11707 and n11351_not n11360 ; n11899
g11708 and n11349_not n11899 ; n11900
g11709 and asqrt[20] n11900 ; n11901
g11710 nor n11349 n11351 ; n11902
g11711 and asqrt[20] n11902 ; n11903
g11712 nor n11360 n11903 ; n11904
g11713 nor n11901 n11904 ; n11905
g11714 nor asqrt[24] n11887 ; n11906
g11715 and n11896_not n11906 ; n11907
g11716 nor n11905 n11907 ; n11908
g11717 nor n11898 n11908 ; n11909
g11718 and asqrt[25] n11909_not ; n11910
g11719 and n11363_not n11369 ; n11911
g11720 and n11371_not n11911 ; n11912
g11721 and asqrt[20] n11912 ; n11913
g11722 nor n11363 n11371 ; n11914
g11723 and asqrt[20] n11914 ; n11915
g11724 nor n11369 n11915 ; n11916
g11725 nor n11913 n11916 ; n11917
g11726 nor asqrt[25] n11898 ; n11918
g11727 and n11908_not n11918 ; n11919
g11728 nor n11917 n11919 ; n11920
g11729 nor n11910 n11920 ; n11921
g11730 and asqrt[26] n11921_not ; n11922
g11731 and n11381 n11383_not ; n11923
g11732 and n11374_not n11923 ; n11924
g11733 and asqrt[20] n11924 ; n11925
g11734 nor n11374 n11383 ; n11926
g11735 and asqrt[20] n11926 ; n11927
g11736 nor n11381 n11927 ; n11928
g11737 nor n11925 n11928 ; n11929
g11738 nor asqrt[26] n11910 ; n11930
g11739 and n11920_not n11930 ; n11931
g11740 nor n11929 n11931 ; n11932
g11741 nor n11922 n11932 ; n11933
g11742 and asqrt[27] n11933_not ; n11934
g11743 and n11386_not n11393 ; n11935
g11744 and n11395_not n11935 ; n11936
g11745 and asqrt[20] n11936 ; n11937
g11746 nor n11386 n11395 ; n11938
g11747 and asqrt[20] n11938 ; n11939
g11748 nor n11393 n11939 ; n11940
g11749 nor n11937 n11940 ; n11941
g11750 nor asqrt[27] n11922 ; n11942
g11751 and n11932_not n11942 ; n11943
g11752 nor n11941 n11943 ; n11944
g11753 nor n11934 n11944 ; n11945
g11754 and asqrt[28] n11945_not ; n11946
g11755 and n11405 n11407_not ; n11947
g11756 and n11398_not n11947 ; n11948
g11757 and asqrt[20] n11948 ; n11949
g11758 nor n11398 n11407 ; n11950
g11759 and asqrt[20] n11950 ; n11951
g11760 nor n11405 n11951 ; n11952
g11761 nor n11949 n11952 ; n11953
g11762 nor asqrt[28] n11934 ; n11954
g11763 and n11944_not n11954 ; n11955
g11764 nor n11953 n11955 ; n11956
g11765 nor n11946 n11956 ; n11957
g11766 and asqrt[29] n11957_not ; n11958
g11767 and n11410_not n11417 ; n11959
g11768 and n11419_not n11959 ; n11960
g11769 and asqrt[20] n11960 ; n11961
g11770 nor n11410 n11419 ; n11962
g11771 and asqrt[20] n11962 ; n11963
g11772 nor n11417 n11963 ; n11964
g11773 nor n11961 n11964 ; n11965
g11774 nor asqrt[29] n11946 ; n11966
g11775 and n11956_not n11966 ; n11967
g11776 nor n11965 n11967 ; n11968
g11777 nor n11958 n11968 ; n11969
g11778 and asqrt[30] n11969_not ; n11970
g11779 and n11429 n11431_not ; n11971
g11780 and n11422_not n11971 ; n11972
g11781 and asqrt[20] n11972 ; n11973
g11782 nor n11422 n11431 ; n11974
g11783 and asqrt[20] n11974 ; n11975
g11784 nor n11429 n11975 ; n11976
g11785 nor n11973 n11976 ; n11977
g11786 nor asqrt[30] n11958 ; n11978
g11787 and n11968_not n11978 ; n11979
g11788 nor n11977 n11979 ; n11980
g11789 nor n11970 n11980 ; n11981
g11790 and asqrt[31] n11981_not ; n11982
g11791 and n11434_not n11441 ; n11983
g11792 and n11443_not n11983 ; n11984
g11793 and asqrt[20] n11984 ; n11985
g11794 nor n11434 n11443 ; n11986
g11795 and asqrt[20] n11986 ; n11987
g11796 nor n11441 n11987 ; n11988
g11797 nor n11985 n11988 ; n11989
g11798 nor asqrt[31] n11970 ; n11990
g11799 and n11980_not n11990 ; n11991
g11800 nor n11989 n11991 ; n11992
g11801 nor n11982 n11992 ; n11993
g11802 and asqrt[32] n11993_not ; n11994
g11803 and n11453 n11455_not ; n11995
g11804 and n11446_not n11995 ; n11996
g11805 and asqrt[20] n11996 ; n11997
g11806 nor n11446 n11455 ; n11998
g11807 and asqrt[20] n11998 ; n11999
g11808 nor n11453 n11999 ; n12000
g11809 nor n11997 n12000 ; n12001
g11810 nor asqrt[32] n11982 ; n12002
g11811 and n11992_not n12002 ; n12003
g11812 nor n12001 n12003 ; n12004
g11813 nor n11994 n12004 ; n12005
g11814 and asqrt[33] n12005_not ; n12006
g11815 and n11458_not n11465 ; n12007
g11816 and n11467_not n12007 ; n12008
g11817 and asqrt[20] n12008 ; n12009
g11818 nor n11458 n11467 ; n12010
g11819 and asqrt[20] n12010 ; n12011
g11820 nor n11465 n12011 ; n12012
g11821 nor n12009 n12012 ; n12013
g11822 nor asqrt[33] n11994 ; n12014
g11823 and n12004_not n12014 ; n12015
g11824 nor n12013 n12015 ; n12016
g11825 nor n12006 n12016 ; n12017
g11826 and asqrt[34] n12017_not ; n12018
g11827 and n11477 n11479_not ; n12019
g11828 and n11470_not n12019 ; n12020
g11829 and asqrt[20] n12020 ; n12021
g11830 nor n11470 n11479 ; n12022
g11831 and asqrt[20] n12022 ; n12023
g11832 nor n11477 n12023 ; n12024
g11833 nor n12021 n12024 ; n12025
g11834 nor asqrt[34] n12006 ; n12026
g11835 and n12016_not n12026 ; n12027
g11836 nor n12025 n12027 ; n12028
g11837 nor n12018 n12028 ; n12029
g11838 and asqrt[35] n12029_not ; n12030
g11839 and n11482_not n11489 ; n12031
g11840 and n11491_not n12031 ; n12032
g11841 and asqrt[20] n12032 ; n12033
g11842 nor n11482 n11491 ; n12034
g11843 and asqrt[20] n12034 ; n12035
g11844 nor n11489 n12035 ; n12036
g11845 nor n12033 n12036 ; n12037
g11846 nor asqrt[35] n12018 ; n12038
g11847 and n12028_not n12038 ; n12039
g11848 nor n12037 n12039 ; n12040
g11849 nor n12030 n12040 ; n12041
g11850 and asqrt[36] n12041_not ; n12042
g11851 and n11501 n11503_not ; n12043
g11852 and n11494_not n12043 ; n12044
g11853 and asqrt[20] n12044 ; n12045
g11854 nor n11494 n11503 ; n12046
g11855 and asqrt[20] n12046 ; n12047
g11856 nor n11501 n12047 ; n12048
g11857 nor n12045 n12048 ; n12049
g11858 nor asqrt[36] n12030 ; n12050
g11859 and n12040_not n12050 ; n12051
g11860 nor n12049 n12051 ; n12052
g11861 nor n12042 n12052 ; n12053
g11862 and asqrt[37] n12053_not ; n12054
g11863 and n11506_not n11513 ; n12055
g11864 and n11515_not n12055 ; n12056
g11865 and asqrt[20] n12056 ; n12057
g11866 nor n11506 n11515 ; n12058
g11867 and asqrt[20] n12058 ; n12059
g11868 nor n11513 n12059 ; n12060
g11869 nor n12057 n12060 ; n12061
g11870 nor asqrt[37] n12042 ; n12062
g11871 and n12052_not n12062 ; n12063
g11872 nor n12061 n12063 ; n12064
g11873 nor n12054 n12064 ; n12065
g11874 and asqrt[38] n12065_not ; n12066
g11875 and n11525 n11527_not ; n12067
g11876 and n11518_not n12067 ; n12068
g11877 and asqrt[20] n12068 ; n12069
g11878 nor n11518 n11527 ; n12070
g11879 and asqrt[20] n12070 ; n12071
g11880 nor n11525 n12071 ; n12072
g11881 nor n12069 n12072 ; n12073
g11882 nor asqrt[38] n12054 ; n12074
g11883 and n12064_not n12074 ; n12075
g11884 nor n12073 n12075 ; n12076
g11885 nor n12066 n12076 ; n12077
g11886 and asqrt[39] n12077_not ; n12078
g11887 and n11530_not n11537 ; n12079
g11888 and n11539_not n12079 ; n12080
g11889 and asqrt[20] n12080 ; n12081
g11890 nor n11530 n11539 ; n12082
g11891 and asqrt[20] n12082 ; n12083
g11892 nor n11537 n12083 ; n12084
g11893 nor n12081 n12084 ; n12085
g11894 nor asqrt[39] n12066 ; n12086
g11895 and n12076_not n12086 ; n12087
g11896 nor n12085 n12087 ; n12088
g11897 nor n12078 n12088 ; n12089
g11898 and asqrt[40] n12089_not ; n12090
g11899 and n11549 n11551_not ; n12091
g11900 and n11542_not n12091 ; n12092
g11901 and asqrt[20] n12092 ; n12093
g11902 nor n11542 n11551 ; n12094
g11903 and asqrt[20] n12094 ; n12095
g11904 nor n11549 n12095 ; n12096
g11905 nor n12093 n12096 ; n12097
g11906 nor asqrt[40] n12078 ; n12098
g11907 and n12088_not n12098 ; n12099
g11908 nor n12097 n12099 ; n12100
g11909 nor n12090 n12100 ; n12101
g11910 and asqrt[41] n12101_not ; n12102
g11911 and n11554_not n11561 ; n12103
g11912 and n11563_not n12103 ; n12104
g11913 and asqrt[20] n12104 ; n12105
g11914 nor n11554 n11563 ; n12106
g11915 and asqrt[20] n12106 ; n12107
g11916 nor n11561 n12107 ; n12108
g11917 nor n12105 n12108 ; n12109
g11918 nor asqrt[41] n12090 ; n12110
g11919 and n12100_not n12110 ; n12111
g11920 nor n12109 n12111 ; n12112
g11921 nor n12102 n12112 ; n12113
g11922 and asqrt[42] n12113_not ; n12114
g11923 and n11573 n11575_not ; n12115
g11924 and n11566_not n12115 ; n12116
g11925 and asqrt[20] n12116 ; n12117
g11926 nor n11566 n11575 ; n12118
g11927 and asqrt[20] n12118 ; n12119
g11928 nor n11573 n12119 ; n12120
g11929 nor n12117 n12120 ; n12121
g11930 nor asqrt[42] n12102 ; n12122
g11931 and n12112_not n12122 ; n12123
g11932 nor n12121 n12123 ; n12124
g11933 nor n12114 n12124 ; n12125
g11934 and asqrt[43] n12125_not ; n12126
g11935 and n11578_not n11585 ; n12127
g11936 and n11587_not n12127 ; n12128
g11937 and asqrt[20] n12128 ; n12129
g11938 nor n11578 n11587 ; n12130
g11939 and asqrt[20] n12130 ; n12131
g11940 nor n11585 n12131 ; n12132
g11941 nor n12129 n12132 ; n12133
g11942 nor asqrt[43] n12114 ; n12134
g11943 and n12124_not n12134 ; n12135
g11944 nor n12133 n12135 ; n12136
g11945 nor n12126 n12136 ; n12137
g11946 and asqrt[44] n12137_not ; n12138
g11947 and n11597 n11599_not ; n12139
g11948 and n11590_not n12139 ; n12140
g11949 and asqrt[20] n12140 ; n12141
g11950 nor n11590 n11599 ; n12142
g11951 and asqrt[20] n12142 ; n12143
g11952 nor n11597 n12143 ; n12144
g11953 nor n12141 n12144 ; n12145
g11954 nor asqrt[44] n12126 ; n12146
g11955 and n12136_not n12146 ; n12147
g11956 nor n12145 n12147 ; n12148
g11957 nor n12138 n12148 ; n12149
g11958 and asqrt[45] n12149_not ; n12150
g11959 nor asqrt[45] n12138 ; n12151
g11960 and n12148_not n12151 ; n12152
g11961 and n11602_not n11611 ; n12153
g11962 and n11604_not n12153 ; n12154
g11963 and asqrt[20] n12154 ; n12155
g11964 nor n11602 n11604 ; n12156
g11965 and asqrt[20] n12156 ; n12157
g11966 nor n11611 n12157 ; n12158
g11967 nor n12155 n12158 ; n12159
g11968 nor n12152 n12159 ; n12160
g11969 nor n12150 n12160 ; n12161
g11970 and asqrt[46] n12161_not ; n12162
g11971 and n11621 n11623_not ; n12163
g11972 and n11614_not n12163 ; n12164
g11973 and asqrt[20] n12164 ; n12165
g11974 nor n11614 n11623 ; n12166
g11975 and asqrt[20] n12166 ; n12167
g11976 nor n11621 n12167 ; n12168
g11977 nor n12165 n12168 ; n12169
g11978 nor asqrt[46] n12150 ; n12170
g11979 and n12160_not n12170 ; n12171
g11980 nor n12169 n12171 ; n12172
g11981 nor n12162 n12172 ; n12173
g11982 and asqrt[47] n12173_not ; n12174
g11983 and n11626_not n11633 ; n12175
g11984 and n11635_not n12175 ; n12176
g11985 and asqrt[20] n12176 ; n12177
g11986 nor n11626 n11635 ; n12178
g11987 and asqrt[20] n12178 ; n12179
g11988 nor n11633 n12179 ; n12180
g11989 nor n12177 n12180 ; n12181
g11990 nor asqrt[47] n12162 ; n12182
g11991 and n12172_not n12182 ; n12183
g11992 nor n12181 n12183 ; n12184
g11993 nor n12174 n12184 ; n12185
g11994 and asqrt[48] n12185_not ; n12186
g11995 and n11645 n11647_not ; n12187
g11996 and n11638_not n12187 ; n12188
g11997 and asqrt[20] n12188 ; n12189
g11998 nor n11638 n11647 ; n12190
g11999 and asqrt[20] n12190 ; n12191
g12000 nor n11645 n12191 ; n12192
g12001 nor n12189 n12192 ; n12193
g12002 nor asqrt[48] n12174 ; n12194
g12003 and n12184_not n12194 ; n12195
g12004 nor n12193 n12195 ; n12196
g12005 nor n12186 n12196 ; n12197
g12006 and asqrt[49] n12197_not ; n12198
g12007 and n11650_not n11657 ; n12199
g12008 and n11659_not n12199 ; n12200
g12009 and asqrt[20] n12200 ; n12201
g12010 nor n11650 n11659 ; n12202
g12011 and asqrt[20] n12202 ; n12203
g12012 nor n11657 n12203 ; n12204
g12013 nor n12201 n12204 ; n12205
g12014 nor asqrt[49] n12186 ; n12206
g12015 and n12196_not n12206 ; n12207
g12016 nor n12205 n12207 ; n12208
g12017 nor n12198 n12208 ; n12209
g12018 and asqrt[50] n12209_not ; n12210
g12019 and n11669 n11671_not ; n12211
g12020 and n11662_not n12211 ; n12212
g12021 and asqrt[20] n12212 ; n12213
g12022 nor n11662 n11671 ; n12214
g12023 and asqrt[20] n12214 ; n12215
g12024 nor n11669 n12215 ; n12216
g12025 nor n12213 n12216 ; n12217
g12026 nor asqrt[50] n12198 ; n12218
g12027 and n12208_not n12218 ; n12219
g12028 nor n12217 n12219 ; n12220
g12029 nor n12210 n12220 ; n12221
g12030 and asqrt[51] n12221_not ; n12222
g12031 and n11674_not n11681 ; n12223
g12032 and n11683_not n12223 ; n12224
g12033 and asqrt[20] n12224 ; n12225
g12034 nor n11674 n11683 ; n12226
g12035 and asqrt[20] n12226 ; n12227
g12036 nor n11681 n12227 ; n12228
g12037 nor n12225 n12228 ; n12229
g12038 nor asqrt[51] n12210 ; n12230
g12039 and n12220_not n12230 ; n12231
g12040 nor n12229 n12231 ; n12232
g12041 nor n12222 n12232 ; n12233
g12042 and asqrt[52] n12233_not ; n12234
g12043 and n11693 n11695_not ; n12235
g12044 and n11686_not n12235 ; n12236
g12045 and asqrt[20] n12236 ; n12237
g12046 nor n11686 n11695 ; n12238
g12047 and asqrt[20] n12238 ; n12239
g12048 nor n11693 n12239 ; n12240
g12049 nor n12237 n12240 ; n12241
g12050 nor asqrt[52] n12222 ; n12242
g12051 and n12232_not n12242 ; n12243
g12052 nor n12241 n12243 ; n12244
g12053 nor n12234 n12244 ; n12245
g12054 and asqrt[53] n12245_not ; n12246
g12055 and n11698_not n11705 ; n12247
g12056 and n11707_not n12247 ; n12248
g12057 and asqrt[20] n12248 ; n12249
g12058 nor n11698 n11707 ; n12250
g12059 and asqrt[20] n12250 ; n12251
g12060 nor n11705 n12251 ; n12252
g12061 nor n12249 n12252 ; n12253
g12062 nor asqrt[53] n12234 ; n12254
g12063 and n12244_not n12254 ; n12255
g12064 nor n12253 n12255 ; n12256
g12065 nor n12246 n12256 ; n12257
g12066 and asqrt[54] n12257_not ; n12258
g12067 and n11717 n11719_not ; n12259
g12068 and n11710_not n12259 ; n12260
g12069 and asqrt[20] n12260 ; n12261
g12070 nor n11710 n11719 ; n12262
g12071 and asqrt[20] n12262 ; n12263
g12072 nor n11717 n12263 ; n12264
g12073 nor n12261 n12264 ; n12265
g12074 nor asqrt[54] n12246 ; n12266
g12075 and n12256_not n12266 ; n12267
g12076 nor n12265 n12267 ; n12268
g12077 nor n12258 n12268 ; n12269
g12078 and asqrt[55] n12269_not ; n12270
g12079 and n11722_not n11729 ; n12271
g12080 and n11731_not n12271 ; n12272
g12081 and asqrt[20] n12272 ; n12273
g12082 nor n11722 n11731 ; n12274
g12083 and asqrt[20] n12274 ; n12275
g12084 nor n11729 n12275 ; n12276
g12085 nor n12273 n12276 ; n12277
g12086 nor asqrt[55] n12258 ; n12278
g12087 and n12268_not n12278 ; n12279
g12088 nor n12277 n12279 ; n12280
g12089 nor n12270 n12280 ; n12281
g12090 and asqrt[56] n12281_not ; n12282
g12091 and n11741 n11743_not ; n12283
g12092 and n11734_not n12283 ; n12284
g12093 and asqrt[20] n12284 ; n12285
g12094 nor n11734 n11743 ; n12286
g12095 and asqrt[20] n12286 ; n12287
g12096 nor n11741 n12287 ; n12288
g12097 nor n12285 n12288 ; n12289
g12098 nor asqrt[56] n12270 ; n12290
g12099 and n12280_not n12290 ; n12291
g12100 nor n12289 n12291 ; n12292
g12101 nor n12282 n12292 ; n12293
g12102 and asqrt[57] n12293_not ; n12294
g12103 and n11746_not n11753 ; n12295
g12104 and n11755_not n12295 ; n12296
g12105 and asqrt[20] n12296 ; n12297
g12106 nor n11746 n11755 ; n12298
g12107 and asqrt[20] n12298 ; n12299
g12108 nor n11753 n12299 ; n12300
g12109 nor n12297 n12300 ; n12301
g12110 nor asqrt[57] n12282 ; n12302
g12111 and n12292_not n12302 ; n12303
g12112 nor n12301 n12303 ; n12304
g12113 nor n12294 n12304 ; n12305
g12114 and asqrt[58] n12305_not ; n12306
g12115 and n11765 n11767_not ; n12307
g12116 and n11758_not n12307 ; n12308
g12117 and asqrt[20] n12308 ; n12309
g12118 nor n11758 n11767 ; n12310
g12119 and asqrt[20] n12310 ; n12311
g12120 nor n11765 n12311 ; n12312
g12121 nor n12309 n12312 ; n12313
g12122 nor asqrt[58] n12294 ; n12314
g12123 and n12304_not n12314 ; n12315
g12124 nor n12313 n12315 ; n12316
g12125 nor n12306 n12316 ; n12317
g12126 and asqrt[59] n12317_not ; n12318
g12127 and n11770_not n11777 ; n12319
g12128 and n11779_not n12319 ; n12320
g12129 and asqrt[20] n12320 ; n12321
g12130 nor n11770 n11779 ; n12322
g12131 and asqrt[20] n12322 ; n12323
g12132 nor n11777 n12323 ; n12324
g12133 nor n12321 n12324 ; n12325
g12134 nor asqrt[59] n12306 ; n12326
g12135 and n12316_not n12326 ; n12327
g12136 nor n12325 n12327 ; n12328
g12137 nor n12318 n12328 ; n12329
g12138 and asqrt[60] n12329_not ; n12330
g12139 and n11789 n11791_not ; n12331
g12140 and n11782_not n12331 ; n12332
g12141 and asqrt[20] n12332 ; n12333
g12142 nor n11782 n11791 ; n12334
g12143 and asqrt[20] n12334 ; n12335
g12144 nor n11789 n12335 ; n12336
g12145 nor n12333 n12336 ; n12337
g12146 nor asqrt[60] n12318 ; n12338
g12147 and n12328_not n12338 ; n12339
g12148 nor n12337 n12339 ; n12340
g12149 nor n12330 n12340 ; n12341
g12150 and asqrt[61] n12341_not ; n12342
g12151 and n11794_not n11801 ; n12343
g12152 and n11803_not n12343 ; n12344
g12153 and asqrt[20] n12344 ; n12345
g12154 nor n11794 n11803 ; n12346
g12155 and asqrt[20] n12346 ; n12347
g12156 nor n11801 n12347 ; n12348
g12157 nor n12345 n12348 ; n12349
g12158 nor asqrt[61] n12330 ; n12350
g12159 and n12340_not n12350 ; n12351
g12160 nor n12349 n12351 ; n12352
g12161 nor n12342 n12352 ; n12353
g12162 and asqrt[62] n12353_not ; n12354
g12163 and n11813 n11815_not ; n12355
g12164 and n11806_not n12355 ; n12356
g12165 and asqrt[20] n12356 ; n12357
g12166 nor n11806 n11815 ; n12358
g12167 and asqrt[20] n12358 ; n12359
g12168 nor n11813 n12359 ; n12360
g12169 nor n12357 n12360 ; n12361
g12170 nor asqrt[62] n12342 ; n12362
g12171 and n12352_not n12362 ; n12363
g12172 nor n12361 n12363 ; n12364
g12173 nor n12354 n12364 ; n12365
g12174 and n11818_not n11825 ; n12366
g12175 and n11827_not n12366 ; n12367
g12176 and asqrt[20] n12367 ; n12368
g12177 nor n11818 n11827 ; n12369
g12178 and asqrt[20] n12369 ; n12370
g12179 nor n11825 n12370 ; n12371
g12180 nor n12368 n12371 ; n12372
g12181 nor n11829 n11836 ; n12373
g12182 and asqrt[20] n12373 ; n12374
g12183 nor n11844 n12374 ; n12375
g12184 and n12372_not n12375 ; n12376
g12185 and n12365_not n12376 ; n12377
g12186 nor asqrt[63] n12377 ; n12378
g12187 and n12354_not n12372 ; n12379
g12188 and n12364_not n12379 ; n12380
g12189 and n11836_not asqrt[20] ; n12381
g12190 and n11829 n12381_not ; n12382
g12191 and asqrt[63] n12373_not ; n12383
g12192 and n12382_not n12383 ; n12384
g12193 nor n11832 n11853 ; n12385
g12194 and n11835_not n12385 ; n12386
g12195 and n11848_not n12386 ; n12387
g12196 and n11844_not n12387 ; n12388
g12197 and n11842_not n12388 ; n12389
g12198 nor n12384 n12389 ; n12390
g12199 and n12380_not n12390 ; n12391
g12200 nand n12378_not n12391 ; asqrt[19]
g12201 and a[38] asqrt[19] ; n12393
g12202 nor a[36] a[37] ; n12394
g12203 and a[38]_not n12394 ; n12395
g12204 nor n12393 n12395 ; n12396
g12205 and asqrt[20] n12396_not ; n12397
g12206 nor n11853 n12395 ; n12398
g12207 and n11848_not n12398 ; n12399
g12208 and n11844_not n12399 ; n12400
g12209 and n11842_not n12400 ; n12401
g12210 and n12393_not n12401 ; n12402
g12211 and a[38]_not asqrt[19] ; n12403
g12212 and a[39] n12403_not ; n12404
g12213 and n11858 asqrt[19] ; n12405
g12214 nor n12404 n12405 ; n12406
g12215 and n12402_not n12406 ; n12407
g12216 nor n12397 n12407 ; n12408
g12217 and asqrt[21] n12408_not ; n12409
g12218 nor asqrt[21] n12397 ; n12410
g12219 and n12407_not n12410 ; n12411
g12220 and asqrt[20] n12389_not ; n12412
g12221 and n12384_not n12412 ; n12413
g12222 and n12380_not n12413 ; n12414
g12223 and n12378_not n12414 ; n12415
g12224 nor n12405 n12415 ; n12416
g12225 and a[40] n12416_not ; n12417
g12226 nor a[40] n12415 ; n12418
g12227 and n12405_not n12418 ; n12419
g12228 nor n12417 n12419 ; n12420
g12229 nor n12411 n12420 ; n12421
g12230 nor n12409 n12421 ; n12422
g12231 and asqrt[22] n12422_not ; n12423
g12232 nor n11861 n11866 ; n12424
g12233 and n11870_not n12424 ; n12425
g12234 and asqrt[19] n12425 ; n12426
g12235 and asqrt[19] n12424 ; n12427
g12236 and n11870 n12427_not ; n12428
g12237 nor n12426 n12428 ; n12429
g12238 nor asqrt[22] n12409 ; n12430
g12239 and n12421_not n12430 ; n12431
g12240 nor n12429 n12431 ; n12432
g12241 nor n12423 n12432 ; n12433
g12242 and asqrt[23] n12433_not ; n12434
g12243 and n11875_not n11884 ; n12435
g12244 and n11873_not n12435 ; n12436
g12245 and asqrt[19] n12436 ; n12437
g12246 nor n11873 n11875 ; n12438
g12247 and asqrt[19] n12438 ; n12439
g12248 nor n11884 n12439 ; n12440
g12249 nor n12437 n12440 ; n12441
g12250 nor asqrt[23] n12423 ; n12442
g12251 and n12432_not n12442 ; n12443
g12252 nor n12441 n12443 ; n12444
g12253 nor n12434 n12444 ; n12445
g12254 and asqrt[24] n12445_not ; n12446
g12255 and n11887_not n11893 ; n12447
g12256 and n11895_not n12447 ; n12448
g12257 and asqrt[19] n12448 ; n12449
g12258 nor n11887 n11895 ; n12450
g12259 and asqrt[19] n12450 ; n12451
g12260 nor n11893 n12451 ; n12452
g12261 nor n12449 n12452 ; n12453
g12262 nor asqrt[24] n12434 ; n12454
g12263 and n12444_not n12454 ; n12455
g12264 nor n12453 n12455 ; n12456
g12265 nor n12446 n12456 ; n12457
g12266 and asqrt[25] n12457_not ; n12458
g12267 and n11905 n11907_not ; n12459
g12268 and n11898_not n12459 ; n12460
g12269 and asqrt[19] n12460 ; n12461
g12270 nor n11898 n11907 ; n12462
g12271 and asqrt[19] n12462 ; n12463
g12272 nor n11905 n12463 ; n12464
g12273 nor n12461 n12464 ; n12465
g12274 nor asqrt[25] n12446 ; n12466
g12275 and n12456_not n12466 ; n12467
g12276 nor n12465 n12467 ; n12468
g12277 nor n12458 n12468 ; n12469
g12278 and asqrt[26] n12469_not ; n12470
g12279 and n11910_not n11917 ; n12471
g12280 and n11919_not n12471 ; n12472
g12281 and asqrt[19] n12472 ; n12473
g12282 nor n11910 n11919 ; n12474
g12283 and asqrt[19] n12474 ; n12475
g12284 nor n11917 n12475 ; n12476
g12285 nor n12473 n12476 ; n12477
g12286 nor asqrt[26] n12458 ; n12478
g12287 and n12468_not n12478 ; n12479
g12288 nor n12477 n12479 ; n12480
g12289 nor n12470 n12480 ; n12481
g12290 and asqrt[27] n12481_not ; n12482
g12291 and n11929 n11931_not ; n12483
g12292 and n11922_not n12483 ; n12484
g12293 and asqrt[19] n12484 ; n12485
g12294 nor n11922 n11931 ; n12486
g12295 and asqrt[19] n12486 ; n12487
g12296 nor n11929 n12487 ; n12488
g12297 nor n12485 n12488 ; n12489
g12298 nor asqrt[27] n12470 ; n12490
g12299 and n12480_not n12490 ; n12491
g12300 nor n12489 n12491 ; n12492
g12301 nor n12482 n12492 ; n12493
g12302 and asqrt[28] n12493_not ; n12494
g12303 and n11934_not n11941 ; n12495
g12304 and n11943_not n12495 ; n12496
g12305 and asqrt[19] n12496 ; n12497
g12306 nor n11934 n11943 ; n12498
g12307 and asqrt[19] n12498 ; n12499
g12308 nor n11941 n12499 ; n12500
g12309 nor n12497 n12500 ; n12501
g12310 nor asqrt[28] n12482 ; n12502
g12311 and n12492_not n12502 ; n12503
g12312 nor n12501 n12503 ; n12504
g12313 nor n12494 n12504 ; n12505
g12314 and asqrt[29] n12505_not ; n12506
g12315 and n11953 n11955_not ; n12507
g12316 and n11946_not n12507 ; n12508
g12317 and asqrt[19] n12508 ; n12509
g12318 nor n11946 n11955 ; n12510
g12319 and asqrt[19] n12510 ; n12511
g12320 nor n11953 n12511 ; n12512
g12321 nor n12509 n12512 ; n12513
g12322 nor asqrt[29] n12494 ; n12514
g12323 and n12504_not n12514 ; n12515
g12324 nor n12513 n12515 ; n12516
g12325 nor n12506 n12516 ; n12517
g12326 and asqrt[30] n12517_not ; n12518
g12327 and n11958_not n11965 ; n12519
g12328 and n11967_not n12519 ; n12520
g12329 and asqrt[19] n12520 ; n12521
g12330 nor n11958 n11967 ; n12522
g12331 and asqrt[19] n12522 ; n12523
g12332 nor n11965 n12523 ; n12524
g12333 nor n12521 n12524 ; n12525
g12334 nor asqrt[30] n12506 ; n12526
g12335 and n12516_not n12526 ; n12527
g12336 nor n12525 n12527 ; n12528
g12337 nor n12518 n12528 ; n12529
g12338 and asqrt[31] n12529_not ; n12530
g12339 and n11977 n11979_not ; n12531
g12340 and n11970_not n12531 ; n12532
g12341 and asqrt[19] n12532 ; n12533
g12342 nor n11970 n11979 ; n12534
g12343 and asqrt[19] n12534 ; n12535
g12344 nor n11977 n12535 ; n12536
g12345 nor n12533 n12536 ; n12537
g12346 nor asqrt[31] n12518 ; n12538
g12347 and n12528_not n12538 ; n12539
g12348 nor n12537 n12539 ; n12540
g12349 nor n12530 n12540 ; n12541
g12350 and asqrt[32] n12541_not ; n12542
g12351 and n11982_not n11989 ; n12543
g12352 and n11991_not n12543 ; n12544
g12353 and asqrt[19] n12544 ; n12545
g12354 nor n11982 n11991 ; n12546
g12355 and asqrt[19] n12546 ; n12547
g12356 nor n11989 n12547 ; n12548
g12357 nor n12545 n12548 ; n12549
g12358 nor asqrt[32] n12530 ; n12550
g12359 and n12540_not n12550 ; n12551
g12360 nor n12549 n12551 ; n12552
g12361 nor n12542 n12552 ; n12553
g12362 and asqrt[33] n12553_not ; n12554
g12363 and n12001 n12003_not ; n12555
g12364 and n11994_not n12555 ; n12556
g12365 and asqrt[19] n12556 ; n12557
g12366 nor n11994 n12003 ; n12558
g12367 and asqrt[19] n12558 ; n12559
g12368 nor n12001 n12559 ; n12560
g12369 nor n12557 n12560 ; n12561
g12370 nor asqrt[33] n12542 ; n12562
g12371 and n12552_not n12562 ; n12563
g12372 nor n12561 n12563 ; n12564
g12373 nor n12554 n12564 ; n12565
g12374 and asqrt[34] n12565_not ; n12566
g12375 and n12006_not n12013 ; n12567
g12376 and n12015_not n12567 ; n12568
g12377 and asqrt[19] n12568 ; n12569
g12378 nor n12006 n12015 ; n12570
g12379 and asqrt[19] n12570 ; n12571
g12380 nor n12013 n12571 ; n12572
g12381 nor n12569 n12572 ; n12573
g12382 nor asqrt[34] n12554 ; n12574
g12383 and n12564_not n12574 ; n12575
g12384 nor n12573 n12575 ; n12576
g12385 nor n12566 n12576 ; n12577
g12386 and asqrt[35] n12577_not ; n12578
g12387 and n12025 n12027_not ; n12579
g12388 and n12018_not n12579 ; n12580
g12389 and asqrt[19] n12580 ; n12581
g12390 nor n12018 n12027 ; n12582
g12391 and asqrt[19] n12582 ; n12583
g12392 nor n12025 n12583 ; n12584
g12393 nor n12581 n12584 ; n12585
g12394 nor asqrt[35] n12566 ; n12586
g12395 and n12576_not n12586 ; n12587
g12396 nor n12585 n12587 ; n12588
g12397 nor n12578 n12588 ; n12589
g12398 and asqrt[36] n12589_not ; n12590
g12399 and n12030_not n12037 ; n12591
g12400 and n12039_not n12591 ; n12592
g12401 and asqrt[19] n12592 ; n12593
g12402 nor n12030 n12039 ; n12594
g12403 and asqrt[19] n12594 ; n12595
g12404 nor n12037 n12595 ; n12596
g12405 nor n12593 n12596 ; n12597
g12406 nor asqrt[36] n12578 ; n12598
g12407 and n12588_not n12598 ; n12599
g12408 nor n12597 n12599 ; n12600
g12409 nor n12590 n12600 ; n12601
g12410 and asqrt[37] n12601_not ; n12602
g12411 and n12049 n12051_not ; n12603
g12412 and n12042_not n12603 ; n12604
g12413 and asqrt[19] n12604 ; n12605
g12414 nor n12042 n12051 ; n12606
g12415 and asqrt[19] n12606 ; n12607
g12416 nor n12049 n12607 ; n12608
g12417 nor n12605 n12608 ; n12609
g12418 nor asqrt[37] n12590 ; n12610
g12419 and n12600_not n12610 ; n12611
g12420 nor n12609 n12611 ; n12612
g12421 nor n12602 n12612 ; n12613
g12422 and asqrt[38] n12613_not ; n12614
g12423 and n12054_not n12061 ; n12615
g12424 and n12063_not n12615 ; n12616
g12425 and asqrt[19] n12616 ; n12617
g12426 nor n12054 n12063 ; n12618
g12427 and asqrt[19] n12618 ; n12619
g12428 nor n12061 n12619 ; n12620
g12429 nor n12617 n12620 ; n12621
g12430 nor asqrt[38] n12602 ; n12622
g12431 and n12612_not n12622 ; n12623
g12432 nor n12621 n12623 ; n12624
g12433 nor n12614 n12624 ; n12625
g12434 and asqrt[39] n12625_not ; n12626
g12435 and n12073 n12075_not ; n12627
g12436 and n12066_not n12627 ; n12628
g12437 and asqrt[19] n12628 ; n12629
g12438 nor n12066 n12075 ; n12630
g12439 and asqrt[19] n12630 ; n12631
g12440 nor n12073 n12631 ; n12632
g12441 nor n12629 n12632 ; n12633
g12442 nor asqrt[39] n12614 ; n12634
g12443 and n12624_not n12634 ; n12635
g12444 nor n12633 n12635 ; n12636
g12445 nor n12626 n12636 ; n12637
g12446 and asqrt[40] n12637_not ; n12638
g12447 and n12078_not n12085 ; n12639
g12448 and n12087_not n12639 ; n12640
g12449 and asqrt[19] n12640 ; n12641
g12450 nor n12078 n12087 ; n12642
g12451 and asqrt[19] n12642 ; n12643
g12452 nor n12085 n12643 ; n12644
g12453 nor n12641 n12644 ; n12645
g12454 nor asqrt[40] n12626 ; n12646
g12455 and n12636_not n12646 ; n12647
g12456 nor n12645 n12647 ; n12648
g12457 nor n12638 n12648 ; n12649
g12458 and asqrt[41] n12649_not ; n12650
g12459 and n12097 n12099_not ; n12651
g12460 and n12090_not n12651 ; n12652
g12461 and asqrt[19] n12652 ; n12653
g12462 nor n12090 n12099 ; n12654
g12463 and asqrt[19] n12654 ; n12655
g12464 nor n12097 n12655 ; n12656
g12465 nor n12653 n12656 ; n12657
g12466 nor asqrt[41] n12638 ; n12658
g12467 and n12648_not n12658 ; n12659
g12468 nor n12657 n12659 ; n12660
g12469 nor n12650 n12660 ; n12661
g12470 and asqrt[42] n12661_not ; n12662
g12471 and n12102_not n12109 ; n12663
g12472 and n12111_not n12663 ; n12664
g12473 and asqrt[19] n12664 ; n12665
g12474 nor n12102 n12111 ; n12666
g12475 and asqrt[19] n12666 ; n12667
g12476 nor n12109 n12667 ; n12668
g12477 nor n12665 n12668 ; n12669
g12478 nor asqrt[42] n12650 ; n12670
g12479 and n12660_not n12670 ; n12671
g12480 nor n12669 n12671 ; n12672
g12481 nor n12662 n12672 ; n12673
g12482 and asqrt[43] n12673_not ; n12674
g12483 and n12121 n12123_not ; n12675
g12484 and n12114_not n12675 ; n12676
g12485 and asqrt[19] n12676 ; n12677
g12486 nor n12114 n12123 ; n12678
g12487 and asqrt[19] n12678 ; n12679
g12488 nor n12121 n12679 ; n12680
g12489 nor n12677 n12680 ; n12681
g12490 nor asqrt[43] n12662 ; n12682
g12491 and n12672_not n12682 ; n12683
g12492 nor n12681 n12683 ; n12684
g12493 nor n12674 n12684 ; n12685
g12494 and asqrt[44] n12685_not ; n12686
g12495 and n12126_not n12133 ; n12687
g12496 and n12135_not n12687 ; n12688
g12497 and asqrt[19] n12688 ; n12689
g12498 nor n12126 n12135 ; n12690
g12499 and asqrt[19] n12690 ; n12691
g12500 nor n12133 n12691 ; n12692
g12501 nor n12689 n12692 ; n12693
g12502 nor asqrt[44] n12674 ; n12694
g12503 and n12684_not n12694 ; n12695
g12504 nor n12693 n12695 ; n12696
g12505 nor n12686 n12696 ; n12697
g12506 and asqrt[45] n12697_not ; n12698
g12507 and n12145 n12147_not ; n12699
g12508 and n12138_not n12699 ; n12700
g12509 and asqrt[19] n12700 ; n12701
g12510 nor n12138 n12147 ; n12702
g12511 and asqrt[19] n12702 ; n12703
g12512 nor n12145 n12703 ; n12704
g12513 nor n12701 n12704 ; n12705
g12514 nor asqrt[45] n12686 ; n12706
g12515 and n12696_not n12706 ; n12707
g12516 nor n12705 n12707 ; n12708
g12517 nor n12698 n12708 ; n12709
g12518 and asqrt[46] n12709_not ; n12710
g12519 nor asqrt[46] n12698 ; n12711
g12520 and n12708_not n12711 ; n12712
g12521 and n12150_not n12159 ; n12713
g12522 and n12152_not n12713 ; n12714
g12523 and asqrt[19] n12714 ; n12715
g12524 nor n12150 n12152 ; n12716
g12525 and asqrt[19] n12716 ; n12717
g12526 nor n12159 n12717 ; n12718
g12527 nor n12715 n12718 ; n12719
g12528 nor n12712 n12719 ; n12720
g12529 nor n12710 n12720 ; n12721
g12530 and asqrt[47] n12721_not ; n12722
g12531 and n12169 n12171_not ; n12723
g12532 and n12162_not n12723 ; n12724
g12533 and asqrt[19] n12724 ; n12725
g12534 nor n12162 n12171 ; n12726
g12535 and asqrt[19] n12726 ; n12727
g12536 nor n12169 n12727 ; n12728
g12537 nor n12725 n12728 ; n12729
g12538 nor asqrt[47] n12710 ; n12730
g12539 and n12720_not n12730 ; n12731
g12540 nor n12729 n12731 ; n12732
g12541 nor n12722 n12732 ; n12733
g12542 and asqrt[48] n12733_not ; n12734
g12543 and n12174_not n12181 ; n12735
g12544 and n12183_not n12735 ; n12736
g12545 and asqrt[19] n12736 ; n12737
g12546 nor n12174 n12183 ; n12738
g12547 and asqrt[19] n12738 ; n12739
g12548 nor n12181 n12739 ; n12740
g12549 nor n12737 n12740 ; n12741
g12550 nor asqrt[48] n12722 ; n12742
g12551 and n12732_not n12742 ; n12743
g12552 nor n12741 n12743 ; n12744
g12553 nor n12734 n12744 ; n12745
g12554 and asqrt[49] n12745_not ; n12746
g12555 and n12193 n12195_not ; n12747
g12556 and n12186_not n12747 ; n12748
g12557 and asqrt[19] n12748 ; n12749
g12558 nor n12186 n12195 ; n12750
g12559 and asqrt[19] n12750 ; n12751
g12560 nor n12193 n12751 ; n12752
g12561 nor n12749 n12752 ; n12753
g12562 nor asqrt[49] n12734 ; n12754
g12563 and n12744_not n12754 ; n12755
g12564 nor n12753 n12755 ; n12756
g12565 nor n12746 n12756 ; n12757
g12566 and asqrt[50] n12757_not ; n12758
g12567 and n12198_not n12205 ; n12759
g12568 and n12207_not n12759 ; n12760
g12569 and asqrt[19] n12760 ; n12761
g12570 nor n12198 n12207 ; n12762
g12571 and asqrt[19] n12762 ; n12763
g12572 nor n12205 n12763 ; n12764
g12573 nor n12761 n12764 ; n12765
g12574 nor asqrt[50] n12746 ; n12766
g12575 and n12756_not n12766 ; n12767
g12576 nor n12765 n12767 ; n12768
g12577 nor n12758 n12768 ; n12769
g12578 and asqrt[51] n12769_not ; n12770
g12579 and n12217 n12219_not ; n12771
g12580 and n12210_not n12771 ; n12772
g12581 and asqrt[19] n12772 ; n12773
g12582 nor n12210 n12219 ; n12774
g12583 and asqrt[19] n12774 ; n12775
g12584 nor n12217 n12775 ; n12776
g12585 nor n12773 n12776 ; n12777
g12586 nor asqrt[51] n12758 ; n12778
g12587 and n12768_not n12778 ; n12779
g12588 nor n12777 n12779 ; n12780
g12589 nor n12770 n12780 ; n12781
g12590 and asqrt[52] n12781_not ; n12782
g12591 and n12222_not n12229 ; n12783
g12592 and n12231_not n12783 ; n12784
g12593 and asqrt[19] n12784 ; n12785
g12594 nor n12222 n12231 ; n12786
g12595 and asqrt[19] n12786 ; n12787
g12596 nor n12229 n12787 ; n12788
g12597 nor n12785 n12788 ; n12789
g12598 nor asqrt[52] n12770 ; n12790
g12599 and n12780_not n12790 ; n12791
g12600 nor n12789 n12791 ; n12792
g12601 nor n12782 n12792 ; n12793
g12602 and asqrt[53] n12793_not ; n12794
g12603 and n12241 n12243_not ; n12795
g12604 and n12234_not n12795 ; n12796
g12605 and asqrt[19] n12796 ; n12797
g12606 nor n12234 n12243 ; n12798
g12607 and asqrt[19] n12798 ; n12799
g12608 nor n12241 n12799 ; n12800
g12609 nor n12797 n12800 ; n12801
g12610 nor asqrt[53] n12782 ; n12802
g12611 and n12792_not n12802 ; n12803
g12612 nor n12801 n12803 ; n12804
g12613 nor n12794 n12804 ; n12805
g12614 and asqrt[54] n12805_not ; n12806
g12615 and n12246_not n12253 ; n12807
g12616 and n12255_not n12807 ; n12808
g12617 and asqrt[19] n12808 ; n12809
g12618 nor n12246 n12255 ; n12810
g12619 and asqrt[19] n12810 ; n12811
g12620 nor n12253 n12811 ; n12812
g12621 nor n12809 n12812 ; n12813
g12622 nor asqrt[54] n12794 ; n12814
g12623 and n12804_not n12814 ; n12815
g12624 nor n12813 n12815 ; n12816
g12625 nor n12806 n12816 ; n12817
g12626 and asqrt[55] n12817_not ; n12818
g12627 and n12265 n12267_not ; n12819
g12628 and n12258_not n12819 ; n12820
g12629 and asqrt[19] n12820 ; n12821
g12630 nor n12258 n12267 ; n12822
g12631 and asqrt[19] n12822 ; n12823
g12632 nor n12265 n12823 ; n12824
g12633 nor n12821 n12824 ; n12825
g12634 nor asqrt[55] n12806 ; n12826
g12635 and n12816_not n12826 ; n12827
g12636 nor n12825 n12827 ; n12828
g12637 nor n12818 n12828 ; n12829
g12638 and asqrt[56] n12829_not ; n12830
g12639 and n12270_not n12277 ; n12831
g12640 and n12279_not n12831 ; n12832
g12641 and asqrt[19] n12832 ; n12833
g12642 nor n12270 n12279 ; n12834
g12643 and asqrt[19] n12834 ; n12835
g12644 nor n12277 n12835 ; n12836
g12645 nor n12833 n12836 ; n12837
g12646 nor asqrt[56] n12818 ; n12838
g12647 and n12828_not n12838 ; n12839
g12648 nor n12837 n12839 ; n12840
g12649 nor n12830 n12840 ; n12841
g12650 and asqrt[57] n12841_not ; n12842
g12651 and n12289 n12291_not ; n12843
g12652 and n12282_not n12843 ; n12844
g12653 and asqrt[19] n12844 ; n12845
g12654 nor n12282 n12291 ; n12846
g12655 and asqrt[19] n12846 ; n12847
g12656 nor n12289 n12847 ; n12848
g12657 nor n12845 n12848 ; n12849
g12658 nor asqrt[57] n12830 ; n12850
g12659 and n12840_not n12850 ; n12851
g12660 nor n12849 n12851 ; n12852
g12661 nor n12842 n12852 ; n12853
g12662 and asqrt[58] n12853_not ; n12854
g12663 and n12294_not n12301 ; n12855
g12664 and n12303_not n12855 ; n12856
g12665 and asqrt[19] n12856 ; n12857
g12666 nor n12294 n12303 ; n12858
g12667 and asqrt[19] n12858 ; n12859
g12668 nor n12301 n12859 ; n12860
g12669 nor n12857 n12860 ; n12861
g12670 nor asqrt[58] n12842 ; n12862
g12671 and n12852_not n12862 ; n12863
g12672 nor n12861 n12863 ; n12864
g12673 nor n12854 n12864 ; n12865
g12674 and asqrt[59] n12865_not ; n12866
g12675 and n12313 n12315_not ; n12867
g12676 and n12306_not n12867 ; n12868
g12677 and asqrt[19] n12868 ; n12869
g12678 nor n12306 n12315 ; n12870
g12679 and asqrt[19] n12870 ; n12871
g12680 nor n12313 n12871 ; n12872
g12681 nor n12869 n12872 ; n12873
g12682 nor asqrt[59] n12854 ; n12874
g12683 and n12864_not n12874 ; n12875
g12684 nor n12873 n12875 ; n12876
g12685 nor n12866 n12876 ; n12877
g12686 and asqrt[60] n12877_not ; n12878
g12687 and n12318_not n12325 ; n12879
g12688 and n12327_not n12879 ; n12880
g12689 and asqrt[19] n12880 ; n12881
g12690 nor n12318 n12327 ; n12882
g12691 and asqrt[19] n12882 ; n12883
g12692 nor n12325 n12883 ; n12884
g12693 nor n12881 n12884 ; n12885
g12694 nor asqrt[60] n12866 ; n12886
g12695 and n12876_not n12886 ; n12887
g12696 nor n12885 n12887 ; n12888
g12697 nor n12878 n12888 ; n12889
g12698 and asqrt[61] n12889_not ; n12890
g12699 and n12337 n12339_not ; n12891
g12700 and n12330_not n12891 ; n12892
g12701 and asqrt[19] n12892 ; n12893
g12702 nor n12330 n12339 ; n12894
g12703 and asqrt[19] n12894 ; n12895
g12704 nor n12337 n12895 ; n12896
g12705 nor n12893 n12896 ; n12897
g12706 nor asqrt[61] n12878 ; n12898
g12707 and n12888_not n12898 ; n12899
g12708 nor n12897 n12899 ; n12900
g12709 nor n12890 n12900 ; n12901
g12710 and asqrt[62] n12901_not ; n12902
g12711 and n12342_not n12349 ; n12903
g12712 and n12351_not n12903 ; n12904
g12713 and asqrt[19] n12904 ; n12905
g12714 nor n12342 n12351 ; n12906
g12715 and asqrt[19] n12906 ; n12907
g12716 nor n12349 n12907 ; n12908
g12717 nor n12905 n12908 ; n12909
g12718 nor asqrt[62] n12890 ; n12910
g12719 and n12900_not n12910 ; n12911
g12720 nor n12909 n12911 ; n12912
g12721 nor n12902 n12912 ; n12913
g12722 and n12361 n12363_not ; n12914
g12723 and n12354_not n12914 ; n12915
g12724 and asqrt[19] n12915 ; n12916
g12725 nor n12354 n12363 ; n12917
g12726 and asqrt[19] n12917 ; n12918
g12727 nor n12361 n12918 ; n12919
g12728 nor n12916 n12919 ; n12920
g12729 nor n12365 n12372 ; n12921
g12730 and asqrt[19] n12921 ; n12922
g12731 nor n12380 n12922 ; n12923
g12732 and n12920_not n12923 ; n12924
g12733 and n12913_not n12924 ; n12925
g12734 nor asqrt[63] n12925 ; n12926
g12735 and n12902_not n12920 ; n12927
g12736 and n12912_not n12927 ; n12928
g12737 and n12372_not asqrt[19] ; n12929
g12738 and n12365 n12929_not ; n12930
g12739 and asqrt[63] n12921_not ; n12931
g12740 and n12930_not n12931 ; n12932
g12741 nor n12368 n12389 ; n12933
g12742 and n12371_not n12933 ; n12934
g12743 and n12384_not n12934 ; n12935
g12744 and n12380_not n12935 ; n12936
g12745 and n12378_not n12936 ; n12937
g12746 nor n12932 n12937 ; n12938
g12747 and n12928_not n12938 ; n12939
g12748 nand n12926_not n12939 ; asqrt[18]
g12749 and a[36] asqrt[18] ; n12941
g12750 nor a[34] a[35] ; n12942
g12751 and a[36]_not n12942 ; n12943
g12752 nor n12941 n12943 ; n12944
g12753 and asqrt[19] n12944_not ; n12945
g12754 nor n12389 n12943 ; n12946
g12755 and n12384_not n12946 ; n12947
g12756 and n12380_not n12947 ; n12948
g12757 and n12378_not n12948 ; n12949
g12758 and n12941_not n12949 ; n12950
g12759 and a[36]_not asqrt[18] ; n12951
g12760 and a[37] n12951_not ; n12952
g12761 and n12394 asqrt[18] ; n12953
g12762 nor n12952 n12953 ; n12954
g12763 and n12950_not n12954 ; n12955
g12764 nor n12945 n12955 ; n12956
g12765 and asqrt[20] n12956_not ; n12957
g12766 nor asqrt[20] n12945 ; n12958
g12767 and n12955_not n12958 ; n12959
g12768 and asqrt[19] n12937_not ; n12960
g12769 and n12932_not n12960 ; n12961
g12770 and n12928_not n12961 ; n12962
g12771 and n12926_not n12962 ; n12963
g12772 nor n12953 n12963 ; n12964
g12773 and a[38] n12964_not ; n12965
g12774 nor a[38] n12963 ; n12966
g12775 and n12953_not n12966 ; n12967
g12776 nor n12965 n12967 ; n12968
g12777 nor n12959 n12968 ; n12969
g12778 nor n12957 n12969 ; n12970
g12779 and asqrt[21] n12970_not ; n12971
g12780 nor n12397 n12402 ; n12972
g12781 and n12406_not n12972 ; n12973
g12782 and asqrt[18] n12973 ; n12974
g12783 and asqrt[18] n12972 ; n12975
g12784 and n12406 n12975_not ; n12976
g12785 nor n12974 n12976 ; n12977
g12786 nor asqrt[21] n12957 ; n12978
g12787 and n12969_not n12978 ; n12979
g12788 nor n12977 n12979 ; n12980
g12789 nor n12971 n12980 ; n12981
g12790 and asqrt[22] n12981_not ; n12982
g12791 and n12411_not n12420 ; n12983
g12792 and n12409_not n12983 ; n12984
g12793 and asqrt[18] n12984 ; n12985
g12794 nor n12409 n12411 ; n12986
g12795 and asqrt[18] n12986 ; n12987
g12796 nor n12420 n12987 ; n12988
g12797 nor n12985 n12988 ; n12989
g12798 nor asqrt[22] n12971 ; n12990
g12799 and n12980_not n12990 ; n12991
g12800 nor n12989 n12991 ; n12992
g12801 nor n12982 n12992 ; n12993
g12802 and asqrt[23] n12993_not ; n12994
g12803 and n12423_not n12429 ; n12995
g12804 and n12431_not n12995 ; n12996
g12805 and asqrt[18] n12996 ; n12997
g12806 nor n12423 n12431 ; n12998
g12807 and asqrt[18] n12998 ; n12999
g12808 nor n12429 n12999 ; n13000
g12809 nor n12997 n13000 ; n13001
g12810 nor asqrt[23] n12982 ; n13002
g12811 and n12992_not n13002 ; n13003
g12812 nor n13001 n13003 ; n13004
g12813 nor n12994 n13004 ; n13005
g12814 and asqrt[24] n13005_not ; n13006
g12815 and n12441 n12443_not ; n13007
g12816 and n12434_not n13007 ; n13008
g12817 and asqrt[18] n13008 ; n13009
g12818 nor n12434 n12443 ; n13010
g12819 and asqrt[18] n13010 ; n13011
g12820 nor n12441 n13011 ; n13012
g12821 nor n13009 n13012 ; n13013
g12822 nor asqrt[24] n12994 ; n13014
g12823 and n13004_not n13014 ; n13015
g12824 nor n13013 n13015 ; n13016
g12825 nor n13006 n13016 ; n13017
g12826 and asqrt[25] n13017_not ; n13018
g12827 and n12446_not n12453 ; n13019
g12828 and n12455_not n13019 ; n13020
g12829 and asqrt[18] n13020 ; n13021
g12830 nor n12446 n12455 ; n13022
g12831 and asqrt[18] n13022 ; n13023
g12832 nor n12453 n13023 ; n13024
g12833 nor n13021 n13024 ; n13025
g12834 nor asqrt[25] n13006 ; n13026
g12835 and n13016_not n13026 ; n13027
g12836 nor n13025 n13027 ; n13028
g12837 nor n13018 n13028 ; n13029
g12838 and asqrt[26] n13029_not ; n13030
g12839 and n12465 n12467_not ; n13031
g12840 and n12458_not n13031 ; n13032
g12841 and asqrt[18] n13032 ; n13033
g12842 nor n12458 n12467 ; n13034
g12843 and asqrt[18] n13034 ; n13035
g12844 nor n12465 n13035 ; n13036
g12845 nor n13033 n13036 ; n13037
g12846 nor asqrt[26] n13018 ; n13038
g12847 and n13028_not n13038 ; n13039
g12848 nor n13037 n13039 ; n13040
g12849 nor n13030 n13040 ; n13041
g12850 and asqrt[27] n13041_not ; n13042
g12851 and n12470_not n12477 ; n13043
g12852 and n12479_not n13043 ; n13044
g12853 and asqrt[18] n13044 ; n13045
g12854 nor n12470 n12479 ; n13046
g12855 and asqrt[18] n13046 ; n13047
g12856 nor n12477 n13047 ; n13048
g12857 nor n13045 n13048 ; n13049
g12858 nor asqrt[27] n13030 ; n13050
g12859 and n13040_not n13050 ; n13051
g12860 nor n13049 n13051 ; n13052
g12861 nor n13042 n13052 ; n13053
g12862 and asqrt[28] n13053_not ; n13054
g12863 and n12489 n12491_not ; n13055
g12864 and n12482_not n13055 ; n13056
g12865 and asqrt[18] n13056 ; n13057
g12866 nor n12482 n12491 ; n13058
g12867 and asqrt[18] n13058 ; n13059
g12868 nor n12489 n13059 ; n13060
g12869 nor n13057 n13060 ; n13061
g12870 nor asqrt[28] n13042 ; n13062
g12871 and n13052_not n13062 ; n13063
g12872 nor n13061 n13063 ; n13064
g12873 nor n13054 n13064 ; n13065
g12874 and asqrt[29] n13065_not ; n13066
g12875 and n12494_not n12501 ; n13067
g12876 and n12503_not n13067 ; n13068
g12877 and asqrt[18] n13068 ; n13069
g12878 nor n12494 n12503 ; n13070
g12879 and asqrt[18] n13070 ; n13071
g12880 nor n12501 n13071 ; n13072
g12881 nor n13069 n13072 ; n13073
g12882 nor asqrt[29] n13054 ; n13074
g12883 and n13064_not n13074 ; n13075
g12884 nor n13073 n13075 ; n13076
g12885 nor n13066 n13076 ; n13077
g12886 and asqrt[30] n13077_not ; n13078
g12887 and n12513 n12515_not ; n13079
g12888 and n12506_not n13079 ; n13080
g12889 and asqrt[18] n13080 ; n13081
g12890 nor n12506 n12515 ; n13082
g12891 and asqrt[18] n13082 ; n13083
g12892 nor n12513 n13083 ; n13084
g12893 nor n13081 n13084 ; n13085
g12894 nor asqrt[30] n13066 ; n13086
g12895 and n13076_not n13086 ; n13087
g12896 nor n13085 n13087 ; n13088
g12897 nor n13078 n13088 ; n13089
g12898 and asqrt[31] n13089_not ; n13090
g12899 and n12518_not n12525 ; n13091
g12900 and n12527_not n13091 ; n13092
g12901 and asqrt[18] n13092 ; n13093
g12902 nor n12518 n12527 ; n13094
g12903 and asqrt[18] n13094 ; n13095
g12904 nor n12525 n13095 ; n13096
g12905 nor n13093 n13096 ; n13097
g12906 nor asqrt[31] n13078 ; n13098
g12907 and n13088_not n13098 ; n13099
g12908 nor n13097 n13099 ; n13100
g12909 nor n13090 n13100 ; n13101
g12910 and asqrt[32] n13101_not ; n13102
g12911 and n12537 n12539_not ; n13103
g12912 and n12530_not n13103 ; n13104
g12913 and asqrt[18] n13104 ; n13105
g12914 nor n12530 n12539 ; n13106
g12915 and asqrt[18] n13106 ; n13107
g12916 nor n12537 n13107 ; n13108
g12917 nor n13105 n13108 ; n13109
g12918 nor asqrt[32] n13090 ; n13110
g12919 and n13100_not n13110 ; n13111
g12920 nor n13109 n13111 ; n13112
g12921 nor n13102 n13112 ; n13113
g12922 and asqrt[33] n13113_not ; n13114
g12923 and n12542_not n12549 ; n13115
g12924 and n12551_not n13115 ; n13116
g12925 and asqrt[18] n13116 ; n13117
g12926 nor n12542 n12551 ; n13118
g12927 and asqrt[18] n13118 ; n13119
g12928 nor n12549 n13119 ; n13120
g12929 nor n13117 n13120 ; n13121
g12930 nor asqrt[33] n13102 ; n13122
g12931 and n13112_not n13122 ; n13123
g12932 nor n13121 n13123 ; n13124
g12933 nor n13114 n13124 ; n13125
g12934 and asqrt[34] n13125_not ; n13126
g12935 and n12561 n12563_not ; n13127
g12936 and n12554_not n13127 ; n13128
g12937 and asqrt[18] n13128 ; n13129
g12938 nor n12554 n12563 ; n13130
g12939 and asqrt[18] n13130 ; n13131
g12940 nor n12561 n13131 ; n13132
g12941 nor n13129 n13132 ; n13133
g12942 nor asqrt[34] n13114 ; n13134
g12943 and n13124_not n13134 ; n13135
g12944 nor n13133 n13135 ; n13136
g12945 nor n13126 n13136 ; n13137
g12946 and asqrt[35] n13137_not ; n13138
g12947 and n12566_not n12573 ; n13139
g12948 and n12575_not n13139 ; n13140
g12949 and asqrt[18] n13140 ; n13141
g12950 nor n12566 n12575 ; n13142
g12951 and asqrt[18] n13142 ; n13143
g12952 nor n12573 n13143 ; n13144
g12953 nor n13141 n13144 ; n13145
g12954 nor asqrt[35] n13126 ; n13146
g12955 and n13136_not n13146 ; n13147
g12956 nor n13145 n13147 ; n13148
g12957 nor n13138 n13148 ; n13149
g12958 and asqrt[36] n13149_not ; n13150
g12959 and n12585 n12587_not ; n13151
g12960 and n12578_not n13151 ; n13152
g12961 and asqrt[18] n13152 ; n13153
g12962 nor n12578 n12587 ; n13154
g12963 and asqrt[18] n13154 ; n13155
g12964 nor n12585 n13155 ; n13156
g12965 nor n13153 n13156 ; n13157
g12966 nor asqrt[36] n13138 ; n13158
g12967 and n13148_not n13158 ; n13159
g12968 nor n13157 n13159 ; n13160
g12969 nor n13150 n13160 ; n13161
g12970 and asqrt[37] n13161_not ; n13162
g12971 and n12590_not n12597 ; n13163
g12972 and n12599_not n13163 ; n13164
g12973 and asqrt[18] n13164 ; n13165
g12974 nor n12590 n12599 ; n13166
g12975 and asqrt[18] n13166 ; n13167
g12976 nor n12597 n13167 ; n13168
g12977 nor n13165 n13168 ; n13169
g12978 nor asqrt[37] n13150 ; n13170
g12979 and n13160_not n13170 ; n13171
g12980 nor n13169 n13171 ; n13172
g12981 nor n13162 n13172 ; n13173
g12982 and asqrt[38] n13173_not ; n13174
g12983 and n12609 n12611_not ; n13175
g12984 and n12602_not n13175 ; n13176
g12985 and asqrt[18] n13176 ; n13177
g12986 nor n12602 n12611 ; n13178
g12987 and asqrt[18] n13178 ; n13179
g12988 nor n12609 n13179 ; n13180
g12989 nor n13177 n13180 ; n13181
g12990 nor asqrt[38] n13162 ; n13182
g12991 and n13172_not n13182 ; n13183
g12992 nor n13181 n13183 ; n13184
g12993 nor n13174 n13184 ; n13185
g12994 and asqrt[39] n13185_not ; n13186
g12995 and n12614_not n12621 ; n13187
g12996 and n12623_not n13187 ; n13188
g12997 and asqrt[18] n13188 ; n13189
g12998 nor n12614 n12623 ; n13190
g12999 and asqrt[18] n13190 ; n13191
g13000 nor n12621 n13191 ; n13192
g13001 nor n13189 n13192 ; n13193
g13002 nor asqrt[39] n13174 ; n13194
g13003 and n13184_not n13194 ; n13195
g13004 nor n13193 n13195 ; n13196
g13005 nor n13186 n13196 ; n13197
g13006 and asqrt[40] n13197_not ; n13198
g13007 and n12633 n12635_not ; n13199
g13008 and n12626_not n13199 ; n13200
g13009 and asqrt[18] n13200 ; n13201
g13010 nor n12626 n12635 ; n13202
g13011 and asqrt[18] n13202 ; n13203
g13012 nor n12633 n13203 ; n13204
g13013 nor n13201 n13204 ; n13205
g13014 nor asqrt[40] n13186 ; n13206
g13015 and n13196_not n13206 ; n13207
g13016 nor n13205 n13207 ; n13208
g13017 nor n13198 n13208 ; n13209
g13018 and asqrt[41] n13209_not ; n13210
g13019 and n12638_not n12645 ; n13211
g13020 and n12647_not n13211 ; n13212
g13021 and asqrt[18] n13212 ; n13213
g13022 nor n12638 n12647 ; n13214
g13023 and asqrt[18] n13214 ; n13215
g13024 nor n12645 n13215 ; n13216
g13025 nor n13213 n13216 ; n13217
g13026 nor asqrt[41] n13198 ; n13218
g13027 and n13208_not n13218 ; n13219
g13028 nor n13217 n13219 ; n13220
g13029 nor n13210 n13220 ; n13221
g13030 and asqrt[42] n13221_not ; n13222
g13031 and n12657 n12659_not ; n13223
g13032 and n12650_not n13223 ; n13224
g13033 and asqrt[18] n13224 ; n13225
g13034 nor n12650 n12659 ; n13226
g13035 and asqrt[18] n13226 ; n13227
g13036 nor n12657 n13227 ; n13228
g13037 nor n13225 n13228 ; n13229
g13038 nor asqrt[42] n13210 ; n13230
g13039 and n13220_not n13230 ; n13231
g13040 nor n13229 n13231 ; n13232
g13041 nor n13222 n13232 ; n13233
g13042 and asqrt[43] n13233_not ; n13234
g13043 and n12662_not n12669 ; n13235
g13044 and n12671_not n13235 ; n13236
g13045 and asqrt[18] n13236 ; n13237
g13046 nor n12662 n12671 ; n13238
g13047 and asqrt[18] n13238 ; n13239
g13048 nor n12669 n13239 ; n13240
g13049 nor n13237 n13240 ; n13241
g13050 nor asqrt[43] n13222 ; n13242
g13051 and n13232_not n13242 ; n13243
g13052 nor n13241 n13243 ; n13244
g13053 nor n13234 n13244 ; n13245
g13054 and asqrt[44] n13245_not ; n13246
g13055 and n12681 n12683_not ; n13247
g13056 and n12674_not n13247 ; n13248
g13057 and asqrt[18] n13248 ; n13249
g13058 nor n12674 n12683 ; n13250
g13059 and asqrt[18] n13250 ; n13251
g13060 nor n12681 n13251 ; n13252
g13061 nor n13249 n13252 ; n13253
g13062 nor asqrt[44] n13234 ; n13254
g13063 and n13244_not n13254 ; n13255
g13064 nor n13253 n13255 ; n13256
g13065 nor n13246 n13256 ; n13257
g13066 and asqrt[45] n13257_not ; n13258
g13067 and n12686_not n12693 ; n13259
g13068 and n12695_not n13259 ; n13260
g13069 and asqrt[18] n13260 ; n13261
g13070 nor n12686 n12695 ; n13262
g13071 and asqrt[18] n13262 ; n13263
g13072 nor n12693 n13263 ; n13264
g13073 nor n13261 n13264 ; n13265
g13074 nor asqrt[45] n13246 ; n13266
g13075 and n13256_not n13266 ; n13267
g13076 nor n13265 n13267 ; n13268
g13077 nor n13258 n13268 ; n13269
g13078 and asqrt[46] n13269_not ; n13270
g13079 and n12705 n12707_not ; n13271
g13080 and n12698_not n13271 ; n13272
g13081 and asqrt[18] n13272 ; n13273
g13082 nor n12698 n12707 ; n13274
g13083 and asqrt[18] n13274 ; n13275
g13084 nor n12705 n13275 ; n13276
g13085 nor n13273 n13276 ; n13277
g13086 nor asqrt[46] n13258 ; n13278
g13087 and n13268_not n13278 ; n13279
g13088 nor n13277 n13279 ; n13280
g13089 nor n13270 n13280 ; n13281
g13090 and asqrt[47] n13281_not ; n13282
g13091 nor asqrt[47] n13270 ; n13283
g13092 and n13280_not n13283 ; n13284
g13093 and n12710_not n12719 ; n13285
g13094 and n12712_not n13285 ; n13286
g13095 and asqrt[18] n13286 ; n13287
g13096 nor n12710 n12712 ; n13288
g13097 and asqrt[18] n13288 ; n13289
g13098 nor n12719 n13289 ; n13290
g13099 nor n13287 n13290 ; n13291
g13100 nor n13284 n13291 ; n13292
g13101 nor n13282 n13292 ; n13293
g13102 and asqrt[48] n13293_not ; n13294
g13103 and n12729 n12731_not ; n13295
g13104 and n12722_not n13295 ; n13296
g13105 and asqrt[18] n13296 ; n13297
g13106 nor n12722 n12731 ; n13298
g13107 and asqrt[18] n13298 ; n13299
g13108 nor n12729 n13299 ; n13300
g13109 nor n13297 n13300 ; n13301
g13110 nor asqrt[48] n13282 ; n13302
g13111 and n13292_not n13302 ; n13303
g13112 nor n13301 n13303 ; n13304
g13113 nor n13294 n13304 ; n13305
g13114 and asqrt[49] n13305_not ; n13306
g13115 and n12734_not n12741 ; n13307
g13116 and n12743_not n13307 ; n13308
g13117 and asqrt[18] n13308 ; n13309
g13118 nor n12734 n12743 ; n13310
g13119 and asqrt[18] n13310 ; n13311
g13120 nor n12741 n13311 ; n13312
g13121 nor n13309 n13312 ; n13313
g13122 nor asqrt[49] n13294 ; n13314
g13123 and n13304_not n13314 ; n13315
g13124 nor n13313 n13315 ; n13316
g13125 nor n13306 n13316 ; n13317
g13126 and asqrt[50] n13317_not ; n13318
g13127 and n12753 n12755_not ; n13319
g13128 and n12746_not n13319 ; n13320
g13129 and asqrt[18] n13320 ; n13321
g13130 nor n12746 n12755 ; n13322
g13131 and asqrt[18] n13322 ; n13323
g13132 nor n12753 n13323 ; n13324
g13133 nor n13321 n13324 ; n13325
g13134 nor asqrt[50] n13306 ; n13326
g13135 and n13316_not n13326 ; n13327
g13136 nor n13325 n13327 ; n13328
g13137 nor n13318 n13328 ; n13329
g13138 and asqrt[51] n13329_not ; n13330
g13139 and n12758_not n12765 ; n13331
g13140 and n12767_not n13331 ; n13332
g13141 and asqrt[18] n13332 ; n13333
g13142 nor n12758 n12767 ; n13334
g13143 and asqrt[18] n13334 ; n13335
g13144 nor n12765 n13335 ; n13336
g13145 nor n13333 n13336 ; n13337
g13146 nor asqrt[51] n13318 ; n13338
g13147 and n13328_not n13338 ; n13339
g13148 nor n13337 n13339 ; n13340
g13149 nor n13330 n13340 ; n13341
g13150 and asqrt[52] n13341_not ; n13342
g13151 and n12777 n12779_not ; n13343
g13152 and n12770_not n13343 ; n13344
g13153 and asqrt[18] n13344 ; n13345
g13154 nor n12770 n12779 ; n13346
g13155 and asqrt[18] n13346 ; n13347
g13156 nor n12777 n13347 ; n13348
g13157 nor n13345 n13348 ; n13349
g13158 nor asqrt[52] n13330 ; n13350
g13159 and n13340_not n13350 ; n13351
g13160 nor n13349 n13351 ; n13352
g13161 nor n13342 n13352 ; n13353
g13162 and asqrt[53] n13353_not ; n13354
g13163 and n12782_not n12789 ; n13355
g13164 and n12791_not n13355 ; n13356
g13165 and asqrt[18] n13356 ; n13357
g13166 nor n12782 n12791 ; n13358
g13167 and asqrt[18] n13358 ; n13359
g13168 nor n12789 n13359 ; n13360
g13169 nor n13357 n13360 ; n13361
g13170 nor asqrt[53] n13342 ; n13362
g13171 and n13352_not n13362 ; n13363
g13172 nor n13361 n13363 ; n13364
g13173 nor n13354 n13364 ; n13365
g13174 and asqrt[54] n13365_not ; n13366
g13175 and n12801 n12803_not ; n13367
g13176 and n12794_not n13367 ; n13368
g13177 and asqrt[18] n13368 ; n13369
g13178 nor n12794 n12803 ; n13370
g13179 and asqrt[18] n13370 ; n13371
g13180 nor n12801 n13371 ; n13372
g13181 nor n13369 n13372 ; n13373
g13182 nor asqrt[54] n13354 ; n13374
g13183 and n13364_not n13374 ; n13375
g13184 nor n13373 n13375 ; n13376
g13185 nor n13366 n13376 ; n13377
g13186 and asqrt[55] n13377_not ; n13378
g13187 and n12806_not n12813 ; n13379
g13188 and n12815_not n13379 ; n13380
g13189 and asqrt[18] n13380 ; n13381
g13190 nor n12806 n12815 ; n13382
g13191 and asqrt[18] n13382 ; n13383
g13192 nor n12813 n13383 ; n13384
g13193 nor n13381 n13384 ; n13385
g13194 nor asqrt[55] n13366 ; n13386
g13195 and n13376_not n13386 ; n13387
g13196 nor n13385 n13387 ; n13388
g13197 nor n13378 n13388 ; n13389
g13198 and asqrt[56] n13389_not ; n13390
g13199 and n12825 n12827_not ; n13391
g13200 and n12818_not n13391 ; n13392
g13201 and asqrt[18] n13392 ; n13393
g13202 nor n12818 n12827 ; n13394
g13203 and asqrt[18] n13394 ; n13395
g13204 nor n12825 n13395 ; n13396
g13205 nor n13393 n13396 ; n13397
g13206 nor asqrt[56] n13378 ; n13398
g13207 and n13388_not n13398 ; n13399
g13208 nor n13397 n13399 ; n13400
g13209 nor n13390 n13400 ; n13401
g13210 and asqrt[57] n13401_not ; n13402
g13211 and n12830_not n12837 ; n13403
g13212 and n12839_not n13403 ; n13404
g13213 and asqrt[18] n13404 ; n13405
g13214 nor n12830 n12839 ; n13406
g13215 and asqrt[18] n13406 ; n13407
g13216 nor n12837 n13407 ; n13408
g13217 nor n13405 n13408 ; n13409
g13218 nor asqrt[57] n13390 ; n13410
g13219 and n13400_not n13410 ; n13411
g13220 nor n13409 n13411 ; n13412
g13221 nor n13402 n13412 ; n13413
g13222 and asqrt[58] n13413_not ; n13414
g13223 and n12849 n12851_not ; n13415
g13224 and n12842_not n13415 ; n13416
g13225 and asqrt[18] n13416 ; n13417
g13226 nor n12842 n12851 ; n13418
g13227 and asqrt[18] n13418 ; n13419
g13228 nor n12849 n13419 ; n13420
g13229 nor n13417 n13420 ; n13421
g13230 nor asqrt[58] n13402 ; n13422
g13231 and n13412_not n13422 ; n13423
g13232 nor n13421 n13423 ; n13424
g13233 nor n13414 n13424 ; n13425
g13234 and asqrt[59] n13425_not ; n13426
g13235 and n12854_not n12861 ; n13427
g13236 and n12863_not n13427 ; n13428
g13237 and asqrt[18] n13428 ; n13429
g13238 nor n12854 n12863 ; n13430
g13239 and asqrt[18] n13430 ; n13431
g13240 nor n12861 n13431 ; n13432
g13241 nor n13429 n13432 ; n13433
g13242 nor asqrt[59] n13414 ; n13434
g13243 and n13424_not n13434 ; n13435
g13244 nor n13433 n13435 ; n13436
g13245 nor n13426 n13436 ; n13437
g13246 and asqrt[60] n13437_not ; n13438
g13247 and n12873 n12875_not ; n13439
g13248 and n12866_not n13439 ; n13440
g13249 and asqrt[18] n13440 ; n13441
g13250 nor n12866 n12875 ; n13442
g13251 and asqrt[18] n13442 ; n13443
g13252 nor n12873 n13443 ; n13444
g13253 nor n13441 n13444 ; n13445
g13254 nor asqrt[60] n13426 ; n13446
g13255 and n13436_not n13446 ; n13447
g13256 nor n13445 n13447 ; n13448
g13257 nor n13438 n13448 ; n13449
g13258 and asqrt[61] n13449_not ; n13450
g13259 and n12878_not n12885 ; n13451
g13260 and n12887_not n13451 ; n13452
g13261 and asqrt[18] n13452 ; n13453
g13262 nor n12878 n12887 ; n13454
g13263 and asqrt[18] n13454 ; n13455
g13264 nor n12885 n13455 ; n13456
g13265 nor n13453 n13456 ; n13457
g13266 nor asqrt[61] n13438 ; n13458
g13267 and n13448_not n13458 ; n13459
g13268 nor n13457 n13459 ; n13460
g13269 nor n13450 n13460 ; n13461
g13270 and asqrt[62] n13461_not ; n13462
g13271 and n12897 n12899_not ; n13463
g13272 and n12890_not n13463 ; n13464
g13273 and asqrt[18] n13464 ; n13465
g13274 nor n12890 n12899 ; n13466
g13275 and asqrt[18] n13466 ; n13467
g13276 nor n12897 n13467 ; n13468
g13277 nor n13465 n13468 ; n13469
g13278 nor asqrt[62] n13450 ; n13470
g13279 and n13460_not n13470 ; n13471
g13280 nor n13469 n13471 ; n13472
g13281 nor n13462 n13472 ; n13473
g13282 and n12902_not n12909 ; n13474
g13283 and n12911_not n13474 ; n13475
g13284 and asqrt[18] n13475 ; n13476
g13285 nor n12902 n12911 ; n13477
g13286 and asqrt[18] n13477 ; n13478
g13287 nor n12909 n13478 ; n13479
g13288 nor n13476 n13479 ; n13480
g13289 nor n12913 n12920 ; n13481
g13290 and asqrt[18] n13481 ; n13482
g13291 nor n12928 n13482 ; n13483
g13292 and n13480_not n13483 ; n13484
g13293 and n13473_not n13484 ; n13485
g13294 nor asqrt[63] n13485 ; n13486
g13295 and n13462_not n13480 ; n13487
g13296 and n13472_not n13487 ; n13488
g13297 and n12920_not asqrt[18] ; n13489
g13298 and n12913 n13489_not ; n13490
g13299 and asqrt[63] n13481_not ; n13491
g13300 and n13490_not n13491 ; n13492
g13301 nor n12916 n12937 ; n13493
g13302 and n12919_not n13493 ; n13494
g13303 and n12932_not n13494 ; n13495
g13304 and n12928_not n13495 ; n13496
g13305 and n12926_not n13496 ; n13497
g13306 nor n13492 n13497 ; n13498
g13307 and n13488_not n13498 ; n13499
g13308 nand n13486_not n13499 ; asqrt[17]
g13309 and a[34] asqrt[17] ; n13501
g13310 nor a[32] a[33] ; n13502
g13311 and a[34]_not n13502 ; n13503
g13312 nor n13501 n13503 ; n13504
g13313 and asqrt[18] n13504_not ; n13505
g13314 nor n12937 n13503 ; n13506
g13315 and n12932_not n13506 ; n13507
g13316 and n12928_not n13507 ; n13508
g13317 and n12926_not n13508 ; n13509
g13318 and n13501_not n13509 ; n13510
g13319 and a[34]_not asqrt[17] ; n13511
g13320 and a[35] n13511_not ; n13512
g13321 and n12942 asqrt[17] ; n13513
g13322 nor n13512 n13513 ; n13514
g13323 and n13510_not n13514 ; n13515
g13324 nor n13505 n13515 ; n13516
g13325 and asqrt[19] n13516_not ; n13517
g13326 nor asqrt[19] n13505 ; n13518
g13327 and n13515_not n13518 ; n13519
g13328 and asqrt[18] n13497_not ; n13520
g13329 and n13492_not n13520 ; n13521
g13330 and n13488_not n13521 ; n13522
g13331 and n13486_not n13522 ; n13523
g13332 nor n13513 n13523 ; n13524
g13333 and a[36] n13524_not ; n13525
g13334 nor a[36] n13523 ; n13526
g13335 and n13513_not n13526 ; n13527
g13336 nor n13525 n13527 ; n13528
g13337 nor n13519 n13528 ; n13529
g13338 nor n13517 n13529 ; n13530
g13339 and asqrt[20] n13530_not ; n13531
g13340 nor n12945 n12950 ; n13532
g13341 and n12954_not n13532 ; n13533
g13342 and asqrt[17] n13533 ; n13534
g13343 and asqrt[17] n13532 ; n13535
g13344 and n12954 n13535_not ; n13536
g13345 nor n13534 n13536 ; n13537
g13346 nor asqrt[20] n13517 ; n13538
g13347 and n13529_not n13538 ; n13539
g13348 nor n13537 n13539 ; n13540
g13349 nor n13531 n13540 ; n13541
g13350 and asqrt[21] n13541_not ; n13542
g13351 and n12959_not n12968 ; n13543
g13352 and n12957_not n13543 ; n13544
g13353 and asqrt[17] n13544 ; n13545
g13354 nor n12957 n12959 ; n13546
g13355 and asqrt[17] n13546 ; n13547
g13356 nor n12968 n13547 ; n13548
g13357 nor n13545 n13548 ; n13549
g13358 nor asqrt[21] n13531 ; n13550
g13359 and n13540_not n13550 ; n13551
g13360 nor n13549 n13551 ; n13552
g13361 nor n13542 n13552 ; n13553
g13362 and asqrt[22] n13553_not ; n13554
g13363 and n12971_not n12977 ; n13555
g13364 and n12979_not n13555 ; n13556
g13365 and asqrt[17] n13556 ; n13557
g13366 nor n12971 n12979 ; n13558
g13367 and asqrt[17] n13558 ; n13559
g13368 nor n12977 n13559 ; n13560
g13369 nor n13557 n13560 ; n13561
g13370 nor asqrt[22] n13542 ; n13562
g13371 and n13552_not n13562 ; n13563
g13372 nor n13561 n13563 ; n13564
g13373 nor n13554 n13564 ; n13565
g13374 and asqrt[23] n13565_not ; n13566
g13375 and n12989 n12991_not ; n13567
g13376 and n12982_not n13567 ; n13568
g13377 and asqrt[17] n13568 ; n13569
g13378 nor n12982 n12991 ; n13570
g13379 and asqrt[17] n13570 ; n13571
g13380 nor n12989 n13571 ; n13572
g13381 nor n13569 n13572 ; n13573
g13382 nor asqrt[23] n13554 ; n13574
g13383 and n13564_not n13574 ; n13575
g13384 nor n13573 n13575 ; n13576
g13385 nor n13566 n13576 ; n13577
g13386 and asqrt[24] n13577_not ; n13578
g13387 and n12994_not n13001 ; n13579
g13388 and n13003_not n13579 ; n13580
g13389 and asqrt[17] n13580 ; n13581
g13390 nor n12994 n13003 ; n13582
g13391 and asqrt[17] n13582 ; n13583
g13392 nor n13001 n13583 ; n13584
g13393 nor n13581 n13584 ; n13585
g13394 nor asqrt[24] n13566 ; n13586
g13395 and n13576_not n13586 ; n13587
g13396 nor n13585 n13587 ; n13588
g13397 nor n13578 n13588 ; n13589
g13398 and asqrt[25] n13589_not ; n13590
g13399 and n13013 n13015_not ; n13591
g13400 and n13006_not n13591 ; n13592
g13401 and asqrt[17] n13592 ; n13593
g13402 nor n13006 n13015 ; n13594
g13403 and asqrt[17] n13594 ; n13595
g13404 nor n13013 n13595 ; n13596
g13405 nor n13593 n13596 ; n13597
g13406 nor asqrt[25] n13578 ; n13598
g13407 and n13588_not n13598 ; n13599
g13408 nor n13597 n13599 ; n13600
g13409 nor n13590 n13600 ; n13601
g13410 and asqrt[26] n13601_not ; n13602
g13411 and n13018_not n13025 ; n13603
g13412 and n13027_not n13603 ; n13604
g13413 and asqrt[17] n13604 ; n13605
g13414 nor n13018 n13027 ; n13606
g13415 and asqrt[17] n13606 ; n13607
g13416 nor n13025 n13607 ; n13608
g13417 nor n13605 n13608 ; n13609
g13418 nor asqrt[26] n13590 ; n13610
g13419 and n13600_not n13610 ; n13611
g13420 nor n13609 n13611 ; n13612
g13421 nor n13602 n13612 ; n13613
g13422 and asqrt[27] n13613_not ; n13614
g13423 and n13037 n13039_not ; n13615
g13424 and n13030_not n13615 ; n13616
g13425 and asqrt[17] n13616 ; n13617
g13426 nor n13030 n13039 ; n13618
g13427 and asqrt[17] n13618 ; n13619
g13428 nor n13037 n13619 ; n13620
g13429 nor n13617 n13620 ; n13621
g13430 nor asqrt[27] n13602 ; n13622
g13431 and n13612_not n13622 ; n13623
g13432 nor n13621 n13623 ; n13624
g13433 nor n13614 n13624 ; n13625
g13434 and asqrt[28] n13625_not ; n13626
g13435 and n13042_not n13049 ; n13627
g13436 and n13051_not n13627 ; n13628
g13437 and asqrt[17] n13628 ; n13629
g13438 nor n13042 n13051 ; n13630
g13439 and asqrt[17] n13630 ; n13631
g13440 nor n13049 n13631 ; n13632
g13441 nor n13629 n13632 ; n13633
g13442 nor asqrt[28] n13614 ; n13634
g13443 and n13624_not n13634 ; n13635
g13444 nor n13633 n13635 ; n13636
g13445 nor n13626 n13636 ; n13637
g13446 and asqrt[29] n13637_not ; n13638
g13447 and n13061 n13063_not ; n13639
g13448 and n13054_not n13639 ; n13640
g13449 and asqrt[17] n13640 ; n13641
g13450 nor n13054 n13063 ; n13642
g13451 and asqrt[17] n13642 ; n13643
g13452 nor n13061 n13643 ; n13644
g13453 nor n13641 n13644 ; n13645
g13454 nor asqrt[29] n13626 ; n13646
g13455 and n13636_not n13646 ; n13647
g13456 nor n13645 n13647 ; n13648
g13457 nor n13638 n13648 ; n13649
g13458 and asqrt[30] n13649_not ; n13650
g13459 and n13066_not n13073 ; n13651
g13460 and n13075_not n13651 ; n13652
g13461 and asqrt[17] n13652 ; n13653
g13462 nor n13066 n13075 ; n13654
g13463 and asqrt[17] n13654 ; n13655
g13464 nor n13073 n13655 ; n13656
g13465 nor n13653 n13656 ; n13657
g13466 nor asqrt[30] n13638 ; n13658
g13467 and n13648_not n13658 ; n13659
g13468 nor n13657 n13659 ; n13660
g13469 nor n13650 n13660 ; n13661
g13470 and asqrt[31] n13661_not ; n13662
g13471 and n13085 n13087_not ; n13663
g13472 and n13078_not n13663 ; n13664
g13473 and asqrt[17] n13664 ; n13665
g13474 nor n13078 n13087 ; n13666
g13475 and asqrt[17] n13666 ; n13667
g13476 nor n13085 n13667 ; n13668
g13477 nor n13665 n13668 ; n13669
g13478 nor asqrt[31] n13650 ; n13670
g13479 and n13660_not n13670 ; n13671
g13480 nor n13669 n13671 ; n13672
g13481 nor n13662 n13672 ; n13673
g13482 and asqrt[32] n13673_not ; n13674
g13483 and n13090_not n13097 ; n13675
g13484 and n13099_not n13675 ; n13676
g13485 and asqrt[17] n13676 ; n13677
g13486 nor n13090 n13099 ; n13678
g13487 and asqrt[17] n13678 ; n13679
g13488 nor n13097 n13679 ; n13680
g13489 nor n13677 n13680 ; n13681
g13490 nor asqrt[32] n13662 ; n13682
g13491 and n13672_not n13682 ; n13683
g13492 nor n13681 n13683 ; n13684
g13493 nor n13674 n13684 ; n13685
g13494 and asqrt[33] n13685_not ; n13686
g13495 and n13109 n13111_not ; n13687
g13496 and n13102_not n13687 ; n13688
g13497 and asqrt[17] n13688 ; n13689
g13498 nor n13102 n13111 ; n13690
g13499 and asqrt[17] n13690 ; n13691
g13500 nor n13109 n13691 ; n13692
g13501 nor n13689 n13692 ; n13693
g13502 nor asqrt[33] n13674 ; n13694
g13503 and n13684_not n13694 ; n13695
g13504 nor n13693 n13695 ; n13696
g13505 nor n13686 n13696 ; n13697
g13506 and asqrt[34] n13697_not ; n13698
g13507 and n13114_not n13121 ; n13699
g13508 and n13123_not n13699 ; n13700
g13509 and asqrt[17] n13700 ; n13701
g13510 nor n13114 n13123 ; n13702
g13511 and asqrt[17] n13702 ; n13703
g13512 nor n13121 n13703 ; n13704
g13513 nor n13701 n13704 ; n13705
g13514 nor asqrt[34] n13686 ; n13706
g13515 and n13696_not n13706 ; n13707
g13516 nor n13705 n13707 ; n13708
g13517 nor n13698 n13708 ; n13709
g13518 and asqrt[35] n13709_not ; n13710
g13519 and n13133 n13135_not ; n13711
g13520 and n13126_not n13711 ; n13712
g13521 and asqrt[17] n13712 ; n13713
g13522 nor n13126 n13135 ; n13714
g13523 and asqrt[17] n13714 ; n13715
g13524 nor n13133 n13715 ; n13716
g13525 nor n13713 n13716 ; n13717
g13526 nor asqrt[35] n13698 ; n13718
g13527 and n13708_not n13718 ; n13719
g13528 nor n13717 n13719 ; n13720
g13529 nor n13710 n13720 ; n13721
g13530 and asqrt[36] n13721_not ; n13722
g13531 and n13138_not n13145 ; n13723
g13532 and n13147_not n13723 ; n13724
g13533 and asqrt[17] n13724 ; n13725
g13534 nor n13138 n13147 ; n13726
g13535 and asqrt[17] n13726 ; n13727
g13536 nor n13145 n13727 ; n13728
g13537 nor n13725 n13728 ; n13729
g13538 nor asqrt[36] n13710 ; n13730
g13539 and n13720_not n13730 ; n13731
g13540 nor n13729 n13731 ; n13732
g13541 nor n13722 n13732 ; n13733
g13542 and asqrt[37] n13733_not ; n13734
g13543 and n13157 n13159_not ; n13735
g13544 and n13150_not n13735 ; n13736
g13545 and asqrt[17] n13736 ; n13737
g13546 nor n13150 n13159 ; n13738
g13547 and asqrt[17] n13738 ; n13739
g13548 nor n13157 n13739 ; n13740
g13549 nor n13737 n13740 ; n13741
g13550 nor asqrt[37] n13722 ; n13742
g13551 and n13732_not n13742 ; n13743
g13552 nor n13741 n13743 ; n13744
g13553 nor n13734 n13744 ; n13745
g13554 and asqrt[38] n13745_not ; n13746
g13555 and n13162_not n13169 ; n13747
g13556 and n13171_not n13747 ; n13748
g13557 and asqrt[17] n13748 ; n13749
g13558 nor n13162 n13171 ; n13750
g13559 and asqrt[17] n13750 ; n13751
g13560 nor n13169 n13751 ; n13752
g13561 nor n13749 n13752 ; n13753
g13562 nor asqrt[38] n13734 ; n13754
g13563 and n13744_not n13754 ; n13755
g13564 nor n13753 n13755 ; n13756
g13565 nor n13746 n13756 ; n13757
g13566 and asqrt[39] n13757_not ; n13758
g13567 and n13181 n13183_not ; n13759
g13568 and n13174_not n13759 ; n13760
g13569 and asqrt[17] n13760 ; n13761
g13570 nor n13174 n13183 ; n13762
g13571 and asqrt[17] n13762 ; n13763
g13572 nor n13181 n13763 ; n13764
g13573 nor n13761 n13764 ; n13765
g13574 nor asqrt[39] n13746 ; n13766
g13575 and n13756_not n13766 ; n13767
g13576 nor n13765 n13767 ; n13768
g13577 nor n13758 n13768 ; n13769
g13578 and asqrt[40] n13769_not ; n13770
g13579 and n13186_not n13193 ; n13771
g13580 and n13195_not n13771 ; n13772
g13581 and asqrt[17] n13772 ; n13773
g13582 nor n13186 n13195 ; n13774
g13583 and asqrt[17] n13774 ; n13775
g13584 nor n13193 n13775 ; n13776
g13585 nor n13773 n13776 ; n13777
g13586 nor asqrt[40] n13758 ; n13778
g13587 and n13768_not n13778 ; n13779
g13588 nor n13777 n13779 ; n13780
g13589 nor n13770 n13780 ; n13781
g13590 and asqrt[41] n13781_not ; n13782
g13591 and n13205 n13207_not ; n13783
g13592 and n13198_not n13783 ; n13784
g13593 and asqrt[17] n13784 ; n13785
g13594 nor n13198 n13207 ; n13786
g13595 and asqrt[17] n13786 ; n13787
g13596 nor n13205 n13787 ; n13788
g13597 nor n13785 n13788 ; n13789
g13598 nor asqrt[41] n13770 ; n13790
g13599 and n13780_not n13790 ; n13791
g13600 nor n13789 n13791 ; n13792
g13601 nor n13782 n13792 ; n13793
g13602 and asqrt[42] n13793_not ; n13794
g13603 and n13210_not n13217 ; n13795
g13604 and n13219_not n13795 ; n13796
g13605 and asqrt[17] n13796 ; n13797
g13606 nor n13210 n13219 ; n13798
g13607 and asqrt[17] n13798 ; n13799
g13608 nor n13217 n13799 ; n13800
g13609 nor n13797 n13800 ; n13801
g13610 nor asqrt[42] n13782 ; n13802
g13611 and n13792_not n13802 ; n13803
g13612 nor n13801 n13803 ; n13804
g13613 nor n13794 n13804 ; n13805
g13614 and asqrt[43] n13805_not ; n13806
g13615 and n13229 n13231_not ; n13807
g13616 and n13222_not n13807 ; n13808
g13617 and asqrt[17] n13808 ; n13809
g13618 nor n13222 n13231 ; n13810
g13619 and asqrt[17] n13810 ; n13811
g13620 nor n13229 n13811 ; n13812
g13621 nor n13809 n13812 ; n13813
g13622 nor asqrt[43] n13794 ; n13814
g13623 and n13804_not n13814 ; n13815
g13624 nor n13813 n13815 ; n13816
g13625 nor n13806 n13816 ; n13817
g13626 and asqrt[44] n13817_not ; n13818
g13627 and n13234_not n13241 ; n13819
g13628 and n13243_not n13819 ; n13820
g13629 and asqrt[17] n13820 ; n13821
g13630 nor n13234 n13243 ; n13822
g13631 and asqrt[17] n13822 ; n13823
g13632 nor n13241 n13823 ; n13824
g13633 nor n13821 n13824 ; n13825
g13634 nor asqrt[44] n13806 ; n13826
g13635 and n13816_not n13826 ; n13827
g13636 nor n13825 n13827 ; n13828
g13637 nor n13818 n13828 ; n13829
g13638 and asqrt[45] n13829_not ; n13830
g13639 and n13253 n13255_not ; n13831
g13640 and n13246_not n13831 ; n13832
g13641 and asqrt[17] n13832 ; n13833
g13642 nor n13246 n13255 ; n13834
g13643 and asqrt[17] n13834 ; n13835
g13644 nor n13253 n13835 ; n13836
g13645 nor n13833 n13836 ; n13837
g13646 nor asqrt[45] n13818 ; n13838
g13647 and n13828_not n13838 ; n13839
g13648 nor n13837 n13839 ; n13840
g13649 nor n13830 n13840 ; n13841
g13650 and asqrt[46] n13841_not ; n13842
g13651 and n13258_not n13265 ; n13843
g13652 and n13267_not n13843 ; n13844
g13653 and asqrt[17] n13844 ; n13845
g13654 nor n13258 n13267 ; n13846
g13655 and asqrt[17] n13846 ; n13847
g13656 nor n13265 n13847 ; n13848
g13657 nor n13845 n13848 ; n13849
g13658 nor asqrt[46] n13830 ; n13850
g13659 and n13840_not n13850 ; n13851
g13660 nor n13849 n13851 ; n13852
g13661 nor n13842 n13852 ; n13853
g13662 and asqrt[47] n13853_not ; n13854
g13663 and n13277 n13279_not ; n13855
g13664 and n13270_not n13855 ; n13856
g13665 and asqrt[17] n13856 ; n13857
g13666 nor n13270 n13279 ; n13858
g13667 and asqrt[17] n13858 ; n13859
g13668 nor n13277 n13859 ; n13860
g13669 nor n13857 n13860 ; n13861
g13670 nor asqrt[47] n13842 ; n13862
g13671 and n13852_not n13862 ; n13863
g13672 nor n13861 n13863 ; n13864
g13673 nor n13854 n13864 ; n13865
g13674 and asqrt[48] n13865_not ; n13866
g13675 nor asqrt[48] n13854 ; n13867
g13676 and n13864_not n13867 ; n13868
g13677 and n13282_not n13291 ; n13869
g13678 and n13284_not n13869 ; n13870
g13679 and asqrt[17] n13870 ; n13871
g13680 nor n13282 n13284 ; n13872
g13681 and asqrt[17] n13872 ; n13873
g13682 nor n13291 n13873 ; n13874
g13683 nor n13871 n13874 ; n13875
g13684 nor n13868 n13875 ; n13876
g13685 nor n13866 n13876 ; n13877
g13686 and asqrt[49] n13877_not ; n13878
g13687 and n13301 n13303_not ; n13879
g13688 and n13294_not n13879 ; n13880
g13689 and asqrt[17] n13880 ; n13881
g13690 nor n13294 n13303 ; n13882
g13691 and asqrt[17] n13882 ; n13883
g13692 nor n13301 n13883 ; n13884
g13693 nor n13881 n13884 ; n13885
g13694 nor asqrt[49] n13866 ; n13886
g13695 and n13876_not n13886 ; n13887
g13696 nor n13885 n13887 ; n13888
g13697 nor n13878 n13888 ; n13889
g13698 and asqrt[50] n13889_not ; n13890
g13699 and n13306_not n13313 ; n13891
g13700 and n13315_not n13891 ; n13892
g13701 and asqrt[17] n13892 ; n13893
g13702 nor n13306 n13315 ; n13894
g13703 and asqrt[17] n13894 ; n13895
g13704 nor n13313 n13895 ; n13896
g13705 nor n13893 n13896 ; n13897
g13706 nor asqrt[50] n13878 ; n13898
g13707 and n13888_not n13898 ; n13899
g13708 nor n13897 n13899 ; n13900
g13709 nor n13890 n13900 ; n13901
g13710 and asqrt[51] n13901_not ; n13902
g13711 and n13325 n13327_not ; n13903
g13712 and n13318_not n13903 ; n13904
g13713 and asqrt[17] n13904 ; n13905
g13714 nor n13318 n13327 ; n13906
g13715 and asqrt[17] n13906 ; n13907
g13716 nor n13325 n13907 ; n13908
g13717 nor n13905 n13908 ; n13909
g13718 nor asqrt[51] n13890 ; n13910
g13719 and n13900_not n13910 ; n13911
g13720 nor n13909 n13911 ; n13912
g13721 nor n13902 n13912 ; n13913
g13722 and asqrt[52] n13913_not ; n13914
g13723 and n13330_not n13337 ; n13915
g13724 and n13339_not n13915 ; n13916
g13725 and asqrt[17] n13916 ; n13917
g13726 nor n13330 n13339 ; n13918
g13727 and asqrt[17] n13918 ; n13919
g13728 nor n13337 n13919 ; n13920
g13729 nor n13917 n13920 ; n13921
g13730 nor asqrt[52] n13902 ; n13922
g13731 and n13912_not n13922 ; n13923
g13732 nor n13921 n13923 ; n13924
g13733 nor n13914 n13924 ; n13925
g13734 and asqrt[53] n13925_not ; n13926
g13735 and n13349 n13351_not ; n13927
g13736 and n13342_not n13927 ; n13928
g13737 and asqrt[17] n13928 ; n13929
g13738 nor n13342 n13351 ; n13930
g13739 and asqrt[17] n13930 ; n13931
g13740 nor n13349 n13931 ; n13932
g13741 nor n13929 n13932 ; n13933
g13742 nor asqrt[53] n13914 ; n13934
g13743 and n13924_not n13934 ; n13935
g13744 nor n13933 n13935 ; n13936
g13745 nor n13926 n13936 ; n13937
g13746 and asqrt[54] n13937_not ; n13938
g13747 and n13354_not n13361 ; n13939
g13748 and n13363_not n13939 ; n13940
g13749 and asqrt[17] n13940 ; n13941
g13750 nor n13354 n13363 ; n13942
g13751 and asqrt[17] n13942 ; n13943
g13752 nor n13361 n13943 ; n13944
g13753 nor n13941 n13944 ; n13945
g13754 nor asqrt[54] n13926 ; n13946
g13755 and n13936_not n13946 ; n13947
g13756 nor n13945 n13947 ; n13948
g13757 nor n13938 n13948 ; n13949
g13758 and asqrt[55] n13949_not ; n13950
g13759 and n13373 n13375_not ; n13951
g13760 and n13366_not n13951 ; n13952
g13761 and asqrt[17] n13952 ; n13953
g13762 nor n13366 n13375 ; n13954
g13763 and asqrt[17] n13954 ; n13955
g13764 nor n13373 n13955 ; n13956
g13765 nor n13953 n13956 ; n13957
g13766 nor asqrt[55] n13938 ; n13958
g13767 and n13948_not n13958 ; n13959
g13768 nor n13957 n13959 ; n13960
g13769 nor n13950 n13960 ; n13961
g13770 and asqrt[56] n13961_not ; n13962
g13771 and n13378_not n13385 ; n13963
g13772 and n13387_not n13963 ; n13964
g13773 and asqrt[17] n13964 ; n13965
g13774 nor n13378 n13387 ; n13966
g13775 and asqrt[17] n13966 ; n13967
g13776 nor n13385 n13967 ; n13968
g13777 nor n13965 n13968 ; n13969
g13778 nor asqrt[56] n13950 ; n13970
g13779 and n13960_not n13970 ; n13971
g13780 nor n13969 n13971 ; n13972
g13781 nor n13962 n13972 ; n13973
g13782 and asqrt[57] n13973_not ; n13974
g13783 and n13397 n13399_not ; n13975
g13784 and n13390_not n13975 ; n13976
g13785 and asqrt[17] n13976 ; n13977
g13786 nor n13390 n13399 ; n13978
g13787 and asqrt[17] n13978 ; n13979
g13788 nor n13397 n13979 ; n13980
g13789 nor n13977 n13980 ; n13981
g13790 nor asqrt[57] n13962 ; n13982
g13791 and n13972_not n13982 ; n13983
g13792 nor n13981 n13983 ; n13984
g13793 nor n13974 n13984 ; n13985
g13794 and asqrt[58] n13985_not ; n13986
g13795 and n13402_not n13409 ; n13987
g13796 and n13411_not n13987 ; n13988
g13797 and asqrt[17] n13988 ; n13989
g13798 nor n13402 n13411 ; n13990
g13799 and asqrt[17] n13990 ; n13991
g13800 nor n13409 n13991 ; n13992
g13801 nor n13989 n13992 ; n13993
g13802 nor asqrt[58] n13974 ; n13994
g13803 and n13984_not n13994 ; n13995
g13804 nor n13993 n13995 ; n13996
g13805 nor n13986 n13996 ; n13997
g13806 and asqrt[59] n13997_not ; n13998
g13807 and n13421 n13423_not ; n13999
g13808 and n13414_not n13999 ; n14000
g13809 and asqrt[17] n14000 ; n14001
g13810 nor n13414 n13423 ; n14002
g13811 and asqrt[17] n14002 ; n14003
g13812 nor n13421 n14003 ; n14004
g13813 nor n14001 n14004 ; n14005
g13814 nor asqrt[59] n13986 ; n14006
g13815 and n13996_not n14006 ; n14007
g13816 nor n14005 n14007 ; n14008
g13817 nor n13998 n14008 ; n14009
g13818 and asqrt[60] n14009_not ; n14010
g13819 and n13426_not n13433 ; n14011
g13820 and n13435_not n14011 ; n14012
g13821 and asqrt[17] n14012 ; n14013
g13822 nor n13426 n13435 ; n14014
g13823 and asqrt[17] n14014 ; n14015
g13824 nor n13433 n14015 ; n14016
g13825 nor n14013 n14016 ; n14017
g13826 nor asqrt[60] n13998 ; n14018
g13827 and n14008_not n14018 ; n14019
g13828 nor n14017 n14019 ; n14020
g13829 nor n14010 n14020 ; n14021
g13830 and asqrt[61] n14021_not ; n14022
g13831 and n13445 n13447_not ; n14023
g13832 and n13438_not n14023 ; n14024
g13833 and asqrt[17] n14024 ; n14025
g13834 nor n13438 n13447 ; n14026
g13835 and asqrt[17] n14026 ; n14027
g13836 nor n13445 n14027 ; n14028
g13837 nor n14025 n14028 ; n14029
g13838 nor asqrt[61] n14010 ; n14030
g13839 and n14020_not n14030 ; n14031
g13840 nor n14029 n14031 ; n14032
g13841 nor n14022 n14032 ; n14033
g13842 and asqrt[62] n14033_not ; n14034
g13843 and n13450_not n13457 ; n14035
g13844 and n13459_not n14035 ; n14036
g13845 and asqrt[17] n14036 ; n14037
g13846 nor n13450 n13459 ; n14038
g13847 and asqrt[17] n14038 ; n14039
g13848 nor n13457 n14039 ; n14040
g13849 nor n14037 n14040 ; n14041
g13850 nor asqrt[62] n14022 ; n14042
g13851 and n14032_not n14042 ; n14043
g13852 nor n14041 n14043 ; n14044
g13853 nor n14034 n14044 ; n14045
g13854 and n13469 n13471_not ; n14046
g13855 and n13462_not n14046 ; n14047
g13856 and asqrt[17] n14047 ; n14048
g13857 nor n13462 n13471 ; n14049
g13858 and asqrt[17] n14049 ; n14050
g13859 nor n13469 n14050 ; n14051
g13860 nor n14048 n14051 ; n14052
g13861 nor n13473 n13480 ; n14053
g13862 and asqrt[17] n14053 ; n14054
g13863 nor n13488 n14054 ; n14055
g13864 and n14052_not n14055 ; n14056
g13865 and n14045_not n14056 ; n14057
g13866 nor asqrt[63] n14057 ; n14058
g13867 and n14034_not n14052 ; n14059
g13868 and n14044_not n14059 ; n14060
g13869 and n13480_not asqrt[17] ; n14061
g13870 and n13473 n14061_not ; n14062
g13871 and asqrt[63] n14053_not ; n14063
g13872 and n14062_not n14063 ; n14064
g13873 nor n13476 n13497 ; n14065
g13874 and n13479_not n14065 ; n14066
g13875 and n13492_not n14066 ; n14067
g13876 and n13488_not n14067 ; n14068
g13877 and n13486_not n14068 ; n14069
g13878 nor n14064 n14069 ; n14070
g13879 and n14060_not n14070 ; n14071
g13880 nand n14058_not n14071 ; asqrt[16]
g13881 and a[32] asqrt[16] ; n14073
g13882 nor a[30] a[31] ; n14074
g13883 and a[32]_not n14074 ; n14075
g13884 nor n14073 n14075 ; n14076
g13885 and asqrt[17] n14076_not ; n14077
g13886 nor n13497 n14075 ; n14078
g13887 and n13492_not n14078 ; n14079
g13888 and n13488_not n14079 ; n14080
g13889 and n13486_not n14080 ; n14081
g13890 and n14073_not n14081 ; n14082
g13891 and a[32]_not asqrt[16] ; n14083
g13892 and a[33] n14083_not ; n14084
g13893 and n13502 asqrt[16] ; n14085
g13894 nor n14084 n14085 ; n14086
g13895 and n14082_not n14086 ; n14087
g13896 nor n14077 n14087 ; n14088
g13897 and asqrt[18] n14088_not ; n14089
g13898 nor asqrt[18] n14077 ; n14090
g13899 and n14087_not n14090 ; n14091
g13900 and asqrt[17] n14069_not ; n14092
g13901 and n14064_not n14092 ; n14093
g13902 and n14060_not n14093 ; n14094
g13903 and n14058_not n14094 ; n14095
g13904 nor n14085 n14095 ; n14096
g13905 and a[34] n14096_not ; n14097
g13906 nor a[34] n14095 ; n14098
g13907 and n14085_not n14098 ; n14099
g13908 nor n14097 n14099 ; n14100
g13909 nor n14091 n14100 ; n14101
g13910 nor n14089 n14101 ; n14102
g13911 and asqrt[19] n14102_not ; n14103
g13912 nor n13505 n13510 ; n14104
g13913 and n13514_not n14104 ; n14105
g13914 and asqrt[16] n14105 ; n14106
g13915 and asqrt[16] n14104 ; n14107
g13916 and n13514 n14107_not ; n14108
g13917 nor n14106 n14108 ; n14109
g13918 nor asqrt[19] n14089 ; n14110
g13919 and n14101_not n14110 ; n14111
g13920 nor n14109 n14111 ; n14112
g13921 nor n14103 n14112 ; n14113
g13922 and asqrt[20] n14113_not ; n14114
g13923 and n13519_not n13528 ; n14115
g13924 and n13517_not n14115 ; n14116
g13925 and asqrt[16] n14116 ; n14117
g13926 nor n13517 n13519 ; n14118
g13927 and asqrt[16] n14118 ; n14119
g13928 nor n13528 n14119 ; n14120
g13929 nor n14117 n14120 ; n14121
g13930 nor asqrt[20] n14103 ; n14122
g13931 and n14112_not n14122 ; n14123
g13932 nor n14121 n14123 ; n14124
g13933 nor n14114 n14124 ; n14125
g13934 and asqrt[21] n14125_not ; n14126
g13935 and n13531_not n13537 ; n14127
g13936 and n13539_not n14127 ; n14128
g13937 and asqrt[16] n14128 ; n14129
g13938 nor n13531 n13539 ; n14130
g13939 and asqrt[16] n14130 ; n14131
g13940 nor n13537 n14131 ; n14132
g13941 nor n14129 n14132 ; n14133
g13942 nor asqrt[21] n14114 ; n14134
g13943 and n14124_not n14134 ; n14135
g13944 nor n14133 n14135 ; n14136
g13945 nor n14126 n14136 ; n14137
g13946 and asqrt[22] n14137_not ; n14138
g13947 and n13549 n13551_not ; n14139
g13948 and n13542_not n14139 ; n14140
g13949 and asqrt[16] n14140 ; n14141
g13950 nor n13542 n13551 ; n14142
g13951 and asqrt[16] n14142 ; n14143
g13952 nor n13549 n14143 ; n14144
g13953 nor n14141 n14144 ; n14145
g13954 nor asqrt[22] n14126 ; n14146
g13955 and n14136_not n14146 ; n14147
g13956 nor n14145 n14147 ; n14148
g13957 nor n14138 n14148 ; n14149
g13958 and asqrt[23] n14149_not ; n14150
g13959 and n13554_not n13561 ; n14151
g13960 and n13563_not n14151 ; n14152
g13961 and asqrt[16] n14152 ; n14153
g13962 nor n13554 n13563 ; n14154
g13963 and asqrt[16] n14154 ; n14155
g13964 nor n13561 n14155 ; n14156
g13965 nor n14153 n14156 ; n14157
g13966 nor asqrt[23] n14138 ; n14158
g13967 and n14148_not n14158 ; n14159
g13968 nor n14157 n14159 ; n14160
g13969 nor n14150 n14160 ; n14161
g13970 and asqrt[24] n14161_not ; n14162
g13971 and n13573 n13575_not ; n14163
g13972 and n13566_not n14163 ; n14164
g13973 and asqrt[16] n14164 ; n14165
g13974 nor n13566 n13575 ; n14166
g13975 and asqrt[16] n14166 ; n14167
g13976 nor n13573 n14167 ; n14168
g13977 nor n14165 n14168 ; n14169
g13978 nor asqrt[24] n14150 ; n14170
g13979 and n14160_not n14170 ; n14171
g13980 nor n14169 n14171 ; n14172
g13981 nor n14162 n14172 ; n14173
g13982 and asqrt[25] n14173_not ; n14174
g13983 and n13578_not n13585 ; n14175
g13984 and n13587_not n14175 ; n14176
g13985 and asqrt[16] n14176 ; n14177
g13986 nor n13578 n13587 ; n14178
g13987 and asqrt[16] n14178 ; n14179
g13988 nor n13585 n14179 ; n14180
g13989 nor n14177 n14180 ; n14181
g13990 nor asqrt[25] n14162 ; n14182
g13991 and n14172_not n14182 ; n14183
g13992 nor n14181 n14183 ; n14184
g13993 nor n14174 n14184 ; n14185
g13994 and asqrt[26] n14185_not ; n14186
g13995 and n13597 n13599_not ; n14187
g13996 and n13590_not n14187 ; n14188
g13997 and asqrt[16] n14188 ; n14189
g13998 nor n13590 n13599 ; n14190
g13999 and asqrt[16] n14190 ; n14191
g14000 nor n13597 n14191 ; n14192
g14001 nor n14189 n14192 ; n14193
g14002 nor asqrt[26] n14174 ; n14194
g14003 and n14184_not n14194 ; n14195
g14004 nor n14193 n14195 ; n14196
g14005 nor n14186 n14196 ; n14197
g14006 and asqrt[27] n14197_not ; n14198
g14007 and n13602_not n13609 ; n14199
g14008 and n13611_not n14199 ; n14200
g14009 and asqrt[16] n14200 ; n14201
g14010 nor n13602 n13611 ; n14202
g14011 and asqrt[16] n14202 ; n14203
g14012 nor n13609 n14203 ; n14204
g14013 nor n14201 n14204 ; n14205
g14014 nor asqrt[27] n14186 ; n14206
g14015 and n14196_not n14206 ; n14207
g14016 nor n14205 n14207 ; n14208
g14017 nor n14198 n14208 ; n14209
g14018 and asqrt[28] n14209_not ; n14210
g14019 and n13621 n13623_not ; n14211
g14020 and n13614_not n14211 ; n14212
g14021 and asqrt[16] n14212 ; n14213
g14022 nor n13614 n13623 ; n14214
g14023 and asqrt[16] n14214 ; n14215
g14024 nor n13621 n14215 ; n14216
g14025 nor n14213 n14216 ; n14217
g14026 nor asqrt[28] n14198 ; n14218
g14027 and n14208_not n14218 ; n14219
g14028 nor n14217 n14219 ; n14220
g14029 nor n14210 n14220 ; n14221
g14030 and asqrt[29] n14221_not ; n14222
g14031 and n13626_not n13633 ; n14223
g14032 and n13635_not n14223 ; n14224
g14033 and asqrt[16] n14224 ; n14225
g14034 nor n13626 n13635 ; n14226
g14035 and asqrt[16] n14226 ; n14227
g14036 nor n13633 n14227 ; n14228
g14037 nor n14225 n14228 ; n14229
g14038 nor asqrt[29] n14210 ; n14230
g14039 and n14220_not n14230 ; n14231
g14040 nor n14229 n14231 ; n14232
g14041 nor n14222 n14232 ; n14233
g14042 and asqrt[30] n14233_not ; n14234
g14043 and n13645 n13647_not ; n14235
g14044 and n13638_not n14235 ; n14236
g14045 and asqrt[16] n14236 ; n14237
g14046 nor n13638 n13647 ; n14238
g14047 and asqrt[16] n14238 ; n14239
g14048 nor n13645 n14239 ; n14240
g14049 nor n14237 n14240 ; n14241
g14050 nor asqrt[30] n14222 ; n14242
g14051 and n14232_not n14242 ; n14243
g14052 nor n14241 n14243 ; n14244
g14053 nor n14234 n14244 ; n14245
g14054 and asqrt[31] n14245_not ; n14246
g14055 and n13650_not n13657 ; n14247
g14056 and n13659_not n14247 ; n14248
g14057 and asqrt[16] n14248 ; n14249
g14058 nor n13650 n13659 ; n14250
g14059 and asqrt[16] n14250 ; n14251
g14060 nor n13657 n14251 ; n14252
g14061 nor n14249 n14252 ; n14253
g14062 nor asqrt[31] n14234 ; n14254
g14063 and n14244_not n14254 ; n14255
g14064 nor n14253 n14255 ; n14256
g14065 nor n14246 n14256 ; n14257
g14066 and asqrt[32] n14257_not ; n14258
g14067 and n13669 n13671_not ; n14259
g14068 and n13662_not n14259 ; n14260
g14069 and asqrt[16] n14260 ; n14261
g14070 nor n13662 n13671 ; n14262
g14071 and asqrt[16] n14262 ; n14263
g14072 nor n13669 n14263 ; n14264
g14073 nor n14261 n14264 ; n14265
g14074 nor asqrt[32] n14246 ; n14266
g14075 and n14256_not n14266 ; n14267
g14076 nor n14265 n14267 ; n14268
g14077 nor n14258 n14268 ; n14269
g14078 and asqrt[33] n14269_not ; n14270
g14079 and n13674_not n13681 ; n14271
g14080 and n13683_not n14271 ; n14272
g14081 and asqrt[16] n14272 ; n14273
g14082 nor n13674 n13683 ; n14274
g14083 and asqrt[16] n14274 ; n14275
g14084 nor n13681 n14275 ; n14276
g14085 nor n14273 n14276 ; n14277
g14086 nor asqrt[33] n14258 ; n14278
g14087 and n14268_not n14278 ; n14279
g14088 nor n14277 n14279 ; n14280
g14089 nor n14270 n14280 ; n14281
g14090 and asqrt[34] n14281_not ; n14282
g14091 and n13693 n13695_not ; n14283
g14092 and n13686_not n14283 ; n14284
g14093 and asqrt[16] n14284 ; n14285
g14094 nor n13686 n13695 ; n14286
g14095 and asqrt[16] n14286 ; n14287
g14096 nor n13693 n14287 ; n14288
g14097 nor n14285 n14288 ; n14289
g14098 nor asqrt[34] n14270 ; n14290
g14099 and n14280_not n14290 ; n14291
g14100 nor n14289 n14291 ; n14292
g14101 nor n14282 n14292 ; n14293
g14102 and asqrt[35] n14293_not ; n14294
g14103 and n13698_not n13705 ; n14295
g14104 and n13707_not n14295 ; n14296
g14105 and asqrt[16] n14296 ; n14297
g14106 nor n13698 n13707 ; n14298
g14107 and asqrt[16] n14298 ; n14299
g14108 nor n13705 n14299 ; n14300
g14109 nor n14297 n14300 ; n14301
g14110 nor asqrt[35] n14282 ; n14302
g14111 and n14292_not n14302 ; n14303
g14112 nor n14301 n14303 ; n14304
g14113 nor n14294 n14304 ; n14305
g14114 and asqrt[36] n14305_not ; n14306
g14115 and n13717 n13719_not ; n14307
g14116 and n13710_not n14307 ; n14308
g14117 and asqrt[16] n14308 ; n14309
g14118 nor n13710 n13719 ; n14310
g14119 and asqrt[16] n14310 ; n14311
g14120 nor n13717 n14311 ; n14312
g14121 nor n14309 n14312 ; n14313
g14122 nor asqrt[36] n14294 ; n14314
g14123 and n14304_not n14314 ; n14315
g14124 nor n14313 n14315 ; n14316
g14125 nor n14306 n14316 ; n14317
g14126 and asqrt[37] n14317_not ; n14318
g14127 and n13722_not n13729 ; n14319
g14128 and n13731_not n14319 ; n14320
g14129 and asqrt[16] n14320 ; n14321
g14130 nor n13722 n13731 ; n14322
g14131 and asqrt[16] n14322 ; n14323
g14132 nor n13729 n14323 ; n14324
g14133 nor n14321 n14324 ; n14325
g14134 nor asqrt[37] n14306 ; n14326
g14135 and n14316_not n14326 ; n14327
g14136 nor n14325 n14327 ; n14328
g14137 nor n14318 n14328 ; n14329
g14138 and asqrt[38] n14329_not ; n14330
g14139 and n13741 n13743_not ; n14331
g14140 and n13734_not n14331 ; n14332
g14141 and asqrt[16] n14332 ; n14333
g14142 nor n13734 n13743 ; n14334
g14143 and asqrt[16] n14334 ; n14335
g14144 nor n13741 n14335 ; n14336
g14145 nor n14333 n14336 ; n14337
g14146 nor asqrt[38] n14318 ; n14338
g14147 and n14328_not n14338 ; n14339
g14148 nor n14337 n14339 ; n14340
g14149 nor n14330 n14340 ; n14341
g14150 and asqrt[39] n14341_not ; n14342
g14151 and n13746_not n13753 ; n14343
g14152 and n13755_not n14343 ; n14344
g14153 and asqrt[16] n14344 ; n14345
g14154 nor n13746 n13755 ; n14346
g14155 and asqrt[16] n14346 ; n14347
g14156 nor n13753 n14347 ; n14348
g14157 nor n14345 n14348 ; n14349
g14158 nor asqrt[39] n14330 ; n14350
g14159 and n14340_not n14350 ; n14351
g14160 nor n14349 n14351 ; n14352
g14161 nor n14342 n14352 ; n14353
g14162 and asqrt[40] n14353_not ; n14354
g14163 and n13765 n13767_not ; n14355
g14164 and n13758_not n14355 ; n14356
g14165 and asqrt[16] n14356 ; n14357
g14166 nor n13758 n13767 ; n14358
g14167 and asqrt[16] n14358 ; n14359
g14168 nor n13765 n14359 ; n14360
g14169 nor n14357 n14360 ; n14361
g14170 nor asqrt[40] n14342 ; n14362
g14171 and n14352_not n14362 ; n14363
g14172 nor n14361 n14363 ; n14364
g14173 nor n14354 n14364 ; n14365
g14174 and asqrt[41] n14365_not ; n14366
g14175 and n13770_not n13777 ; n14367
g14176 and n13779_not n14367 ; n14368
g14177 and asqrt[16] n14368 ; n14369
g14178 nor n13770 n13779 ; n14370
g14179 and asqrt[16] n14370 ; n14371
g14180 nor n13777 n14371 ; n14372
g14181 nor n14369 n14372 ; n14373
g14182 nor asqrt[41] n14354 ; n14374
g14183 and n14364_not n14374 ; n14375
g14184 nor n14373 n14375 ; n14376
g14185 nor n14366 n14376 ; n14377
g14186 and asqrt[42] n14377_not ; n14378
g14187 and n13789 n13791_not ; n14379
g14188 and n13782_not n14379 ; n14380
g14189 and asqrt[16] n14380 ; n14381
g14190 nor n13782 n13791 ; n14382
g14191 and asqrt[16] n14382 ; n14383
g14192 nor n13789 n14383 ; n14384
g14193 nor n14381 n14384 ; n14385
g14194 nor asqrt[42] n14366 ; n14386
g14195 and n14376_not n14386 ; n14387
g14196 nor n14385 n14387 ; n14388
g14197 nor n14378 n14388 ; n14389
g14198 and asqrt[43] n14389_not ; n14390
g14199 and n13794_not n13801 ; n14391
g14200 and n13803_not n14391 ; n14392
g14201 and asqrt[16] n14392 ; n14393
g14202 nor n13794 n13803 ; n14394
g14203 and asqrt[16] n14394 ; n14395
g14204 nor n13801 n14395 ; n14396
g14205 nor n14393 n14396 ; n14397
g14206 nor asqrt[43] n14378 ; n14398
g14207 and n14388_not n14398 ; n14399
g14208 nor n14397 n14399 ; n14400
g14209 nor n14390 n14400 ; n14401
g14210 and asqrt[44] n14401_not ; n14402
g14211 and n13813 n13815_not ; n14403
g14212 and n13806_not n14403 ; n14404
g14213 and asqrt[16] n14404 ; n14405
g14214 nor n13806 n13815 ; n14406
g14215 and asqrt[16] n14406 ; n14407
g14216 nor n13813 n14407 ; n14408
g14217 nor n14405 n14408 ; n14409
g14218 nor asqrt[44] n14390 ; n14410
g14219 and n14400_not n14410 ; n14411
g14220 nor n14409 n14411 ; n14412
g14221 nor n14402 n14412 ; n14413
g14222 and asqrt[45] n14413_not ; n14414
g14223 and n13818_not n13825 ; n14415
g14224 and n13827_not n14415 ; n14416
g14225 and asqrt[16] n14416 ; n14417
g14226 nor n13818 n13827 ; n14418
g14227 and asqrt[16] n14418 ; n14419
g14228 nor n13825 n14419 ; n14420
g14229 nor n14417 n14420 ; n14421
g14230 nor asqrt[45] n14402 ; n14422
g14231 and n14412_not n14422 ; n14423
g14232 nor n14421 n14423 ; n14424
g14233 nor n14414 n14424 ; n14425
g14234 and asqrt[46] n14425_not ; n14426
g14235 and n13837 n13839_not ; n14427
g14236 and n13830_not n14427 ; n14428
g14237 and asqrt[16] n14428 ; n14429
g14238 nor n13830 n13839 ; n14430
g14239 and asqrt[16] n14430 ; n14431
g14240 nor n13837 n14431 ; n14432
g14241 nor n14429 n14432 ; n14433
g14242 nor asqrt[46] n14414 ; n14434
g14243 and n14424_not n14434 ; n14435
g14244 nor n14433 n14435 ; n14436
g14245 nor n14426 n14436 ; n14437
g14246 and asqrt[47] n14437_not ; n14438
g14247 and n13842_not n13849 ; n14439
g14248 and n13851_not n14439 ; n14440
g14249 and asqrt[16] n14440 ; n14441
g14250 nor n13842 n13851 ; n14442
g14251 and asqrt[16] n14442 ; n14443
g14252 nor n13849 n14443 ; n14444
g14253 nor n14441 n14444 ; n14445
g14254 nor asqrt[47] n14426 ; n14446
g14255 and n14436_not n14446 ; n14447
g14256 nor n14445 n14447 ; n14448
g14257 nor n14438 n14448 ; n14449
g14258 and asqrt[48] n14449_not ; n14450
g14259 and n13861 n13863_not ; n14451
g14260 and n13854_not n14451 ; n14452
g14261 and asqrt[16] n14452 ; n14453
g14262 nor n13854 n13863 ; n14454
g14263 and asqrt[16] n14454 ; n14455
g14264 nor n13861 n14455 ; n14456
g14265 nor n14453 n14456 ; n14457
g14266 nor asqrt[48] n14438 ; n14458
g14267 and n14448_not n14458 ; n14459
g14268 nor n14457 n14459 ; n14460
g14269 nor n14450 n14460 ; n14461
g14270 and asqrt[49] n14461_not ; n14462
g14271 nor asqrt[49] n14450 ; n14463
g14272 and n14460_not n14463 ; n14464
g14273 and n13866_not n13875 ; n14465
g14274 and n13868_not n14465 ; n14466
g14275 and asqrt[16] n14466 ; n14467
g14276 nor n13866 n13868 ; n14468
g14277 and asqrt[16] n14468 ; n14469
g14278 nor n13875 n14469 ; n14470
g14279 nor n14467 n14470 ; n14471
g14280 nor n14464 n14471 ; n14472
g14281 nor n14462 n14472 ; n14473
g14282 and asqrt[50] n14473_not ; n14474
g14283 and n13885 n13887_not ; n14475
g14284 and n13878_not n14475 ; n14476
g14285 and asqrt[16] n14476 ; n14477
g14286 nor n13878 n13887 ; n14478
g14287 and asqrt[16] n14478 ; n14479
g14288 nor n13885 n14479 ; n14480
g14289 nor n14477 n14480 ; n14481
g14290 nor asqrt[50] n14462 ; n14482
g14291 and n14472_not n14482 ; n14483
g14292 nor n14481 n14483 ; n14484
g14293 nor n14474 n14484 ; n14485
g14294 and asqrt[51] n14485_not ; n14486
g14295 and n13890_not n13897 ; n14487
g14296 and n13899_not n14487 ; n14488
g14297 and asqrt[16] n14488 ; n14489
g14298 nor n13890 n13899 ; n14490
g14299 and asqrt[16] n14490 ; n14491
g14300 nor n13897 n14491 ; n14492
g14301 nor n14489 n14492 ; n14493
g14302 nor asqrt[51] n14474 ; n14494
g14303 and n14484_not n14494 ; n14495
g14304 nor n14493 n14495 ; n14496
g14305 nor n14486 n14496 ; n14497
g14306 and asqrt[52] n14497_not ; n14498
g14307 and n13909 n13911_not ; n14499
g14308 and n13902_not n14499 ; n14500
g14309 and asqrt[16] n14500 ; n14501
g14310 nor n13902 n13911 ; n14502
g14311 and asqrt[16] n14502 ; n14503
g14312 nor n13909 n14503 ; n14504
g14313 nor n14501 n14504 ; n14505
g14314 nor asqrt[52] n14486 ; n14506
g14315 and n14496_not n14506 ; n14507
g14316 nor n14505 n14507 ; n14508
g14317 nor n14498 n14508 ; n14509
g14318 and asqrt[53] n14509_not ; n14510
g14319 and n13914_not n13921 ; n14511
g14320 and n13923_not n14511 ; n14512
g14321 and asqrt[16] n14512 ; n14513
g14322 nor n13914 n13923 ; n14514
g14323 and asqrt[16] n14514 ; n14515
g14324 nor n13921 n14515 ; n14516
g14325 nor n14513 n14516 ; n14517
g14326 nor asqrt[53] n14498 ; n14518
g14327 and n14508_not n14518 ; n14519
g14328 nor n14517 n14519 ; n14520
g14329 nor n14510 n14520 ; n14521
g14330 and asqrt[54] n14521_not ; n14522
g14331 and n13933 n13935_not ; n14523
g14332 and n13926_not n14523 ; n14524
g14333 and asqrt[16] n14524 ; n14525
g14334 nor n13926 n13935 ; n14526
g14335 and asqrt[16] n14526 ; n14527
g14336 nor n13933 n14527 ; n14528
g14337 nor n14525 n14528 ; n14529
g14338 nor asqrt[54] n14510 ; n14530
g14339 and n14520_not n14530 ; n14531
g14340 nor n14529 n14531 ; n14532
g14341 nor n14522 n14532 ; n14533
g14342 and asqrt[55] n14533_not ; n14534
g14343 and n13938_not n13945 ; n14535
g14344 and n13947_not n14535 ; n14536
g14345 and asqrt[16] n14536 ; n14537
g14346 nor n13938 n13947 ; n14538
g14347 and asqrt[16] n14538 ; n14539
g14348 nor n13945 n14539 ; n14540
g14349 nor n14537 n14540 ; n14541
g14350 nor asqrt[55] n14522 ; n14542
g14351 and n14532_not n14542 ; n14543
g14352 nor n14541 n14543 ; n14544
g14353 nor n14534 n14544 ; n14545
g14354 and asqrt[56] n14545_not ; n14546
g14355 and n13957 n13959_not ; n14547
g14356 and n13950_not n14547 ; n14548
g14357 and asqrt[16] n14548 ; n14549
g14358 nor n13950 n13959 ; n14550
g14359 and asqrt[16] n14550 ; n14551
g14360 nor n13957 n14551 ; n14552
g14361 nor n14549 n14552 ; n14553
g14362 nor asqrt[56] n14534 ; n14554
g14363 and n14544_not n14554 ; n14555
g14364 nor n14553 n14555 ; n14556
g14365 nor n14546 n14556 ; n14557
g14366 and asqrt[57] n14557_not ; n14558
g14367 and n13962_not n13969 ; n14559
g14368 and n13971_not n14559 ; n14560
g14369 and asqrt[16] n14560 ; n14561
g14370 nor n13962 n13971 ; n14562
g14371 and asqrt[16] n14562 ; n14563
g14372 nor n13969 n14563 ; n14564
g14373 nor n14561 n14564 ; n14565
g14374 nor asqrt[57] n14546 ; n14566
g14375 and n14556_not n14566 ; n14567
g14376 nor n14565 n14567 ; n14568
g14377 nor n14558 n14568 ; n14569
g14378 and asqrt[58] n14569_not ; n14570
g14379 and n13981 n13983_not ; n14571
g14380 and n13974_not n14571 ; n14572
g14381 and asqrt[16] n14572 ; n14573
g14382 nor n13974 n13983 ; n14574
g14383 and asqrt[16] n14574 ; n14575
g14384 nor n13981 n14575 ; n14576
g14385 nor n14573 n14576 ; n14577
g14386 nor asqrt[58] n14558 ; n14578
g14387 and n14568_not n14578 ; n14579
g14388 nor n14577 n14579 ; n14580
g14389 nor n14570 n14580 ; n14581
g14390 and asqrt[59] n14581_not ; n14582
g14391 and n13986_not n13993 ; n14583
g14392 and n13995_not n14583 ; n14584
g14393 and asqrt[16] n14584 ; n14585
g14394 nor n13986 n13995 ; n14586
g14395 and asqrt[16] n14586 ; n14587
g14396 nor n13993 n14587 ; n14588
g14397 nor n14585 n14588 ; n14589
g14398 nor asqrt[59] n14570 ; n14590
g14399 and n14580_not n14590 ; n14591
g14400 nor n14589 n14591 ; n14592
g14401 nor n14582 n14592 ; n14593
g14402 and asqrt[60] n14593_not ; n14594
g14403 and n14005 n14007_not ; n14595
g14404 and n13998_not n14595 ; n14596
g14405 and asqrt[16] n14596 ; n14597
g14406 nor n13998 n14007 ; n14598
g14407 and asqrt[16] n14598 ; n14599
g14408 nor n14005 n14599 ; n14600
g14409 nor n14597 n14600 ; n14601
g14410 nor asqrt[60] n14582 ; n14602
g14411 and n14592_not n14602 ; n14603
g14412 nor n14601 n14603 ; n14604
g14413 nor n14594 n14604 ; n14605
g14414 and asqrt[61] n14605_not ; n14606
g14415 and n14010_not n14017 ; n14607
g14416 and n14019_not n14607 ; n14608
g14417 and asqrt[16] n14608 ; n14609
g14418 nor n14010 n14019 ; n14610
g14419 and asqrt[16] n14610 ; n14611
g14420 nor n14017 n14611 ; n14612
g14421 nor n14609 n14612 ; n14613
g14422 nor asqrt[61] n14594 ; n14614
g14423 and n14604_not n14614 ; n14615
g14424 nor n14613 n14615 ; n14616
g14425 nor n14606 n14616 ; n14617
g14426 and asqrt[62] n14617_not ; n14618
g14427 and n14029 n14031_not ; n14619
g14428 and n14022_not n14619 ; n14620
g14429 and asqrt[16] n14620 ; n14621
g14430 nor n14022 n14031 ; n14622
g14431 and asqrt[16] n14622 ; n14623
g14432 nor n14029 n14623 ; n14624
g14433 nor n14621 n14624 ; n14625
g14434 nor asqrt[62] n14606 ; n14626
g14435 and n14616_not n14626 ; n14627
g14436 nor n14625 n14627 ; n14628
g14437 nor n14618 n14628 ; n14629
g14438 and n14034_not n14041 ; n14630
g14439 and n14043_not n14630 ; n14631
g14440 and asqrt[16] n14631 ; n14632
g14441 nor n14034 n14043 ; n14633
g14442 and asqrt[16] n14633 ; n14634
g14443 nor n14041 n14634 ; n14635
g14444 nor n14632 n14635 ; n14636
g14445 nor n14045 n14052 ; n14637
g14446 and asqrt[16] n14637 ; n14638
g14447 nor n14060 n14638 ; n14639
g14448 and n14636_not n14639 ; n14640
g14449 and n14629_not n14640 ; n14641
g14450 nor asqrt[63] n14641 ; n14642
g14451 and n14618_not n14636 ; n14643
g14452 and n14628_not n14643 ; n14644
g14453 and n14052_not asqrt[16] ; n14645
g14454 and n14045 n14645_not ; n14646
g14455 and asqrt[63] n14637_not ; n14647
g14456 and n14646_not n14647 ; n14648
g14457 nor n14048 n14069 ; n14649
g14458 and n14051_not n14649 ; n14650
g14459 and n14064_not n14650 ; n14651
g14460 and n14060_not n14651 ; n14652
g14461 and n14058_not n14652 ; n14653
g14462 nor n14648 n14653 ; n14654
g14463 and n14644_not n14654 ; n14655
g14464 nand n14642_not n14655 ; asqrt[15]
g14465 and a[30] asqrt[15] ; n14657
g14466 nor a[28] a[29] ; n14658
g14467 and a[30]_not n14658 ; n14659
g14468 nor n14657 n14659 ; n14660
g14469 and asqrt[16] n14660_not ; n14661
g14470 nor n14069 n14659 ; n14662
g14471 and n14064_not n14662 ; n14663
g14472 and n14060_not n14663 ; n14664
g14473 and n14058_not n14664 ; n14665
g14474 and n14657_not n14665 ; n14666
g14475 and a[30]_not asqrt[15] ; n14667
g14476 and a[31] n14667_not ; n14668
g14477 and n14074 asqrt[15] ; n14669
g14478 nor n14668 n14669 ; n14670
g14479 and n14666_not n14670 ; n14671
g14480 nor n14661 n14671 ; n14672
g14481 and asqrt[17] n14672_not ; n14673
g14482 nor asqrt[17] n14661 ; n14674
g14483 and n14671_not n14674 ; n14675
g14484 and asqrt[16] n14653_not ; n14676
g14485 and n14648_not n14676 ; n14677
g14486 and n14644_not n14677 ; n14678
g14487 and n14642_not n14678 ; n14679
g14488 nor n14669 n14679 ; n14680
g14489 and a[32] n14680_not ; n14681
g14490 nor a[32] n14679 ; n14682
g14491 and n14669_not n14682 ; n14683
g14492 nor n14681 n14683 ; n14684
g14493 nor n14675 n14684 ; n14685
g14494 nor n14673 n14685 ; n14686
g14495 and asqrt[18] n14686_not ; n14687
g14496 nor n14077 n14082 ; n14688
g14497 and n14086_not n14688 ; n14689
g14498 and asqrt[15] n14689 ; n14690
g14499 and asqrt[15] n14688 ; n14691
g14500 and n14086 n14691_not ; n14692
g14501 nor n14690 n14692 ; n14693
g14502 nor asqrt[18] n14673 ; n14694
g14503 and n14685_not n14694 ; n14695
g14504 nor n14693 n14695 ; n14696
g14505 nor n14687 n14696 ; n14697
g14506 and asqrt[19] n14697_not ; n14698
g14507 and n14091_not n14100 ; n14699
g14508 and n14089_not n14699 ; n14700
g14509 and asqrt[15] n14700 ; n14701
g14510 nor n14089 n14091 ; n14702
g14511 and asqrt[15] n14702 ; n14703
g14512 nor n14100 n14703 ; n14704
g14513 nor n14701 n14704 ; n14705
g14514 nor asqrt[19] n14687 ; n14706
g14515 and n14696_not n14706 ; n14707
g14516 nor n14705 n14707 ; n14708
g14517 nor n14698 n14708 ; n14709
g14518 and asqrt[20] n14709_not ; n14710
g14519 and n14103_not n14109 ; n14711
g14520 and n14111_not n14711 ; n14712
g14521 and asqrt[15] n14712 ; n14713
g14522 nor n14103 n14111 ; n14714
g14523 and asqrt[15] n14714 ; n14715
g14524 nor n14109 n14715 ; n14716
g14525 nor n14713 n14716 ; n14717
g14526 nor asqrt[20] n14698 ; n14718
g14527 and n14708_not n14718 ; n14719
g14528 nor n14717 n14719 ; n14720
g14529 nor n14710 n14720 ; n14721
g14530 and asqrt[21] n14721_not ; n14722
g14531 and n14121 n14123_not ; n14723
g14532 and n14114_not n14723 ; n14724
g14533 and asqrt[15] n14724 ; n14725
g14534 nor n14114 n14123 ; n14726
g14535 and asqrt[15] n14726 ; n14727
g14536 nor n14121 n14727 ; n14728
g14537 nor n14725 n14728 ; n14729
g14538 nor asqrt[21] n14710 ; n14730
g14539 and n14720_not n14730 ; n14731
g14540 nor n14729 n14731 ; n14732
g14541 nor n14722 n14732 ; n14733
g14542 and asqrt[22] n14733_not ; n14734
g14543 and n14126_not n14133 ; n14735
g14544 and n14135_not n14735 ; n14736
g14545 and asqrt[15] n14736 ; n14737
g14546 nor n14126 n14135 ; n14738
g14547 and asqrt[15] n14738 ; n14739
g14548 nor n14133 n14739 ; n14740
g14549 nor n14737 n14740 ; n14741
g14550 nor asqrt[22] n14722 ; n14742
g14551 and n14732_not n14742 ; n14743
g14552 nor n14741 n14743 ; n14744
g14553 nor n14734 n14744 ; n14745
g14554 and asqrt[23] n14745_not ; n14746
g14555 and n14145 n14147_not ; n14747
g14556 and n14138_not n14747 ; n14748
g14557 and asqrt[15] n14748 ; n14749
g14558 nor n14138 n14147 ; n14750
g14559 and asqrt[15] n14750 ; n14751
g14560 nor n14145 n14751 ; n14752
g14561 nor n14749 n14752 ; n14753
g14562 nor asqrt[23] n14734 ; n14754
g14563 and n14744_not n14754 ; n14755
g14564 nor n14753 n14755 ; n14756
g14565 nor n14746 n14756 ; n14757
g14566 and asqrt[24] n14757_not ; n14758
g14567 and n14150_not n14157 ; n14759
g14568 and n14159_not n14759 ; n14760
g14569 and asqrt[15] n14760 ; n14761
g14570 nor n14150 n14159 ; n14762
g14571 and asqrt[15] n14762 ; n14763
g14572 nor n14157 n14763 ; n14764
g14573 nor n14761 n14764 ; n14765
g14574 nor asqrt[24] n14746 ; n14766
g14575 and n14756_not n14766 ; n14767
g14576 nor n14765 n14767 ; n14768
g14577 nor n14758 n14768 ; n14769
g14578 and asqrt[25] n14769_not ; n14770
g14579 and n14169 n14171_not ; n14771
g14580 and n14162_not n14771 ; n14772
g14581 and asqrt[15] n14772 ; n14773
g14582 nor n14162 n14171 ; n14774
g14583 and asqrt[15] n14774 ; n14775
g14584 nor n14169 n14775 ; n14776
g14585 nor n14773 n14776 ; n14777
g14586 nor asqrt[25] n14758 ; n14778
g14587 and n14768_not n14778 ; n14779
g14588 nor n14777 n14779 ; n14780
g14589 nor n14770 n14780 ; n14781
g14590 and asqrt[26] n14781_not ; n14782
g14591 and n14174_not n14181 ; n14783
g14592 and n14183_not n14783 ; n14784
g14593 and asqrt[15] n14784 ; n14785
g14594 nor n14174 n14183 ; n14786
g14595 and asqrt[15] n14786 ; n14787
g14596 nor n14181 n14787 ; n14788
g14597 nor n14785 n14788 ; n14789
g14598 nor asqrt[26] n14770 ; n14790
g14599 and n14780_not n14790 ; n14791
g14600 nor n14789 n14791 ; n14792
g14601 nor n14782 n14792 ; n14793
g14602 and asqrt[27] n14793_not ; n14794
g14603 and n14193 n14195_not ; n14795
g14604 and n14186_not n14795 ; n14796
g14605 and asqrt[15] n14796 ; n14797
g14606 nor n14186 n14195 ; n14798
g14607 and asqrt[15] n14798 ; n14799
g14608 nor n14193 n14799 ; n14800
g14609 nor n14797 n14800 ; n14801
g14610 nor asqrt[27] n14782 ; n14802
g14611 and n14792_not n14802 ; n14803
g14612 nor n14801 n14803 ; n14804
g14613 nor n14794 n14804 ; n14805
g14614 and asqrt[28] n14805_not ; n14806
g14615 and n14198_not n14205 ; n14807
g14616 and n14207_not n14807 ; n14808
g14617 and asqrt[15] n14808 ; n14809
g14618 nor n14198 n14207 ; n14810
g14619 and asqrt[15] n14810 ; n14811
g14620 nor n14205 n14811 ; n14812
g14621 nor n14809 n14812 ; n14813
g14622 nor asqrt[28] n14794 ; n14814
g14623 and n14804_not n14814 ; n14815
g14624 nor n14813 n14815 ; n14816
g14625 nor n14806 n14816 ; n14817
g14626 and asqrt[29] n14817_not ; n14818
g14627 and n14217 n14219_not ; n14819
g14628 and n14210_not n14819 ; n14820
g14629 and asqrt[15] n14820 ; n14821
g14630 nor n14210 n14219 ; n14822
g14631 and asqrt[15] n14822 ; n14823
g14632 nor n14217 n14823 ; n14824
g14633 nor n14821 n14824 ; n14825
g14634 nor asqrt[29] n14806 ; n14826
g14635 and n14816_not n14826 ; n14827
g14636 nor n14825 n14827 ; n14828
g14637 nor n14818 n14828 ; n14829
g14638 and asqrt[30] n14829_not ; n14830
g14639 and n14222_not n14229 ; n14831
g14640 and n14231_not n14831 ; n14832
g14641 and asqrt[15] n14832 ; n14833
g14642 nor n14222 n14231 ; n14834
g14643 and asqrt[15] n14834 ; n14835
g14644 nor n14229 n14835 ; n14836
g14645 nor n14833 n14836 ; n14837
g14646 nor asqrt[30] n14818 ; n14838
g14647 and n14828_not n14838 ; n14839
g14648 nor n14837 n14839 ; n14840
g14649 nor n14830 n14840 ; n14841
g14650 and asqrt[31] n14841_not ; n14842
g14651 and n14241 n14243_not ; n14843
g14652 and n14234_not n14843 ; n14844
g14653 and asqrt[15] n14844 ; n14845
g14654 nor n14234 n14243 ; n14846
g14655 and asqrt[15] n14846 ; n14847
g14656 nor n14241 n14847 ; n14848
g14657 nor n14845 n14848 ; n14849
g14658 nor asqrt[31] n14830 ; n14850
g14659 and n14840_not n14850 ; n14851
g14660 nor n14849 n14851 ; n14852
g14661 nor n14842 n14852 ; n14853
g14662 and asqrt[32] n14853_not ; n14854
g14663 and n14246_not n14253 ; n14855
g14664 and n14255_not n14855 ; n14856
g14665 and asqrt[15] n14856 ; n14857
g14666 nor n14246 n14255 ; n14858
g14667 and asqrt[15] n14858 ; n14859
g14668 nor n14253 n14859 ; n14860
g14669 nor n14857 n14860 ; n14861
g14670 nor asqrt[32] n14842 ; n14862
g14671 and n14852_not n14862 ; n14863
g14672 nor n14861 n14863 ; n14864
g14673 nor n14854 n14864 ; n14865
g14674 and asqrt[33] n14865_not ; n14866
g14675 and n14265 n14267_not ; n14867
g14676 and n14258_not n14867 ; n14868
g14677 and asqrt[15] n14868 ; n14869
g14678 nor n14258 n14267 ; n14870
g14679 and asqrt[15] n14870 ; n14871
g14680 nor n14265 n14871 ; n14872
g14681 nor n14869 n14872 ; n14873
g14682 nor asqrt[33] n14854 ; n14874
g14683 and n14864_not n14874 ; n14875
g14684 nor n14873 n14875 ; n14876
g14685 nor n14866 n14876 ; n14877
g14686 and asqrt[34] n14877_not ; n14878
g14687 and n14270_not n14277 ; n14879
g14688 and n14279_not n14879 ; n14880
g14689 and asqrt[15] n14880 ; n14881
g14690 nor n14270 n14279 ; n14882
g14691 and asqrt[15] n14882 ; n14883
g14692 nor n14277 n14883 ; n14884
g14693 nor n14881 n14884 ; n14885
g14694 nor asqrt[34] n14866 ; n14886
g14695 and n14876_not n14886 ; n14887
g14696 nor n14885 n14887 ; n14888
g14697 nor n14878 n14888 ; n14889
g14698 and asqrt[35] n14889_not ; n14890
g14699 and n14289 n14291_not ; n14891
g14700 and n14282_not n14891 ; n14892
g14701 and asqrt[15] n14892 ; n14893
g14702 nor n14282 n14291 ; n14894
g14703 and asqrt[15] n14894 ; n14895
g14704 nor n14289 n14895 ; n14896
g14705 nor n14893 n14896 ; n14897
g14706 nor asqrt[35] n14878 ; n14898
g14707 and n14888_not n14898 ; n14899
g14708 nor n14897 n14899 ; n14900
g14709 nor n14890 n14900 ; n14901
g14710 and asqrt[36] n14901_not ; n14902
g14711 and n14294_not n14301 ; n14903
g14712 and n14303_not n14903 ; n14904
g14713 and asqrt[15] n14904 ; n14905
g14714 nor n14294 n14303 ; n14906
g14715 and asqrt[15] n14906 ; n14907
g14716 nor n14301 n14907 ; n14908
g14717 nor n14905 n14908 ; n14909
g14718 nor asqrt[36] n14890 ; n14910
g14719 and n14900_not n14910 ; n14911
g14720 nor n14909 n14911 ; n14912
g14721 nor n14902 n14912 ; n14913
g14722 and asqrt[37] n14913_not ; n14914
g14723 and n14313 n14315_not ; n14915
g14724 and n14306_not n14915 ; n14916
g14725 and asqrt[15] n14916 ; n14917
g14726 nor n14306 n14315 ; n14918
g14727 and asqrt[15] n14918 ; n14919
g14728 nor n14313 n14919 ; n14920
g14729 nor n14917 n14920 ; n14921
g14730 nor asqrt[37] n14902 ; n14922
g14731 and n14912_not n14922 ; n14923
g14732 nor n14921 n14923 ; n14924
g14733 nor n14914 n14924 ; n14925
g14734 and asqrt[38] n14925_not ; n14926
g14735 and n14318_not n14325 ; n14927
g14736 and n14327_not n14927 ; n14928
g14737 and asqrt[15] n14928 ; n14929
g14738 nor n14318 n14327 ; n14930
g14739 and asqrt[15] n14930 ; n14931
g14740 nor n14325 n14931 ; n14932
g14741 nor n14929 n14932 ; n14933
g14742 nor asqrt[38] n14914 ; n14934
g14743 and n14924_not n14934 ; n14935
g14744 nor n14933 n14935 ; n14936
g14745 nor n14926 n14936 ; n14937
g14746 and asqrt[39] n14937_not ; n14938
g14747 and n14337 n14339_not ; n14939
g14748 and n14330_not n14939 ; n14940
g14749 and asqrt[15] n14940 ; n14941
g14750 nor n14330 n14339 ; n14942
g14751 and asqrt[15] n14942 ; n14943
g14752 nor n14337 n14943 ; n14944
g14753 nor n14941 n14944 ; n14945
g14754 nor asqrt[39] n14926 ; n14946
g14755 and n14936_not n14946 ; n14947
g14756 nor n14945 n14947 ; n14948
g14757 nor n14938 n14948 ; n14949
g14758 and asqrt[40] n14949_not ; n14950
g14759 and n14342_not n14349 ; n14951
g14760 and n14351_not n14951 ; n14952
g14761 and asqrt[15] n14952 ; n14953
g14762 nor n14342 n14351 ; n14954
g14763 and asqrt[15] n14954 ; n14955
g14764 nor n14349 n14955 ; n14956
g14765 nor n14953 n14956 ; n14957
g14766 nor asqrt[40] n14938 ; n14958
g14767 and n14948_not n14958 ; n14959
g14768 nor n14957 n14959 ; n14960
g14769 nor n14950 n14960 ; n14961
g14770 and asqrt[41] n14961_not ; n14962
g14771 and n14361 n14363_not ; n14963
g14772 and n14354_not n14963 ; n14964
g14773 and asqrt[15] n14964 ; n14965
g14774 nor n14354 n14363 ; n14966
g14775 and asqrt[15] n14966 ; n14967
g14776 nor n14361 n14967 ; n14968
g14777 nor n14965 n14968 ; n14969
g14778 nor asqrt[41] n14950 ; n14970
g14779 and n14960_not n14970 ; n14971
g14780 nor n14969 n14971 ; n14972
g14781 nor n14962 n14972 ; n14973
g14782 and asqrt[42] n14973_not ; n14974
g14783 and n14366_not n14373 ; n14975
g14784 and n14375_not n14975 ; n14976
g14785 and asqrt[15] n14976 ; n14977
g14786 nor n14366 n14375 ; n14978
g14787 and asqrt[15] n14978 ; n14979
g14788 nor n14373 n14979 ; n14980
g14789 nor n14977 n14980 ; n14981
g14790 nor asqrt[42] n14962 ; n14982
g14791 and n14972_not n14982 ; n14983
g14792 nor n14981 n14983 ; n14984
g14793 nor n14974 n14984 ; n14985
g14794 and asqrt[43] n14985_not ; n14986
g14795 and n14385 n14387_not ; n14987
g14796 and n14378_not n14987 ; n14988
g14797 and asqrt[15] n14988 ; n14989
g14798 nor n14378 n14387 ; n14990
g14799 and asqrt[15] n14990 ; n14991
g14800 nor n14385 n14991 ; n14992
g14801 nor n14989 n14992 ; n14993
g14802 nor asqrt[43] n14974 ; n14994
g14803 and n14984_not n14994 ; n14995
g14804 nor n14993 n14995 ; n14996
g14805 nor n14986 n14996 ; n14997
g14806 and asqrt[44] n14997_not ; n14998
g14807 and n14390_not n14397 ; n14999
g14808 and n14399_not n14999 ; n15000
g14809 and asqrt[15] n15000 ; n15001
g14810 nor n14390 n14399 ; n15002
g14811 and asqrt[15] n15002 ; n15003
g14812 nor n14397 n15003 ; n15004
g14813 nor n15001 n15004 ; n15005
g14814 nor asqrt[44] n14986 ; n15006
g14815 and n14996_not n15006 ; n15007
g14816 nor n15005 n15007 ; n15008
g14817 nor n14998 n15008 ; n15009
g14818 and asqrt[45] n15009_not ; n15010
g14819 and n14409 n14411_not ; n15011
g14820 and n14402_not n15011 ; n15012
g14821 and asqrt[15] n15012 ; n15013
g14822 nor n14402 n14411 ; n15014
g14823 and asqrt[15] n15014 ; n15015
g14824 nor n14409 n15015 ; n15016
g14825 nor n15013 n15016 ; n15017
g14826 nor asqrt[45] n14998 ; n15018
g14827 and n15008_not n15018 ; n15019
g14828 nor n15017 n15019 ; n15020
g14829 nor n15010 n15020 ; n15021
g14830 and asqrt[46] n15021_not ; n15022
g14831 and n14414_not n14421 ; n15023
g14832 and n14423_not n15023 ; n15024
g14833 and asqrt[15] n15024 ; n15025
g14834 nor n14414 n14423 ; n15026
g14835 and asqrt[15] n15026 ; n15027
g14836 nor n14421 n15027 ; n15028
g14837 nor n15025 n15028 ; n15029
g14838 nor asqrt[46] n15010 ; n15030
g14839 and n15020_not n15030 ; n15031
g14840 nor n15029 n15031 ; n15032
g14841 nor n15022 n15032 ; n15033
g14842 and asqrt[47] n15033_not ; n15034
g14843 and n14433 n14435_not ; n15035
g14844 and n14426_not n15035 ; n15036
g14845 and asqrt[15] n15036 ; n15037
g14846 nor n14426 n14435 ; n15038
g14847 and asqrt[15] n15038 ; n15039
g14848 nor n14433 n15039 ; n15040
g14849 nor n15037 n15040 ; n15041
g14850 nor asqrt[47] n15022 ; n15042
g14851 and n15032_not n15042 ; n15043
g14852 nor n15041 n15043 ; n15044
g14853 nor n15034 n15044 ; n15045
g14854 and asqrt[48] n15045_not ; n15046
g14855 and n14438_not n14445 ; n15047
g14856 and n14447_not n15047 ; n15048
g14857 and asqrt[15] n15048 ; n15049
g14858 nor n14438 n14447 ; n15050
g14859 and asqrt[15] n15050 ; n15051
g14860 nor n14445 n15051 ; n15052
g14861 nor n15049 n15052 ; n15053
g14862 nor asqrt[48] n15034 ; n15054
g14863 and n15044_not n15054 ; n15055
g14864 nor n15053 n15055 ; n15056
g14865 nor n15046 n15056 ; n15057
g14866 and asqrt[49] n15057_not ; n15058
g14867 and n14457 n14459_not ; n15059
g14868 and n14450_not n15059 ; n15060
g14869 and asqrt[15] n15060 ; n15061
g14870 nor n14450 n14459 ; n15062
g14871 and asqrt[15] n15062 ; n15063
g14872 nor n14457 n15063 ; n15064
g14873 nor n15061 n15064 ; n15065
g14874 nor asqrt[49] n15046 ; n15066
g14875 and n15056_not n15066 ; n15067
g14876 nor n15065 n15067 ; n15068
g14877 nor n15058 n15068 ; n15069
g14878 and asqrt[50] n15069_not ; n15070
g14879 nor asqrt[50] n15058 ; n15071
g14880 and n15068_not n15071 ; n15072
g14881 and n14462_not n14471 ; n15073
g14882 and n14464_not n15073 ; n15074
g14883 and asqrt[15] n15074 ; n15075
g14884 nor n14462 n14464 ; n15076
g14885 and asqrt[15] n15076 ; n15077
g14886 nor n14471 n15077 ; n15078
g14887 nor n15075 n15078 ; n15079
g14888 nor n15072 n15079 ; n15080
g14889 nor n15070 n15080 ; n15081
g14890 and asqrt[51] n15081_not ; n15082
g14891 and n14481 n14483_not ; n15083
g14892 and n14474_not n15083 ; n15084
g14893 and asqrt[15] n15084 ; n15085
g14894 nor n14474 n14483 ; n15086
g14895 and asqrt[15] n15086 ; n15087
g14896 nor n14481 n15087 ; n15088
g14897 nor n15085 n15088 ; n15089
g14898 nor asqrt[51] n15070 ; n15090
g14899 and n15080_not n15090 ; n15091
g14900 nor n15089 n15091 ; n15092
g14901 nor n15082 n15092 ; n15093
g14902 and asqrt[52] n15093_not ; n15094
g14903 and n14486_not n14493 ; n15095
g14904 and n14495_not n15095 ; n15096
g14905 and asqrt[15] n15096 ; n15097
g14906 nor n14486 n14495 ; n15098
g14907 and asqrt[15] n15098 ; n15099
g14908 nor n14493 n15099 ; n15100
g14909 nor n15097 n15100 ; n15101
g14910 nor asqrt[52] n15082 ; n15102
g14911 and n15092_not n15102 ; n15103
g14912 nor n15101 n15103 ; n15104
g14913 nor n15094 n15104 ; n15105
g14914 and asqrt[53] n15105_not ; n15106
g14915 and n14505 n14507_not ; n15107
g14916 and n14498_not n15107 ; n15108
g14917 and asqrt[15] n15108 ; n15109
g14918 nor n14498 n14507 ; n15110
g14919 and asqrt[15] n15110 ; n15111
g14920 nor n14505 n15111 ; n15112
g14921 nor n15109 n15112 ; n15113
g14922 nor asqrt[53] n15094 ; n15114
g14923 and n15104_not n15114 ; n15115
g14924 nor n15113 n15115 ; n15116
g14925 nor n15106 n15116 ; n15117
g14926 and asqrt[54] n15117_not ; n15118
g14927 and n14510_not n14517 ; n15119
g14928 and n14519_not n15119 ; n15120
g14929 and asqrt[15] n15120 ; n15121
g14930 nor n14510 n14519 ; n15122
g14931 and asqrt[15] n15122 ; n15123
g14932 nor n14517 n15123 ; n15124
g14933 nor n15121 n15124 ; n15125
g14934 nor asqrt[54] n15106 ; n15126
g14935 and n15116_not n15126 ; n15127
g14936 nor n15125 n15127 ; n15128
g14937 nor n15118 n15128 ; n15129
g14938 and asqrt[55] n15129_not ; n15130
g14939 and n14529 n14531_not ; n15131
g14940 and n14522_not n15131 ; n15132
g14941 and asqrt[15] n15132 ; n15133
g14942 nor n14522 n14531 ; n15134
g14943 and asqrt[15] n15134 ; n15135
g14944 nor n14529 n15135 ; n15136
g14945 nor n15133 n15136 ; n15137
g14946 nor asqrt[55] n15118 ; n15138
g14947 and n15128_not n15138 ; n15139
g14948 nor n15137 n15139 ; n15140
g14949 nor n15130 n15140 ; n15141
g14950 and asqrt[56] n15141_not ; n15142
g14951 and n14534_not n14541 ; n15143
g14952 and n14543_not n15143 ; n15144
g14953 and asqrt[15] n15144 ; n15145
g14954 nor n14534 n14543 ; n15146
g14955 and asqrt[15] n15146 ; n15147
g14956 nor n14541 n15147 ; n15148
g14957 nor n15145 n15148 ; n15149
g14958 nor asqrt[56] n15130 ; n15150
g14959 and n15140_not n15150 ; n15151
g14960 nor n15149 n15151 ; n15152
g14961 nor n15142 n15152 ; n15153
g14962 and asqrt[57] n15153_not ; n15154
g14963 and n14553 n14555_not ; n15155
g14964 and n14546_not n15155 ; n15156
g14965 and asqrt[15] n15156 ; n15157
g14966 nor n14546 n14555 ; n15158
g14967 and asqrt[15] n15158 ; n15159
g14968 nor n14553 n15159 ; n15160
g14969 nor n15157 n15160 ; n15161
g14970 nor asqrt[57] n15142 ; n15162
g14971 and n15152_not n15162 ; n15163
g14972 nor n15161 n15163 ; n15164
g14973 nor n15154 n15164 ; n15165
g14974 and asqrt[58] n15165_not ; n15166
g14975 and n14558_not n14565 ; n15167
g14976 and n14567_not n15167 ; n15168
g14977 and asqrt[15] n15168 ; n15169
g14978 nor n14558 n14567 ; n15170
g14979 and asqrt[15] n15170 ; n15171
g14980 nor n14565 n15171 ; n15172
g14981 nor n15169 n15172 ; n15173
g14982 nor asqrt[58] n15154 ; n15174
g14983 and n15164_not n15174 ; n15175
g14984 nor n15173 n15175 ; n15176
g14985 nor n15166 n15176 ; n15177
g14986 and asqrt[59] n15177_not ; n15178
g14987 and n14577 n14579_not ; n15179
g14988 and n14570_not n15179 ; n15180
g14989 and asqrt[15] n15180 ; n15181
g14990 nor n14570 n14579 ; n15182
g14991 and asqrt[15] n15182 ; n15183
g14992 nor n14577 n15183 ; n15184
g14993 nor n15181 n15184 ; n15185
g14994 nor asqrt[59] n15166 ; n15186
g14995 and n15176_not n15186 ; n15187
g14996 nor n15185 n15187 ; n15188
g14997 nor n15178 n15188 ; n15189
g14998 and asqrt[60] n15189_not ; n15190
g14999 and n14582_not n14589 ; n15191
g15000 and n14591_not n15191 ; n15192
g15001 and asqrt[15] n15192 ; n15193
g15002 nor n14582 n14591 ; n15194
g15003 and asqrt[15] n15194 ; n15195
g15004 nor n14589 n15195 ; n15196
g15005 nor n15193 n15196 ; n15197
g15006 nor asqrt[60] n15178 ; n15198
g15007 and n15188_not n15198 ; n15199
g15008 nor n15197 n15199 ; n15200
g15009 nor n15190 n15200 ; n15201
g15010 and asqrt[61] n15201_not ; n15202
g15011 and n14601 n14603_not ; n15203
g15012 and n14594_not n15203 ; n15204
g15013 and asqrt[15] n15204 ; n15205
g15014 nor n14594 n14603 ; n15206
g15015 and asqrt[15] n15206 ; n15207
g15016 nor n14601 n15207 ; n15208
g15017 nor n15205 n15208 ; n15209
g15018 nor asqrt[61] n15190 ; n15210
g15019 and n15200_not n15210 ; n15211
g15020 nor n15209 n15211 ; n15212
g15021 nor n15202 n15212 ; n15213
g15022 and asqrt[62] n15213_not ; n15214
g15023 and n14606_not n14613 ; n15215
g15024 and n14615_not n15215 ; n15216
g15025 and asqrt[15] n15216 ; n15217
g15026 nor n14606 n14615 ; n15218
g15027 and asqrt[15] n15218 ; n15219
g15028 nor n14613 n15219 ; n15220
g15029 nor n15217 n15220 ; n15221
g15030 nor asqrt[62] n15202 ; n15222
g15031 and n15212_not n15222 ; n15223
g15032 nor n15221 n15223 ; n15224
g15033 nor n15214 n15224 ; n15225
g15034 and n14625 n14627_not ; n15226
g15035 and n14618_not n15226 ; n15227
g15036 and asqrt[15] n15227 ; n15228
g15037 nor n14618 n14627 ; n15229
g15038 and asqrt[15] n15229 ; n15230
g15039 nor n14625 n15230 ; n15231
g15040 nor n15228 n15231 ; n15232
g15041 nor n14629 n14636 ; n15233
g15042 and asqrt[15] n15233 ; n15234
g15043 nor n14644 n15234 ; n15235
g15044 and n15232_not n15235 ; n15236
g15045 and n15225_not n15236 ; n15237
g15046 nor asqrt[63] n15237 ; n15238
g15047 and n15214_not n15232 ; n15239
g15048 and n15224_not n15239 ; n15240
g15049 and n14636_not asqrt[15] ; n15241
g15050 and n14629 n15241_not ; n15242
g15051 and asqrt[63] n15233_not ; n15243
g15052 and n15242_not n15243 ; n15244
g15053 nor n14632 n14653 ; n15245
g15054 and n14635_not n15245 ; n15246
g15055 and n14648_not n15246 ; n15247
g15056 and n14644_not n15247 ; n15248
g15057 and n14642_not n15248 ; n15249
g15058 nor n15244 n15249 ; n15250
g15059 and n15240_not n15250 ; n15251
g15060 nand n15238_not n15251 ; asqrt[14]
g15061 and a[28] asqrt[14] ; n15253
g15062 nor a[26] a[27] ; n15254
g15063 and a[28]_not n15254 ; n15255
g15064 nor n15253 n15255 ; n15256
g15065 and asqrt[15] n15256_not ; n15257
g15066 nor n14653 n15255 ; n15258
g15067 and n14648_not n15258 ; n15259
g15068 and n14644_not n15259 ; n15260
g15069 and n14642_not n15260 ; n15261
g15070 and n15253_not n15261 ; n15262
g15071 and a[28]_not asqrt[14] ; n15263
g15072 and a[29] n15263_not ; n15264
g15073 and n14658 asqrt[14] ; n15265
g15074 nor n15264 n15265 ; n15266
g15075 and n15262_not n15266 ; n15267
g15076 nor n15257 n15267 ; n15268
g15077 and asqrt[16] n15268_not ; n15269
g15078 nor asqrt[16] n15257 ; n15270
g15079 and n15267_not n15270 ; n15271
g15080 and asqrt[15] n15249_not ; n15272
g15081 and n15244_not n15272 ; n15273
g15082 and n15240_not n15273 ; n15274
g15083 and n15238_not n15274 ; n15275
g15084 nor n15265 n15275 ; n15276
g15085 and a[30] n15276_not ; n15277
g15086 nor a[30] n15275 ; n15278
g15087 and n15265_not n15278 ; n15279
g15088 nor n15277 n15279 ; n15280
g15089 nor n15271 n15280 ; n15281
g15090 nor n15269 n15281 ; n15282
g15091 and asqrt[17] n15282_not ; n15283
g15092 nor n14661 n14666 ; n15284
g15093 and n14670_not n15284 ; n15285
g15094 and asqrt[14] n15285 ; n15286
g15095 and asqrt[14] n15284 ; n15287
g15096 and n14670 n15287_not ; n15288
g15097 nor n15286 n15288 ; n15289
g15098 nor asqrt[17] n15269 ; n15290
g15099 and n15281_not n15290 ; n15291
g15100 nor n15289 n15291 ; n15292
g15101 nor n15283 n15292 ; n15293
g15102 and asqrt[18] n15293_not ; n15294
g15103 and n14675_not n14684 ; n15295
g15104 and n14673_not n15295 ; n15296
g15105 and asqrt[14] n15296 ; n15297
g15106 nor n14673 n14675 ; n15298
g15107 and asqrt[14] n15298 ; n15299
g15108 nor n14684 n15299 ; n15300
g15109 nor n15297 n15300 ; n15301
g15110 nor asqrt[18] n15283 ; n15302
g15111 and n15292_not n15302 ; n15303
g15112 nor n15301 n15303 ; n15304
g15113 nor n15294 n15304 ; n15305
g15114 and asqrt[19] n15305_not ; n15306
g15115 and n14687_not n14693 ; n15307
g15116 and n14695_not n15307 ; n15308
g15117 and asqrt[14] n15308 ; n15309
g15118 nor n14687 n14695 ; n15310
g15119 and asqrt[14] n15310 ; n15311
g15120 nor n14693 n15311 ; n15312
g15121 nor n15309 n15312 ; n15313
g15122 nor asqrt[19] n15294 ; n15314
g15123 and n15304_not n15314 ; n15315
g15124 nor n15313 n15315 ; n15316
g15125 nor n15306 n15316 ; n15317
g15126 and asqrt[20] n15317_not ; n15318
g15127 and n14705 n14707_not ; n15319
g15128 and n14698_not n15319 ; n15320
g15129 and asqrt[14] n15320 ; n15321
g15130 nor n14698 n14707 ; n15322
g15131 and asqrt[14] n15322 ; n15323
g15132 nor n14705 n15323 ; n15324
g15133 nor n15321 n15324 ; n15325
g15134 nor asqrt[20] n15306 ; n15326
g15135 and n15316_not n15326 ; n15327
g15136 nor n15325 n15327 ; n15328
g15137 nor n15318 n15328 ; n15329
g15138 and asqrt[21] n15329_not ; n15330
g15139 and n14710_not n14717 ; n15331
g15140 and n14719_not n15331 ; n15332
g15141 and asqrt[14] n15332 ; n15333
g15142 nor n14710 n14719 ; n15334
g15143 and asqrt[14] n15334 ; n15335
g15144 nor n14717 n15335 ; n15336
g15145 nor n15333 n15336 ; n15337
g15146 nor asqrt[21] n15318 ; n15338
g15147 and n15328_not n15338 ; n15339
g15148 nor n15337 n15339 ; n15340
g15149 nor n15330 n15340 ; n15341
g15150 and asqrt[22] n15341_not ; n15342
g15151 and n14729 n14731_not ; n15343
g15152 and n14722_not n15343 ; n15344
g15153 and asqrt[14] n15344 ; n15345
g15154 nor n14722 n14731 ; n15346
g15155 and asqrt[14] n15346 ; n15347
g15156 nor n14729 n15347 ; n15348
g15157 nor n15345 n15348 ; n15349
g15158 nor asqrt[22] n15330 ; n15350
g15159 and n15340_not n15350 ; n15351
g15160 nor n15349 n15351 ; n15352
g15161 nor n15342 n15352 ; n15353
g15162 and asqrt[23] n15353_not ; n15354
g15163 and n14734_not n14741 ; n15355
g15164 and n14743_not n15355 ; n15356
g15165 and asqrt[14] n15356 ; n15357
g15166 nor n14734 n14743 ; n15358
g15167 and asqrt[14] n15358 ; n15359
g15168 nor n14741 n15359 ; n15360
g15169 nor n15357 n15360 ; n15361
g15170 nor asqrt[23] n15342 ; n15362
g15171 and n15352_not n15362 ; n15363
g15172 nor n15361 n15363 ; n15364
g15173 nor n15354 n15364 ; n15365
g15174 and asqrt[24] n15365_not ; n15366
g15175 and n14753 n14755_not ; n15367
g15176 and n14746_not n15367 ; n15368
g15177 and asqrt[14] n15368 ; n15369
g15178 nor n14746 n14755 ; n15370
g15179 and asqrt[14] n15370 ; n15371
g15180 nor n14753 n15371 ; n15372
g15181 nor n15369 n15372 ; n15373
g15182 nor asqrt[24] n15354 ; n15374
g15183 and n15364_not n15374 ; n15375
g15184 nor n15373 n15375 ; n15376
g15185 nor n15366 n15376 ; n15377
g15186 and asqrt[25] n15377_not ; n15378
g15187 and n14758_not n14765 ; n15379
g15188 and n14767_not n15379 ; n15380
g15189 and asqrt[14] n15380 ; n15381
g15190 nor n14758 n14767 ; n15382
g15191 and asqrt[14] n15382 ; n15383
g15192 nor n14765 n15383 ; n15384
g15193 nor n15381 n15384 ; n15385
g15194 nor asqrt[25] n15366 ; n15386
g15195 and n15376_not n15386 ; n15387
g15196 nor n15385 n15387 ; n15388
g15197 nor n15378 n15388 ; n15389
g15198 and asqrt[26] n15389_not ; n15390
g15199 and n14777 n14779_not ; n15391
g15200 and n14770_not n15391 ; n15392
g15201 and asqrt[14] n15392 ; n15393
g15202 nor n14770 n14779 ; n15394
g15203 and asqrt[14] n15394 ; n15395
g15204 nor n14777 n15395 ; n15396
g15205 nor n15393 n15396 ; n15397
g15206 nor asqrt[26] n15378 ; n15398
g15207 and n15388_not n15398 ; n15399
g15208 nor n15397 n15399 ; n15400
g15209 nor n15390 n15400 ; n15401
g15210 and asqrt[27] n15401_not ; n15402
g15211 and n14782_not n14789 ; n15403
g15212 and n14791_not n15403 ; n15404
g15213 and asqrt[14] n15404 ; n15405
g15214 nor n14782 n14791 ; n15406
g15215 and asqrt[14] n15406 ; n15407
g15216 nor n14789 n15407 ; n15408
g15217 nor n15405 n15408 ; n15409
g15218 nor asqrt[27] n15390 ; n15410
g15219 and n15400_not n15410 ; n15411
g15220 nor n15409 n15411 ; n15412
g15221 nor n15402 n15412 ; n15413
g15222 and asqrt[28] n15413_not ; n15414
g15223 and n14801 n14803_not ; n15415
g15224 and n14794_not n15415 ; n15416
g15225 and asqrt[14] n15416 ; n15417
g15226 nor n14794 n14803 ; n15418
g15227 and asqrt[14] n15418 ; n15419
g15228 nor n14801 n15419 ; n15420
g15229 nor n15417 n15420 ; n15421
g15230 nor asqrt[28] n15402 ; n15422
g15231 and n15412_not n15422 ; n15423
g15232 nor n15421 n15423 ; n15424
g15233 nor n15414 n15424 ; n15425
g15234 and asqrt[29] n15425_not ; n15426
g15235 and n14806_not n14813 ; n15427
g15236 and n14815_not n15427 ; n15428
g15237 and asqrt[14] n15428 ; n15429
g15238 nor n14806 n14815 ; n15430
g15239 and asqrt[14] n15430 ; n15431
g15240 nor n14813 n15431 ; n15432
g15241 nor n15429 n15432 ; n15433
g15242 nor asqrt[29] n15414 ; n15434
g15243 and n15424_not n15434 ; n15435
g15244 nor n15433 n15435 ; n15436
g15245 nor n15426 n15436 ; n15437
g15246 and asqrt[30] n15437_not ; n15438
g15247 and n14825 n14827_not ; n15439
g15248 and n14818_not n15439 ; n15440
g15249 and asqrt[14] n15440 ; n15441
g15250 nor n14818 n14827 ; n15442
g15251 and asqrt[14] n15442 ; n15443
g15252 nor n14825 n15443 ; n15444
g15253 nor n15441 n15444 ; n15445
g15254 nor asqrt[30] n15426 ; n15446
g15255 and n15436_not n15446 ; n15447
g15256 nor n15445 n15447 ; n15448
g15257 nor n15438 n15448 ; n15449
g15258 and asqrt[31] n15449_not ; n15450
g15259 and n14830_not n14837 ; n15451
g15260 and n14839_not n15451 ; n15452
g15261 and asqrt[14] n15452 ; n15453
g15262 nor n14830 n14839 ; n15454
g15263 and asqrt[14] n15454 ; n15455
g15264 nor n14837 n15455 ; n15456
g15265 nor n15453 n15456 ; n15457
g15266 nor asqrt[31] n15438 ; n15458
g15267 and n15448_not n15458 ; n15459
g15268 nor n15457 n15459 ; n15460
g15269 nor n15450 n15460 ; n15461
g15270 and asqrt[32] n15461_not ; n15462
g15271 and n14849 n14851_not ; n15463
g15272 and n14842_not n15463 ; n15464
g15273 and asqrt[14] n15464 ; n15465
g15274 nor n14842 n14851 ; n15466
g15275 and asqrt[14] n15466 ; n15467
g15276 nor n14849 n15467 ; n15468
g15277 nor n15465 n15468 ; n15469
g15278 nor asqrt[32] n15450 ; n15470
g15279 and n15460_not n15470 ; n15471
g15280 nor n15469 n15471 ; n15472
g15281 nor n15462 n15472 ; n15473
g15282 and asqrt[33] n15473_not ; n15474
g15283 and n14854_not n14861 ; n15475
g15284 and n14863_not n15475 ; n15476
g15285 and asqrt[14] n15476 ; n15477
g15286 nor n14854 n14863 ; n15478
g15287 and asqrt[14] n15478 ; n15479
g15288 nor n14861 n15479 ; n15480
g15289 nor n15477 n15480 ; n15481
g15290 nor asqrt[33] n15462 ; n15482
g15291 and n15472_not n15482 ; n15483
g15292 nor n15481 n15483 ; n15484
g15293 nor n15474 n15484 ; n15485
g15294 and asqrt[34] n15485_not ; n15486
g15295 and n14873 n14875_not ; n15487
g15296 and n14866_not n15487 ; n15488
g15297 and asqrt[14] n15488 ; n15489
g15298 nor n14866 n14875 ; n15490
g15299 and asqrt[14] n15490 ; n15491
g15300 nor n14873 n15491 ; n15492
g15301 nor n15489 n15492 ; n15493
g15302 nor asqrt[34] n15474 ; n15494
g15303 and n15484_not n15494 ; n15495
g15304 nor n15493 n15495 ; n15496
g15305 nor n15486 n15496 ; n15497
g15306 and asqrt[35] n15497_not ; n15498
g15307 and n14878_not n14885 ; n15499
g15308 and n14887_not n15499 ; n15500
g15309 and asqrt[14] n15500 ; n15501
g15310 nor n14878 n14887 ; n15502
g15311 and asqrt[14] n15502 ; n15503
g15312 nor n14885 n15503 ; n15504
g15313 nor n15501 n15504 ; n15505
g15314 nor asqrt[35] n15486 ; n15506
g15315 and n15496_not n15506 ; n15507
g15316 nor n15505 n15507 ; n15508
g15317 nor n15498 n15508 ; n15509
g15318 and asqrt[36] n15509_not ; n15510
g15319 and n14897 n14899_not ; n15511
g15320 and n14890_not n15511 ; n15512
g15321 and asqrt[14] n15512 ; n15513
g15322 nor n14890 n14899 ; n15514
g15323 and asqrt[14] n15514 ; n15515
g15324 nor n14897 n15515 ; n15516
g15325 nor n15513 n15516 ; n15517
g15326 nor asqrt[36] n15498 ; n15518
g15327 and n15508_not n15518 ; n15519
g15328 nor n15517 n15519 ; n15520
g15329 nor n15510 n15520 ; n15521
g15330 and asqrt[37] n15521_not ; n15522
g15331 and n14902_not n14909 ; n15523
g15332 and n14911_not n15523 ; n15524
g15333 and asqrt[14] n15524 ; n15525
g15334 nor n14902 n14911 ; n15526
g15335 and asqrt[14] n15526 ; n15527
g15336 nor n14909 n15527 ; n15528
g15337 nor n15525 n15528 ; n15529
g15338 nor asqrt[37] n15510 ; n15530
g15339 and n15520_not n15530 ; n15531
g15340 nor n15529 n15531 ; n15532
g15341 nor n15522 n15532 ; n15533
g15342 and asqrt[38] n15533_not ; n15534
g15343 and n14921 n14923_not ; n15535
g15344 and n14914_not n15535 ; n15536
g15345 and asqrt[14] n15536 ; n15537
g15346 nor n14914 n14923 ; n15538
g15347 and asqrt[14] n15538 ; n15539
g15348 nor n14921 n15539 ; n15540
g15349 nor n15537 n15540 ; n15541
g15350 nor asqrt[38] n15522 ; n15542
g15351 and n15532_not n15542 ; n15543
g15352 nor n15541 n15543 ; n15544
g15353 nor n15534 n15544 ; n15545
g15354 and asqrt[39] n15545_not ; n15546
g15355 and n14926_not n14933 ; n15547
g15356 and n14935_not n15547 ; n15548
g15357 and asqrt[14] n15548 ; n15549
g15358 nor n14926 n14935 ; n15550
g15359 and asqrt[14] n15550 ; n15551
g15360 nor n14933 n15551 ; n15552
g15361 nor n15549 n15552 ; n15553
g15362 nor asqrt[39] n15534 ; n15554
g15363 and n15544_not n15554 ; n15555
g15364 nor n15553 n15555 ; n15556
g15365 nor n15546 n15556 ; n15557
g15366 and asqrt[40] n15557_not ; n15558
g15367 and n14945 n14947_not ; n15559
g15368 and n14938_not n15559 ; n15560
g15369 and asqrt[14] n15560 ; n15561
g15370 nor n14938 n14947 ; n15562
g15371 and asqrt[14] n15562 ; n15563
g15372 nor n14945 n15563 ; n15564
g15373 nor n15561 n15564 ; n15565
g15374 nor asqrt[40] n15546 ; n15566
g15375 and n15556_not n15566 ; n15567
g15376 nor n15565 n15567 ; n15568
g15377 nor n15558 n15568 ; n15569
g15378 and asqrt[41] n15569_not ; n15570
g15379 and n14950_not n14957 ; n15571
g15380 and n14959_not n15571 ; n15572
g15381 and asqrt[14] n15572 ; n15573
g15382 nor n14950 n14959 ; n15574
g15383 and asqrt[14] n15574 ; n15575
g15384 nor n14957 n15575 ; n15576
g15385 nor n15573 n15576 ; n15577
g15386 nor asqrt[41] n15558 ; n15578
g15387 and n15568_not n15578 ; n15579
g15388 nor n15577 n15579 ; n15580
g15389 nor n15570 n15580 ; n15581
g15390 and asqrt[42] n15581_not ; n15582
g15391 and n14969 n14971_not ; n15583
g15392 and n14962_not n15583 ; n15584
g15393 and asqrt[14] n15584 ; n15585
g15394 nor n14962 n14971 ; n15586
g15395 and asqrt[14] n15586 ; n15587
g15396 nor n14969 n15587 ; n15588
g15397 nor n15585 n15588 ; n15589
g15398 nor asqrt[42] n15570 ; n15590
g15399 and n15580_not n15590 ; n15591
g15400 nor n15589 n15591 ; n15592
g15401 nor n15582 n15592 ; n15593
g15402 and asqrt[43] n15593_not ; n15594
g15403 and n14974_not n14981 ; n15595
g15404 and n14983_not n15595 ; n15596
g15405 and asqrt[14] n15596 ; n15597
g15406 nor n14974 n14983 ; n15598
g15407 and asqrt[14] n15598 ; n15599
g15408 nor n14981 n15599 ; n15600
g15409 nor n15597 n15600 ; n15601
g15410 nor asqrt[43] n15582 ; n15602
g15411 and n15592_not n15602 ; n15603
g15412 nor n15601 n15603 ; n15604
g15413 nor n15594 n15604 ; n15605
g15414 and asqrt[44] n15605_not ; n15606
g15415 and n14993 n14995_not ; n15607
g15416 and n14986_not n15607 ; n15608
g15417 and asqrt[14] n15608 ; n15609
g15418 nor n14986 n14995 ; n15610
g15419 and asqrt[14] n15610 ; n15611
g15420 nor n14993 n15611 ; n15612
g15421 nor n15609 n15612 ; n15613
g15422 nor asqrt[44] n15594 ; n15614
g15423 and n15604_not n15614 ; n15615
g15424 nor n15613 n15615 ; n15616
g15425 nor n15606 n15616 ; n15617
g15426 and asqrt[45] n15617_not ; n15618
g15427 and n14998_not n15005 ; n15619
g15428 and n15007_not n15619 ; n15620
g15429 and asqrt[14] n15620 ; n15621
g15430 nor n14998 n15007 ; n15622
g15431 and asqrt[14] n15622 ; n15623
g15432 nor n15005 n15623 ; n15624
g15433 nor n15621 n15624 ; n15625
g15434 nor asqrt[45] n15606 ; n15626
g15435 and n15616_not n15626 ; n15627
g15436 nor n15625 n15627 ; n15628
g15437 nor n15618 n15628 ; n15629
g15438 and asqrt[46] n15629_not ; n15630
g15439 and n15017 n15019_not ; n15631
g15440 and n15010_not n15631 ; n15632
g15441 and asqrt[14] n15632 ; n15633
g15442 nor n15010 n15019 ; n15634
g15443 and asqrt[14] n15634 ; n15635
g15444 nor n15017 n15635 ; n15636
g15445 nor n15633 n15636 ; n15637
g15446 nor asqrt[46] n15618 ; n15638
g15447 and n15628_not n15638 ; n15639
g15448 nor n15637 n15639 ; n15640
g15449 nor n15630 n15640 ; n15641
g15450 and asqrt[47] n15641_not ; n15642
g15451 and n15022_not n15029 ; n15643
g15452 and n15031_not n15643 ; n15644
g15453 and asqrt[14] n15644 ; n15645
g15454 nor n15022 n15031 ; n15646
g15455 and asqrt[14] n15646 ; n15647
g15456 nor n15029 n15647 ; n15648
g15457 nor n15645 n15648 ; n15649
g15458 nor asqrt[47] n15630 ; n15650
g15459 and n15640_not n15650 ; n15651
g15460 nor n15649 n15651 ; n15652
g15461 nor n15642 n15652 ; n15653
g15462 and asqrt[48] n15653_not ; n15654
g15463 and n15041 n15043_not ; n15655
g15464 and n15034_not n15655 ; n15656
g15465 and asqrt[14] n15656 ; n15657
g15466 nor n15034 n15043 ; n15658
g15467 and asqrt[14] n15658 ; n15659
g15468 nor n15041 n15659 ; n15660
g15469 nor n15657 n15660 ; n15661
g15470 nor asqrt[48] n15642 ; n15662
g15471 and n15652_not n15662 ; n15663
g15472 nor n15661 n15663 ; n15664
g15473 nor n15654 n15664 ; n15665
g15474 and asqrt[49] n15665_not ; n15666
g15475 and n15046_not n15053 ; n15667
g15476 and n15055_not n15667 ; n15668
g15477 and asqrt[14] n15668 ; n15669
g15478 nor n15046 n15055 ; n15670
g15479 and asqrt[14] n15670 ; n15671
g15480 nor n15053 n15671 ; n15672
g15481 nor n15669 n15672 ; n15673
g15482 nor asqrt[49] n15654 ; n15674
g15483 and n15664_not n15674 ; n15675
g15484 nor n15673 n15675 ; n15676
g15485 nor n15666 n15676 ; n15677
g15486 and asqrt[50] n15677_not ; n15678
g15487 and n15065 n15067_not ; n15679
g15488 and n15058_not n15679 ; n15680
g15489 and asqrt[14] n15680 ; n15681
g15490 nor n15058 n15067 ; n15682
g15491 and asqrt[14] n15682 ; n15683
g15492 nor n15065 n15683 ; n15684
g15493 nor n15681 n15684 ; n15685
g15494 nor asqrt[50] n15666 ; n15686
g15495 and n15676_not n15686 ; n15687
g15496 nor n15685 n15687 ; n15688
g15497 nor n15678 n15688 ; n15689
g15498 and asqrt[51] n15689_not ; n15690
g15499 nor asqrt[51] n15678 ; n15691
g15500 and n15688_not n15691 ; n15692
g15501 and n15070_not n15079 ; n15693
g15502 and n15072_not n15693 ; n15694
g15503 and asqrt[14] n15694 ; n15695
g15504 nor n15070 n15072 ; n15696
g15505 and asqrt[14] n15696 ; n15697
g15506 nor n15079 n15697 ; n15698
g15507 nor n15695 n15698 ; n15699
g15508 nor n15692 n15699 ; n15700
g15509 nor n15690 n15700 ; n15701
g15510 and asqrt[52] n15701_not ; n15702
g15511 and n15089 n15091_not ; n15703
g15512 and n15082_not n15703 ; n15704
g15513 and asqrt[14] n15704 ; n15705
g15514 nor n15082 n15091 ; n15706
g15515 and asqrt[14] n15706 ; n15707
g15516 nor n15089 n15707 ; n15708
g15517 nor n15705 n15708 ; n15709
g15518 nor asqrt[52] n15690 ; n15710
g15519 and n15700_not n15710 ; n15711
g15520 nor n15709 n15711 ; n15712
g15521 nor n15702 n15712 ; n15713
g15522 and asqrt[53] n15713_not ; n15714
g15523 and n15094_not n15101 ; n15715
g15524 and n15103_not n15715 ; n15716
g15525 and asqrt[14] n15716 ; n15717
g15526 nor n15094 n15103 ; n15718
g15527 and asqrt[14] n15718 ; n15719
g15528 nor n15101 n15719 ; n15720
g15529 nor n15717 n15720 ; n15721
g15530 nor asqrt[53] n15702 ; n15722
g15531 and n15712_not n15722 ; n15723
g15532 nor n15721 n15723 ; n15724
g15533 nor n15714 n15724 ; n15725
g15534 and asqrt[54] n15725_not ; n15726
g15535 and n15113 n15115_not ; n15727
g15536 and n15106_not n15727 ; n15728
g15537 and asqrt[14] n15728 ; n15729
g15538 nor n15106 n15115 ; n15730
g15539 and asqrt[14] n15730 ; n15731
g15540 nor n15113 n15731 ; n15732
g15541 nor n15729 n15732 ; n15733
g15542 nor asqrt[54] n15714 ; n15734
g15543 and n15724_not n15734 ; n15735
g15544 nor n15733 n15735 ; n15736
g15545 nor n15726 n15736 ; n15737
g15546 and asqrt[55] n15737_not ; n15738
g15547 and n15118_not n15125 ; n15739
g15548 and n15127_not n15739 ; n15740
g15549 and asqrt[14] n15740 ; n15741
g15550 nor n15118 n15127 ; n15742
g15551 and asqrt[14] n15742 ; n15743
g15552 nor n15125 n15743 ; n15744
g15553 nor n15741 n15744 ; n15745
g15554 nor asqrt[55] n15726 ; n15746
g15555 and n15736_not n15746 ; n15747
g15556 nor n15745 n15747 ; n15748
g15557 nor n15738 n15748 ; n15749
g15558 and asqrt[56] n15749_not ; n15750
g15559 and n15137 n15139_not ; n15751
g15560 and n15130_not n15751 ; n15752
g15561 and asqrt[14] n15752 ; n15753
g15562 nor n15130 n15139 ; n15754
g15563 and asqrt[14] n15754 ; n15755
g15564 nor n15137 n15755 ; n15756
g15565 nor n15753 n15756 ; n15757
g15566 nor asqrt[56] n15738 ; n15758
g15567 and n15748_not n15758 ; n15759
g15568 nor n15757 n15759 ; n15760
g15569 nor n15750 n15760 ; n15761
g15570 and asqrt[57] n15761_not ; n15762
g15571 and n15142_not n15149 ; n15763
g15572 and n15151_not n15763 ; n15764
g15573 and asqrt[14] n15764 ; n15765
g15574 nor n15142 n15151 ; n15766
g15575 and asqrt[14] n15766 ; n15767
g15576 nor n15149 n15767 ; n15768
g15577 nor n15765 n15768 ; n15769
g15578 nor asqrt[57] n15750 ; n15770
g15579 and n15760_not n15770 ; n15771
g15580 nor n15769 n15771 ; n15772
g15581 nor n15762 n15772 ; n15773
g15582 and asqrt[58] n15773_not ; n15774
g15583 and n15161 n15163_not ; n15775
g15584 and n15154_not n15775 ; n15776
g15585 and asqrt[14] n15776 ; n15777
g15586 nor n15154 n15163 ; n15778
g15587 and asqrt[14] n15778 ; n15779
g15588 nor n15161 n15779 ; n15780
g15589 nor n15777 n15780 ; n15781
g15590 nor asqrt[58] n15762 ; n15782
g15591 and n15772_not n15782 ; n15783
g15592 nor n15781 n15783 ; n15784
g15593 nor n15774 n15784 ; n15785
g15594 and asqrt[59] n15785_not ; n15786
g15595 and n15166_not n15173 ; n15787
g15596 and n15175_not n15787 ; n15788
g15597 and asqrt[14] n15788 ; n15789
g15598 nor n15166 n15175 ; n15790
g15599 and asqrt[14] n15790 ; n15791
g15600 nor n15173 n15791 ; n15792
g15601 nor n15789 n15792 ; n15793
g15602 nor asqrt[59] n15774 ; n15794
g15603 and n15784_not n15794 ; n15795
g15604 nor n15793 n15795 ; n15796
g15605 nor n15786 n15796 ; n15797
g15606 and asqrt[60] n15797_not ; n15798
g15607 and n15185 n15187_not ; n15799
g15608 and n15178_not n15799 ; n15800
g15609 and asqrt[14] n15800 ; n15801
g15610 nor n15178 n15187 ; n15802
g15611 and asqrt[14] n15802 ; n15803
g15612 nor n15185 n15803 ; n15804
g15613 nor n15801 n15804 ; n15805
g15614 nor asqrt[60] n15786 ; n15806
g15615 and n15796_not n15806 ; n15807
g15616 nor n15805 n15807 ; n15808
g15617 nor n15798 n15808 ; n15809
g15618 and asqrt[61] n15809_not ; n15810
g15619 and n15190_not n15197 ; n15811
g15620 and n15199_not n15811 ; n15812
g15621 and asqrt[14] n15812 ; n15813
g15622 nor n15190 n15199 ; n15814
g15623 and asqrt[14] n15814 ; n15815
g15624 nor n15197 n15815 ; n15816
g15625 nor n15813 n15816 ; n15817
g15626 nor asqrt[61] n15798 ; n15818
g15627 and n15808_not n15818 ; n15819
g15628 nor n15817 n15819 ; n15820
g15629 nor n15810 n15820 ; n15821
g15630 and asqrt[62] n15821_not ; n15822
g15631 and n15209 n15211_not ; n15823
g15632 and n15202_not n15823 ; n15824
g15633 and asqrt[14] n15824 ; n15825
g15634 nor n15202 n15211 ; n15826
g15635 and asqrt[14] n15826 ; n15827
g15636 nor n15209 n15827 ; n15828
g15637 nor n15825 n15828 ; n15829
g15638 nor asqrt[62] n15810 ; n15830
g15639 and n15820_not n15830 ; n15831
g15640 nor n15829 n15831 ; n15832
g15641 nor n15822 n15832 ; n15833
g15642 and n15214_not n15221 ; n15834
g15643 and n15223_not n15834 ; n15835
g15644 and asqrt[14] n15835 ; n15836
g15645 nor n15214 n15223 ; n15837
g15646 and asqrt[14] n15837 ; n15838
g15647 nor n15221 n15838 ; n15839
g15648 nor n15836 n15839 ; n15840
g15649 nor n15225 n15232 ; n15841
g15650 and asqrt[14] n15841 ; n15842
g15651 nor n15240 n15842 ; n15843
g15652 and n15840_not n15843 ; n15844
g15653 and n15833_not n15844 ; n15845
g15654 nor asqrt[63] n15845 ; n15846
g15655 and n15822_not n15840 ; n15847
g15656 and n15832_not n15847 ; n15848
g15657 and n15232_not asqrt[14] ; n15849
g15658 and n15225 n15849_not ; n15850
g15659 and asqrt[63] n15841_not ; n15851
g15660 and n15850_not n15851 ; n15852
g15661 nor n15228 n15249 ; n15853
g15662 and n15231_not n15853 ; n15854
g15663 and n15244_not n15854 ; n15855
g15664 and n15240_not n15855 ; n15856
g15665 and n15238_not n15856 ; n15857
g15666 nor n15852 n15857 ; n15858
g15667 and n15848_not n15858 ; n15859
g15668 nand n15846_not n15859 ; asqrt[13]
g15669 and a[26] asqrt[13] ; n15861
g15670 nor a[24] a[25] ; n15862
g15671 and a[26]_not n15862 ; n15863
g15672 nor n15861 n15863 ; n15864
g15673 and asqrt[14] n15864_not ; n15865
g15674 nor n15249 n15863 ; n15866
g15675 and n15244_not n15866 ; n15867
g15676 and n15240_not n15867 ; n15868
g15677 and n15238_not n15868 ; n15869
g15678 and n15861_not n15869 ; n15870
g15679 and a[26]_not asqrt[13] ; n15871
g15680 and a[27] n15871_not ; n15872
g15681 and n15254 asqrt[13] ; n15873
g15682 nor n15872 n15873 ; n15874
g15683 and n15870_not n15874 ; n15875
g15684 nor n15865 n15875 ; n15876
g15685 and asqrt[15] n15876_not ; n15877
g15686 nor asqrt[15] n15865 ; n15878
g15687 and n15875_not n15878 ; n15879
g15688 and asqrt[14] n15857_not ; n15880
g15689 and n15852_not n15880 ; n15881
g15690 and n15848_not n15881 ; n15882
g15691 and n15846_not n15882 ; n15883
g15692 nor n15873 n15883 ; n15884
g15693 and a[28] n15884_not ; n15885
g15694 nor a[28] n15883 ; n15886
g15695 and n15873_not n15886 ; n15887
g15696 nor n15885 n15887 ; n15888
g15697 nor n15879 n15888 ; n15889
g15698 nor n15877 n15889 ; n15890
g15699 and asqrt[16] n15890_not ; n15891
g15700 nor n15257 n15262 ; n15892
g15701 and n15266_not n15892 ; n15893
g15702 and asqrt[13] n15893 ; n15894
g15703 and asqrt[13] n15892 ; n15895
g15704 and n15266 n15895_not ; n15896
g15705 nor n15894 n15896 ; n15897
g15706 nor asqrt[16] n15877 ; n15898
g15707 and n15889_not n15898 ; n15899
g15708 nor n15897 n15899 ; n15900
g15709 nor n15891 n15900 ; n15901
g15710 and asqrt[17] n15901_not ; n15902
g15711 and n15271_not n15280 ; n15903
g15712 and n15269_not n15903 ; n15904
g15713 and asqrt[13] n15904 ; n15905
g15714 nor n15269 n15271 ; n15906
g15715 and asqrt[13] n15906 ; n15907
g15716 nor n15280 n15907 ; n15908
g15717 nor n15905 n15908 ; n15909
g15718 nor asqrt[17] n15891 ; n15910
g15719 and n15900_not n15910 ; n15911
g15720 nor n15909 n15911 ; n15912
g15721 nor n15902 n15912 ; n15913
g15722 and asqrt[18] n15913_not ; n15914
g15723 and n15283_not n15289 ; n15915
g15724 and n15291_not n15915 ; n15916
g15725 and asqrt[13] n15916 ; n15917
g15726 nor n15283 n15291 ; n15918
g15727 and asqrt[13] n15918 ; n15919
g15728 nor n15289 n15919 ; n15920
g15729 nor n15917 n15920 ; n15921
g15730 nor asqrt[18] n15902 ; n15922
g15731 and n15912_not n15922 ; n15923
g15732 nor n15921 n15923 ; n15924
g15733 nor n15914 n15924 ; n15925
g15734 and asqrt[19] n15925_not ; n15926
g15735 and n15301 n15303_not ; n15927
g15736 and n15294_not n15927 ; n15928
g15737 and asqrt[13] n15928 ; n15929
g15738 nor n15294 n15303 ; n15930
g15739 and asqrt[13] n15930 ; n15931
g15740 nor n15301 n15931 ; n15932
g15741 nor n15929 n15932 ; n15933
g15742 nor asqrt[19] n15914 ; n15934
g15743 and n15924_not n15934 ; n15935
g15744 nor n15933 n15935 ; n15936
g15745 nor n15926 n15936 ; n15937
g15746 and asqrt[20] n15937_not ; n15938
g15747 and n15306_not n15313 ; n15939
g15748 and n15315_not n15939 ; n15940
g15749 and asqrt[13] n15940 ; n15941
g15750 nor n15306 n15315 ; n15942
g15751 and asqrt[13] n15942 ; n15943
g15752 nor n15313 n15943 ; n15944
g15753 nor n15941 n15944 ; n15945
g15754 nor asqrt[20] n15926 ; n15946
g15755 and n15936_not n15946 ; n15947
g15756 nor n15945 n15947 ; n15948
g15757 nor n15938 n15948 ; n15949
g15758 and asqrt[21] n15949_not ; n15950
g15759 and n15325 n15327_not ; n15951
g15760 and n15318_not n15951 ; n15952
g15761 and asqrt[13] n15952 ; n15953
g15762 nor n15318 n15327 ; n15954
g15763 and asqrt[13] n15954 ; n15955
g15764 nor n15325 n15955 ; n15956
g15765 nor n15953 n15956 ; n15957
g15766 nor asqrt[21] n15938 ; n15958
g15767 and n15948_not n15958 ; n15959
g15768 nor n15957 n15959 ; n15960
g15769 nor n15950 n15960 ; n15961
g15770 and asqrt[22] n15961_not ; n15962
g15771 and n15330_not n15337 ; n15963
g15772 and n15339_not n15963 ; n15964
g15773 and asqrt[13] n15964 ; n15965
g15774 nor n15330 n15339 ; n15966
g15775 and asqrt[13] n15966 ; n15967
g15776 nor n15337 n15967 ; n15968
g15777 nor n15965 n15968 ; n15969
g15778 nor asqrt[22] n15950 ; n15970
g15779 and n15960_not n15970 ; n15971
g15780 nor n15969 n15971 ; n15972
g15781 nor n15962 n15972 ; n15973
g15782 and asqrt[23] n15973_not ; n15974
g15783 and n15349 n15351_not ; n15975
g15784 and n15342_not n15975 ; n15976
g15785 and asqrt[13] n15976 ; n15977
g15786 nor n15342 n15351 ; n15978
g15787 and asqrt[13] n15978 ; n15979
g15788 nor n15349 n15979 ; n15980
g15789 nor n15977 n15980 ; n15981
g15790 nor asqrt[23] n15962 ; n15982
g15791 and n15972_not n15982 ; n15983
g15792 nor n15981 n15983 ; n15984
g15793 nor n15974 n15984 ; n15985
g15794 and asqrt[24] n15985_not ; n15986
g15795 and n15354_not n15361 ; n15987
g15796 and n15363_not n15987 ; n15988
g15797 and asqrt[13] n15988 ; n15989
g15798 nor n15354 n15363 ; n15990
g15799 and asqrt[13] n15990 ; n15991
g15800 nor n15361 n15991 ; n15992
g15801 nor n15989 n15992 ; n15993
g15802 nor asqrt[24] n15974 ; n15994
g15803 and n15984_not n15994 ; n15995
g15804 nor n15993 n15995 ; n15996
g15805 nor n15986 n15996 ; n15997
g15806 and asqrt[25] n15997_not ; n15998
g15807 and n15373 n15375_not ; n15999
g15808 and n15366_not n15999 ; n16000
g15809 and asqrt[13] n16000 ; n16001
g15810 nor n15366 n15375 ; n16002
g15811 and asqrt[13] n16002 ; n16003
g15812 nor n15373 n16003 ; n16004
g15813 nor n16001 n16004 ; n16005
g15814 nor asqrt[25] n15986 ; n16006
g15815 and n15996_not n16006 ; n16007
g15816 nor n16005 n16007 ; n16008
g15817 nor n15998 n16008 ; n16009
g15818 and asqrt[26] n16009_not ; n16010
g15819 and n15378_not n15385 ; n16011
g15820 and n15387_not n16011 ; n16012
g15821 and asqrt[13] n16012 ; n16013
g15822 nor n15378 n15387 ; n16014
g15823 and asqrt[13] n16014 ; n16015
g15824 nor n15385 n16015 ; n16016
g15825 nor n16013 n16016 ; n16017
g15826 nor asqrt[26] n15998 ; n16018
g15827 and n16008_not n16018 ; n16019
g15828 nor n16017 n16019 ; n16020
g15829 nor n16010 n16020 ; n16021
g15830 and asqrt[27] n16021_not ; n16022
g15831 and n15397 n15399_not ; n16023
g15832 and n15390_not n16023 ; n16024
g15833 and asqrt[13] n16024 ; n16025
g15834 nor n15390 n15399 ; n16026
g15835 and asqrt[13] n16026 ; n16027
g15836 nor n15397 n16027 ; n16028
g15837 nor n16025 n16028 ; n16029
g15838 nor asqrt[27] n16010 ; n16030
g15839 and n16020_not n16030 ; n16031
g15840 nor n16029 n16031 ; n16032
g15841 nor n16022 n16032 ; n16033
g15842 and asqrt[28] n16033_not ; n16034
g15843 and n15402_not n15409 ; n16035
g15844 and n15411_not n16035 ; n16036
g15845 and asqrt[13] n16036 ; n16037
g15846 nor n15402 n15411 ; n16038
g15847 and asqrt[13] n16038 ; n16039
g15848 nor n15409 n16039 ; n16040
g15849 nor n16037 n16040 ; n16041
g15850 nor asqrt[28] n16022 ; n16042
g15851 and n16032_not n16042 ; n16043
g15852 nor n16041 n16043 ; n16044
g15853 nor n16034 n16044 ; n16045
g15854 and asqrt[29] n16045_not ; n16046
g15855 and n15421 n15423_not ; n16047
g15856 and n15414_not n16047 ; n16048
g15857 and asqrt[13] n16048 ; n16049
g15858 nor n15414 n15423 ; n16050
g15859 and asqrt[13] n16050 ; n16051
g15860 nor n15421 n16051 ; n16052
g15861 nor n16049 n16052 ; n16053
g15862 nor asqrt[29] n16034 ; n16054
g15863 and n16044_not n16054 ; n16055
g15864 nor n16053 n16055 ; n16056
g15865 nor n16046 n16056 ; n16057
g15866 and asqrt[30] n16057_not ; n16058
g15867 and n15426_not n15433 ; n16059
g15868 and n15435_not n16059 ; n16060
g15869 and asqrt[13] n16060 ; n16061
g15870 nor n15426 n15435 ; n16062
g15871 and asqrt[13] n16062 ; n16063
g15872 nor n15433 n16063 ; n16064
g15873 nor n16061 n16064 ; n16065
g15874 nor asqrt[30] n16046 ; n16066
g15875 and n16056_not n16066 ; n16067
g15876 nor n16065 n16067 ; n16068
g15877 nor n16058 n16068 ; n16069
g15878 and asqrt[31] n16069_not ; n16070
g15879 and n15445 n15447_not ; n16071
g15880 and n15438_not n16071 ; n16072
g15881 and asqrt[13] n16072 ; n16073
g15882 nor n15438 n15447 ; n16074
g15883 and asqrt[13] n16074 ; n16075
g15884 nor n15445 n16075 ; n16076
g15885 nor n16073 n16076 ; n16077
g15886 nor asqrt[31] n16058 ; n16078
g15887 and n16068_not n16078 ; n16079
g15888 nor n16077 n16079 ; n16080
g15889 nor n16070 n16080 ; n16081
g15890 and asqrt[32] n16081_not ; n16082
g15891 and n15450_not n15457 ; n16083
g15892 and n15459_not n16083 ; n16084
g15893 and asqrt[13] n16084 ; n16085
g15894 nor n15450 n15459 ; n16086
g15895 and asqrt[13] n16086 ; n16087
g15896 nor n15457 n16087 ; n16088
g15897 nor n16085 n16088 ; n16089
g15898 nor asqrt[32] n16070 ; n16090
g15899 and n16080_not n16090 ; n16091
g15900 nor n16089 n16091 ; n16092
g15901 nor n16082 n16092 ; n16093
g15902 and asqrt[33] n16093_not ; n16094
g15903 and n15469 n15471_not ; n16095
g15904 and n15462_not n16095 ; n16096
g15905 and asqrt[13] n16096 ; n16097
g15906 nor n15462 n15471 ; n16098
g15907 and asqrt[13] n16098 ; n16099
g15908 nor n15469 n16099 ; n16100
g15909 nor n16097 n16100 ; n16101
g15910 nor asqrt[33] n16082 ; n16102
g15911 and n16092_not n16102 ; n16103
g15912 nor n16101 n16103 ; n16104
g15913 nor n16094 n16104 ; n16105
g15914 and asqrt[34] n16105_not ; n16106
g15915 and n15474_not n15481 ; n16107
g15916 and n15483_not n16107 ; n16108
g15917 and asqrt[13] n16108 ; n16109
g15918 nor n15474 n15483 ; n16110
g15919 and asqrt[13] n16110 ; n16111
g15920 nor n15481 n16111 ; n16112
g15921 nor n16109 n16112 ; n16113
g15922 nor asqrt[34] n16094 ; n16114
g15923 and n16104_not n16114 ; n16115
g15924 nor n16113 n16115 ; n16116
g15925 nor n16106 n16116 ; n16117
g15926 and asqrt[35] n16117_not ; n16118
g15927 and n15493 n15495_not ; n16119
g15928 and n15486_not n16119 ; n16120
g15929 and asqrt[13] n16120 ; n16121
g15930 nor n15486 n15495 ; n16122
g15931 and asqrt[13] n16122 ; n16123
g15932 nor n15493 n16123 ; n16124
g15933 nor n16121 n16124 ; n16125
g15934 nor asqrt[35] n16106 ; n16126
g15935 and n16116_not n16126 ; n16127
g15936 nor n16125 n16127 ; n16128
g15937 nor n16118 n16128 ; n16129
g15938 and asqrt[36] n16129_not ; n16130
g15939 and n15498_not n15505 ; n16131
g15940 and n15507_not n16131 ; n16132
g15941 and asqrt[13] n16132 ; n16133
g15942 nor n15498 n15507 ; n16134
g15943 and asqrt[13] n16134 ; n16135
g15944 nor n15505 n16135 ; n16136
g15945 nor n16133 n16136 ; n16137
g15946 nor asqrt[36] n16118 ; n16138
g15947 and n16128_not n16138 ; n16139
g15948 nor n16137 n16139 ; n16140
g15949 nor n16130 n16140 ; n16141
g15950 and asqrt[37] n16141_not ; n16142
g15951 and n15517 n15519_not ; n16143
g15952 and n15510_not n16143 ; n16144
g15953 and asqrt[13] n16144 ; n16145
g15954 nor n15510 n15519 ; n16146
g15955 and asqrt[13] n16146 ; n16147
g15956 nor n15517 n16147 ; n16148
g15957 nor n16145 n16148 ; n16149
g15958 nor asqrt[37] n16130 ; n16150
g15959 and n16140_not n16150 ; n16151
g15960 nor n16149 n16151 ; n16152
g15961 nor n16142 n16152 ; n16153
g15962 and asqrt[38] n16153_not ; n16154
g15963 and n15522_not n15529 ; n16155
g15964 and n15531_not n16155 ; n16156
g15965 and asqrt[13] n16156 ; n16157
g15966 nor n15522 n15531 ; n16158
g15967 and asqrt[13] n16158 ; n16159
g15968 nor n15529 n16159 ; n16160
g15969 nor n16157 n16160 ; n16161
g15970 nor asqrt[38] n16142 ; n16162
g15971 and n16152_not n16162 ; n16163
g15972 nor n16161 n16163 ; n16164
g15973 nor n16154 n16164 ; n16165
g15974 and asqrt[39] n16165_not ; n16166
g15975 and n15541 n15543_not ; n16167
g15976 and n15534_not n16167 ; n16168
g15977 and asqrt[13] n16168 ; n16169
g15978 nor n15534 n15543 ; n16170
g15979 and asqrt[13] n16170 ; n16171
g15980 nor n15541 n16171 ; n16172
g15981 nor n16169 n16172 ; n16173
g15982 nor asqrt[39] n16154 ; n16174
g15983 and n16164_not n16174 ; n16175
g15984 nor n16173 n16175 ; n16176
g15985 nor n16166 n16176 ; n16177
g15986 and asqrt[40] n16177_not ; n16178
g15987 and n15546_not n15553 ; n16179
g15988 and n15555_not n16179 ; n16180
g15989 and asqrt[13] n16180 ; n16181
g15990 nor n15546 n15555 ; n16182
g15991 and asqrt[13] n16182 ; n16183
g15992 nor n15553 n16183 ; n16184
g15993 nor n16181 n16184 ; n16185
g15994 nor asqrt[40] n16166 ; n16186
g15995 and n16176_not n16186 ; n16187
g15996 nor n16185 n16187 ; n16188
g15997 nor n16178 n16188 ; n16189
g15998 and asqrt[41] n16189_not ; n16190
g15999 and n15565 n15567_not ; n16191
g16000 and n15558_not n16191 ; n16192
g16001 and asqrt[13] n16192 ; n16193
g16002 nor n15558 n15567 ; n16194
g16003 and asqrt[13] n16194 ; n16195
g16004 nor n15565 n16195 ; n16196
g16005 nor n16193 n16196 ; n16197
g16006 nor asqrt[41] n16178 ; n16198
g16007 and n16188_not n16198 ; n16199
g16008 nor n16197 n16199 ; n16200
g16009 nor n16190 n16200 ; n16201
g16010 and asqrt[42] n16201_not ; n16202
g16011 and n15570_not n15577 ; n16203
g16012 and n15579_not n16203 ; n16204
g16013 and asqrt[13] n16204 ; n16205
g16014 nor n15570 n15579 ; n16206
g16015 and asqrt[13] n16206 ; n16207
g16016 nor n15577 n16207 ; n16208
g16017 nor n16205 n16208 ; n16209
g16018 nor asqrt[42] n16190 ; n16210
g16019 and n16200_not n16210 ; n16211
g16020 nor n16209 n16211 ; n16212
g16021 nor n16202 n16212 ; n16213
g16022 and asqrt[43] n16213_not ; n16214
g16023 and n15589 n15591_not ; n16215
g16024 and n15582_not n16215 ; n16216
g16025 and asqrt[13] n16216 ; n16217
g16026 nor n15582 n15591 ; n16218
g16027 and asqrt[13] n16218 ; n16219
g16028 nor n15589 n16219 ; n16220
g16029 nor n16217 n16220 ; n16221
g16030 nor asqrt[43] n16202 ; n16222
g16031 and n16212_not n16222 ; n16223
g16032 nor n16221 n16223 ; n16224
g16033 nor n16214 n16224 ; n16225
g16034 and asqrt[44] n16225_not ; n16226
g16035 and n15594_not n15601 ; n16227
g16036 and n15603_not n16227 ; n16228
g16037 and asqrt[13] n16228 ; n16229
g16038 nor n15594 n15603 ; n16230
g16039 and asqrt[13] n16230 ; n16231
g16040 nor n15601 n16231 ; n16232
g16041 nor n16229 n16232 ; n16233
g16042 nor asqrt[44] n16214 ; n16234
g16043 and n16224_not n16234 ; n16235
g16044 nor n16233 n16235 ; n16236
g16045 nor n16226 n16236 ; n16237
g16046 and asqrt[45] n16237_not ; n16238
g16047 and n15613 n15615_not ; n16239
g16048 and n15606_not n16239 ; n16240
g16049 and asqrt[13] n16240 ; n16241
g16050 nor n15606 n15615 ; n16242
g16051 and asqrt[13] n16242 ; n16243
g16052 nor n15613 n16243 ; n16244
g16053 nor n16241 n16244 ; n16245
g16054 nor asqrt[45] n16226 ; n16246
g16055 and n16236_not n16246 ; n16247
g16056 nor n16245 n16247 ; n16248
g16057 nor n16238 n16248 ; n16249
g16058 and asqrt[46] n16249_not ; n16250
g16059 and n15618_not n15625 ; n16251
g16060 and n15627_not n16251 ; n16252
g16061 and asqrt[13] n16252 ; n16253
g16062 nor n15618 n15627 ; n16254
g16063 and asqrt[13] n16254 ; n16255
g16064 nor n15625 n16255 ; n16256
g16065 nor n16253 n16256 ; n16257
g16066 nor asqrt[46] n16238 ; n16258
g16067 and n16248_not n16258 ; n16259
g16068 nor n16257 n16259 ; n16260
g16069 nor n16250 n16260 ; n16261
g16070 and asqrt[47] n16261_not ; n16262
g16071 and n15637 n15639_not ; n16263
g16072 and n15630_not n16263 ; n16264
g16073 and asqrt[13] n16264 ; n16265
g16074 nor n15630 n15639 ; n16266
g16075 and asqrt[13] n16266 ; n16267
g16076 nor n15637 n16267 ; n16268
g16077 nor n16265 n16268 ; n16269
g16078 nor asqrt[47] n16250 ; n16270
g16079 and n16260_not n16270 ; n16271
g16080 nor n16269 n16271 ; n16272
g16081 nor n16262 n16272 ; n16273
g16082 and asqrt[48] n16273_not ; n16274
g16083 and n15642_not n15649 ; n16275
g16084 and n15651_not n16275 ; n16276
g16085 and asqrt[13] n16276 ; n16277
g16086 nor n15642 n15651 ; n16278
g16087 and asqrt[13] n16278 ; n16279
g16088 nor n15649 n16279 ; n16280
g16089 nor n16277 n16280 ; n16281
g16090 nor asqrt[48] n16262 ; n16282
g16091 and n16272_not n16282 ; n16283
g16092 nor n16281 n16283 ; n16284
g16093 nor n16274 n16284 ; n16285
g16094 and asqrt[49] n16285_not ; n16286
g16095 and n15661 n15663_not ; n16287
g16096 and n15654_not n16287 ; n16288
g16097 and asqrt[13] n16288 ; n16289
g16098 nor n15654 n15663 ; n16290
g16099 and asqrt[13] n16290 ; n16291
g16100 nor n15661 n16291 ; n16292
g16101 nor n16289 n16292 ; n16293
g16102 nor asqrt[49] n16274 ; n16294
g16103 and n16284_not n16294 ; n16295
g16104 nor n16293 n16295 ; n16296
g16105 nor n16286 n16296 ; n16297
g16106 and asqrt[50] n16297_not ; n16298
g16107 and n15666_not n15673 ; n16299
g16108 and n15675_not n16299 ; n16300
g16109 and asqrt[13] n16300 ; n16301
g16110 nor n15666 n15675 ; n16302
g16111 and asqrt[13] n16302 ; n16303
g16112 nor n15673 n16303 ; n16304
g16113 nor n16301 n16304 ; n16305
g16114 nor asqrt[50] n16286 ; n16306
g16115 and n16296_not n16306 ; n16307
g16116 nor n16305 n16307 ; n16308
g16117 nor n16298 n16308 ; n16309
g16118 and asqrt[51] n16309_not ; n16310
g16119 and n15685 n15687_not ; n16311
g16120 and n15678_not n16311 ; n16312
g16121 and asqrt[13] n16312 ; n16313
g16122 nor n15678 n15687 ; n16314
g16123 and asqrt[13] n16314 ; n16315
g16124 nor n15685 n16315 ; n16316
g16125 nor n16313 n16316 ; n16317
g16126 nor asqrt[51] n16298 ; n16318
g16127 and n16308_not n16318 ; n16319
g16128 nor n16317 n16319 ; n16320
g16129 nor n16310 n16320 ; n16321
g16130 and asqrt[52] n16321_not ; n16322
g16131 nor asqrt[52] n16310 ; n16323
g16132 and n16320_not n16323 ; n16324
g16133 and n15690_not n15699 ; n16325
g16134 and n15692_not n16325 ; n16326
g16135 and asqrt[13] n16326 ; n16327
g16136 nor n15690 n15692 ; n16328
g16137 and asqrt[13] n16328 ; n16329
g16138 nor n15699 n16329 ; n16330
g16139 nor n16327 n16330 ; n16331
g16140 nor n16324 n16331 ; n16332
g16141 nor n16322 n16332 ; n16333
g16142 and asqrt[53] n16333_not ; n16334
g16143 and n15709 n15711_not ; n16335
g16144 and n15702_not n16335 ; n16336
g16145 and asqrt[13] n16336 ; n16337
g16146 nor n15702 n15711 ; n16338
g16147 and asqrt[13] n16338 ; n16339
g16148 nor n15709 n16339 ; n16340
g16149 nor n16337 n16340 ; n16341
g16150 nor asqrt[53] n16322 ; n16342
g16151 and n16332_not n16342 ; n16343
g16152 nor n16341 n16343 ; n16344
g16153 nor n16334 n16344 ; n16345
g16154 and asqrt[54] n16345_not ; n16346
g16155 and n15714_not n15721 ; n16347
g16156 and n15723_not n16347 ; n16348
g16157 and asqrt[13] n16348 ; n16349
g16158 nor n15714 n15723 ; n16350
g16159 and asqrt[13] n16350 ; n16351
g16160 nor n15721 n16351 ; n16352
g16161 nor n16349 n16352 ; n16353
g16162 nor asqrt[54] n16334 ; n16354
g16163 and n16344_not n16354 ; n16355
g16164 nor n16353 n16355 ; n16356
g16165 nor n16346 n16356 ; n16357
g16166 and asqrt[55] n16357_not ; n16358
g16167 and n15733 n15735_not ; n16359
g16168 and n15726_not n16359 ; n16360
g16169 and asqrt[13] n16360 ; n16361
g16170 nor n15726 n15735 ; n16362
g16171 and asqrt[13] n16362 ; n16363
g16172 nor n15733 n16363 ; n16364
g16173 nor n16361 n16364 ; n16365
g16174 nor asqrt[55] n16346 ; n16366
g16175 and n16356_not n16366 ; n16367
g16176 nor n16365 n16367 ; n16368
g16177 nor n16358 n16368 ; n16369
g16178 and asqrt[56] n16369_not ; n16370
g16179 and n15738_not n15745 ; n16371
g16180 and n15747_not n16371 ; n16372
g16181 and asqrt[13] n16372 ; n16373
g16182 nor n15738 n15747 ; n16374
g16183 and asqrt[13] n16374 ; n16375
g16184 nor n15745 n16375 ; n16376
g16185 nor n16373 n16376 ; n16377
g16186 nor asqrt[56] n16358 ; n16378
g16187 and n16368_not n16378 ; n16379
g16188 nor n16377 n16379 ; n16380
g16189 nor n16370 n16380 ; n16381
g16190 and asqrt[57] n16381_not ; n16382
g16191 and n15757 n15759_not ; n16383
g16192 and n15750_not n16383 ; n16384
g16193 and asqrt[13] n16384 ; n16385
g16194 nor n15750 n15759 ; n16386
g16195 and asqrt[13] n16386 ; n16387
g16196 nor n15757 n16387 ; n16388
g16197 nor n16385 n16388 ; n16389
g16198 nor asqrt[57] n16370 ; n16390
g16199 and n16380_not n16390 ; n16391
g16200 nor n16389 n16391 ; n16392
g16201 nor n16382 n16392 ; n16393
g16202 and asqrt[58] n16393_not ; n16394
g16203 and n15762_not n15769 ; n16395
g16204 and n15771_not n16395 ; n16396
g16205 and asqrt[13] n16396 ; n16397
g16206 nor n15762 n15771 ; n16398
g16207 and asqrt[13] n16398 ; n16399
g16208 nor n15769 n16399 ; n16400
g16209 nor n16397 n16400 ; n16401
g16210 nor asqrt[58] n16382 ; n16402
g16211 and n16392_not n16402 ; n16403
g16212 nor n16401 n16403 ; n16404
g16213 nor n16394 n16404 ; n16405
g16214 and asqrt[59] n16405_not ; n16406
g16215 and n15781 n15783_not ; n16407
g16216 and n15774_not n16407 ; n16408
g16217 and asqrt[13] n16408 ; n16409
g16218 nor n15774 n15783 ; n16410
g16219 and asqrt[13] n16410 ; n16411
g16220 nor n15781 n16411 ; n16412
g16221 nor n16409 n16412 ; n16413
g16222 nor asqrt[59] n16394 ; n16414
g16223 and n16404_not n16414 ; n16415
g16224 nor n16413 n16415 ; n16416
g16225 nor n16406 n16416 ; n16417
g16226 and asqrt[60] n16417_not ; n16418
g16227 and n15786_not n15793 ; n16419
g16228 and n15795_not n16419 ; n16420
g16229 and asqrt[13] n16420 ; n16421
g16230 nor n15786 n15795 ; n16422
g16231 and asqrt[13] n16422 ; n16423
g16232 nor n15793 n16423 ; n16424
g16233 nor n16421 n16424 ; n16425
g16234 nor asqrt[60] n16406 ; n16426
g16235 and n16416_not n16426 ; n16427
g16236 nor n16425 n16427 ; n16428
g16237 nor n16418 n16428 ; n16429
g16238 and asqrt[61] n16429_not ; n16430
g16239 and n15805 n15807_not ; n16431
g16240 and n15798_not n16431 ; n16432
g16241 and asqrt[13] n16432 ; n16433
g16242 nor n15798 n15807 ; n16434
g16243 and asqrt[13] n16434 ; n16435
g16244 nor n15805 n16435 ; n16436
g16245 nor n16433 n16436 ; n16437
g16246 nor asqrt[61] n16418 ; n16438
g16247 and n16428_not n16438 ; n16439
g16248 nor n16437 n16439 ; n16440
g16249 nor n16430 n16440 ; n16441
g16250 and asqrt[62] n16441_not ; n16442
g16251 and n15810_not n15817 ; n16443
g16252 and n15819_not n16443 ; n16444
g16253 and asqrt[13] n16444 ; n16445
g16254 nor n15810 n15819 ; n16446
g16255 and asqrt[13] n16446 ; n16447
g16256 nor n15817 n16447 ; n16448
g16257 nor n16445 n16448 ; n16449
g16258 nor asqrt[62] n16430 ; n16450
g16259 and n16440_not n16450 ; n16451
g16260 nor n16449 n16451 ; n16452
g16261 nor n16442 n16452 ; n16453
g16262 and n15829 n15831_not ; n16454
g16263 and n15822_not n16454 ; n16455
g16264 and asqrt[13] n16455 ; n16456
g16265 nor n15822 n15831 ; n16457
g16266 and asqrt[13] n16457 ; n16458
g16267 nor n15829 n16458 ; n16459
g16268 nor n16456 n16459 ; n16460
g16269 nor n15833 n15840 ; n16461
g16270 and asqrt[13] n16461 ; n16462
g16271 nor n15848 n16462 ; n16463
g16272 and n16460_not n16463 ; n16464
g16273 and n16453_not n16464 ; n16465
g16274 nor asqrt[63] n16465 ; n16466
g16275 and n16442_not n16460 ; n16467
g16276 and n16452_not n16467 ; n16468
g16277 and n15840_not asqrt[13] ; n16469
g16278 and n15833 n16469_not ; n16470
g16279 and asqrt[63] n16461_not ; n16471
g16280 and n16470_not n16471 ; n16472
g16281 nor n15836 n15857 ; n16473
g16282 and n15839_not n16473 ; n16474
g16283 and n15852_not n16474 ; n16475
g16284 and n15848_not n16475 ; n16476
g16285 and n15846_not n16476 ; n16477
g16286 nor n16472 n16477 ; n16478
g16287 and n16468_not n16478 ; n16479
g16288 nand n16466_not n16479 ; asqrt[12]
g16289 and a[24] asqrt[12] ; n16481
g16290 nor a[22] a[23] ; n16482
g16291 and a[24]_not n16482 ; n16483
g16292 nor n16481 n16483 ; n16484
g16293 and asqrt[13] n16484_not ; n16485
g16294 nor n15857 n16483 ; n16486
g16295 and n15852_not n16486 ; n16487
g16296 and n15848_not n16487 ; n16488
g16297 and n15846_not n16488 ; n16489
g16298 and n16481_not n16489 ; n16490
g16299 and a[24]_not asqrt[12] ; n16491
g16300 and a[25] n16491_not ; n16492
g16301 and n15862 asqrt[12] ; n16493
g16302 nor n16492 n16493 ; n16494
g16303 and n16490_not n16494 ; n16495
g16304 nor n16485 n16495 ; n16496
g16305 and asqrt[14] n16496_not ; n16497
g16306 nor asqrt[14] n16485 ; n16498
g16307 and n16495_not n16498 ; n16499
g16308 and asqrt[13] n16477_not ; n16500
g16309 and n16472_not n16500 ; n16501
g16310 and n16468_not n16501 ; n16502
g16311 and n16466_not n16502 ; n16503
g16312 nor n16493 n16503 ; n16504
g16313 and a[26] n16504_not ; n16505
g16314 nor a[26] n16503 ; n16506
g16315 and n16493_not n16506 ; n16507
g16316 nor n16505 n16507 ; n16508
g16317 nor n16499 n16508 ; n16509
g16318 nor n16497 n16509 ; n16510
g16319 and asqrt[15] n16510_not ; n16511
g16320 nor n15865 n15870 ; n16512
g16321 and n15874_not n16512 ; n16513
g16322 and asqrt[12] n16513 ; n16514
g16323 and asqrt[12] n16512 ; n16515
g16324 and n15874 n16515_not ; n16516
g16325 nor n16514 n16516 ; n16517
g16326 nor asqrt[15] n16497 ; n16518
g16327 and n16509_not n16518 ; n16519
g16328 nor n16517 n16519 ; n16520
g16329 nor n16511 n16520 ; n16521
g16330 and asqrt[16] n16521_not ; n16522
g16331 and n15879_not n15888 ; n16523
g16332 and n15877_not n16523 ; n16524
g16333 and asqrt[12] n16524 ; n16525
g16334 nor n15877 n15879 ; n16526
g16335 and asqrt[12] n16526 ; n16527
g16336 nor n15888 n16527 ; n16528
g16337 nor n16525 n16528 ; n16529
g16338 nor asqrt[16] n16511 ; n16530
g16339 and n16520_not n16530 ; n16531
g16340 nor n16529 n16531 ; n16532
g16341 nor n16522 n16532 ; n16533
g16342 and asqrt[17] n16533_not ; n16534
g16343 and n15891_not n15897 ; n16535
g16344 and n15899_not n16535 ; n16536
g16345 and asqrt[12] n16536 ; n16537
g16346 nor n15891 n15899 ; n16538
g16347 and asqrt[12] n16538 ; n16539
g16348 nor n15897 n16539 ; n16540
g16349 nor n16537 n16540 ; n16541
g16350 nor asqrt[17] n16522 ; n16542
g16351 and n16532_not n16542 ; n16543
g16352 nor n16541 n16543 ; n16544
g16353 nor n16534 n16544 ; n16545
g16354 and asqrt[18] n16545_not ; n16546
g16355 and n15909 n15911_not ; n16547
g16356 and n15902_not n16547 ; n16548
g16357 and asqrt[12] n16548 ; n16549
g16358 nor n15902 n15911 ; n16550
g16359 and asqrt[12] n16550 ; n16551
g16360 nor n15909 n16551 ; n16552
g16361 nor n16549 n16552 ; n16553
g16362 nor asqrt[18] n16534 ; n16554
g16363 and n16544_not n16554 ; n16555
g16364 nor n16553 n16555 ; n16556
g16365 nor n16546 n16556 ; n16557
g16366 and asqrt[19] n16557_not ; n16558
g16367 and n15914_not n15921 ; n16559
g16368 and n15923_not n16559 ; n16560
g16369 and asqrt[12] n16560 ; n16561
g16370 nor n15914 n15923 ; n16562
g16371 and asqrt[12] n16562 ; n16563
g16372 nor n15921 n16563 ; n16564
g16373 nor n16561 n16564 ; n16565
g16374 nor asqrt[19] n16546 ; n16566
g16375 and n16556_not n16566 ; n16567
g16376 nor n16565 n16567 ; n16568
g16377 nor n16558 n16568 ; n16569
g16378 and asqrt[20] n16569_not ; n16570
g16379 and n15933 n15935_not ; n16571
g16380 and n15926_not n16571 ; n16572
g16381 and asqrt[12] n16572 ; n16573
g16382 nor n15926 n15935 ; n16574
g16383 and asqrt[12] n16574 ; n16575
g16384 nor n15933 n16575 ; n16576
g16385 nor n16573 n16576 ; n16577
g16386 nor asqrt[20] n16558 ; n16578
g16387 and n16568_not n16578 ; n16579
g16388 nor n16577 n16579 ; n16580
g16389 nor n16570 n16580 ; n16581
g16390 and asqrt[21] n16581_not ; n16582
g16391 and n15938_not n15945 ; n16583
g16392 and n15947_not n16583 ; n16584
g16393 and asqrt[12] n16584 ; n16585
g16394 nor n15938 n15947 ; n16586
g16395 and asqrt[12] n16586 ; n16587
g16396 nor n15945 n16587 ; n16588
g16397 nor n16585 n16588 ; n16589
g16398 nor asqrt[21] n16570 ; n16590
g16399 and n16580_not n16590 ; n16591
g16400 nor n16589 n16591 ; n16592
g16401 nor n16582 n16592 ; n16593
g16402 and asqrt[22] n16593_not ; n16594
g16403 and n15957 n15959_not ; n16595
g16404 and n15950_not n16595 ; n16596
g16405 and asqrt[12] n16596 ; n16597
g16406 nor n15950 n15959 ; n16598
g16407 and asqrt[12] n16598 ; n16599
g16408 nor n15957 n16599 ; n16600
g16409 nor n16597 n16600 ; n16601
g16410 nor asqrt[22] n16582 ; n16602
g16411 and n16592_not n16602 ; n16603
g16412 nor n16601 n16603 ; n16604
g16413 nor n16594 n16604 ; n16605
g16414 and asqrt[23] n16605_not ; n16606
g16415 and n15962_not n15969 ; n16607
g16416 and n15971_not n16607 ; n16608
g16417 and asqrt[12] n16608 ; n16609
g16418 nor n15962 n15971 ; n16610
g16419 and asqrt[12] n16610 ; n16611
g16420 nor n15969 n16611 ; n16612
g16421 nor n16609 n16612 ; n16613
g16422 nor asqrt[23] n16594 ; n16614
g16423 and n16604_not n16614 ; n16615
g16424 nor n16613 n16615 ; n16616
g16425 nor n16606 n16616 ; n16617
g16426 and asqrt[24] n16617_not ; n16618
g16427 and n15981 n15983_not ; n16619
g16428 and n15974_not n16619 ; n16620
g16429 and asqrt[12] n16620 ; n16621
g16430 nor n15974 n15983 ; n16622
g16431 and asqrt[12] n16622 ; n16623
g16432 nor n15981 n16623 ; n16624
g16433 nor n16621 n16624 ; n16625
g16434 nor asqrt[24] n16606 ; n16626
g16435 and n16616_not n16626 ; n16627
g16436 nor n16625 n16627 ; n16628
g16437 nor n16618 n16628 ; n16629
g16438 and asqrt[25] n16629_not ; n16630
g16439 and n15986_not n15993 ; n16631
g16440 and n15995_not n16631 ; n16632
g16441 and asqrt[12] n16632 ; n16633
g16442 nor n15986 n15995 ; n16634
g16443 and asqrt[12] n16634 ; n16635
g16444 nor n15993 n16635 ; n16636
g16445 nor n16633 n16636 ; n16637
g16446 nor asqrt[25] n16618 ; n16638
g16447 and n16628_not n16638 ; n16639
g16448 nor n16637 n16639 ; n16640
g16449 nor n16630 n16640 ; n16641
g16450 and asqrt[26] n16641_not ; n16642
g16451 and n16005 n16007_not ; n16643
g16452 and n15998_not n16643 ; n16644
g16453 and asqrt[12] n16644 ; n16645
g16454 nor n15998 n16007 ; n16646
g16455 and asqrt[12] n16646 ; n16647
g16456 nor n16005 n16647 ; n16648
g16457 nor n16645 n16648 ; n16649
g16458 nor asqrt[26] n16630 ; n16650
g16459 and n16640_not n16650 ; n16651
g16460 nor n16649 n16651 ; n16652
g16461 nor n16642 n16652 ; n16653
g16462 and asqrt[27] n16653_not ; n16654
g16463 and n16010_not n16017 ; n16655
g16464 and n16019_not n16655 ; n16656
g16465 and asqrt[12] n16656 ; n16657
g16466 nor n16010 n16019 ; n16658
g16467 and asqrt[12] n16658 ; n16659
g16468 nor n16017 n16659 ; n16660
g16469 nor n16657 n16660 ; n16661
g16470 nor asqrt[27] n16642 ; n16662
g16471 and n16652_not n16662 ; n16663
g16472 nor n16661 n16663 ; n16664
g16473 nor n16654 n16664 ; n16665
g16474 and asqrt[28] n16665_not ; n16666
g16475 and n16029 n16031_not ; n16667
g16476 and n16022_not n16667 ; n16668
g16477 and asqrt[12] n16668 ; n16669
g16478 nor n16022 n16031 ; n16670
g16479 and asqrt[12] n16670 ; n16671
g16480 nor n16029 n16671 ; n16672
g16481 nor n16669 n16672 ; n16673
g16482 nor asqrt[28] n16654 ; n16674
g16483 and n16664_not n16674 ; n16675
g16484 nor n16673 n16675 ; n16676
g16485 nor n16666 n16676 ; n16677
g16486 and asqrt[29] n16677_not ; n16678
g16487 and n16034_not n16041 ; n16679
g16488 and n16043_not n16679 ; n16680
g16489 and asqrt[12] n16680 ; n16681
g16490 nor n16034 n16043 ; n16682
g16491 and asqrt[12] n16682 ; n16683
g16492 nor n16041 n16683 ; n16684
g16493 nor n16681 n16684 ; n16685
g16494 nor asqrt[29] n16666 ; n16686
g16495 and n16676_not n16686 ; n16687
g16496 nor n16685 n16687 ; n16688
g16497 nor n16678 n16688 ; n16689
g16498 and asqrt[30] n16689_not ; n16690
g16499 and n16053 n16055_not ; n16691
g16500 and n16046_not n16691 ; n16692
g16501 and asqrt[12] n16692 ; n16693
g16502 nor n16046 n16055 ; n16694
g16503 and asqrt[12] n16694 ; n16695
g16504 nor n16053 n16695 ; n16696
g16505 nor n16693 n16696 ; n16697
g16506 nor asqrt[30] n16678 ; n16698
g16507 and n16688_not n16698 ; n16699
g16508 nor n16697 n16699 ; n16700
g16509 nor n16690 n16700 ; n16701
g16510 and asqrt[31] n16701_not ; n16702
g16511 and n16058_not n16065 ; n16703
g16512 and n16067_not n16703 ; n16704
g16513 and asqrt[12] n16704 ; n16705
g16514 nor n16058 n16067 ; n16706
g16515 and asqrt[12] n16706 ; n16707
g16516 nor n16065 n16707 ; n16708
g16517 nor n16705 n16708 ; n16709
g16518 nor asqrt[31] n16690 ; n16710
g16519 and n16700_not n16710 ; n16711
g16520 nor n16709 n16711 ; n16712
g16521 nor n16702 n16712 ; n16713
g16522 and asqrt[32] n16713_not ; n16714
g16523 and n16077 n16079_not ; n16715
g16524 and n16070_not n16715 ; n16716
g16525 and asqrt[12] n16716 ; n16717
g16526 nor n16070 n16079 ; n16718
g16527 and asqrt[12] n16718 ; n16719
g16528 nor n16077 n16719 ; n16720
g16529 nor n16717 n16720 ; n16721
g16530 nor asqrt[32] n16702 ; n16722
g16531 and n16712_not n16722 ; n16723
g16532 nor n16721 n16723 ; n16724
g16533 nor n16714 n16724 ; n16725
g16534 and asqrt[33] n16725_not ; n16726
g16535 and n16082_not n16089 ; n16727
g16536 and n16091_not n16727 ; n16728
g16537 and asqrt[12] n16728 ; n16729
g16538 nor n16082 n16091 ; n16730
g16539 and asqrt[12] n16730 ; n16731
g16540 nor n16089 n16731 ; n16732
g16541 nor n16729 n16732 ; n16733
g16542 nor asqrt[33] n16714 ; n16734
g16543 and n16724_not n16734 ; n16735
g16544 nor n16733 n16735 ; n16736
g16545 nor n16726 n16736 ; n16737
g16546 and asqrt[34] n16737_not ; n16738
g16547 and n16101 n16103_not ; n16739
g16548 and n16094_not n16739 ; n16740
g16549 and asqrt[12] n16740 ; n16741
g16550 nor n16094 n16103 ; n16742
g16551 and asqrt[12] n16742 ; n16743
g16552 nor n16101 n16743 ; n16744
g16553 nor n16741 n16744 ; n16745
g16554 nor asqrt[34] n16726 ; n16746
g16555 and n16736_not n16746 ; n16747
g16556 nor n16745 n16747 ; n16748
g16557 nor n16738 n16748 ; n16749
g16558 and asqrt[35] n16749_not ; n16750
g16559 and n16106_not n16113 ; n16751
g16560 and n16115_not n16751 ; n16752
g16561 and asqrt[12] n16752 ; n16753
g16562 nor n16106 n16115 ; n16754
g16563 and asqrt[12] n16754 ; n16755
g16564 nor n16113 n16755 ; n16756
g16565 nor n16753 n16756 ; n16757
g16566 nor asqrt[35] n16738 ; n16758
g16567 and n16748_not n16758 ; n16759
g16568 nor n16757 n16759 ; n16760
g16569 nor n16750 n16760 ; n16761
g16570 and asqrt[36] n16761_not ; n16762
g16571 and n16125 n16127_not ; n16763
g16572 and n16118_not n16763 ; n16764
g16573 and asqrt[12] n16764 ; n16765
g16574 nor n16118 n16127 ; n16766
g16575 and asqrt[12] n16766 ; n16767
g16576 nor n16125 n16767 ; n16768
g16577 nor n16765 n16768 ; n16769
g16578 nor asqrt[36] n16750 ; n16770
g16579 and n16760_not n16770 ; n16771
g16580 nor n16769 n16771 ; n16772
g16581 nor n16762 n16772 ; n16773
g16582 and asqrt[37] n16773_not ; n16774
g16583 and n16130_not n16137 ; n16775
g16584 and n16139_not n16775 ; n16776
g16585 and asqrt[12] n16776 ; n16777
g16586 nor n16130 n16139 ; n16778
g16587 and asqrt[12] n16778 ; n16779
g16588 nor n16137 n16779 ; n16780
g16589 nor n16777 n16780 ; n16781
g16590 nor asqrt[37] n16762 ; n16782
g16591 and n16772_not n16782 ; n16783
g16592 nor n16781 n16783 ; n16784
g16593 nor n16774 n16784 ; n16785
g16594 and asqrt[38] n16785_not ; n16786
g16595 and n16149 n16151_not ; n16787
g16596 and n16142_not n16787 ; n16788
g16597 and asqrt[12] n16788 ; n16789
g16598 nor n16142 n16151 ; n16790
g16599 and asqrt[12] n16790 ; n16791
g16600 nor n16149 n16791 ; n16792
g16601 nor n16789 n16792 ; n16793
g16602 nor asqrt[38] n16774 ; n16794
g16603 and n16784_not n16794 ; n16795
g16604 nor n16793 n16795 ; n16796
g16605 nor n16786 n16796 ; n16797
g16606 and asqrt[39] n16797_not ; n16798
g16607 and n16154_not n16161 ; n16799
g16608 and n16163_not n16799 ; n16800
g16609 and asqrt[12] n16800 ; n16801
g16610 nor n16154 n16163 ; n16802
g16611 and asqrt[12] n16802 ; n16803
g16612 nor n16161 n16803 ; n16804
g16613 nor n16801 n16804 ; n16805
g16614 nor asqrt[39] n16786 ; n16806
g16615 and n16796_not n16806 ; n16807
g16616 nor n16805 n16807 ; n16808
g16617 nor n16798 n16808 ; n16809
g16618 and asqrt[40] n16809_not ; n16810
g16619 and n16173 n16175_not ; n16811
g16620 and n16166_not n16811 ; n16812
g16621 and asqrt[12] n16812 ; n16813
g16622 nor n16166 n16175 ; n16814
g16623 and asqrt[12] n16814 ; n16815
g16624 nor n16173 n16815 ; n16816
g16625 nor n16813 n16816 ; n16817
g16626 nor asqrt[40] n16798 ; n16818
g16627 and n16808_not n16818 ; n16819
g16628 nor n16817 n16819 ; n16820
g16629 nor n16810 n16820 ; n16821
g16630 and asqrt[41] n16821_not ; n16822
g16631 and n16178_not n16185 ; n16823
g16632 and n16187_not n16823 ; n16824
g16633 and asqrt[12] n16824 ; n16825
g16634 nor n16178 n16187 ; n16826
g16635 and asqrt[12] n16826 ; n16827
g16636 nor n16185 n16827 ; n16828
g16637 nor n16825 n16828 ; n16829
g16638 nor asqrt[41] n16810 ; n16830
g16639 and n16820_not n16830 ; n16831
g16640 nor n16829 n16831 ; n16832
g16641 nor n16822 n16832 ; n16833
g16642 and asqrt[42] n16833_not ; n16834
g16643 and n16197 n16199_not ; n16835
g16644 and n16190_not n16835 ; n16836
g16645 and asqrt[12] n16836 ; n16837
g16646 nor n16190 n16199 ; n16838
g16647 and asqrt[12] n16838 ; n16839
g16648 nor n16197 n16839 ; n16840
g16649 nor n16837 n16840 ; n16841
g16650 nor asqrt[42] n16822 ; n16842
g16651 and n16832_not n16842 ; n16843
g16652 nor n16841 n16843 ; n16844
g16653 nor n16834 n16844 ; n16845
g16654 and asqrt[43] n16845_not ; n16846
g16655 and n16202_not n16209 ; n16847
g16656 and n16211_not n16847 ; n16848
g16657 and asqrt[12] n16848 ; n16849
g16658 nor n16202 n16211 ; n16850
g16659 and asqrt[12] n16850 ; n16851
g16660 nor n16209 n16851 ; n16852
g16661 nor n16849 n16852 ; n16853
g16662 nor asqrt[43] n16834 ; n16854
g16663 and n16844_not n16854 ; n16855
g16664 nor n16853 n16855 ; n16856
g16665 nor n16846 n16856 ; n16857
g16666 and asqrt[44] n16857_not ; n16858
g16667 and n16221 n16223_not ; n16859
g16668 and n16214_not n16859 ; n16860
g16669 and asqrt[12] n16860 ; n16861
g16670 nor n16214 n16223 ; n16862
g16671 and asqrt[12] n16862 ; n16863
g16672 nor n16221 n16863 ; n16864
g16673 nor n16861 n16864 ; n16865
g16674 nor asqrt[44] n16846 ; n16866
g16675 and n16856_not n16866 ; n16867
g16676 nor n16865 n16867 ; n16868
g16677 nor n16858 n16868 ; n16869
g16678 and asqrt[45] n16869_not ; n16870
g16679 and n16226_not n16233 ; n16871
g16680 and n16235_not n16871 ; n16872
g16681 and asqrt[12] n16872 ; n16873
g16682 nor n16226 n16235 ; n16874
g16683 and asqrt[12] n16874 ; n16875
g16684 nor n16233 n16875 ; n16876
g16685 nor n16873 n16876 ; n16877
g16686 nor asqrt[45] n16858 ; n16878
g16687 and n16868_not n16878 ; n16879
g16688 nor n16877 n16879 ; n16880
g16689 nor n16870 n16880 ; n16881
g16690 and asqrt[46] n16881_not ; n16882
g16691 and n16245 n16247_not ; n16883
g16692 and n16238_not n16883 ; n16884
g16693 and asqrt[12] n16884 ; n16885
g16694 nor n16238 n16247 ; n16886
g16695 and asqrt[12] n16886 ; n16887
g16696 nor n16245 n16887 ; n16888
g16697 nor n16885 n16888 ; n16889
g16698 nor asqrt[46] n16870 ; n16890
g16699 and n16880_not n16890 ; n16891
g16700 nor n16889 n16891 ; n16892
g16701 nor n16882 n16892 ; n16893
g16702 and asqrt[47] n16893_not ; n16894
g16703 and n16250_not n16257 ; n16895
g16704 and n16259_not n16895 ; n16896
g16705 and asqrt[12] n16896 ; n16897
g16706 nor n16250 n16259 ; n16898
g16707 and asqrt[12] n16898 ; n16899
g16708 nor n16257 n16899 ; n16900
g16709 nor n16897 n16900 ; n16901
g16710 nor asqrt[47] n16882 ; n16902
g16711 and n16892_not n16902 ; n16903
g16712 nor n16901 n16903 ; n16904
g16713 nor n16894 n16904 ; n16905
g16714 and asqrt[48] n16905_not ; n16906
g16715 and n16269 n16271_not ; n16907
g16716 and n16262_not n16907 ; n16908
g16717 and asqrt[12] n16908 ; n16909
g16718 nor n16262 n16271 ; n16910
g16719 and asqrt[12] n16910 ; n16911
g16720 nor n16269 n16911 ; n16912
g16721 nor n16909 n16912 ; n16913
g16722 nor asqrt[48] n16894 ; n16914
g16723 and n16904_not n16914 ; n16915
g16724 nor n16913 n16915 ; n16916
g16725 nor n16906 n16916 ; n16917
g16726 and asqrt[49] n16917_not ; n16918
g16727 and n16274_not n16281 ; n16919
g16728 and n16283_not n16919 ; n16920
g16729 and asqrt[12] n16920 ; n16921
g16730 nor n16274 n16283 ; n16922
g16731 and asqrt[12] n16922 ; n16923
g16732 nor n16281 n16923 ; n16924
g16733 nor n16921 n16924 ; n16925
g16734 nor asqrt[49] n16906 ; n16926
g16735 and n16916_not n16926 ; n16927
g16736 nor n16925 n16927 ; n16928
g16737 nor n16918 n16928 ; n16929
g16738 and asqrt[50] n16929_not ; n16930
g16739 and n16293 n16295_not ; n16931
g16740 and n16286_not n16931 ; n16932
g16741 and asqrt[12] n16932 ; n16933
g16742 nor n16286 n16295 ; n16934
g16743 and asqrt[12] n16934 ; n16935
g16744 nor n16293 n16935 ; n16936
g16745 nor n16933 n16936 ; n16937
g16746 nor asqrt[50] n16918 ; n16938
g16747 and n16928_not n16938 ; n16939
g16748 nor n16937 n16939 ; n16940
g16749 nor n16930 n16940 ; n16941
g16750 and asqrt[51] n16941_not ; n16942
g16751 and n16298_not n16305 ; n16943
g16752 and n16307_not n16943 ; n16944
g16753 and asqrt[12] n16944 ; n16945
g16754 nor n16298 n16307 ; n16946
g16755 and asqrt[12] n16946 ; n16947
g16756 nor n16305 n16947 ; n16948
g16757 nor n16945 n16948 ; n16949
g16758 nor asqrt[51] n16930 ; n16950
g16759 and n16940_not n16950 ; n16951
g16760 nor n16949 n16951 ; n16952
g16761 nor n16942 n16952 ; n16953
g16762 and asqrt[52] n16953_not ; n16954
g16763 and n16317 n16319_not ; n16955
g16764 and n16310_not n16955 ; n16956
g16765 and asqrt[12] n16956 ; n16957
g16766 nor n16310 n16319 ; n16958
g16767 and asqrt[12] n16958 ; n16959
g16768 nor n16317 n16959 ; n16960
g16769 nor n16957 n16960 ; n16961
g16770 nor asqrt[52] n16942 ; n16962
g16771 and n16952_not n16962 ; n16963
g16772 nor n16961 n16963 ; n16964
g16773 nor n16954 n16964 ; n16965
g16774 and asqrt[53] n16965_not ; n16966
g16775 nor asqrt[53] n16954 ; n16967
g16776 and n16964_not n16967 ; n16968
g16777 and n16322_not n16331 ; n16969
g16778 and n16324_not n16969 ; n16970
g16779 and asqrt[12] n16970 ; n16971
g16780 nor n16322 n16324 ; n16972
g16781 and asqrt[12] n16972 ; n16973
g16782 nor n16331 n16973 ; n16974
g16783 nor n16971 n16974 ; n16975
g16784 nor n16968 n16975 ; n16976
g16785 nor n16966 n16976 ; n16977
g16786 and asqrt[54] n16977_not ; n16978
g16787 and n16341 n16343_not ; n16979
g16788 and n16334_not n16979 ; n16980
g16789 and asqrt[12] n16980 ; n16981
g16790 nor n16334 n16343 ; n16982
g16791 and asqrt[12] n16982 ; n16983
g16792 nor n16341 n16983 ; n16984
g16793 nor n16981 n16984 ; n16985
g16794 nor asqrt[54] n16966 ; n16986
g16795 and n16976_not n16986 ; n16987
g16796 nor n16985 n16987 ; n16988
g16797 nor n16978 n16988 ; n16989
g16798 and asqrt[55] n16989_not ; n16990
g16799 and n16346_not n16353 ; n16991
g16800 and n16355_not n16991 ; n16992
g16801 and asqrt[12] n16992 ; n16993
g16802 nor n16346 n16355 ; n16994
g16803 and asqrt[12] n16994 ; n16995
g16804 nor n16353 n16995 ; n16996
g16805 nor n16993 n16996 ; n16997
g16806 nor asqrt[55] n16978 ; n16998
g16807 and n16988_not n16998 ; n16999
g16808 nor n16997 n16999 ; n17000
g16809 nor n16990 n17000 ; n17001
g16810 and asqrt[56] n17001_not ; n17002
g16811 and n16365 n16367_not ; n17003
g16812 and n16358_not n17003 ; n17004
g16813 and asqrt[12] n17004 ; n17005
g16814 nor n16358 n16367 ; n17006
g16815 and asqrt[12] n17006 ; n17007
g16816 nor n16365 n17007 ; n17008
g16817 nor n17005 n17008 ; n17009
g16818 nor asqrt[56] n16990 ; n17010
g16819 and n17000_not n17010 ; n17011
g16820 nor n17009 n17011 ; n17012
g16821 nor n17002 n17012 ; n17013
g16822 and asqrt[57] n17013_not ; n17014
g16823 and n16370_not n16377 ; n17015
g16824 and n16379_not n17015 ; n17016
g16825 and asqrt[12] n17016 ; n17017
g16826 nor n16370 n16379 ; n17018
g16827 and asqrt[12] n17018 ; n17019
g16828 nor n16377 n17019 ; n17020
g16829 nor n17017 n17020 ; n17021
g16830 nor asqrt[57] n17002 ; n17022
g16831 and n17012_not n17022 ; n17023
g16832 nor n17021 n17023 ; n17024
g16833 nor n17014 n17024 ; n17025
g16834 and asqrt[58] n17025_not ; n17026
g16835 and n16389 n16391_not ; n17027
g16836 and n16382_not n17027 ; n17028
g16837 and asqrt[12] n17028 ; n17029
g16838 nor n16382 n16391 ; n17030
g16839 and asqrt[12] n17030 ; n17031
g16840 nor n16389 n17031 ; n17032
g16841 nor n17029 n17032 ; n17033
g16842 nor asqrt[58] n17014 ; n17034
g16843 and n17024_not n17034 ; n17035
g16844 nor n17033 n17035 ; n17036
g16845 nor n17026 n17036 ; n17037
g16846 and asqrt[59] n17037_not ; n17038
g16847 and n16394_not n16401 ; n17039
g16848 and n16403_not n17039 ; n17040
g16849 and asqrt[12] n17040 ; n17041
g16850 nor n16394 n16403 ; n17042
g16851 and asqrt[12] n17042 ; n17043
g16852 nor n16401 n17043 ; n17044
g16853 nor n17041 n17044 ; n17045
g16854 nor asqrt[59] n17026 ; n17046
g16855 and n17036_not n17046 ; n17047
g16856 nor n17045 n17047 ; n17048
g16857 nor n17038 n17048 ; n17049
g16858 and asqrt[60] n17049_not ; n17050
g16859 and n16413 n16415_not ; n17051
g16860 and n16406_not n17051 ; n17052
g16861 and asqrt[12] n17052 ; n17053
g16862 nor n16406 n16415 ; n17054
g16863 and asqrt[12] n17054 ; n17055
g16864 nor n16413 n17055 ; n17056
g16865 nor n17053 n17056 ; n17057
g16866 nor asqrt[60] n17038 ; n17058
g16867 and n17048_not n17058 ; n17059
g16868 nor n17057 n17059 ; n17060
g16869 nor n17050 n17060 ; n17061
g16870 and asqrt[61] n17061_not ; n17062
g16871 and n16418_not n16425 ; n17063
g16872 and n16427_not n17063 ; n17064
g16873 and asqrt[12] n17064 ; n17065
g16874 nor n16418 n16427 ; n17066
g16875 and asqrt[12] n17066 ; n17067
g16876 nor n16425 n17067 ; n17068
g16877 nor n17065 n17068 ; n17069
g16878 nor asqrt[61] n17050 ; n17070
g16879 and n17060_not n17070 ; n17071
g16880 nor n17069 n17071 ; n17072
g16881 nor n17062 n17072 ; n17073
g16882 and asqrt[62] n17073_not ; n17074
g16883 and n16437 n16439_not ; n17075
g16884 and n16430_not n17075 ; n17076
g16885 and asqrt[12] n17076 ; n17077
g16886 nor n16430 n16439 ; n17078
g16887 and asqrt[12] n17078 ; n17079
g16888 nor n16437 n17079 ; n17080
g16889 nor n17077 n17080 ; n17081
g16890 nor asqrt[62] n17062 ; n17082
g16891 and n17072_not n17082 ; n17083
g16892 nor n17081 n17083 ; n17084
g16893 nor n17074 n17084 ; n17085
g16894 and n16442_not n16449 ; n17086
g16895 and n16451_not n17086 ; n17087
g16896 and asqrt[12] n17087 ; n17088
g16897 nor n16442 n16451 ; n17089
g16898 and asqrt[12] n17089 ; n17090
g16899 nor n16449 n17090 ; n17091
g16900 nor n17088 n17091 ; n17092
g16901 nor n16453 n16460 ; n17093
g16902 and asqrt[12] n17093 ; n17094
g16903 nor n16468 n17094 ; n17095
g16904 and n17092_not n17095 ; n17096
g16905 and n17085_not n17096 ; n17097
g16906 nor asqrt[63] n17097 ; n17098
g16907 and n17074_not n17092 ; n17099
g16908 and n17084_not n17099 ; n17100
g16909 and n16460_not asqrt[12] ; n17101
g16910 and n16453 n17101_not ; n17102
g16911 and asqrt[63] n17093_not ; n17103
g16912 and n17102_not n17103 ; n17104
g16913 nor n16456 n16477 ; n17105
g16914 and n16459_not n17105 ; n17106
g16915 and n16472_not n17106 ; n17107
g16916 and n16468_not n17107 ; n17108
g16917 and n16466_not n17108 ; n17109
g16918 nor n17104 n17109 ; n17110
g16919 and n17100_not n17110 ; n17111
g16920 nand n17098_not n17111 ; asqrt[11]
g16921 and a[22] asqrt[11] ; n17113
g16922 nor a[20] a[21] ; n17114
g16923 and a[22]_not n17114 ; n17115
g16924 nor n17113 n17115 ; n17116
g16925 and asqrt[12] n17116_not ; n17117
g16926 nor n16477 n17115 ; n17118
g16927 and n16472_not n17118 ; n17119
g16928 and n16468_not n17119 ; n17120
g16929 and n16466_not n17120 ; n17121
g16930 and n17113_not n17121 ; n17122
g16931 and a[22]_not asqrt[11] ; n17123
g16932 and a[23] n17123_not ; n17124
g16933 and n16482 asqrt[11] ; n17125
g16934 nor n17124 n17125 ; n17126
g16935 and n17122_not n17126 ; n17127
g16936 nor n17117 n17127 ; n17128
g16937 and asqrt[13] n17128_not ; n17129
g16938 nor asqrt[13] n17117 ; n17130
g16939 and n17127_not n17130 ; n17131
g16940 and asqrt[12] n17109_not ; n17132
g16941 and n17104_not n17132 ; n17133
g16942 and n17100_not n17133 ; n17134
g16943 and n17098_not n17134 ; n17135
g16944 nor n17125 n17135 ; n17136
g16945 and a[24] n17136_not ; n17137
g16946 nor a[24] n17135 ; n17138
g16947 and n17125_not n17138 ; n17139
g16948 nor n17137 n17139 ; n17140
g16949 nor n17131 n17140 ; n17141
g16950 nor n17129 n17141 ; n17142
g16951 and asqrt[14] n17142_not ; n17143
g16952 nor n16485 n16490 ; n17144
g16953 and n16494_not n17144 ; n17145
g16954 and asqrt[11] n17145 ; n17146
g16955 and asqrt[11] n17144 ; n17147
g16956 and n16494 n17147_not ; n17148
g16957 nor n17146 n17148 ; n17149
g16958 nor asqrt[14] n17129 ; n17150
g16959 and n17141_not n17150 ; n17151
g16960 nor n17149 n17151 ; n17152
g16961 nor n17143 n17152 ; n17153
g16962 and asqrt[15] n17153_not ; n17154
g16963 and n16499_not n16508 ; n17155
g16964 and n16497_not n17155 ; n17156
g16965 and asqrt[11] n17156 ; n17157
g16966 nor n16497 n16499 ; n17158
g16967 and asqrt[11] n17158 ; n17159
g16968 nor n16508 n17159 ; n17160
g16969 nor n17157 n17160 ; n17161
g16970 nor asqrt[15] n17143 ; n17162
g16971 and n17152_not n17162 ; n17163
g16972 nor n17161 n17163 ; n17164
g16973 nor n17154 n17164 ; n17165
g16974 and asqrt[16] n17165_not ; n17166
g16975 and n16511_not n16517 ; n17167
g16976 and n16519_not n17167 ; n17168
g16977 and asqrt[11] n17168 ; n17169
g16978 nor n16511 n16519 ; n17170
g16979 and asqrt[11] n17170 ; n17171
g16980 nor n16517 n17171 ; n17172
g16981 nor n17169 n17172 ; n17173
g16982 nor asqrt[16] n17154 ; n17174
g16983 and n17164_not n17174 ; n17175
g16984 nor n17173 n17175 ; n17176
g16985 nor n17166 n17176 ; n17177
g16986 and asqrt[17] n17177_not ; n17178
g16987 and n16529 n16531_not ; n17179
g16988 and n16522_not n17179 ; n17180
g16989 and asqrt[11] n17180 ; n17181
g16990 nor n16522 n16531 ; n17182
g16991 and asqrt[11] n17182 ; n17183
g16992 nor n16529 n17183 ; n17184
g16993 nor n17181 n17184 ; n17185
g16994 nor asqrt[17] n17166 ; n17186
g16995 and n17176_not n17186 ; n17187
g16996 nor n17185 n17187 ; n17188
g16997 nor n17178 n17188 ; n17189
g16998 and asqrt[18] n17189_not ; n17190
g16999 and n16534_not n16541 ; n17191
g17000 and n16543_not n17191 ; n17192
g17001 and asqrt[11] n17192 ; n17193
g17002 nor n16534 n16543 ; n17194
g17003 and asqrt[11] n17194 ; n17195
g17004 nor n16541 n17195 ; n17196
g17005 nor n17193 n17196 ; n17197
g17006 nor asqrt[18] n17178 ; n17198
g17007 and n17188_not n17198 ; n17199
g17008 nor n17197 n17199 ; n17200
g17009 nor n17190 n17200 ; n17201
g17010 and asqrt[19] n17201_not ; n17202
g17011 and n16553 n16555_not ; n17203
g17012 and n16546_not n17203 ; n17204
g17013 and asqrt[11] n17204 ; n17205
g17014 nor n16546 n16555 ; n17206
g17015 and asqrt[11] n17206 ; n17207
g17016 nor n16553 n17207 ; n17208
g17017 nor n17205 n17208 ; n17209
g17018 nor asqrt[19] n17190 ; n17210
g17019 and n17200_not n17210 ; n17211
g17020 nor n17209 n17211 ; n17212
g17021 nor n17202 n17212 ; n17213
g17022 and asqrt[20] n17213_not ; n17214
g17023 and n16558_not n16565 ; n17215
g17024 and n16567_not n17215 ; n17216
g17025 and asqrt[11] n17216 ; n17217
g17026 nor n16558 n16567 ; n17218
g17027 and asqrt[11] n17218 ; n17219
g17028 nor n16565 n17219 ; n17220
g17029 nor n17217 n17220 ; n17221
g17030 nor asqrt[20] n17202 ; n17222
g17031 and n17212_not n17222 ; n17223
g17032 nor n17221 n17223 ; n17224
g17033 nor n17214 n17224 ; n17225
g17034 and asqrt[21] n17225_not ; n17226
g17035 and n16577 n16579_not ; n17227
g17036 and n16570_not n17227 ; n17228
g17037 and asqrt[11] n17228 ; n17229
g17038 nor n16570 n16579 ; n17230
g17039 and asqrt[11] n17230 ; n17231
g17040 nor n16577 n17231 ; n17232
g17041 nor n17229 n17232 ; n17233
g17042 nor asqrt[21] n17214 ; n17234
g17043 and n17224_not n17234 ; n17235
g17044 nor n17233 n17235 ; n17236
g17045 nor n17226 n17236 ; n17237
g17046 and asqrt[22] n17237_not ; n17238
g17047 and n16582_not n16589 ; n17239
g17048 and n16591_not n17239 ; n17240
g17049 and asqrt[11] n17240 ; n17241
g17050 nor n16582 n16591 ; n17242
g17051 and asqrt[11] n17242 ; n17243
g17052 nor n16589 n17243 ; n17244
g17053 nor n17241 n17244 ; n17245
g17054 nor asqrt[22] n17226 ; n17246
g17055 and n17236_not n17246 ; n17247
g17056 nor n17245 n17247 ; n17248
g17057 nor n17238 n17248 ; n17249
g17058 and asqrt[23] n17249_not ; n17250
g17059 and n16601 n16603_not ; n17251
g17060 and n16594_not n17251 ; n17252
g17061 and asqrt[11] n17252 ; n17253
g17062 nor n16594 n16603 ; n17254
g17063 and asqrt[11] n17254 ; n17255
g17064 nor n16601 n17255 ; n17256
g17065 nor n17253 n17256 ; n17257
g17066 nor asqrt[23] n17238 ; n17258
g17067 and n17248_not n17258 ; n17259
g17068 nor n17257 n17259 ; n17260
g17069 nor n17250 n17260 ; n17261
g17070 and asqrt[24] n17261_not ; n17262
g17071 and n16606_not n16613 ; n17263
g17072 and n16615_not n17263 ; n17264
g17073 and asqrt[11] n17264 ; n17265
g17074 nor n16606 n16615 ; n17266
g17075 and asqrt[11] n17266 ; n17267
g17076 nor n16613 n17267 ; n17268
g17077 nor n17265 n17268 ; n17269
g17078 nor asqrt[24] n17250 ; n17270
g17079 and n17260_not n17270 ; n17271
g17080 nor n17269 n17271 ; n17272
g17081 nor n17262 n17272 ; n17273
g17082 and asqrt[25] n17273_not ; n17274
g17083 and n16625 n16627_not ; n17275
g17084 and n16618_not n17275 ; n17276
g17085 and asqrt[11] n17276 ; n17277
g17086 nor n16618 n16627 ; n17278
g17087 and asqrt[11] n17278 ; n17279
g17088 nor n16625 n17279 ; n17280
g17089 nor n17277 n17280 ; n17281
g17090 nor asqrt[25] n17262 ; n17282
g17091 and n17272_not n17282 ; n17283
g17092 nor n17281 n17283 ; n17284
g17093 nor n17274 n17284 ; n17285
g17094 and asqrt[26] n17285_not ; n17286
g17095 and n16630_not n16637 ; n17287
g17096 and n16639_not n17287 ; n17288
g17097 and asqrt[11] n17288 ; n17289
g17098 nor n16630 n16639 ; n17290
g17099 and asqrt[11] n17290 ; n17291
g17100 nor n16637 n17291 ; n17292
g17101 nor n17289 n17292 ; n17293
g17102 nor asqrt[26] n17274 ; n17294
g17103 and n17284_not n17294 ; n17295
g17104 nor n17293 n17295 ; n17296
g17105 nor n17286 n17296 ; n17297
g17106 and asqrt[27] n17297_not ; n17298
g17107 and n16649 n16651_not ; n17299
g17108 and n16642_not n17299 ; n17300
g17109 and asqrt[11] n17300 ; n17301
g17110 nor n16642 n16651 ; n17302
g17111 and asqrt[11] n17302 ; n17303
g17112 nor n16649 n17303 ; n17304
g17113 nor n17301 n17304 ; n17305
g17114 nor asqrt[27] n17286 ; n17306
g17115 and n17296_not n17306 ; n17307
g17116 nor n17305 n17307 ; n17308
g17117 nor n17298 n17308 ; n17309
g17118 and asqrt[28] n17309_not ; n17310
g17119 and n16654_not n16661 ; n17311
g17120 and n16663_not n17311 ; n17312
g17121 and asqrt[11] n17312 ; n17313
g17122 nor n16654 n16663 ; n17314
g17123 and asqrt[11] n17314 ; n17315
g17124 nor n16661 n17315 ; n17316
g17125 nor n17313 n17316 ; n17317
g17126 nor asqrt[28] n17298 ; n17318
g17127 and n17308_not n17318 ; n17319
g17128 nor n17317 n17319 ; n17320
g17129 nor n17310 n17320 ; n17321
g17130 and asqrt[29] n17321_not ; n17322
g17131 and n16673 n16675_not ; n17323
g17132 and n16666_not n17323 ; n17324
g17133 and asqrt[11] n17324 ; n17325
g17134 nor n16666 n16675 ; n17326
g17135 and asqrt[11] n17326 ; n17327
g17136 nor n16673 n17327 ; n17328
g17137 nor n17325 n17328 ; n17329
g17138 nor asqrt[29] n17310 ; n17330
g17139 and n17320_not n17330 ; n17331
g17140 nor n17329 n17331 ; n17332
g17141 nor n17322 n17332 ; n17333
g17142 and asqrt[30] n17333_not ; n17334
g17143 and n16678_not n16685 ; n17335
g17144 and n16687_not n17335 ; n17336
g17145 and asqrt[11] n17336 ; n17337
g17146 nor n16678 n16687 ; n17338
g17147 and asqrt[11] n17338 ; n17339
g17148 nor n16685 n17339 ; n17340
g17149 nor n17337 n17340 ; n17341
g17150 nor asqrt[30] n17322 ; n17342
g17151 and n17332_not n17342 ; n17343
g17152 nor n17341 n17343 ; n17344
g17153 nor n17334 n17344 ; n17345
g17154 and asqrt[31] n17345_not ; n17346
g17155 and n16697 n16699_not ; n17347
g17156 and n16690_not n17347 ; n17348
g17157 and asqrt[11] n17348 ; n17349
g17158 nor n16690 n16699 ; n17350
g17159 and asqrt[11] n17350 ; n17351
g17160 nor n16697 n17351 ; n17352
g17161 nor n17349 n17352 ; n17353
g17162 nor asqrt[31] n17334 ; n17354
g17163 and n17344_not n17354 ; n17355
g17164 nor n17353 n17355 ; n17356
g17165 nor n17346 n17356 ; n17357
g17166 and asqrt[32] n17357_not ; n17358
g17167 and n16702_not n16709 ; n17359
g17168 and n16711_not n17359 ; n17360
g17169 and asqrt[11] n17360 ; n17361
g17170 nor n16702 n16711 ; n17362
g17171 and asqrt[11] n17362 ; n17363
g17172 nor n16709 n17363 ; n17364
g17173 nor n17361 n17364 ; n17365
g17174 nor asqrt[32] n17346 ; n17366
g17175 and n17356_not n17366 ; n17367
g17176 nor n17365 n17367 ; n17368
g17177 nor n17358 n17368 ; n17369
g17178 and asqrt[33] n17369_not ; n17370
g17179 and n16721 n16723_not ; n17371
g17180 and n16714_not n17371 ; n17372
g17181 and asqrt[11] n17372 ; n17373
g17182 nor n16714 n16723 ; n17374
g17183 and asqrt[11] n17374 ; n17375
g17184 nor n16721 n17375 ; n17376
g17185 nor n17373 n17376 ; n17377
g17186 nor asqrt[33] n17358 ; n17378
g17187 and n17368_not n17378 ; n17379
g17188 nor n17377 n17379 ; n17380
g17189 nor n17370 n17380 ; n17381
g17190 and asqrt[34] n17381_not ; n17382
g17191 and n16726_not n16733 ; n17383
g17192 and n16735_not n17383 ; n17384
g17193 and asqrt[11] n17384 ; n17385
g17194 nor n16726 n16735 ; n17386
g17195 and asqrt[11] n17386 ; n17387
g17196 nor n16733 n17387 ; n17388
g17197 nor n17385 n17388 ; n17389
g17198 nor asqrt[34] n17370 ; n17390
g17199 and n17380_not n17390 ; n17391
g17200 nor n17389 n17391 ; n17392
g17201 nor n17382 n17392 ; n17393
g17202 and asqrt[35] n17393_not ; n17394
g17203 and n16745 n16747_not ; n17395
g17204 and n16738_not n17395 ; n17396
g17205 and asqrt[11] n17396 ; n17397
g17206 nor n16738 n16747 ; n17398
g17207 and asqrt[11] n17398 ; n17399
g17208 nor n16745 n17399 ; n17400
g17209 nor n17397 n17400 ; n17401
g17210 nor asqrt[35] n17382 ; n17402
g17211 and n17392_not n17402 ; n17403
g17212 nor n17401 n17403 ; n17404
g17213 nor n17394 n17404 ; n17405
g17214 and asqrt[36] n17405_not ; n17406
g17215 and n16750_not n16757 ; n17407
g17216 and n16759_not n17407 ; n17408
g17217 and asqrt[11] n17408 ; n17409
g17218 nor n16750 n16759 ; n17410
g17219 and asqrt[11] n17410 ; n17411
g17220 nor n16757 n17411 ; n17412
g17221 nor n17409 n17412 ; n17413
g17222 nor asqrt[36] n17394 ; n17414
g17223 and n17404_not n17414 ; n17415
g17224 nor n17413 n17415 ; n17416
g17225 nor n17406 n17416 ; n17417
g17226 and asqrt[37] n17417_not ; n17418
g17227 and n16769 n16771_not ; n17419
g17228 and n16762_not n17419 ; n17420
g17229 and asqrt[11] n17420 ; n17421
g17230 nor n16762 n16771 ; n17422
g17231 and asqrt[11] n17422 ; n17423
g17232 nor n16769 n17423 ; n17424
g17233 nor n17421 n17424 ; n17425
g17234 nor asqrt[37] n17406 ; n17426
g17235 and n17416_not n17426 ; n17427
g17236 nor n17425 n17427 ; n17428
g17237 nor n17418 n17428 ; n17429
g17238 and asqrt[38] n17429_not ; n17430
g17239 and n16774_not n16781 ; n17431
g17240 and n16783_not n17431 ; n17432
g17241 and asqrt[11] n17432 ; n17433
g17242 nor n16774 n16783 ; n17434
g17243 and asqrt[11] n17434 ; n17435
g17244 nor n16781 n17435 ; n17436
g17245 nor n17433 n17436 ; n17437
g17246 nor asqrt[38] n17418 ; n17438
g17247 and n17428_not n17438 ; n17439
g17248 nor n17437 n17439 ; n17440
g17249 nor n17430 n17440 ; n17441
g17250 and asqrt[39] n17441_not ; n17442
g17251 and n16793 n16795_not ; n17443
g17252 and n16786_not n17443 ; n17444
g17253 and asqrt[11] n17444 ; n17445
g17254 nor n16786 n16795 ; n17446
g17255 and asqrt[11] n17446 ; n17447
g17256 nor n16793 n17447 ; n17448
g17257 nor n17445 n17448 ; n17449
g17258 nor asqrt[39] n17430 ; n17450
g17259 and n17440_not n17450 ; n17451
g17260 nor n17449 n17451 ; n17452
g17261 nor n17442 n17452 ; n17453
g17262 and asqrt[40] n17453_not ; n17454
g17263 and n16798_not n16805 ; n17455
g17264 and n16807_not n17455 ; n17456
g17265 and asqrt[11] n17456 ; n17457
g17266 nor n16798 n16807 ; n17458
g17267 and asqrt[11] n17458 ; n17459
g17268 nor n16805 n17459 ; n17460
g17269 nor n17457 n17460 ; n17461
g17270 nor asqrt[40] n17442 ; n17462
g17271 and n17452_not n17462 ; n17463
g17272 nor n17461 n17463 ; n17464
g17273 nor n17454 n17464 ; n17465
g17274 and asqrt[41] n17465_not ; n17466
g17275 and n16817 n16819_not ; n17467
g17276 and n16810_not n17467 ; n17468
g17277 and asqrt[11] n17468 ; n17469
g17278 nor n16810 n16819 ; n17470
g17279 and asqrt[11] n17470 ; n17471
g17280 nor n16817 n17471 ; n17472
g17281 nor n17469 n17472 ; n17473
g17282 nor asqrt[41] n17454 ; n17474
g17283 and n17464_not n17474 ; n17475
g17284 nor n17473 n17475 ; n17476
g17285 nor n17466 n17476 ; n17477
g17286 and asqrt[42] n17477_not ; n17478
g17287 and n16822_not n16829 ; n17479
g17288 and n16831_not n17479 ; n17480
g17289 and asqrt[11] n17480 ; n17481
g17290 nor n16822 n16831 ; n17482
g17291 and asqrt[11] n17482 ; n17483
g17292 nor n16829 n17483 ; n17484
g17293 nor n17481 n17484 ; n17485
g17294 nor asqrt[42] n17466 ; n17486
g17295 and n17476_not n17486 ; n17487
g17296 nor n17485 n17487 ; n17488
g17297 nor n17478 n17488 ; n17489
g17298 and asqrt[43] n17489_not ; n17490
g17299 and n16841 n16843_not ; n17491
g17300 and n16834_not n17491 ; n17492
g17301 and asqrt[11] n17492 ; n17493
g17302 nor n16834 n16843 ; n17494
g17303 and asqrt[11] n17494 ; n17495
g17304 nor n16841 n17495 ; n17496
g17305 nor n17493 n17496 ; n17497
g17306 nor asqrt[43] n17478 ; n17498
g17307 and n17488_not n17498 ; n17499
g17308 nor n17497 n17499 ; n17500
g17309 nor n17490 n17500 ; n17501
g17310 and asqrt[44] n17501_not ; n17502
g17311 and n16846_not n16853 ; n17503
g17312 and n16855_not n17503 ; n17504
g17313 and asqrt[11] n17504 ; n17505
g17314 nor n16846 n16855 ; n17506
g17315 and asqrt[11] n17506 ; n17507
g17316 nor n16853 n17507 ; n17508
g17317 nor n17505 n17508 ; n17509
g17318 nor asqrt[44] n17490 ; n17510
g17319 and n17500_not n17510 ; n17511
g17320 nor n17509 n17511 ; n17512
g17321 nor n17502 n17512 ; n17513
g17322 and asqrt[45] n17513_not ; n17514
g17323 and n16865 n16867_not ; n17515
g17324 and n16858_not n17515 ; n17516
g17325 and asqrt[11] n17516 ; n17517
g17326 nor n16858 n16867 ; n17518
g17327 and asqrt[11] n17518 ; n17519
g17328 nor n16865 n17519 ; n17520
g17329 nor n17517 n17520 ; n17521
g17330 nor asqrt[45] n17502 ; n17522
g17331 and n17512_not n17522 ; n17523
g17332 nor n17521 n17523 ; n17524
g17333 nor n17514 n17524 ; n17525
g17334 and asqrt[46] n17525_not ; n17526
g17335 and n16870_not n16877 ; n17527
g17336 and n16879_not n17527 ; n17528
g17337 and asqrt[11] n17528 ; n17529
g17338 nor n16870 n16879 ; n17530
g17339 and asqrt[11] n17530 ; n17531
g17340 nor n16877 n17531 ; n17532
g17341 nor n17529 n17532 ; n17533
g17342 nor asqrt[46] n17514 ; n17534
g17343 and n17524_not n17534 ; n17535
g17344 nor n17533 n17535 ; n17536
g17345 nor n17526 n17536 ; n17537
g17346 and asqrt[47] n17537_not ; n17538
g17347 and n16889 n16891_not ; n17539
g17348 and n16882_not n17539 ; n17540
g17349 and asqrt[11] n17540 ; n17541
g17350 nor n16882 n16891 ; n17542
g17351 and asqrt[11] n17542 ; n17543
g17352 nor n16889 n17543 ; n17544
g17353 nor n17541 n17544 ; n17545
g17354 nor asqrt[47] n17526 ; n17546
g17355 and n17536_not n17546 ; n17547
g17356 nor n17545 n17547 ; n17548
g17357 nor n17538 n17548 ; n17549
g17358 and asqrt[48] n17549_not ; n17550
g17359 and n16894_not n16901 ; n17551
g17360 and n16903_not n17551 ; n17552
g17361 and asqrt[11] n17552 ; n17553
g17362 nor n16894 n16903 ; n17554
g17363 and asqrt[11] n17554 ; n17555
g17364 nor n16901 n17555 ; n17556
g17365 nor n17553 n17556 ; n17557
g17366 nor asqrt[48] n17538 ; n17558
g17367 and n17548_not n17558 ; n17559
g17368 nor n17557 n17559 ; n17560
g17369 nor n17550 n17560 ; n17561
g17370 and asqrt[49] n17561_not ; n17562
g17371 and n16913 n16915_not ; n17563
g17372 and n16906_not n17563 ; n17564
g17373 and asqrt[11] n17564 ; n17565
g17374 nor n16906 n16915 ; n17566
g17375 and asqrt[11] n17566 ; n17567
g17376 nor n16913 n17567 ; n17568
g17377 nor n17565 n17568 ; n17569
g17378 nor asqrt[49] n17550 ; n17570
g17379 and n17560_not n17570 ; n17571
g17380 nor n17569 n17571 ; n17572
g17381 nor n17562 n17572 ; n17573
g17382 and asqrt[50] n17573_not ; n17574
g17383 and n16918_not n16925 ; n17575
g17384 and n16927_not n17575 ; n17576
g17385 and asqrt[11] n17576 ; n17577
g17386 nor n16918 n16927 ; n17578
g17387 and asqrt[11] n17578 ; n17579
g17388 nor n16925 n17579 ; n17580
g17389 nor n17577 n17580 ; n17581
g17390 nor asqrt[50] n17562 ; n17582
g17391 and n17572_not n17582 ; n17583
g17392 nor n17581 n17583 ; n17584
g17393 nor n17574 n17584 ; n17585
g17394 and asqrt[51] n17585_not ; n17586
g17395 and n16937 n16939_not ; n17587
g17396 and n16930_not n17587 ; n17588
g17397 and asqrt[11] n17588 ; n17589
g17398 nor n16930 n16939 ; n17590
g17399 and asqrt[11] n17590 ; n17591
g17400 nor n16937 n17591 ; n17592
g17401 nor n17589 n17592 ; n17593
g17402 nor asqrt[51] n17574 ; n17594
g17403 and n17584_not n17594 ; n17595
g17404 nor n17593 n17595 ; n17596
g17405 nor n17586 n17596 ; n17597
g17406 and asqrt[52] n17597_not ; n17598
g17407 and n16942_not n16949 ; n17599
g17408 and n16951_not n17599 ; n17600
g17409 and asqrt[11] n17600 ; n17601
g17410 nor n16942 n16951 ; n17602
g17411 and asqrt[11] n17602 ; n17603
g17412 nor n16949 n17603 ; n17604
g17413 nor n17601 n17604 ; n17605
g17414 nor asqrt[52] n17586 ; n17606
g17415 and n17596_not n17606 ; n17607
g17416 nor n17605 n17607 ; n17608
g17417 nor n17598 n17608 ; n17609
g17418 and asqrt[53] n17609_not ; n17610
g17419 and n16961 n16963_not ; n17611
g17420 and n16954_not n17611 ; n17612
g17421 and asqrt[11] n17612 ; n17613
g17422 nor n16954 n16963 ; n17614
g17423 and asqrt[11] n17614 ; n17615
g17424 nor n16961 n17615 ; n17616
g17425 nor n17613 n17616 ; n17617
g17426 nor asqrt[53] n17598 ; n17618
g17427 and n17608_not n17618 ; n17619
g17428 nor n17617 n17619 ; n17620
g17429 nor n17610 n17620 ; n17621
g17430 and asqrt[54] n17621_not ; n17622
g17431 nor asqrt[54] n17610 ; n17623
g17432 and n17620_not n17623 ; n17624
g17433 and n16966_not n16975 ; n17625
g17434 and n16968_not n17625 ; n17626
g17435 and asqrt[11] n17626 ; n17627
g17436 nor n16966 n16968 ; n17628
g17437 and asqrt[11] n17628 ; n17629
g17438 nor n16975 n17629 ; n17630
g17439 nor n17627 n17630 ; n17631
g17440 nor n17624 n17631 ; n17632
g17441 nor n17622 n17632 ; n17633
g17442 and asqrt[55] n17633_not ; n17634
g17443 and n16985 n16987_not ; n17635
g17444 and n16978_not n17635 ; n17636
g17445 and asqrt[11] n17636 ; n17637
g17446 nor n16978 n16987 ; n17638
g17447 and asqrt[11] n17638 ; n17639
g17448 nor n16985 n17639 ; n17640
g17449 nor n17637 n17640 ; n17641
g17450 nor asqrt[55] n17622 ; n17642
g17451 and n17632_not n17642 ; n17643
g17452 nor n17641 n17643 ; n17644
g17453 nor n17634 n17644 ; n17645
g17454 and asqrt[56] n17645_not ; n17646
g17455 and n16990_not n16997 ; n17647
g17456 and n16999_not n17647 ; n17648
g17457 and asqrt[11] n17648 ; n17649
g17458 nor n16990 n16999 ; n17650
g17459 and asqrt[11] n17650 ; n17651
g17460 nor n16997 n17651 ; n17652
g17461 nor n17649 n17652 ; n17653
g17462 nor asqrt[56] n17634 ; n17654
g17463 and n17644_not n17654 ; n17655
g17464 nor n17653 n17655 ; n17656
g17465 nor n17646 n17656 ; n17657
g17466 and asqrt[57] n17657_not ; n17658
g17467 and n17009 n17011_not ; n17659
g17468 and n17002_not n17659 ; n17660
g17469 and asqrt[11] n17660 ; n17661
g17470 nor n17002 n17011 ; n17662
g17471 and asqrt[11] n17662 ; n17663
g17472 nor n17009 n17663 ; n17664
g17473 nor n17661 n17664 ; n17665
g17474 nor asqrt[57] n17646 ; n17666
g17475 and n17656_not n17666 ; n17667
g17476 nor n17665 n17667 ; n17668
g17477 nor n17658 n17668 ; n17669
g17478 and asqrt[58] n17669_not ; n17670
g17479 and n17014_not n17021 ; n17671
g17480 and n17023_not n17671 ; n17672
g17481 and asqrt[11] n17672 ; n17673
g17482 nor n17014 n17023 ; n17674
g17483 and asqrt[11] n17674 ; n17675
g17484 nor n17021 n17675 ; n17676
g17485 nor n17673 n17676 ; n17677
g17486 nor asqrt[58] n17658 ; n17678
g17487 and n17668_not n17678 ; n17679
g17488 nor n17677 n17679 ; n17680
g17489 nor n17670 n17680 ; n17681
g17490 and asqrt[59] n17681_not ; n17682
g17491 and n17033 n17035_not ; n17683
g17492 and n17026_not n17683 ; n17684
g17493 and asqrt[11] n17684 ; n17685
g17494 nor n17026 n17035 ; n17686
g17495 and asqrt[11] n17686 ; n17687
g17496 nor n17033 n17687 ; n17688
g17497 nor n17685 n17688 ; n17689
g17498 nor asqrt[59] n17670 ; n17690
g17499 and n17680_not n17690 ; n17691
g17500 nor n17689 n17691 ; n17692
g17501 nor n17682 n17692 ; n17693
g17502 and asqrt[60] n17693_not ; n17694
g17503 and n17038_not n17045 ; n17695
g17504 and n17047_not n17695 ; n17696
g17505 and asqrt[11] n17696 ; n17697
g17506 nor n17038 n17047 ; n17698
g17507 and asqrt[11] n17698 ; n17699
g17508 nor n17045 n17699 ; n17700
g17509 nor n17697 n17700 ; n17701
g17510 nor asqrt[60] n17682 ; n17702
g17511 and n17692_not n17702 ; n17703
g17512 nor n17701 n17703 ; n17704
g17513 nor n17694 n17704 ; n17705
g17514 and asqrt[61] n17705_not ; n17706
g17515 and n17057 n17059_not ; n17707
g17516 and n17050_not n17707 ; n17708
g17517 and asqrt[11] n17708 ; n17709
g17518 nor n17050 n17059 ; n17710
g17519 and asqrt[11] n17710 ; n17711
g17520 nor n17057 n17711 ; n17712
g17521 nor n17709 n17712 ; n17713
g17522 nor asqrt[61] n17694 ; n17714
g17523 and n17704_not n17714 ; n17715
g17524 nor n17713 n17715 ; n17716
g17525 nor n17706 n17716 ; n17717
g17526 and asqrt[62] n17717_not ; n17718
g17527 and n17062_not n17069 ; n17719
g17528 and n17071_not n17719 ; n17720
g17529 and asqrt[11] n17720 ; n17721
g17530 nor n17062 n17071 ; n17722
g17531 and asqrt[11] n17722 ; n17723
g17532 nor n17069 n17723 ; n17724
g17533 nor n17721 n17724 ; n17725
g17534 nor asqrt[62] n17706 ; n17726
g17535 and n17716_not n17726 ; n17727
g17536 nor n17725 n17727 ; n17728
g17537 nor n17718 n17728 ; n17729
g17538 and n17081 n17083_not ; n17730
g17539 and n17074_not n17730 ; n17731
g17540 and asqrt[11] n17731 ; n17732
g17541 nor n17074 n17083 ; n17733
g17542 and asqrt[11] n17733 ; n17734
g17543 nor n17081 n17734 ; n17735
g17544 nor n17732 n17735 ; n17736
g17545 nor n17085 n17092 ; n17737
g17546 and asqrt[11] n17737 ; n17738
g17547 nor n17100 n17738 ; n17739
g17548 and n17736_not n17739 ; n17740
g17549 and n17729_not n17740 ; n17741
g17550 nor asqrt[63] n17741 ; n17742
g17551 and n17718_not n17736 ; n17743
g17552 and n17728_not n17743 ; n17744
g17553 and n17092_not asqrt[11] ; n17745
g17554 and n17085 n17745_not ; n17746
g17555 and asqrt[63] n17737_not ; n17747
g17556 and n17746_not n17747 ; n17748
g17557 nor n17088 n17109 ; n17749
g17558 and n17091_not n17749 ; n17750
g17559 and n17104_not n17750 ; n17751
g17560 and n17100_not n17751 ; n17752
g17561 and n17098_not n17752 ; n17753
g17562 nor n17748 n17753 ; n17754
g17563 and n17744_not n17754 ; n17755
g17564 nand n17742_not n17755 ; asqrt[10]
g17565 and a[20] asqrt[10] ; n17757
g17566 nor a[18] a[19] ; n17758
g17567 and a[20]_not n17758 ; n17759
g17568 nor n17757 n17759 ; n17760
g17569 and asqrt[11] n17760_not ; n17761
g17570 nor n17109 n17759 ; n17762
g17571 and n17104_not n17762 ; n17763
g17572 and n17100_not n17763 ; n17764
g17573 and n17098_not n17764 ; n17765
g17574 and n17757_not n17765 ; n17766
g17575 and a[20]_not asqrt[10] ; n17767
g17576 and a[21] n17767_not ; n17768
g17577 and n17114 asqrt[10] ; n17769
g17578 nor n17768 n17769 ; n17770
g17579 and n17766_not n17770 ; n17771
g17580 nor n17761 n17771 ; n17772
g17581 and asqrt[12] n17772_not ; n17773
g17582 nor asqrt[12] n17761 ; n17774
g17583 and n17771_not n17774 ; n17775
g17584 and asqrt[11] n17753_not ; n17776
g17585 and n17748_not n17776 ; n17777
g17586 and n17744_not n17777 ; n17778
g17587 and n17742_not n17778 ; n17779
g17588 nor n17769 n17779 ; n17780
g17589 and a[22] n17780_not ; n17781
g17590 nor a[22] n17779 ; n17782
g17591 and n17769_not n17782 ; n17783
g17592 nor n17781 n17783 ; n17784
g17593 nor n17775 n17784 ; n17785
g17594 nor n17773 n17785 ; n17786
g17595 and asqrt[13] n17786_not ; n17787
g17596 nor n17117 n17122 ; n17788
g17597 and n17126_not n17788 ; n17789
g17598 and asqrt[10] n17789 ; n17790
g17599 and asqrt[10] n17788 ; n17791
g17600 and n17126 n17791_not ; n17792
g17601 nor n17790 n17792 ; n17793
g17602 nor asqrt[13] n17773 ; n17794
g17603 and n17785_not n17794 ; n17795
g17604 nor n17793 n17795 ; n17796
g17605 nor n17787 n17796 ; n17797
g17606 and asqrt[14] n17797_not ; n17798
g17607 and n17131_not n17140 ; n17799
g17608 and n17129_not n17799 ; n17800
g17609 and asqrt[10] n17800 ; n17801
g17610 nor n17129 n17131 ; n17802
g17611 and asqrt[10] n17802 ; n17803
g17612 nor n17140 n17803 ; n17804
g17613 nor n17801 n17804 ; n17805
g17614 nor asqrt[14] n17787 ; n17806
g17615 and n17796_not n17806 ; n17807
g17616 nor n17805 n17807 ; n17808
g17617 nor n17798 n17808 ; n17809
g17618 and asqrt[15] n17809_not ; n17810
g17619 and n17143_not n17149 ; n17811
g17620 and n17151_not n17811 ; n17812
g17621 and asqrt[10] n17812 ; n17813
g17622 nor n17143 n17151 ; n17814
g17623 and asqrt[10] n17814 ; n17815
g17624 nor n17149 n17815 ; n17816
g17625 nor n17813 n17816 ; n17817
g17626 nor asqrt[15] n17798 ; n17818
g17627 and n17808_not n17818 ; n17819
g17628 nor n17817 n17819 ; n17820
g17629 nor n17810 n17820 ; n17821
g17630 and asqrt[16] n17821_not ; n17822
g17631 and n17161 n17163_not ; n17823
g17632 and n17154_not n17823 ; n17824
g17633 and asqrt[10] n17824 ; n17825
g17634 nor n17154 n17163 ; n17826
g17635 and asqrt[10] n17826 ; n17827
g17636 nor n17161 n17827 ; n17828
g17637 nor n17825 n17828 ; n17829
g17638 nor asqrt[16] n17810 ; n17830
g17639 and n17820_not n17830 ; n17831
g17640 nor n17829 n17831 ; n17832
g17641 nor n17822 n17832 ; n17833
g17642 and asqrt[17] n17833_not ; n17834
g17643 and n17166_not n17173 ; n17835
g17644 and n17175_not n17835 ; n17836
g17645 and asqrt[10] n17836 ; n17837
g17646 nor n17166 n17175 ; n17838
g17647 and asqrt[10] n17838 ; n17839
g17648 nor n17173 n17839 ; n17840
g17649 nor n17837 n17840 ; n17841
g17650 nor asqrt[17] n17822 ; n17842
g17651 and n17832_not n17842 ; n17843
g17652 nor n17841 n17843 ; n17844
g17653 nor n17834 n17844 ; n17845
g17654 and asqrt[18] n17845_not ; n17846
g17655 and n17185 n17187_not ; n17847
g17656 and n17178_not n17847 ; n17848
g17657 and asqrt[10] n17848 ; n17849
g17658 nor n17178 n17187 ; n17850
g17659 and asqrt[10] n17850 ; n17851
g17660 nor n17185 n17851 ; n17852
g17661 nor n17849 n17852 ; n17853
g17662 nor asqrt[18] n17834 ; n17854
g17663 and n17844_not n17854 ; n17855
g17664 nor n17853 n17855 ; n17856
g17665 nor n17846 n17856 ; n17857
g17666 and asqrt[19] n17857_not ; n17858
g17667 and n17190_not n17197 ; n17859
g17668 and n17199_not n17859 ; n17860
g17669 and asqrt[10] n17860 ; n17861
g17670 nor n17190 n17199 ; n17862
g17671 and asqrt[10] n17862 ; n17863
g17672 nor n17197 n17863 ; n17864
g17673 nor n17861 n17864 ; n17865
g17674 nor asqrt[19] n17846 ; n17866
g17675 and n17856_not n17866 ; n17867
g17676 nor n17865 n17867 ; n17868
g17677 nor n17858 n17868 ; n17869
g17678 and asqrt[20] n17869_not ; n17870
g17679 and n17209 n17211_not ; n17871
g17680 and n17202_not n17871 ; n17872
g17681 and asqrt[10] n17872 ; n17873
g17682 nor n17202 n17211 ; n17874
g17683 and asqrt[10] n17874 ; n17875
g17684 nor n17209 n17875 ; n17876
g17685 nor n17873 n17876 ; n17877
g17686 nor asqrt[20] n17858 ; n17878
g17687 and n17868_not n17878 ; n17879
g17688 nor n17877 n17879 ; n17880
g17689 nor n17870 n17880 ; n17881
g17690 and asqrt[21] n17881_not ; n17882
g17691 and n17214_not n17221 ; n17883
g17692 and n17223_not n17883 ; n17884
g17693 and asqrt[10] n17884 ; n17885
g17694 nor n17214 n17223 ; n17886
g17695 and asqrt[10] n17886 ; n17887
g17696 nor n17221 n17887 ; n17888
g17697 nor n17885 n17888 ; n17889
g17698 nor asqrt[21] n17870 ; n17890
g17699 and n17880_not n17890 ; n17891
g17700 nor n17889 n17891 ; n17892
g17701 nor n17882 n17892 ; n17893
g17702 and asqrt[22] n17893_not ; n17894
g17703 and n17233 n17235_not ; n17895
g17704 and n17226_not n17895 ; n17896
g17705 and asqrt[10] n17896 ; n17897
g17706 nor n17226 n17235 ; n17898
g17707 and asqrt[10] n17898 ; n17899
g17708 nor n17233 n17899 ; n17900
g17709 nor n17897 n17900 ; n17901
g17710 nor asqrt[22] n17882 ; n17902
g17711 and n17892_not n17902 ; n17903
g17712 nor n17901 n17903 ; n17904
g17713 nor n17894 n17904 ; n17905
g17714 and asqrt[23] n17905_not ; n17906
g17715 and n17238_not n17245 ; n17907
g17716 and n17247_not n17907 ; n17908
g17717 and asqrt[10] n17908 ; n17909
g17718 nor n17238 n17247 ; n17910
g17719 and asqrt[10] n17910 ; n17911
g17720 nor n17245 n17911 ; n17912
g17721 nor n17909 n17912 ; n17913
g17722 nor asqrt[23] n17894 ; n17914
g17723 and n17904_not n17914 ; n17915
g17724 nor n17913 n17915 ; n17916
g17725 nor n17906 n17916 ; n17917
g17726 and asqrt[24] n17917_not ; n17918
g17727 and n17257 n17259_not ; n17919
g17728 and n17250_not n17919 ; n17920
g17729 and asqrt[10] n17920 ; n17921
g17730 nor n17250 n17259 ; n17922
g17731 and asqrt[10] n17922 ; n17923
g17732 nor n17257 n17923 ; n17924
g17733 nor n17921 n17924 ; n17925
g17734 nor asqrt[24] n17906 ; n17926
g17735 and n17916_not n17926 ; n17927
g17736 nor n17925 n17927 ; n17928
g17737 nor n17918 n17928 ; n17929
g17738 and asqrt[25] n17929_not ; n17930
g17739 and n17262_not n17269 ; n17931
g17740 and n17271_not n17931 ; n17932
g17741 and asqrt[10] n17932 ; n17933
g17742 nor n17262 n17271 ; n17934
g17743 and asqrt[10] n17934 ; n17935
g17744 nor n17269 n17935 ; n17936
g17745 nor n17933 n17936 ; n17937
g17746 nor asqrt[25] n17918 ; n17938
g17747 and n17928_not n17938 ; n17939
g17748 nor n17937 n17939 ; n17940
g17749 nor n17930 n17940 ; n17941
g17750 and asqrt[26] n17941_not ; n17942
g17751 and n17281 n17283_not ; n17943
g17752 and n17274_not n17943 ; n17944
g17753 and asqrt[10] n17944 ; n17945
g17754 nor n17274 n17283 ; n17946
g17755 and asqrt[10] n17946 ; n17947
g17756 nor n17281 n17947 ; n17948
g17757 nor n17945 n17948 ; n17949
g17758 nor asqrt[26] n17930 ; n17950
g17759 and n17940_not n17950 ; n17951
g17760 nor n17949 n17951 ; n17952
g17761 nor n17942 n17952 ; n17953
g17762 and asqrt[27] n17953_not ; n17954
g17763 and n17286_not n17293 ; n17955
g17764 and n17295_not n17955 ; n17956
g17765 and asqrt[10] n17956 ; n17957
g17766 nor n17286 n17295 ; n17958
g17767 and asqrt[10] n17958 ; n17959
g17768 nor n17293 n17959 ; n17960
g17769 nor n17957 n17960 ; n17961
g17770 nor asqrt[27] n17942 ; n17962
g17771 and n17952_not n17962 ; n17963
g17772 nor n17961 n17963 ; n17964
g17773 nor n17954 n17964 ; n17965
g17774 and asqrt[28] n17965_not ; n17966
g17775 and n17305 n17307_not ; n17967
g17776 and n17298_not n17967 ; n17968
g17777 and asqrt[10] n17968 ; n17969
g17778 nor n17298 n17307 ; n17970
g17779 and asqrt[10] n17970 ; n17971
g17780 nor n17305 n17971 ; n17972
g17781 nor n17969 n17972 ; n17973
g17782 nor asqrt[28] n17954 ; n17974
g17783 and n17964_not n17974 ; n17975
g17784 nor n17973 n17975 ; n17976
g17785 nor n17966 n17976 ; n17977
g17786 and asqrt[29] n17977_not ; n17978
g17787 and n17310_not n17317 ; n17979
g17788 and n17319_not n17979 ; n17980
g17789 and asqrt[10] n17980 ; n17981
g17790 nor n17310 n17319 ; n17982
g17791 and asqrt[10] n17982 ; n17983
g17792 nor n17317 n17983 ; n17984
g17793 nor n17981 n17984 ; n17985
g17794 nor asqrt[29] n17966 ; n17986
g17795 and n17976_not n17986 ; n17987
g17796 nor n17985 n17987 ; n17988
g17797 nor n17978 n17988 ; n17989
g17798 and asqrt[30] n17989_not ; n17990
g17799 and n17329 n17331_not ; n17991
g17800 and n17322_not n17991 ; n17992
g17801 and asqrt[10] n17992 ; n17993
g17802 nor n17322 n17331 ; n17994
g17803 and asqrt[10] n17994 ; n17995
g17804 nor n17329 n17995 ; n17996
g17805 nor n17993 n17996 ; n17997
g17806 nor asqrt[30] n17978 ; n17998
g17807 and n17988_not n17998 ; n17999
g17808 nor n17997 n17999 ; n18000
g17809 nor n17990 n18000 ; n18001
g17810 and asqrt[31] n18001_not ; n18002
g17811 and n17334_not n17341 ; n18003
g17812 and n17343_not n18003 ; n18004
g17813 and asqrt[10] n18004 ; n18005
g17814 nor n17334 n17343 ; n18006
g17815 and asqrt[10] n18006 ; n18007
g17816 nor n17341 n18007 ; n18008
g17817 nor n18005 n18008 ; n18009
g17818 nor asqrt[31] n17990 ; n18010
g17819 and n18000_not n18010 ; n18011
g17820 nor n18009 n18011 ; n18012
g17821 nor n18002 n18012 ; n18013
g17822 and asqrt[32] n18013_not ; n18014
g17823 and n17353 n17355_not ; n18015
g17824 and n17346_not n18015 ; n18016
g17825 and asqrt[10] n18016 ; n18017
g17826 nor n17346 n17355 ; n18018
g17827 and asqrt[10] n18018 ; n18019
g17828 nor n17353 n18019 ; n18020
g17829 nor n18017 n18020 ; n18021
g17830 nor asqrt[32] n18002 ; n18022
g17831 and n18012_not n18022 ; n18023
g17832 nor n18021 n18023 ; n18024
g17833 nor n18014 n18024 ; n18025
g17834 and asqrt[33] n18025_not ; n18026
g17835 and n17358_not n17365 ; n18027
g17836 and n17367_not n18027 ; n18028
g17837 and asqrt[10] n18028 ; n18029
g17838 nor n17358 n17367 ; n18030
g17839 and asqrt[10] n18030 ; n18031
g17840 nor n17365 n18031 ; n18032
g17841 nor n18029 n18032 ; n18033
g17842 nor asqrt[33] n18014 ; n18034
g17843 and n18024_not n18034 ; n18035
g17844 nor n18033 n18035 ; n18036
g17845 nor n18026 n18036 ; n18037
g17846 and asqrt[34] n18037_not ; n18038
g17847 and n17377 n17379_not ; n18039
g17848 and n17370_not n18039 ; n18040
g17849 and asqrt[10] n18040 ; n18041
g17850 nor n17370 n17379 ; n18042
g17851 and asqrt[10] n18042 ; n18043
g17852 nor n17377 n18043 ; n18044
g17853 nor n18041 n18044 ; n18045
g17854 nor asqrt[34] n18026 ; n18046
g17855 and n18036_not n18046 ; n18047
g17856 nor n18045 n18047 ; n18048
g17857 nor n18038 n18048 ; n18049
g17858 and asqrt[35] n18049_not ; n18050
g17859 and n17382_not n17389 ; n18051
g17860 and n17391_not n18051 ; n18052
g17861 and asqrt[10] n18052 ; n18053
g17862 nor n17382 n17391 ; n18054
g17863 and asqrt[10] n18054 ; n18055
g17864 nor n17389 n18055 ; n18056
g17865 nor n18053 n18056 ; n18057
g17866 nor asqrt[35] n18038 ; n18058
g17867 and n18048_not n18058 ; n18059
g17868 nor n18057 n18059 ; n18060
g17869 nor n18050 n18060 ; n18061
g17870 and asqrt[36] n18061_not ; n18062
g17871 and n17401 n17403_not ; n18063
g17872 and n17394_not n18063 ; n18064
g17873 and asqrt[10] n18064 ; n18065
g17874 nor n17394 n17403 ; n18066
g17875 and asqrt[10] n18066 ; n18067
g17876 nor n17401 n18067 ; n18068
g17877 nor n18065 n18068 ; n18069
g17878 nor asqrt[36] n18050 ; n18070
g17879 and n18060_not n18070 ; n18071
g17880 nor n18069 n18071 ; n18072
g17881 nor n18062 n18072 ; n18073
g17882 and asqrt[37] n18073_not ; n18074
g17883 and n17406_not n17413 ; n18075
g17884 and n17415_not n18075 ; n18076
g17885 and asqrt[10] n18076 ; n18077
g17886 nor n17406 n17415 ; n18078
g17887 and asqrt[10] n18078 ; n18079
g17888 nor n17413 n18079 ; n18080
g17889 nor n18077 n18080 ; n18081
g17890 nor asqrt[37] n18062 ; n18082
g17891 and n18072_not n18082 ; n18083
g17892 nor n18081 n18083 ; n18084
g17893 nor n18074 n18084 ; n18085
g17894 and asqrt[38] n18085_not ; n18086
g17895 and n17425 n17427_not ; n18087
g17896 and n17418_not n18087 ; n18088
g17897 and asqrt[10] n18088 ; n18089
g17898 nor n17418 n17427 ; n18090
g17899 and asqrt[10] n18090 ; n18091
g17900 nor n17425 n18091 ; n18092
g17901 nor n18089 n18092 ; n18093
g17902 nor asqrt[38] n18074 ; n18094
g17903 and n18084_not n18094 ; n18095
g17904 nor n18093 n18095 ; n18096
g17905 nor n18086 n18096 ; n18097
g17906 and asqrt[39] n18097_not ; n18098
g17907 and n17430_not n17437 ; n18099
g17908 and n17439_not n18099 ; n18100
g17909 and asqrt[10] n18100 ; n18101
g17910 nor n17430 n17439 ; n18102
g17911 and asqrt[10] n18102 ; n18103
g17912 nor n17437 n18103 ; n18104
g17913 nor n18101 n18104 ; n18105
g17914 nor asqrt[39] n18086 ; n18106
g17915 and n18096_not n18106 ; n18107
g17916 nor n18105 n18107 ; n18108
g17917 nor n18098 n18108 ; n18109
g17918 and asqrt[40] n18109_not ; n18110
g17919 and n17449 n17451_not ; n18111
g17920 and n17442_not n18111 ; n18112
g17921 and asqrt[10] n18112 ; n18113
g17922 nor n17442 n17451 ; n18114
g17923 and asqrt[10] n18114 ; n18115
g17924 nor n17449 n18115 ; n18116
g17925 nor n18113 n18116 ; n18117
g17926 nor asqrt[40] n18098 ; n18118
g17927 and n18108_not n18118 ; n18119
g17928 nor n18117 n18119 ; n18120
g17929 nor n18110 n18120 ; n18121
g17930 and asqrt[41] n18121_not ; n18122
g17931 and n17454_not n17461 ; n18123
g17932 and n17463_not n18123 ; n18124
g17933 and asqrt[10] n18124 ; n18125
g17934 nor n17454 n17463 ; n18126
g17935 and asqrt[10] n18126 ; n18127
g17936 nor n17461 n18127 ; n18128
g17937 nor n18125 n18128 ; n18129
g17938 nor asqrt[41] n18110 ; n18130
g17939 and n18120_not n18130 ; n18131
g17940 nor n18129 n18131 ; n18132
g17941 nor n18122 n18132 ; n18133
g17942 and asqrt[42] n18133_not ; n18134
g17943 and n17473 n17475_not ; n18135
g17944 and n17466_not n18135 ; n18136
g17945 and asqrt[10] n18136 ; n18137
g17946 nor n17466 n17475 ; n18138
g17947 and asqrt[10] n18138 ; n18139
g17948 nor n17473 n18139 ; n18140
g17949 nor n18137 n18140 ; n18141
g17950 nor asqrt[42] n18122 ; n18142
g17951 and n18132_not n18142 ; n18143
g17952 nor n18141 n18143 ; n18144
g17953 nor n18134 n18144 ; n18145
g17954 and asqrt[43] n18145_not ; n18146
g17955 and n17478_not n17485 ; n18147
g17956 and n17487_not n18147 ; n18148
g17957 and asqrt[10] n18148 ; n18149
g17958 nor n17478 n17487 ; n18150
g17959 and asqrt[10] n18150 ; n18151
g17960 nor n17485 n18151 ; n18152
g17961 nor n18149 n18152 ; n18153
g17962 nor asqrt[43] n18134 ; n18154
g17963 and n18144_not n18154 ; n18155
g17964 nor n18153 n18155 ; n18156
g17965 nor n18146 n18156 ; n18157
g17966 and asqrt[44] n18157_not ; n18158
g17967 and n17497 n17499_not ; n18159
g17968 and n17490_not n18159 ; n18160
g17969 and asqrt[10] n18160 ; n18161
g17970 nor n17490 n17499 ; n18162
g17971 and asqrt[10] n18162 ; n18163
g17972 nor n17497 n18163 ; n18164
g17973 nor n18161 n18164 ; n18165
g17974 nor asqrt[44] n18146 ; n18166
g17975 and n18156_not n18166 ; n18167
g17976 nor n18165 n18167 ; n18168
g17977 nor n18158 n18168 ; n18169
g17978 and asqrt[45] n18169_not ; n18170
g17979 and n17502_not n17509 ; n18171
g17980 and n17511_not n18171 ; n18172
g17981 and asqrt[10] n18172 ; n18173
g17982 nor n17502 n17511 ; n18174
g17983 and asqrt[10] n18174 ; n18175
g17984 nor n17509 n18175 ; n18176
g17985 nor n18173 n18176 ; n18177
g17986 nor asqrt[45] n18158 ; n18178
g17987 and n18168_not n18178 ; n18179
g17988 nor n18177 n18179 ; n18180
g17989 nor n18170 n18180 ; n18181
g17990 and asqrt[46] n18181_not ; n18182
g17991 and n17521 n17523_not ; n18183
g17992 and n17514_not n18183 ; n18184
g17993 and asqrt[10] n18184 ; n18185
g17994 nor n17514 n17523 ; n18186
g17995 and asqrt[10] n18186 ; n18187
g17996 nor n17521 n18187 ; n18188
g17997 nor n18185 n18188 ; n18189
g17998 nor asqrt[46] n18170 ; n18190
g17999 and n18180_not n18190 ; n18191
g18000 nor n18189 n18191 ; n18192
g18001 nor n18182 n18192 ; n18193
g18002 and asqrt[47] n18193_not ; n18194
g18003 and n17526_not n17533 ; n18195
g18004 and n17535_not n18195 ; n18196
g18005 and asqrt[10] n18196 ; n18197
g18006 nor n17526 n17535 ; n18198
g18007 and asqrt[10] n18198 ; n18199
g18008 nor n17533 n18199 ; n18200
g18009 nor n18197 n18200 ; n18201
g18010 nor asqrt[47] n18182 ; n18202
g18011 and n18192_not n18202 ; n18203
g18012 nor n18201 n18203 ; n18204
g18013 nor n18194 n18204 ; n18205
g18014 and asqrt[48] n18205_not ; n18206
g18015 and n17545 n17547_not ; n18207
g18016 and n17538_not n18207 ; n18208
g18017 and asqrt[10] n18208 ; n18209
g18018 nor n17538 n17547 ; n18210
g18019 and asqrt[10] n18210 ; n18211
g18020 nor n17545 n18211 ; n18212
g18021 nor n18209 n18212 ; n18213
g18022 nor asqrt[48] n18194 ; n18214
g18023 and n18204_not n18214 ; n18215
g18024 nor n18213 n18215 ; n18216
g18025 nor n18206 n18216 ; n18217
g18026 and asqrt[49] n18217_not ; n18218
g18027 and n17550_not n17557 ; n18219
g18028 and n17559_not n18219 ; n18220
g18029 and asqrt[10] n18220 ; n18221
g18030 nor n17550 n17559 ; n18222
g18031 and asqrt[10] n18222 ; n18223
g18032 nor n17557 n18223 ; n18224
g18033 nor n18221 n18224 ; n18225
g18034 nor asqrt[49] n18206 ; n18226
g18035 and n18216_not n18226 ; n18227
g18036 nor n18225 n18227 ; n18228
g18037 nor n18218 n18228 ; n18229
g18038 and asqrt[50] n18229_not ; n18230
g18039 and n17569 n17571_not ; n18231
g18040 and n17562_not n18231 ; n18232
g18041 and asqrt[10] n18232 ; n18233
g18042 nor n17562 n17571 ; n18234
g18043 and asqrt[10] n18234 ; n18235
g18044 nor n17569 n18235 ; n18236
g18045 nor n18233 n18236 ; n18237
g18046 nor asqrt[50] n18218 ; n18238
g18047 and n18228_not n18238 ; n18239
g18048 nor n18237 n18239 ; n18240
g18049 nor n18230 n18240 ; n18241
g18050 and asqrt[51] n18241_not ; n18242
g18051 and n17574_not n17581 ; n18243
g18052 and n17583_not n18243 ; n18244
g18053 and asqrt[10] n18244 ; n18245
g18054 nor n17574 n17583 ; n18246
g18055 and asqrt[10] n18246 ; n18247
g18056 nor n17581 n18247 ; n18248
g18057 nor n18245 n18248 ; n18249
g18058 nor asqrt[51] n18230 ; n18250
g18059 and n18240_not n18250 ; n18251
g18060 nor n18249 n18251 ; n18252
g18061 nor n18242 n18252 ; n18253
g18062 and asqrt[52] n18253_not ; n18254
g18063 and n17593 n17595_not ; n18255
g18064 and n17586_not n18255 ; n18256
g18065 and asqrt[10] n18256 ; n18257
g18066 nor n17586 n17595 ; n18258
g18067 and asqrt[10] n18258 ; n18259
g18068 nor n17593 n18259 ; n18260
g18069 nor n18257 n18260 ; n18261
g18070 nor asqrt[52] n18242 ; n18262
g18071 and n18252_not n18262 ; n18263
g18072 nor n18261 n18263 ; n18264
g18073 nor n18254 n18264 ; n18265
g18074 and asqrt[53] n18265_not ; n18266
g18075 and n17598_not n17605 ; n18267
g18076 and n17607_not n18267 ; n18268
g18077 and asqrt[10] n18268 ; n18269
g18078 nor n17598 n17607 ; n18270
g18079 and asqrt[10] n18270 ; n18271
g18080 nor n17605 n18271 ; n18272
g18081 nor n18269 n18272 ; n18273
g18082 nor asqrt[53] n18254 ; n18274
g18083 and n18264_not n18274 ; n18275
g18084 nor n18273 n18275 ; n18276
g18085 nor n18266 n18276 ; n18277
g18086 and asqrt[54] n18277_not ; n18278
g18087 and n17617 n17619_not ; n18279
g18088 and n17610_not n18279 ; n18280
g18089 and asqrt[10] n18280 ; n18281
g18090 nor n17610 n17619 ; n18282
g18091 and asqrt[10] n18282 ; n18283
g18092 nor n17617 n18283 ; n18284
g18093 nor n18281 n18284 ; n18285
g18094 nor asqrt[54] n18266 ; n18286
g18095 and n18276_not n18286 ; n18287
g18096 nor n18285 n18287 ; n18288
g18097 nor n18278 n18288 ; n18289
g18098 and asqrt[55] n18289_not ; n18290
g18099 nor asqrt[55] n18278 ; n18291
g18100 and n18288_not n18291 ; n18292
g18101 and n17622_not n17631 ; n18293
g18102 and n17624_not n18293 ; n18294
g18103 and asqrt[10] n18294 ; n18295
g18104 nor n17622 n17624 ; n18296
g18105 and asqrt[10] n18296 ; n18297
g18106 nor n17631 n18297 ; n18298
g18107 nor n18295 n18298 ; n18299
g18108 nor n18292 n18299 ; n18300
g18109 nor n18290 n18300 ; n18301
g18110 and asqrt[56] n18301_not ; n18302
g18111 and n17641 n17643_not ; n18303
g18112 and n17634_not n18303 ; n18304
g18113 and asqrt[10] n18304 ; n18305
g18114 nor n17634 n17643 ; n18306
g18115 and asqrt[10] n18306 ; n18307
g18116 nor n17641 n18307 ; n18308
g18117 nor n18305 n18308 ; n18309
g18118 nor asqrt[56] n18290 ; n18310
g18119 and n18300_not n18310 ; n18311
g18120 nor n18309 n18311 ; n18312
g18121 nor n18302 n18312 ; n18313
g18122 and asqrt[57] n18313_not ; n18314
g18123 and n17646_not n17653 ; n18315
g18124 and n17655_not n18315 ; n18316
g18125 and asqrt[10] n18316 ; n18317
g18126 nor n17646 n17655 ; n18318
g18127 and asqrt[10] n18318 ; n18319
g18128 nor n17653 n18319 ; n18320
g18129 nor n18317 n18320 ; n18321
g18130 nor asqrt[57] n18302 ; n18322
g18131 and n18312_not n18322 ; n18323
g18132 nor n18321 n18323 ; n18324
g18133 nor n18314 n18324 ; n18325
g18134 and asqrt[58] n18325_not ; n18326
g18135 and n17665 n17667_not ; n18327
g18136 and n17658_not n18327 ; n18328
g18137 and asqrt[10] n18328 ; n18329
g18138 nor n17658 n17667 ; n18330
g18139 and asqrt[10] n18330 ; n18331
g18140 nor n17665 n18331 ; n18332
g18141 nor n18329 n18332 ; n18333
g18142 nor asqrt[58] n18314 ; n18334
g18143 and n18324_not n18334 ; n18335
g18144 nor n18333 n18335 ; n18336
g18145 nor n18326 n18336 ; n18337
g18146 and asqrt[59] n18337_not ; n18338
g18147 and n17670_not n17677 ; n18339
g18148 and n17679_not n18339 ; n18340
g18149 and asqrt[10] n18340 ; n18341
g18150 nor n17670 n17679 ; n18342
g18151 and asqrt[10] n18342 ; n18343
g18152 nor n17677 n18343 ; n18344
g18153 nor n18341 n18344 ; n18345
g18154 nor asqrt[59] n18326 ; n18346
g18155 and n18336_not n18346 ; n18347
g18156 nor n18345 n18347 ; n18348
g18157 nor n18338 n18348 ; n18349
g18158 and asqrt[60] n18349_not ; n18350
g18159 and n17689 n17691_not ; n18351
g18160 and n17682_not n18351 ; n18352
g18161 and asqrt[10] n18352 ; n18353
g18162 nor n17682 n17691 ; n18354
g18163 and asqrt[10] n18354 ; n18355
g18164 nor n17689 n18355 ; n18356
g18165 nor n18353 n18356 ; n18357
g18166 nor asqrt[60] n18338 ; n18358
g18167 and n18348_not n18358 ; n18359
g18168 nor n18357 n18359 ; n18360
g18169 nor n18350 n18360 ; n18361
g18170 and asqrt[61] n18361_not ; n18362
g18171 and n17694_not n17701 ; n18363
g18172 and n17703_not n18363 ; n18364
g18173 and asqrt[10] n18364 ; n18365
g18174 nor n17694 n17703 ; n18366
g18175 and asqrt[10] n18366 ; n18367
g18176 nor n17701 n18367 ; n18368
g18177 nor n18365 n18368 ; n18369
g18178 nor asqrt[61] n18350 ; n18370
g18179 and n18360_not n18370 ; n18371
g18180 nor n18369 n18371 ; n18372
g18181 nor n18362 n18372 ; n18373
g18182 and asqrt[62] n18373_not ; n18374
g18183 and n17713 n17715_not ; n18375
g18184 and n17706_not n18375 ; n18376
g18185 and asqrt[10] n18376 ; n18377
g18186 nor n17706 n17715 ; n18378
g18187 and asqrt[10] n18378 ; n18379
g18188 nor n17713 n18379 ; n18380
g18189 nor n18377 n18380 ; n18381
g18190 nor asqrt[62] n18362 ; n18382
g18191 and n18372_not n18382 ; n18383
g18192 nor n18381 n18383 ; n18384
g18193 nor n18374 n18384 ; n18385
g18194 and n17718_not n17725 ; n18386
g18195 and n17727_not n18386 ; n18387
g18196 and asqrt[10] n18387 ; n18388
g18197 nor n17718 n17727 ; n18389
g18198 and asqrt[10] n18389 ; n18390
g18199 nor n17725 n18390 ; n18391
g18200 nor n18388 n18391 ; n18392
g18201 nor n17729 n17736 ; n18393
g18202 and asqrt[10] n18393 ; n18394
g18203 nor n17744 n18394 ; n18395
g18204 and n18392_not n18395 ; n18396
g18205 and n18385_not n18396 ; n18397
g18206 nor asqrt[63] n18397 ; n18398
g18207 and n18374_not n18392 ; n18399
g18208 and n18384_not n18399 ; n18400
g18209 and n17736_not asqrt[10] ; n18401
g18210 and n17729 n18401_not ; n18402
g18211 and asqrt[63] n18393_not ; n18403
g18212 and n18402_not n18403 ; n18404
g18213 nor n17732 n17753 ; n18405
g18214 and n17735_not n18405 ; n18406
g18215 and n17748_not n18406 ; n18407
g18216 and n17744_not n18407 ; n18408
g18217 and n17742_not n18408 ; n18409
g18218 nor n18404 n18409 ; n18410
g18219 and n18400_not n18410 ; n18411
g18220 nand n18398_not n18411 ; asqrt[9]
g18221 and a[18] asqrt[9] ; n18413
g18222 nor a[16] a[17] ; n18414
g18223 and a[18]_not n18414 ; n18415
g18224 nor n18413 n18415 ; n18416
g18225 and asqrt[10] n18416_not ; n18417
g18226 nor n17753 n18415 ; n18418
g18227 and n17748_not n18418 ; n18419
g18228 and n17744_not n18419 ; n18420
g18229 and n17742_not n18420 ; n18421
g18230 and n18413_not n18421 ; n18422
g18231 and a[18]_not asqrt[9] ; n18423
g18232 and a[19] n18423_not ; n18424
g18233 and n17758 asqrt[9] ; n18425
g18234 nor n18424 n18425 ; n18426
g18235 and n18422_not n18426 ; n18427
g18236 nor n18417 n18427 ; n18428
g18237 and asqrt[11] n18428_not ; n18429
g18238 nor asqrt[11] n18417 ; n18430
g18239 and n18427_not n18430 ; n18431
g18240 and asqrt[10] n18409_not ; n18432
g18241 and n18404_not n18432 ; n18433
g18242 and n18400_not n18433 ; n18434
g18243 and n18398_not n18434 ; n18435
g18244 nor n18425 n18435 ; n18436
g18245 and a[20] n18436_not ; n18437
g18246 nor a[20] n18435 ; n18438
g18247 and n18425_not n18438 ; n18439
g18248 nor n18437 n18439 ; n18440
g18249 nor n18431 n18440 ; n18441
g18250 nor n18429 n18441 ; n18442
g18251 and asqrt[12] n18442_not ; n18443
g18252 nor n17761 n17766 ; n18444
g18253 and n17770_not n18444 ; n18445
g18254 and asqrt[9] n18445 ; n18446
g18255 and asqrt[9] n18444 ; n18447
g18256 and n17770 n18447_not ; n18448
g18257 nor n18446 n18448 ; n18449
g18258 nor asqrt[12] n18429 ; n18450
g18259 and n18441_not n18450 ; n18451
g18260 nor n18449 n18451 ; n18452
g18261 nor n18443 n18452 ; n18453
g18262 and asqrt[13] n18453_not ; n18454
g18263 and n17775_not n17784 ; n18455
g18264 and n17773_not n18455 ; n18456
g18265 and asqrt[9] n18456 ; n18457
g18266 nor n17773 n17775 ; n18458
g18267 and asqrt[9] n18458 ; n18459
g18268 nor n17784 n18459 ; n18460
g18269 nor n18457 n18460 ; n18461
g18270 nor asqrt[13] n18443 ; n18462
g18271 and n18452_not n18462 ; n18463
g18272 nor n18461 n18463 ; n18464
g18273 nor n18454 n18464 ; n18465
g18274 and asqrt[14] n18465_not ; n18466
g18275 and n17787_not n17793 ; n18467
g18276 and n17795_not n18467 ; n18468
g18277 and asqrt[9] n18468 ; n18469
g18278 nor n17787 n17795 ; n18470
g18279 and asqrt[9] n18470 ; n18471
g18280 nor n17793 n18471 ; n18472
g18281 nor n18469 n18472 ; n18473
g18282 nor asqrt[14] n18454 ; n18474
g18283 and n18464_not n18474 ; n18475
g18284 nor n18473 n18475 ; n18476
g18285 nor n18466 n18476 ; n18477
g18286 and asqrt[15] n18477_not ; n18478
g18287 and n17805 n17807_not ; n18479
g18288 and n17798_not n18479 ; n18480
g18289 and asqrt[9] n18480 ; n18481
g18290 nor n17798 n17807 ; n18482
g18291 and asqrt[9] n18482 ; n18483
g18292 nor n17805 n18483 ; n18484
g18293 nor n18481 n18484 ; n18485
g18294 nor asqrt[15] n18466 ; n18486
g18295 and n18476_not n18486 ; n18487
g18296 nor n18485 n18487 ; n18488
g18297 nor n18478 n18488 ; n18489
g18298 and asqrt[16] n18489_not ; n18490
g18299 and n17810_not n17817 ; n18491
g18300 and n17819_not n18491 ; n18492
g18301 and asqrt[9] n18492 ; n18493
g18302 nor n17810 n17819 ; n18494
g18303 and asqrt[9] n18494 ; n18495
g18304 nor n17817 n18495 ; n18496
g18305 nor n18493 n18496 ; n18497
g18306 nor asqrt[16] n18478 ; n18498
g18307 and n18488_not n18498 ; n18499
g18308 nor n18497 n18499 ; n18500
g18309 nor n18490 n18500 ; n18501
g18310 and asqrt[17] n18501_not ; n18502
g18311 and n17829 n17831_not ; n18503
g18312 and n17822_not n18503 ; n18504
g18313 and asqrt[9] n18504 ; n18505
g18314 nor n17822 n17831 ; n18506
g18315 and asqrt[9] n18506 ; n18507
g18316 nor n17829 n18507 ; n18508
g18317 nor n18505 n18508 ; n18509
g18318 nor asqrt[17] n18490 ; n18510
g18319 and n18500_not n18510 ; n18511
g18320 nor n18509 n18511 ; n18512
g18321 nor n18502 n18512 ; n18513
g18322 and asqrt[18] n18513_not ; n18514
g18323 and n17834_not n17841 ; n18515
g18324 and n17843_not n18515 ; n18516
g18325 and asqrt[9] n18516 ; n18517
g18326 nor n17834 n17843 ; n18518
g18327 and asqrt[9] n18518 ; n18519
g18328 nor n17841 n18519 ; n18520
g18329 nor n18517 n18520 ; n18521
g18330 nor asqrt[18] n18502 ; n18522
g18331 and n18512_not n18522 ; n18523
g18332 nor n18521 n18523 ; n18524
g18333 nor n18514 n18524 ; n18525
g18334 and asqrt[19] n18525_not ; n18526
g18335 and n17853 n17855_not ; n18527
g18336 and n17846_not n18527 ; n18528
g18337 and asqrt[9] n18528 ; n18529
g18338 nor n17846 n17855 ; n18530
g18339 and asqrt[9] n18530 ; n18531
g18340 nor n17853 n18531 ; n18532
g18341 nor n18529 n18532 ; n18533
g18342 nor asqrt[19] n18514 ; n18534
g18343 and n18524_not n18534 ; n18535
g18344 nor n18533 n18535 ; n18536
g18345 nor n18526 n18536 ; n18537
g18346 and asqrt[20] n18537_not ; n18538
g18347 and n17858_not n17865 ; n18539
g18348 and n17867_not n18539 ; n18540
g18349 and asqrt[9] n18540 ; n18541
g18350 nor n17858 n17867 ; n18542
g18351 and asqrt[9] n18542 ; n18543
g18352 nor n17865 n18543 ; n18544
g18353 nor n18541 n18544 ; n18545
g18354 nor asqrt[20] n18526 ; n18546
g18355 and n18536_not n18546 ; n18547
g18356 nor n18545 n18547 ; n18548
g18357 nor n18538 n18548 ; n18549
g18358 and asqrt[21] n18549_not ; n18550
g18359 and n17877 n17879_not ; n18551
g18360 and n17870_not n18551 ; n18552
g18361 and asqrt[9] n18552 ; n18553
g18362 nor n17870 n17879 ; n18554
g18363 and asqrt[9] n18554 ; n18555
g18364 nor n17877 n18555 ; n18556
g18365 nor n18553 n18556 ; n18557
g18366 nor asqrt[21] n18538 ; n18558
g18367 and n18548_not n18558 ; n18559
g18368 nor n18557 n18559 ; n18560
g18369 nor n18550 n18560 ; n18561
g18370 and asqrt[22] n18561_not ; n18562
g18371 and n17882_not n17889 ; n18563
g18372 and n17891_not n18563 ; n18564
g18373 and asqrt[9] n18564 ; n18565
g18374 nor n17882 n17891 ; n18566
g18375 and asqrt[9] n18566 ; n18567
g18376 nor n17889 n18567 ; n18568
g18377 nor n18565 n18568 ; n18569
g18378 nor asqrt[22] n18550 ; n18570
g18379 and n18560_not n18570 ; n18571
g18380 nor n18569 n18571 ; n18572
g18381 nor n18562 n18572 ; n18573
g18382 and asqrt[23] n18573_not ; n18574
g18383 and n17901 n17903_not ; n18575
g18384 and n17894_not n18575 ; n18576
g18385 and asqrt[9] n18576 ; n18577
g18386 nor n17894 n17903 ; n18578
g18387 and asqrt[9] n18578 ; n18579
g18388 nor n17901 n18579 ; n18580
g18389 nor n18577 n18580 ; n18581
g18390 nor asqrt[23] n18562 ; n18582
g18391 and n18572_not n18582 ; n18583
g18392 nor n18581 n18583 ; n18584
g18393 nor n18574 n18584 ; n18585
g18394 and asqrt[24] n18585_not ; n18586
g18395 and n17906_not n17913 ; n18587
g18396 and n17915_not n18587 ; n18588
g18397 and asqrt[9] n18588 ; n18589
g18398 nor n17906 n17915 ; n18590
g18399 and asqrt[9] n18590 ; n18591
g18400 nor n17913 n18591 ; n18592
g18401 nor n18589 n18592 ; n18593
g18402 nor asqrt[24] n18574 ; n18594
g18403 and n18584_not n18594 ; n18595
g18404 nor n18593 n18595 ; n18596
g18405 nor n18586 n18596 ; n18597
g18406 and asqrt[25] n18597_not ; n18598
g18407 and n17925 n17927_not ; n18599
g18408 and n17918_not n18599 ; n18600
g18409 and asqrt[9] n18600 ; n18601
g18410 nor n17918 n17927 ; n18602
g18411 and asqrt[9] n18602 ; n18603
g18412 nor n17925 n18603 ; n18604
g18413 nor n18601 n18604 ; n18605
g18414 nor asqrt[25] n18586 ; n18606
g18415 and n18596_not n18606 ; n18607
g18416 nor n18605 n18607 ; n18608
g18417 nor n18598 n18608 ; n18609
g18418 and asqrt[26] n18609_not ; n18610
g18419 and n17930_not n17937 ; n18611
g18420 and n17939_not n18611 ; n18612
g18421 and asqrt[9] n18612 ; n18613
g18422 nor n17930 n17939 ; n18614
g18423 and asqrt[9] n18614 ; n18615
g18424 nor n17937 n18615 ; n18616
g18425 nor n18613 n18616 ; n18617
g18426 nor asqrt[26] n18598 ; n18618
g18427 and n18608_not n18618 ; n18619
g18428 nor n18617 n18619 ; n18620
g18429 nor n18610 n18620 ; n18621
g18430 and asqrt[27] n18621_not ; n18622
g18431 and n17949 n17951_not ; n18623
g18432 and n17942_not n18623 ; n18624
g18433 and asqrt[9] n18624 ; n18625
g18434 nor n17942 n17951 ; n18626
g18435 and asqrt[9] n18626 ; n18627
g18436 nor n17949 n18627 ; n18628
g18437 nor n18625 n18628 ; n18629
g18438 nor asqrt[27] n18610 ; n18630
g18439 and n18620_not n18630 ; n18631
g18440 nor n18629 n18631 ; n18632
g18441 nor n18622 n18632 ; n18633
g18442 and asqrt[28] n18633_not ; n18634
g18443 and n17954_not n17961 ; n18635
g18444 and n17963_not n18635 ; n18636
g18445 and asqrt[9] n18636 ; n18637
g18446 nor n17954 n17963 ; n18638
g18447 and asqrt[9] n18638 ; n18639
g18448 nor n17961 n18639 ; n18640
g18449 nor n18637 n18640 ; n18641
g18450 nor asqrt[28] n18622 ; n18642
g18451 and n18632_not n18642 ; n18643
g18452 nor n18641 n18643 ; n18644
g18453 nor n18634 n18644 ; n18645
g18454 and asqrt[29] n18645_not ; n18646
g18455 and n17973 n17975_not ; n18647
g18456 and n17966_not n18647 ; n18648
g18457 and asqrt[9] n18648 ; n18649
g18458 nor n17966 n17975 ; n18650
g18459 and asqrt[9] n18650 ; n18651
g18460 nor n17973 n18651 ; n18652
g18461 nor n18649 n18652 ; n18653
g18462 nor asqrt[29] n18634 ; n18654
g18463 and n18644_not n18654 ; n18655
g18464 nor n18653 n18655 ; n18656
g18465 nor n18646 n18656 ; n18657
g18466 and asqrt[30] n18657_not ; n18658
g18467 and n17978_not n17985 ; n18659
g18468 and n17987_not n18659 ; n18660
g18469 and asqrt[9] n18660 ; n18661
g18470 nor n17978 n17987 ; n18662
g18471 and asqrt[9] n18662 ; n18663
g18472 nor n17985 n18663 ; n18664
g18473 nor n18661 n18664 ; n18665
g18474 nor asqrt[30] n18646 ; n18666
g18475 and n18656_not n18666 ; n18667
g18476 nor n18665 n18667 ; n18668
g18477 nor n18658 n18668 ; n18669
g18478 and asqrt[31] n18669_not ; n18670
g18479 and n17997 n17999_not ; n18671
g18480 and n17990_not n18671 ; n18672
g18481 and asqrt[9] n18672 ; n18673
g18482 nor n17990 n17999 ; n18674
g18483 and asqrt[9] n18674 ; n18675
g18484 nor n17997 n18675 ; n18676
g18485 nor n18673 n18676 ; n18677
g18486 nor asqrt[31] n18658 ; n18678
g18487 and n18668_not n18678 ; n18679
g18488 nor n18677 n18679 ; n18680
g18489 nor n18670 n18680 ; n18681
g18490 and asqrt[32] n18681_not ; n18682
g18491 and n18002_not n18009 ; n18683
g18492 and n18011_not n18683 ; n18684
g18493 and asqrt[9] n18684 ; n18685
g18494 nor n18002 n18011 ; n18686
g18495 and asqrt[9] n18686 ; n18687
g18496 nor n18009 n18687 ; n18688
g18497 nor n18685 n18688 ; n18689
g18498 nor asqrt[32] n18670 ; n18690
g18499 and n18680_not n18690 ; n18691
g18500 nor n18689 n18691 ; n18692
g18501 nor n18682 n18692 ; n18693
g18502 and asqrt[33] n18693_not ; n18694
g18503 and n18021 n18023_not ; n18695
g18504 and n18014_not n18695 ; n18696
g18505 and asqrt[9] n18696 ; n18697
g18506 nor n18014 n18023 ; n18698
g18507 and asqrt[9] n18698 ; n18699
g18508 nor n18021 n18699 ; n18700
g18509 nor n18697 n18700 ; n18701
g18510 nor asqrt[33] n18682 ; n18702
g18511 and n18692_not n18702 ; n18703
g18512 nor n18701 n18703 ; n18704
g18513 nor n18694 n18704 ; n18705
g18514 and asqrt[34] n18705_not ; n18706
g18515 and n18026_not n18033 ; n18707
g18516 and n18035_not n18707 ; n18708
g18517 and asqrt[9] n18708 ; n18709
g18518 nor n18026 n18035 ; n18710
g18519 and asqrt[9] n18710 ; n18711
g18520 nor n18033 n18711 ; n18712
g18521 nor n18709 n18712 ; n18713
g18522 nor asqrt[34] n18694 ; n18714
g18523 and n18704_not n18714 ; n18715
g18524 nor n18713 n18715 ; n18716
g18525 nor n18706 n18716 ; n18717
g18526 and asqrt[35] n18717_not ; n18718
g18527 and n18045 n18047_not ; n18719
g18528 and n18038_not n18719 ; n18720
g18529 and asqrt[9] n18720 ; n18721
g18530 nor n18038 n18047 ; n18722
g18531 and asqrt[9] n18722 ; n18723
g18532 nor n18045 n18723 ; n18724
g18533 nor n18721 n18724 ; n18725
g18534 nor asqrt[35] n18706 ; n18726
g18535 and n18716_not n18726 ; n18727
g18536 nor n18725 n18727 ; n18728
g18537 nor n18718 n18728 ; n18729
g18538 and asqrt[36] n18729_not ; n18730
g18539 and n18050_not n18057 ; n18731
g18540 and n18059_not n18731 ; n18732
g18541 and asqrt[9] n18732 ; n18733
g18542 nor n18050 n18059 ; n18734
g18543 and asqrt[9] n18734 ; n18735
g18544 nor n18057 n18735 ; n18736
g18545 nor n18733 n18736 ; n18737
g18546 nor asqrt[36] n18718 ; n18738
g18547 and n18728_not n18738 ; n18739
g18548 nor n18737 n18739 ; n18740
g18549 nor n18730 n18740 ; n18741
g18550 and asqrt[37] n18741_not ; n18742
g18551 and n18069 n18071_not ; n18743
g18552 and n18062_not n18743 ; n18744
g18553 and asqrt[9] n18744 ; n18745
g18554 nor n18062 n18071 ; n18746
g18555 and asqrt[9] n18746 ; n18747
g18556 nor n18069 n18747 ; n18748
g18557 nor n18745 n18748 ; n18749
g18558 nor asqrt[37] n18730 ; n18750
g18559 and n18740_not n18750 ; n18751
g18560 nor n18749 n18751 ; n18752
g18561 nor n18742 n18752 ; n18753
g18562 and asqrt[38] n18753_not ; n18754
g18563 and n18074_not n18081 ; n18755
g18564 and n18083_not n18755 ; n18756
g18565 and asqrt[9] n18756 ; n18757
g18566 nor n18074 n18083 ; n18758
g18567 and asqrt[9] n18758 ; n18759
g18568 nor n18081 n18759 ; n18760
g18569 nor n18757 n18760 ; n18761
g18570 nor asqrt[38] n18742 ; n18762
g18571 and n18752_not n18762 ; n18763
g18572 nor n18761 n18763 ; n18764
g18573 nor n18754 n18764 ; n18765
g18574 and asqrt[39] n18765_not ; n18766
g18575 and n18093 n18095_not ; n18767
g18576 and n18086_not n18767 ; n18768
g18577 and asqrt[9] n18768 ; n18769
g18578 nor n18086 n18095 ; n18770
g18579 and asqrt[9] n18770 ; n18771
g18580 nor n18093 n18771 ; n18772
g18581 nor n18769 n18772 ; n18773
g18582 nor asqrt[39] n18754 ; n18774
g18583 and n18764_not n18774 ; n18775
g18584 nor n18773 n18775 ; n18776
g18585 nor n18766 n18776 ; n18777
g18586 and asqrt[40] n18777_not ; n18778
g18587 and n18098_not n18105 ; n18779
g18588 and n18107_not n18779 ; n18780
g18589 and asqrt[9] n18780 ; n18781
g18590 nor n18098 n18107 ; n18782
g18591 and asqrt[9] n18782 ; n18783
g18592 nor n18105 n18783 ; n18784
g18593 nor n18781 n18784 ; n18785
g18594 nor asqrt[40] n18766 ; n18786
g18595 and n18776_not n18786 ; n18787
g18596 nor n18785 n18787 ; n18788
g18597 nor n18778 n18788 ; n18789
g18598 and asqrt[41] n18789_not ; n18790
g18599 and n18117 n18119_not ; n18791
g18600 and n18110_not n18791 ; n18792
g18601 and asqrt[9] n18792 ; n18793
g18602 nor n18110 n18119 ; n18794
g18603 and asqrt[9] n18794 ; n18795
g18604 nor n18117 n18795 ; n18796
g18605 nor n18793 n18796 ; n18797
g18606 nor asqrt[41] n18778 ; n18798
g18607 and n18788_not n18798 ; n18799
g18608 nor n18797 n18799 ; n18800
g18609 nor n18790 n18800 ; n18801
g18610 and asqrt[42] n18801_not ; n18802
g18611 and n18122_not n18129 ; n18803
g18612 and n18131_not n18803 ; n18804
g18613 and asqrt[9] n18804 ; n18805
g18614 nor n18122 n18131 ; n18806
g18615 and asqrt[9] n18806 ; n18807
g18616 nor n18129 n18807 ; n18808
g18617 nor n18805 n18808 ; n18809
g18618 nor asqrt[42] n18790 ; n18810
g18619 and n18800_not n18810 ; n18811
g18620 nor n18809 n18811 ; n18812
g18621 nor n18802 n18812 ; n18813
g18622 and asqrt[43] n18813_not ; n18814
g18623 and n18141 n18143_not ; n18815
g18624 and n18134_not n18815 ; n18816
g18625 and asqrt[9] n18816 ; n18817
g18626 nor n18134 n18143 ; n18818
g18627 and asqrt[9] n18818 ; n18819
g18628 nor n18141 n18819 ; n18820
g18629 nor n18817 n18820 ; n18821
g18630 nor asqrt[43] n18802 ; n18822
g18631 and n18812_not n18822 ; n18823
g18632 nor n18821 n18823 ; n18824
g18633 nor n18814 n18824 ; n18825
g18634 and asqrt[44] n18825_not ; n18826
g18635 and n18146_not n18153 ; n18827
g18636 and n18155_not n18827 ; n18828
g18637 and asqrt[9] n18828 ; n18829
g18638 nor n18146 n18155 ; n18830
g18639 and asqrt[9] n18830 ; n18831
g18640 nor n18153 n18831 ; n18832
g18641 nor n18829 n18832 ; n18833
g18642 nor asqrt[44] n18814 ; n18834
g18643 and n18824_not n18834 ; n18835
g18644 nor n18833 n18835 ; n18836
g18645 nor n18826 n18836 ; n18837
g18646 and asqrt[45] n18837_not ; n18838
g18647 and n18165 n18167_not ; n18839
g18648 and n18158_not n18839 ; n18840
g18649 and asqrt[9] n18840 ; n18841
g18650 nor n18158 n18167 ; n18842
g18651 and asqrt[9] n18842 ; n18843
g18652 nor n18165 n18843 ; n18844
g18653 nor n18841 n18844 ; n18845
g18654 nor asqrt[45] n18826 ; n18846
g18655 and n18836_not n18846 ; n18847
g18656 nor n18845 n18847 ; n18848
g18657 nor n18838 n18848 ; n18849
g18658 and asqrt[46] n18849_not ; n18850
g18659 and n18170_not n18177 ; n18851
g18660 and n18179_not n18851 ; n18852
g18661 and asqrt[9] n18852 ; n18853
g18662 nor n18170 n18179 ; n18854
g18663 and asqrt[9] n18854 ; n18855
g18664 nor n18177 n18855 ; n18856
g18665 nor n18853 n18856 ; n18857
g18666 nor asqrt[46] n18838 ; n18858
g18667 and n18848_not n18858 ; n18859
g18668 nor n18857 n18859 ; n18860
g18669 nor n18850 n18860 ; n18861
g18670 and asqrt[47] n18861_not ; n18862
g18671 and n18189 n18191_not ; n18863
g18672 and n18182_not n18863 ; n18864
g18673 and asqrt[9] n18864 ; n18865
g18674 nor n18182 n18191 ; n18866
g18675 and asqrt[9] n18866 ; n18867
g18676 nor n18189 n18867 ; n18868
g18677 nor n18865 n18868 ; n18869
g18678 nor asqrt[47] n18850 ; n18870
g18679 and n18860_not n18870 ; n18871
g18680 nor n18869 n18871 ; n18872
g18681 nor n18862 n18872 ; n18873
g18682 and asqrt[48] n18873_not ; n18874
g18683 and n18194_not n18201 ; n18875
g18684 and n18203_not n18875 ; n18876
g18685 and asqrt[9] n18876 ; n18877
g18686 nor n18194 n18203 ; n18878
g18687 and asqrt[9] n18878 ; n18879
g18688 nor n18201 n18879 ; n18880
g18689 nor n18877 n18880 ; n18881
g18690 nor asqrt[48] n18862 ; n18882
g18691 and n18872_not n18882 ; n18883
g18692 nor n18881 n18883 ; n18884
g18693 nor n18874 n18884 ; n18885
g18694 and asqrt[49] n18885_not ; n18886
g18695 and n18213 n18215_not ; n18887
g18696 and n18206_not n18887 ; n18888
g18697 and asqrt[9] n18888 ; n18889
g18698 nor n18206 n18215 ; n18890
g18699 and asqrt[9] n18890 ; n18891
g18700 nor n18213 n18891 ; n18892
g18701 nor n18889 n18892 ; n18893
g18702 nor asqrt[49] n18874 ; n18894
g18703 and n18884_not n18894 ; n18895
g18704 nor n18893 n18895 ; n18896
g18705 nor n18886 n18896 ; n18897
g18706 and asqrt[50] n18897_not ; n18898
g18707 and n18218_not n18225 ; n18899
g18708 and n18227_not n18899 ; n18900
g18709 and asqrt[9] n18900 ; n18901
g18710 nor n18218 n18227 ; n18902
g18711 and asqrt[9] n18902 ; n18903
g18712 nor n18225 n18903 ; n18904
g18713 nor n18901 n18904 ; n18905
g18714 nor asqrt[50] n18886 ; n18906
g18715 and n18896_not n18906 ; n18907
g18716 nor n18905 n18907 ; n18908
g18717 nor n18898 n18908 ; n18909
g18718 and asqrt[51] n18909_not ; n18910
g18719 and n18237 n18239_not ; n18911
g18720 and n18230_not n18911 ; n18912
g18721 and asqrt[9] n18912 ; n18913
g18722 nor n18230 n18239 ; n18914
g18723 and asqrt[9] n18914 ; n18915
g18724 nor n18237 n18915 ; n18916
g18725 nor n18913 n18916 ; n18917
g18726 nor asqrt[51] n18898 ; n18918
g18727 and n18908_not n18918 ; n18919
g18728 nor n18917 n18919 ; n18920
g18729 nor n18910 n18920 ; n18921
g18730 and asqrt[52] n18921_not ; n18922
g18731 and n18242_not n18249 ; n18923
g18732 and n18251_not n18923 ; n18924
g18733 and asqrt[9] n18924 ; n18925
g18734 nor n18242 n18251 ; n18926
g18735 and asqrt[9] n18926 ; n18927
g18736 nor n18249 n18927 ; n18928
g18737 nor n18925 n18928 ; n18929
g18738 nor asqrt[52] n18910 ; n18930
g18739 and n18920_not n18930 ; n18931
g18740 nor n18929 n18931 ; n18932
g18741 nor n18922 n18932 ; n18933
g18742 and asqrt[53] n18933_not ; n18934
g18743 and n18261 n18263_not ; n18935
g18744 and n18254_not n18935 ; n18936
g18745 and asqrt[9] n18936 ; n18937
g18746 nor n18254 n18263 ; n18938
g18747 and asqrt[9] n18938 ; n18939
g18748 nor n18261 n18939 ; n18940
g18749 nor n18937 n18940 ; n18941
g18750 nor asqrt[53] n18922 ; n18942
g18751 and n18932_not n18942 ; n18943
g18752 nor n18941 n18943 ; n18944
g18753 nor n18934 n18944 ; n18945
g18754 and asqrt[54] n18945_not ; n18946
g18755 and n18266_not n18273 ; n18947
g18756 and n18275_not n18947 ; n18948
g18757 and asqrt[9] n18948 ; n18949
g18758 nor n18266 n18275 ; n18950
g18759 and asqrt[9] n18950 ; n18951
g18760 nor n18273 n18951 ; n18952
g18761 nor n18949 n18952 ; n18953
g18762 nor asqrt[54] n18934 ; n18954
g18763 and n18944_not n18954 ; n18955
g18764 nor n18953 n18955 ; n18956
g18765 nor n18946 n18956 ; n18957
g18766 and asqrt[55] n18957_not ; n18958
g18767 and n18285 n18287_not ; n18959
g18768 and n18278_not n18959 ; n18960
g18769 and asqrt[9] n18960 ; n18961
g18770 nor n18278 n18287 ; n18962
g18771 and asqrt[9] n18962 ; n18963
g18772 nor n18285 n18963 ; n18964
g18773 nor n18961 n18964 ; n18965
g18774 nor asqrt[55] n18946 ; n18966
g18775 and n18956_not n18966 ; n18967
g18776 nor n18965 n18967 ; n18968
g18777 nor n18958 n18968 ; n18969
g18778 and asqrt[56] n18969_not ; n18970
g18779 nor asqrt[56] n18958 ; n18971
g18780 and n18968_not n18971 ; n18972
g18781 and n18290_not n18299 ; n18973
g18782 and n18292_not n18973 ; n18974
g18783 and asqrt[9] n18974 ; n18975
g18784 nor n18290 n18292 ; n18976
g18785 and asqrt[9] n18976 ; n18977
g18786 nor n18299 n18977 ; n18978
g18787 nor n18975 n18978 ; n18979
g18788 nor n18972 n18979 ; n18980
g18789 nor n18970 n18980 ; n18981
g18790 and asqrt[57] n18981_not ; n18982
g18791 and n18309 n18311_not ; n18983
g18792 and n18302_not n18983 ; n18984
g18793 and asqrt[9] n18984 ; n18985
g18794 nor n18302 n18311 ; n18986
g18795 and asqrt[9] n18986 ; n18987
g18796 nor n18309 n18987 ; n18988
g18797 nor n18985 n18988 ; n18989
g18798 nor asqrt[57] n18970 ; n18990
g18799 and n18980_not n18990 ; n18991
g18800 nor n18989 n18991 ; n18992
g18801 nor n18982 n18992 ; n18993
g18802 and asqrt[58] n18993_not ; n18994
g18803 and n18314_not n18321 ; n18995
g18804 and n18323_not n18995 ; n18996
g18805 and asqrt[9] n18996 ; n18997
g18806 nor n18314 n18323 ; n18998
g18807 and asqrt[9] n18998 ; n18999
g18808 nor n18321 n18999 ; n19000
g18809 nor n18997 n19000 ; n19001
g18810 nor asqrt[58] n18982 ; n19002
g18811 and n18992_not n19002 ; n19003
g18812 nor n19001 n19003 ; n19004
g18813 nor n18994 n19004 ; n19005
g18814 and asqrt[59] n19005_not ; n19006
g18815 and n18333 n18335_not ; n19007
g18816 and n18326_not n19007 ; n19008
g18817 and asqrt[9] n19008 ; n19009
g18818 nor n18326 n18335 ; n19010
g18819 and asqrt[9] n19010 ; n19011
g18820 nor n18333 n19011 ; n19012
g18821 nor n19009 n19012 ; n19013
g18822 nor asqrt[59] n18994 ; n19014
g18823 and n19004_not n19014 ; n19015
g18824 nor n19013 n19015 ; n19016
g18825 nor n19006 n19016 ; n19017
g18826 and asqrt[60] n19017_not ; n19018
g18827 and n18338_not n18345 ; n19019
g18828 and n18347_not n19019 ; n19020
g18829 and asqrt[9] n19020 ; n19021
g18830 nor n18338 n18347 ; n19022
g18831 and asqrt[9] n19022 ; n19023
g18832 nor n18345 n19023 ; n19024
g18833 nor n19021 n19024 ; n19025
g18834 nor asqrt[60] n19006 ; n19026
g18835 and n19016_not n19026 ; n19027
g18836 nor n19025 n19027 ; n19028
g18837 nor n19018 n19028 ; n19029
g18838 and asqrt[61] n19029_not ; n19030
g18839 and n18357 n18359_not ; n19031
g18840 and n18350_not n19031 ; n19032
g18841 and asqrt[9] n19032 ; n19033
g18842 nor n18350 n18359 ; n19034
g18843 and asqrt[9] n19034 ; n19035
g18844 nor n18357 n19035 ; n19036
g18845 nor n19033 n19036 ; n19037
g18846 nor asqrt[61] n19018 ; n19038
g18847 and n19028_not n19038 ; n19039
g18848 nor n19037 n19039 ; n19040
g18849 nor n19030 n19040 ; n19041
g18850 and asqrt[62] n19041_not ; n19042
g18851 and n18362_not n18369 ; n19043
g18852 and n18371_not n19043 ; n19044
g18853 and asqrt[9] n19044 ; n19045
g18854 nor n18362 n18371 ; n19046
g18855 and asqrt[9] n19046 ; n19047
g18856 nor n18369 n19047 ; n19048
g18857 nor n19045 n19048 ; n19049
g18858 nor asqrt[62] n19030 ; n19050
g18859 and n19040_not n19050 ; n19051
g18860 nor n19049 n19051 ; n19052
g18861 nor n19042 n19052 ; n19053
g18862 and n18381 n18383_not ; n19054
g18863 and n18374_not n19054 ; n19055
g18864 and asqrt[9] n19055 ; n19056
g18865 nor n18374 n18383 ; n19057
g18866 and asqrt[9] n19057 ; n19058
g18867 nor n18381 n19058 ; n19059
g18868 nor n19056 n19059 ; n19060
g18869 nor n18385 n18392 ; n19061
g18870 and asqrt[9] n19061 ; n19062
g18871 nor n18400 n19062 ; n19063
g18872 and n19060_not n19063 ; n19064
g18873 and n19053_not n19064 ; n19065
g18874 nor asqrt[63] n19065 ; n19066
g18875 and n19042_not n19060 ; n19067
g18876 and n19052_not n19067 ; n19068
g18877 and n18392_not asqrt[9] ; n19069
g18878 and n18385 n19069_not ; n19070
g18879 and asqrt[63] n19061_not ; n19071
g18880 and n19070_not n19071 ; n19072
g18881 nor n18388 n18409 ; n19073
g18882 and n18391_not n19073 ; n19074
g18883 and n18404_not n19074 ; n19075
g18884 and n18400_not n19075 ; n19076
g18885 and n18398_not n19076 ; n19077
g18886 nor n19072 n19077 ; n19078
g18887 and n19068_not n19078 ; n19079
g18888 nand n19066_not n19079 ; asqrt[8]
g18889 and a[16] asqrt[8] ; n19081
g18890 nor a[14] a[15] ; n19082
g18891 and a[16]_not n19082 ; n19083
g18892 nor n19081 n19083 ; n19084
g18893 and asqrt[9] n19084_not ; n19085
g18894 nor n18409 n19083 ; n19086
g18895 and n18404_not n19086 ; n19087
g18896 and n18400_not n19087 ; n19088
g18897 and n18398_not n19088 ; n19089
g18898 and n19081_not n19089 ; n19090
g18899 and a[16]_not asqrt[8] ; n19091
g18900 and a[17] n19091_not ; n19092
g18901 and n18414 asqrt[8] ; n19093
g18902 nor n19092 n19093 ; n19094
g18903 and n19090_not n19094 ; n19095
g18904 nor n19085 n19095 ; n19096
g18905 and asqrt[10] n19096_not ; n19097
g18906 nor asqrt[10] n19085 ; n19098
g18907 and n19095_not n19098 ; n19099
g18908 and asqrt[9] n19077_not ; n19100
g18909 and n19072_not n19100 ; n19101
g18910 and n19068_not n19101 ; n19102
g18911 and n19066_not n19102 ; n19103
g18912 nor n19093 n19103 ; n19104
g18913 and a[18] n19104_not ; n19105
g18914 nor a[18] n19103 ; n19106
g18915 and n19093_not n19106 ; n19107
g18916 nor n19105 n19107 ; n19108
g18917 nor n19099 n19108 ; n19109
g18918 nor n19097 n19109 ; n19110
g18919 and asqrt[11] n19110_not ; n19111
g18920 nor n18417 n18422 ; n19112
g18921 and n18426_not n19112 ; n19113
g18922 and asqrt[8] n19113 ; n19114
g18923 and asqrt[8] n19112 ; n19115
g18924 and n18426 n19115_not ; n19116
g18925 nor n19114 n19116 ; n19117
g18926 nor asqrt[11] n19097 ; n19118
g18927 and n19109_not n19118 ; n19119
g18928 nor n19117 n19119 ; n19120
g18929 nor n19111 n19120 ; n19121
g18930 and asqrt[12] n19121_not ; n19122
g18931 and n18431_not n18440 ; n19123
g18932 and n18429_not n19123 ; n19124
g18933 and asqrt[8] n19124 ; n19125
g18934 nor n18429 n18431 ; n19126
g18935 and asqrt[8] n19126 ; n19127
g18936 nor n18440 n19127 ; n19128
g18937 nor n19125 n19128 ; n19129
g18938 nor asqrt[12] n19111 ; n19130
g18939 and n19120_not n19130 ; n19131
g18940 nor n19129 n19131 ; n19132
g18941 nor n19122 n19132 ; n19133
g18942 and asqrt[13] n19133_not ; n19134
g18943 and n18443_not n18449 ; n19135
g18944 and n18451_not n19135 ; n19136
g18945 and asqrt[8] n19136 ; n19137
g18946 nor n18443 n18451 ; n19138
g18947 and asqrt[8] n19138 ; n19139
g18948 nor n18449 n19139 ; n19140
g18949 nor n19137 n19140 ; n19141
g18950 nor asqrt[13] n19122 ; n19142
g18951 and n19132_not n19142 ; n19143
g18952 nor n19141 n19143 ; n19144
g18953 nor n19134 n19144 ; n19145
g18954 and asqrt[14] n19145_not ; n19146
g18955 and n18461 n18463_not ; n19147
g18956 and n18454_not n19147 ; n19148
g18957 and asqrt[8] n19148 ; n19149
g18958 nor n18454 n18463 ; n19150
g18959 and asqrt[8] n19150 ; n19151
g18960 nor n18461 n19151 ; n19152
g18961 nor n19149 n19152 ; n19153
g18962 nor asqrt[14] n19134 ; n19154
g18963 and n19144_not n19154 ; n19155
g18964 nor n19153 n19155 ; n19156
g18965 nor n19146 n19156 ; n19157
g18966 and asqrt[15] n19157_not ; n19158
g18967 and n18466_not n18473 ; n19159
g18968 and n18475_not n19159 ; n19160
g18969 and asqrt[8] n19160 ; n19161
g18970 nor n18466 n18475 ; n19162
g18971 and asqrt[8] n19162 ; n19163
g18972 nor n18473 n19163 ; n19164
g18973 nor n19161 n19164 ; n19165
g18974 nor asqrt[15] n19146 ; n19166
g18975 and n19156_not n19166 ; n19167
g18976 nor n19165 n19167 ; n19168
g18977 nor n19158 n19168 ; n19169
g18978 and asqrt[16] n19169_not ; n19170
g18979 and n18485 n18487_not ; n19171
g18980 and n18478_not n19171 ; n19172
g18981 and asqrt[8] n19172 ; n19173
g18982 nor n18478 n18487 ; n19174
g18983 and asqrt[8] n19174 ; n19175
g18984 nor n18485 n19175 ; n19176
g18985 nor n19173 n19176 ; n19177
g18986 nor asqrt[16] n19158 ; n19178
g18987 and n19168_not n19178 ; n19179
g18988 nor n19177 n19179 ; n19180
g18989 nor n19170 n19180 ; n19181
g18990 and asqrt[17] n19181_not ; n19182
g18991 and n18490_not n18497 ; n19183
g18992 and n18499_not n19183 ; n19184
g18993 and asqrt[8] n19184 ; n19185
g18994 nor n18490 n18499 ; n19186
g18995 and asqrt[8] n19186 ; n19187
g18996 nor n18497 n19187 ; n19188
g18997 nor n19185 n19188 ; n19189
g18998 nor asqrt[17] n19170 ; n19190
g18999 and n19180_not n19190 ; n19191
g19000 nor n19189 n19191 ; n19192
g19001 nor n19182 n19192 ; n19193
g19002 and asqrt[18] n19193_not ; n19194
g19003 and n18509 n18511_not ; n19195
g19004 and n18502_not n19195 ; n19196
g19005 and asqrt[8] n19196 ; n19197
g19006 nor n18502 n18511 ; n19198
g19007 and asqrt[8] n19198 ; n19199
g19008 nor n18509 n19199 ; n19200
g19009 nor n19197 n19200 ; n19201
g19010 nor asqrt[18] n19182 ; n19202
g19011 and n19192_not n19202 ; n19203
g19012 nor n19201 n19203 ; n19204
g19013 nor n19194 n19204 ; n19205
g19014 and asqrt[19] n19205_not ; n19206
g19015 and n18514_not n18521 ; n19207
g19016 and n18523_not n19207 ; n19208
g19017 and asqrt[8] n19208 ; n19209
g19018 nor n18514 n18523 ; n19210
g19019 and asqrt[8] n19210 ; n19211
g19020 nor n18521 n19211 ; n19212
g19021 nor n19209 n19212 ; n19213
g19022 nor asqrt[19] n19194 ; n19214
g19023 and n19204_not n19214 ; n19215
g19024 nor n19213 n19215 ; n19216
g19025 nor n19206 n19216 ; n19217
g19026 and asqrt[20] n19217_not ; n19218
g19027 and n18533 n18535_not ; n19219
g19028 and n18526_not n19219 ; n19220
g19029 and asqrt[8] n19220 ; n19221
g19030 nor n18526 n18535 ; n19222
g19031 and asqrt[8] n19222 ; n19223
g19032 nor n18533 n19223 ; n19224
g19033 nor n19221 n19224 ; n19225
g19034 nor asqrt[20] n19206 ; n19226
g19035 and n19216_not n19226 ; n19227
g19036 nor n19225 n19227 ; n19228
g19037 nor n19218 n19228 ; n19229
g19038 and asqrt[21] n19229_not ; n19230
g19039 and n18538_not n18545 ; n19231
g19040 and n18547_not n19231 ; n19232
g19041 and asqrt[8] n19232 ; n19233
g19042 nor n18538 n18547 ; n19234
g19043 and asqrt[8] n19234 ; n19235
g19044 nor n18545 n19235 ; n19236
g19045 nor n19233 n19236 ; n19237
g19046 nor asqrt[21] n19218 ; n19238
g19047 and n19228_not n19238 ; n19239
g19048 nor n19237 n19239 ; n19240
g19049 nor n19230 n19240 ; n19241
g19050 and asqrt[22] n19241_not ; n19242
g19051 and n18557 n18559_not ; n19243
g19052 and n18550_not n19243 ; n19244
g19053 and asqrt[8] n19244 ; n19245
g19054 nor n18550 n18559 ; n19246
g19055 and asqrt[8] n19246 ; n19247
g19056 nor n18557 n19247 ; n19248
g19057 nor n19245 n19248 ; n19249
g19058 nor asqrt[22] n19230 ; n19250
g19059 and n19240_not n19250 ; n19251
g19060 nor n19249 n19251 ; n19252
g19061 nor n19242 n19252 ; n19253
g19062 and asqrt[23] n19253_not ; n19254
g19063 and n18562_not n18569 ; n19255
g19064 and n18571_not n19255 ; n19256
g19065 and asqrt[8] n19256 ; n19257
g19066 nor n18562 n18571 ; n19258
g19067 and asqrt[8] n19258 ; n19259
g19068 nor n18569 n19259 ; n19260
g19069 nor n19257 n19260 ; n19261
g19070 nor asqrt[23] n19242 ; n19262
g19071 and n19252_not n19262 ; n19263
g19072 nor n19261 n19263 ; n19264
g19073 nor n19254 n19264 ; n19265
g19074 and asqrt[24] n19265_not ; n19266
g19075 and n18581 n18583_not ; n19267
g19076 and n18574_not n19267 ; n19268
g19077 and asqrt[8] n19268 ; n19269
g19078 nor n18574 n18583 ; n19270
g19079 and asqrt[8] n19270 ; n19271
g19080 nor n18581 n19271 ; n19272
g19081 nor n19269 n19272 ; n19273
g19082 nor asqrt[24] n19254 ; n19274
g19083 and n19264_not n19274 ; n19275
g19084 nor n19273 n19275 ; n19276
g19085 nor n19266 n19276 ; n19277
g19086 and asqrt[25] n19277_not ; n19278
g19087 and n18586_not n18593 ; n19279
g19088 and n18595_not n19279 ; n19280
g19089 and asqrt[8] n19280 ; n19281
g19090 nor n18586 n18595 ; n19282
g19091 and asqrt[8] n19282 ; n19283
g19092 nor n18593 n19283 ; n19284
g19093 nor n19281 n19284 ; n19285
g19094 nor asqrt[25] n19266 ; n19286
g19095 and n19276_not n19286 ; n19287
g19096 nor n19285 n19287 ; n19288
g19097 nor n19278 n19288 ; n19289
g19098 and asqrt[26] n19289_not ; n19290
g19099 and n18605 n18607_not ; n19291
g19100 and n18598_not n19291 ; n19292
g19101 and asqrt[8] n19292 ; n19293
g19102 nor n18598 n18607 ; n19294
g19103 and asqrt[8] n19294 ; n19295
g19104 nor n18605 n19295 ; n19296
g19105 nor n19293 n19296 ; n19297
g19106 nor asqrt[26] n19278 ; n19298
g19107 and n19288_not n19298 ; n19299
g19108 nor n19297 n19299 ; n19300
g19109 nor n19290 n19300 ; n19301
g19110 and asqrt[27] n19301_not ; n19302
g19111 and n18610_not n18617 ; n19303
g19112 and n18619_not n19303 ; n19304
g19113 and asqrt[8] n19304 ; n19305
g19114 nor n18610 n18619 ; n19306
g19115 and asqrt[8] n19306 ; n19307
g19116 nor n18617 n19307 ; n19308
g19117 nor n19305 n19308 ; n19309
g19118 nor asqrt[27] n19290 ; n19310
g19119 and n19300_not n19310 ; n19311
g19120 nor n19309 n19311 ; n19312
g19121 nor n19302 n19312 ; n19313
g19122 and asqrt[28] n19313_not ; n19314
g19123 and n18629 n18631_not ; n19315
g19124 and n18622_not n19315 ; n19316
g19125 and asqrt[8] n19316 ; n19317
g19126 nor n18622 n18631 ; n19318
g19127 and asqrt[8] n19318 ; n19319
g19128 nor n18629 n19319 ; n19320
g19129 nor n19317 n19320 ; n19321
g19130 nor asqrt[28] n19302 ; n19322
g19131 and n19312_not n19322 ; n19323
g19132 nor n19321 n19323 ; n19324
g19133 nor n19314 n19324 ; n19325
g19134 and asqrt[29] n19325_not ; n19326
g19135 and n18634_not n18641 ; n19327
g19136 and n18643_not n19327 ; n19328
g19137 and asqrt[8] n19328 ; n19329
g19138 nor n18634 n18643 ; n19330
g19139 and asqrt[8] n19330 ; n19331
g19140 nor n18641 n19331 ; n19332
g19141 nor n19329 n19332 ; n19333
g19142 nor asqrt[29] n19314 ; n19334
g19143 and n19324_not n19334 ; n19335
g19144 nor n19333 n19335 ; n19336
g19145 nor n19326 n19336 ; n19337
g19146 and asqrt[30] n19337_not ; n19338
g19147 and n18653 n18655_not ; n19339
g19148 and n18646_not n19339 ; n19340
g19149 and asqrt[8] n19340 ; n19341
g19150 nor n18646 n18655 ; n19342
g19151 and asqrt[8] n19342 ; n19343
g19152 nor n18653 n19343 ; n19344
g19153 nor n19341 n19344 ; n19345
g19154 nor asqrt[30] n19326 ; n19346
g19155 and n19336_not n19346 ; n19347
g19156 nor n19345 n19347 ; n19348
g19157 nor n19338 n19348 ; n19349
g19158 and asqrt[31] n19349_not ; n19350
g19159 and n18658_not n18665 ; n19351
g19160 and n18667_not n19351 ; n19352
g19161 and asqrt[8] n19352 ; n19353
g19162 nor n18658 n18667 ; n19354
g19163 and asqrt[8] n19354 ; n19355
g19164 nor n18665 n19355 ; n19356
g19165 nor n19353 n19356 ; n19357
g19166 nor asqrt[31] n19338 ; n19358
g19167 and n19348_not n19358 ; n19359
g19168 nor n19357 n19359 ; n19360
g19169 nor n19350 n19360 ; n19361
g19170 and asqrt[32] n19361_not ; n19362
g19171 and n18677 n18679_not ; n19363
g19172 and n18670_not n19363 ; n19364
g19173 and asqrt[8] n19364 ; n19365
g19174 nor n18670 n18679 ; n19366
g19175 and asqrt[8] n19366 ; n19367
g19176 nor n18677 n19367 ; n19368
g19177 nor n19365 n19368 ; n19369
g19178 nor asqrt[32] n19350 ; n19370
g19179 and n19360_not n19370 ; n19371
g19180 nor n19369 n19371 ; n19372
g19181 nor n19362 n19372 ; n19373
g19182 and asqrt[33] n19373_not ; n19374
g19183 and n18682_not n18689 ; n19375
g19184 and n18691_not n19375 ; n19376
g19185 and asqrt[8] n19376 ; n19377
g19186 nor n18682 n18691 ; n19378
g19187 and asqrt[8] n19378 ; n19379
g19188 nor n18689 n19379 ; n19380
g19189 nor n19377 n19380 ; n19381
g19190 nor asqrt[33] n19362 ; n19382
g19191 and n19372_not n19382 ; n19383
g19192 nor n19381 n19383 ; n19384
g19193 nor n19374 n19384 ; n19385
g19194 and asqrt[34] n19385_not ; n19386
g19195 and n18701 n18703_not ; n19387
g19196 and n18694_not n19387 ; n19388
g19197 and asqrt[8] n19388 ; n19389
g19198 nor n18694 n18703 ; n19390
g19199 and asqrt[8] n19390 ; n19391
g19200 nor n18701 n19391 ; n19392
g19201 nor n19389 n19392 ; n19393
g19202 nor asqrt[34] n19374 ; n19394
g19203 and n19384_not n19394 ; n19395
g19204 nor n19393 n19395 ; n19396
g19205 nor n19386 n19396 ; n19397
g19206 and asqrt[35] n19397_not ; n19398
g19207 and n18706_not n18713 ; n19399
g19208 and n18715_not n19399 ; n19400
g19209 and asqrt[8] n19400 ; n19401
g19210 nor n18706 n18715 ; n19402
g19211 and asqrt[8] n19402 ; n19403
g19212 nor n18713 n19403 ; n19404
g19213 nor n19401 n19404 ; n19405
g19214 nor asqrt[35] n19386 ; n19406
g19215 and n19396_not n19406 ; n19407
g19216 nor n19405 n19407 ; n19408
g19217 nor n19398 n19408 ; n19409
g19218 and asqrt[36] n19409_not ; n19410
g19219 and n18725 n18727_not ; n19411
g19220 and n18718_not n19411 ; n19412
g19221 and asqrt[8] n19412 ; n19413
g19222 nor n18718 n18727 ; n19414
g19223 and asqrt[8] n19414 ; n19415
g19224 nor n18725 n19415 ; n19416
g19225 nor n19413 n19416 ; n19417
g19226 nor asqrt[36] n19398 ; n19418
g19227 and n19408_not n19418 ; n19419
g19228 nor n19417 n19419 ; n19420
g19229 nor n19410 n19420 ; n19421
g19230 and asqrt[37] n19421_not ; n19422
g19231 and n18730_not n18737 ; n19423
g19232 and n18739_not n19423 ; n19424
g19233 and asqrt[8] n19424 ; n19425
g19234 nor n18730 n18739 ; n19426
g19235 and asqrt[8] n19426 ; n19427
g19236 nor n18737 n19427 ; n19428
g19237 nor n19425 n19428 ; n19429
g19238 nor asqrt[37] n19410 ; n19430
g19239 and n19420_not n19430 ; n19431
g19240 nor n19429 n19431 ; n19432
g19241 nor n19422 n19432 ; n19433
g19242 and asqrt[38] n19433_not ; n19434
g19243 and n18749 n18751_not ; n19435
g19244 and n18742_not n19435 ; n19436
g19245 and asqrt[8] n19436 ; n19437
g19246 nor n18742 n18751 ; n19438
g19247 and asqrt[8] n19438 ; n19439
g19248 nor n18749 n19439 ; n19440
g19249 nor n19437 n19440 ; n19441
g19250 nor asqrt[38] n19422 ; n19442
g19251 and n19432_not n19442 ; n19443
g19252 nor n19441 n19443 ; n19444
g19253 nor n19434 n19444 ; n19445
g19254 and asqrt[39] n19445_not ; n19446
g19255 and n18754_not n18761 ; n19447
g19256 and n18763_not n19447 ; n19448
g19257 and asqrt[8] n19448 ; n19449
g19258 nor n18754 n18763 ; n19450
g19259 and asqrt[8] n19450 ; n19451
g19260 nor n18761 n19451 ; n19452
g19261 nor n19449 n19452 ; n19453
g19262 nor asqrt[39] n19434 ; n19454
g19263 and n19444_not n19454 ; n19455
g19264 nor n19453 n19455 ; n19456
g19265 nor n19446 n19456 ; n19457
g19266 and asqrt[40] n19457_not ; n19458
g19267 and n18773 n18775_not ; n19459
g19268 and n18766_not n19459 ; n19460
g19269 and asqrt[8] n19460 ; n19461
g19270 nor n18766 n18775 ; n19462
g19271 and asqrt[8] n19462 ; n19463
g19272 nor n18773 n19463 ; n19464
g19273 nor n19461 n19464 ; n19465
g19274 nor asqrt[40] n19446 ; n19466
g19275 and n19456_not n19466 ; n19467
g19276 nor n19465 n19467 ; n19468
g19277 nor n19458 n19468 ; n19469
g19278 and asqrt[41] n19469_not ; n19470
g19279 and n18778_not n18785 ; n19471
g19280 and n18787_not n19471 ; n19472
g19281 and asqrt[8] n19472 ; n19473
g19282 nor n18778 n18787 ; n19474
g19283 and asqrt[8] n19474 ; n19475
g19284 nor n18785 n19475 ; n19476
g19285 nor n19473 n19476 ; n19477
g19286 nor asqrt[41] n19458 ; n19478
g19287 and n19468_not n19478 ; n19479
g19288 nor n19477 n19479 ; n19480
g19289 nor n19470 n19480 ; n19481
g19290 and asqrt[42] n19481_not ; n19482
g19291 and n18797 n18799_not ; n19483
g19292 and n18790_not n19483 ; n19484
g19293 and asqrt[8] n19484 ; n19485
g19294 nor n18790 n18799 ; n19486
g19295 and asqrt[8] n19486 ; n19487
g19296 nor n18797 n19487 ; n19488
g19297 nor n19485 n19488 ; n19489
g19298 nor asqrt[42] n19470 ; n19490
g19299 and n19480_not n19490 ; n19491
g19300 nor n19489 n19491 ; n19492
g19301 nor n19482 n19492 ; n19493
g19302 and asqrt[43] n19493_not ; n19494
g19303 and n18802_not n18809 ; n19495
g19304 and n18811_not n19495 ; n19496
g19305 and asqrt[8] n19496 ; n19497
g19306 nor n18802 n18811 ; n19498
g19307 and asqrt[8] n19498 ; n19499
g19308 nor n18809 n19499 ; n19500
g19309 nor n19497 n19500 ; n19501
g19310 nor asqrt[43] n19482 ; n19502
g19311 and n19492_not n19502 ; n19503
g19312 nor n19501 n19503 ; n19504
g19313 nor n19494 n19504 ; n19505
g19314 and asqrt[44] n19505_not ; n19506
g19315 and n18821 n18823_not ; n19507
g19316 and n18814_not n19507 ; n19508
g19317 and asqrt[8] n19508 ; n19509
g19318 nor n18814 n18823 ; n19510
g19319 and asqrt[8] n19510 ; n19511
g19320 nor n18821 n19511 ; n19512
g19321 nor n19509 n19512 ; n19513
g19322 nor asqrt[44] n19494 ; n19514
g19323 and n19504_not n19514 ; n19515
g19324 nor n19513 n19515 ; n19516
g19325 nor n19506 n19516 ; n19517
g19326 and asqrt[45] n19517_not ; n19518
g19327 and n18826_not n18833 ; n19519
g19328 and n18835_not n19519 ; n19520
g19329 and asqrt[8] n19520 ; n19521
g19330 nor n18826 n18835 ; n19522
g19331 and asqrt[8] n19522 ; n19523
g19332 nor n18833 n19523 ; n19524
g19333 nor n19521 n19524 ; n19525
g19334 nor asqrt[45] n19506 ; n19526
g19335 and n19516_not n19526 ; n19527
g19336 nor n19525 n19527 ; n19528
g19337 nor n19518 n19528 ; n19529
g19338 and asqrt[46] n19529_not ; n19530
g19339 and n18845 n18847_not ; n19531
g19340 and n18838_not n19531 ; n19532
g19341 and asqrt[8] n19532 ; n19533
g19342 nor n18838 n18847 ; n19534
g19343 and asqrt[8] n19534 ; n19535
g19344 nor n18845 n19535 ; n19536
g19345 nor n19533 n19536 ; n19537
g19346 nor asqrt[46] n19518 ; n19538
g19347 and n19528_not n19538 ; n19539
g19348 nor n19537 n19539 ; n19540
g19349 nor n19530 n19540 ; n19541
g19350 and asqrt[47] n19541_not ; n19542
g19351 and n18850_not n18857 ; n19543
g19352 and n18859_not n19543 ; n19544
g19353 and asqrt[8] n19544 ; n19545
g19354 nor n18850 n18859 ; n19546
g19355 and asqrt[8] n19546 ; n19547
g19356 nor n18857 n19547 ; n19548
g19357 nor n19545 n19548 ; n19549
g19358 nor asqrt[47] n19530 ; n19550
g19359 and n19540_not n19550 ; n19551
g19360 nor n19549 n19551 ; n19552
g19361 nor n19542 n19552 ; n19553
g19362 and asqrt[48] n19553_not ; n19554
g19363 and n18869 n18871_not ; n19555
g19364 and n18862_not n19555 ; n19556
g19365 and asqrt[8] n19556 ; n19557
g19366 nor n18862 n18871 ; n19558
g19367 and asqrt[8] n19558 ; n19559
g19368 nor n18869 n19559 ; n19560
g19369 nor n19557 n19560 ; n19561
g19370 nor asqrt[48] n19542 ; n19562
g19371 and n19552_not n19562 ; n19563
g19372 nor n19561 n19563 ; n19564
g19373 nor n19554 n19564 ; n19565
g19374 and asqrt[49] n19565_not ; n19566
g19375 and n18874_not n18881 ; n19567
g19376 and n18883_not n19567 ; n19568
g19377 and asqrt[8] n19568 ; n19569
g19378 nor n18874 n18883 ; n19570
g19379 and asqrt[8] n19570 ; n19571
g19380 nor n18881 n19571 ; n19572
g19381 nor n19569 n19572 ; n19573
g19382 nor asqrt[49] n19554 ; n19574
g19383 and n19564_not n19574 ; n19575
g19384 nor n19573 n19575 ; n19576
g19385 nor n19566 n19576 ; n19577
g19386 and asqrt[50] n19577_not ; n19578
g19387 and n18893 n18895_not ; n19579
g19388 and n18886_not n19579 ; n19580
g19389 and asqrt[8] n19580 ; n19581
g19390 nor n18886 n18895 ; n19582
g19391 and asqrt[8] n19582 ; n19583
g19392 nor n18893 n19583 ; n19584
g19393 nor n19581 n19584 ; n19585
g19394 nor asqrt[50] n19566 ; n19586
g19395 and n19576_not n19586 ; n19587
g19396 nor n19585 n19587 ; n19588
g19397 nor n19578 n19588 ; n19589
g19398 and asqrt[51] n19589_not ; n19590
g19399 and n18898_not n18905 ; n19591
g19400 and n18907_not n19591 ; n19592
g19401 and asqrt[8] n19592 ; n19593
g19402 nor n18898 n18907 ; n19594
g19403 and asqrt[8] n19594 ; n19595
g19404 nor n18905 n19595 ; n19596
g19405 nor n19593 n19596 ; n19597
g19406 nor asqrt[51] n19578 ; n19598
g19407 and n19588_not n19598 ; n19599
g19408 nor n19597 n19599 ; n19600
g19409 nor n19590 n19600 ; n19601
g19410 and asqrt[52] n19601_not ; n19602
g19411 and n18917 n18919_not ; n19603
g19412 and n18910_not n19603 ; n19604
g19413 and asqrt[8] n19604 ; n19605
g19414 nor n18910 n18919 ; n19606
g19415 and asqrt[8] n19606 ; n19607
g19416 nor n18917 n19607 ; n19608
g19417 nor n19605 n19608 ; n19609
g19418 nor asqrt[52] n19590 ; n19610
g19419 and n19600_not n19610 ; n19611
g19420 nor n19609 n19611 ; n19612
g19421 nor n19602 n19612 ; n19613
g19422 and asqrt[53] n19613_not ; n19614
g19423 and n18922_not n18929 ; n19615
g19424 and n18931_not n19615 ; n19616
g19425 and asqrt[8] n19616 ; n19617
g19426 nor n18922 n18931 ; n19618
g19427 and asqrt[8] n19618 ; n19619
g19428 nor n18929 n19619 ; n19620
g19429 nor n19617 n19620 ; n19621
g19430 nor asqrt[53] n19602 ; n19622
g19431 and n19612_not n19622 ; n19623
g19432 nor n19621 n19623 ; n19624
g19433 nor n19614 n19624 ; n19625
g19434 and asqrt[54] n19625_not ; n19626
g19435 and n18941 n18943_not ; n19627
g19436 and n18934_not n19627 ; n19628
g19437 and asqrt[8] n19628 ; n19629
g19438 nor n18934 n18943 ; n19630
g19439 and asqrt[8] n19630 ; n19631
g19440 nor n18941 n19631 ; n19632
g19441 nor n19629 n19632 ; n19633
g19442 nor asqrt[54] n19614 ; n19634
g19443 and n19624_not n19634 ; n19635
g19444 nor n19633 n19635 ; n19636
g19445 nor n19626 n19636 ; n19637
g19446 and asqrt[55] n19637_not ; n19638
g19447 and n18946_not n18953 ; n19639
g19448 and n18955_not n19639 ; n19640
g19449 and asqrt[8] n19640 ; n19641
g19450 nor n18946 n18955 ; n19642
g19451 and asqrt[8] n19642 ; n19643
g19452 nor n18953 n19643 ; n19644
g19453 nor n19641 n19644 ; n19645
g19454 nor asqrt[55] n19626 ; n19646
g19455 and n19636_not n19646 ; n19647
g19456 nor n19645 n19647 ; n19648
g19457 nor n19638 n19648 ; n19649
g19458 and asqrt[56] n19649_not ; n19650
g19459 and n18965 n18967_not ; n19651
g19460 and n18958_not n19651 ; n19652
g19461 and asqrt[8] n19652 ; n19653
g19462 nor n18958 n18967 ; n19654
g19463 and asqrt[8] n19654 ; n19655
g19464 nor n18965 n19655 ; n19656
g19465 nor n19653 n19656 ; n19657
g19466 nor asqrt[56] n19638 ; n19658
g19467 and n19648_not n19658 ; n19659
g19468 nor n19657 n19659 ; n19660
g19469 nor n19650 n19660 ; n19661
g19470 and asqrt[57] n19661_not ; n19662
g19471 nor asqrt[57] n19650 ; n19663
g19472 and n19660_not n19663 ; n19664
g19473 and n18970_not n18979 ; n19665
g19474 and n18972_not n19665 ; n19666
g19475 and asqrt[8] n19666 ; n19667
g19476 nor n18970 n18972 ; n19668
g19477 and asqrt[8] n19668 ; n19669
g19478 nor n18979 n19669 ; n19670
g19479 nor n19667 n19670 ; n19671
g19480 nor n19664 n19671 ; n19672
g19481 nor n19662 n19672 ; n19673
g19482 and asqrt[58] n19673_not ; n19674
g19483 and n18989 n18991_not ; n19675
g19484 and n18982_not n19675 ; n19676
g19485 and asqrt[8] n19676 ; n19677
g19486 nor n18982 n18991 ; n19678
g19487 and asqrt[8] n19678 ; n19679
g19488 nor n18989 n19679 ; n19680
g19489 nor n19677 n19680 ; n19681
g19490 nor asqrt[58] n19662 ; n19682
g19491 and n19672_not n19682 ; n19683
g19492 nor n19681 n19683 ; n19684
g19493 nor n19674 n19684 ; n19685
g19494 and asqrt[59] n19685_not ; n19686
g19495 and n18994_not n19001 ; n19687
g19496 and n19003_not n19687 ; n19688
g19497 and asqrt[8] n19688 ; n19689
g19498 nor n18994 n19003 ; n19690
g19499 and asqrt[8] n19690 ; n19691
g19500 nor n19001 n19691 ; n19692
g19501 nor n19689 n19692 ; n19693
g19502 nor asqrt[59] n19674 ; n19694
g19503 and n19684_not n19694 ; n19695
g19504 nor n19693 n19695 ; n19696
g19505 nor n19686 n19696 ; n19697
g19506 and asqrt[60] n19697_not ; n19698
g19507 and n19013 n19015_not ; n19699
g19508 and n19006_not n19699 ; n19700
g19509 and asqrt[8] n19700 ; n19701
g19510 nor n19006 n19015 ; n19702
g19511 and asqrt[8] n19702 ; n19703
g19512 nor n19013 n19703 ; n19704
g19513 nor n19701 n19704 ; n19705
g19514 nor asqrt[60] n19686 ; n19706
g19515 and n19696_not n19706 ; n19707
g19516 nor n19705 n19707 ; n19708
g19517 nor n19698 n19708 ; n19709
g19518 and asqrt[61] n19709_not ; n19710
g19519 and n19018_not n19025 ; n19711
g19520 and n19027_not n19711 ; n19712
g19521 and asqrt[8] n19712 ; n19713
g19522 nor n19018 n19027 ; n19714
g19523 and asqrt[8] n19714 ; n19715
g19524 nor n19025 n19715 ; n19716
g19525 nor n19713 n19716 ; n19717
g19526 nor asqrt[61] n19698 ; n19718
g19527 and n19708_not n19718 ; n19719
g19528 nor n19717 n19719 ; n19720
g19529 nor n19710 n19720 ; n19721
g19530 and asqrt[62] n19721_not ; n19722
g19531 and n19037 n19039_not ; n19723
g19532 and n19030_not n19723 ; n19724
g19533 and asqrt[8] n19724 ; n19725
g19534 nor n19030 n19039 ; n19726
g19535 and asqrt[8] n19726 ; n19727
g19536 nor n19037 n19727 ; n19728
g19537 nor n19725 n19728 ; n19729
g19538 nor asqrt[62] n19710 ; n19730
g19539 and n19720_not n19730 ; n19731
g19540 nor n19729 n19731 ; n19732
g19541 nor n19722 n19732 ; n19733
g19542 and n19042_not n19049 ; n19734
g19543 and n19051_not n19734 ; n19735
g19544 and asqrt[8] n19735 ; n19736
g19545 nor n19042 n19051 ; n19737
g19546 and asqrt[8] n19737 ; n19738
g19547 nor n19049 n19738 ; n19739
g19548 nor n19736 n19739 ; n19740
g19549 nor n19053 n19060 ; n19741
g19550 and asqrt[8] n19741 ; n19742
g19551 nor n19068 n19742 ; n19743
g19552 and n19740_not n19743 ; n19744
g19553 and n19733_not n19744 ; n19745
g19554 nor asqrt[63] n19745 ; n19746
g19555 and n19722_not n19740 ; n19747
g19556 and n19732_not n19747 ; n19748
g19557 and n19060_not asqrt[8] ; n19749
g19558 and n19053 n19749_not ; n19750
g19559 and asqrt[63] n19741_not ; n19751
g19560 and n19750_not n19751 ; n19752
g19561 nor n19056 n19077 ; n19753
g19562 and n19059_not n19753 ; n19754
g19563 and n19072_not n19754 ; n19755
g19564 and n19068_not n19755 ; n19756
g19565 and n19066_not n19756 ; n19757
g19566 nor n19752 n19757 ; n19758
g19567 and n19748_not n19758 ; n19759
g19568 nand n19746_not n19759 ; asqrt[7]
g19569 and a[14] asqrt[7] ; n19761
g19570 nor a[12] a[13] ; n19762
g19571 and a[14]_not n19762 ; n19763
g19572 nor n19761 n19763 ; n19764
g19573 and asqrt[8] n19764_not ; n19765
g19574 nor n19077 n19763 ; n19766
g19575 and n19072_not n19766 ; n19767
g19576 and n19068_not n19767 ; n19768
g19577 and n19066_not n19768 ; n19769
g19578 and n19761_not n19769 ; n19770
g19579 and a[14]_not asqrt[7] ; n19771
g19580 and a[15] n19771_not ; n19772
g19581 and n19082 asqrt[7] ; n19773
g19582 nor n19772 n19773 ; n19774
g19583 and n19770_not n19774 ; n19775
g19584 nor n19765 n19775 ; n19776
g19585 and asqrt[9] n19776_not ; n19777
g19586 nor asqrt[9] n19765 ; n19778
g19587 and n19775_not n19778 ; n19779
g19588 and asqrt[8] n19757_not ; n19780
g19589 and n19752_not n19780 ; n19781
g19590 and n19748_not n19781 ; n19782
g19591 and n19746_not n19782 ; n19783
g19592 nor n19773 n19783 ; n19784
g19593 and a[16] n19784_not ; n19785
g19594 nor a[16] n19783 ; n19786
g19595 and n19773_not n19786 ; n19787
g19596 nor n19785 n19787 ; n19788
g19597 nor n19779 n19788 ; n19789
g19598 nor n19777 n19789 ; n19790
g19599 and asqrt[10] n19790_not ; n19791
g19600 nor n19085 n19090 ; n19792
g19601 and n19094_not n19792 ; n19793
g19602 and asqrt[7] n19793 ; n19794
g19603 and asqrt[7] n19792 ; n19795
g19604 and n19094 n19795_not ; n19796
g19605 nor n19794 n19796 ; n19797
g19606 nor asqrt[10] n19777 ; n19798
g19607 and n19789_not n19798 ; n19799
g19608 nor n19797 n19799 ; n19800
g19609 nor n19791 n19800 ; n19801
g19610 and asqrt[11] n19801_not ; n19802
g19611 and n19099_not n19108 ; n19803
g19612 and n19097_not n19803 ; n19804
g19613 and asqrt[7] n19804 ; n19805
g19614 nor n19097 n19099 ; n19806
g19615 and asqrt[7] n19806 ; n19807
g19616 nor n19108 n19807 ; n19808
g19617 nor n19805 n19808 ; n19809
g19618 nor asqrt[11] n19791 ; n19810
g19619 and n19800_not n19810 ; n19811
g19620 nor n19809 n19811 ; n19812
g19621 nor n19802 n19812 ; n19813
g19622 and asqrt[12] n19813_not ; n19814
g19623 and n19111_not n19117 ; n19815
g19624 and n19119_not n19815 ; n19816
g19625 and asqrt[7] n19816 ; n19817
g19626 nor n19111 n19119 ; n19818
g19627 and asqrt[7] n19818 ; n19819
g19628 nor n19117 n19819 ; n19820
g19629 nor n19817 n19820 ; n19821
g19630 nor asqrt[12] n19802 ; n19822
g19631 and n19812_not n19822 ; n19823
g19632 nor n19821 n19823 ; n19824
g19633 nor n19814 n19824 ; n19825
g19634 and asqrt[13] n19825_not ; n19826
g19635 and n19129 n19131_not ; n19827
g19636 and n19122_not n19827 ; n19828
g19637 and asqrt[7] n19828 ; n19829
g19638 nor n19122 n19131 ; n19830
g19639 and asqrt[7] n19830 ; n19831
g19640 nor n19129 n19831 ; n19832
g19641 nor n19829 n19832 ; n19833
g19642 nor asqrt[13] n19814 ; n19834
g19643 and n19824_not n19834 ; n19835
g19644 nor n19833 n19835 ; n19836
g19645 nor n19826 n19836 ; n19837
g19646 and asqrt[14] n19837_not ; n19838
g19647 and n19134_not n19141 ; n19839
g19648 and n19143_not n19839 ; n19840
g19649 and asqrt[7] n19840 ; n19841
g19650 nor n19134 n19143 ; n19842
g19651 and asqrt[7] n19842 ; n19843
g19652 nor n19141 n19843 ; n19844
g19653 nor n19841 n19844 ; n19845
g19654 nor asqrt[14] n19826 ; n19846
g19655 and n19836_not n19846 ; n19847
g19656 nor n19845 n19847 ; n19848
g19657 nor n19838 n19848 ; n19849
g19658 and asqrt[15] n19849_not ; n19850
g19659 and n19153 n19155_not ; n19851
g19660 and n19146_not n19851 ; n19852
g19661 and asqrt[7] n19852 ; n19853
g19662 nor n19146 n19155 ; n19854
g19663 and asqrt[7] n19854 ; n19855
g19664 nor n19153 n19855 ; n19856
g19665 nor n19853 n19856 ; n19857
g19666 nor asqrt[15] n19838 ; n19858
g19667 and n19848_not n19858 ; n19859
g19668 nor n19857 n19859 ; n19860
g19669 nor n19850 n19860 ; n19861
g19670 and asqrt[16] n19861_not ; n19862
g19671 and n19158_not n19165 ; n19863
g19672 and n19167_not n19863 ; n19864
g19673 and asqrt[7] n19864 ; n19865
g19674 nor n19158 n19167 ; n19866
g19675 and asqrt[7] n19866 ; n19867
g19676 nor n19165 n19867 ; n19868
g19677 nor n19865 n19868 ; n19869
g19678 nor asqrt[16] n19850 ; n19870
g19679 and n19860_not n19870 ; n19871
g19680 nor n19869 n19871 ; n19872
g19681 nor n19862 n19872 ; n19873
g19682 and asqrt[17] n19873_not ; n19874
g19683 and n19177 n19179_not ; n19875
g19684 and n19170_not n19875 ; n19876
g19685 and asqrt[7] n19876 ; n19877
g19686 nor n19170 n19179 ; n19878
g19687 and asqrt[7] n19878 ; n19879
g19688 nor n19177 n19879 ; n19880
g19689 nor n19877 n19880 ; n19881
g19690 nor asqrt[17] n19862 ; n19882
g19691 and n19872_not n19882 ; n19883
g19692 nor n19881 n19883 ; n19884
g19693 nor n19874 n19884 ; n19885
g19694 and asqrt[18] n19885_not ; n19886
g19695 and n19182_not n19189 ; n19887
g19696 and n19191_not n19887 ; n19888
g19697 and asqrt[7] n19888 ; n19889
g19698 nor n19182 n19191 ; n19890
g19699 and asqrt[7] n19890 ; n19891
g19700 nor n19189 n19891 ; n19892
g19701 nor n19889 n19892 ; n19893
g19702 nor asqrt[18] n19874 ; n19894
g19703 and n19884_not n19894 ; n19895
g19704 nor n19893 n19895 ; n19896
g19705 nor n19886 n19896 ; n19897
g19706 and asqrt[19] n19897_not ; n19898
g19707 and n19201 n19203_not ; n19899
g19708 and n19194_not n19899 ; n19900
g19709 and asqrt[7] n19900 ; n19901
g19710 nor n19194 n19203 ; n19902
g19711 and asqrt[7] n19902 ; n19903
g19712 nor n19201 n19903 ; n19904
g19713 nor n19901 n19904 ; n19905
g19714 nor asqrt[19] n19886 ; n19906
g19715 and n19896_not n19906 ; n19907
g19716 nor n19905 n19907 ; n19908
g19717 nor n19898 n19908 ; n19909
g19718 and asqrt[20] n19909_not ; n19910
g19719 and n19206_not n19213 ; n19911
g19720 and n19215_not n19911 ; n19912
g19721 and asqrt[7] n19912 ; n19913
g19722 nor n19206 n19215 ; n19914
g19723 and asqrt[7] n19914 ; n19915
g19724 nor n19213 n19915 ; n19916
g19725 nor n19913 n19916 ; n19917
g19726 nor asqrt[20] n19898 ; n19918
g19727 and n19908_not n19918 ; n19919
g19728 nor n19917 n19919 ; n19920
g19729 nor n19910 n19920 ; n19921
g19730 and asqrt[21] n19921_not ; n19922
g19731 and n19225 n19227_not ; n19923
g19732 and n19218_not n19923 ; n19924
g19733 and asqrt[7] n19924 ; n19925
g19734 nor n19218 n19227 ; n19926
g19735 and asqrt[7] n19926 ; n19927
g19736 nor n19225 n19927 ; n19928
g19737 nor n19925 n19928 ; n19929
g19738 nor asqrt[21] n19910 ; n19930
g19739 and n19920_not n19930 ; n19931
g19740 nor n19929 n19931 ; n19932
g19741 nor n19922 n19932 ; n19933
g19742 and asqrt[22] n19933_not ; n19934
g19743 and n19230_not n19237 ; n19935
g19744 and n19239_not n19935 ; n19936
g19745 and asqrt[7] n19936 ; n19937
g19746 nor n19230 n19239 ; n19938
g19747 and asqrt[7] n19938 ; n19939
g19748 nor n19237 n19939 ; n19940
g19749 nor n19937 n19940 ; n19941
g19750 nor asqrt[22] n19922 ; n19942
g19751 and n19932_not n19942 ; n19943
g19752 nor n19941 n19943 ; n19944
g19753 nor n19934 n19944 ; n19945
g19754 and asqrt[23] n19945_not ; n19946
g19755 and n19249 n19251_not ; n19947
g19756 and n19242_not n19947 ; n19948
g19757 and asqrt[7] n19948 ; n19949
g19758 nor n19242 n19251 ; n19950
g19759 and asqrt[7] n19950 ; n19951
g19760 nor n19249 n19951 ; n19952
g19761 nor n19949 n19952 ; n19953
g19762 nor asqrt[23] n19934 ; n19954
g19763 and n19944_not n19954 ; n19955
g19764 nor n19953 n19955 ; n19956
g19765 nor n19946 n19956 ; n19957
g19766 and asqrt[24] n19957_not ; n19958
g19767 and n19254_not n19261 ; n19959
g19768 and n19263_not n19959 ; n19960
g19769 and asqrt[7] n19960 ; n19961
g19770 nor n19254 n19263 ; n19962
g19771 and asqrt[7] n19962 ; n19963
g19772 nor n19261 n19963 ; n19964
g19773 nor n19961 n19964 ; n19965
g19774 nor asqrt[24] n19946 ; n19966
g19775 and n19956_not n19966 ; n19967
g19776 nor n19965 n19967 ; n19968
g19777 nor n19958 n19968 ; n19969
g19778 and asqrt[25] n19969_not ; n19970
g19779 and n19273 n19275_not ; n19971
g19780 and n19266_not n19971 ; n19972
g19781 and asqrt[7] n19972 ; n19973
g19782 nor n19266 n19275 ; n19974
g19783 and asqrt[7] n19974 ; n19975
g19784 nor n19273 n19975 ; n19976
g19785 nor n19973 n19976 ; n19977
g19786 nor asqrt[25] n19958 ; n19978
g19787 and n19968_not n19978 ; n19979
g19788 nor n19977 n19979 ; n19980
g19789 nor n19970 n19980 ; n19981
g19790 and asqrt[26] n19981_not ; n19982
g19791 and n19278_not n19285 ; n19983
g19792 and n19287_not n19983 ; n19984
g19793 and asqrt[7] n19984 ; n19985
g19794 nor n19278 n19287 ; n19986
g19795 and asqrt[7] n19986 ; n19987
g19796 nor n19285 n19987 ; n19988
g19797 nor n19985 n19988 ; n19989
g19798 nor asqrt[26] n19970 ; n19990
g19799 and n19980_not n19990 ; n19991
g19800 nor n19989 n19991 ; n19992
g19801 nor n19982 n19992 ; n19993
g19802 and asqrt[27] n19993_not ; n19994
g19803 and n19297 n19299_not ; n19995
g19804 and n19290_not n19995 ; n19996
g19805 and asqrt[7] n19996 ; n19997
g19806 nor n19290 n19299 ; n19998
g19807 and asqrt[7] n19998 ; n19999
g19808 nor n19297 n19999 ; n20000
g19809 nor n19997 n20000 ; n20001
g19810 nor asqrt[27] n19982 ; n20002
g19811 and n19992_not n20002 ; n20003
g19812 nor n20001 n20003 ; n20004
g19813 nor n19994 n20004 ; n20005
g19814 and asqrt[28] n20005_not ; n20006
g19815 and n19302_not n19309 ; n20007
g19816 and n19311_not n20007 ; n20008
g19817 and asqrt[7] n20008 ; n20009
g19818 nor n19302 n19311 ; n20010
g19819 and asqrt[7] n20010 ; n20011
g19820 nor n19309 n20011 ; n20012
g19821 nor n20009 n20012 ; n20013
g19822 nor asqrt[28] n19994 ; n20014
g19823 and n20004_not n20014 ; n20015
g19824 nor n20013 n20015 ; n20016
g19825 nor n20006 n20016 ; n20017
g19826 and asqrt[29] n20017_not ; n20018
g19827 and n19321 n19323_not ; n20019
g19828 and n19314_not n20019 ; n20020
g19829 and asqrt[7] n20020 ; n20021
g19830 nor n19314 n19323 ; n20022
g19831 and asqrt[7] n20022 ; n20023
g19832 nor n19321 n20023 ; n20024
g19833 nor n20021 n20024 ; n20025
g19834 nor asqrt[29] n20006 ; n20026
g19835 and n20016_not n20026 ; n20027
g19836 nor n20025 n20027 ; n20028
g19837 nor n20018 n20028 ; n20029
g19838 and asqrt[30] n20029_not ; n20030
g19839 and n19326_not n19333 ; n20031
g19840 and n19335_not n20031 ; n20032
g19841 and asqrt[7] n20032 ; n20033
g19842 nor n19326 n19335 ; n20034
g19843 and asqrt[7] n20034 ; n20035
g19844 nor n19333 n20035 ; n20036
g19845 nor n20033 n20036 ; n20037
g19846 nor asqrt[30] n20018 ; n20038
g19847 and n20028_not n20038 ; n20039
g19848 nor n20037 n20039 ; n20040
g19849 nor n20030 n20040 ; n20041
g19850 and asqrt[31] n20041_not ; n20042
g19851 and n19345 n19347_not ; n20043
g19852 and n19338_not n20043 ; n20044
g19853 and asqrt[7] n20044 ; n20045
g19854 nor n19338 n19347 ; n20046
g19855 and asqrt[7] n20046 ; n20047
g19856 nor n19345 n20047 ; n20048
g19857 nor n20045 n20048 ; n20049
g19858 nor asqrt[31] n20030 ; n20050
g19859 and n20040_not n20050 ; n20051
g19860 nor n20049 n20051 ; n20052
g19861 nor n20042 n20052 ; n20053
g19862 and asqrt[32] n20053_not ; n20054
g19863 and n19350_not n19357 ; n20055
g19864 and n19359_not n20055 ; n20056
g19865 and asqrt[7] n20056 ; n20057
g19866 nor n19350 n19359 ; n20058
g19867 and asqrt[7] n20058 ; n20059
g19868 nor n19357 n20059 ; n20060
g19869 nor n20057 n20060 ; n20061
g19870 nor asqrt[32] n20042 ; n20062
g19871 and n20052_not n20062 ; n20063
g19872 nor n20061 n20063 ; n20064
g19873 nor n20054 n20064 ; n20065
g19874 and asqrt[33] n20065_not ; n20066
g19875 and n19369 n19371_not ; n20067
g19876 and n19362_not n20067 ; n20068
g19877 and asqrt[7] n20068 ; n20069
g19878 nor n19362 n19371 ; n20070
g19879 and asqrt[7] n20070 ; n20071
g19880 nor n19369 n20071 ; n20072
g19881 nor n20069 n20072 ; n20073
g19882 nor asqrt[33] n20054 ; n20074
g19883 and n20064_not n20074 ; n20075
g19884 nor n20073 n20075 ; n20076
g19885 nor n20066 n20076 ; n20077
g19886 and asqrt[34] n20077_not ; n20078
g19887 and n19374_not n19381 ; n20079
g19888 and n19383_not n20079 ; n20080
g19889 and asqrt[7] n20080 ; n20081
g19890 nor n19374 n19383 ; n20082
g19891 and asqrt[7] n20082 ; n20083
g19892 nor n19381 n20083 ; n20084
g19893 nor n20081 n20084 ; n20085
g19894 nor asqrt[34] n20066 ; n20086
g19895 and n20076_not n20086 ; n20087
g19896 nor n20085 n20087 ; n20088
g19897 nor n20078 n20088 ; n20089
g19898 and asqrt[35] n20089_not ; n20090
g19899 and n19393 n19395_not ; n20091
g19900 and n19386_not n20091 ; n20092
g19901 and asqrt[7] n20092 ; n20093
g19902 nor n19386 n19395 ; n20094
g19903 and asqrt[7] n20094 ; n20095
g19904 nor n19393 n20095 ; n20096
g19905 nor n20093 n20096 ; n20097
g19906 nor asqrt[35] n20078 ; n20098
g19907 and n20088_not n20098 ; n20099
g19908 nor n20097 n20099 ; n20100
g19909 nor n20090 n20100 ; n20101
g19910 and asqrt[36] n20101_not ; n20102
g19911 and n19398_not n19405 ; n20103
g19912 and n19407_not n20103 ; n20104
g19913 and asqrt[7] n20104 ; n20105
g19914 nor n19398 n19407 ; n20106
g19915 and asqrt[7] n20106 ; n20107
g19916 nor n19405 n20107 ; n20108
g19917 nor n20105 n20108 ; n20109
g19918 nor asqrt[36] n20090 ; n20110
g19919 and n20100_not n20110 ; n20111
g19920 nor n20109 n20111 ; n20112
g19921 nor n20102 n20112 ; n20113
g19922 and asqrt[37] n20113_not ; n20114
g19923 and n19417 n19419_not ; n20115
g19924 and n19410_not n20115 ; n20116
g19925 and asqrt[7] n20116 ; n20117
g19926 nor n19410 n19419 ; n20118
g19927 and asqrt[7] n20118 ; n20119
g19928 nor n19417 n20119 ; n20120
g19929 nor n20117 n20120 ; n20121
g19930 nor asqrt[37] n20102 ; n20122
g19931 and n20112_not n20122 ; n20123
g19932 nor n20121 n20123 ; n20124
g19933 nor n20114 n20124 ; n20125
g19934 and asqrt[38] n20125_not ; n20126
g19935 and n19422_not n19429 ; n20127
g19936 and n19431_not n20127 ; n20128
g19937 and asqrt[7] n20128 ; n20129
g19938 nor n19422 n19431 ; n20130
g19939 and asqrt[7] n20130 ; n20131
g19940 nor n19429 n20131 ; n20132
g19941 nor n20129 n20132 ; n20133
g19942 nor asqrt[38] n20114 ; n20134
g19943 and n20124_not n20134 ; n20135
g19944 nor n20133 n20135 ; n20136
g19945 nor n20126 n20136 ; n20137
g19946 and asqrt[39] n20137_not ; n20138
g19947 and n19441 n19443_not ; n20139
g19948 and n19434_not n20139 ; n20140
g19949 and asqrt[7] n20140 ; n20141
g19950 nor n19434 n19443 ; n20142
g19951 and asqrt[7] n20142 ; n20143
g19952 nor n19441 n20143 ; n20144
g19953 nor n20141 n20144 ; n20145
g19954 nor asqrt[39] n20126 ; n20146
g19955 and n20136_not n20146 ; n20147
g19956 nor n20145 n20147 ; n20148
g19957 nor n20138 n20148 ; n20149
g19958 and asqrt[40] n20149_not ; n20150
g19959 and n19446_not n19453 ; n20151
g19960 and n19455_not n20151 ; n20152
g19961 and asqrt[7] n20152 ; n20153
g19962 nor n19446 n19455 ; n20154
g19963 and asqrt[7] n20154 ; n20155
g19964 nor n19453 n20155 ; n20156
g19965 nor n20153 n20156 ; n20157
g19966 nor asqrt[40] n20138 ; n20158
g19967 and n20148_not n20158 ; n20159
g19968 nor n20157 n20159 ; n20160
g19969 nor n20150 n20160 ; n20161
g19970 and asqrt[41] n20161_not ; n20162
g19971 and n19465 n19467_not ; n20163
g19972 and n19458_not n20163 ; n20164
g19973 and asqrt[7] n20164 ; n20165
g19974 nor n19458 n19467 ; n20166
g19975 and asqrt[7] n20166 ; n20167
g19976 nor n19465 n20167 ; n20168
g19977 nor n20165 n20168 ; n20169
g19978 nor asqrt[41] n20150 ; n20170
g19979 and n20160_not n20170 ; n20171
g19980 nor n20169 n20171 ; n20172
g19981 nor n20162 n20172 ; n20173
g19982 and asqrt[42] n20173_not ; n20174
g19983 and n19470_not n19477 ; n20175
g19984 and n19479_not n20175 ; n20176
g19985 and asqrt[7] n20176 ; n20177
g19986 nor n19470 n19479 ; n20178
g19987 and asqrt[7] n20178 ; n20179
g19988 nor n19477 n20179 ; n20180
g19989 nor n20177 n20180 ; n20181
g19990 nor asqrt[42] n20162 ; n20182
g19991 and n20172_not n20182 ; n20183
g19992 nor n20181 n20183 ; n20184
g19993 nor n20174 n20184 ; n20185
g19994 and asqrt[43] n20185_not ; n20186
g19995 and n19489 n19491_not ; n20187
g19996 and n19482_not n20187 ; n20188
g19997 and asqrt[7] n20188 ; n20189
g19998 nor n19482 n19491 ; n20190
g19999 and asqrt[7] n20190 ; n20191
g20000 nor n19489 n20191 ; n20192
g20001 nor n20189 n20192 ; n20193
g20002 nor asqrt[43] n20174 ; n20194
g20003 and n20184_not n20194 ; n20195
g20004 nor n20193 n20195 ; n20196
g20005 nor n20186 n20196 ; n20197
g20006 and asqrt[44] n20197_not ; n20198
g20007 and n19494_not n19501 ; n20199
g20008 and n19503_not n20199 ; n20200
g20009 and asqrt[7] n20200 ; n20201
g20010 nor n19494 n19503 ; n20202
g20011 and asqrt[7] n20202 ; n20203
g20012 nor n19501 n20203 ; n20204
g20013 nor n20201 n20204 ; n20205
g20014 nor asqrt[44] n20186 ; n20206
g20015 and n20196_not n20206 ; n20207
g20016 nor n20205 n20207 ; n20208
g20017 nor n20198 n20208 ; n20209
g20018 and asqrt[45] n20209_not ; n20210
g20019 and n19513 n19515_not ; n20211
g20020 and n19506_not n20211 ; n20212
g20021 and asqrt[7] n20212 ; n20213
g20022 nor n19506 n19515 ; n20214
g20023 and asqrt[7] n20214 ; n20215
g20024 nor n19513 n20215 ; n20216
g20025 nor n20213 n20216 ; n20217
g20026 nor asqrt[45] n20198 ; n20218
g20027 and n20208_not n20218 ; n20219
g20028 nor n20217 n20219 ; n20220
g20029 nor n20210 n20220 ; n20221
g20030 and asqrt[46] n20221_not ; n20222
g20031 and n19518_not n19525 ; n20223
g20032 and n19527_not n20223 ; n20224
g20033 and asqrt[7] n20224 ; n20225
g20034 nor n19518 n19527 ; n20226
g20035 and asqrt[7] n20226 ; n20227
g20036 nor n19525 n20227 ; n20228
g20037 nor n20225 n20228 ; n20229
g20038 nor asqrt[46] n20210 ; n20230
g20039 and n20220_not n20230 ; n20231
g20040 nor n20229 n20231 ; n20232
g20041 nor n20222 n20232 ; n20233
g20042 and asqrt[47] n20233_not ; n20234
g20043 and n19537 n19539_not ; n20235
g20044 and n19530_not n20235 ; n20236
g20045 and asqrt[7] n20236 ; n20237
g20046 nor n19530 n19539 ; n20238
g20047 and asqrt[7] n20238 ; n20239
g20048 nor n19537 n20239 ; n20240
g20049 nor n20237 n20240 ; n20241
g20050 nor asqrt[47] n20222 ; n20242
g20051 and n20232_not n20242 ; n20243
g20052 nor n20241 n20243 ; n20244
g20053 nor n20234 n20244 ; n20245
g20054 and asqrt[48] n20245_not ; n20246
g20055 and n19542_not n19549 ; n20247
g20056 and n19551_not n20247 ; n20248
g20057 and asqrt[7] n20248 ; n20249
g20058 nor n19542 n19551 ; n20250
g20059 and asqrt[7] n20250 ; n20251
g20060 nor n19549 n20251 ; n20252
g20061 nor n20249 n20252 ; n20253
g20062 nor asqrt[48] n20234 ; n20254
g20063 and n20244_not n20254 ; n20255
g20064 nor n20253 n20255 ; n20256
g20065 nor n20246 n20256 ; n20257
g20066 and asqrt[49] n20257_not ; n20258
g20067 and n19561 n19563_not ; n20259
g20068 and n19554_not n20259 ; n20260
g20069 and asqrt[7] n20260 ; n20261
g20070 nor n19554 n19563 ; n20262
g20071 and asqrt[7] n20262 ; n20263
g20072 nor n19561 n20263 ; n20264
g20073 nor n20261 n20264 ; n20265
g20074 nor asqrt[49] n20246 ; n20266
g20075 and n20256_not n20266 ; n20267
g20076 nor n20265 n20267 ; n20268
g20077 nor n20258 n20268 ; n20269
g20078 and asqrt[50] n20269_not ; n20270
g20079 and n19566_not n19573 ; n20271
g20080 and n19575_not n20271 ; n20272
g20081 and asqrt[7] n20272 ; n20273
g20082 nor n19566 n19575 ; n20274
g20083 and asqrt[7] n20274 ; n20275
g20084 nor n19573 n20275 ; n20276
g20085 nor n20273 n20276 ; n20277
g20086 nor asqrt[50] n20258 ; n20278
g20087 and n20268_not n20278 ; n20279
g20088 nor n20277 n20279 ; n20280
g20089 nor n20270 n20280 ; n20281
g20090 and asqrt[51] n20281_not ; n20282
g20091 and n19585 n19587_not ; n20283
g20092 and n19578_not n20283 ; n20284
g20093 and asqrt[7] n20284 ; n20285
g20094 nor n19578 n19587 ; n20286
g20095 and asqrt[7] n20286 ; n20287
g20096 nor n19585 n20287 ; n20288
g20097 nor n20285 n20288 ; n20289
g20098 nor asqrt[51] n20270 ; n20290
g20099 and n20280_not n20290 ; n20291
g20100 nor n20289 n20291 ; n20292
g20101 nor n20282 n20292 ; n20293
g20102 and asqrt[52] n20293_not ; n20294
g20103 and n19590_not n19597 ; n20295
g20104 and n19599_not n20295 ; n20296
g20105 and asqrt[7] n20296 ; n20297
g20106 nor n19590 n19599 ; n20298
g20107 and asqrt[7] n20298 ; n20299
g20108 nor n19597 n20299 ; n20300
g20109 nor n20297 n20300 ; n20301
g20110 nor asqrt[52] n20282 ; n20302
g20111 and n20292_not n20302 ; n20303
g20112 nor n20301 n20303 ; n20304
g20113 nor n20294 n20304 ; n20305
g20114 and asqrt[53] n20305_not ; n20306
g20115 and n19609 n19611_not ; n20307
g20116 and n19602_not n20307 ; n20308
g20117 and asqrt[7] n20308 ; n20309
g20118 nor n19602 n19611 ; n20310
g20119 and asqrt[7] n20310 ; n20311
g20120 nor n19609 n20311 ; n20312
g20121 nor n20309 n20312 ; n20313
g20122 nor asqrt[53] n20294 ; n20314
g20123 and n20304_not n20314 ; n20315
g20124 nor n20313 n20315 ; n20316
g20125 nor n20306 n20316 ; n20317
g20126 and asqrt[54] n20317_not ; n20318
g20127 and n19614_not n19621 ; n20319
g20128 and n19623_not n20319 ; n20320
g20129 and asqrt[7] n20320 ; n20321
g20130 nor n19614 n19623 ; n20322
g20131 and asqrt[7] n20322 ; n20323
g20132 nor n19621 n20323 ; n20324
g20133 nor n20321 n20324 ; n20325
g20134 nor asqrt[54] n20306 ; n20326
g20135 and n20316_not n20326 ; n20327
g20136 nor n20325 n20327 ; n20328
g20137 nor n20318 n20328 ; n20329
g20138 and asqrt[55] n20329_not ; n20330
g20139 and n19633 n19635_not ; n20331
g20140 and n19626_not n20331 ; n20332
g20141 and asqrt[7] n20332 ; n20333
g20142 nor n19626 n19635 ; n20334
g20143 and asqrt[7] n20334 ; n20335
g20144 nor n19633 n20335 ; n20336
g20145 nor n20333 n20336 ; n20337
g20146 nor asqrt[55] n20318 ; n20338
g20147 and n20328_not n20338 ; n20339
g20148 nor n20337 n20339 ; n20340
g20149 nor n20330 n20340 ; n20341
g20150 and asqrt[56] n20341_not ; n20342
g20151 and n19638_not n19645 ; n20343
g20152 and n19647_not n20343 ; n20344
g20153 and asqrt[7] n20344 ; n20345
g20154 nor n19638 n19647 ; n20346
g20155 and asqrt[7] n20346 ; n20347
g20156 nor n19645 n20347 ; n20348
g20157 nor n20345 n20348 ; n20349
g20158 nor asqrt[56] n20330 ; n20350
g20159 and n20340_not n20350 ; n20351
g20160 nor n20349 n20351 ; n20352
g20161 nor n20342 n20352 ; n20353
g20162 and asqrt[57] n20353_not ; n20354
g20163 and n19657 n19659_not ; n20355
g20164 and n19650_not n20355 ; n20356
g20165 and asqrt[7] n20356 ; n20357
g20166 nor n19650 n19659 ; n20358
g20167 and asqrt[7] n20358 ; n20359
g20168 nor n19657 n20359 ; n20360
g20169 nor n20357 n20360 ; n20361
g20170 nor asqrt[57] n20342 ; n20362
g20171 and n20352_not n20362 ; n20363
g20172 nor n20361 n20363 ; n20364
g20173 nor n20354 n20364 ; n20365
g20174 and asqrt[58] n20365_not ; n20366
g20175 nor asqrt[58] n20354 ; n20367
g20176 and n20364_not n20367 ; n20368
g20177 and n19662_not n19671 ; n20369
g20178 and n19664_not n20369 ; n20370
g20179 and asqrt[7] n20370 ; n20371
g20180 nor n19662 n19664 ; n20372
g20181 and asqrt[7] n20372 ; n20373
g20182 nor n19671 n20373 ; n20374
g20183 nor n20371 n20374 ; n20375
g20184 nor n20368 n20375 ; n20376
g20185 nor n20366 n20376 ; n20377
g20186 and asqrt[59] n20377_not ; n20378
g20187 and n19681 n19683_not ; n20379
g20188 and n19674_not n20379 ; n20380
g20189 and asqrt[7] n20380 ; n20381
g20190 nor n19674 n19683 ; n20382
g20191 and asqrt[7] n20382 ; n20383
g20192 nor n19681 n20383 ; n20384
g20193 nor n20381 n20384 ; n20385
g20194 nor asqrt[59] n20366 ; n20386
g20195 and n20376_not n20386 ; n20387
g20196 nor n20385 n20387 ; n20388
g20197 nor n20378 n20388 ; n20389
g20198 and asqrt[60] n20389_not ; n20390
g20199 and n19686_not n19693 ; n20391
g20200 and n19695_not n20391 ; n20392
g20201 and asqrt[7] n20392 ; n20393
g20202 nor n19686 n19695 ; n20394
g20203 and asqrt[7] n20394 ; n20395
g20204 nor n19693 n20395 ; n20396
g20205 nor n20393 n20396 ; n20397
g20206 nor asqrt[60] n20378 ; n20398
g20207 and n20388_not n20398 ; n20399
g20208 nor n20397 n20399 ; n20400
g20209 nor n20390 n20400 ; n20401
g20210 and asqrt[61] n20401_not ; n20402
g20211 and n19705 n19707_not ; n20403
g20212 and n19698_not n20403 ; n20404
g20213 and asqrt[7] n20404 ; n20405
g20214 nor n19698 n19707 ; n20406
g20215 and asqrt[7] n20406 ; n20407
g20216 nor n19705 n20407 ; n20408
g20217 nor n20405 n20408 ; n20409
g20218 nor asqrt[61] n20390 ; n20410
g20219 and n20400_not n20410 ; n20411
g20220 nor n20409 n20411 ; n20412
g20221 nor n20402 n20412 ; n20413
g20222 and asqrt[62] n20413_not ; n20414
g20223 and n19710_not n19717 ; n20415
g20224 and n19719_not n20415 ; n20416
g20225 and asqrt[7] n20416 ; n20417
g20226 nor n19710 n19719 ; n20418
g20227 and asqrt[7] n20418 ; n20419
g20228 nor n19717 n20419 ; n20420
g20229 nor n20417 n20420 ; n20421
g20230 nor asqrt[62] n20402 ; n20422
g20231 and n20412_not n20422 ; n20423
g20232 nor n20421 n20423 ; n20424
g20233 nor n20414 n20424 ; n20425
g20234 and n19729 n19731_not ; n20426
g20235 and n19722_not n20426 ; n20427
g20236 and asqrt[7] n20427 ; n20428
g20237 nor n19722 n19731 ; n20429
g20238 and asqrt[7] n20429 ; n20430
g20239 nor n19729 n20430 ; n20431
g20240 nor n20428 n20431 ; n20432
g20241 nor n19733 n19740 ; n20433
g20242 and asqrt[7] n20433 ; n20434
g20243 nor n19748 n20434 ; n20435
g20244 and n20432_not n20435 ; n20436
g20245 and n20425_not n20436 ; n20437
g20246 nor asqrt[63] n20437 ; n20438
g20247 and n20414_not n20432 ; n20439
g20248 and n20424_not n20439 ; n20440
g20249 and n19740_not asqrt[7] ; n20441
g20250 and n19733 n20441_not ; n20442
g20251 and asqrt[63] n20433_not ; n20443
g20252 and n20442_not n20443 ; n20444
g20253 nor n19736 n19757 ; n20445
g20254 and n19739_not n20445 ; n20446
g20255 and n19752_not n20446 ; n20447
g20256 and n19748_not n20447 ; n20448
g20257 and n19746_not n20448 ; n20449
g20258 nor n20444 n20449 ; n20450
g20259 and n20440_not n20450 ; n20451
g20260 nand n20438_not n20451 ; asqrt[6]
g20261 and a[12] asqrt[6] ; n20453
g20262 nor a[10] a[11] ; n20454
g20263 and a[12]_not n20454 ; n20455
g20264 nor n20453 n20455 ; n20456
g20265 and asqrt[7] n20456_not ; n20457
g20266 nor n19757 n20455 ; n20458
g20267 and n19752_not n20458 ; n20459
g20268 and n19748_not n20459 ; n20460
g20269 and n19746_not n20460 ; n20461
g20270 and n20453_not n20461 ; n20462
g20271 and a[12]_not asqrt[6] ; n20463
g20272 and a[13] n20463_not ; n20464
g20273 and n19762 asqrt[6] ; n20465
g20274 nor n20464 n20465 ; n20466
g20275 and n20462_not n20466 ; n20467
g20276 nor n20457 n20467 ; n20468
g20277 and asqrt[8] n20468_not ; n20469
g20278 nor asqrt[8] n20457 ; n20470
g20279 and n20467_not n20470 ; n20471
g20280 and asqrt[7] n20449_not ; n20472
g20281 and n20444_not n20472 ; n20473
g20282 and n20440_not n20473 ; n20474
g20283 and n20438_not n20474 ; n20475
g20284 nor n20465 n20475 ; n20476
g20285 and a[14] n20476_not ; n20477
g20286 nor a[14] n20475 ; n20478
g20287 and n20465_not n20478 ; n20479
g20288 nor n20477 n20479 ; n20480
g20289 nor n20471 n20480 ; n20481
g20290 nor n20469 n20481 ; n20482
g20291 and asqrt[9] n20482_not ; n20483
g20292 nor n19765 n19770 ; n20484
g20293 and n19774_not n20484 ; n20485
g20294 and asqrt[6] n20485 ; n20486
g20295 and asqrt[6] n20484 ; n20487
g20296 and n19774 n20487_not ; n20488
g20297 nor n20486 n20488 ; n20489
g20298 nor asqrt[9] n20469 ; n20490
g20299 and n20481_not n20490 ; n20491
g20300 nor n20489 n20491 ; n20492
g20301 nor n20483 n20492 ; n20493
g20302 and asqrt[10] n20493_not ; n20494
g20303 and n19779_not n19788 ; n20495
g20304 and n19777_not n20495 ; n20496
g20305 and asqrt[6] n20496 ; n20497
g20306 nor n19777 n19779 ; n20498
g20307 and asqrt[6] n20498 ; n20499
g20308 nor n19788 n20499 ; n20500
g20309 nor n20497 n20500 ; n20501
g20310 nor asqrt[10] n20483 ; n20502
g20311 and n20492_not n20502 ; n20503
g20312 nor n20501 n20503 ; n20504
g20313 nor n20494 n20504 ; n20505
g20314 and asqrt[11] n20505_not ; n20506
g20315 and n19791_not n19797 ; n20507
g20316 and n19799_not n20507 ; n20508
g20317 and asqrt[6] n20508 ; n20509
g20318 nor n19791 n19799 ; n20510
g20319 and asqrt[6] n20510 ; n20511
g20320 nor n19797 n20511 ; n20512
g20321 nor n20509 n20512 ; n20513
g20322 nor asqrt[11] n20494 ; n20514
g20323 and n20504_not n20514 ; n20515
g20324 nor n20513 n20515 ; n20516
g20325 nor n20506 n20516 ; n20517
g20326 and asqrt[12] n20517_not ; n20518
g20327 and n19809 n19811_not ; n20519
g20328 and n19802_not n20519 ; n20520
g20329 and asqrt[6] n20520 ; n20521
g20330 nor n19802 n19811 ; n20522
g20331 and asqrt[6] n20522 ; n20523
g20332 nor n19809 n20523 ; n20524
g20333 nor n20521 n20524 ; n20525
g20334 nor asqrt[12] n20506 ; n20526
g20335 and n20516_not n20526 ; n20527
g20336 nor n20525 n20527 ; n20528
g20337 nor n20518 n20528 ; n20529
g20338 and asqrt[13] n20529_not ; n20530
g20339 and n19814_not n19821 ; n20531
g20340 and n19823_not n20531 ; n20532
g20341 and asqrt[6] n20532 ; n20533
g20342 nor n19814 n19823 ; n20534
g20343 and asqrt[6] n20534 ; n20535
g20344 nor n19821 n20535 ; n20536
g20345 nor n20533 n20536 ; n20537
g20346 nor asqrt[13] n20518 ; n20538
g20347 and n20528_not n20538 ; n20539
g20348 nor n20537 n20539 ; n20540
g20349 nor n20530 n20540 ; n20541
g20350 and asqrt[14] n20541_not ; n20542
g20351 and n19833 n19835_not ; n20543
g20352 and n19826_not n20543 ; n20544
g20353 and asqrt[6] n20544 ; n20545
g20354 nor n19826 n19835 ; n20546
g20355 and asqrt[6] n20546 ; n20547
g20356 nor n19833 n20547 ; n20548
g20357 nor n20545 n20548 ; n20549
g20358 nor asqrt[14] n20530 ; n20550
g20359 and n20540_not n20550 ; n20551
g20360 nor n20549 n20551 ; n20552
g20361 nor n20542 n20552 ; n20553
g20362 and asqrt[15] n20553_not ; n20554
g20363 and n19838_not n19845 ; n20555
g20364 and n19847_not n20555 ; n20556
g20365 and asqrt[6] n20556 ; n20557
g20366 nor n19838 n19847 ; n20558
g20367 and asqrt[6] n20558 ; n20559
g20368 nor n19845 n20559 ; n20560
g20369 nor n20557 n20560 ; n20561
g20370 nor asqrt[15] n20542 ; n20562
g20371 and n20552_not n20562 ; n20563
g20372 nor n20561 n20563 ; n20564
g20373 nor n20554 n20564 ; n20565
g20374 and asqrt[16] n20565_not ; n20566
g20375 and n19857 n19859_not ; n20567
g20376 and n19850_not n20567 ; n20568
g20377 and asqrt[6] n20568 ; n20569
g20378 nor n19850 n19859 ; n20570
g20379 and asqrt[6] n20570 ; n20571
g20380 nor n19857 n20571 ; n20572
g20381 nor n20569 n20572 ; n20573
g20382 nor asqrt[16] n20554 ; n20574
g20383 and n20564_not n20574 ; n20575
g20384 nor n20573 n20575 ; n20576
g20385 nor n20566 n20576 ; n20577
g20386 and asqrt[17] n20577_not ; n20578
g20387 and n19862_not n19869 ; n20579
g20388 and n19871_not n20579 ; n20580
g20389 and asqrt[6] n20580 ; n20581
g20390 nor n19862 n19871 ; n20582
g20391 and asqrt[6] n20582 ; n20583
g20392 nor n19869 n20583 ; n20584
g20393 nor n20581 n20584 ; n20585
g20394 nor asqrt[17] n20566 ; n20586
g20395 and n20576_not n20586 ; n20587
g20396 nor n20585 n20587 ; n20588
g20397 nor n20578 n20588 ; n20589
g20398 and asqrt[18] n20589_not ; n20590
g20399 and n19881 n19883_not ; n20591
g20400 and n19874_not n20591 ; n20592
g20401 and asqrt[6] n20592 ; n20593
g20402 nor n19874 n19883 ; n20594
g20403 and asqrt[6] n20594 ; n20595
g20404 nor n19881 n20595 ; n20596
g20405 nor n20593 n20596 ; n20597
g20406 nor asqrt[18] n20578 ; n20598
g20407 and n20588_not n20598 ; n20599
g20408 nor n20597 n20599 ; n20600
g20409 nor n20590 n20600 ; n20601
g20410 and asqrt[19] n20601_not ; n20602
g20411 and n19886_not n19893 ; n20603
g20412 and n19895_not n20603 ; n20604
g20413 and asqrt[6] n20604 ; n20605
g20414 nor n19886 n19895 ; n20606
g20415 and asqrt[6] n20606 ; n20607
g20416 nor n19893 n20607 ; n20608
g20417 nor n20605 n20608 ; n20609
g20418 nor asqrt[19] n20590 ; n20610
g20419 and n20600_not n20610 ; n20611
g20420 nor n20609 n20611 ; n20612
g20421 nor n20602 n20612 ; n20613
g20422 and asqrt[20] n20613_not ; n20614
g20423 and n19905 n19907_not ; n20615
g20424 and n19898_not n20615 ; n20616
g20425 and asqrt[6] n20616 ; n20617
g20426 nor n19898 n19907 ; n20618
g20427 and asqrt[6] n20618 ; n20619
g20428 nor n19905 n20619 ; n20620
g20429 nor n20617 n20620 ; n20621
g20430 nor asqrt[20] n20602 ; n20622
g20431 and n20612_not n20622 ; n20623
g20432 nor n20621 n20623 ; n20624
g20433 nor n20614 n20624 ; n20625
g20434 and asqrt[21] n20625_not ; n20626
g20435 and n19910_not n19917 ; n20627
g20436 and n19919_not n20627 ; n20628
g20437 and asqrt[6] n20628 ; n20629
g20438 nor n19910 n19919 ; n20630
g20439 and asqrt[6] n20630 ; n20631
g20440 nor n19917 n20631 ; n20632
g20441 nor n20629 n20632 ; n20633
g20442 nor asqrt[21] n20614 ; n20634
g20443 and n20624_not n20634 ; n20635
g20444 nor n20633 n20635 ; n20636
g20445 nor n20626 n20636 ; n20637
g20446 and asqrt[22] n20637_not ; n20638
g20447 and n19929 n19931_not ; n20639
g20448 and n19922_not n20639 ; n20640
g20449 and asqrt[6] n20640 ; n20641
g20450 nor n19922 n19931 ; n20642
g20451 and asqrt[6] n20642 ; n20643
g20452 nor n19929 n20643 ; n20644
g20453 nor n20641 n20644 ; n20645
g20454 nor asqrt[22] n20626 ; n20646
g20455 and n20636_not n20646 ; n20647
g20456 nor n20645 n20647 ; n20648
g20457 nor n20638 n20648 ; n20649
g20458 and asqrt[23] n20649_not ; n20650
g20459 and n19934_not n19941 ; n20651
g20460 and n19943_not n20651 ; n20652
g20461 and asqrt[6] n20652 ; n20653
g20462 nor n19934 n19943 ; n20654
g20463 and asqrt[6] n20654 ; n20655
g20464 nor n19941 n20655 ; n20656
g20465 nor n20653 n20656 ; n20657
g20466 nor asqrt[23] n20638 ; n20658
g20467 and n20648_not n20658 ; n20659
g20468 nor n20657 n20659 ; n20660
g20469 nor n20650 n20660 ; n20661
g20470 and asqrt[24] n20661_not ; n20662
g20471 and n19953 n19955_not ; n20663
g20472 and n19946_not n20663 ; n20664
g20473 and asqrt[6] n20664 ; n20665
g20474 nor n19946 n19955 ; n20666
g20475 and asqrt[6] n20666 ; n20667
g20476 nor n19953 n20667 ; n20668
g20477 nor n20665 n20668 ; n20669
g20478 nor asqrt[24] n20650 ; n20670
g20479 and n20660_not n20670 ; n20671
g20480 nor n20669 n20671 ; n20672
g20481 nor n20662 n20672 ; n20673
g20482 and asqrt[25] n20673_not ; n20674
g20483 and n19958_not n19965 ; n20675
g20484 and n19967_not n20675 ; n20676
g20485 and asqrt[6] n20676 ; n20677
g20486 nor n19958 n19967 ; n20678
g20487 and asqrt[6] n20678 ; n20679
g20488 nor n19965 n20679 ; n20680
g20489 nor n20677 n20680 ; n20681
g20490 nor asqrt[25] n20662 ; n20682
g20491 and n20672_not n20682 ; n20683
g20492 nor n20681 n20683 ; n20684
g20493 nor n20674 n20684 ; n20685
g20494 and asqrt[26] n20685_not ; n20686
g20495 and n19977 n19979_not ; n20687
g20496 and n19970_not n20687 ; n20688
g20497 and asqrt[6] n20688 ; n20689
g20498 nor n19970 n19979 ; n20690
g20499 and asqrt[6] n20690 ; n20691
g20500 nor n19977 n20691 ; n20692
g20501 nor n20689 n20692 ; n20693
g20502 nor asqrt[26] n20674 ; n20694
g20503 and n20684_not n20694 ; n20695
g20504 nor n20693 n20695 ; n20696
g20505 nor n20686 n20696 ; n20697
g20506 and asqrt[27] n20697_not ; n20698
g20507 and n19982_not n19989 ; n20699
g20508 and n19991_not n20699 ; n20700
g20509 and asqrt[6] n20700 ; n20701
g20510 nor n19982 n19991 ; n20702
g20511 and asqrt[6] n20702 ; n20703
g20512 nor n19989 n20703 ; n20704
g20513 nor n20701 n20704 ; n20705
g20514 nor asqrt[27] n20686 ; n20706
g20515 and n20696_not n20706 ; n20707
g20516 nor n20705 n20707 ; n20708
g20517 nor n20698 n20708 ; n20709
g20518 and asqrt[28] n20709_not ; n20710
g20519 and n20001 n20003_not ; n20711
g20520 and n19994_not n20711 ; n20712
g20521 and asqrt[6] n20712 ; n20713
g20522 nor n19994 n20003 ; n20714
g20523 and asqrt[6] n20714 ; n20715
g20524 nor n20001 n20715 ; n20716
g20525 nor n20713 n20716 ; n20717
g20526 nor asqrt[28] n20698 ; n20718
g20527 and n20708_not n20718 ; n20719
g20528 nor n20717 n20719 ; n20720
g20529 nor n20710 n20720 ; n20721
g20530 and asqrt[29] n20721_not ; n20722
g20531 and n20006_not n20013 ; n20723
g20532 and n20015_not n20723 ; n20724
g20533 and asqrt[6] n20724 ; n20725
g20534 nor n20006 n20015 ; n20726
g20535 and asqrt[6] n20726 ; n20727
g20536 nor n20013 n20727 ; n20728
g20537 nor n20725 n20728 ; n20729
g20538 nor asqrt[29] n20710 ; n20730
g20539 and n20720_not n20730 ; n20731
g20540 nor n20729 n20731 ; n20732
g20541 nor n20722 n20732 ; n20733
g20542 and asqrt[30] n20733_not ; n20734
g20543 and n20025 n20027_not ; n20735
g20544 and n20018_not n20735 ; n20736
g20545 and asqrt[6] n20736 ; n20737
g20546 nor n20018 n20027 ; n20738
g20547 and asqrt[6] n20738 ; n20739
g20548 nor n20025 n20739 ; n20740
g20549 nor n20737 n20740 ; n20741
g20550 nor asqrt[30] n20722 ; n20742
g20551 and n20732_not n20742 ; n20743
g20552 nor n20741 n20743 ; n20744
g20553 nor n20734 n20744 ; n20745
g20554 and asqrt[31] n20745_not ; n20746
g20555 and n20030_not n20037 ; n20747
g20556 and n20039_not n20747 ; n20748
g20557 and asqrt[6] n20748 ; n20749
g20558 nor n20030 n20039 ; n20750
g20559 and asqrt[6] n20750 ; n20751
g20560 nor n20037 n20751 ; n20752
g20561 nor n20749 n20752 ; n20753
g20562 nor asqrt[31] n20734 ; n20754
g20563 and n20744_not n20754 ; n20755
g20564 nor n20753 n20755 ; n20756
g20565 nor n20746 n20756 ; n20757
g20566 and asqrt[32] n20757_not ; n20758
g20567 and n20049 n20051_not ; n20759
g20568 and n20042_not n20759 ; n20760
g20569 and asqrt[6] n20760 ; n20761
g20570 nor n20042 n20051 ; n20762
g20571 and asqrt[6] n20762 ; n20763
g20572 nor n20049 n20763 ; n20764
g20573 nor n20761 n20764 ; n20765
g20574 nor asqrt[32] n20746 ; n20766
g20575 and n20756_not n20766 ; n20767
g20576 nor n20765 n20767 ; n20768
g20577 nor n20758 n20768 ; n20769
g20578 and asqrt[33] n20769_not ; n20770
g20579 and n20054_not n20061 ; n20771
g20580 and n20063_not n20771 ; n20772
g20581 and asqrt[6] n20772 ; n20773
g20582 nor n20054 n20063 ; n20774
g20583 and asqrt[6] n20774 ; n20775
g20584 nor n20061 n20775 ; n20776
g20585 nor n20773 n20776 ; n20777
g20586 nor asqrt[33] n20758 ; n20778
g20587 and n20768_not n20778 ; n20779
g20588 nor n20777 n20779 ; n20780
g20589 nor n20770 n20780 ; n20781
g20590 and asqrt[34] n20781_not ; n20782
g20591 and n20073 n20075_not ; n20783
g20592 and n20066_not n20783 ; n20784
g20593 and asqrt[6] n20784 ; n20785
g20594 nor n20066 n20075 ; n20786
g20595 and asqrt[6] n20786 ; n20787
g20596 nor n20073 n20787 ; n20788
g20597 nor n20785 n20788 ; n20789
g20598 nor asqrt[34] n20770 ; n20790
g20599 and n20780_not n20790 ; n20791
g20600 nor n20789 n20791 ; n20792
g20601 nor n20782 n20792 ; n20793
g20602 and asqrt[35] n20793_not ; n20794
g20603 and n20078_not n20085 ; n20795
g20604 and n20087_not n20795 ; n20796
g20605 and asqrt[6] n20796 ; n20797
g20606 nor n20078 n20087 ; n20798
g20607 and asqrt[6] n20798 ; n20799
g20608 nor n20085 n20799 ; n20800
g20609 nor n20797 n20800 ; n20801
g20610 nor asqrt[35] n20782 ; n20802
g20611 and n20792_not n20802 ; n20803
g20612 nor n20801 n20803 ; n20804
g20613 nor n20794 n20804 ; n20805
g20614 and asqrt[36] n20805_not ; n20806
g20615 and n20097 n20099_not ; n20807
g20616 and n20090_not n20807 ; n20808
g20617 and asqrt[6] n20808 ; n20809
g20618 nor n20090 n20099 ; n20810
g20619 and asqrt[6] n20810 ; n20811
g20620 nor n20097 n20811 ; n20812
g20621 nor n20809 n20812 ; n20813
g20622 nor asqrt[36] n20794 ; n20814
g20623 and n20804_not n20814 ; n20815
g20624 nor n20813 n20815 ; n20816
g20625 nor n20806 n20816 ; n20817
g20626 and asqrt[37] n20817_not ; n20818
g20627 and n20102_not n20109 ; n20819
g20628 and n20111_not n20819 ; n20820
g20629 and asqrt[6] n20820 ; n20821
g20630 nor n20102 n20111 ; n20822
g20631 and asqrt[6] n20822 ; n20823
g20632 nor n20109 n20823 ; n20824
g20633 nor n20821 n20824 ; n20825
g20634 nor asqrt[37] n20806 ; n20826
g20635 and n20816_not n20826 ; n20827
g20636 nor n20825 n20827 ; n20828
g20637 nor n20818 n20828 ; n20829
g20638 and asqrt[38] n20829_not ; n20830
g20639 and n20121 n20123_not ; n20831
g20640 and n20114_not n20831 ; n20832
g20641 and asqrt[6] n20832 ; n20833
g20642 nor n20114 n20123 ; n20834
g20643 and asqrt[6] n20834 ; n20835
g20644 nor n20121 n20835 ; n20836
g20645 nor n20833 n20836 ; n20837
g20646 nor asqrt[38] n20818 ; n20838
g20647 and n20828_not n20838 ; n20839
g20648 nor n20837 n20839 ; n20840
g20649 nor n20830 n20840 ; n20841
g20650 and asqrt[39] n20841_not ; n20842
g20651 and n20126_not n20133 ; n20843
g20652 and n20135_not n20843 ; n20844
g20653 and asqrt[6] n20844 ; n20845
g20654 nor n20126 n20135 ; n20846
g20655 and asqrt[6] n20846 ; n20847
g20656 nor n20133 n20847 ; n20848
g20657 nor n20845 n20848 ; n20849
g20658 nor asqrt[39] n20830 ; n20850
g20659 and n20840_not n20850 ; n20851
g20660 nor n20849 n20851 ; n20852
g20661 nor n20842 n20852 ; n20853
g20662 and asqrt[40] n20853_not ; n20854
g20663 and n20145 n20147_not ; n20855
g20664 and n20138_not n20855 ; n20856
g20665 and asqrt[6] n20856 ; n20857
g20666 nor n20138 n20147 ; n20858
g20667 and asqrt[6] n20858 ; n20859
g20668 nor n20145 n20859 ; n20860
g20669 nor n20857 n20860 ; n20861
g20670 nor asqrt[40] n20842 ; n20862
g20671 and n20852_not n20862 ; n20863
g20672 nor n20861 n20863 ; n20864
g20673 nor n20854 n20864 ; n20865
g20674 and asqrt[41] n20865_not ; n20866
g20675 and n20150_not n20157 ; n20867
g20676 and n20159_not n20867 ; n20868
g20677 and asqrt[6] n20868 ; n20869
g20678 nor n20150 n20159 ; n20870
g20679 and asqrt[6] n20870 ; n20871
g20680 nor n20157 n20871 ; n20872
g20681 nor n20869 n20872 ; n20873
g20682 nor asqrt[41] n20854 ; n20874
g20683 and n20864_not n20874 ; n20875
g20684 nor n20873 n20875 ; n20876
g20685 nor n20866 n20876 ; n20877
g20686 and asqrt[42] n20877_not ; n20878
g20687 and n20169 n20171_not ; n20879
g20688 and n20162_not n20879 ; n20880
g20689 and asqrt[6] n20880 ; n20881
g20690 nor n20162 n20171 ; n20882
g20691 and asqrt[6] n20882 ; n20883
g20692 nor n20169 n20883 ; n20884
g20693 nor n20881 n20884 ; n20885
g20694 nor asqrt[42] n20866 ; n20886
g20695 and n20876_not n20886 ; n20887
g20696 nor n20885 n20887 ; n20888
g20697 nor n20878 n20888 ; n20889
g20698 and asqrt[43] n20889_not ; n20890
g20699 and n20174_not n20181 ; n20891
g20700 and n20183_not n20891 ; n20892
g20701 and asqrt[6] n20892 ; n20893
g20702 nor n20174 n20183 ; n20894
g20703 and asqrt[6] n20894 ; n20895
g20704 nor n20181 n20895 ; n20896
g20705 nor n20893 n20896 ; n20897
g20706 nor asqrt[43] n20878 ; n20898
g20707 and n20888_not n20898 ; n20899
g20708 nor n20897 n20899 ; n20900
g20709 nor n20890 n20900 ; n20901
g20710 and asqrt[44] n20901_not ; n20902
g20711 and n20193 n20195_not ; n20903
g20712 and n20186_not n20903 ; n20904
g20713 and asqrt[6] n20904 ; n20905
g20714 nor n20186 n20195 ; n20906
g20715 and asqrt[6] n20906 ; n20907
g20716 nor n20193 n20907 ; n20908
g20717 nor n20905 n20908 ; n20909
g20718 nor asqrt[44] n20890 ; n20910
g20719 and n20900_not n20910 ; n20911
g20720 nor n20909 n20911 ; n20912
g20721 nor n20902 n20912 ; n20913
g20722 and asqrt[45] n20913_not ; n20914
g20723 and n20198_not n20205 ; n20915
g20724 and n20207_not n20915 ; n20916
g20725 and asqrt[6] n20916 ; n20917
g20726 nor n20198 n20207 ; n20918
g20727 and asqrt[6] n20918 ; n20919
g20728 nor n20205 n20919 ; n20920
g20729 nor n20917 n20920 ; n20921
g20730 nor asqrt[45] n20902 ; n20922
g20731 and n20912_not n20922 ; n20923
g20732 nor n20921 n20923 ; n20924
g20733 nor n20914 n20924 ; n20925
g20734 and asqrt[46] n20925_not ; n20926
g20735 and n20217 n20219_not ; n20927
g20736 and n20210_not n20927 ; n20928
g20737 and asqrt[6] n20928 ; n20929
g20738 nor n20210 n20219 ; n20930
g20739 and asqrt[6] n20930 ; n20931
g20740 nor n20217 n20931 ; n20932
g20741 nor n20929 n20932 ; n20933
g20742 nor asqrt[46] n20914 ; n20934
g20743 and n20924_not n20934 ; n20935
g20744 nor n20933 n20935 ; n20936
g20745 nor n20926 n20936 ; n20937
g20746 and asqrt[47] n20937_not ; n20938
g20747 and n20222_not n20229 ; n20939
g20748 and n20231_not n20939 ; n20940
g20749 and asqrt[6] n20940 ; n20941
g20750 nor n20222 n20231 ; n20942
g20751 and asqrt[6] n20942 ; n20943
g20752 nor n20229 n20943 ; n20944
g20753 nor n20941 n20944 ; n20945
g20754 nor asqrt[47] n20926 ; n20946
g20755 and n20936_not n20946 ; n20947
g20756 nor n20945 n20947 ; n20948
g20757 nor n20938 n20948 ; n20949
g20758 and asqrt[48] n20949_not ; n20950
g20759 and n20241 n20243_not ; n20951
g20760 and n20234_not n20951 ; n20952
g20761 and asqrt[6] n20952 ; n20953
g20762 nor n20234 n20243 ; n20954
g20763 and asqrt[6] n20954 ; n20955
g20764 nor n20241 n20955 ; n20956
g20765 nor n20953 n20956 ; n20957
g20766 nor asqrt[48] n20938 ; n20958
g20767 and n20948_not n20958 ; n20959
g20768 nor n20957 n20959 ; n20960
g20769 nor n20950 n20960 ; n20961
g20770 and asqrt[49] n20961_not ; n20962
g20771 and n20246_not n20253 ; n20963
g20772 and n20255_not n20963 ; n20964
g20773 and asqrt[6] n20964 ; n20965
g20774 nor n20246 n20255 ; n20966
g20775 and asqrt[6] n20966 ; n20967
g20776 nor n20253 n20967 ; n20968
g20777 nor n20965 n20968 ; n20969
g20778 nor asqrt[49] n20950 ; n20970
g20779 and n20960_not n20970 ; n20971
g20780 nor n20969 n20971 ; n20972
g20781 nor n20962 n20972 ; n20973
g20782 and asqrt[50] n20973_not ; n20974
g20783 and n20265 n20267_not ; n20975
g20784 and n20258_not n20975 ; n20976
g20785 and asqrt[6] n20976 ; n20977
g20786 nor n20258 n20267 ; n20978
g20787 and asqrt[6] n20978 ; n20979
g20788 nor n20265 n20979 ; n20980
g20789 nor n20977 n20980 ; n20981
g20790 nor asqrt[50] n20962 ; n20982
g20791 and n20972_not n20982 ; n20983
g20792 nor n20981 n20983 ; n20984
g20793 nor n20974 n20984 ; n20985
g20794 and asqrt[51] n20985_not ; n20986
g20795 and n20270_not n20277 ; n20987
g20796 and n20279_not n20987 ; n20988
g20797 and asqrt[6] n20988 ; n20989
g20798 nor n20270 n20279 ; n20990
g20799 and asqrt[6] n20990 ; n20991
g20800 nor n20277 n20991 ; n20992
g20801 nor n20989 n20992 ; n20993
g20802 nor asqrt[51] n20974 ; n20994
g20803 and n20984_not n20994 ; n20995
g20804 nor n20993 n20995 ; n20996
g20805 nor n20986 n20996 ; n20997
g20806 and asqrt[52] n20997_not ; n20998
g20807 and n20289 n20291_not ; n20999
g20808 and n20282_not n20999 ; n21000
g20809 and asqrt[6] n21000 ; n21001
g20810 nor n20282 n20291 ; n21002
g20811 and asqrt[6] n21002 ; n21003
g20812 nor n20289 n21003 ; n21004
g20813 nor n21001 n21004 ; n21005
g20814 nor asqrt[52] n20986 ; n21006
g20815 and n20996_not n21006 ; n21007
g20816 nor n21005 n21007 ; n21008
g20817 nor n20998 n21008 ; n21009
g20818 and asqrt[53] n21009_not ; n21010
g20819 and n20294_not n20301 ; n21011
g20820 and n20303_not n21011 ; n21012
g20821 and asqrt[6] n21012 ; n21013
g20822 nor n20294 n20303 ; n21014
g20823 and asqrt[6] n21014 ; n21015
g20824 nor n20301 n21015 ; n21016
g20825 nor n21013 n21016 ; n21017
g20826 nor asqrt[53] n20998 ; n21018
g20827 and n21008_not n21018 ; n21019
g20828 nor n21017 n21019 ; n21020
g20829 nor n21010 n21020 ; n21021
g20830 and asqrt[54] n21021_not ; n21022
g20831 and n20313 n20315_not ; n21023
g20832 and n20306_not n21023 ; n21024
g20833 and asqrt[6] n21024 ; n21025
g20834 nor n20306 n20315 ; n21026
g20835 and asqrt[6] n21026 ; n21027
g20836 nor n20313 n21027 ; n21028
g20837 nor n21025 n21028 ; n21029
g20838 nor asqrt[54] n21010 ; n21030
g20839 and n21020_not n21030 ; n21031
g20840 nor n21029 n21031 ; n21032
g20841 nor n21022 n21032 ; n21033
g20842 and asqrt[55] n21033_not ; n21034
g20843 and n20318_not n20325 ; n21035
g20844 and n20327_not n21035 ; n21036
g20845 and asqrt[6] n21036 ; n21037
g20846 nor n20318 n20327 ; n21038
g20847 and asqrt[6] n21038 ; n21039
g20848 nor n20325 n21039 ; n21040
g20849 nor n21037 n21040 ; n21041
g20850 nor asqrt[55] n21022 ; n21042
g20851 and n21032_not n21042 ; n21043
g20852 nor n21041 n21043 ; n21044
g20853 nor n21034 n21044 ; n21045
g20854 and asqrt[56] n21045_not ; n21046
g20855 and n20337 n20339_not ; n21047
g20856 and n20330_not n21047 ; n21048
g20857 and asqrt[6] n21048 ; n21049
g20858 nor n20330 n20339 ; n21050
g20859 and asqrt[6] n21050 ; n21051
g20860 nor n20337 n21051 ; n21052
g20861 nor n21049 n21052 ; n21053
g20862 nor asqrt[56] n21034 ; n21054
g20863 and n21044_not n21054 ; n21055
g20864 nor n21053 n21055 ; n21056
g20865 nor n21046 n21056 ; n21057
g20866 and asqrt[57] n21057_not ; n21058
g20867 and n20342_not n20349 ; n21059
g20868 and n20351_not n21059 ; n21060
g20869 and asqrt[6] n21060 ; n21061
g20870 nor n20342 n20351 ; n21062
g20871 and asqrt[6] n21062 ; n21063
g20872 nor n20349 n21063 ; n21064
g20873 nor n21061 n21064 ; n21065
g20874 nor asqrt[57] n21046 ; n21066
g20875 and n21056_not n21066 ; n21067
g20876 nor n21065 n21067 ; n21068
g20877 nor n21058 n21068 ; n21069
g20878 and asqrt[58] n21069_not ; n21070
g20879 and n20361 n20363_not ; n21071
g20880 and n20354_not n21071 ; n21072
g20881 and asqrt[6] n21072 ; n21073
g20882 nor n20354 n20363 ; n21074
g20883 and asqrt[6] n21074 ; n21075
g20884 nor n20361 n21075 ; n21076
g20885 nor n21073 n21076 ; n21077
g20886 nor asqrt[58] n21058 ; n21078
g20887 and n21068_not n21078 ; n21079
g20888 nor n21077 n21079 ; n21080
g20889 nor n21070 n21080 ; n21081
g20890 and asqrt[59] n21081_not ; n21082
g20891 nor asqrt[59] n21070 ; n21083
g20892 and n21080_not n21083 ; n21084
g20893 and n20366_not n20375 ; n21085
g20894 and n20368_not n21085 ; n21086
g20895 and asqrt[6] n21086 ; n21087
g20896 nor n20366 n20368 ; n21088
g20897 and asqrt[6] n21088 ; n21089
g20898 nor n20375 n21089 ; n21090
g20899 nor n21087 n21090 ; n21091
g20900 nor n21084 n21091 ; n21092
g20901 nor n21082 n21092 ; n21093
g20902 and asqrt[60] n21093_not ; n21094
g20903 and n20385 n20387_not ; n21095
g20904 and n20378_not n21095 ; n21096
g20905 and asqrt[6] n21096 ; n21097
g20906 nor n20378 n20387 ; n21098
g20907 and asqrt[6] n21098 ; n21099
g20908 nor n20385 n21099 ; n21100
g20909 nor n21097 n21100 ; n21101
g20910 nor asqrt[60] n21082 ; n21102
g20911 and n21092_not n21102 ; n21103
g20912 nor n21101 n21103 ; n21104
g20913 nor n21094 n21104 ; n21105
g20914 and asqrt[61] n21105_not ; n21106
g20915 and n20390_not n20397 ; n21107
g20916 and n20399_not n21107 ; n21108
g20917 and asqrt[6] n21108 ; n21109
g20918 nor n20390 n20399 ; n21110
g20919 and asqrt[6] n21110 ; n21111
g20920 nor n20397 n21111 ; n21112
g20921 nor n21109 n21112 ; n21113
g20922 nor asqrt[61] n21094 ; n21114
g20923 and n21104_not n21114 ; n21115
g20924 nor n21113 n21115 ; n21116
g20925 nor n21106 n21116 ; n21117
g20926 and asqrt[62] n21117_not ; n21118
g20927 and n20409 n20411_not ; n21119
g20928 and n20402_not n21119 ; n21120
g20929 and asqrt[6] n21120 ; n21121
g20930 nor n20402 n20411 ; n21122
g20931 and asqrt[6] n21122 ; n21123
g20932 nor n20409 n21123 ; n21124
g20933 nor n21121 n21124 ; n21125
g20934 nor asqrt[62] n21106 ; n21126
g20935 and n21116_not n21126 ; n21127
g20936 nor n21125 n21127 ; n21128
g20937 nor n21118 n21128 ; n21129
g20938 and n20414_not n20421 ; n21130
g20939 and n20423_not n21130 ; n21131
g20940 and asqrt[6] n21131 ; n21132
g20941 nor n20414 n20423 ; n21133
g20942 and asqrt[6] n21133 ; n21134
g20943 nor n20421 n21134 ; n21135
g20944 nor n21132 n21135 ; n21136
g20945 nor n20425 n20432 ; n21137
g20946 and asqrt[6] n21137 ; n21138
g20947 nor n20440 n21138 ; n21139
g20948 and n21136_not n21139 ; n21140
g20949 and n21129_not n21140 ; n21141
g20950 nor asqrt[63] n21141 ; n21142
g20951 and n21118_not n21136 ; n21143
g20952 and n21128_not n21143 ; n21144
g20953 and n20432_not asqrt[6] ; n21145
g20954 and n20425 n21145_not ; n21146
g20955 and asqrt[63] n21137_not ; n21147
g20956 and n21146_not n21147 ; n21148
g20957 nor n21144 n21148 ; n21149
g20958 nand n21142_not n21149 ; asqrt[5]
g20959 and a[10] asqrt[5] ; n21151
g20960 nor a[8] a[9] ; n21152
g20961 and a[10]_not n21152 ; n21153
g20962 nor n21151 n21153 ; n21154
g20963 and asqrt[6] n21154_not ; n21155
g20964 nor n20449 n21153 ; n21156
g20965 and n20444_not n21156 ; n21157
g20966 and n20440_not n21157 ; n21158
g20967 and n20438_not n21158 ; n21159
g20968 and n21151_not n21159 ; n21160
g20969 and a[10]_not asqrt[5] ; n21161
g20970 and a[11] n21161_not ; n21162
g20971 and n20454 asqrt[5] ; n21163
g20972 nor n21162 n21163 ; n21164
g20973 and n21160_not n21164 ; n21165
g20974 nor n21155 n21165 ; n21166
g20975 and asqrt[7] n21166_not ; n21167
g20976 nor asqrt[7] n21155 ; n21168
g20977 and n21165_not n21168 ; n21169
g20978 and asqrt[6] n21148_not ; n21170
g20979 and n21144_not n21170 ; n21171
g20980 and n21142_not n21171 ; n21172
g20981 nor n21163 n21172 ; n21173
g20982 and a[12] n21173_not ; n21174
g20983 nor a[12] n21172 ; n21175
g20984 and n21163_not n21175 ; n21176
g20985 nor n21174 n21176 ; n21177
g20986 nor n21169 n21177 ; n21178
g20987 nor n21167 n21178 ; n21179
g20988 and asqrt[8] n21179_not ; n21180
g20989 nor n20457 n20462 ; n21181
g20990 and n20466_not n21181 ; n21182
g20991 and asqrt[5] n21182 ; n21183
g20992 and asqrt[5] n21181 ; n21184
g20993 and n20466 n21184_not ; n21185
g20994 nor n21183 n21185 ; n21186
g20995 nor asqrt[8] n21167 ; n21187
g20996 and n21178_not n21187 ; n21188
g20997 nor n21186 n21188 ; n21189
g20998 nor n21180 n21189 ; n21190
g20999 and asqrt[9] n21190_not ; n21191
g21000 and n20471_not n20480 ; n21192
g21001 and n20469_not n21192 ; n21193
g21002 and asqrt[5] n21193 ; n21194
g21003 nor n20469 n20471 ; n21195
g21004 and asqrt[5] n21195 ; n21196
g21005 nor n20480 n21196 ; n21197
g21006 nor n21194 n21197 ; n21198
g21007 nor asqrt[9] n21180 ; n21199
g21008 and n21189_not n21199 ; n21200
g21009 nor n21198 n21200 ; n21201
g21010 nor n21191 n21201 ; n21202
g21011 and asqrt[10] n21202_not ; n21203
g21012 and n20483_not n20489 ; n21204
g21013 and n20491_not n21204 ; n21205
g21014 and asqrt[5] n21205 ; n21206
g21015 nor n20483 n20491 ; n21207
g21016 and asqrt[5] n21207 ; n21208
g21017 nor n20489 n21208 ; n21209
g21018 nor n21206 n21209 ; n21210
g21019 nor asqrt[10] n21191 ; n21211
g21020 and n21201_not n21211 ; n21212
g21021 nor n21210 n21212 ; n21213
g21022 nor n21203 n21213 ; n21214
g21023 and asqrt[11] n21214_not ; n21215
g21024 and n20501 n20503_not ; n21216
g21025 and n20494_not n21216 ; n21217
g21026 and asqrt[5] n21217 ; n21218
g21027 nor n20494 n20503 ; n21219
g21028 and asqrt[5] n21219 ; n21220
g21029 nor n20501 n21220 ; n21221
g21030 nor n21218 n21221 ; n21222
g21031 nor asqrt[11] n21203 ; n21223
g21032 and n21213_not n21223 ; n21224
g21033 nor n21222 n21224 ; n21225
g21034 nor n21215 n21225 ; n21226
g21035 and asqrt[12] n21226_not ; n21227
g21036 and n20506_not n20513 ; n21228
g21037 and n20515_not n21228 ; n21229
g21038 and asqrt[5] n21229 ; n21230
g21039 nor n20506 n20515 ; n21231
g21040 and asqrt[5] n21231 ; n21232
g21041 nor n20513 n21232 ; n21233
g21042 nor n21230 n21233 ; n21234
g21043 nor asqrt[12] n21215 ; n21235
g21044 and n21225_not n21235 ; n21236
g21045 nor n21234 n21236 ; n21237
g21046 nor n21227 n21237 ; n21238
g21047 and asqrt[13] n21238_not ; n21239
g21048 and n20525 n20527_not ; n21240
g21049 and n20518_not n21240 ; n21241
g21050 and asqrt[5] n21241 ; n21242
g21051 nor n20518 n20527 ; n21243
g21052 and asqrt[5] n21243 ; n21244
g21053 nor n20525 n21244 ; n21245
g21054 nor n21242 n21245 ; n21246
g21055 nor asqrt[13] n21227 ; n21247
g21056 and n21237_not n21247 ; n21248
g21057 nor n21246 n21248 ; n21249
g21058 nor n21239 n21249 ; n21250
g21059 and asqrt[14] n21250_not ; n21251
g21060 and n20530_not n20537 ; n21252
g21061 and n20539_not n21252 ; n21253
g21062 and asqrt[5] n21253 ; n21254
g21063 nor n20530 n20539 ; n21255
g21064 and asqrt[5] n21255 ; n21256
g21065 nor n20537 n21256 ; n21257
g21066 nor n21254 n21257 ; n21258
g21067 nor asqrt[14] n21239 ; n21259
g21068 and n21249_not n21259 ; n21260
g21069 nor n21258 n21260 ; n21261
g21070 nor n21251 n21261 ; n21262
g21071 and asqrt[15] n21262_not ; n21263
g21072 and n20549 n20551_not ; n21264
g21073 and n20542_not n21264 ; n21265
g21074 and asqrt[5] n21265 ; n21266
g21075 nor n20542 n20551 ; n21267
g21076 and asqrt[5] n21267 ; n21268
g21077 nor n20549 n21268 ; n21269
g21078 nor n21266 n21269 ; n21270
g21079 nor asqrt[15] n21251 ; n21271
g21080 and n21261_not n21271 ; n21272
g21081 nor n21270 n21272 ; n21273
g21082 nor n21263 n21273 ; n21274
g21083 and asqrt[16] n21274_not ; n21275
g21084 and n20554_not n20561 ; n21276
g21085 and n20563_not n21276 ; n21277
g21086 and asqrt[5] n21277 ; n21278
g21087 nor n20554 n20563 ; n21279
g21088 and asqrt[5] n21279 ; n21280
g21089 nor n20561 n21280 ; n21281
g21090 nor n21278 n21281 ; n21282
g21091 nor asqrt[16] n21263 ; n21283
g21092 and n21273_not n21283 ; n21284
g21093 nor n21282 n21284 ; n21285
g21094 nor n21275 n21285 ; n21286
g21095 and asqrt[17] n21286_not ; n21287
g21096 and n20573 n20575_not ; n21288
g21097 and n20566_not n21288 ; n21289
g21098 and asqrt[5] n21289 ; n21290
g21099 nor n20566 n20575 ; n21291
g21100 and asqrt[5] n21291 ; n21292
g21101 nor n20573 n21292 ; n21293
g21102 nor n21290 n21293 ; n21294
g21103 nor asqrt[17] n21275 ; n21295
g21104 and n21285_not n21295 ; n21296
g21105 nor n21294 n21296 ; n21297
g21106 nor n21287 n21297 ; n21298
g21107 and asqrt[18] n21298_not ; n21299
g21108 and n20578_not n20585 ; n21300
g21109 and n20587_not n21300 ; n21301
g21110 and asqrt[5] n21301 ; n21302
g21111 nor n20578 n20587 ; n21303
g21112 and asqrt[5] n21303 ; n21304
g21113 nor n20585 n21304 ; n21305
g21114 nor n21302 n21305 ; n21306
g21115 nor asqrt[18] n21287 ; n21307
g21116 and n21297_not n21307 ; n21308
g21117 nor n21306 n21308 ; n21309
g21118 nor n21299 n21309 ; n21310
g21119 and asqrt[19] n21310_not ; n21311
g21120 and n20597 n20599_not ; n21312
g21121 and n20590_not n21312 ; n21313
g21122 and asqrt[5] n21313 ; n21314
g21123 nor n20590 n20599 ; n21315
g21124 and asqrt[5] n21315 ; n21316
g21125 nor n20597 n21316 ; n21317
g21126 nor n21314 n21317 ; n21318
g21127 nor asqrt[19] n21299 ; n21319
g21128 and n21309_not n21319 ; n21320
g21129 nor n21318 n21320 ; n21321
g21130 nor n21311 n21321 ; n21322
g21131 and asqrt[20] n21322_not ; n21323
g21132 and n20602_not n20609 ; n21324
g21133 and n20611_not n21324 ; n21325
g21134 and asqrt[5] n21325 ; n21326
g21135 nor n20602 n20611 ; n21327
g21136 and asqrt[5] n21327 ; n21328
g21137 nor n20609 n21328 ; n21329
g21138 nor n21326 n21329 ; n21330
g21139 nor asqrt[20] n21311 ; n21331
g21140 and n21321_not n21331 ; n21332
g21141 nor n21330 n21332 ; n21333
g21142 nor n21323 n21333 ; n21334
g21143 and asqrt[21] n21334_not ; n21335
g21144 and n20621 n20623_not ; n21336
g21145 and n20614_not n21336 ; n21337
g21146 and asqrt[5] n21337 ; n21338
g21147 nor n20614 n20623 ; n21339
g21148 and asqrt[5] n21339 ; n21340
g21149 nor n20621 n21340 ; n21341
g21150 nor n21338 n21341 ; n21342
g21151 nor asqrt[21] n21323 ; n21343
g21152 and n21333_not n21343 ; n21344
g21153 nor n21342 n21344 ; n21345
g21154 nor n21335 n21345 ; n21346
g21155 and asqrt[22] n21346_not ; n21347
g21156 and n20626_not n20633 ; n21348
g21157 and n20635_not n21348 ; n21349
g21158 and asqrt[5] n21349 ; n21350
g21159 nor n20626 n20635 ; n21351
g21160 and asqrt[5] n21351 ; n21352
g21161 nor n20633 n21352 ; n21353
g21162 nor n21350 n21353 ; n21354
g21163 nor asqrt[22] n21335 ; n21355
g21164 and n21345_not n21355 ; n21356
g21165 nor n21354 n21356 ; n21357
g21166 nor n21347 n21357 ; n21358
g21167 and asqrt[23] n21358_not ; n21359
g21168 and n20645 n20647_not ; n21360
g21169 and n20638_not n21360 ; n21361
g21170 and asqrt[5] n21361 ; n21362
g21171 nor n20638 n20647 ; n21363
g21172 and asqrt[5] n21363 ; n21364
g21173 nor n20645 n21364 ; n21365
g21174 nor n21362 n21365 ; n21366
g21175 nor asqrt[23] n21347 ; n21367
g21176 and n21357_not n21367 ; n21368
g21177 nor n21366 n21368 ; n21369
g21178 nor n21359 n21369 ; n21370
g21179 and asqrt[24] n21370_not ; n21371
g21180 and n20650_not n20657 ; n21372
g21181 and n20659_not n21372 ; n21373
g21182 and asqrt[5] n21373 ; n21374
g21183 nor n20650 n20659 ; n21375
g21184 and asqrt[5] n21375 ; n21376
g21185 nor n20657 n21376 ; n21377
g21186 nor n21374 n21377 ; n21378
g21187 nor asqrt[24] n21359 ; n21379
g21188 and n21369_not n21379 ; n21380
g21189 nor n21378 n21380 ; n21381
g21190 nor n21371 n21381 ; n21382
g21191 and asqrt[25] n21382_not ; n21383
g21192 and n20669 n20671_not ; n21384
g21193 and n20662_not n21384 ; n21385
g21194 and asqrt[5] n21385 ; n21386
g21195 nor n20662 n20671 ; n21387
g21196 and asqrt[5] n21387 ; n21388
g21197 nor n20669 n21388 ; n21389
g21198 nor n21386 n21389 ; n21390
g21199 nor asqrt[25] n21371 ; n21391
g21200 and n21381_not n21391 ; n21392
g21201 nor n21390 n21392 ; n21393
g21202 nor n21383 n21393 ; n21394
g21203 and asqrt[26] n21394_not ; n21395
g21204 and n20674_not n20681 ; n21396
g21205 and n20683_not n21396 ; n21397
g21206 and asqrt[5] n21397 ; n21398
g21207 nor n20674 n20683 ; n21399
g21208 and asqrt[5] n21399 ; n21400
g21209 nor n20681 n21400 ; n21401
g21210 nor n21398 n21401 ; n21402
g21211 nor asqrt[26] n21383 ; n21403
g21212 and n21393_not n21403 ; n21404
g21213 nor n21402 n21404 ; n21405
g21214 nor n21395 n21405 ; n21406
g21215 and asqrt[27] n21406_not ; n21407
g21216 and n20693 n20695_not ; n21408
g21217 and n20686_not n21408 ; n21409
g21218 and asqrt[5] n21409 ; n21410
g21219 nor n20686 n20695 ; n21411
g21220 and asqrt[5] n21411 ; n21412
g21221 nor n20693 n21412 ; n21413
g21222 nor n21410 n21413 ; n21414
g21223 nor asqrt[27] n21395 ; n21415
g21224 and n21405_not n21415 ; n21416
g21225 nor n21414 n21416 ; n21417
g21226 nor n21407 n21417 ; n21418
g21227 and asqrt[28] n21418_not ; n21419
g21228 and n20698_not n20705 ; n21420
g21229 and n20707_not n21420 ; n21421
g21230 and asqrt[5] n21421 ; n21422
g21231 nor n20698 n20707 ; n21423
g21232 and asqrt[5] n21423 ; n21424
g21233 nor n20705 n21424 ; n21425
g21234 nor n21422 n21425 ; n21426
g21235 nor asqrt[28] n21407 ; n21427
g21236 and n21417_not n21427 ; n21428
g21237 nor n21426 n21428 ; n21429
g21238 nor n21419 n21429 ; n21430
g21239 and asqrt[29] n21430_not ; n21431
g21240 and n20717 n20719_not ; n21432
g21241 and n20710_not n21432 ; n21433
g21242 and asqrt[5] n21433 ; n21434
g21243 nor n20710 n20719 ; n21435
g21244 and asqrt[5] n21435 ; n21436
g21245 nor n20717 n21436 ; n21437
g21246 nor n21434 n21437 ; n21438
g21247 nor asqrt[29] n21419 ; n21439
g21248 and n21429_not n21439 ; n21440
g21249 nor n21438 n21440 ; n21441
g21250 nor n21431 n21441 ; n21442
g21251 and asqrt[30] n21442_not ; n21443
g21252 and n20722_not n20729 ; n21444
g21253 and n20731_not n21444 ; n21445
g21254 and asqrt[5] n21445 ; n21446
g21255 nor n20722 n20731 ; n21447
g21256 and asqrt[5] n21447 ; n21448
g21257 nor n20729 n21448 ; n21449
g21258 nor n21446 n21449 ; n21450
g21259 nor asqrt[30] n21431 ; n21451
g21260 and n21441_not n21451 ; n21452
g21261 nor n21450 n21452 ; n21453
g21262 nor n21443 n21453 ; n21454
g21263 and asqrt[31] n21454_not ; n21455
g21264 and n20741 n20743_not ; n21456
g21265 and n20734_not n21456 ; n21457
g21266 and asqrt[5] n21457 ; n21458
g21267 nor n20734 n20743 ; n21459
g21268 and asqrt[5] n21459 ; n21460
g21269 nor n20741 n21460 ; n21461
g21270 nor n21458 n21461 ; n21462
g21271 nor asqrt[31] n21443 ; n21463
g21272 and n21453_not n21463 ; n21464
g21273 nor n21462 n21464 ; n21465
g21274 nor n21455 n21465 ; n21466
g21275 and asqrt[32] n21466_not ; n21467
g21276 and n20746_not n20753 ; n21468
g21277 and n20755_not n21468 ; n21469
g21278 and asqrt[5] n21469 ; n21470
g21279 nor n20746 n20755 ; n21471
g21280 and asqrt[5] n21471 ; n21472
g21281 nor n20753 n21472 ; n21473
g21282 nor n21470 n21473 ; n21474
g21283 nor asqrt[32] n21455 ; n21475
g21284 and n21465_not n21475 ; n21476
g21285 nor n21474 n21476 ; n21477
g21286 nor n21467 n21477 ; n21478
g21287 and asqrt[33] n21478_not ; n21479
g21288 and n20765 n20767_not ; n21480
g21289 and n20758_not n21480 ; n21481
g21290 and asqrt[5] n21481 ; n21482
g21291 nor n20758 n20767 ; n21483
g21292 and asqrt[5] n21483 ; n21484
g21293 nor n20765 n21484 ; n21485
g21294 nor n21482 n21485 ; n21486
g21295 nor asqrt[33] n21467 ; n21487
g21296 and n21477_not n21487 ; n21488
g21297 nor n21486 n21488 ; n21489
g21298 nor n21479 n21489 ; n21490
g21299 and asqrt[34] n21490_not ; n21491
g21300 and n20770_not n20777 ; n21492
g21301 and n20779_not n21492 ; n21493
g21302 and asqrt[5] n21493 ; n21494
g21303 nor n20770 n20779 ; n21495
g21304 and asqrt[5] n21495 ; n21496
g21305 nor n20777 n21496 ; n21497
g21306 nor n21494 n21497 ; n21498
g21307 nor asqrt[34] n21479 ; n21499
g21308 and n21489_not n21499 ; n21500
g21309 nor n21498 n21500 ; n21501
g21310 nor n21491 n21501 ; n21502
g21311 and asqrt[35] n21502_not ; n21503
g21312 and n20789 n20791_not ; n21504
g21313 and n20782_not n21504 ; n21505
g21314 and asqrt[5] n21505 ; n21506
g21315 nor n20782 n20791 ; n21507
g21316 and asqrt[5] n21507 ; n21508
g21317 nor n20789 n21508 ; n21509
g21318 nor n21506 n21509 ; n21510
g21319 nor asqrt[35] n21491 ; n21511
g21320 and n21501_not n21511 ; n21512
g21321 nor n21510 n21512 ; n21513
g21322 nor n21503 n21513 ; n21514
g21323 and asqrt[36] n21514_not ; n21515
g21324 and n20794_not n20801 ; n21516
g21325 and n20803_not n21516 ; n21517
g21326 and asqrt[5] n21517 ; n21518
g21327 nor n20794 n20803 ; n21519
g21328 and asqrt[5] n21519 ; n21520
g21329 nor n20801 n21520 ; n21521
g21330 nor n21518 n21521 ; n21522
g21331 nor asqrt[36] n21503 ; n21523
g21332 and n21513_not n21523 ; n21524
g21333 nor n21522 n21524 ; n21525
g21334 nor n21515 n21525 ; n21526
g21335 and asqrt[37] n21526_not ; n21527
g21336 and n20813 n20815_not ; n21528
g21337 and n20806_not n21528 ; n21529
g21338 and asqrt[5] n21529 ; n21530
g21339 nor n20806 n20815 ; n21531
g21340 and asqrt[5] n21531 ; n21532
g21341 nor n20813 n21532 ; n21533
g21342 nor n21530 n21533 ; n21534
g21343 nor asqrt[37] n21515 ; n21535
g21344 and n21525_not n21535 ; n21536
g21345 nor n21534 n21536 ; n21537
g21346 nor n21527 n21537 ; n21538
g21347 and asqrt[38] n21538_not ; n21539
g21348 and n20818_not n20825 ; n21540
g21349 and n20827_not n21540 ; n21541
g21350 and asqrt[5] n21541 ; n21542
g21351 nor n20818 n20827 ; n21543
g21352 and asqrt[5] n21543 ; n21544
g21353 nor n20825 n21544 ; n21545
g21354 nor n21542 n21545 ; n21546
g21355 nor asqrt[38] n21527 ; n21547
g21356 and n21537_not n21547 ; n21548
g21357 nor n21546 n21548 ; n21549
g21358 nor n21539 n21549 ; n21550
g21359 and asqrt[39] n21550_not ; n21551
g21360 and n20837 n20839_not ; n21552
g21361 and n20830_not n21552 ; n21553
g21362 and asqrt[5] n21553 ; n21554
g21363 nor n20830 n20839 ; n21555
g21364 and asqrt[5] n21555 ; n21556
g21365 nor n20837 n21556 ; n21557
g21366 nor n21554 n21557 ; n21558
g21367 nor asqrt[39] n21539 ; n21559
g21368 and n21549_not n21559 ; n21560
g21369 nor n21558 n21560 ; n21561
g21370 nor n21551 n21561 ; n21562
g21371 and asqrt[40] n21562_not ; n21563
g21372 and n20842_not n20849 ; n21564
g21373 and n20851_not n21564 ; n21565
g21374 and asqrt[5] n21565 ; n21566
g21375 nor n20842 n20851 ; n21567
g21376 and asqrt[5] n21567 ; n21568
g21377 nor n20849 n21568 ; n21569
g21378 nor n21566 n21569 ; n21570
g21379 nor asqrt[40] n21551 ; n21571
g21380 and n21561_not n21571 ; n21572
g21381 nor n21570 n21572 ; n21573
g21382 nor n21563 n21573 ; n21574
g21383 and asqrt[41] n21574_not ; n21575
g21384 and n20861 n20863_not ; n21576
g21385 and n20854_not n21576 ; n21577
g21386 and asqrt[5] n21577 ; n21578
g21387 nor n20854 n20863 ; n21579
g21388 and asqrt[5] n21579 ; n21580
g21389 nor n20861 n21580 ; n21581
g21390 nor n21578 n21581 ; n21582
g21391 nor asqrt[41] n21563 ; n21583
g21392 and n21573_not n21583 ; n21584
g21393 nor n21582 n21584 ; n21585
g21394 nor n21575 n21585 ; n21586
g21395 and asqrt[42] n21586_not ; n21587
g21396 and n20866_not n20873 ; n21588
g21397 and n20875_not n21588 ; n21589
g21398 and asqrt[5] n21589 ; n21590
g21399 nor n20866 n20875 ; n21591
g21400 and asqrt[5] n21591 ; n21592
g21401 nor n20873 n21592 ; n21593
g21402 nor n21590 n21593 ; n21594
g21403 nor asqrt[42] n21575 ; n21595
g21404 and n21585_not n21595 ; n21596
g21405 nor n21594 n21596 ; n21597
g21406 nor n21587 n21597 ; n21598
g21407 and asqrt[43] n21598_not ; n21599
g21408 and n20885 n20887_not ; n21600
g21409 and n20878_not n21600 ; n21601
g21410 and asqrt[5] n21601 ; n21602
g21411 nor n20878 n20887 ; n21603
g21412 and asqrt[5] n21603 ; n21604
g21413 nor n20885 n21604 ; n21605
g21414 nor n21602 n21605 ; n21606
g21415 nor asqrt[43] n21587 ; n21607
g21416 and n21597_not n21607 ; n21608
g21417 nor n21606 n21608 ; n21609
g21418 nor n21599 n21609 ; n21610
g21419 and asqrt[44] n21610_not ; n21611
g21420 and n20890_not n20897 ; n21612
g21421 and n20899_not n21612 ; n21613
g21422 and asqrt[5] n21613 ; n21614
g21423 nor n20890 n20899 ; n21615
g21424 and asqrt[5] n21615 ; n21616
g21425 nor n20897 n21616 ; n21617
g21426 nor n21614 n21617 ; n21618
g21427 nor asqrt[44] n21599 ; n21619
g21428 and n21609_not n21619 ; n21620
g21429 nor n21618 n21620 ; n21621
g21430 nor n21611 n21621 ; n21622
g21431 and asqrt[45] n21622_not ; n21623
g21432 and n20909 n20911_not ; n21624
g21433 and n20902_not n21624 ; n21625
g21434 and asqrt[5] n21625 ; n21626
g21435 nor n20902 n20911 ; n21627
g21436 and asqrt[5] n21627 ; n21628
g21437 nor n20909 n21628 ; n21629
g21438 nor n21626 n21629 ; n21630
g21439 nor asqrt[45] n21611 ; n21631
g21440 and n21621_not n21631 ; n21632
g21441 nor n21630 n21632 ; n21633
g21442 nor n21623 n21633 ; n21634
g21443 and asqrt[46] n21634_not ; n21635
g21444 and n20914_not n20921 ; n21636
g21445 and n20923_not n21636 ; n21637
g21446 and asqrt[5] n21637 ; n21638
g21447 nor n20914 n20923 ; n21639
g21448 and asqrt[5] n21639 ; n21640
g21449 nor n20921 n21640 ; n21641
g21450 nor n21638 n21641 ; n21642
g21451 nor asqrt[46] n21623 ; n21643
g21452 and n21633_not n21643 ; n21644
g21453 nor n21642 n21644 ; n21645
g21454 nor n21635 n21645 ; n21646
g21455 and asqrt[47] n21646_not ; n21647
g21456 and n20933 n20935_not ; n21648
g21457 and n20926_not n21648 ; n21649
g21458 and asqrt[5] n21649 ; n21650
g21459 nor n20926 n20935 ; n21651
g21460 and asqrt[5] n21651 ; n21652
g21461 nor n20933 n21652 ; n21653
g21462 nor n21650 n21653 ; n21654
g21463 nor asqrt[47] n21635 ; n21655
g21464 and n21645_not n21655 ; n21656
g21465 nor n21654 n21656 ; n21657
g21466 nor n21647 n21657 ; n21658
g21467 and asqrt[48] n21658_not ; n21659
g21468 and n20938_not n20945 ; n21660
g21469 and n20947_not n21660 ; n21661
g21470 and asqrt[5] n21661 ; n21662
g21471 nor n20938 n20947 ; n21663
g21472 and asqrt[5] n21663 ; n21664
g21473 nor n20945 n21664 ; n21665
g21474 nor n21662 n21665 ; n21666
g21475 nor asqrt[48] n21647 ; n21667
g21476 and n21657_not n21667 ; n21668
g21477 nor n21666 n21668 ; n21669
g21478 nor n21659 n21669 ; n21670
g21479 and asqrt[49] n21670_not ; n21671
g21480 and n20957 n20959_not ; n21672
g21481 and n20950_not n21672 ; n21673
g21482 and asqrt[5] n21673 ; n21674
g21483 nor n20950 n20959 ; n21675
g21484 and asqrt[5] n21675 ; n21676
g21485 nor n20957 n21676 ; n21677
g21486 nor n21674 n21677 ; n21678
g21487 nor asqrt[49] n21659 ; n21679
g21488 and n21669_not n21679 ; n21680
g21489 nor n21678 n21680 ; n21681
g21490 nor n21671 n21681 ; n21682
g21491 and asqrt[50] n21682_not ; n21683
g21492 and n20962_not n20969 ; n21684
g21493 and n20971_not n21684 ; n21685
g21494 and asqrt[5] n21685 ; n21686
g21495 nor n20962 n20971 ; n21687
g21496 and asqrt[5] n21687 ; n21688
g21497 nor n20969 n21688 ; n21689
g21498 nor n21686 n21689 ; n21690
g21499 nor asqrt[50] n21671 ; n21691
g21500 and n21681_not n21691 ; n21692
g21501 nor n21690 n21692 ; n21693
g21502 nor n21683 n21693 ; n21694
g21503 and asqrt[51] n21694_not ; n21695
g21504 and n20981 n20983_not ; n21696
g21505 and n20974_not n21696 ; n21697
g21506 and asqrt[5] n21697 ; n21698
g21507 nor n20974 n20983 ; n21699
g21508 and asqrt[5] n21699 ; n21700
g21509 nor n20981 n21700 ; n21701
g21510 nor n21698 n21701 ; n21702
g21511 nor asqrt[51] n21683 ; n21703
g21512 and n21693_not n21703 ; n21704
g21513 nor n21702 n21704 ; n21705
g21514 nor n21695 n21705 ; n21706
g21515 and asqrt[52] n21706_not ; n21707
g21516 and n20986_not n20993 ; n21708
g21517 and n20995_not n21708 ; n21709
g21518 and asqrt[5] n21709 ; n21710
g21519 nor n20986 n20995 ; n21711
g21520 and asqrt[5] n21711 ; n21712
g21521 nor n20993 n21712 ; n21713
g21522 nor n21710 n21713 ; n21714
g21523 nor asqrt[52] n21695 ; n21715
g21524 and n21705_not n21715 ; n21716
g21525 nor n21714 n21716 ; n21717
g21526 nor n21707 n21717 ; n21718
g21527 and asqrt[53] n21718_not ; n21719
g21528 and n21005 n21007_not ; n21720
g21529 and n20998_not n21720 ; n21721
g21530 and asqrt[5] n21721 ; n21722
g21531 nor n20998 n21007 ; n21723
g21532 and asqrt[5] n21723 ; n21724
g21533 nor n21005 n21724 ; n21725
g21534 nor n21722 n21725 ; n21726
g21535 nor asqrt[53] n21707 ; n21727
g21536 and n21717_not n21727 ; n21728
g21537 nor n21726 n21728 ; n21729
g21538 nor n21719 n21729 ; n21730
g21539 and asqrt[54] n21730_not ; n21731
g21540 and n21010_not n21017 ; n21732
g21541 and n21019_not n21732 ; n21733
g21542 and asqrt[5] n21733 ; n21734
g21543 nor n21010 n21019 ; n21735
g21544 and asqrt[5] n21735 ; n21736
g21545 nor n21017 n21736 ; n21737
g21546 nor n21734 n21737 ; n21738
g21547 nor asqrt[54] n21719 ; n21739
g21548 and n21729_not n21739 ; n21740
g21549 nor n21738 n21740 ; n21741
g21550 nor n21731 n21741 ; n21742
g21551 and asqrt[55] n21742_not ; n21743
g21552 and n21029 n21031_not ; n21744
g21553 and n21022_not n21744 ; n21745
g21554 and asqrt[5] n21745 ; n21746
g21555 nor n21022 n21031 ; n21747
g21556 and asqrt[5] n21747 ; n21748
g21557 nor n21029 n21748 ; n21749
g21558 nor n21746 n21749 ; n21750
g21559 nor asqrt[55] n21731 ; n21751
g21560 and n21741_not n21751 ; n21752
g21561 nor n21750 n21752 ; n21753
g21562 nor n21743 n21753 ; n21754
g21563 and asqrt[56] n21754_not ; n21755
g21564 and n21034_not n21041 ; n21756
g21565 and n21043_not n21756 ; n21757
g21566 and asqrt[5] n21757 ; n21758
g21567 nor n21034 n21043 ; n21759
g21568 and asqrt[5] n21759 ; n21760
g21569 nor n21041 n21760 ; n21761
g21570 nor n21758 n21761 ; n21762
g21571 nor asqrt[56] n21743 ; n21763
g21572 and n21753_not n21763 ; n21764
g21573 nor n21762 n21764 ; n21765
g21574 nor n21755 n21765 ; n21766
g21575 and asqrt[57] n21766_not ; n21767
g21576 and n21053 n21055_not ; n21768
g21577 and n21046_not n21768 ; n21769
g21578 and asqrt[5] n21769 ; n21770
g21579 nor n21046 n21055 ; n21771
g21580 and asqrt[5] n21771 ; n21772
g21581 nor n21053 n21772 ; n21773
g21582 nor n21770 n21773 ; n21774
g21583 nor asqrt[57] n21755 ; n21775
g21584 and n21765_not n21775 ; n21776
g21585 nor n21774 n21776 ; n21777
g21586 nor n21767 n21777 ; n21778
g21587 and asqrt[58] n21778_not ; n21779
g21588 and n21058_not n21065 ; n21780
g21589 and n21067_not n21780 ; n21781
g21590 and asqrt[5] n21781 ; n21782
g21591 nor n21058 n21067 ; n21783
g21592 and asqrt[5] n21783 ; n21784
g21593 nor n21065 n21784 ; n21785
g21594 nor n21782 n21785 ; n21786
g21595 nor asqrt[58] n21767 ; n21787
g21596 and n21777_not n21787 ; n21788
g21597 nor n21786 n21788 ; n21789
g21598 nor n21779 n21789 ; n21790
g21599 and asqrt[59] n21790_not ; n21791
g21600 and n21077 n21079_not ; n21792
g21601 and n21070_not n21792 ; n21793
g21602 and asqrt[5] n21793 ; n21794
g21603 nor n21070 n21079 ; n21795
g21604 and asqrt[5] n21795 ; n21796
g21605 nor n21077 n21796 ; n21797
g21606 nor n21794 n21797 ; n21798
g21607 nor asqrt[59] n21779 ; n21799
g21608 and n21789_not n21799 ; n21800
g21609 nor n21798 n21800 ; n21801
g21610 nor n21791 n21801 ; n21802
g21611 and asqrt[60] n21802_not ; n21803
g21612 nor asqrt[60] n21791 ; n21804
g21613 and n21801_not n21804 ; n21805
g21614 and n21082_not n21091 ; n21806
g21615 and n21084_not n21806 ; n21807
g21616 and asqrt[5] n21807 ; n21808
g21617 nor n21082 n21084 ; n21809
g21618 and asqrt[5] n21809 ; n21810
g21619 nor n21091 n21810 ; n21811
g21620 nor n21808 n21811 ; n21812
g21621 nor n21805 n21812 ; n21813
g21622 nor n21803 n21813 ; n21814
g21623 and asqrt[61] n21814_not ; n21815
g21624 and n21101 n21103_not ; n21816
g21625 and n21094_not n21816 ; n21817
g21626 and asqrt[5] n21817 ; n21818
g21627 nor n21094 n21103 ; n21819
g21628 and asqrt[5] n21819 ; n21820
g21629 nor n21101 n21820 ; n21821
g21630 nor n21818 n21821 ; n21822
g21631 nor asqrt[61] n21803 ; n21823
g21632 and n21813_not n21823 ; n21824
g21633 nor n21822 n21824 ; n21825
g21634 nor n21815 n21825 ; n21826
g21635 and asqrt[62] n21826_not ; n21827
g21636 and n21106_not n21113 ; n21828
g21637 and n21115_not n21828 ; n21829
g21638 and asqrt[5] n21829 ; n21830
g21639 nor n21106 n21115 ; n21831
g21640 and asqrt[5] n21831 ; n21832
g21641 nor n21113 n21832 ; n21833
g21642 nor n21830 n21833 ; n21834
g21643 nor asqrt[62] n21815 ; n21835
g21644 and n21825_not n21835 ; n21836
g21645 nor n21834 n21836 ; n21837
g21646 nor n21827 n21837 ; n21838
g21647 and n21125 n21127_not ; n21839
g21648 and n21118_not n21839 ; n21840
g21649 and asqrt[5] n21840 ; n21841
g21650 nor n21118 n21127 ; n21842
g21651 and asqrt[5] n21842 ; n21843
g21652 nor n21125 n21843 ; n21844
g21653 nor n21841 n21844 ; n21845
g21654 nor n21129 n21136 ; n21846
g21655 and asqrt[5] n21846 ; n21847
g21656 nor n21144 n21847 ; n21848
g21657 and n21845_not n21848 ; n21849
g21658 and n21838_not n21849 ; n21850
g21659 nor asqrt[63] n21850 ; n21851
g21660 and n21827_not n21845 ; n21852
g21661 and n21837_not n21852 ; n21853
g21662 and n21136_not asqrt[5] ; n21854
g21663 and n21129 n21854_not ; n21855
g21664 and asqrt[63] n21846_not ; n21856
g21665 and n21855_not n21856 ; n21857
g21666 nor n21853 n21857 ; n21858
g21667 nand n21851_not n21858 ; asqrt[4]
g21668 and a[8] asqrt[4] ; n21860
g21669 nor a[6] a[7] ; n21861
g21670 and a[8]_not n21861 ; n21862
g21671 nor n21860 n21862 ; n21863
g21672 and asqrt[5] n21863_not ; n21864
g21673 nor n21148 n21862 ; n21865
g21674 and n21144_not n21865 ; n21866
g21675 and n21142_not n21866 ; n21867
g21676 and n21860_not n21867 ; n21868
g21677 and a[8]_not asqrt[4] ; n21869
g21678 and a[9] n21869_not ; n21870
g21679 and n21152 asqrt[4] ; n21871
g21680 nor n21870 n21871 ; n21872
g21681 and n21868_not n21872 ; n21873
g21682 nor n21864 n21873 ; n21874
g21683 and asqrt[6] n21874_not ; n21875
g21684 nor asqrt[6] n21864 ; n21876
g21685 and n21873_not n21876 ; n21877
g21686 and asqrt[5] n21857_not ; n21878
g21687 and n21853_not n21878 ; n21879
g21688 and n21851_not n21879 ; n21880
g21689 nor n21871 n21880 ; n21881
g21690 and a[10] n21881_not ; n21882
g21691 nor a[10] n21880 ; n21883
g21692 and n21871_not n21883 ; n21884
g21693 nor n21882 n21884 ; n21885
g21694 nor n21877 n21885 ; n21886
g21695 nor n21875 n21886 ; n21887
g21696 and asqrt[7] n21887_not ; n21888
g21697 nor n21155 n21160 ; n21889
g21698 and n21164_not n21889 ; n21890
g21699 and asqrt[4] n21890 ; n21891
g21700 and asqrt[4] n21889 ; n21892
g21701 and n21164 n21892_not ; n21893
g21702 nor n21891 n21893 ; n21894
g21703 nor asqrt[7] n21875 ; n21895
g21704 and n21886_not n21895 ; n21896
g21705 nor n21894 n21896 ; n21897
g21706 nor n21888 n21897 ; n21898
g21707 and asqrt[8] n21898_not ; n21899
g21708 and n21169_not n21177 ; n21900
g21709 and n21167_not n21900 ; n21901
g21710 and asqrt[4] n21901 ; n21902
g21711 nor n21167 n21169 ; n21903
g21712 and asqrt[4] n21903 ; n21904
g21713 nor n21177 n21904 ; n21905
g21714 nor n21902 n21905 ; n21906
g21715 nor asqrt[8] n21888 ; n21907
g21716 and n21897_not n21907 ; n21908
g21717 nor n21906 n21908 ; n21909
g21718 nor n21899 n21909 ; n21910
g21719 and asqrt[9] n21910_not ; n21911
g21720 and n21180_not n21186 ; n21912
g21721 and n21188_not n21912 ; n21913
g21722 and asqrt[4] n21913 ; n21914
g21723 nor n21180 n21188 ; n21915
g21724 and asqrt[4] n21915 ; n21916
g21725 nor n21186 n21916 ; n21917
g21726 nor n21914 n21917 ; n21918
g21727 nor asqrt[9] n21899 ; n21919
g21728 and n21909_not n21919 ; n21920
g21729 nor n21918 n21920 ; n21921
g21730 nor n21911 n21921 ; n21922
g21731 and asqrt[10] n21922_not ; n21923
g21732 and n21198 n21200_not ; n21924
g21733 and n21191_not n21924 ; n21925
g21734 and asqrt[4] n21925 ; n21926
g21735 nor n21191 n21200 ; n21927
g21736 and asqrt[4] n21927 ; n21928
g21737 nor n21198 n21928 ; n21929
g21738 nor n21926 n21929 ; n21930
g21739 nor asqrt[10] n21911 ; n21931
g21740 and n21921_not n21931 ; n21932
g21741 nor n21930 n21932 ; n21933
g21742 nor n21923 n21933 ; n21934
g21743 and asqrt[11] n21934_not ; n21935
g21744 and n21203_not n21210 ; n21936
g21745 and n21212_not n21936 ; n21937
g21746 and asqrt[4] n21937 ; n21938
g21747 nor n21203 n21212 ; n21939
g21748 and asqrt[4] n21939 ; n21940
g21749 nor n21210 n21940 ; n21941
g21750 nor n21938 n21941 ; n21942
g21751 nor asqrt[11] n21923 ; n21943
g21752 and n21933_not n21943 ; n21944
g21753 nor n21942 n21944 ; n21945
g21754 nor n21935 n21945 ; n21946
g21755 and asqrt[12] n21946_not ; n21947
g21756 and n21222 n21224_not ; n21948
g21757 and n21215_not n21948 ; n21949
g21758 and asqrt[4] n21949 ; n21950
g21759 nor n21215 n21224 ; n21951
g21760 and asqrt[4] n21951 ; n21952
g21761 nor n21222 n21952 ; n21953
g21762 nor n21950 n21953 ; n21954
g21763 nor asqrt[12] n21935 ; n21955
g21764 and n21945_not n21955 ; n21956
g21765 nor n21954 n21956 ; n21957
g21766 nor n21947 n21957 ; n21958
g21767 and asqrt[13] n21958_not ; n21959
g21768 and n21227_not n21234 ; n21960
g21769 and n21236_not n21960 ; n21961
g21770 and asqrt[4] n21961 ; n21962
g21771 nor n21227 n21236 ; n21963
g21772 and asqrt[4] n21963 ; n21964
g21773 nor n21234 n21964 ; n21965
g21774 nor n21962 n21965 ; n21966
g21775 nor asqrt[13] n21947 ; n21967
g21776 and n21957_not n21967 ; n21968
g21777 nor n21966 n21968 ; n21969
g21778 nor n21959 n21969 ; n21970
g21779 and asqrt[14] n21970_not ; n21971
g21780 and n21246 n21248_not ; n21972
g21781 and n21239_not n21972 ; n21973
g21782 and asqrt[4] n21973 ; n21974
g21783 nor n21239 n21248 ; n21975
g21784 and asqrt[4] n21975 ; n21976
g21785 nor n21246 n21976 ; n21977
g21786 nor n21974 n21977 ; n21978
g21787 nor asqrt[14] n21959 ; n21979
g21788 and n21969_not n21979 ; n21980
g21789 nor n21978 n21980 ; n21981
g21790 nor n21971 n21981 ; n21982
g21791 and asqrt[15] n21982_not ; n21983
g21792 and n21251_not n21258 ; n21984
g21793 and n21260_not n21984 ; n21985
g21794 and asqrt[4] n21985 ; n21986
g21795 nor n21251 n21260 ; n21987
g21796 and asqrt[4] n21987 ; n21988
g21797 nor n21258 n21988 ; n21989
g21798 nor n21986 n21989 ; n21990
g21799 nor asqrt[15] n21971 ; n21991
g21800 and n21981_not n21991 ; n21992
g21801 nor n21990 n21992 ; n21993
g21802 nor n21983 n21993 ; n21994
g21803 and asqrt[16] n21994_not ; n21995
g21804 and n21270 n21272_not ; n21996
g21805 and n21263_not n21996 ; n21997
g21806 and asqrt[4] n21997 ; n21998
g21807 nor n21263 n21272 ; n21999
g21808 and asqrt[4] n21999 ; n22000
g21809 nor n21270 n22000 ; n22001
g21810 nor n21998 n22001 ; n22002
g21811 nor asqrt[16] n21983 ; n22003
g21812 and n21993_not n22003 ; n22004
g21813 nor n22002 n22004 ; n22005
g21814 nor n21995 n22005 ; n22006
g21815 and asqrt[17] n22006_not ; n22007
g21816 and n21275_not n21282 ; n22008
g21817 and n21284_not n22008 ; n22009
g21818 and asqrt[4] n22009 ; n22010
g21819 nor n21275 n21284 ; n22011
g21820 and asqrt[4] n22011 ; n22012
g21821 nor n21282 n22012 ; n22013
g21822 nor n22010 n22013 ; n22014
g21823 nor asqrt[17] n21995 ; n22015
g21824 and n22005_not n22015 ; n22016
g21825 nor n22014 n22016 ; n22017
g21826 nor n22007 n22017 ; n22018
g21827 and asqrt[18] n22018_not ; n22019
g21828 and n21294 n21296_not ; n22020
g21829 and n21287_not n22020 ; n22021
g21830 and asqrt[4] n22021 ; n22022
g21831 nor n21287 n21296 ; n22023
g21832 and asqrt[4] n22023 ; n22024
g21833 nor n21294 n22024 ; n22025
g21834 nor n22022 n22025 ; n22026
g21835 nor asqrt[18] n22007 ; n22027
g21836 and n22017_not n22027 ; n22028
g21837 nor n22026 n22028 ; n22029
g21838 nor n22019 n22029 ; n22030
g21839 and asqrt[19] n22030_not ; n22031
g21840 and n21299_not n21306 ; n22032
g21841 and n21308_not n22032 ; n22033
g21842 and asqrt[4] n22033 ; n22034
g21843 nor n21299 n21308 ; n22035
g21844 and asqrt[4] n22035 ; n22036
g21845 nor n21306 n22036 ; n22037
g21846 nor n22034 n22037 ; n22038
g21847 nor asqrt[19] n22019 ; n22039
g21848 and n22029_not n22039 ; n22040
g21849 nor n22038 n22040 ; n22041
g21850 nor n22031 n22041 ; n22042
g21851 and asqrt[20] n22042_not ; n22043
g21852 and n21318 n21320_not ; n22044
g21853 and n21311_not n22044 ; n22045
g21854 and asqrt[4] n22045 ; n22046
g21855 nor n21311 n21320 ; n22047
g21856 and asqrt[4] n22047 ; n22048
g21857 nor n21318 n22048 ; n22049
g21858 nor n22046 n22049 ; n22050
g21859 nor asqrt[20] n22031 ; n22051
g21860 and n22041_not n22051 ; n22052
g21861 nor n22050 n22052 ; n22053
g21862 nor n22043 n22053 ; n22054
g21863 and asqrt[21] n22054_not ; n22055
g21864 and n21323_not n21330 ; n22056
g21865 and n21332_not n22056 ; n22057
g21866 and asqrt[4] n22057 ; n22058
g21867 nor n21323 n21332 ; n22059
g21868 and asqrt[4] n22059 ; n22060
g21869 nor n21330 n22060 ; n22061
g21870 nor n22058 n22061 ; n22062
g21871 nor asqrt[21] n22043 ; n22063
g21872 and n22053_not n22063 ; n22064
g21873 nor n22062 n22064 ; n22065
g21874 nor n22055 n22065 ; n22066
g21875 and asqrt[22] n22066_not ; n22067
g21876 and n21342 n21344_not ; n22068
g21877 and n21335_not n22068 ; n22069
g21878 and asqrt[4] n22069 ; n22070
g21879 nor n21335 n21344 ; n22071
g21880 and asqrt[4] n22071 ; n22072
g21881 nor n21342 n22072 ; n22073
g21882 nor n22070 n22073 ; n22074
g21883 nor asqrt[22] n22055 ; n22075
g21884 and n22065_not n22075 ; n22076
g21885 nor n22074 n22076 ; n22077
g21886 nor n22067 n22077 ; n22078
g21887 and asqrt[23] n22078_not ; n22079
g21888 and n21347_not n21354 ; n22080
g21889 and n21356_not n22080 ; n22081
g21890 and asqrt[4] n22081 ; n22082
g21891 nor n21347 n21356 ; n22083
g21892 and asqrt[4] n22083 ; n22084
g21893 nor n21354 n22084 ; n22085
g21894 nor n22082 n22085 ; n22086
g21895 nor asqrt[23] n22067 ; n22087
g21896 and n22077_not n22087 ; n22088
g21897 nor n22086 n22088 ; n22089
g21898 nor n22079 n22089 ; n22090
g21899 and asqrt[24] n22090_not ; n22091
g21900 and n21366 n21368_not ; n22092
g21901 and n21359_not n22092 ; n22093
g21902 and asqrt[4] n22093 ; n22094
g21903 nor n21359 n21368 ; n22095
g21904 and asqrt[4] n22095 ; n22096
g21905 nor n21366 n22096 ; n22097
g21906 nor n22094 n22097 ; n22098
g21907 nor asqrt[24] n22079 ; n22099
g21908 and n22089_not n22099 ; n22100
g21909 nor n22098 n22100 ; n22101
g21910 nor n22091 n22101 ; n22102
g21911 and asqrt[25] n22102_not ; n22103
g21912 and n21371_not n21378 ; n22104
g21913 and n21380_not n22104 ; n22105
g21914 and asqrt[4] n22105 ; n22106
g21915 nor n21371 n21380 ; n22107
g21916 and asqrt[4] n22107 ; n22108
g21917 nor n21378 n22108 ; n22109
g21918 nor n22106 n22109 ; n22110
g21919 nor asqrt[25] n22091 ; n22111
g21920 and n22101_not n22111 ; n22112
g21921 nor n22110 n22112 ; n22113
g21922 nor n22103 n22113 ; n22114
g21923 and asqrt[26] n22114_not ; n22115
g21924 and n21390 n21392_not ; n22116
g21925 and n21383_not n22116 ; n22117
g21926 and asqrt[4] n22117 ; n22118
g21927 nor n21383 n21392 ; n22119
g21928 and asqrt[4] n22119 ; n22120
g21929 nor n21390 n22120 ; n22121
g21930 nor n22118 n22121 ; n22122
g21931 nor asqrt[26] n22103 ; n22123
g21932 and n22113_not n22123 ; n22124
g21933 nor n22122 n22124 ; n22125
g21934 nor n22115 n22125 ; n22126
g21935 and asqrt[27] n22126_not ; n22127
g21936 and n21395_not n21402 ; n22128
g21937 and n21404_not n22128 ; n22129
g21938 and asqrt[4] n22129 ; n22130
g21939 nor n21395 n21404 ; n22131
g21940 and asqrt[4] n22131 ; n22132
g21941 nor n21402 n22132 ; n22133
g21942 nor n22130 n22133 ; n22134
g21943 nor asqrt[27] n22115 ; n22135
g21944 and n22125_not n22135 ; n22136
g21945 nor n22134 n22136 ; n22137
g21946 nor n22127 n22137 ; n22138
g21947 and asqrt[28] n22138_not ; n22139
g21948 and n21414 n21416_not ; n22140
g21949 and n21407_not n22140 ; n22141
g21950 and asqrt[4] n22141 ; n22142
g21951 nor n21407 n21416 ; n22143
g21952 and asqrt[4] n22143 ; n22144
g21953 nor n21414 n22144 ; n22145
g21954 nor n22142 n22145 ; n22146
g21955 nor asqrt[28] n22127 ; n22147
g21956 and n22137_not n22147 ; n22148
g21957 nor n22146 n22148 ; n22149
g21958 nor n22139 n22149 ; n22150
g21959 and asqrt[29] n22150_not ; n22151
g21960 and n21419_not n21426 ; n22152
g21961 and n21428_not n22152 ; n22153
g21962 and asqrt[4] n22153 ; n22154
g21963 nor n21419 n21428 ; n22155
g21964 and asqrt[4] n22155 ; n22156
g21965 nor n21426 n22156 ; n22157
g21966 nor n22154 n22157 ; n22158
g21967 nor asqrt[29] n22139 ; n22159
g21968 and n22149_not n22159 ; n22160
g21969 nor n22158 n22160 ; n22161
g21970 nor n22151 n22161 ; n22162
g21971 and asqrt[30] n22162_not ; n22163
g21972 and n21438 n21440_not ; n22164
g21973 and n21431_not n22164 ; n22165
g21974 and asqrt[4] n22165 ; n22166
g21975 nor n21431 n21440 ; n22167
g21976 and asqrt[4] n22167 ; n22168
g21977 nor n21438 n22168 ; n22169
g21978 nor n22166 n22169 ; n22170
g21979 nor asqrt[30] n22151 ; n22171
g21980 and n22161_not n22171 ; n22172
g21981 nor n22170 n22172 ; n22173
g21982 nor n22163 n22173 ; n22174
g21983 and asqrt[31] n22174_not ; n22175
g21984 and n21443_not n21450 ; n22176
g21985 and n21452_not n22176 ; n22177
g21986 and asqrt[4] n22177 ; n22178
g21987 nor n21443 n21452 ; n22179
g21988 and asqrt[4] n22179 ; n22180
g21989 nor n21450 n22180 ; n22181
g21990 nor n22178 n22181 ; n22182
g21991 nor asqrt[31] n22163 ; n22183
g21992 and n22173_not n22183 ; n22184
g21993 nor n22182 n22184 ; n22185
g21994 nor n22175 n22185 ; n22186
g21995 and asqrt[32] n22186_not ; n22187
g21996 and n21462 n21464_not ; n22188
g21997 and n21455_not n22188 ; n22189
g21998 and asqrt[4] n22189 ; n22190
g21999 nor n21455 n21464 ; n22191
g22000 and asqrt[4] n22191 ; n22192
g22001 nor n21462 n22192 ; n22193
g22002 nor n22190 n22193 ; n22194
g22003 nor asqrt[32] n22175 ; n22195
g22004 and n22185_not n22195 ; n22196
g22005 nor n22194 n22196 ; n22197
g22006 nor n22187 n22197 ; n22198
g22007 and asqrt[33] n22198_not ; n22199
g22008 and n21467_not n21474 ; n22200
g22009 and n21476_not n22200 ; n22201
g22010 and asqrt[4] n22201 ; n22202
g22011 nor n21467 n21476 ; n22203
g22012 and asqrt[4] n22203 ; n22204
g22013 nor n21474 n22204 ; n22205
g22014 nor n22202 n22205 ; n22206
g22015 nor asqrt[33] n22187 ; n22207
g22016 and n22197_not n22207 ; n22208
g22017 nor n22206 n22208 ; n22209
g22018 nor n22199 n22209 ; n22210
g22019 and asqrt[34] n22210_not ; n22211
g22020 and n21486 n21488_not ; n22212
g22021 and n21479_not n22212 ; n22213
g22022 and asqrt[4] n22213 ; n22214
g22023 nor n21479 n21488 ; n22215
g22024 and asqrt[4] n22215 ; n22216
g22025 nor n21486 n22216 ; n22217
g22026 nor n22214 n22217 ; n22218
g22027 nor asqrt[34] n22199 ; n22219
g22028 and n22209_not n22219 ; n22220
g22029 nor n22218 n22220 ; n22221
g22030 nor n22211 n22221 ; n22222
g22031 and asqrt[35] n22222_not ; n22223
g22032 and n21491_not n21498 ; n22224
g22033 and n21500_not n22224 ; n22225
g22034 and asqrt[4] n22225 ; n22226
g22035 nor n21491 n21500 ; n22227
g22036 and asqrt[4] n22227 ; n22228
g22037 nor n21498 n22228 ; n22229
g22038 nor n22226 n22229 ; n22230
g22039 nor asqrt[35] n22211 ; n22231
g22040 and n22221_not n22231 ; n22232
g22041 nor n22230 n22232 ; n22233
g22042 nor n22223 n22233 ; n22234
g22043 and asqrt[36] n22234_not ; n22235
g22044 and n21510 n21512_not ; n22236
g22045 and n21503_not n22236 ; n22237
g22046 and asqrt[4] n22237 ; n22238
g22047 nor n21503 n21512 ; n22239
g22048 and asqrt[4] n22239 ; n22240
g22049 nor n21510 n22240 ; n22241
g22050 nor n22238 n22241 ; n22242
g22051 nor asqrt[36] n22223 ; n22243
g22052 and n22233_not n22243 ; n22244
g22053 nor n22242 n22244 ; n22245
g22054 nor n22235 n22245 ; n22246
g22055 and asqrt[37] n22246_not ; n22247
g22056 and n21515_not n21522 ; n22248
g22057 and n21524_not n22248 ; n22249
g22058 and asqrt[4] n22249 ; n22250
g22059 nor n21515 n21524 ; n22251
g22060 and asqrt[4] n22251 ; n22252
g22061 nor n21522 n22252 ; n22253
g22062 nor n22250 n22253 ; n22254
g22063 nor asqrt[37] n22235 ; n22255
g22064 and n22245_not n22255 ; n22256
g22065 nor n22254 n22256 ; n22257
g22066 nor n22247 n22257 ; n22258
g22067 and asqrt[38] n22258_not ; n22259
g22068 and n21534 n21536_not ; n22260
g22069 and n21527_not n22260 ; n22261
g22070 and asqrt[4] n22261 ; n22262
g22071 nor n21527 n21536 ; n22263
g22072 and asqrt[4] n22263 ; n22264
g22073 nor n21534 n22264 ; n22265
g22074 nor n22262 n22265 ; n22266
g22075 nor asqrt[38] n22247 ; n22267
g22076 and n22257_not n22267 ; n22268
g22077 nor n22266 n22268 ; n22269
g22078 nor n22259 n22269 ; n22270
g22079 and asqrt[39] n22270_not ; n22271
g22080 and n21539_not n21546 ; n22272
g22081 and n21548_not n22272 ; n22273
g22082 and asqrt[4] n22273 ; n22274
g22083 nor n21539 n21548 ; n22275
g22084 and asqrt[4] n22275 ; n22276
g22085 nor n21546 n22276 ; n22277
g22086 nor n22274 n22277 ; n22278
g22087 nor asqrt[39] n22259 ; n22279
g22088 and n22269_not n22279 ; n22280
g22089 nor n22278 n22280 ; n22281
g22090 nor n22271 n22281 ; n22282
g22091 and asqrt[40] n22282_not ; n22283
g22092 and n21558 n21560_not ; n22284
g22093 and n21551_not n22284 ; n22285
g22094 and asqrt[4] n22285 ; n22286
g22095 nor n21551 n21560 ; n22287
g22096 and asqrt[4] n22287 ; n22288
g22097 nor n21558 n22288 ; n22289
g22098 nor n22286 n22289 ; n22290
g22099 nor asqrt[40] n22271 ; n22291
g22100 and n22281_not n22291 ; n22292
g22101 nor n22290 n22292 ; n22293
g22102 nor n22283 n22293 ; n22294
g22103 and asqrt[41] n22294_not ; n22295
g22104 and n21563_not n21570 ; n22296
g22105 and n21572_not n22296 ; n22297
g22106 and asqrt[4] n22297 ; n22298
g22107 nor n21563 n21572 ; n22299
g22108 and asqrt[4] n22299 ; n22300
g22109 nor n21570 n22300 ; n22301
g22110 nor n22298 n22301 ; n22302
g22111 nor asqrt[41] n22283 ; n22303
g22112 and n22293_not n22303 ; n22304
g22113 nor n22302 n22304 ; n22305
g22114 nor n22295 n22305 ; n22306
g22115 and asqrt[42] n22306_not ; n22307
g22116 and n21582 n21584_not ; n22308
g22117 and n21575_not n22308 ; n22309
g22118 and asqrt[4] n22309 ; n22310
g22119 nor n21575 n21584 ; n22311
g22120 and asqrt[4] n22311 ; n22312
g22121 nor n21582 n22312 ; n22313
g22122 nor n22310 n22313 ; n22314
g22123 nor asqrt[42] n22295 ; n22315
g22124 and n22305_not n22315 ; n22316
g22125 nor n22314 n22316 ; n22317
g22126 nor n22307 n22317 ; n22318
g22127 and asqrt[43] n22318_not ; n22319
g22128 and n21587_not n21594 ; n22320
g22129 and n21596_not n22320 ; n22321
g22130 and asqrt[4] n22321 ; n22322
g22131 nor n21587 n21596 ; n22323
g22132 and asqrt[4] n22323 ; n22324
g22133 nor n21594 n22324 ; n22325
g22134 nor n22322 n22325 ; n22326
g22135 nor asqrt[43] n22307 ; n22327
g22136 and n22317_not n22327 ; n22328
g22137 nor n22326 n22328 ; n22329
g22138 nor n22319 n22329 ; n22330
g22139 and asqrt[44] n22330_not ; n22331
g22140 and n21606 n21608_not ; n22332
g22141 and n21599_not n22332 ; n22333
g22142 and asqrt[4] n22333 ; n22334
g22143 nor n21599 n21608 ; n22335
g22144 and asqrt[4] n22335 ; n22336
g22145 nor n21606 n22336 ; n22337
g22146 nor n22334 n22337 ; n22338
g22147 nor asqrt[44] n22319 ; n22339
g22148 and n22329_not n22339 ; n22340
g22149 nor n22338 n22340 ; n22341
g22150 nor n22331 n22341 ; n22342
g22151 and asqrt[45] n22342_not ; n22343
g22152 and n21611_not n21618 ; n22344
g22153 and n21620_not n22344 ; n22345
g22154 and asqrt[4] n22345 ; n22346
g22155 nor n21611 n21620 ; n22347
g22156 and asqrt[4] n22347 ; n22348
g22157 nor n21618 n22348 ; n22349
g22158 nor n22346 n22349 ; n22350
g22159 nor asqrt[45] n22331 ; n22351
g22160 and n22341_not n22351 ; n22352
g22161 nor n22350 n22352 ; n22353
g22162 nor n22343 n22353 ; n22354
g22163 and asqrt[46] n22354_not ; n22355
g22164 and n21630 n21632_not ; n22356
g22165 and n21623_not n22356 ; n22357
g22166 and asqrt[4] n22357 ; n22358
g22167 nor n21623 n21632 ; n22359
g22168 and asqrt[4] n22359 ; n22360
g22169 nor n21630 n22360 ; n22361
g22170 nor n22358 n22361 ; n22362
g22171 nor asqrt[46] n22343 ; n22363
g22172 and n22353_not n22363 ; n22364
g22173 nor n22362 n22364 ; n22365
g22174 nor n22355 n22365 ; n22366
g22175 and asqrt[47] n22366_not ; n22367
g22176 and n21635_not n21642 ; n22368
g22177 and n21644_not n22368 ; n22369
g22178 and asqrt[4] n22369 ; n22370
g22179 nor n21635 n21644 ; n22371
g22180 and asqrt[4] n22371 ; n22372
g22181 nor n21642 n22372 ; n22373
g22182 nor n22370 n22373 ; n22374
g22183 nor asqrt[47] n22355 ; n22375
g22184 and n22365_not n22375 ; n22376
g22185 nor n22374 n22376 ; n22377
g22186 nor n22367 n22377 ; n22378
g22187 and asqrt[48] n22378_not ; n22379
g22188 and n21654 n21656_not ; n22380
g22189 and n21647_not n22380 ; n22381
g22190 and asqrt[4] n22381 ; n22382
g22191 nor n21647 n21656 ; n22383
g22192 and asqrt[4] n22383 ; n22384
g22193 nor n21654 n22384 ; n22385
g22194 nor n22382 n22385 ; n22386
g22195 nor asqrt[48] n22367 ; n22387
g22196 and n22377_not n22387 ; n22388
g22197 nor n22386 n22388 ; n22389
g22198 nor n22379 n22389 ; n22390
g22199 and asqrt[49] n22390_not ; n22391
g22200 and n21659_not n21666 ; n22392
g22201 and n21668_not n22392 ; n22393
g22202 and asqrt[4] n22393 ; n22394
g22203 nor n21659 n21668 ; n22395
g22204 and asqrt[4] n22395 ; n22396
g22205 nor n21666 n22396 ; n22397
g22206 nor n22394 n22397 ; n22398
g22207 nor asqrt[49] n22379 ; n22399
g22208 and n22389_not n22399 ; n22400
g22209 nor n22398 n22400 ; n22401
g22210 nor n22391 n22401 ; n22402
g22211 and asqrt[50] n22402_not ; n22403
g22212 and n21678 n21680_not ; n22404
g22213 and n21671_not n22404 ; n22405
g22214 and asqrt[4] n22405 ; n22406
g22215 nor n21671 n21680 ; n22407
g22216 and asqrt[4] n22407 ; n22408
g22217 nor n21678 n22408 ; n22409
g22218 nor n22406 n22409 ; n22410
g22219 nor asqrt[50] n22391 ; n22411
g22220 and n22401_not n22411 ; n22412
g22221 nor n22410 n22412 ; n22413
g22222 nor n22403 n22413 ; n22414
g22223 and asqrt[51] n22414_not ; n22415
g22224 and n21683_not n21690 ; n22416
g22225 and n21692_not n22416 ; n22417
g22226 and asqrt[4] n22417 ; n22418
g22227 nor n21683 n21692 ; n22419
g22228 and asqrt[4] n22419 ; n22420
g22229 nor n21690 n22420 ; n22421
g22230 nor n22418 n22421 ; n22422
g22231 nor asqrt[51] n22403 ; n22423
g22232 and n22413_not n22423 ; n22424
g22233 nor n22422 n22424 ; n22425
g22234 nor n22415 n22425 ; n22426
g22235 and asqrt[52] n22426_not ; n22427
g22236 and n21702 n21704_not ; n22428
g22237 and n21695_not n22428 ; n22429
g22238 and asqrt[4] n22429 ; n22430
g22239 nor n21695 n21704 ; n22431
g22240 and asqrt[4] n22431 ; n22432
g22241 nor n21702 n22432 ; n22433
g22242 nor n22430 n22433 ; n22434
g22243 nor asqrt[52] n22415 ; n22435
g22244 and n22425_not n22435 ; n22436
g22245 nor n22434 n22436 ; n22437
g22246 nor n22427 n22437 ; n22438
g22247 and asqrt[53] n22438_not ; n22439
g22248 and n21707_not n21714 ; n22440
g22249 and n21716_not n22440 ; n22441
g22250 and asqrt[4] n22441 ; n22442
g22251 nor n21707 n21716 ; n22443
g22252 and asqrt[4] n22443 ; n22444
g22253 nor n21714 n22444 ; n22445
g22254 nor n22442 n22445 ; n22446
g22255 nor asqrt[53] n22427 ; n22447
g22256 and n22437_not n22447 ; n22448
g22257 nor n22446 n22448 ; n22449
g22258 nor n22439 n22449 ; n22450
g22259 and asqrt[54] n22450_not ; n22451
g22260 and n21726 n21728_not ; n22452
g22261 and n21719_not n22452 ; n22453
g22262 and asqrt[4] n22453 ; n22454
g22263 nor n21719 n21728 ; n22455
g22264 and asqrt[4] n22455 ; n22456
g22265 nor n21726 n22456 ; n22457
g22266 nor n22454 n22457 ; n22458
g22267 nor asqrt[54] n22439 ; n22459
g22268 and n22449_not n22459 ; n22460
g22269 nor n22458 n22460 ; n22461
g22270 nor n22451 n22461 ; n22462
g22271 and asqrt[55] n22462_not ; n22463
g22272 and n21731_not n21738 ; n22464
g22273 and n21740_not n22464 ; n22465
g22274 and asqrt[4] n22465 ; n22466
g22275 nor n21731 n21740 ; n22467
g22276 and asqrt[4] n22467 ; n22468
g22277 nor n21738 n22468 ; n22469
g22278 nor n22466 n22469 ; n22470
g22279 nor asqrt[55] n22451 ; n22471
g22280 and n22461_not n22471 ; n22472
g22281 nor n22470 n22472 ; n22473
g22282 nor n22463 n22473 ; n22474
g22283 and asqrt[56] n22474_not ; n22475
g22284 and n21750 n21752_not ; n22476
g22285 and n21743_not n22476 ; n22477
g22286 and asqrt[4] n22477 ; n22478
g22287 nor n21743 n21752 ; n22479
g22288 and asqrt[4] n22479 ; n22480
g22289 nor n21750 n22480 ; n22481
g22290 nor n22478 n22481 ; n22482
g22291 nor asqrt[56] n22463 ; n22483
g22292 and n22473_not n22483 ; n22484
g22293 nor n22482 n22484 ; n22485
g22294 nor n22475 n22485 ; n22486
g22295 and asqrt[57] n22486_not ; n22487
g22296 and n21755_not n21762 ; n22488
g22297 and n21764_not n22488 ; n22489
g22298 and asqrt[4] n22489 ; n22490
g22299 nor n21755 n21764 ; n22491
g22300 and asqrt[4] n22491 ; n22492
g22301 nor n21762 n22492 ; n22493
g22302 nor n22490 n22493 ; n22494
g22303 nor asqrt[57] n22475 ; n22495
g22304 and n22485_not n22495 ; n22496
g22305 nor n22494 n22496 ; n22497
g22306 nor n22487 n22497 ; n22498
g22307 and asqrt[58] n22498_not ; n22499
g22308 and n21774 n21776_not ; n22500
g22309 and n21767_not n22500 ; n22501
g22310 and asqrt[4] n22501 ; n22502
g22311 nor n21767 n21776 ; n22503
g22312 and asqrt[4] n22503 ; n22504
g22313 nor n21774 n22504 ; n22505
g22314 nor n22502 n22505 ; n22506
g22315 nor asqrt[58] n22487 ; n22507
g22316 and n22497_not n22507 ; n22508
g22317 nor n22506 n22508 ; n22509
g22318 nor n22499 n22509 ; n22510
g22319 and asqrt[59] n22510_not ; n22511
g22320 and n21779_not n21786 ; n22512
g22321 and n21788_not n22512 ; n22513
g22322 and asqrt[4] n22513 ; n22514
g22323 nor n21779 n21788 ; n22515
g22324 and asqrt[4] n22515 ; n22516
g22325 nor n21786 n22516 ; n22517
g22326 nor n22514 n22517 ; n22518
g22327 nor asqrt[59] n22499 ; n22519
g22328 and n22509_not n22519 ; n22520
g22329 nor n22518 n22520 ; n22521
g22330 nor n22511 n22521 ; n22522
g22331 and asqrt[60] n22522_not ; n22523
g22332 and n21798 n21800_not ; n22524
g22333 and n21791_not n22524 ; n22525
g22334 and asqrt[4] n22525 ; n22526
g22335 nor n21791 n21800 ; n22527
g22336 and asqrt[4] n22527 ; n22528
g22337 nor n21798 n22528 ; n22529
g22338 nor n22526 n22529 ; n22530
g22339 nor asqrt[60] n22511 ; n22531
g22340 and n22521_not n22531 ; n22532
g22341 nor n22530 n22532 ; n22533
g22342 nor n22523 n22533 ; n22534
g22343 and asqrt[61] n22534_not ; n22535
g22344 nor asqrt[61] n22523 ; n22536
g22345 and n22533_not n22536 ; n22537
g22346 and n21803_not n21812 ; n22538
g22347 and n21805_not n22538 ; n22539
g22348 and asqrt[4] n22539 ; n22540
g22349 nor n21803 n21805 ; n22541
g22350 and asqrt[4] n22541 ; n22542
g22351 nor n21812 n22542 ; n22543
g22352 nor n22540 n22543 ; n22544
g22353 nor n22537 n22544 ; n22545
g22354 nor n22535 n22545 ; n22546
g22355 and asqrt[62] n22546_not ; n22547
g22356 and n21822 n21824_not ; n22548
g22357 and n21815_not n22548 ; n22549
g22358 and asqrt[4] n22549 ; n22550
g22359 nor n21815 n21824 ; n22551
g22360 and asqrt[4] n22551 ; n22552
g22361 nor n21822 n22552 ; n22553
g22362 nor n22550 n22553 ; n22554
g22363 nor asqrt[62] n22535 ; n22555
g22364 and n22545_not n22555 ; n22556
g22365 nor n22554 n22556 ; n22557
g22366 nor n22547 n22557 ; n22558
g22367 and n21827_not n21834 ; n22559
g22368 and n21836_not n22559 ; n22560
g22369 and asqrt[4] n22560 ; n22561
g22370 nor n21827 n21836 ; n22562
g22371 and asqrt[4] n22562 ; n22563
g22372 nor n21834 n22563 ; n22564
g22373 nor n22561 n22564 ; n22565
g22374 nor n21838 n21845 ; n22566
g22375 and asqrt[4] n22566 ; n22567
g22376 nor n21853 n22567 ; n22568
g22377 and n22565_not n22568 ; n22569
g22378 and n22558_not n22569 ; n22570
g22379 nor asqrt[63] n22570 ; n22571
g22380 and n22547_not n22565 ; n22572
g22381 and n22557_not n22572 ; n22573
g22382 and n21845_not asqrt[4] ; n22574
g22383 and n21838 n22574_not ; n22575
g22384 and asqrt[63] n22566_not ; n22576
g22385 and n22575_not n22576 ; n22577
g22386 nor n22573 n22577 ; n22578
g22387 nand n22571_not n22578 ; asqrt[3]
g22388 and a[6] asqrt[3] ; n22580
g22389 nor a[4] a[5] ; n22581
g22390 and a[6]_not n22581 ; n22582
g22391 nor n22580 n22582 ; n22583
g22392 and asqrt[4] n22583_not ; n22584
g22393 nor n21857 n22582 ; n22585
g22394 and n21853_not n22585 ; n22586
g22395 and n21851_not n22586 ; n22587
g22396 and n22580_not n22587 ; n22588
g22397 and a[6]_not asqrt[3] ; n22589
g22398 and a[7] n22589_not ; n22590
g22399 and n21861 asqrt[3] ; n22591
g22400 nor n22590 n22591 ; n22592
g22401 and n22588_not n22592 ; n22593
g22402 nor n22584 n22593 ; n22594
g22403 and asqrt[5] n22594_not ; n22595
g22404 nor asqrt[5] n22584 ; n22596
g22405 and n22593_not n22596 ; n22597
g22406 and asqrt[4] n22577_not ; n22598
g22407 and n22573_not n22598 ; n22599
g22408 and n22571_not n22599 ; n22600
g22409 nor n22591 n22600 ; n22601
g22410 and a[8] n22601_not ; n22602
g22411 nor a[8] n22600 ; n22603
g22412 and n22591_not n22603 ; n22604
g22413 nor n22602 n22604 ; n22605
g22414 nor n22597 n22605 ; n22606
g22415 nor n22595 n22606 ; n22607
g22416 and asqrt[6] n22607_not ; n22608
g22417 nor n21864 n21868 ; n22609
g22418 and n21872_not n22609 ; n22610
g22419 and asqrt[3] n22610 ; n22611
g22420 and asqrt[3] n22609 ; n22612
g22421 and n21872 n22612_not ; n22613
g22422 nor n22611 n22613 ; n22614
g22423 nor asqrt[6] n22595 ; n22615
g22424 and n22606_not n22615 ; n22616
g22425 nor n22614 n22616 ; n22617
g22426 nor n22608 n22617 ; n22618
g22427 and asqrt[7] n22618_not ; n22619
g22428 and n21877_not n21885 ; n22620
g22429 and n21875_not n22620 ; n22621
g22430 and asqrt[3] n22621 ; n22622
g22431 nor n21875 n21877 ; n22623
g22432 and asqrt[3] n22623 ; n22624
g22433 nor n21885 n22624 ; n22625
g22434 nor n22622 n22625 ; n22626
g22435 nor asqrt[7] n22608 ; n22627
g22436 and n22617_not n22627 ; n22628
g22437 nor n22626 n22628 ; n22629
g22438 nor n22619 n22629 ; n22630
g22439 and asqrt[8] n22630_not ; n22631
g22440 and n21888_not n21894 ; n22632
g22441 and n21896_not n22632 ; n22633
g22442 and asqrt[3] n22633 ; n22634
g22443 nor n21888 n21896 ; n22635
g22444 and asqrt[3] n22635 ; n22636
g22445 nor n21894 n22636 ; n22637
g22446 nor n22634 n22637 ; n22638
g22447 nor asqrt[8] n22619 ; n22639
g22448 and n22629_not n22639 ; n22640
g22449 nor n22638 n22640 ; n22641
g22450 nor n22631 n22641 ; n22642
g22451 and asqrt[9] n22642_not ; n22643
g22452 and n21906 n21908_not ; n22644
g22453 and n21899_not n22644 ; n22645
g22454 and asqrt[3] n22645 ; n22646
g22455 nor n21899 n21908 ; n22647
g22456 and asqrt[3] n22647 ; n22648
g22457 nor n21906 n22648 ; n22649
g22458 nor n22646 n22649 ; n22650
g22459 nor asqrt[9] n22631 ; n22651
g22460 and n22641_not n22651 ; n22652
g22461 nor n22650 n22652 ; n22653
g22462 nor n22643 n22653 ; n22654
g22463 and asqrt[10] n22654_not ; n22655
g22464 and n21911_not n21918 ; n22656
g22465 and n21920_not n22656 ; n22657
g22466 and asqrt[3] n22657 ; n22658
g22467 nor n21911 n21920 ; n22659
g22468 and asqrt[3] n22659 ; n22660
g22469 nor n21918 n22660 ; n22661
g22470 nor n22658 n22661 ; n22662
g22471 nor asqrt[10] n22643 ; n22663
g22472 and n22653_not n22663 ; n22664
g22473 nor n22662 n22664 ; n22665
g22474 nor n22655 n22665 ; n22666
g22475 and asqrt[11] n22666_not ; n22667
g22476 and n21930 n21932_not ; n22668
g22477 and n21923_not n22668 ; n22669
g22478 and asqrt[3] n22669 ; n22670
g22479 nor n21923 n21932 ; n22671
g22480 and asqrt[3] n22671 ; n22672
g22481 nor n21930 n22672 ; n22673
g22482 nor n22670 n22673 ; n22674
g22483 nor asqrt[11] n22655 ; n22675
g22484 and n22665_not n22675 ; n22676
g22485 nor n22674 n22676 ; n22677
g22486 nor n22667 n22677 ; n22678
g22487 and asqrt[12] n22678_not ; n22679
g22488 and n21935_not n21942 ; n22680
g22489 and n21944_not n22680 ; n22681
g22490 and asqrt[3] n22681 ; n22682
g22491 nor n21935 n21944 ; n22683
g22492 and asqrt[3] n22683 ; n22684
g22493 nor n21942 n22684 ; n22685
g22494 nor n22682 n22685 ; n22686
g22495 nor asqrt[12] n22667 ; n22687
g22496 and n22677_not n22687 ; n22688
g22497 nor n22686 n22688 ; n22689
g22498 nor n22679 n22689 ; n22690
g22499 and asqrt[13] n22690_not ; n22691
g22500 and n21954 n21956_not ; n22692
g22501 and n21947_not n22692 ; n22693
g22502 and asqrt[3] n22693 ; n22694
g22503 nor n21947 n21956 ; n22695
g22504 and asqrt[3] n22695 ; n22696
g22505 nor n21954 n22696 ; n22697
g22506 nor n22694 n22697 ; n22698
g22507 nor asqrt[13] n22679 ; n22699
g22508 and n22689_not n22699 ; n22700
g22509 nor n22698 n22700 ; n22701
g22510 nor n22691 n22701 ; n22702
g22511 and asqrt[14] n22702_not ; n22703
g22512 and n21959_not n21966 ; n22704
g22513 and n21968_not n22704 ; n22705
g22514 and asqrt[3] n22705 ; n22706
g22515 nor n21959 n21968 ; n22707
g22516 and asqrt[3] n22707 ; n22708
g22517 nor n21966 n22708 ; n22709
g22518 nor n22706 n22709 ; n22710
g22519 nor asqrt[14] n22691 ; n22711
g22520 and n22701_not n22711 ; n22712
g22521 nor n22710 n22712 ; n22713
g22522 nor n22703 n22713 ; n22714
g22523 and asqrt[15] n22714_not ; n22715
g22524 and n21978 n21980_not ; n22716
g22525 and n21971_not n22716 ; n22717
g22526 and asqrt[3] n22717 ; n22718
g22527 nor n21971 n21980 ; n22719
g22528 and asqrt[3] n22719 ; n22720
g22529 nor n21978 n22720 ; n22721
g22530 nor n22718 n22721 ; n22722
g22531 nor asqrt[15] n22703 ; n22723
g22532 and n22713_not n22723 ; n22724
g22533 nor n22722 n22724 ; n22725
g22534 nor n22715 n22725 ; n22726
g22535 and asqrt[16] n22726_not ; n22727
g22536 and n21983_not n21990 ; n22728
g22537 and n21992_not n22728 ; n22729
g22538 and asqrt[3] n22729 ; n22730
g22539 nor n21983 n21992 ; n22731
g22540 and asqrt[3] n22731 ; n22732
g22541 nor n21990 n22732 ; n22733
g22542 nor n22730 n22733 ; n22734
g22543 nor asqrt[16] n22715 ; n22735
g22544 and n22725_not n22735 ; n22736
g22545 nor n22734 n22736 ; n22737
g22546 nor n22727 n22737 ; n22738
g22547 and asqrt[17] n22738_not ; n22739
g22548 and n22002 n22004_not ; n22740
g22549 and n21995_not n22740 ; n22741
g22550 and asqrt[3] n22741 ; n22742
g22551 nor n21995 n22004 ; n22743
g22552 and asqrt[3] n22743 ; n22744
g22553 nor n22002 n22744 ; n22745
g22554 nor n22742 n22745 ; n22746
g22555 nor asqrt[17] n22727 ; n22747
g22556 and n22737_not n22747 ; n22748
g22557 nor n22746 n22748 ; n22749
g22558 nor n22739 n22749 ; n22750
g22559 and asqrt[18] n22750_not ; n22751
g22560 and n22007_not n22014 ; n22752
g22561 and n22016_not n22752 ; n22753
g22562 and asqrt[3] n22753 ; n22754
g22563 nor n22007 n22016 ; n22755
g22564 and asqrt[3] n22755 ; n22756
g22565 nor n22014 n22756 ; n22757
g22566 nor n22754 n22757 ; n22758
g22567 nor asqrt[18] n22739 ; n22759
g22568 and n22749_not n22759 ; n22760
g22569 nor n22758 n22760 ; n22761
g22570 nor n22751 n22761 ; n22762
g22571 and asqrt[19] n22762_not ; n22763
g22572 and n22026 n22028_not ; n22764
g22573 and n22019_not n22764 ; n22765
g22574 and asqrt[3] n22765 ; n22766
g22575 nor n22019 n22028 ; n22767
g22576 and asqrt[3] n22767 ; n22768
g22577 nor n22026 n22768 ; n22769
g22578 nor n22766 n22769 ; n22770
g22579 nor asqrt[19] n22751 ; n22771
g22580 and n22761_not n22771 ; n22772
g22581 nor n22770 n22772 ; n22773
g22582 nor n22763 n22773 ; n22774
g22583 and asqrt[20] n22774_not ; n22775
g22584 and n22031_not n22038 ; n22776
g22585 and n22040_not n22776 ; n22777
g22586 and asqrt[3] n22777 ; n22778
g22587 nor n22031 n22040 ; n22779
g22588 and asqrt[3] n22779 ; n22780
g22589 nor n22038 n22780 ; n22781
g22590 nor n22778 n22781 ; n22782
g22591 nor asqrt[20] n22763 ; n22783
g22592 and n22773_not n22783 ; n22784
g22593 nor n22782 n22784 ; n22785
g22594 nor n22775 n22785 ; n22786
g22595 and asqrt[21] n22786_not ; n22787
g22596 and n22050 n22052_not ; n22788
g22597 and n22043_not n22788 ; n22789
g22598 and asqrt[3] n22789 ; n22790
g22599 nor n22043 n22052 ; n22791
g22600 and asqrt[3] n22791 ; n22792
g22601 nor n22050 n22792 ; n22793
g22602 nor n22790 n22793 ; n22794
g22603 nor asqrt[21] n22775 ; n22795
g22604 and n22785_not n22795 ; n22796
g22605 nor n22794 n22796 ; n22797
g22606 nor n22787 n22797 ; n22798
g22607 and asqrt[22] n22798_not ; n22799
g22608 and n22055_not n22062 ; n22800
g22609 and n22064_not n22800 ; n22801
g22610 and asqrt[3] n22801 ; n22802
g22611 nor n22055 n22064 ; n22803
g22612 and asqrt[3] n22803 ; n22804
g22613 nor n22062 n22804 ; n22805
g22614 nor n22802 n22805 ; n22806
g22615 nor asqrt[22] n22787 ; n22807
g22616 and n22797_not n22807 ; n22808
g22617 nor n22806 n22808 ; n22809
g22618 nor n22799 n22809 ; n22810
g22619 and asqrt[23] n22810_not ; n22811
g22620 and n22074 n22076_not ; n22812
g22621 and n22067_not n22812 ; n22813
g22622 and asqrt[3] n22813 ; n22814
g22623 nor n22067 n22076 ; n22815
g22624 and asqrt[3] n22815 ; n22816
g22625 nor n22074 n22816 ; n22817
g22626 nor n22814 n22817 ; n22818
g22627 nor asqrt[23] n22799 ; n22819
g22628 and n22809_not n22819 ; n22820
g22629 nor n22818 n22820 ; n22821
g22630 nor n22811 n22821 ; n22822
g22631 and asqrt[24] n22822_not ; n22823
g22632 and n22079_not n22086 ; n22824
g22633 and n22088_not n22824 ; n22825
g22634 and asqrt[3] n22825 ; n22826
g22635 nor n22079 n22088 ; n22827
g22636 and asqrt[3] n22827 ; n22828
g22637 nor n22086 n22828 ; n22829
g22638 nor n22826 n22829 ; n22830
g22639 nor asqrt[24] n22811 ; n22831
g22640 and n22821_not n22831 ; n22832
g22641 nor n22830 n22832 ; n22833
g22642 nor n22823 n22833 ; n22834
g22643 and asqrt[25] n22834_not ; n22835
g22644 and n22098 n22100_not ; n22836
g22645 and n22091_not n22836 ; n22837
g22646 and asqrt[3] n22837 ; n22838
g22647 nor n22091 n22100 ; n22839
g22648 and asqrt[3] n22839 ; n22840
g22649 nor n22098 n22840 ; n22841
g22650 nor n22838 n22841 ; n22842
g22651 nor asqrt[25] n22823 ; n22843
g22652 and n22833_not n22843 ; n22844
g22653 nor n22842 n22844 ; n22845
g22654 nor n22835 n22845 ; n22846
g22655 and asqrt[26] n22846_not ; n22847
g22656 and n22103_not n22110 ; n22848
g22657 and n22112_not n22848 ; n22849
g22658 and asqrt[3] n22849 ; n22850
g22659 nor n22103 n22112 ; n22851
g22660 and asqrt[3] n22851 ; n22852
g22661 nor n22110 n22852 ; n22853
g22662 nor n22850 n22853 ; n22854
g22663 nor asqrt[26] n22835 ; n22855
g22664 and n22845_not n22855 ; n22856
g22665 nor n22854 n22856 ; n22857
g22666 nor n22847 n22857 ; n22858
g22667 and asqrt[27] n22858_not ; n22859
g22668 and n22122 n22124_not ; n22860
g22669 and n22115_not n22860 ; n22861
g22670 and asqrt[3] n22861 ; n22862
g22671 nor n22115 n22124 ; n22863
g22672 and asqrt[3] n22863 ; n22864
g22673 nor n22122 n22864 ; n22865
g22674 nor n22862 n22865 ; n22866
g22675 nor asqrt[27] n22847 ; n22867
g22676 and n22857_not n22867 ; n22868
g22677 nor n22866 n22868 ; n22869
g22678 nor n22859 n22869 ; n22870
g22679 and asqrt[28] n22870_not ; n22871
g22680 and n22127_not n22134 ; n22872
g22681 and n22136_not n22872 ; n22873
g22682 and asqrt[3] n22873 ; n22874
g22683 nor n22127 n22136 ; n22875
g22684 and asqrt[3] n22875 ; n22876
g22685 nor n22134 n22876 ; n22877
g22686 nor n22874 n22877 ; n22878
g22687 nor asqrt[28] n22859 ; n22879
g22688 and n22869_not n22879 ; n22880
g22689 nor n22878 n22880 ; n22881
g22690 nor n22871 n22881 ; n22882
g22691 and asqrt[29] n22882_not ; n22883
g22692 and n22146 n22148_not ; n22884
g22693 and n22139_not n22884 ; n22885
g22694 and asqrt[3] n22885 ; n22886
g22695 nor n22139 n22148 ; n22887
g22696 and asqrt[3] n22887 ; n22888
g22697 nor n22146 n22888 ; n22889
g22698 nor n22886 n22889 ; n22890
g22699 nor asqrt[29] n22871 ; n22891
g22700 and n22881_not n22891 ; n22892
g22701 nor n22890 n22892 ; n22893
g22702 nor n22883 n22893 ; n22894
g22703 and asqrt[30] n22894_not ; n22895
g22704 and n22151_not n22158 ; n22896
g22705 and n22160_not n22896 ; n22897
g22706 and asqrt[3] n22897 ; n22898
g22707 nor n22151 n22160 ; n22899
g22708 and asqrt[3] n22899 ; n22900
g22709 nor n22158 n22900 ; n22901
g22710 nor n22898 n22901 ; n22902
g22711 nor asqrt[30] n22883 ; n22903
g22712 and n22893_not n22903 ; n22904
g22713 nor n22902 n22904 ; n22905
g22714 nor n22895 n22905 ; n22906
g22715 and asqrt[31] n22906_not ; n22907
g22716 and n22170 n22172_not ; n22908
g22717 and n22163_not n22908 ; n22909
g22718 and asqrt[3] n22909 ; n22910
g22719 nor n22163 n22172 ; n22911
g22720 and asqrt[3] n22911 ; n22912
g22721 nor n22170 n22912 ; n22913
g22722 nor n22910 n22913 ; n22914
g22723 nor asqrt[31] n22895 ; n22915
g22724 and n22905_not n22915 ; n22916
g22725 nor n22914 n22916 ; n22917
g22726 nor n22907 n22917 ; n22918
g22727 and asqrt[32] n22918_not ; n22919
g22728 and n22175_not n22182 ; n22920
g22729 and n22184_not n22920 ; n22921
g22730 and asqrt[3] n22921 ; n22922
g22731 nor n22175 n22184 ; n22923
g22732 and asqrt[3] n22923 ; n22924
g22733 nor n22182 n22924 ; n22925
g22734 nor n22922 n22925 ; n22926
g22735 nor asqrt[32] n22907 ; n22927
g22736 and n22917_not n22927 ; n22928
g22737 nor n22926 n22928 ; n22929
g22738 nor n22919 n22929 ; n22930
g22739 and asqrt[33] n22930_not ; n22931
g22740 and n22194 n22196_not ; n22932
g22741 and n22187_not n22932 ; n22933
g22742 and asqrt[3] n22933 ; n22934
g22743 nor n22187 n22196 ; n22935
g22744 and asqrt[3] n22935 ; n22936
g22745 nor n22194 n22936 ; n22937
g22746 nor n22934 n22937 ; n22938
g22747 nor asqrt[33] n22919 ; n22939
g22748 and n22929_not n22939 ; n22940
g22749 nor n22938 n22940 ; n22941
g22750 nor n22931 n22941 ; n22942
g22751 and asqrt[34] n22942_not ; n22943
g22752 and n22199_not n22206 ; n22944
g22753 and n22208_not n22944 ; n22945
g22754 and asqrt[3] n22945 ; n22946
g22755 nor n22199 n22208 ; n22947
g22756 and asqrt[3] n22947 ; n22948
g22757 nor n22206 n22948 ; n22949
g22758 nor n22946 n22949 ; n22950
g22759 nor asqrt[34] n22931 ; n22951
g22760 and n22941_not n22951 ; n22952
g22761 nor n22950 n22952 ; n22953
g22762 nor n22943 n22953 ; n22954
g22763 and asqrt[35] n22954_not ; n22955
g22764 and n22218 n22220_not ; n22956
g22765 and n22211_not n22956 ; n22957
g22766 and asqrt[3] n22957 ; n22958
g22767 nor n22211 n22220 ; n22959
g22768 and asqrt[3] n22959 ; n22960
g22769 nor n22218 n22960 ; n22961
g22770 nor n22958 n22961 ; n22962
g22771 nor asqrt[35] n22943 ; n22963
g22772 and n22953_not n22963 ; n22964
g22773 nor n22962 n22964 ; n22965
g22774 nor n22955 n22965 ; n22966
g22775 and asqrt[36] n22966_not ; n22967
g22776 and n22223_not n22230 ; n22968
g22777 and n22232_not n22968 ; n22969
g22778 and asqrt[3] n22969 ; n22970
g22779 nor n22223 n22232 ; n22971
g22780 and asqrt[3] n22971 ; n22972
g22781 nor n22230 n22972 ; n22973
g22782 nor n22970 n22973 ; n22974
g22783 nor asqrt[36] n22955 ; n22975
g22784 and n22965_not n22975 ; n22976
g22785 nor n22974 n22976 ; n22977
g22786 nor n22967 n22977 ; n22978
g22787 and asqrt[37] n22978_not ; n22979
g22788 and n22242 n22244_not ; n22980
g22789 and n22235_not n22980 ; n22981
g22790 and asqrt[3] n22981 ; n22982
g22791 nor n22235 n22244 ; n22983
g22792 and asqrt[3] n22983 ; n22984
g22793 nor n22242 n22984 ; n22985
g22794 nor n22982 n22985 ; n22986
g22795 nor asqrt[37] n22967 ; n22987
g22796 and n22977_not n22987 ; n22988
g22797 nor n22986 n22988 ; n22989
g22798 nor n22979 n22989 ; n22990
g22799 and asqrt[38] n22990_not ; n22991
g22800 and n22247_not n22254 ; n22992
g22801 and n22256_not n22992 ; n22993
g22802 and asqrt[3] n22993 ; n22994
g22803 nor n22247 n22256 ; n22995
g22804 and asqrt[3] n22995 ; n22996
g22805 nor n22254 n22996 ; n22997
g22806 nor n22994 n22997 ; n22998
g22807 nor asqrt[38] n22979 ; n22999
g22808 and n22989_not n22999 ; n23000
g22809 nor n22998 n23000 ; n23001
g22810 nor n22991 n23001 ; n23002
g22811 and asqrt[39] n23002_not ; n23003
g22812 and n22266 n22268_not ; n23004
g22813 and n22259_not n23004 ; n23005
g22814 and asqrt[3] n23005 ; n23006
g22815 nor n22259 n22268 ; n23007
g22816 and asqrt[3] n23007 ; n23008
g22817 nor n22266 n23008 ; n23009
g22818 nor n23006 n23009 ; n23010
g22819 nor asqrt[39] n22991 ; n23011
g22820 and n23001_not n23011 ; n23012
g22821 nor n23010 n23012 ; n23013
g22822 nor n23003 n23013 ; n23014
g22823 and asqrt[40] n23014_not ; n23015
g22824 and n22271_not n22278 ; n23016
g22825 and n22280_not n23016 ; n23017
g22826 and asqrt[3] n23017 ; n23018
g22827 nor n22271 n22280 ; n23019
g22828 and asqrt[3] n23019 ; n23020
g22829 nor n22278 n23020 ; n23021
g22830 nor n23018 n23021 ; n23022
g22831 nor asqrt[40] n23003 ; n23023
g22832 and n23013_not n23023 ; n23024
g22833 nor n23022 n23024 ; n23025
g22834 nor n23015 n23025 ; n23026
g22835 and asqrt[41] n23026_not ; n23027
g22836 and n22290 n22292_not ; n23028
g22837 and n22283_not n23028 ; n23029
g22838 and asqrt[3] n23029 ; n23030
g22839 nor n22283 n22292 ; n23031
g22840 and asqrt[3] n23031 ; n23032
g22841 nor n22290 n23032 ; n23033
g22842 nor n23030 n23033 ; n23034
g22843 nor asqrt[41] n23015 ; n23035
g22844 and n23025_not n23035 ; n23036
g22845 nor n23034 n23036 ; n23037
g22846 nor n23027 n23037 ; n23038
g22847 and asqrt[42] n23038_not ; n23039
g22848 and n22295_not n22302 ; n23040
g22849 and n22304_not n23040 ; n23041
g22850 and asqrt[3] n23041 ; n23042
g22851 nor n22295 n22304 ; n23043
g22852 and asqrt[3] n23043 ; n23044
g22853 nor n22302 n23044 ; n23045
g22854 nor n23042 n23045 ; n23046
g22855 nor asqrt[42] n23027 ; n23047
g22856 and n23037_not n23047 ; n23048
g22857 nor n23046 n23048 ; n23049
g22858 nor n23039 n23049 ; n23050
g22859 and asqrt[43] n23050_not ; n23051
g22860 and n22314 n22316_not ; n23052
g22861 and n22307_not n23052 ; n23053
g22862 and asqrt[3] n23053 ; n23054
g22863 nor n22307 n22316 ; n23055
g22864 and asqrt[3] n23055 ; n23056
g22865 nor n22314 n23056 ; n23057
g22866 nor n23054 n23057 ; n23058
g22867 nor asqrt[43] n23039 ; n23059
g22868 and n23049_not n23059 ; n23060
g22869 nor n23058 n23060 ; n23061
g22870 nor n23051 n23061 ; n23062
g22871 and asqrt[44] n23062_not ; n23063
g22872 and n22319_not n22326 ; n23064
g22873 and n22328_not n23064 ; n23065
g22874 and asqrt[3] n23065 ; n23066
g22875 nor n22319 n22328 ; n23067
g22876 and asqrt[3] n23067 ; n23068
g22877 nor n22326 n23068 ; n23069
g22878 nor n23066 n23069 ; n23070
g22879 nor asqrt[44] n23051 ; n23071
g22880 and n23061_not n23071 ; n23072
g22881 nor n23070 n23072 ; n23073
g22882 nor n23063 n23073 ; n23074
g22883 and asqrt[45] n23074_not ; n23075
g22884 and n22338 n22340_not ; n23076
g22885 and n22331_not n23076 ; n23077
g22886 and asqrt[3] n23077 ; n23078
g22887 nor n22331 n22340 ; n23079
g22888 and asqrt[3] n23079 ; n23080
g22889 nor n22338 n23080 ; n23081
g22890 nor n23078 n23081 ; n23082
g22891 nor asqrt[45] n23063 ; n23083
g22892 and n23073_not n23083 ; n23084
g22893 nor n23082 n23084 ; n23085
g22894 nor n23075 n23085 ; n23086
g22895 and asqrt[46] n23086_not ; n23087
g22896 and n22343_not n22350 ; n23088
g22897 and n22352_not n23088 ; n23089
g22898 and asqrt[3] n23089 ; n23090
g22899 nor n22343 n22352 ; n23091
g22900 and asqrt[3] n23091 ; n23092
g22901 nor n22350 n23092 ; n23093
g22902 nor n23090 n23093 ; n23094
g22903 nor asqrt[46] n23075 ; n23095
g22904 and n23085_not n23095 ; n23096
g22905 nor n23094 n23096 ; n23097
g22906 nor n23087 n23097 ; n23098
g22907 and asqrt[47] n23098_not ; n23099
g22908 and n22362 n22364_not ; n23100
g22909 and n22355_not n23100 ; n23101
g22910 and asqrt[3] n23101 ; n23102
g22911 nor n22355 n22364 ; n23103
g22912 and asqrt[3] n23103 ; n23104
g22913 nor n22362 n23104 ; n23105
g22914 nor n23102 n23105 ; n23106
g22915 nor asqrt[47] n23087 ; n23107
g22916 and n23097_not n23107 ; n23108
g22917 nor n23106 n23108 ; n23109
g22918 nor n23099 n23109 ; n23110
g22919 and asqrt[48] n23110_not ; n23111
g22920 and n22367_not n22374 ; n23112
g22921 and n22376_not n23112 ; n23113
g22922 and asqrt[3] n23113 ; n23114
g22923 nor n22367 n22376 ; n23115
g22924 and asqrt[3] n23115 ; n23116
g22925 nor n22374 n23116 ; n23117
g22926 nor n23114 n23117 ; n23118
g22927 nor asqrt[48] n23099 ; n23119
g22928 and n23109_not n23119 ; n23120
g22929 nor n23118 n23120 ; n23121
g22930 nor n23111 n23121 ; n23122
g22931 and asqrt[49] n23122_not ; n23123
g22932 and n22386 n22388_not ; n23124
g22933 and n22379_not n23124 ; n23125
g22934 and asqrt[3] n23125 ; n23126
g22935 nor n22379 n22388 ; n23127
g22936 and asqrt[3] n23127 ; n23128
g22937 nor n22386 n23128 ; n23129
g22938 nor n23126 n23129 ; n23130
g22939 nor asqrt[49] n23111 ; n23131
g22940 and n23121_not n23131 ; n23132
g22941 nor n23130 n23132 ; n23133
g22942 nor n23123 n23133 ; n23134
g22943 and asqrt[50] n23134_not ; n23135
g22944 and n22391_not n22398 ; n23136
g22945 and n22400_not n23136 ; n23137
g22946 and asqrt[3] n23137 ; n23138
g22947 nor n22391 n22400 ; n23139
g22948 and asqrt[3] n23139 ; n23140
g22949 nor n22398 n23140 ; n23141
g22950 nor n23138 n23141 ; n23142
g22951 nor asqrt[50] n23123 ; n23143
g22952 and n23133_not n23143 ; n23144
g22953 nor n23142 n23144 ; n23145
g22954 nor n23135 n23145 ; n23146
g22955 and asqrt[51] n23146_not ; n23147
g22956 and n22410 n22412_not ; n23148
g22957 and n22403_not n23148 ; n23149
g22958 and asqrt[3] n23149 ; n23150
g22959 nor n22403 n22412 ; n23151
g22960 and asqrt[3] n23151 ; n23152
g22961 nor n22410 n23152 ; n23153
g22962 nor n23150 n23153 ; n23154
g22963 nor asqrt[51] n23135 ; n23155
g22964 and n23145_not n23155 ; n23156
g22965 nor n23154 n23156 ; n23157
g22966 nor n23147 n23157 ; n23158
g22967 and asqrt[52] n23158_not ; n23159
g22968 and n22415_not n22422 ; n23160
g22969 and n22424_not n23160 ; n23161
g22970 and asqrt[3] n23161 ; n23162
g22971 nor n22415 n22424 ; n23163
g22972 and asqrt[3] n23163 ; n23164
g22973 nor n22422 n23164 ; n23165
g22974 nor n23162 n23165 ; n23166
g22975 nor asqrt[52] n23147 ; n23167
g22976 and n23157_not n23167 ; n23168
g22977 nor n23166 n23168 ; n23169
g22978 nor n23159 n23169 ; n23170
g22979 and asqrt[53] n23170_not ; n23171
g22980 and n22434 n22436_not ; n23172
g22981 and n22427_not n23172 ; n23173
g22982 and asqrt[3] n23173 ; n23174
g22983 nor n22427 n22436 ; n23175
g22984 and asqrt[3] n23175 ; n23176
g22985 nor n22434 n23176 ; n23177
g22986 nor n23174 n23177 ; n23178
g22987 nor asqrt[53] n23159 ; n23179
g22988 and n23169_not n23179 ; n23180
g22989 nor n23178 n23180 ; n23181
g22990 nor n23171 n23181 ; n23182
g22991 and asqrt[54] n23182_not ; n23183
g22992 and n22439_not n22446 ; n23184
g22993 and n22448_not n23184 ; n23185
g22994 and asqrt[3] n23185 ; n23186
g22995 nor n22439 n22448 ; n23187
g22996 and asqrt[3] n23187 ; n23188
g22997 nor n22446 n23188 ; n23189
g22998 nor n23186 n23189 ; n23190
g22999 nor asqrt[54] n23171 ; n23191
g23000 and n23181_not n23191 ; n23192
g23001 nor n23190 n23192 ; n23193
g23002 nor n23183 n23193 ; n23194
g23003 and asqrt[55] n23194_not ; n23195
g23004 and n22458 n22460_not ; n23196
g23005 and n22451_not n23196 ; n23197
g23006 and asqrt[3] n23197 ; n23198
g23007 nor n22451 n22460 ; n23199
g23008 and asqrt[3] n23199 ; n23200
g23009 nor n22458 n23200 ; n23201
g23010 nor n23198 n23201 ; n23202
g23011 nor asqrt[55] n23183 ; n23203
g23012 and n23193_not n23203 ; n23204
g23013 nor n23202 n23204 ; n23205
g23014 nor n23195 n23205 ; n23206
g23015 and asqrt[56] n23206_not ; n23207
g23016 and n22463_not n22470 ; n23208
g23017 and n22472_not n23208 ; n23209
g23018 and asqrt[3] n23209 ; n23210
g23019 nor n22463 n22472 ; n23211
g23020 and asqrt[3] n23211 ; n23212
g23021 nor n22470 n23212 ; n23213
g23022 nor n23210 n23213 ; n23214
g23023 nor asqrt[56] n23195 ; n23215
g23024 and n23205_not n23215 ; n23216
g23025 nor n23214 n23216 ; n23217
g23026 nor n23207 n23217 ; n23218
g23027 and asqrt[57] n23218_not ; n23219
g23028 and n22482 n22484_not ; n23220
g23029 and n22475_not n23220 ; n23221
g23030 and asqrt[3] n23221 ; n23222
g23031 nor n22475 n22484 ; n23223
g23032 and asqrt[3] n23223 ; n23224
g23033 nor n22482 n23224 ; n23225
g23034 nor n23222 n23225 ; n23226
g23035 nor asqrt[57] n23207 ; n23227
g23036 and n23217_not n23227 ; n23228
g23037 nor n23226 n23228 ; n23229
g23038 nor n23219 n23229 ; n23230
g23039 and asqrt[58] n23230_not ; n23231
g23040 and n22487_not n22494 ; n23232
g23041 and n22496_not n23232 ; n23233
g23042 and asqrt[3] n23233 ; n23234
g23043 nor n22487 n22496 ; n23235
g23044 and asqrt[3] n23235 ; n23236
g23045 nor n22494 n23236 ; n23237
g23046 nor n23234 n23237 ; n23238
g23047 nor asqrt[58] n23219 ; n23239
g23048 and n23229_not n23239 ; n23240
g23049 nor n23238 n23240 ; n23241
g23050 nor n23231 n23241 ; n23242
g23051 and asqrt[59] n23242_not ; n23243
g23052 and n22506 n22508_not ; n23244
g23053 and n22499_not n23244 ; n23245
g23054 and asqrt[3] n23245 ; n23246
g23055 nor n22499 n22508 ; n23247
g23056 and asqrt[3] n23247 ; n23248
g23057 nor n22506 n23248 ; n23249
g23058 nor n23246 n23249 ; n23250
g23059 nor asqrt[59] n23231 ; n23251
g23060 and n23241_not n23251 ; n23252
g23061 nor n23250 n23252 ; n23253
g23062 nor n23243 n23253 ; n23254
g23063 and asqrt[60] n23254_not ; n23255
g23064 and n22511_not n22518 ; n23256
g23065 and n22520_not n23256 ; n23257
g23066 and asqrt[3] n23257 ; n23258
g23067 nor n22511 n22520 ; n23259
g23068 and asqrt[3] n23259 ; n23260
g23069 nor n22518 n23260 ; n23261
g23070 nor n23258 n23261 ; n23262
g23071 nor asqrt[60] n23243 ; n23263
g23072 and n23253_not n23263 ; n23264
g23073 nor n23262 n23264 ; n23265
g23074 nor n23255 n23265 ; n23266
g23075 and asqrt[61] n23266_not ; n23267
g23076 and n22530 n22532_not ; n23268
g23077 and n22523_not n23268 ; n23269
g23078 and asqrt[3] n23269 ; n23270
g23079 nor n22523 n22532 ; n23271
g23080 and asqrt[3] n23271 ; n23272
g23081 nor n22530 n23272 ; n23273
g23082 nor n23270 n23273 ; n23274
g23083 nor asqrt[61] n23255 ; n23275
g23084 and n23265_not n23275 ; n23276
g23085 nor n23274 n23276 ; n23277
g23086 nor n23267 n23277 ; n23278
g23087 and asqrt[62] n23278_not ; n23279
g23088 nor asqrt[62] n23267 ; n23280
g23089 and n23277_not n23280 ; n23281
g23090 and n22535_not n22544 ; n23282
g23091 and n22537_not n23282 ; n23283
g23092 and asqrt[3] n23283 ; n23284
g23093 nor n22535 n22537 ; n23285
g23094 and asqrt[3] n23285 ; n23286
g23095 nor n22544 n23286 ; n23287
g23096 nor n23284 n23287 ; n23288
g23097 nor n23281 n23288 ; n23289
g23098 nor n23279 n23289 ; n23290
g23099 and n22554 n22556_not ; n23291
g23100 and n22547_not n23291 ; n23292
g23101 and asqrt[3] n23292 ; n23293
g23102 nor n22547 n22556 ; n23294
g23103 and asqrt[3] n23294 ; n23295
g23104 nor n22554 n23295 ; n23296
g23105 nor n23293 n23296 ; n23297
g23106 nor n22558 n22565 ; n23298
g23107 and asqrt[3] n23298 ; n23299
g23108 nor n22573 n23299 ; n23300
g23109 and n23297_not n23300 ; n23301
g23110 and n23290_not n23301 ; n23302
g23111 nor asqrt[63] n23302 ; n23303
g23112 and n23279_not n23297 ; n23304
g23113 and n23289_not n23304 ; n23305
g23114 and n22565_not asqrt[3] ; n23306
g23115 and n22558 n23306_not ; n23307
g23116 and asqrt[63] n23298_not ; n23308
g23117 and n23307_not n23308 ; n23309
g23118 nor n23305 n23309 ; n23310
g23119 nand n23303_not n23310 ; asqrt[2]
g23120 and n23255_not n23262 ; n23312
g23121 and n23264_not n23312 ; n23313
g23122 and asqrt[2] n23313 ; n23314
g23123 nor n23255 n23264 ; n23315
g23124 and asqrt[2] n23315 ; n23316
g23125 nor n23262 n23316 ; n23317
g23126 nor n23314 n23317 ; n23318
g23127 and a[4] asqrt[2] ; n23319
g23128 nor a[2] a[3] ; n23320
g23129 and a[4]_not n23320 ; n23321
g23130 nor n23319 n23321 ; n23322
g23131 and asqrt[3] n23322_not ; n23323
g23132 nor n22577 n23321 ; n23324
g23133 and n22573_not n23324 ; n23325
g23134 and n22571_not n23325 ; n23326
g23135 and n23319_not n23326 ; n23327
g23136 and a[4]_not asqrt[2] ; n23328
g23137 and a[5] n23328_not ; n23329
g23138 and n22581 asqrt[2] ; n23330
g23139 nor n23329 n23330 ; n23331
g23140 and n23327_not n23331 ; n23332
g23141 nor n23323 n23332 ; n23333
g23142 and asqrt[4] n23333_not ; n23334
g23143 nor asqrt[4] n23323 ; n23335
g23144 and n23332_not n23335 ; n23336
g23145 and asqrt[3] n23309_not ; n23337
g23146 and n23305_not n23337 ; n23338
g23147 and n23303_not n23338 ; n23339
g23148 nor n23330 n23339 ; n23340
g23149 and a[6] n23340_not ; n23341
g23150 nor a[6] n23339 ; n23342
g23151 and n23330_not n23342 ; n23343
g23152 nor n23341 n23343 ; n23344
g23153 nor n23336 n23344 ; n23345
g23154 nor n23334 n23345 ; n23346
g23155 and asqrt[5] n23346_not ; n23347
g23156 nor n22584 n22588 ; n23348
g23157 and n22592_not n23348 ; n23349
g23158 and asqrt[2] n23349 ; n23350
g23159 and asqrt[2] n23348 ; n23351
g23160 and n22592 n23351_not ; n23352
g23161 nor n23350 n23352 ; n23353
g23162 nor asqrt[5] n23334 ; n23354
g23163 and n23345_not n23354 ; n23355
g23164 nor n23353 n23355 ; n23356
g23165 nor n23347 n23356 ; n23357
g23166 and asqrt[6] n23357_not ; n23358
g23167 and n22597_not n22605 ; n23359
g23168 and n22595_not n23359 ; n23360
g23169 and asqrt[2] n23360 ; n23361
g23170 nor n22595 n22597 ; n23362
g23171 and asqrt[2] n23362 ; n23363
g23172 nor n22605 n23363 ; n23364
g23173 nor n23361 n23364 ; n23365
g23174 nor asqrt[6] n23347 ; n23366
g23175 and n23356_not n23366 ; n23367
g23176 nor n23365 n23367 ; n23368
g23177 nor n23358 n23368 ; n23369
g23178 and asqrt[7] n23369_not ; n23370
g23179 and n22608_not n22614 ; n23371
g23180 and n22616_not n23371 ; n23372
g23181 and asqrt[2] n23372 ; n23373
g23182 nor n22608 n22616 ; n23374
g23183 and asqrt[2] n23374 ; n23375
g23184 nor n22614 n23375 ; n23376
g23185 nor n23373 n23376 ; n23377
g23186 nor asqrt[7] n23358 ; n23378
g23187 and n23368_not n23378 ; n23379
g23188 nor n23377 n23379 ; n23380
g23189 nor n23370 n23380 ; n23381
g23190 and asqrt[8] n23381_not ; n23382
g23191 and n22626 n22628_not ; n23383
g23192 and n22619_not n23383 ; n23384
g23193 and asqrt[2] n23384 ; n23385
g23194 nor n22619 n22628 ; n23386
g23195 and asqrt[2] n23386 ; n23387
g23196 nor n22626 n23387 ; n23388
g23197 nor n23385 n23388 ; n23389
g23198 nor asqrt[8] n23370 ; n23390
g23199 and n23380_not n23390 ; n23391
g23200 nor n23389 n23391 ; n23392
g23201 nor n23382 n23392 ; n23393
g23202 and asqrt[9] n23393_not ; n23394
g23203 and n22631_not n22638 ; n23395
g23204 and n22640_not n23395 ; n23396
g23205 and asqrt[2] n23396 ; n23397
g23206 nor n22631 n22640 ; n23398
g23207 and asqrt[2] n23398 ; n23399
g23208 nor n22638 n23399 ; n23400
g23209 nor n23397 n23400 ; n23401
g23210 nor asqrt[9] n23382 ; n23402
g23211 and n23392_not n23402 ; n23403
g23212 nor n23401 n23403 ; n23404
g23213 nor n23394 n23404 ; n23405
g23214 and asqrt[10] n23405_not ; n23406
g23215 and n22650 n22652_not ; n23407
g23216 and n22643_not n23407 ; n23408
g23217 and asqrt[2] n23408 ; n23409
g23218 nor n22643 n22652 ; n23410
g23219 and asqrt[2] n23410 ; n23411
g23220 nor n22650 n23411 ; n23412
g23221 nor n23409 n23412 ; n23413
g23222 nor asqrt[10] n23394 ; n23414
g23223 and n23404_not n23414 ; n23415
g23224 nor n23413 n23415 ; n23416
g23225 nor n23406 n23416 ; n23417
g23226 and asqrt[11] n23417_not ; n23418
g23227 and n22655_not n22662 ; n23419
g23228 and n22664_not n23419 ; n23420
g23229 and asqrt[2] n23420 ; n23421
g23230 nor n22655 n22664 ; n23422
g23231 and asqrt[2] n23422 ; n23423
g23232 nor n22662 n23423 ; n23424
g23233 nor n23421 n23424 ; n23425
g23234 nor asqrt[11] n23406 ; n23426
g23235 and n23416_not n23426 ; n23427
g23236 nor n23425 n23427 ; n23428
g23237 nor n23418 n23428 ; n23429
g23238 and asqrt[12] n23429_not ; n23430
g23239 and n22674 n22676_not ; n23431
g23240 and n22667_not n23431 ; n23432
g23241 and asqrt[2] n23432 ; n23433
g23242 nor n22667 n22676 ; n23434
g23243 and asqrt[2] n23434 ; n23435
g23244 nor n22674 n23435 ; n23436
g23245 nor n23433 n23436 ; n23437
g23246 nor asqrt[12] n23418 ; n23438
g23247 and n23428_not n23438 ; n23439
g23248 nor n23437 n23439 ; n23440
g23249 nor n23430 n23440 ; n23441
g23250 and asqrt[13] n23441_not ; n23442
g23251 and n22679_not n22686 ; n23443
g23252 and n22688_not n23443 ; n23444
g23253 and asqrt[2] n23444 ; n23445
g23254 nor n22679 n22688 ; n23446
g23255 and asqrt[2] n23446 ; n23447
g23256 nor n22686 n23447 ; n23448
g23257 nor n23445 n23448 ; n23449
g23258 nor asqrt[13] n23430 ; n23450
g23259 and n23440_not n23450 ; n23451
g23260 nor n23449 n23451 ; n23452
g23261 nor n23442 n23452 ; n23453
g23262 and asqrt[14] n23453_not ; n23454
g23263 and n22698 n22700_not ; n23455
g23264 and n22691_not n23455 ; n23456
g23265 and asqrt[2] n23456 ; n23457
g23266 nor n22691 n22700 ; n23458
g23267 and asqrt[2] n23458 ; n23459
g23268 nor n22698 n23459 ; n23460
g23269 nor n23457 n23460 ; n23461
g23270 nor asqrt[14] n23442 ; n23462
g23271 and n23452_not n23462 ; n23463
g23272 nor n23461 n23463 ; n23464
g23273 nor n23454 n23464 ; n23465
g23274 and asqrt[15] n23465_not ; n23466
g23275 and n22703_not n22710 ; n23467
g23276 and n22712_not n23467 ; n23468
g23277 and asqrt[2] n23468 ; n23469
g23278 nor n22703 n22712 ; n23470
g23279 and asqrt[2] n23470 ; n23471
g23280 nor n22710 n23471 ; n23472
g23281 nor n23469 n23472 ; n23473
g23282 nor asqrt[15] n23454 ; n23474
g23283 and n23464_not n23474 ; n23475
g23284 nor n23473 n23475 ; n23476
g23285 nor n23466 n23476 ; n23477
g23286 and asqrt[16] n23477_not ; n23478
g23287 and n22722 n22724_not ; n23479
g23288 and n22715_not n23479 ; n23480
g23289 and asqrt[2] n23480 ; n23481
g23290 nor n22715 n22724 ; n23482
g23291 and asqrt[2] n23482 ; n23483
g23292 nor n22722 n23483 ; n23484
g23293 nor n23481 n23484 ; n23485
g23294 nor asqrt[16] n23466 ; n23486
g23295 and n23476_not n23486 ; n23487
g23296 nor n23485 n23487 ; n23488
g23297 nor n23478 n23488 ; n23489
g23298 and asqrt[17] n23489_not ; n23490
g23299 and n22727_not n22734 ; n23491
g23300 and n22736_not n23491 ; n23492
g23301 and asqrt[2] n23492 ; n23493
g23302 nor n22727 n22736 ; n23494
g23303 and asqrt[2] n23494 ; n23495
g23304 nor n22734 n23495 ; n23496
g23305 nor n23493 n23496 ; n23497
g23306 nor asqrt[17] n23478 ; n23498
g23307 and n23488_not n23498 ; n23499
g23308 nor n23497 n23499 ; n23500
g23309 nor n23490 n23500 ; n23501
g23310 and asqrt[18] n23501_not ; n23502
g23311 and n22746 n22748_not ; n23503
g23312 and n22739_not n23503 ; n23504
g23313 and asqrt[2] n23504 ; n23505
g23314 nor n22739 n22748 ; n23506
g23315 and asqrt[2] n23506 ; n23507
g23316 nor n22746 n23507 ; n23508
g23317 nor n23505 n23508 ; n23509
g23318 nor asqrt[18] n23490 ; n23510
g23319 and n23500_not n23510 ; n23511
g23320 nor n23509 n23511 ; n23512
g23321 nor n23502 n23512 ; n23513
g23322 and asqrt[19] n23513_not ; n23514
g23323 and n22751_not n22758 ; n23515
g23324 and n22760_not n23515 ; n23516
g23325 and asqrt[2] n23516 ; n23517
g23326 nor n22751 n22760 ; n23518
g23327 and asqrt[2] n23518 ; n23519
g23328 nor n22758 n23519 ; n23520
g23329 nor n23517 n23520 ; n23521
g23330 nor asqrt[19] n23502 ; n23522
g23331 and n23512_not n23522 ; n23523
g23332 nor n23521 n23523 ; n23524
g23333 nor n23514 n23524 ; n23525
g23334 and asqrt[20] n23525_not ; n23526
g23335 and n22770 n22772_not ; n23527
g23336 and n22763_not n23527 ; n23528
g23337 and asqrt[2] n23528 ; n23529
g23338 nor n22763 n22772 ; n23530
g23339 and asqrt[2] n23530 ; n23531
g23340 nor n22770 n23531 ; n23532
g23341 nor n23529 n23532 ; n23533
g23342 nor asqrt[20] n23514 ; n23534
g23343 and n23524_not n23534 ; n23535
g23344 nor n23533 n23535 ; n23536
g23345 nor n23526 n23536 ; n23537
g23346 and asqrt[21] n23537_not ; n23538
g23347 and n22775_not n22782 ; n23539
g23348 and n22784_not n23539 ; n23540
g23349 and asqrt[2] n23540 ; n23541
g23350 nor n22775 n22784 ; n23542
g23351 and asqrt[2] n23542 ; n23543
g23352 nor n22782 n23543 ; n23544
g23353 nor n23541 n23544 ; n23545
g23354 nor asqrt[21] n23526 ; n23546
g23355 and n23536_not n23546 ; n23547
g23356 nor n23545 n23547 ; n23548
g23357 nor n23538 n23548 ; n23549
g23358 and asqrt[22] n23549_not ; n23550
g23359 and n22794 n22796_not ; n23551
g23360 and n22787_not n23551 ; n23552
g23361 and asqrt[2] n23552 ; n23553
g23362 nor n22787 n22796 ; n23554
g23363 and asqrt[2] n23554 ; n23555
g23364 nor n22794 n23555 ; n23556
g23365 nor n23553 n23556 ; n23557
g23366 nor asqrt[22] n23538 ; n23558
g23367 and n23548_not n23558 ; n23559
g23368 nor n23557 n23559 ; n23560
g23369 nor n23550 n23560 ; n23561
g23370 and asqrt[23] n23561_not ; n23562
g23371 and n22799_not n22806 ; n23563
g23372 and n22808_not n23563 ; n23564
g23373 and asqrt[2] n23564 ; n23565
g23374 nor n22799 n22808 ; n23566
g23375 and asqrt[2] n23566 ; n23567
g23376 nor n22806 n23567 ; n23568
g23377 nor n23565 n23568 ; n23569
g23378 nor asqrt[23] n23550 ; n23570
g23379 and n23560_not n23570 ; n23571
g23380 nor n23569 n23571 ; n23572
g23381 nor n23562 n23572 ; n23573
g23382 and asqrt[24] n23573_not ; n23574
g23383 and n22818 n22820_not ; n23575
g23384 and n22811_not n23575 ; n23576
g23385 and asqrt[2] n23576 ; n23577
g23386 nor n22811 n22820 ; n23578
g23387 and asqrt[2] n23578 ; n23579
g23388 nor n22818 n23579 ; n23580
g23389 nor n23577 n23580 ; n23581
g23390 nor asqrt[24] n23562 ; n23582
g23391 and n23572_not n23582 ; n23583
g23392 nor n23581 n23583 ; n23584
g23393 nor n23574 n23584 ; n23585
g23394 and asqrt[25] n23585_not ; n23586
g23395 and n22823_not n22830 ; n23587
g23396 and n22832_not n23587 ; n23588
g23397 and asqrt[2] n23588 ; n23589
g23398 nor n22823 n22832 ; n23590
g23399 and asqrt[2] n23590 ; n23591
g23400 nor n22830 n23591 ; n23592
g23401 nor n23589 n23592 ; n23593
g23402 nor asqrt[25] n23574 ; n23594
g23403 and n23584_not n23594 ; n23595
g23404 nor n23593 n23595 ; n23596
g23405 nor n23586 n23596 ; n23597
g23406 and asqrt[26] n23597_not ; n23598
g23407 and n22842 n22844_not ; n23599
g23408 and n22835_not n23599 ; n23600
g23409 and asqrt[2] n23600 ; n23601
g23410 nor n22835 n22844 ; n23602
g23411 and asqrt[2] n23602 ; n23603
g23412 nor n22842 n23603 ; n23604
g23413 nor n23601 n23604 ; n23605
g23414 nor asqrt[26] n23586 ; n23606
g23415 and n23596_not n23606 ; n23607
g23416 nor n23605 n23607 ; n23608
g23417 nor n23598 n23608 ; n23609
g23418 and asqrt[27] n23609_not ; n23610
g23419 and n22847_not n22854 ; n23611
g23420 and n22856_not n23611 ; n23612
g23421 and asqrt[2] n23612 ; n23613
g23422 nor n22847 n22856 ; n23614
g23423 and asqrt[2] n23614 ; n23615
g23424 nor n22854 n23615 ; n23616
g23425 nor n23613 n23616 ; n23617
g23426 nor asqrt[27] n23598 ; n23618
g23427 and n23608_not n23618 ; n23619
g23428 nor n23617 n23619 ; n23620
g23429 nor n23610 n23620 ; n23621
g23430 and asqrt[28] n23621_not ; n23622
g23431 and n22866 n22868_not ; n23623
g23432 and n22859_not n23623 ; n23624
g23433 and asqrt[2] n23624 ; n23625
g23434 nor n22859 n22868 ; n23626
g23435 and asqrt[2] n23626 ; n23627
g23436 nor n22866 n23627 ; n23628
g23437 nor n23625 n23628 ; n23629
g23438 nor asqrt[28] n23610 ; n23630
g23439 and n23620_not n23630 ; n23631
g23440 nor n23629 n23631 ; n23632
g23441 nor n23622 n23632 ; n23633
g23442 and asqrt[29] n23633_not ; n23634
g23443 and n22871_not n22878 ; n23635
g23444 and n22880_not n23635 ; n23636
g23445 and asqrt[2] n23636 ; n23637
g23446 nor n22871 n22880 ; n23638
g23447 and asqrt[2] n23638 ; n23639
g23448 nor n22878 n23639 ; n23640
g23449 nor n23637 n23640 ; n23641
g23450 nor asqrt[29] n23622 ; n23642
g23451 and n23632_not n23642 ; n23643
g23452 nor n23641 n23643 ; n23644
g23453 nor n23634 n23644 ; n23645
g23454 and asqrt[30] n23645_not ; n23646
g23455 and n22890 n22892_not ; n23647
g23456 and n22883_not n23647 ; n23648
g23457 and asqrt[2] n23648 ; n23649
g23458 nor n22883 n22892 ; n23650
g23459 and asqrt[2] n23650 ; n23651
g23460 nor n22890 n23651 ; n23652
g23461 nor n23649 n23652 ; n23653
g23462 nor asqrt[30] n23634 ; n23654
g23463 and n23644_not n23654 ; n23655
g23464 nor n23653 n23655 ; n23656
g23465 nor n23646 n23656 ; n23657
g23466 and asqrt[31] n23657_not ; n23658
g23467 and n22895_not n22902 ; n23659
g23468 and n22904_not n23659 ; n23660
g23469 and asqrt[2] n23660 ; n23661
g23470 nor n22895 n22904 ; n23662
g23471 and asqrt[2] n23662 ; n23663
g23472 nor n22902 n23663 ; n23664
g23473 nor n23661 n23664 ; n23665
g23474 nor asqrt[31] n23646 ; n23666
g23475 and n23656_not n23666 ; n23667
g23476 nor n23665 n23667 ; n23668
g23477 nor n23658 n23668 ; n23669
g23478 and asqrt[32] n23669_not ; n23670
g23479 and n22914 n22916_not ; n23671
g23480 and n22907_not n23671 ; n23672
g23481 and asqrt[2] n23672 ; n23673
g23482 nor n22907 n22916 ; n23674
g23483 and asqrt[2] n23674 ; n23675
g23484 nor n22914 n23675 ; n23676
g23485 nor n23673 n23676 ; n23677
g23486 nor asqrt[32] n23658 ; n23678
g23487 and n23668_not n23678 ; n23679
g23488 nor n23677 n23679 ; n23680
g23489 nor n23670 n23680 ; n23681
g23490 and asqrt[33] n23681_not ; n23682
g23491 and n22919_not n22926 ; n23683
g23492 and n22928_not n23683 ; n23684
g23493 and asqrt[2] n23684 ; n23685
g23494 nor n22919 n22928 ; n23686
g23495 and asqrt[2] n23686 ; n23687
g23496 nor n22926 n23687 ; n23688
g23497 nor n23685 n23688 ; n23689
g23498 nor asqrt[33] n23670 ; n23690
g23499 and n23680_not n23690 ; n23691
g23500 nor n23689 n23691 ; n23692
g23501 nor n23682 n23692 ; n23693
g23502 and asqrt[34] n23693_not ; n23694
g23503 and n22938 n22940_not ; n23695
g23504 and n22931_not n23695 ; n23696
g23505 and asqrt[2] n23696 ; n23697
g23506 nor n22931 n22940 ; n23698
g23507 and asqrt[2] n23698 ; n23699
g23508 nor n22938 n23699 ; n23700
g23509 nor n23697 n23700 ; n23701
g23510 nor asqrt[34] n23682 ; n23702
g23511 and n23692_not n23702 ; n23703
g23512 nor n23701 n23703 ; n23704
g23513 nor n23694 n23704 ; n23705
g23514 and asqrt[35] n23705_not ; n23706
g23515 and n22943_not n22950 ; n23707
g23516 and n22952_not n23707 ; n23708
g23517 and asqrt[2] n23708 ; n23709
g23518 nor n22943 n22952 ; n23710
g23519 and asqrt[2] n23710 ; n23711
g23520 nor n22950 n23711 ; n23712
g23521 nor n23709 n23712 ; n23713
g23522 nor asqrt[35] n23694 ; n23714
g23523 and n23704_not n23714 ; n23715
g23524 nor n23713 n23715 ; n23716
g23525 nor n23706 n23716 ; n23717
g23526 and asqrt[36] n23717_not ; n23718
g23527 and n22962 n22964_not ; n23719
g23528 and n22955_not n23719 ; n23720
g23529 and asqrt[2] n23720 ; n23721
g23530 nor n22955 n22964 ; n23722
g23531 and asqrt[2] n23722 ; n23723
g23532 nor n22962 n23723 ; n23724
g23533 nor n23721 n23724 ; n23725
g23534 nor asqrt[36] n23706 ; n23726
g23535 and n23716_not n23726 ; n23727
g23536 nor n23725 n23727 ; n23728
g23537 nor n23718 n23728 ; n23729
g23538 and asqrt[37] n23729_not ; n23730
g23539 and n22967_not n22974 ; n23731
g23540 and n22976_not n23731 ; n23732
g23541 and asqrt[2] n23732 ; n23733
g23542 nor n22967 n22976 ; n23734
g23543 and asqrt[2] n23734 ; n23735
g23544 nor n22974 n23735 ; n23736
g23545 nor n23733 n23736 ; n23737
g23546 nor asqrt[37] n23718 ; n23738
g23547 and n23728_not n23738 ; n23739
g23548 nor n23737 n23739 ; n23740
g23549 nor n23730 n23740 ; n23741
g23550 and asqrt[38] n23741_not ; n23742
g23551 and n22986 n22988_not ; n23743
g23552 and n22979_not n23743 ; n23744
g23553 and asqrt[2] n23744 ; n23745
g23554 nor n22979 n22988 ; n23746
g23555 and asqrt[2] n23746 ; n23747
g23556 nor n22986 n23747 ; n23748
g23557 nor n23745 n23748 ; n23749
g23558 nor asqrt[38] n23730 ; n23750
g23559 and n23740_not n23750 ; n23751
g23560 nor n23749 n23751 ; n23752
g23561 nor n23742 n23752 ; n23753
g23562 and asqrt[39] n23753_not ; n23754
g23563 and n22991_not n22998 ; n23755
g23564 and n23000_not n23755 ; n23756
g23565 and asqrt[2] n23756 ; n23757
g23566 nor n22991 n23000 ; n23758
g23567 and asqrt[2] n23758 ; n23759
g23568 nor n22998 n23759 ; n23760
g23569 nor n23757 n23760 ; n23761
g23570 nor asqrt[39] n23742 ; n23762
g23571 and n23752_not n23762 ; n23763
g23572 nor n23761 n23763 ; n23764
g23573 nor n23754 n23764 ; n23765
g23574 and asqrt[40] n23765_not ; n23766
g23575 and n23010 n23012_not ; n23767
g23576 and n23003_not n23767 ; n23768
g23577 and asqrt[2] n23768 ; n23769
g23578 nor n23003 n23012 ; n23770
g23579 and asqrt[2] n23770 ; n23771
g23580 nor n23010 n23771 ; n23772
g23581 nor n23769 n23772 ; n23773
g23582 nor asqrt[40] n23754 ; n23774
g23583 and n23764_not n23774 ; n23775
g23584 nor n23773 n23775 ; n23776
g23585 nor n23766 n23776 ; n23777
g23586 and asqrt[41] n23777_not ; n23778
g23587 and n23015_not n23022 ; n23779
g23588 and n23024_not n23779 ; n23780
g23589 and asqrt[2] n23780 ; n23781
g23590 nor n23015 n23024 ; n23782
g23591 and asqrt[2] n23782 ; n23783
g23592 nor n23022 n23783 ; n23784
g23593 nor n23781 n23784 ; n23785
g23594 nor asqrt[41] n23766 ; n23786
g23595 and n23776_not n23786 ; n23787
g23596 nor n23785 n23787 ; n23788
g23597 nor n23778 n23788 ; n23789
g23598 and asqrt[42] n23789_not ; n23790
g23599 and n23034 n23036_not ; n23791
g23600 and n23027_not n23791 ; n23792
g23601 and asqrt[2] n23792 ; n23793
g23602 nor n23027 n23036 ; n23794
g23603 and asqrt[2] n23794 ; n23795
g23604 nor n23034 n23795 ; n23796
g23605 nor n23793 n23796 ; n23797
g23606 nor asqrt[42] n23778 ; n23798
g23607 and n23788_not n23798 ; n23799
g23608 nor n23797 n23799 ; n23800
g23609 nor n23790 n23800 ; n23801
g23610 and asqrt[43] n23801_not ; n23802
g23611 and n23039_not n23046 ; n23803
g23612 and n23048_not n23803 ; n23804
g23613 and asqrt[2] n23804 ; n23805
g23614 nor n23039 n23048 ; n23806
g23615 and asqrt[2] n23806 ; n23807
g23616 nor n23046 n23807 ; n23808
g23617 nor n23805 n23808 ; n23809
g23618 nor asqrt[43] n23790 ; n23810
g23619 and n23800_not n23810 ; n23811
g23620 nor n23809 n23811 ; n23812
g23621 nor n23802 n23812 ; n23813
g23622 and asqrt[44] n23813_not ; n23814
g23623 and n23058 n23060_not ; n23815
g23624 and n23051_not n23815 ; n23816
g23625 and asqrt[2] n23816 ; n23817
g23626 nor n23051 n23060 ; n23818
g23627 and asqrt[2] n23818 ; n23819
g23628 nor n23058 n23819 ; n23820
g23629 nor n23817 n23820 ; n23821
g23630 nor asqrt[44] n23802 ; n23822
g23631 and n23812_not n23822 ; n23823
g23632 nor n23821 n23823 ; n23824
g23633 nor n23814 n23824 ; n23825
g23634 and asqrt[45] n23825_not ; n23826
g23635 and n23063_not n23070 ; n23827
g23636 and n23072_not n23827 ; n23828
g23637 and asqrt[2] n23828 ; n23829
g23638 nor n23063 n23072 ; n23830
g23639 and asqrt[2] n23830 ; n23831
g23640 nor n23070 n23831 ; n23832
g23641 nor n23829 n23832 ; n23833
g23642 nor asqrt[45] n23814 ; n23834
g23643 and n23824_not n23834 ; n23835
g23644 nor n23833 n23835 ; n23836
g23645 nor n23826 n23836 ; n23837
g23646 and asqrt[46] n23837_not ; n23838
g23647 and n23082 n23084_not ; n23839
g23648 and n23075_not n23839 ; n23840
g23649 and asqrt[2] n23840 ; n23841
g23650 nor n23075 n23084 ; n23842
g23651 and asqrt[2] n23842 ; n23843
g23652 nor n23082 n23843 ; n23844
g23653 nor n23841 n23844 ; n23845
g23654 nor asqrt[46] n23826 ; n23846
g23655 and n23836_not n23846 ; n23847
g23656 nor n23845 n23847 ; n23848
g23657 nor n23838 n23848 ; n23849
g23658 and asqrt[47] n23849_not ; n23850
g23659 and n23087_not n23094 ; n23851
g23660 and n23096_not n23851 ; n23852
g23661 and asqrt[2] n23852 ; n23853
g23662 nor n23087 n23096 ; n23854
g23663 and asqrt[2] n23854 ; n23855
g23664 nor n23094 n23855 ; n23856
g23665 nor n23853 n23856 ; n23857
g23666 nor asqrt[47] n23838 ; n23858
g23667 and n23848_not n23858 ; n23859
g23668 nor n23857 n23859 ; n23860
g23669 nor n23850 n23860 ; n23861
g23670 and asqrt[48] n23861_not ; n23862
g23671 and n23106 n23108_not ; n23863
g23672 and n23099_not n23863 ; n23864
g23673 and asqrt[2] n23864 ; n23865
g23674 nor n23099 n23108 ; n23866
g23675 and asqrt[2] n23866 ; n23867
g23676 nor n23106 n23867 ; n23868
g23677 nor n23865 n23868 ; n23869
g23678 nor asqrt[48] n23850 ; n23870
g23679 and n23860_not n23870 ; n23871
g23680 nor n23869 n23871 ; n23872
g23681 nor n23862 n23872 ; n23873
g23682 and asqrt[49] n23873_not ; n23874
g23683 and n23111_not n23118 ; n23875
g23684 and n23120_not n23875 ; n23876
g23685 and asqrt[2] n23876 ; n23877
g23686 nor n23111 n23120 ; n23878
g23687 and asqrt[2] n23878 ; n23879
g23688 nor n23118 n23879 ; n23880
g23689 nor n23877 n23880 ; n23881
g23690 nor asqrt[49] n23862 ; n23882
g23691 and n23872_not n23882 ; n23883
g23692 nor n23881 n23883 ; n23884
g23693 nor n23874 n23884 ; n23885
g23694 and asqrt[50] n23885_not ; n23886
g23695 and n23130 n23132_not ; n23887
g23696 and n23123_not n23887 ; n23888
g23697 and asqrt[2] n23888 ; n23889
g23698 nor n23123 n23132 ; n23890
g23699 and asqrt[2] n23890 ; n23891
g23700 nor n23130 n23891 ; n23892
g23701 nor n23889 n23892 ; n23893
g23702 nor asqrt[50] n23874 ; n23894
g23703 and n23884_not n23894 ; n23895
g23704 nor n23893 n23895 ; n23896
g23705 nor n23886 n23896 ; n23897
g23706 and asqrt[51] n23897_not ; n23898
g23707 and n23135_not n23142 ; n23899
g23708 and n23144_not n23899 ; n23900
g23709 and asqrt[2] n23900 ; n23901
g23710 nor n23135 n23144 ; n23902
g23711 and asqrt[2] n23902 ; n23903
g23712 nor n23142 n23903 ; n23904
g23713 nor n23901 n23904 ; n23905
g23714 nor asqrt[51] n23886 ; n23906
g23715 and n23896_not n23906 ; n23907
g23716 nor n23905 n23907 ; n23908
g23717 nor n23898 n23908 ; n23909
g23718 and asqrt[52] n23909_not ; n23910
g23719 and n23154 n23156_not ; n23911
g23720 and n23147_not n23911 ; n23912
g23721 and asqrt[2] n23912 ; n23913
g23722 nor n23147 n23156 ; n23914
g23723 and asqrt[2] n23914 ; n23915
g23724 nor n23154 n23915 ; n23916
g23725 nor n23913 n23916 ; n23917
g23726 nor asqrt[52] n23898 ; n23918
g23727 and n23908_not n23918 ; n23919
g23728 nor n23917 n23919 ; n23920
g23729 nor n23910 n23920 ; n23921
g23730 and asqrt[53] n23921_not ; n23922
g23731 and n23159_not n23166 ; n23923
g23732 and n23168_not n23923 ; n23924
g23733 and asqrt[2] n23924 ; n23925
g23734 nor n23159 n23168 ; n23926
g23735 and asqrt[2] n23926 ; n23927
g23736 nor n23166 n23927 ; n23928
g23737 nor n23925 n23928 ; n23929
g23738 nor asqrt[53] n23910 ; n23930
g23739 and n23920_not n23930 ; n23931
g23740 nor n23929 n23931 ; n23932
g23741 nor n23922 n23932 ; n23933
g23742 and asqrt[54] n23933_not ; n23934
g23743 and n23178 n23180_not ; n23935
g23744 and n23171_not n23935 ; n23936
g23745 and asqrt[2] n23936 ; n23937
g23746 nor n23171 n23180 ; n23938
g23747 and asqrt[2] n23938 ; n23939
g23748 nor n23178 n23939 ; n23940
g23749 nor n23937 n23940 ; n23941
g23750 nor asqrt[54] n23922 ; n23942
g23751 and n23932_not n23942 ; n23943
g23752 nor n23941 n23943 ; n23944
g23753 nor n23934 n23944 ; n23945
g23754 and asqrt[55] n23945_not ; n23946
g23755 and n23183_not n23190 ; n23947
g23756 and n23192_not n23947 ; n23948
g23757 and asqrt[2] n23948 ; n23949
g23758 nor n23183 n23192 ; n23950
g23759 and asqrt[2] n23950 ; n23951
g23760 nor n23190 n23951 ; n23952
g23761 nor n23949 n23952 ; n23953
g23762 nor asqrt[55] n23934 ; n23954
g23763 and n23944_not n23954 ; n23955
g23764 nor n23953 n23955 ; n23956
g23765 nor n23946 n23956 ; n23957
g23766 and asqrt[56] n23957_not ; n23958
g23767 and n23202 n23204_not ; n23959
g23768 and n23195_not n23959 ; n23960
g23769 and asqrt[2] n23960 ; n23961
g23770 nor n23195 n23204 ; n23962
g23771 and asqrt[2] n23962 ; n23963
g23772 nor n23202 n23963 ; n23964
g23773 nor n23961 n23964 ; n23965
g23774 nor asqrt[56] n23946 ; n23966
g23775 and n23956_not n23966 ; n23967
g23776 nor n23965 n23967 ; n23968
g23777 nor n23958 n23968 ; n23969
g23778 and asqrt[57] n23969_not ; n23970
g23779 and n23207_not n23214 ; n23971
g23780 and n23216_not n23971 ; n23972
g23781 and asqrt[2] n23972 ; n23973
g23782 nor n23207 n23216 ; n23974
g23783 and asqrt[2] n23974 ; n23975
g23784 nor n23214 n23975 ; n23976
g23785 nor n23973 n23976 ; n23977
g23786 nor asqrt[57] n23958 ; n23978
g23787 and n23968_not n23978 ; n23979
g23788 nor n23977 n23979 ; n23980
g23789 nor n23970 n23980 ; n23981
g23790 and asqrt[58] n23981_not ; n23982
g23791 and n23226 n23228_not ; n23983
g23792 and n23219_not n23983 ; n23984
g23793 and asqrt[2] n23984 ; n23985
g23794 nor n23219 n23228 ; n23986
g23795 and asqrt[2] n23986 ; n23987
g23796 nor n23226 n23987 ; n23988
g23797 nor n23985 n23988 ; n23989
g23798 nor asqrt[58] n23970 ; n23990
g23799 and n23980_not n23990 ; n23991
g23800 nor n23989 n23991 ; n23992
g23801 nor n23982 n23992 ; n23993
g23802 and asqrt[59] n23993_not ; n23994
g23803 and n23231_not n23238 ; n23995
g23804 and n23240_not n23995 ; n23996
g23805 and asqrt[2] n23996 ; n23997
g23806 nor n23231 n23240 ; n23998
g23807 and asqrt[2] n23998 ; n23999
g23808 nor n23238 n23999 ; n24000
g23809 nor n23997 n24000 ; n24001
g23810 nor asqrt[59] n23982 ; n24002
g23811 and n23992_not n24002 ; n24003
g23812 nor n24001 n24003 ; n24004
g23813 nor n23994 n24004 ; n24005
g23814 and asqrt[60] n24005_not ; n24006
g23815 and n23250 n23252_not ; n24007
g23816 and n23243_not n24007 ; n24008
g23817 and asqrt[2] n24008 ; n24009
g23818 nor n23243 n23252 ; n24010
g23819 and asqrt[2] n24010 ; n24011
g23820 nor n23250 n24011 ; n24012
g23821 nor n24009 n24012 ; n24013
g23822 nor asqrt[60] n23994 ; n24014
g23823 and n24004_not n24014 ; n24015
g23824 nor n24013 n24015 ; n24016
g23825 nor n24006 n24016 ; n24017
g23826 and asqrt[61] n24017_not ; n24018
g23827 nor asqrt[61] n24006 ; n24019
g23828 and n24016_not n24019 ; n24020
g23829 nor n23318 n24020 ; n24021
g23830 nor n24018 n24021 ; n24022
g23831 and asqrt[62] n24022_not ; n24023
g23832 and n23274 n23276_not ; n24024
g23833 and n23267_not n24024 ; n24025
g23834 and asqrt[2] n24025 ; n24026
g23835 nor n23267 n23276 ; n24027
g23836 and asqrt[2] n24027 ; n24028
g23837 nor n23274 n24028 ; n24029
g23838 nor n24026 n24029 ; n24030
g23839 nor asqrt[62] n24018 ; n24031
g23840 and n24021_not n24031 ; n24032
g23841 nor n24030 n24032 ; n24033
g23842 nor n24023 n24033 ; n24034
g23843 and n23279_not n23288 ; n24035
g23844 and n23281_not n24035 ; n24036
g23845 and asqrt[2] n24036 ; n24037
g23846 nor n23279 n23281 ; n24038
g23847 and asqrt[2] n24038 ; n24039
g23848 nor n23288 n24039 ; n24040
g23849 nor n24037 n24040 ; n24041
g23850 nor n23290 n23297 ; n24042
g23851 and asqrt[2] n24042 ; n24043
g23852 nor n23305 n24043 ; n24044
g23853 and n24041_not n24044 ; n24045
g23854 and n24034_not n24045 ; n24046
g23855 nor asqrt[63] n24046 ; n24047
g23856 and n24023_not n24041 ; n24048
g23857 and n24033_not n24048 ; n24049
g23858 and n23297_not asqrt[2] ; n24050
g23859 and n23290 n24050_not ; n24051
g23860 and asqrt[63] n24042_not ; n24052
g23861 and n24051_not n24052 ; n24053
g23862 nor n24049 n24053 ; n24054
g23863 nand n24047_not n24054 ; asqrt[1]
g23864 nor n24018 n24020 ; n24056
g23865 and asqrt[1] n24056 ; n24057
g23866 nor n23318 n24057 ; n24058
g23867 and n23318 n24018_not ; n24059
g23868 and n24020_not n24059 ; n24060
g23869 and asqrt[1] n24060 ; n24061
g23870 nor n24058 n24061 ; n24062
g23871 nor n23994 n24003 ; n24063
g23872 and asqrt[1] n24063 ; n24064
g23873 nor n24001 n24064 ; n24065
g23874 and n23994_not n24001 ; n24066
g23875 and n24003_not n24066 ; n24067
g23876 and asqrt[1] n24067 ; n24068
g23877 nor n24065 n24068 ; n24069
g23878 nor n23970 n23979 ; n24070
g23879 and asqrt[1] n24070 ; n24071
g23880 nor n23977 n24071 ; n24072
g23881 and n23970_not n23977 ; n24073
g23882 and n23979_not n24073 ; n24074
g23883 and asqrt[1] n24074 ; n24075
g23884 nor n24072 n24075 ; n24076
g23885 nor n23946 n23955 ; n24077
g23886 and asqrt[1] n24077 ; n24078
g23887 nor n23953 n24078 ; n24079
g23888 and n23946_not n23953 ; n24080
g23889 and n23955_not n24080 ; n24081
g23890 and asqrt[1] n24081 ; n24082
g23891 nor n24079 n24082 ; n24083
g23892 nor n23922 n23931 ; n24084
g23893 and asqrt[1] n24084 ; n24085
g23894 nor n23929 n24085 ; n24086
g23895 and n23922_not n23929 ; n24087
g23896 and n23931_not n24087 ; n24088
g23897 and asqrt[1] n24088 ; n24089
g23898 nor n24086 n24089 ; n24090
g23899 nor n23898 n23907 ; n24091
g23900 and asqrt[1] n24091 ; n24092
g23901 nor n23905 n24092 ; n24093
g23902 and n23898_not n23905 ; n24094
g23903 and n23907_not n24094 ; n24095
g23904 and asqrt[1] n24095 ; n24096
g23905 nor n24093 n24096 ; n24097
g23906 nor n23874 n23883 ; n24098
g23907 and asqrt[1] n24098 ; n24099
g23908 nor n23881 n24099 ; n24100
g23909 and n23874_not n23881 ; n24101
g23910 and n23883_not n24101 ; n24102
g23911 and asqrt[1] n24102 ; n24103
g23912 nor n24100 n24103 ; n24104
g23913 nor n23850 n23859 ; n24105
g23914 and asqrt[1] n24105 ; n24106
g23915 nor n23857 n24106 ; n24107
g23916 and n23850_not n23857 ; n24108
g23917 and n23859_not n24108 ; n24109
g23918 and asqrt[1] n24109 ; n24110
g23919 nor n24107 n24110 ; n24111
g23920 nor n23826 n23835 ; n24112
g23921 and asqrt[1] n24112 ; n24113
g23922 nor n23833 n24113 ; n24114
g23923 and n23826_not n23833 ; n24115
g23924 and n23835_not n24115 ; n24116
g23925 and asqrt[1] n24116 ; n24117
g23926 nor n24114 n24117 ; n24118
g23927 nor n23802 n23811 ; n24119
g23928 and asqrt[1] n24119 ; n24120
g23929 nor n23809 n24120 ; n24121
g23930 and n23802_not n23809 ; n24122
g23931 and n23811_not n24122 ; n24123
g23932 and asqrt[1] n24123 ; n24124
g23933 nor n24121 n24124 ; n24125
g23934 nor n23778 n23787 ; n24126
g23935 and asqrt[1] n24126 ; n24127
g23936 nor n23785 n24127 ; n24128
g23937 and n23778_not n23785 ; n24129
g23938 and n23787_not n24129 ; n24130
g23939 and asqrt[1] n24130 ; n24131
g23940 nor n24128 n24131 ; n24132
g23941 nor n23754 n23763 ; n24133
g23942 and asqrt[1] n24133 ; n24134
g23943 nor n23761 n24134 ; n24135
g23944 and n23754_not n23761 ; n24136
g23945 and n23763_not n24136 ; n24137
g23946 and asqrt[1] n24137 ; n24138
g23947 nor n24135 n24138 ; n24139
g23948 nor n23730 n23739 ; n24140
g23949 and asqrt[1] n24140 ; n24141
g23950 nor n23737 n24141 ; n24142
g23951 and n23730_not n23737 ; n24143
g23952 and n23739_not n24143 ; n24144
g23953 and asqrt[1] n24144 ; n24145
g23954 nor n24142 n24145 ; n24146
g23955 nor n23706 n23715 ; n24147
g23956 and asqrt[1] n24147 ; n24148
g23957 nor n23713 n24148 ; n24149
g23958 and n23706_not n23713 ; n24150
g23959 and n23715_not n24150 ; n24151
g23960 and asqrt[1] n24151 ; n24152
g23961 nor n24149 n24152 ; n24153
g23962 nor n23682 n23691 ; n24154
g23963 and asqrt[1] n24154 ; n24155
g23964 nor n23689 n24155 ; n24156
g23965 and n23682_not n23689 ; n24157
g23966 and n23691_not n24157 ; n24158
g23967 and asqrt[1] n24158 ; n24159
g23968 nor n24156 n24159 ; n24160
g23969 nor n23658 n23667 ; n24161
g23970 and asqrt[1] n24161 ; n24162
g23971 nor n23665 n24162 ; n24163
g23972 and n23658_not n23665 ; n24164
g23973 and n23667_not n24164 ; n24165
g23974 and asqrt[1] n24165 ; n24166
g23975 nor n24163 n24166 ; n24167
g23976 nor n23634 n23643 ; n24168
g23977 and asqrt[1] n24168 ; n24169
g23978 nor n23641 n24169 ; n24170
g23979 and n23634_not n23641 ; n24171
g23980 and n23643_not n24171 ; n24172
g23981 and asqrt[1] n24172 ; n24173
g23982 nor n24170 n24173 ; n24174
g23983 nor n23610 n23619 ; n24175
g23984 and asqrt[1] n24175 ; n24176
g23985 nor n23617 n24176 ; n24177
g23986 and n23610_not n23617 ; n24178
g23987 and n23619_not n24178 ; n24179
g23988 and asqrt[1] n24179 ; n24180
g23989 nor n24177 n24180 ; n24181
g23990 nor n23586 n23595 ; n24182
g23991 and asqrt[1] n24182 ; n24183
g23992 nor n23593 n24183 ; n24184
g23993 and n23586_not n23593 ; n24185
g23994 and n23595_not n24185 ; n24186
g23995 and asqrt[1] n24186 ; n24187
g23996 nor n24184 n24187 ; n24188
g23997 nor n23562 n23571 ; n24189
g23998 and asqrt[1] n24189 ; n24190
g23999 nor n23569 n24190 ; n24191
g24000 and n23562_not n23569 ; n24192
g24001 and n23571_not n24192 ; n24193
g24002 and asqrt[1] n24193 ; n24194
g24003 nor n24191 n24194 ; n24195
g24004 nor n23538 n23547 ; n24196
g24005 and asqrt[1] n24196 ; n24197
g24006 nor n23545 n24197 ; n24198
g24007 and n23538_not n23545 ; n24199
g24008 and n23547_not n24199 ; n24200
g24009 and asqrt[1] n24200 ; n24201
g24010 nor n24198 n24201 ; n24202
g24011 nor n23514 n23523 ; n24203
g24012 and asqrt[1] n24203 ; n24204
g24013 nor n23521 n24204 ; n24205
g24014 and n23514_not n23521 ; n24206
g24015 and n23523_not n24206 ; n24207
g24016 and asqrt[1] n24207 ; n24208
g24017 nor n24205 n24208 ; n24209
g24018 nor n23490 n23499 ; n24210
g24019 and asqrt[1] n24210 ; n24211
g24020 nor n23497 n24211 ; n24212
g24021 and n23490_not n23497 ; n24213
g24022 and n23499_not n24213 ; n24214
g24023 and asqrt[1] n24214 ; n24215
g24024 nor n24212 n24215 ; n24216
g24025 nor n23466 n23475 ; n24217
g24026 and asqrt[1] n24217 ; n24218
g24027 nor n23473 n24218 ; n24219
g24028 and n23466_not n23473 ; n24220
g24029 and n23475_not n24220 ; n24221
g24030 and asqrt[1] n24221 ; n24222
g24031 nor n24219 n24222 ; n24223
g24032 nor n23442 n23451 ; n24224
g24033 and asqrt[1] n24224 ; n24225
g24034 nor n23449 n24225 ; n24226
g24035 and n23442_not n23449 ; n24227
g24036 and n23451_not n24227 ; n24228
g24037 and asqrt[1] n24228 ; n24229
g24038 nor n24226 n24229 ; n24230
g24039 nor n23418 n23427 ; n24231
g24040 and asqrt[1] n24231 ; n24232
g24041 nor n23425 n24232 ; n24233
g24042 and n23418_not n23425 ; n24234
g24043 and n23427_not n24234 ; n24235
g24044 and asqrt[1] n24235 ; n24236
g24045 nor n24233 n24236 ; n24237
g24046 nor n23394 n23403 ; n24238
g24047 and asqrt[1] n24238 ; n24239
g24048 nor n23401 n24239 ; n24240
g24049 and n23394_not n23401 ; n24241
g24050 and n23403_not n24241 ; n24242
g24051 and asqrt[1] n24242 ; n24243
g24052 nor n24240 n24243 ; n24244
g24053 nor n23370 n23379 ; n24245
g24054 and asqrt[1] n24245 ; n24246
g24055 nor n23377 n24246 ; n24247
g24056 and n23370_not n23377 ; n24248
g24057 and n23379_not n24248 ; n24249
g24058 and asqrt[1] n24249 ; n24250
g24059 nor n24247 n24250 ; n24251
g24060 and n23347_not n23353 ; n24252
g24061 and n23355_not n24252 ; n24253
g24062 and asqrt[1] n24253 ; n24254
g24063 nor n23347 n23355 ; n24255
g24064 and asqrt[1] n24255 ; n24256
g24065 nor n23353 n24256 ; n24257
g24066 nor n24254 n24257 ; n24258
g24067 nor n23323 n23327 ; n24259
g24068 and n23331_not n24259 ; n24260
g24069 and asqrt[1] n24260 ; n24261
g24070 and asqrt[1] n24259 ; n24262
g24071 and n23331 n24262_not ; n24263
g24072 nor n24261 n24263 ; n24264
g24073 and n23320 asqrt[1] ; n24265
g24074 and asqrt[2] n24053_not ; n24266
g24075 and n24049_not n24266 ; n24267
g24076 and n24047_not n24267 ; n24268
g24077 nor n24265 n24268 ; n24269
g24078 and a[4] n24269_not ; n24270
g24079 nor a[4] n24268 ; n24271
g24080 and n24265_not n24271 ; n24272
g24081 nor n24270 n24272 ; n24273
g24082 and a[2]_not asqrt[1] ; n24274
g24083 and a[3] n24274_not ; n24275
g24084 nor a[0] a[1] ; n24276
g24085 nor a[2] n24276 ; n24277
g24086 and a[2] n24053_not ; n24278
g24087 and n24049_not n24278 ; n24279
g24088 and n24047_not n24279 ; n24280
g24089 nor n24277 n24280 ; n24281
g24090 and n24265_not n24281 ; n24282
g24091 and n24275_not n24282 ; n24283
g24092 nor asqrt[2] n24283 ; n24284
g24093 nor n24265 n24275 ; n24285
g24094 nor n24281 n24285 ; n24286
g24095 nor n24284 n24286 ; n24287
g24096 and n24273_not n24287 ; n24288
g24097 nor asqrt[3] n24288 ; n24289
g24098 and n24273 n24287_not ; n24290
g24099 nor n24289 n24290 ; n24291
g24100 and n24264 n24291_not ; n24292
g24101 nor n24264 n24290 ; n24293
g24102 and n24289_not n24293 ; n24294
g24103 nor asqrt[4] n24294 ; n24295
g24104 nor n23334 n23336 ; n24296
g24105 and asqrt[1] n24296 ; n24297
g24106 nor n23344 n24297 ; n24298
g24107 and n23336_not n23344 ; n24299
g24108 and n23334_not n24299 ; n24300
g24109 and asqrt[1] n24300 ; n24301
g24110 nor n24298 n24301 ; n24302
g24111 nor n24295 n24302 ; n24303
g24112 and n24292_not n24303 ; n24304
g24113 nor asqrt[5] n24304 ; n24305
g24114 nor n24292 n24295 ; n24306
g24115 and n24302 n24306_not ; n24307
g24116 nor n24305 n24307 ; n24308
g24117 and n24258 n24308_not ; n24309
g24118 nor n24258 n24307 ; n24310
g24119 and n24305_not n24310 ; n24311
g24120 nor asqrt[6] n24311 ; n24312
g24121 nor n23358 n23367 ; n24313
g24122 and asqrt[1] n24313 ; n24314
g24123 nor n23365 n24314 ; n24315
g24124 and n23365 n23367_not ; n24316
g24125 and n23358_not n24316 ; n24317
g24126 and asqrt[1] n24317 ; n24318
g24127 nor n24315 n24318 ; n24319
g24128 nor n24312 n24319 ; n24320
g24129 and n24309_not n24320 ; n24321
g24130 nor asqrt[7] n24321 ; n24322
g24131 nor n24309 n24312 ; n24323
g24132 and n24319 n24323_not ; n24324
g24133 nor n24322 n24324 ; n24325
g24134 and n24251 n24325_not ; n24326
g24135 nor n24251 n24324 ; n24327
g24136 and n24322_not n24327 ; n24328
g24137 nor asqrt[8] n24328 ; n24329
g24138 nor n23382 n23391 ; n24330
g24139 and asqrt[1] n24330 ; n24331
g24140 nor n23389 n24331 ; n24332
g24141 and n23389 n23391_not ; n24333
g24142 and n23382_not n24333 ; n24334
g24143 and asqrt[1] n24334 ; n24335
g24144 nor n24332 n24335 ; n24336
g24145 nor n24329 n24336 ; n24337
g24146 and n24326_not n24337 ; n24338
g24147 nor asqrt[9] n24338 ; n24339
g24148 nor n24326 n24329 ; n24340
g24149 and n24336 n24340_not ; n24341
g24150 nor n24339 n24341 ; n24342
g24151 and n24244 n24342_not ; n24343
g24152 nor n24244 n24341 ; n24344
g24153 and n24339_not n24344 ; n24345
g24154 nor asqrt[10] n24345 ; n24346
g24155 nor n23406 n23415 ; n24347
g24156 and asqrt[1] n24347 ; n24348
g24157 nor n23413 n24348 ; n24349
g24158 and n23413 n23415_not ; n24350
g24159 and n23406_not n24350 ; n24351
g24160 and asqrt[1] n24351 ; n24352
g24161 nor n24349 n24352 ; n24353
g24162 nor n24346 n24353 ; n24354
g24163 and n24343_not n24354 ; n24355
g24164 nor asqrt[11] n24355 ; n24356
g24165 nor n24343 n24346 ; n24357
g24166 and n24353 n24357_not ; n24358
g24167 nor n24356 n24358 ; n24359
g24168 and n24237 n24359_not ; n24360
g24169 nor n24237 n24358 ; n24361
g24170 and n24356_not n24361 ; n24362
g24171 nor asqrt[12] n24362 ; n24363
g24172 nor n23430 n23439 ; n24364
g24173 and asqrt[1] n24364 ; n24365
g24174 nor n23437 n24365 ; n24366
g24175 and n23437 n23439_not ; n24367
g24176 and n23430_not n24367 ; n24368
g24177 and asqrt[1] n24368 ; n24369
g24178 nor n24366 n24369 ; n24370
g24179 nor n24363 n24370 ; n24371
g24180 and n24360_not n24371 ; n24372
g24181 nor asqrt[13] n24372 ; n24373
g24182 nor n24360 n24363 ; n24374
g24183 and n24370 n24374_not ; n24375
g24184 nor n24373 n24375 ; n24376
g24185 and n24230 n24376_not ; n24377
g24186 nor n24230 n24375 ; n24378
g24187 and n24373_not n24378 ; n24379
g24188 nor asqrt[14] n24379 ; n24380
g24189 nor n23454 n23463 ; n24381
g24190 and asqrt[1] n24381 ; n24382
g24191 nor n23461 n24382 ; n24383
g24192 and n23461 n23463_not ; n24384
g24193 and n23454_not n24384 ; n24385
g24194 and asqrt[1] n24385 ; n24386
g24195 nor n24383 n24386 ; n24387
g24196 nor n24380 n24387 ; n24388
g24197 and n24377_not n24388 ; n24389
g24198 nor asqrt[15] n24389 ; n24390
g24199 nor n24377 n24380 ; n24391
g24200 and n24387 n24391_not ; n24392
g24201 nor n24390 n24392 ; n24393
g24202 and n24223 n24393_not ; n24394
g24203 nor n24223 n24392 ; n24395
g24204 and n24390_not n24395 ; n24396
g24205 nor asqrt[16] n24396 ; n24397
g24206 nor n23478 n23487 ; n24398
g24207 and asqrt[1] n24398 ; n24399
g24208 nor n23485 n24399 ; n24400
g24209 and n23485 n23487_not ; n24401
g24210 and n23478_not n24401 ; n24402
g24211 and asqrt[1] n24402 ; n24403
g24212 nor n24400 n24403 ; n24404
g24213 nor n24397 n24404 ; n24405
g24214 and n24394_not n24405 ; n24406
g24215 nor asqrt[17] n24406 ; n24407
g24216 nor n24394 n24397 ; n24408
g24217 and n24404 n24408_not ; n24409
g24218 nor n24407 n24409 ; n24410
g24219 and n24216 n24410_not ; n24411
g24220 nor n24216 n24409 ; n24412
g24221 and n24407_not n24412 ; n24413
g24222 nor asqrt[18] n24413 ; n24414
g24223 nor n23502 n23511 ; n24415
g24224 and asqrt[1] n24415 ; n24416
g24225 nor n23509 n24416 ; n24417
g24226 and n23509 n23511_not ; n24418
g24227 and n23502_not n24418 ; n24419
g24228 and asqrt[1] n24419 ; n24420
g24229 nor n24417 n24420 ; n24421
g24230 nor n24414 n24421 ; n24422
g24231 and n24411_not n24422 ; n24423
g24232 nor asqrt[19] n24423 ; n24424
g24233 nor n24411 n24414 ; n24425
g24234 and n24421 n24425_not ; n24426
g24235 nor n24424 n24426 ; n24427
g24236 and n24209 n24427_not ; n24428
g24237 nor n24209 n24426 ; n24429
g24238 and n24424_not n24429 ; n24430
g24239 nor asqrt[20] n24430 ; n24431
g24240 nor n23526 n23535 ; n24432
g24241 and asqrt[1] n24432 ; n24433
g24242 nor n23533 n24433 ; n24434
g24243 and n23533 n23535_not ; n24435
g24244 and n23526_not n24435 ; n24436
g24245 and asqrt[1] n24436 ; n24437
g24246 nor n24434 n24437 ; n24438
g24247 nor n24431 n24438 ; n24439
g24248 and n24428_not n24439 ; n24440
g24249 nor asqrt[21] n24440 ; n24441
g24250 nor n24428 n24431 ; n24442
g24251 and n24438 n24442_not ; n24443
g24252 nor n24441 n24443 ; n24444
g24253 and n24202 n24444_not ; n24445
g24254 nor n24202 n24443 ; n24446
g24255 and n24441_not n24446 ; n24447
g24256 nor asqrt[22] n24447 ; n24448
g24257 nor n23550 n23559 ; n24449
g24258 and asqrt[1] n24449 ; n24450
g24259 nor n23557 n24450 ; n24451
g24260 and n23557 n23559_not ; n24452
g24261 and n23550_not n24452 ; n24453
g24262 and asqrt[1] n24453 ; n24454
g24263 nor n24451 n24454 ; n24455
g24264 nor n24448 n24455 ; n24456
g24265 and n24445_not n24456 ; n24457
g24266 nor asqrt[23] n24457 ; n24458
g24267 nor n24445 n24448 ; n24459
g24268 and n24455 n24459_not ; n24460
g24269 nor n24458 n24460 ; n24461
g24270 and n24195 n24461_not ; n24462
g24271 nor n24195 n24460 ; n24463
g24272 and n24458_not n24463 ; n24464
g24273 nor asqrt[24] n24464 ; n24465
g24274 nor n23574 n23583 ; n24466
g24275 and asqrt[1] n24466 ; n24467
g24276 nor n23581 n24467 ; n24468
g24277 and n23581 n23583_not ; n24469
g24278 and n23574_not n24469 ; n24470
g24279 and asqrt[1] n24470 ; n24471
g24280 nor n24468 n24471 ; n24472
g24281 nor n24465 n24472 ; n24473
g24282 and n24462_not n24473 ; n24474
g24283 nor asqrt[25] n24474 ; n24475
g24284 nor n24462 n24465 ; n24476
g24285 and n24472 n24476_not ; n24477
g24286 nor n24475 n24477 ; n24478
g24287 and n24188 n24478_not ; n24479
g24288 nor n24188 n24477 ; n24480
g24289 and n24475_not n24480 ; n24481
g24290 nor asqrt[26] n24481 ; n24482
g24291 nor n23598 n23607 ; n24483
g24292 and asqrt[1] n24483 ; n24484
g24293 nor n23605 n24484 ; n24485
g24294 and n23605 n23607_not ; n24486
g24295 and n23598_not n24486 ; n24487
g24296 and asqrt[1] n24487 ; n24488
g24297 nor n24485 n24488 ; n24489
g24298 nor n24482 n24489 ; n24490
g24299 and n24479_not n24490 ; n24491
g24300 nor asqrt[27] n24491 ; n24492
g24301 nor n24479 n24482 ; n24493
g24302 and n24489 n24493_not ; n24494
g24303 nor n24492 n24494 ; n24495
g24304 and n24181 n24495_not ; n24496
g24305 nor n24181 n24494 ; n24497
g24306 and n24492_not n24497 ; n24498
g24307 nor asqrt[28] n24498 ; n24499
g24308 nor n23622 n23631 ; n24500
g24309 and asqrt[1] n24500 ; n24501
g24310 nor n23629 n24501 ; n24502
g24311 and n23629 n23631_not ; n24503
g24312 and n23622_not n24503 ; n24504
g24313 and asqrt[1] n24504 ; n24505
g24314 nor n24502 n24505 ; n24506
g24315 nor n24499 n24506 ; n24507
g24316 and n24496_not n24507 ; n24508
g24317 nor asqrt[29] n24508 ; n24509
g24318 nor n24496 n24499 ; n24510
g24319 and n24506 n24510_not ; n24511
g24320 nor n24509 n24511 ; n24512
g24321 and n24174 n24512_not ; n24513
g24322 nor n24174 n24511 ; n24514
g24323 and n24509_not n24514 ; n24515
g24324 nor asqrt[30] n24515 ; n24516
g24325 nor n23646 n23655 ; n24517
g24326 and asqrt[1] n24517 ; n24518
g24327 nor n23653 n24518 ; n24519
g24328 and n23653 n23655_not ; n24520
g24329 and n23646_not n24520 ; n24521
g24330 and asqrt[1] n24521 ; n24522
g24331 nor n24519 n24522 ; n24523
g24332 nor n24516 n24523 ; n24524
g24333 and n24513_not n24524 ; n24525
g24334 nor asqrt[31] n24525 ; n24526
g24335 nor n24513 n24516 ; n24527
g24336 and n24523 n24527_not ; n24528
g24337 nor n24526 n24528 ; n24529
g24338 and n24167 n24529_not ; n24530
g24339 nor n24167 n24528 ; n24531
g24340 and n24526_not n24531 ; n24532
g24341 nor asqrt[32] n24532 ; n24533
g24342 nor n23670 n23679 ; n24534
g24343 and asqrt[1] n24534 ; n24535
g24344 nor n23677 n24535 ; n24536
g24345 and n23677 n23679_not ; n24537
g24346 and n23670_not n24537 ; n24538
g24347 and asqrt[1] n24538 ; n24539
g24348 nor n24536 n24539 ; n24540
g24349 nor n24533 n24540 ; n24541
g24350 and n24530_not n24541 ; n24542
g24351 nor asqrt[33] n24542 ; n24543
g24352 nor n24530 n24533 ; n24544
g24353 and n24540 n24544_not ; n24545
g24354 nor n24543 n24545 ; n24546
g24355 and n24160 n24546_not ; n24547
g24356 nor n24160 n24545 ; n24548
g24357 and n24543_not n24548 ; n24549
g24358 nor asqrt[34] n24549 ; n24550
g24359 nor n23694 n23703 ; n24551
g24360 and asqrt[1] n24551 ; n24552
g24361 nor n23701 n24552 ; n24553
g24362 and n23701 n23703_not ; n24554
g24363 and n23694_not n24554 ; n24555
g24364 and asqrt[1] n24555 ; n24556
g24365 nor n24553 n24556 ; n24557
g24366 nor n24550 n24557 ; n24558
g24367 and n24547_not n24558 ; n24559
g24368 nor asqrt[35] n24559 ; n24560
g24369 nor n24547 n24550 ; n24561
g24370 and n24557 n24561_not ; n24562
g24371 nor n24560 n24562 ; n24563
g24372 and n24153 n24563_not ; n24564
g24373 nor n24153 n24562 ; n24565
g24374 and n24560_not n24565 ; n24566
g24375 nor asqrt[36] n24566 ; n24567
g24376 nor n23718 n23727 ; n24568
g24377 and asqrt[1] n24568 ; n24569
g24378 nor n23725 n24569 ; n24570
g24379 and n23725 n23727_not ; n24571
g24380 and n23718_not n24571 ; n24572
g24381 and asqrt[1] n24572 ; n24573
g24382 nor n24570 n24573 ; n24574
g24383 nor n24567 n24574 ; n24575
g24384 and n24564_not n24575 ; n24576
g24385 nor asqrt[37] n24576 ; n24577
g24386 nor n24564 n24567 ; n24578
g24387 and n24574 n24578_not ; n24579
g24388 nor n24577 n24579 ; n24580
g24389 and n24146 n24580_not ; n24581
g24390 nor n24146 n24579 ; n24582
g24391 and n24577_not n24582 ; n24583
g24392 nor asqrt[38] n24583 ; n24584
g24393 nor n23742 n23751 ; n24585
g24394 and asqrt[1] n24585 ; n24586
g24395 nor n23749 n24586 ; n24587
g24396 and n23749 n23751_not ; n24588
g24397 and n23742_not n24588 ; n24589
g24398 and asqrt[1] n24589 ; n24590
g24399 nor n24587 n24590 ; n24591
g24400 nor n24584 n24591 ; n24592
g24401 and n24581_not n24592 ; n24593
g24402 nor asqrt[39] n24593 ; n24594
g24403 nor n24581 n24584 ; n24595
g24404 and n24591 n24595_not ; n24596
g24405 nor n24594 n24596 ; n24597
g24406 and n24139 n24597_not ; n24598
g24407 nor n24139 n24596 ; n24599
g24408 and n24594_not n24599 ; n24600
g24409 nor asqrt[40] n24600 ; n24601
g24410 nor n23766 n23775 ; n24602
g24411 and asqrt[1] n24602 ; n24603
g24412 nor n23773 n24603 ; n24604
g24413 and n23773 n23775_not ; n24605
g24414 and n23766_not n24605 ; n24606
g24415 and asqrt[1] n24606 ; n24607
g24416 nor n24604 n24607 ; n24608
g24417 nor n24601 n24608 ; n24609
g24418 and n24598_not n24609 ; n24610
g24419 nor asqrt[41] n24610 ; n24611
g24420 nor n24598 n24601 ; n24612
g24421 and n24608 n24612_not ; n24613
g24422 nor n24611 n24613 ; n24614
g24423 and n24132 n24614_not ; n24615
g24424 nor n24132 n24613 ; n24616
g24425 and n24611_not n24616 ; n24617
g24426 nor asqrt[42] n24617 ; n24618
g24427 nor n23790 n23799 ; n24619
g24428 and asqrt[1] n24619 ; n24620
g24429 nor n23797 n24620 ; n24621
g24430 and n23797 n23799_not ; n24622
g24431 and n23790_not n24622 ; n24623
g24432 and asqrt[1] n24623 ; n24624
g24433 nor n24621 n24624 ; n24625
g24434 nor n24618 n24625 ; n24626
g24435 and n24615_not n24626 ; n24627
g24436 nor asqrt[43] n24627 ; n24628
g24437 nor n24615 n24618 ; n24629
g24438 and n24625 n24629_not ; n24630
g24439 nor n24628 n24630 ; n24631
g24440 and n24125 n24631_not ; n24632
g24441 nor n24125 n24630 ; n24633
g24442 and n24628_not n24633 ; n24634
g24443 nor asqrt[44] n24634 ; n24635
g24444 nor n23814 n23823 ; n24636
g24445 and asqrt[1] n24636 ; n24637
g24446 nor n23821 n24637 ; n24638
g24447 and n23821 n23823_not ; n24639
g24448 and n23814_not n24639 ; n24640
g24449 and asqrt[1] n24640 ; n24641
g24450 nor n24638 n24641 ; n24642
g24451 nor n24635 n24642 ; n24643
g24452 and n24632_not n24643 ; n24644
g24453 nor asqrt[45] n24644 ; n24645
g24454 nor n24632 n24635 ; n24646
g24455 and n24642 n24646_not ; n24647
g24456 nor n24645 n24647 ; n24648
g24457 and n24118 n24648_not ; n24649
g24458 nor n24118 n24647 ; n24650
g24459 and n24645_not n24650 ; n24651
g24460 nor asqrt[46] n24651 ; n24652
g24461 nor n23838 n23847 ; n24653
g24462 and asqrt[1] n24653 ; n24654
g24463 nor n23845 n24654 ; n24655
g24464 and n23845 n23847_not ; n24656
g24465 and n23838_not n24656 ; n24657
g24466 and asqrt[1] n24657 ; n24658
g24467 nor n24655 n24658 ; n24659
g24468 nor n24652 n24659 ; n24660
g24469 and n24649_not n24660 ; n24661
g24470 nor asqrt[47] n24661 ; n24662
g24471 nor n24649 n24652 ; n24663
g24472 and n24659 n24663_not ; n24664
g24473 nor n24662 n24664 ; n24665
g24474 and n24111 n24665_not ; n24666
g24475 nor n24111 n24664 ; n24667
g24476 and n24662_not n24667 ; n24668
g24477 nor asqrt[48] n24668 ; n24669
g24478 nor n23862 n23871 ; n24670
g24479 and asqrt[1] n24670 ; n24671
g24480 nor n23869 n24671 ; n24672
g24481 and n23869 n23871_not ; n24673
g24482 and n23862_not n24673 ; n24674
g24483 and asqrt[1] n24674 ; n24675
g24484 nor n24672 n24675 ; n24676
g24485 nor n24669 n24676 ; n24677
g24486 and n24666_not n24677 ; n24678
g24487 nor asqrt[49] n24678 ; n24679
g24488 nor n24666 n24669 ; n24680
g24489 and n24676 n24680_not ; n24681
g24490 nor n24679 n24681 ; n24682
g24491 and n24104 n24682_not ; n24683
g24492 nor n24104 n24681 ; n24684
g24493 and n24679_not n24684 ; n24685
g24494 nor asqrt[50] n24685 ; n24686
g24495 nor n23886 n23895 ; n24687
g24496 and asqrt[1] n24687 ; n24688
g24497 nor n23893 n24688 ; n24689
g24498 and n23893 n23895_not ; n24690
g24499 and n23886_not n24690 ; n24691
g24500 and asqrt[1] n24691 ; n24692
g24501 nor n24689 n24692 ; n24693
g24502 nor n24686 n24693 ; n24694
g24503 and n24683_not n24694 ; n24695
g24504 nor asqrt[51] n24695 ; n24696
g24505 nor n24683 n24686 ; n24697
g24506 and n24693 n24697_not ; n24698
g24507 nor n24696 n24698 ; n24699
g24508 and n24097 n24699_not ; n24700
g24509 nor n24097 n24698 ; n24701
g24510 and n24696_not n24701 ; n24702
g24511 nor asqrt[52] n24702 ; n24703
g24512 nor n23910 n23919 ; n24704
g24513 and asqrt[1] n24704 ; n24705
g24514 nor n23917 n24705 ; n24706
g24515 and n23917 n23919_not ; n24707
g24516 and n23910_not n24707 ; n24708
g24517 and asqrt[1] n24708 ; n24709
g24518 nor n24706 n24709 ; n24710
g24519 nor n24703 n24710 ; n24711
g24520 and n24700_not n24711 ; n24712
g24521 nor asqrt[53] n24712 ; n24713
g24522 nor n24700 n24703 ; n24714
g24523 and n24710 n24714_not ; n24715
g24524 nor n24713 n24715 ; n24716
g24525 and n24090 n24716_not ; n24717
g24526 nor n24090 n24715 ; n24718
g24527 and n24713_not n24718 ; n24719
g24528 nor asqrt[54] n24719 ; n24720
g24529 nor n23934 n23943 ; n24721
g24530 and asqrt[1] n24721 ; n24722
g24531 nor n23941 n24722 ; n24723
g24532 and n23941 n23943_not ; n24724
g24533 and n23934_not n24724 ; n24725
g24534 and asqrt[1] n24725 ; n24726
g24535 nor n24723 n24726 ; n24727
g24536 nor n24720 n24727 ; n24728
g24537 and n24717_not n24728 ; n24729
g24538 nor asqrt[55] n24729 ; n24730
g24539 nor n24717 n24720 ; n24731
g24540 and n24727 n24731_not ; n24732
g24541 nor n24730 n24732 ; n24733
g24542 and n24083 n24733_not ; n24734
g24543 nor n24083 n24732 ; n24735
g24544 and n24730_not n24735 ; n24736
g24545 nor asqrt[56] n24736 ; n24737
g24546 nor n23958 n23967 ; n24738
g24547 and asqrt[1] n24738 ; n24739
g24548 nor n23965 n24739 ; n24740
g24549 and n23965 n23967_not ; n24741
g24550 and n23958_not n24741 ; n24742
g24551 and asqrt[1] n24742 ; n24743
g24552 nor n24740 n24743 ; n24744
g24553 nor n24737 n24744 ; n24745
g24554 and n24734_not n24745 ; n24746
g24555 nor asqrt[57] n24746 ; n24747
g24556 nor n24734 n24737 ; n24748
g24557 and n24744 n24748_not ; n24749
g24558 nor n24747 n24749 ; n24750
g24559 and n24076 n24750_not ; n24751
g24560 nor n24076 n24749 ; n24752
g24561 and n24747_not n24752 ; n24753
g24562 nor asqrt[58] n24753 ; n24754
g24563 nor n23982 n23991 ; n24755
g24564 and asqrt[1] n24755 ; n24756
g24565 nor n23989 n24756 ; n24757
g24566 and n23989 n23991_not ; n24758
g24567 and n23982_not n24758 ; n24759
g24568 and asqrt[1] n24759 ; n24760
g24569 nor n24757 n24760 ; n24761
g24570 nor n24754 n24761 ; n24762
g24571 and n24751_not n24762 ; n24763
g24572 nor asqrt[59] n24763 ; n24764
g24573 nor n24751 n24754 ; n24765
g24574 and n24761 n24765_not ; n24766
g24575 nor n24764 n24766 ; n24767
g24576 and n24069 n24767_not ; n24768
g24577 nor n24069 n24766 ; n24769
g24578 and n24764_not n24769 ; n24770
g24579 nor asqrt[60] n24770 ; n24771
g24580 nor n24006 n24015 ; n24772
g24581 and asqrt[1] n24772 ; n24773
g24582 nor n24013 n24773 ; n24774
g24583 and n24013 n24015_not ; n24775
g24584 and n24006_not n24775 ; n24776
g24585 and asqrt[1] n24776 ; n24777
g24586 nor n24774 n24777 ; n24778
g24587 nor n24771 n24778 ; n24779
g24588 and n24768_not n24779 ; n24780
g24589 nor asqrt[61] n24780 ; n24781
g24590 nor n24768 n24771 ; n24782
g24591 and n24778 n24782_not ; n24783
g24592 nor n24781 n24783 ; n24784
g24593 and n24062 n24784_not ; n24785
g24594 nor n24062 n24783 ; n24786
g24595 and n24781_not n24786 ; n24787
g24596 nor asqrt[62] n24787 ; n24788
g24597 nor n24023 n24032 ; n24789
g24598 and asqrt[1] n24789 ; n24790
g24599 nor n24030 n24790 ; n24791
g24600 and n24030 n24032_not ; n24792
g24601 and n24023_not n24792 ; n24793
g24602 and asqrt[1] n24793 ; n24794
g24603 nor n24791 n24794 ; n24795
g24604 nor n24034 n24041 ; n24796
g24605 and asqrt[1] n24796 ; n24797
g24606 nor n24049 n24797 ; n24798
g24607 and n24795_not n24798 ; n24799
g24608 and n24788_not n24799 ; n24800
g24609 and n24785_not n24800 ; n24801
g24610 nor asqrt[63] n24801 ; n24802
g24611 nor n24785 n24788 ; n24803
g24612 and n24795 n24803_not ; n24804
g24613 and n24041_not asqrt[1] ; n24805
g24614 and n24034 n24805_not ; n24806
g24615 and asqrt[63] n24796_not ; n24807
g24616 and n24806_not n24807 ; n24808
g24617 nor n24804 n24808 ; n24809
g24618 nand n24802_not n24809 ; asqrt[0]
g24619 not n300 ; n300_not
g24620 not n210 ; n210_not
g24621 not n202 ; n202_not
g24622 not n211 ; n211_not
g24623 not n203 ; n203_not
g24624 not n401 ; n401_not
g24625 not n510 ; n510_not
g24626 not n600 ; n600_not
g24627 not n321 ; n321_not
g24628 not n213 ; n213_not
g24629 not n312 ; n312_not
g24630 not n250 ; n250_not
g24631 not n223 ; n223_not
g24632 not n520 ; n520_not
g24633 not n322 ; n322_not
g24634 not n601 ; n601_not
g24635 not n412 ; n412_not
g24636 not n430 ; n430_not
g24637 not n511 ; n511_not
g24638 not n350 ; n350_not
g24639 not n341 ; n341_not
g24640 not n242 ; n242_not
g24641 not n800 ; n800_not
g24642 not n332 ; n332_not
g24643 not n521 ; n521_not
g24644 not n206 ; n206_not
g24645 not n530 ; n530_not
g24646 not n602 ; n602_not
g24647 not n224 ; n224_not
g24648 not n233 ; n233_not
g24649 not n305 ; n305_not
g24650 not n323 ; n323_not
g24651 not n324 ; n324_not
g24652 not n243 ; n243_not
g24653 not n810 ; n810_not
g24654 not n720 ; n720_not
g24655 not n234 ; n234_not
g24656 not n801 ; n801_not
g24657 not n216 ; n216_not
g24658 not n225 ; n225_not
g24659 not n207 ; n207_not
g24660 not n522 ; n522_not
g24661 not n603 ; n603_not
g24662 not n612 ; n612_not
g24663 not n261 ; n261_not
g24664 not n730 ; n730_not
g24665 not n271 ; n271_not
g24666 not n325 ; n325_not
g24667 not n406 ; n406_not
g24668 not n550 ; n550_not
g24669 not n541 ; n541_not
g24670 not n811 ; n811_not
g24671 not n613 ; n613_not
g24672 not n208 ; n208_not
g24673 not n244 ; n244_not
g24674 not n911 ; n911_not
g24675 not n731 ; n731_not
g24676 not n902 ; n902_not
g24677 not n407 ; n407_not
g24678 not n470 ; n470_not
g24679 not n443 ; n443_not
g24680 not n821 ; n821_not
g24681 not n227 ; n227_not
g24682 not n812 ; n812_not
g24683 not n461 ; n461_not
g24684 not n254 ; n254_not
g24685 not n641 ; n641_not
g24686 not n632 ; n632_not
g24687 not n209 ; n209_not
g24688 not n416 ; n416_not
g24689 not n245 ; n245_not
g24690 not n281 ; n281_not
g24691 not n614 ; n614_not
g24692 not n650 ; n650_not
g24693 not n471 ; n471_not
g24694 not n642 ; n642_not
g24695 not n615 ; n615_not
g24696 not n633 ; n633_not
g24697 not n417 ; n417_not
g24698 not n219 ; n219_not
g24699 not n327 ; n327_not
g24700 not n363 ; n363_not
g24701 not n237 ; n237_not
g24702 not n732 ; n732_not
g24703 not n750 ; n750_not
g24704 not n624 ; n624_not
g24705 not n408 ; n408_not
g24706 not n741 ; n741_not
g24707 not n390 ; n390_not
g24708 not n318 ; n318_not
g24709 not n309 ; n309_not
g24710 not n282 ; n282_not
g24711 not n705 ; n705_not
g24712 not n822 ; n822_not
g24713 not n381 ; n381_not
g24714 not n912 ; n912_not
g24715 not n436 ; n436_not
g24716 not n346 ; n346_not
g24717 not n229 ; n229_not
g24718 not n823 ; n823_not
g24719 not n580 ; n580_not
g24720 not n706 ; n706_not
g24721 not n670 ; n670_not
g24722 not n391 ; n391_not
g24723 not n922 ; n922_not
g24724 not n445 ; n445_not
g24725 not n337 ; n337_not
g24726 not n535 ; n535_not
g24727 not n553 ; n553_not
g24728 not n247 ; n247_not
g24729 not n643 ; n643_not
g24730 not n634 ; n634_not
g24731 not n625 ; n625_not
g24732 not n319 ; n319_not
g24733 not n508 ; n508_not
g24734 not n940 ; n940_not
g24735 not n742 ; n742_not
g24736 not n805 ; n805_not
g24737 not n751 ; n751_not
g24738 not n472 ; n472_not
g24739 not n454 ; n454_not
g24740 not n913 ; n913_not
g24741 not n481 ; n481_not
g24742 not n418 ; n418_not
g24743 not n760 ; n760_not
g24744 not n356 ; n356_not
g24745 not n446 ; n446_not
g24746 not n563 ; n563_not
g24747 not n824 ; n824_not
g24748 not n338 ; n338_not
g24749 not n392 ; n392_not
g24750 not n419 ; n419_not
g24751 not n365 ; n365_not
g24752 not n374 ; n374_not
g24753 not n860 ; n860_not
g24754 not n590 ; n590_not
g24755 not n437 ; n437_not
g24756 not n266 ; n266_not
g24757 not n257 ; n257_not
g24758 not n473 ; n473_not
g24759 not n743 ; n743_not
g24760 not n509 ; n509_not
g24761 not n428 ; n428_not
g24762 not n707 ; n707_not
g24763 not n914 ; n914_not
g24764 not n554 ; n554_not
g24765 not n950 ; n950_not
g24766 not n626 ; n626_not
g24767 not n951 ; n951_not
g24768 not n645 ; n645_not
g24769 not n870 ; n870_not
g24770 not n672 ; n672_not
g24771 not n762 ; n762_not
g24772 not n591 ; n591_not
g24773 not n834 ; n834_not
g24774 not n708 ; n708_not
g24775 not n780 ; n780_not
g24776 not n717 ; n717_not
g24777 not n663 ; n663_not
g24778 not n771 ; n771_not
g24779 not n654 ; n654_not
g24780 not n537 ; n537_not
g24781 not n933 ; n933_not
g24782 not n528 ; n528_not
g24783 not n294 ; n294_not
g24784 not n339 ; n339_not
g24785 not n429 ; n429_not
g24786 not n915 ; n915_not
g24787 not n357 ; n357_not
g24788 not n555 ; n555_not
g24789 not n492 ; n492_not
g24790 not n258 ; n258_not
g24791 not n564 ; n564_not
g24792 not n393 ; n393_not
g24793 not n267 ; n267_not
g24794 not n447 ; n447_not
g24795 not n474 ; n474_not
g24796 not n276 ; n276_not
g24797 not n438 ; n438_not
g24798 not n573 ; n573_not
g24799 not n546 ; n546_not
g24800 not n529 ; n529_not
g24801 not n781 ; n781_not
g24802 not n691 ; n691_not
g24803 not n538 ; n538_not
g24804 not n682 ; n682_not
g24805 not n286 ; n286_not
g24806 not n394 ; n394_not
g24807 not n259 ; n259_not
g24808 not n718 ; n718_not
g24809 not n367 ; n367_not
g24810 not n349 ; n349_not
g24811 not n835 ; n835_not
g24812 not n664 ; n664_not
g24813 not n565 ; n565_not
g24814 not n961 ; n961_not
g24815 not n871 ; n871_not
g24816 not n952 ; n952_not
g24817 not n826 ; n826_not
g24818 not n268 ; n268_not
g24819 not n908 ; n908_not
g24820 not n962 ; n962_not
g24821 not n296 ; n296_not
g24822 not n287 ; n287_not
g24823 not n269 ; n269_not
g24824 not n836 ; n836_not
g24825 not n845 ; n845_not
g24826 not n890 ; n890_not
g24827 not n476 ; n476_not
g24828 not n809 ; n809_not
g24829 not n584 ; n584_not
g24830 not n197 ; n197_not
g24831 not n557 ; n557_not
g24832 not n449 ; n449_not
g24833 not n539 ; n539_not
g24834 not n917 ; n917_not
g24835 not n683 ; n683_not
g24836 not n566 ; n566_not
g24837 not n719 ; n719_not
g24838 not n458 ; n458_not
g24839 not n467 ; n467_not
g24840 not n288 ; n288_not
g24841 not n666 ; n666_not
g24842 not n639 ; n639_not
g24843 not n396 ; n396_not
g24844 not n486 ; n486_not
g24845 not n468 ; n468_not
g24846 not n684 ; n684_not
g24847 not n927 ; n927_not
g24848 not n729 ; n729_not
g24849 not n756 ; n756_not
g24850 not n846 ; n846_not
g24851 not n657 ; n657_not
g24852 not n774 ; n774_not
g24853 not n369 ; n369_not
g24854 not n909 ; n909_not
g24855 not n387 ; n387_not
g24856 not n963 ; n963_not
g24857 not n378 ; n378_not
g24858 not n783 ; n783_not
g24859 not n496 ; n496_not
g24860 not n298 ; n298_not
g24861 not n937 ; n937_not
g24862 not n964 ; n964_not
g24863 not n847 ; n847_not
g24864 not n487 ; n487_not
g24865 not n784 ; n784_not
g24866 not n928 ; n928_not
g24867 not n667 ; n667_not
g24868 not n568 ; n568_not
g24869 not n694 ; n694_not
g24870 not n973 ; n973_not
g24871 not n388 ; n388_not
g24872 not n929 ; n929_not
g24873 not n974 ; n974_not
g24874 not n758 ; n758_not
g24875 not n884 ; n884_not
g24876 not n938 ; n938_not
g24877 not n695 ; n695_not
g24878 not n497 ; n497_not
g24879 not n677 ; n677_not
g24880 not n668 ; n668_not
g24881 not n785 ; n785_not
g24882 not n767 ; n767_not
g24883 not n794 ; n794_not
g24884 not n857 ; n857_not
g24885 not n578 ; n578_not
g24886 not n686 ; n686_not
g24887 not n488 ; n488_not
g24888 not n848 ; n848_not
g24889 not n749 ; n749_not
g24890 not n579 ; n579_not
g24891 not n939 ; n939_not
g24892 not n669 ; n669_not
g24893 not n588 ; n588_not
g24894 not n498 ; n498_not
g24895 not n759 ; n759_not
g24896 not n786 ; n786_not
g24897 not n975 ; n975_not
g24898 not n696 ; n696_not
g24899 not n858 ; n858_not
g24900 not n976 ; n976_not
g24901 not n886 ; n886_not
g24902 not n877 ; n877_not
g24903 not n949 ; n949_not
g24904 not n787 ; n787_not
g24905 not n895 ; n895_not
g24906 not n499 ; n499_not
g24907 not n589 ; n589_not
g24908 not n859 ; n859_not
g24909 not n878 ; n878_not
g24910 not n869 ; n869_not
g24911 not n986 ; n986_not
g24912 not n887 ; n887_not
g24913 not n987 ; n987_not
g24914 not n879 ; n879_not
g24915 not n888 ; n888_not
g24916 not n978 ; n978_not
g24917 not n789 ; n789_not
g24918 not n799 ; n799_not
g24919 not n997 ; n997_not
g24920 not n988 ; n988_not
g24921 not n998 ; n998_not
g24922 not n899 ; n899_not
g24923 not n999 ; n999_not
g24924 not n1000 ; n1000_not
g24925 not n1010 ; n1010_not
g24926 not n3000 ; n3000_not
g24927 not n1101 ; n1101_not
g24928 not n1200 ; n1200_not
g24929 not n1011 ; n1011_not
g24930 not n1030 ; n1030_not
g24931 not n2020 ; n2020_not
g24932 not n3001 ; n3001_not
g24933 not n2110 ; n2110_not
g24934 not n1201 ; n1201_not
g24935 not n3010 ; n3010_not
g24936 not n1102 ; n1102_not
g24937 not n3100 ; n3100_not
g24938 not n4100 ; n4100_not
g24939 not n1103 ; n1103_not
g24940 not n1220 ; n1220_not
g24941 not n1301 ; n1301_not
g24942 not n2120 ; n2120_not
g24943 not n2111 ; n2111_not
g24944 not n3110 ; n3110_not
g24945 not n5000 ; n5000_not
g24946 not n3011 ; n3011_not
g24947 not n3200 ; n3200_not
g24948 not n2021 ; n2021_not
g24949 not n2030 ; n2030_not
g24950 not n2102 ; n2102_not
g24951 not n1302 ; n1302_not
g24952 not n1140 ; n1140_not
g24953 not n1104 ; n1104_not
g24954 not n1113 ; n1113_not
g24955 not n1221 ; n1221_not
g24956 not n4002 ; n4002_not
g24957 not n1230 ; n1230_not
g24958 not n3012 ; n3012_not
g24959 not n5001 ; n5001_not
g24960 not n5010 ; n5010_not
g24961 not n1203 ; n1203_not
g24962 not n2031 ; n2031_not
g24963 not n2103 ; n2103_not
g24964 not n2112 ; n2112_not
g24965 not n2121 ; n2121_not
g24966 not n4101 ; n4101_not
g24967 not n2220 ; n2220_not
g24968 not n4110 ; n4110_not
g24969 not n3201 ; n3201_not
g24970 not n3210 ; n3210_not
g24971 not n1024 ; n1024_not
g24972 not n4111 ; n4111_not
g24973 not n1420 ; n1420_not
g24974 not n3103 ; n3103_not
g24975 not n4300 ; n4300_not
g24976 not n1510 ; n1510_not
g24977 not n1231 ; n1231_not
g24978 not n3112 ; n3112_not
g24979 not n2230 ; n2230_not
g24980 not n2221 ; n2221_not
g24981 not n5011 ; n5011_not
g24982 not n2302 ; n2302_not
g24983 not n3130 ; n3130_not
g24984 not n1204 ; n1204_not
g24985 not n3400 ; n3400_not
g24986 not n1303 ; n1303_not
g24987 not n6010 ; n6010_not
g24988 not n2104 ; n2104_not
g24989 not n3211 ; n3211_not
g24990 not n1114 ; n1114_not
g24991 not n2032 ; n2032_not
g24992 not n1051 ; n1051_not
g24993 not n3022 ; n3022_not
g24994 not n1150 ; n1150_not
g24995 not n4003 ; n4003_not
g24996 not n3013 ; n3013_not
g24997 not n1042 ; n1042_not
g24998 not n1501 ; n1501_not
g24999 not n2132 ; n2132_not
g25000 not n4004 ; n4004_not
g25001 not n3140 ; n3140_not
g25002 not n1430 ; n1430_not
g25003 not n6200 ; n6200_not
g25004 not n1232 ; n1232_not
g25005 not n1241 ; n1241_not
g25006 not n3410 ; n3410_not
g25007 not n3023 ; n3023_not
g25008 not n3320 ; n3320_not
g25009 not n1340 ; n1340_not
g25010 not n2231 ; n2231_not
g25011 not n3113 ; n3113_not
g25012 not n3401 ; n3401_not
g25013 not n7010 ; n7010_not
g25014 not n1142 ; n1142_not
g25015 not n4220 ; n4220_not
g25016 not n2006 ; n2006_not
g25017 not n2303 ; n2303_not
g25018 not n4310 ; n4310_not
g25019 not n4301 ; n4301_not
g25020 not n2123 ; n2123_not
g25021 not n2033 ; n2033_not
g25022 not n1520 ; n1520_not
g25023 not n1511 ; n1511_not
g25024 not n1502 ; n1502_not
g25025 not n5012 ; n5012_not
g25026 not n2150 ; n2150_not
g25027 not n6020 ; n6020_not
g25028 not n1304 ; n1304_not
g25029 not n1313 ; n1313_not
g25030 not n2042 ; n2042_not
g25031 not n4112 ; n4112_not
g25032 not n2420 ; n2420_not
g25033 not n2141 ; n2141_not
g25034 not n1205 ; n1205_not
g25035 not n1115 ; n1115_not
g25036 not n1214 ; n1214_not
g25037 not n1151 ; n1151_not
g25038 not n1052 ; n1052_not
g25039 not n3212 ; n3212_not
g25040 not n4040 ; n4040_not
g25041 not n5120 ; n5120_not
g25042 not n5022 ; n5022_not
g25043 not n6210 ; n6210_not
g25044 not n6201 ; n6201_not
g25045 not n2007 ; n2007_not
g25046 not n1431 ; n1431_not
g25047 not n1026 ; n1026_not
g25048 not n2232 ; n2232_not
g25049 not n1503 ; n1503_not
g25050 not n4221 ; n4221_not
g25051 not n3123 ; n3123_not
g25052 not n2043 ; n2043_not
g25053 not n1062 ; n1062_not
g25054 not n3213 ; n3213_not
g25055 not n3222 ; n3222_not
g25056 not n2142 ; n2142_not
g25057 not n1035 ; n1035_not
g25058 not n1053 ; n1053_not
g25059 not n2160 ; n2160_not
g25060 not n2610 ; n2610_not
g25061 not n1242 ; n1242_not
g25062 not n4311 ; n4311_not
g25063 not n7020 ; n7020_not
g25064 not n1017 ; n1017_not
g25065 not n3330 ; n3330_not
g25066 not n3321 ; n3321_not
g25067 not n1710 ; n1710_not
g25068 not n4005 ; n4005_not
g25069 not n4014 ; n4014_not
g25070 not n3060 ; n3060_not
g25071 not n5202 ; n5202_not
g25072 not n6003 ; n6003_not
g25073 not n1620 ; n1620_not
g25074 not n3024 ; n3024_not
g25075 not n1152 ; n1152_not
g25076 not n3114 ; n3114_not
g25077 not n1170 ; n1170_not
g25078 not n8001 ; n8001_not
g25079 not n5013 ; n5013_not
g25080 not n8010 ; n8010_not
g25081 not n4050 ; n4050_not
g25082 not n4041 ; n4041_not
g25083 not n1206 ; n1206_not
g25084 not n4230 ; n4230_not
g25085 not n2601 ; n2601_not
g25086 not n3402 ; n3402_not
g25087 not n5121 ; n5121_not
g25088 not n1116 ; n1116_not
g25089 not n5130 ; n5130_not
g25090 not n3411 ; n3411_not
g25091 not n6102 ; n6102_not
g25092 not n3150 ; n3150_not
g25093 not n3141 ; n3141_not
g25094 not n8100 ; n8100_not
g25095 not n2430 ; n2430_not
g25096 not n2421 ; n2421_not
g25097 not n1161 ; n1161_not
g25098 not n4113 ; n4113_not
g25099 not n1125 ; n1125_not
g25100 not n4122 ; n4122_not
g25101 not n2502 ; n2502_not
g25102 not n1080 ; n1080_not
g25103 not n2304 ; n2304_not
g25104 not n6030 ; n6030_not
g25105 not n1314 ; n1314_not
g25106 not n6021 ; n6021_not
g25107 not n1162 ; n1162_not
g25108 not n8101 ; n8101_not
g25109 not n7210 ; n7210_not
g25110 not n5131 ; n5131_not
g25111 not n1009 ; n1009_not
g25112 not n1630 ; n1630_not
g25113 not n2602 ; n2602_not
g25114 not n1441 ; n1441_not
g25115 not n1018 ; n1018_not
g25116 not n5320 ; n5320_not
g25117 not n4240 ; n4240_not
g25118 not n2620 ; n2620_not
g25119 not n9100 ; n9100_not
g25120 not n1180 ; n1180_not
g25121 not n5500 ; n5500_not
g25122 not n1171 ; n1171_not
g25123 not n4123 ; n4123_not
g25124 not n6400 ; n6400_not
g25125 not n2800 ; n2800_not
g25126 not n1522 ; n1522_not
g25127 not n3061 ; n3061_not
g25128 not n2080 ; n2080_not
g25129 not n4051 ; n4051_not
g25130 not n2206 ; n2206_not
g25131 not n4420 ; n4420_not
g25132 not n2431 ; n2431_not
g25133 not n2170 ; n2170_not
g25134 not n6031 ; n6031_not
g25135 not n3070 ; n3070_not
g25136 not n2341 ; n2341_not
g25137 not n2161 ; n2161_not
g25138 not n1054 ; n1054_not
g25139 not n3223 ; n3223_not
g25140 not n1027 ; n1027_not
g25141 not n3331 ; n3331_not
g25142 not n6103 ; n6103_not
g25143 not n8011 ; n8011_not
g25144 not n3034 ; n3034_not
g25145 not n3412 ; n3412_not
g25146 not n2314 ; n2314_not
g25147 not n2008 ; n2008_not
g25148 not n2305 ; n2305_not
g25149 not n3025 ; n3025_not
g25150 not n1126 ; n1126_not
g25151 not n2503 ; n2503_not
g25152 not n2242 ; n2242_not
g25153 not n1090 ; n1090_not
g25154 not n2044 ; n2044_not
g25155 not n2233 ; n2233_not
g25156 not n4015 ; n4015_not
g25157 not n3520 ; n3520_not
g25158 not n1351 ; n1351_not
g25159 not n4231 ; n4231_not
g25160 not n1342 ; n1342_not
g25161 not n7021 ; n7021_not
g25162 not n5203 ; n5203_not
g25163 not n1207 ; n1207_not
g25164 not n1405 ; n1405_not
g25165 not n4312 ; n4312_not
g25166 not n5023 ; n5023_not
g25167 not n1243 ; n1243_not
g25168 not n1225 ; n1225_not
g25169 not n1333 ; n1333_not
g25170 not n1531 ; n1531_not
g25171 not n1540 ; n1540_not
g25172 not n3115 ; n3115_not
g25173 not n1432 ; n1432_not
g25174 not n1315 ; n1315_not
g25175 not n3151 ; n3151_not
g25176 not n6211 ; n6211_not
g25177 not n1820 ; n1820_not
g25178 not n2621 ; n2621_not
g25179 not n6320 ; n6320_not
g25180 not n8030 ; n8030_not
g25181 not n1091 ; n1091_not
g25182 not n1055 ; n1055_not
g25183 not n3332 ; n3332_not
g25184 not n1073 ; n1073_not
g25185 not n3224 ; n3224_not
g25186 not n2801 ; n2801_not
g25187 not n1910 ; n1910_not
g25188 not n7103 ; n7103_not
g25189 not n2117 ; n2117_not
g25190 not n2135 ; n2135_not
g25191 not n7022 ; n7022_not
g25192 not n1280 ; n1280_not
g25193 not n5024 ; n5024_not
g25194 not n2144 ; n2144_not
g25195 not n6014 ; n6014_not
g25196 not n8210 ; n8210_not
g25197 not n1163 ; n1163_not
g25198 not n4502 ; n4502_not
g25199 not n7400 ; n7400_not
g25200 not n6104 ; n6104_not
g25201 not n1541 ; n1541_not
g25202 not n7220 ; n7220_not
g25203 not n2540 ; n2540_not
g25204 not n1334 ; n1334_not
g25205 not n6212 ; n6212_not
g25206 not n1316 ; n1316_not
g25207 not n4421 ; n4421_not
g25208 not n4430 ; n4430_not
g25209 not n1343 ; n1343_not
g25210 not n5600 ; n5600_not
g25211 not n1127 ; n1127_not
g25212 not n2054 ; n2054_not
g25213 not n2090 ; n2090_not
g25214 not n2081 ; n2081_not
g25215 not n2315 ; n2315_not
g25216 not n3602 ; n3602_not
g25217 not n6140 ; n6140_not
g25218 not n1406 ; n1406_not
g25219 not n3152 ; n3152_not
g25220 not n4016 ; n4016_not
g25221 not n3116 ; n3116_not
g25222 not n6401 ; n6401_not
g25223 not n2162 ; n2162_not
g25224 not n4052 ; n4052_not
g25225 not n2432 ; n2432_not
g25226 not n5204 ; n5204_not
g25227 not n6410 ; n6410_not
g25228 not n1370 ; n1370_not
g25229 not n2504 ; n2504_not
g25230 not n5321 ; n5321_not
g25231 not n3134 ; n3134_not
g25232 not n5060 ; n5060_not
g25233 not n7031 ; n7031_not
g25234 not n2171 ; n2171_not
g25235 not n3260 ; n3260_not
g25236 not n2630 ; n2630_not
g25237 not n4160 ; n4160_not
g25238 not n4322 ; n4322_not
g25239 not n2207 ; n2207_not
g25240 not n6032 ; n6032_not
g25241 not n5132 ; n5132_not
g25242 not n1442 ; n1442_not
g25243 not n4313 ; n4313_not
g25244 not n2018 ; n2018_not
g25245 not n2009 ; n2009_not
g25246 not n2243 ; n2243_not
g25247 not n1028 ; n1028_not
g25248 not n1019 ; n1019_not
g25249 not n1253 ; n1253_not
g25250 not n1244 ; n1244_not
g25251 not n2045 ; n2045_not
g25252 not n5510 ; n5510_not
g25253 not n3080 ; n3080_not
g25254 not n4124 ; n4124_not
g25255 not n9101 ; n9101_not
g25256 not n3071 ; n3071_not
g25257 not n3422 ; n3422_not
g25258 not n4610 ; n4610_not
g25259 not n3521 ; n3521_not
g25260 not n5402 ; n5402_not
g25261 not n5330 ; n5330_not
g25262 not n2810 ; n2810_not
g25263 not n3530 ; n3530_not
g25264 not n5501 ; n5501_not
g25265 not n3251 ; n3251_not
g25266 not n4232 ; n4232_not
g25267 not n8102 ; n8102_not
g25268 not n3413 ; n3413_not
g25269 not n3035 ; n3035_not
g25270 not n1631 ; n1631_not
g25271 not n3350 ; n3350_not
g25272 not n6150 ; n6150_not
g25273 not n3603 ; n3603_not
g25274 not n1092 ; n1092_not
g25275 not n1407 ; n1407_not
g25276 not n1704 ; n1704_not
g25277 not n2370 ; n2370_not
g25278 not n2352 ; n2352_not
g25279 not n5070 ; n5070_not
g25280 not n2343 ; n2343_not
g25281 not n3306 ; n3306_not
g25282 not n1209 ; n1209_not
g25283 not n4620 ; n4620_not
g25284 not n2145 ; n2145_not
g25285 not n4125 ; n4125_not
g25286 not n9111 ; n9111_not
g25287 not n3162 ; n3162_not
g25288 not n4134 ; n4134_not
g25289 not n2172 ; n2172_not
g25290 not n3351 ; n3351_not
g25291 not n7032 ; n7032_not
g25292 not n2244 ; n2244_not
g25293 not n1443 ; n1443_not
g25294 not n8040 ; n8040_not
g25295 not n2208 ; n2208_not
g25296 not n2280 ; n2280_not
g25297 not n6141 ; n6141_not
g25298 not n1254 ; n1254_not
g25299 not n6321 ; n6321_not
g25300 not n5061 ; n5061_not
g25301 not n2316 ; n2316_not
g25302 not n3072 ; n3072_not
g25303 not n2622 ; n2622_not
g25304 not n5241 ; n5241_not
g25305 not n9102 ; n9102_not
g25306 not n4431 ; n4431_not
g25307 not n8400 ; n8400_not
g25308 not n1722 ; n1722_not
g25309 not n2604 ; n2604_not
g25310 not n4206 ; n4206_not
g25311 not n1344 ; n1344_not
g25312 not n1335 ; n1335_not
g25313 not n2631 ; n2631_not
g25314 not n5133 ; n5133_not
g25315 not n5142 ; n5142_not
g25316 not n2406 ; n2406_not
g25317 not n1326 ; n1326_not
g25318 not n2541 ; n2541_not
g25319 not n2550 ; n2550_not
g25320 not n4503 ; n4503_not
g25321 not n6042 ; n6042_not
g25322 not n6033 ; n6033_not
g25323 not n2433 ; n2433_not
g25324 not n8031 ; n8031_not
g25325 not n2703 ; n2703_not
g25326 not n1290 ; n1290_not
g25327 not n4161 ; n4161_not
g25328 not n4170 ; n4170_not
g25329 not n1137 ; n1137_not
g25330 not n6411 ; n6411_not
g25331 not n2505 ; n2505_not
g25332 not n2514 ; n2514_not
g25333 not n1128 ; n1128_not
g25334 not n4323 ; n4323_not
g25335 not n3153 ; n3153_not
g25336 not n3333 ; n3333_not
g25337 not n6114 ; n6114_not
g25338 not n6105 ; n6105_not
g25339 not n3342 ; n3342_not
g25340 not n5106 ; n5106_not
g25341 not n4251 ; n4251_not
g25342 not n3423 ; n3423_not
g25343 not n2820 ; n2820_not
g25344 not n7401 ; n7401_not
g25345 not n5511 ; n5511_not
g25346 not n2334 ; n2334_not
g25347 not n3360 ; n3360_not
g25348 not n1182 ; n1182_not
g25349 not n3900 ; n3900_not
g25350 not n2811 ; n2811_not
g25351 not n9003 ; n9003_not
g25352 not n2019 ; n2019_not
g25353 not n1641 ; n1641_not
g25354 not n8013 ; n8013_not
g25355 not n1632 ; n1632_not
g25356 not n1830 ; n1830_not
g25357 not n2055 ; n2055_not
g25358 not n3225 ; n3225_not
g25359 not n5034 ; n5034_not
g25360 not n5025 ; n5025_not
g25361 not n4017 ; n4017_not
g25362 not n7221 ; n7221_not
g25363 not n7104 ; n7104_not
g25364 not n8112 ; n8112_not
g25365 not n2091 ; n2091_not
g25366 not n5601 ; n5601_not
g25367 not n6330 ; n6330_not
g25368 not n5205 ; n5205_not
g25369 not n1605 ; n1605_not
g25370 not n8220 ; n8220_not
g25371 not n5331 ; n5331_not
g25372 not n7212 ; n7212_not
g25373 not n1191 ; n1191_not
g25374 not n8004 ; n8004_not
g25375 not n3531 ; n3531_not
g25376 not n4800 ; n4800_not
g25377 not n3270 ; n3270_not
g25378 not n9030 ; n9030_not
g25379 not n6213 ; n6213_not
g25380 not n1560 ; n1560_not
g25381 not n4053 ; n4053_not
g25382 not n6222 ; n6222_not
g25383 not n3234 ; n3234_not
g25384 not n3261 ; n3261_not
g25385 not n4062 ; n4062_not
g25386 not n4260 ; n4260_not
g25387 not n1371 ; n1371_not
g25388 not n5403 ; n5403_not
g25389 not n3720 ; n3720_not
g25390 not n9210 ; n9210_not
g25391 not n5700 ; n5700_not
g25392 not n3036 ; n3036_not
g25393 not n4026 ; n4026_not
g25394 not n7330 ; n7330_not
g25395 not n3424 ; n3424_not
g25396 not n2146 ; n2146_not
g25397 not n2335 ; n2335_not
g25398 not n3118 ; n3118_not
g25399 not n2128 ; n2128_not
g25400 not n8041 ; n8041_not
g25401 not n3730 ; n3730_not
g25402 not n3406 ; n3406_not
g25403 not n7033 ; n7033_not
g25404 not n2119 ; n2119_not
g25405 not n1543 ; n1543_not
g25406 not n1516 ; n1516_not
g25407 not n3163 ; n3163_not
g25408 not n1291 ; n1291_not
g25409 not n3532 ; n3532_not
g25410 not n6223 ; n6223_not
g25411 not n2254 ; n2254_not
g25412 not n2245 ; n2245_not
g25413 not n1408 ; n1408_not
g25414 not n7402 ; n7402_not
g25415 not n1417 ; n1417_not
g25416 not n3910 ; n3910_not
g25417 not n1606 ; n1606_not
g25418 not n4135 ; n4135_not
g25419 not n2515 ; n2515_not
g25420 not n2281 ; n2281_not
g25421 not n2290 ; n2290_not
g25422 not n9004 ; n9004_not
g25423 not n4324 ; n4324_not
g25424 not n9220 ; n9220_not
g25425 not n3109 ; n3109_not
g25426 not n1570 ; n1570_not
g25427 not n6331 ; n6331_not
g25428 not n1480 ; n1480_not
g25429 not n2551 ; n2551_not
g25430 not n2326 ; n2326_not
g25431 not n2317 ; n2317_not
g25432 not n4504 ; n4504_not
g25433 not n7231 ; n7231_not
g25434 not n1561 ; n1561_not
g25435 not n2704 ; n2704_not
g25436 not n8401 ; n8401_not
g25437 not n5332 ; n5332_not
g25438 not n5512 ; n5512_not
g25439 not n3091 ; n3091_not
g25440 not n1453 ; n1453_not
g25441 not n6412 ; n6412_not
g25442 not n3802 ; n3802_not
g25443 not n2740 ; n2740_not
g25444 not n5143 ; n5143_not
g25445 not n5710 ; n5710_not
g25446 not n1048 ; n1048_not
g25447 not n5701 ; n5701_not
g25448 not n4207 ; n4207_not
g25449 not n4360 ; n4360_not
g25450 not n8104 ; n8104_not
g25451 not n1534 ; n1534_not
g25452 not n6043 ; n6043_not
g25453 not n4540 ; n4540_not
g25454 not n8014 ; n8014_not
g25455 not n8221 ; n8221_not
g25456 not n1723 ; n1723_not
g25457 not n2632 ; n2632_not
g25458 not n2812 ; n2812_not
g25459 not n3352 ; n3352_not
g25460 not n3361 ; n3361_not
g25461 not n6700 ; n6700_not
g25462 not n3901 ; n3901_not
g25463 not n7222 ; n7222_not
g25464 not n1138 ; n1138_not
g25465 not n1642 ; n1642_not
g25466 not n2155 ; n2155_not
g25467 not n1327 ; n1327_not
g25468 not n1444 ; n1444_not
g25469 not n3046 ; n3046_not
g25470 not n3271 ; n3271_not
g25471 not n4171 ; n4171_not
g25472 not n9040 ; n9040_not
g25473 not n1255 ; n1255_not
g25474 not n5404 ; n5404_not
g25475 not n2092 ; n2092_not
g25476 not n6340 ; n6340_not
g25477 not n2371 ; n2371_not
g25478 not n4621 ; n4621_not
g25479 not n1057 ; n1057_not
g25480 not n1219 ; n1219_not
g25481 not n7411 ; n7411_not
g25482 not n5440 ; n5440_not
g25483 not n1039 ; n1039_not
g25484 not n3460 ; n3460_not
g25485 not n3604 ; n3604_not
g25486 not n1732 ; n1732_not
g25487 not n2605 ; n2605_not
g25488 not n4432 ; n4432_not
g25489 not n4900 ; n4900_not
g25490 not n2902 ; n2902_not
g25491 not n5071 ; n5071_not
g25492 not n5215 ; n5215_not
g25493 not n4630 ; n4630_not
g25494 not n7510 ; n7510_not
g25495 not n4810 ; n4810_not
g25496 not n3721 ; n3721_not
g25497 not n5107 ; n5107_not
g25498 not n2344 ; n2344_not
g25499 not n1831 ; n1831_not
g25500 not n9112 ; n9112_not
g25501 not n2182 ; n2182_not
g25502 not n2173 ; n2173_not
g25503 not n7105 ; n7105_not
g25504 not n1318 ; n1318_not
g25505 not n4270 ; n4270_not
g25506 not n6520 ; n6520_not
g25507 not n8113 ; n8113_not
g25508 not n4027 ; n4027_not
g25509 not n2443 ; n2443_not
g25510 not n4603 ; n4603_not
g25511 not n2209 ; n2209_not
g25512 not n2218 ; n2218_not
g25513 not n4801 ; n4801_not
g25514 not n3235 ; n3235_not
g25515 not n5035 ; n5035_not
g25516 not n4702 ; n4702_not
g25517 not n3307 ; n3307_not
g25518 not n7303 ; n7303_not
g25519 not n3343 ; n3343_not
g25520 not n3037 ; n3037_not
g25521 not n6151 ; n6151_not
g25522 not n4063 ; n4063_not
g25523 not n2407 ; n2407_not
g25524 not n2056 ; n2056_not
g25525 not n6115 ; n6115_not
g25526 not n3272 ; n3272_not
g25527 not n7142 ; n7142_not
g25528 not n2570 ; n2570_not
g25529 not n2642 ; n2642_not
g25530 not n2831 ; n2831_not
g25531 not n3731 ; n3731_not
g25532 not n5243 ; n5243_not
g25533 not n2840 ; n2840_not
g25534 not n3236 ; n3236_not
g25535 not n6224 ; n6224_not
g25536 not n3047 ; n3047_not
g25537 not n4028 ; n4028_not
g25538 not n3470 ; n3470_not
g25539 not n3128 ; n3128_not
g25540 not n8150 ; n8150_not
g25541 not n2741 ; n2741_not
g25542 not n6152 ; n6152_not
g25543 not n8051 ; n8051_not
g25544 not n2903 ; n2903_not
g25545 not n5207 ; n5207_not
g25546 not n7304 ; n7304_not
g25547 not n6332 ; n6332_not
g25548 not n2750 ; n2750_not
g25549 not n8420 ; n8420_not
g25550 not n8114 ; n8114_not
g25551 not n2714 ; n2714_not
g25552 not n7232 ; n7232_not
g25553 not n2705 ; n2705_not
g25554 not n5234 ; n5234_not
g25555 not n2633 ; n2633_not
g25556 not n3461 ; n3461_not
g25557 not n8123 ; n8123_not
g25558 not n3344 ; n3344_not
g25559 not n8600 ; n8600_not
g25560 not n3164 ; n3164_not
g25561 not n6260 ; n6260_not
g25562 not n6116 ; n6116_not
g25563 not n3308 ; n3308_not
g25564 not n7160 ; n7160_not
g25565 not n8042 ; n8042_not
g25566 not n1742 ; n1742_not
g25567 not n1706 ; n1706_not
g25568 not n1715 ; n1715_not
g25569 not n1733 ; n1733_not
g25570 not n1724 ; n1724_not
g25571 not n9113 ; n9113_not
g25572 not n7070 ; n7070_not
g25573 not n7106 ; n7106_not
g25574 not n7115 ; n7115_not
g25575 not n7520 ; n7520_not
g25576 not n1643 ; n1643_not
g25577 not n3641 ; n3641_not
g25578 not n5441 ; n5441_not
g25579 not n1607 ; n1607_not
g25580 not n5450 ; n5450_not
g25581 not n1373 ; n1373_not
g25582 not n1571 ; n1571_not
g25583 not n6602 ; n6602_not
g25584 not n8402 ; n8402_not
g25585 not n4811 ; n4811_not
g25586 not n1922 ; n1922_not
g25587 not n1904 ; n1904_not
g25588 not n5333 ; n5333_not
g25589 not n4505 ; n4505_not
g25590 not n4550 ; n4550_not
g25591 not n4541 ; n4541_not
g25592 not n4901 ; n4901_not
g25593 not n4136 ; n4136_not
g25594 not n3542 ; n3542_not
g25595 not n3533 ; n3533_not
g25596 not n5252 ; n5252_not
g25597 not n5342 ; n5342_not
g25598 not n5270 ; n5270_not
g25599 not n1544 ; n1544_not
g25600 not n5711 ; n5711_not
g25601 not n5306 ; n5306_not
g25602 not n5072 ; n5072_not
g25603 not n5414 ; n5414_not
g25604 not n7007 ; n7007_not
g25605 not n5180 ; n5180_not
g25606 not n9005 ; n9005_not
g25607 not n3614 ; n3614_not
g25608 not n4064 ; n4064_not
g25609 not n3605 ; n3605_not
g25610 not n3911 ; n3911_not
g25611 not n1139 ; n1139_not
g25612 not n1067 ; n1067_not
g25613 not n1049 ; n1049_not
g25614 not n5108 ; n5108_not
g25615 not n6521 ; n6521_not
g25616 not n6530 ; n6530_not
g25617 not n9041 ; n9041_not
g25618 not n5144 ; n5144_not
g25619 not n5603 ; n5603_not
g25620 not n1346 ; n1346_not
g25621 not n1490 ; n1490_not
g25622 not n1292 ; n1292_not
g25623 not n1454 ; n1454_not
g25624 not n5216 ; n5216_not
g25625 not n7412 ; n7412_not
g25626 not n1256 ; n1256_not
g25627 not n1265 ; n1265_not
g25628 not n1418 ; n1418_not
g25629 not n1229 ; n1229_not
g25630 not n5036 ; n5036_not
g25631 not n1364 ; n1364_not
g25632 not n6413 ; n6413_not
g25633 not n1355 ; n1355_not
g25634 not n6422 ; n6422_not
g25635 not n5405 ; n5405_not
g25636 not n4631 ; n4631_not
g25637 not n7340 ; n7340_not
g25638 not n2345 ; n2345_not
g25639 not n2336 ; n2336_not
g25640 not n2327 ; n2327_not
g25641 not n4172 ; n4172_not
g25642 not n2093 ; n2093_not
g25643 not n2291 ; n2291_not
g25644 not n2057 ; n2057_not
g25645 not n6080 ; n6080_not
g25646 not n2066 ; n2066_not
g25647 not n3425 ; n3425_not
g25648 not n2255 ; n2255_not
g25649 not n3434 ; n3434_not
g25650 not n2219 ; n2219_not
g25651 not n8303 ; n8303_not
g25652 not n4334 ; n4334_not
g25653 not n5630 ; n5630_not
g25654 not n4325 ; n4325_not
g25655 not n2552 ; n2552_not
g25656 not n7601 ; n7601_not
g25657 not n9410 ; n9410_not
g25658 not n2516 ; n2516_not
g25659 not n5621 ; n5621_not
g25660 not n7043 ; n7043_not
g25661 not n2480 ; n2480_not
g25662 not n2606 ; n2606_not
g25663 not n6044 ; n6044_not
g25664 not n2444 ; n2444_not
g25665 not n5513 ; n5513_not
g25666 not n2408 ; n2408_not
g25667 not n2615 ; n2615_not
g25668 not n2390 ; n2390_not
g25669 not n5522 ; n5522_not
g25670 not n2372 ; n2372_not
g25671 not n7034 ; n7034_not
g25672 not n1832 ; n1832_not
g25673 not n1841 ; n1841_not
g25674 not n4406 ; n4406_not
g25675 not n1805 ; n1805_not
g25676 not n8231 ; n8231_not
g25677 not n8222 ; n8222_not
g25678 not n4208 ; n4208_not
g25679 not n8024 ; n8024_not
g25680 not n3506 ; n3506_not
g25681 not n8015 ; n8015_not
g25682 not n1760 ; n1760_not
g25683 not n6008 ; n6008_not
g25684 not n9221 ; n9221_not
g25685 not n4433 ; n4433_not
g25686 not n4442 ; n4442_not
g25687 not n8411 ; n8411_not
g25688 not n1931 ; n1931_not
g25689 not n3803 ; n3803_not
g25690 not n5612 ; n5612_not
g25691 not n2183 ; n2183_not
g25692 not n6710 ; n6710_not
g25693 not n2435 ; n2435_not
g25694 not n2147 ; n2147_not
g25695 not n6701 ; n6701_not
g25696 not n4361 ; n4361_not
g25697 not n4370 ; n4370_not
g25698 not n8330 ; n8330_not
g25699 not n4703 ; n4703_not
g25700 not n8430 ; n8430_not
g25701 not n9303 ; n9303_not
g25702 not n8421 ; n8421_not
g25703 not n7341 ; n7341_not
g25704 not n3372 ; n3372_not
g25705 not n3363 ; n3363_not
g25706 not n3381 ; n3381_not
g25707 not n5622 ; n5622_not
g25708 not n3390 ; n3390_not
g25709 not n8412 ; n8412_not
g25710 not n3237 ; n3237_not
g25711 not n3246 ; n3246_not
g25712 not n3543 ; n3543_not
g25713 not n6009 ; n6009_not
g25714 not n3273 ; n3273_not
g25715 not n3282 ; n3282_not
g25716 not n9006 ; n9006_not
g25717 not n3507 ; n3507_not
g25718 not n9015 ; n9015_not
g25719 not n3318 ; n3318_not
g25720 not n3309 ; n3309_not
g25721 not n3615 ; n3615_not
g25722 not n3732 ; n3732_not
g25723 not n3471 ; n3471_not
g25724 not n8232 ; n8232_not
g25725 not n9231 ; n9231_not
g25726 not n9222 ; n9222_not
g25727 not n7413 ; n7413_not
g25728 not n3165 ; n3165_not
g25729 not n3174 ; n3174_not
g25730 not n5640 ; n5640_not
g25731 not n3435 ; n3435_not
g25732 not n3138 ; n3138_not
g25733 not n6225 ; n6225_not
g25734 not n6234 ; n6234_not
g25735 not n4812 ; n4812_not
g25736 not n7080 ; n7080_not
g25737 not n5712 ; n5712_not
g25738 not n6270 ; n6270_not
g25739 not n5343 ; n5343_not
g25740 not n6261 ; n6261_not
g25741 not n1680 ; n1680_not
g25742 not n6306 ; n6306_not
g25743 not n1644 ; n1644_not
g25744 not n1653 ; n1653_not
g25745 not n5307 ; n5307_not
g25746 not n1842 ; n1842_not
g25747 not n6711 ; n6711_not
g25748 not n1617 ; n1617_not
g25749 not n1608 ; n1608_not
g25750 not n1806 ; n1806_not
g25751 not n3840 ; n3840_not
g25752 not n1572 ; n1572_not
g25753 not n1581 ; n1581_not
g25754 not n4290 ; n4290_not
g25755 not n6531 ; n6531_not
g25756 not n2328 ; n2328_not
g25757 not n2292 ; n2292_not
g25758 not n2256 ; n2256_not
g25759 not n6153 ; n6153_not
g25760 not n6162 ; n6162_not
g25761 not n5415 ; n5415_not
g25762 not n7116 ; n7116_not
g25763 not n3804 ; n3804_not
g25764 not n2184 ; n2184_not
g25765 not n2166 ; n2166_not
g25766 not n1932 ; n1932_not
g25767 not n5046 ; n5046_not
g25768 not n5037 ; n5037_not
g25769 not n4704 ; n4704_not
g25770 not n9042 ; n9042_not
g25771 not n2067 ; n2067_not
g25772 not n4740 ; n4740_not
g25773 not n6603 ; n6603_not
g25774 not n8016 ; n8016_not
g25775 not n5217 ; n5217_not
g25776 not n5235 ; n5235_not
g25777 not n1518 ; n1518_not
g25778 not n1491 ; n1491_not
g25779 not n9114 ; n9114_not
g25780 not n1455 ; n1455_not
g25781 not n1419 ; n1419_not
g25782 not n1383 ; n1383_not
g25783 not n1365 ; n1365_not
g25784 not n1176 ; n1176_not
g25785 not n5820 ; n5820_not
g25786 not n1266 ; n1266_not
g25787 not n1077 ; n1077_not
g25788 not n3912 ; n3912_not
g25789 not n1194 ; n1194_not
g25790 not n1068 ; n1068_not
g25791 not n7521 ; n7521_not
g25792 not n6900 ; n6900_not
g25793 not n1770 ; n1770_not
g25794 not n6351 ; n6351_not
g25795 not n7044 ; n7044_not
g25796 not n1734 ; n1734_not
g25797 not n1509 ; n1509_not
g25798 not n5271 ; n5271_not
g25799 not n1707 ; n1707_not
g25800 not n8304 ; n8304_not
g25801 not n9600 ; n9600_not
g25802 not n9123 ; n9123_not
g25803 not n5244 ; n5244_not
g25804 not n7008 ; n7008_not
g25805 not n8340 ; n8340_not
g25806 not n1554 ; n1554_not
g25807 not n1527 ; n1527_not
g25808 not n1545 ; n1545_not
g25809 not n4065 ; n4065_not
g25810 not n2940 ; n2940_not
g25811 not n8601 ; n8601_not
g25812 not n5181 ; n5181_not
g25813 not n4407 ; n4407_not
g25814 not n2904 ; n2904_not
g25815 not n9420 ; n9420_not
g25816 not n5523 ; n5523_not
g25817 not n2850 ; n2850_not
g25818 not n4443 ; n4443_not
g25819 not n9150 ; n9150_not
g25820 not n4146 ; n4146_not
g25821 not n4137 ; n4137_not
g25822 not n6360 ; n6360_not
g25823 not n2571 ; n2571_not
g25824 not n5145 ; n5145_not
g25825 not n2562 ; n2562_not
g25826 not n2553 ; n2553_not
g25827 not n5154 ; n5154_not
g25828 not n2517 ; n2517_not
g25829 not n3930 ; n3930_not
g25830 not n4245 ; n4245_not
g25831 not n4263 ; n4263_not
g25832 not n7305 ; n7305_not
g25833 not n4272 ; n4272_not
g25834 not n8160 ; n8160_not
g25835 not n7710 ; n7710_not
g25836 not n3129 ; n3129_not
g25837 not n5226 ; n5226_not
g25838 not n4335 ; n4335_not
g25839 not n3048 ; n3048_not
g25840 not n4029 ; n4029_not
g25841 not n7233 ; n7233_not
g25842 not n4038 ; n4038_not
g25843 not n8124 ; n8124_not
g25844 not n4371 ; n4371_not
g25845 not n5190 ; n5190_not
g25846 not n4074 ; n4074_not
g25847 not n4209 ; n4209_not
g25848 not n2607 ; n2607_not
g25849 not n6081 ; n6081_not
g25850 not n6090 ; n6090_not
g25851 not n4551 ; n4551_not
g25852 not n2580 ; n2580_not
g25853 not n4560 ; n4560_not
g25854 not n5118 ; n5118_not
g25855 not n5109 ; n5109_not
g25856 not n5451 ; n5451_not
g25857 not n8052 ; n8052_not
g25858 not n7611 ; n7611_not
g25859 not n5073 ; n5073_not
g25860 not n5082 ; n5082_not
g25861 not n6126 ; n6126_not
g25862 not n2148 ; n2148_not
g25863 not n6117 ; n6117_not
g25864 not n4614 ; n4614_not
g25865 not n4632 ; n4632_not
g25866 not n2526 ; n2526_not
g25867 not n6018 ; n6018_not
g25868 not n2751 ; n2751_not
g25869 not n2490 ; n2490_not
g25870 not n2481 ; n2481_not
g25871 not n2715 ; n2715_not
g25872 not n6423 ; n6423_not
g25873 not n7602 ; n7602_not
g25874 not n2445 ; n2445_not
g25875 not n2454 ; n2454_not
g25876 not n4173 ; n4173_not
g25877 not n4218 ; n4218_not
g25878 not n7170 ; n7170_not
g25879 not n4515 ; n4515_not
g25880 not n2643 ; n2643_not
g25881 not n6045 ; n6045_not
g25882 not n6054 ; n6054_not
g25883 not n2409 ; n2409_not
g25884 not n2418 ; n2418_not
g25885 not n8305 ; n8305_not
g25886 not n9304 ; n9304_not
g25887 not n4039 ; n4039_not
g25888 not n3706 ; n3706_not
g25889 not n8341 ; n8341_not
g25890 not n3643 ; n3643_not
g25891 not n3634 ; n3634_not
g25892 not n3940 ; n3940_not
g25893 not n5236 ; n5236_not
g25894 not n7414 ; n7414_not
g25895 not n5245 ; n5245_not
g25896 not n4903 ; n4903_not
g25897 not n7270 ; n7270_not
g25898 not n7450 ; n7450_not
g25899 not n7900 ; n7900_not
g25900 not n4921 ; n4921_not
g25901 not n4912 ; n4912_not
g25902 not n5290 ; n5290_not
g25903 not n7243 ; n7243_not
g25904 not n4930 ; n4930_not
g25905 not n7234 ; n7234_not
g25906 not n5308 ; n5308_not
g25907 not n7522 ; n7522_not
g25908 not n7531 ; n7531_not
g25909 not n4507 ; n4507_not
g25910 not n5344 ; n5344_not
g25911 not n7315 ; n7315_not
g25912 not n5119 ; n5119_not
g25913 not n7351 ; n7351_not
g25914 not n5155 ; n5155_not
g25915 not n4822 ; n4822_not
g25916 not n4741 ; n4741_not
g25917 not n4750 ; n4750_not
g25918 not n4813 ; n4813_not
g25919 not n5083 ; n5083_not
g25920 not n7342 ; n7342_not
g25921 not n7306 ; n7306_not
g25922 not n4714 ; n4714_not
g25923 not n4705 ; n4705_not
g25924 not n5047 ; n5047_not
g25925 not n5191 ; n5191_not
g25926 not n7720 ; n7720_not
g25927 not n4642 ; n4642_not
g25928 not n4633 ; n4633_not
g25929 not n5227 ; n5227_not
g25930 not n7423 ; n7423_not
g25931 not n8161 ; n8161_not
g25932 not n7144 ; n7144_not
g25933 not n3931 ; n3931_not
g25934 not n3913 ; n3913_not
g25935 not n3922 ; n3922_not
g25936 not n4219 ; n4219_not
g25937 not n4183 ; n4183_not
g25938 not n3841 ; n3841_not
g25939 not n3850 ; n3850_not
g25940 not n4147 ; n4147_not
g25941 not n8233 ; n8233_not
g25942 not n5641 ; n5641_not
g25943 not n3814 ; n3814_not
g25944 not n3805 ; n3805_not
g25945 not n7135 ; n7135_not
g25946 not n5272 ; n5272_not
g25947 not n4075 ; n4075_not
g25948 not n3742 ; n3742_not
g25949 not n3733 ; n3733_not
g25950 not n9421 ; n9421_not
g25951 not n7207 ; n7207_not
g25952 not n5380 ; n5380_not
g25953 not n7612 ; n7612_not
g25954 not n5416 ; n5416_not
g25955 not n8035 ; n8035_not
g25956 not n8053 ; n8053_not
g25957 not n7603 ; n7603_not
g25958 not n4273 ; n4273_not
g25959 not n5452 ; n5452_not
g25960 not n4552 ; n4552_not
g25961 not n4516 ; n4516_not
g25962 not n4480 ; n4480_not
g25963 not n5524 ; n5524_not
g25964 not n4444 ; n4444_not
g25965 not n4408 ; n4408_not
g25966 not n8125 ; n8125_not
g25967 not n4372 ; n4372_not
g25968 not n5560 ; n5560_not
g25969 not n4336 ; n4336_not
g25970 not n3472 ; n3472_not
g25971 not n8017 ; n8017_not
g25972 not n3436 ; n3436_not
g25973 not n1807 ; n1807_not
g25974 not n9124 ; n9124_not
g25975 not n6055 ; n6055_not
g25976 not n1843 ; n1843_not
g25977 not n6712 ; n6712_not
g25978 not n3382 ; n3382_not
g25979 not n3085 ; n3085_not
g25980 not n6091 ; n6091_not
g25981 not n5713 ; n5713_not
g25982 not n5722 ; n5722_not
g25983 not n3049 ; n3049_not
g25984 not n3058 ; n3058_not
g25985 not n3319 ; n3319_not
g25986 not n1690 ; n1690_not
g25987 not n1708 ; n1708_not
g25988 not n1726 ; n1726_not
g25989 not n6532 ; n6532_not
g25990 not n3616 ; n3616_not
g25991 not n1753 ; n1753_not
g25992 not n7045 ; n7045_not
g25993 not n2347 ; n2347_not
g25994 not n3580 ; n3580_not
g25995 not n2365 ; n2365_not
g25996 not n1771 ; n1771_not
g25997 not n2356 ; n2356_not
g25998 not n3544 ; n3544_not
g25999 not n3508 ; n3508_not
g26000 not n2608 ; n2608_not
g26001 not n6019 ; n6019_not
g26002 not n5650 ; n5650_not
g26003 not n1942 ; n1942_not
g26004 not n1906 ; n1906_not
g26005 not n1960 ; n1960_not
g26006 not n1735 ; n1735_not
g26007 not n6640 ; n6640_not
g26008 not n8710 ; n8710_not
g26009 not n3139 ; n3139_not
g26010 not n7117 ; n7117_not
g26011 not n5902 ; n5902_not
g26012 not n6271 ; n6271_not
g26013 not n5830 ; n5830_not
g26014 not n5821 ; n5821_not
g26015 not n6604 ; n6604_not
g26016 not n6235 ; n6235_not
g26017 not n2068 ; n2068_not
g26018 not n3283 ; n3283_not
g26019 not n6307 ; n6307_not
g26020 not n1951 ; n1951_not
g26021 not n6127 ; n6127_not
g26022 not n3247 ; n3247_not
g26023 not n9160 ; n9160_not
g26024 not n2950 ; n2950_not
g26025 not n2941 ; n2941_not
g26026 not n7081 ; n7081_not
g26027 not n9232 ; n9232_not
g26028 not n1933 ; n1933_not
g26029 not n1915 ; n1915_not
g26030 not n2905 ; n2905_not
g26031 not n2914 ; n2914_not
g26032 not n3175 ; n3175_not
g26033 not n6163 ; n6163_not
g26034 not n6901 ; n6901_not
g26035 not n7171 ; n7171_not
g26036 not n1519 ; n1519_not
g26037 not n1492 ; n1492_not
g26038 not n2266 ; n2266_not
g26039 not n9052 ; n9052_not
g26040 not n9601 ; n9601_not
g26041 not n2581 ; n2581_not
g26042 not n2572 ; n2572_not
g26043 not n1384 ; n1384_not
g26044 not n2752 ; n2752_not
g26045 not n6424 ; n6424_not
g26046 not n2716 ; n2716_not
g26047 not n2563 ; n2563_not
g26048 not n2680 ; n2680_not
g26049 not n9016 ; n9016_not
g26050 not n2527 ; n2527_not
g26051 not n1267 ; n1267_not
g26052 not n6730 ; n6730_not
g26053 not n1069 ; n1069_not
g26054 not n6460 ; n6460_not
g26055 not n2293 ; n2293_not
g26056 not n2644 ; n2644_not
g26057 not n8530 ; n8530_not
g26058 not n2374 ; n2374_not
g26059 not n2626 ; n2626_not
g26060 not n1078 ; n1078_not
g26061 not n7180 ; n7180_not
g26062 not n8503 ; n8503_not
g26063 not n1654 ; n1654_not
g26064 not n2419 ; n2419_not
g26065 not n1465 ; n1465_not
g26066 not n2185 ; n2185_not
g26067 not n3670 ; n3670_not
g26068 not n1456 ; n1456_not
g26069 not n8611 ; n8611_not
g26070 not n3652 ; n3652_not
g26071 not n1618 ; n1618_not
g26072 not n1429 ; n1429_not
g26073 not n2455 ; n2455_not
g26074 not n7153 ; n7153_not
g26075 not n2257 ; n2257_not
g26076 not n1546 ; n1546_not
g26077 not n8413 ; n8413_not
g26078 not n7009 ; n7009_not
g26079 not n2491 ; n2491_not
g26080 not n1393 ; n1393_not
g26081 not n1582 ; n1582_not
g26082 not n8602 ; n8602_not
g26083 not n4238 ; n4238_not
g26084 not n4247 ; n4247_not
g26085 not n8306 ; n8306_not
g26086 not n2564 ; n2564_not
g26087 not n9530 ; n9530_not
g26088 not n4373 ; n4373_not
g26089 not n8342 ; n8342_not
g26090 not n4715 ; n4715_not
g26091 not n1880 ; n1880_not
g26092 not n4382 ; n4382_not
g26093 not n9044 ; n9044_not
g26094 not n7136 ; n7136_not
g26095 not n2384 ; n2384_not
g26096 not n2366 ; n2366_not
g26097 not n2456 ; n2456_not
g26098 not n2078 ; n2078_not
g26099 not n2069 ; n2069_not
g26100 not n4571 ; n4571_not
g26101 not n2492 ; n2492_not
g26102 not n2267 ; n2267_not
g26103 not n4643 ; n4643_not
g26104 not n6713 ; n6713_not
g26105 not n6722 ; n6722_not
g26106 not n4580 ; n4580_not
g26107 not n2195 ; n2195_not
g26108 not n1961 ; n1961_not
g26109 not n1970 ; n1970_not
g26110 not n7118 ; n7118_not
g26111 not n4337 ; n4337_not
g26112 not n2528 ; n2528_not
g26113 not n4346 ; n4346_not
g26114 not n7613 ; n7613_not
g26115 not n8315 ; n8315_not
g26116 not n1358 ; n1358_not
g26117 not n1178 ; n1178_not
g26118 not n1367 ; n1367_not
g26119 not n5048 ; n5048_not
g26120 not n1394 ; n1394_not
g26121 not n1268 ; n1268_not
g26122 not n1277 ; n1277_not
g26123 not n1466 ; n1466_not
g26124 not n9611 ; n9611_not
g26125 not n5228 ; n5228_not
g26126 not n9602 ; n9602_not
g26127 not n1565 ; n1565_not
g26128 not n1583 ; n1583_not
g26129 not n1385 ; n1385_not
g26130 not n6605 ; n6605_not
g26131 not n1619 ; n1619_not
g26132 not n1655 ; n1655_not
g26133 not n7721 ; n7721_not
g26134 not n6506 ; n6506_not
g26135 not n5156 ; n5156_not
g26136 not n9710 ; n9710_not
g26137 not n9053 ; n9053_not
g26138 not n6470 ; n6470_not
g26139 not n6461 ; n6461_not
g26140 not n6533 ; n6533_not
g26141 not n9017 ; n9017_not
g26142 not n1079 ; n1079_not
g26143 not n6542 ; n6542_not
g26144 not n1187 ; n1187_not
g26145 not n5084 ; n5084_not
g26146 not n5192 ; n5192_not
g26147 not n6425 ; n6425_not
g26148 not n6434 ; n6434_not
g26149 not n1169 ; n1169_not
g26150 not n1907 ; n1907_not
g26151 not n9161 ; n9161_not
g26152 not n4823 ; n4823_not
g26153 not n4490 ; n4490_not
g26154 not n4481 ; n4481_not
g26155 not n1934 ; n1934_not
g26156 not n4445 ; n4445_not
g26157 not n4454 ; n4454_not
g26158 not n1772 ; n1772_not
g26159 not n1781 ; n1781_not
g26160 not n4751 ; n4751_not
g26161 not n4418 ; n4418_not
g26162 not n4409 ; n4409_not
g26163 not n8351 ; n8351_not
g26164 not n1817 ; n1817_not
g26165 not n1808 ; n1808_not
g26166 not n1844 ; n1844_not
g26167 not n1853 ; n1853_not
g26168 not n4940 ; n4940_not
g26169 not n6614 ; n6614_not
g26170 not n1691 ; n1691_not
g26171 not n7901 ; n7901_not
g26172 not n4922 ; n4922_not
g26173 not n1547 ; n1547_not
g26174 not n9125 ; n9125_not
g26175 not n6740 ; n6740_not
g26176 not n6731 ; n6731_not
g26177 not n6650 ; n6650_not
g26178 not n6641 ; n6641_not
g26179 not n8432 ; n8432_not
g26180 not n4517 ; n4517_not
g26181 not n4526 ; n4526_not
g26182 not n4184 ; n4184_not
g26183 not n5642 ; n5642_not
g26184 not n4148 ; n4148_not
g26185 not n7352 ; n7352_not
g26186 not n5624 ; n5624_not
g26187 not n8450 ; n8450_not
g26188 not n3635 ; n3635_not
g26189 not n3617 ; n3617_not
g26190 not n3644 ; n3644_not
g26191 not n8441 ; n8441_not
g26192 not n5651 ; n5651_not
g26193 not n3671 ; n3671_not
g26194 not n5309 ; n5309_not
g26195 not n4076 ; n4076_not
g26196 not n5318 ; n5318_not
g26197 not n7424 ; n7424_not
g26198 not n7019 ; n7019_not
g26199 not n5561 ; n5561_not
g26200 not n4283 ; n4283_not
g26201 not n3176 ; n3176_not
g26202 not n4256 ; n4256_not
g26203 not n4274 ; n4274_not
g26204 not n6164 ; n6164_not
g26205 not n8063 ; n8063_not
g26206 not n8054 ; n8054_not
g26207 not n3248 ; n3248_not
g26208 not n8504 ; n8504_not
g26209 not n5615 ; n5615_not
g26210 not n7316 ; n7316_not
g26211 not n6128 ; n6128_not
g26212 not n3284 ; n3284_not
g26213 not n9431 ; n9431_not
g26214 not n9422 ; n9422_not
g26215 not n6092 ; n6092_not
g26216 not n6902 ; n6902_not
g26217 not n6911 ; n6911_not
g26218 not n6056 ; n6056_not
g26219 not n7532 ; n7532_not
g26220 not n3851 ; n3851_not
g26221 not n3545 ; n3545_not
g26222 not n7091 ; n7091_not
g26223 not n5831 ; n5831_not
g26224 not n5381 ; n5381_not
g26225 not n5462 ; n5462_not
g26226 not n5390 ; n5390_not
g26227 not n5453 ; n5453_not
g26228 not n7082 ; n7082_not
g26229 not n3590 ; n3590_not
g26230 not n3581 ; n3581_not
g26231 not n5417 ; n5417_not
g26232 not n9305 ; n9305_not
g26233 not n3626 ; n3626_not
g26234 not n5426 ; n5426_not
g26235 not n3941 ; n3941_not
g26236 not n3932 ; n3932_not
g26237 not n3923 ; n3923_not
g26238 not n5570 ; n5570_not
g26239 not n3707 ; n3707_not
g26240 not n3446 ; n3446_not
g26241 not n3437 ; n3437_not
g26242 not n3743 ; n3743_not
g26243 not n5903 ; n5903_not
g26244 not n5534 ; n5534_not
g26245 not n5525 ; n5525_not
g26246 not n3473 ; n3473_not
g26247 not n3482 ; n3482_not
g26248 not n7460 ; n7460_not
g26249 not n3518 ; n3518_not
g26250 not n3509 ; n3509_not
g26251 not n3815 ; n3815_not
g26252 not n7046 ; n7046_not
g26253 not n7055 ; n7055_not
g26254 not n5354 ; n5354_not
g26255 not n5345 ; n5345_not
g26256 not n5723 ; n5723_not
g26257 not n7127 ; n7127_not
g26258 not n3059 ; n3059_not
g26259 not n8243 ; n8243_not
g26260 not n8090 ; n8090_not
g26261 not n9503 ; n9503_not
g26262 not n8126 ; n8126_not
g26263 not n2852 ; n2852_not
g26264 not n8207 ; n8207_not
g26265 not n7172 ; n7172_not
g26266 not n6272 ; n6272_not
g26267 not n2753 ; n2753_not
g26268 not n2825 ; n2825_not
g26269 not n2843 ; n2843_not
g26270 not n2690 ; n2690_not
g26271 not n2762 ; n2762_not
g26272 not n2726 ; n2726_not
g26273 not n2717 ; n2717_not
g26274 not n6308 ; n6308_not
g26275 not n8162 ; n8162_not
g26276 not n8171 ; n8171_not
g26277 not n6803 ; n6803_not
g26278 not n2951 ; n2951_not
g26279 not n2681 ; n2681_not
g26280 not n8612 ; n8612_not
g26281 not n8270 ; n8270_not
g26282 not n2870 ; n2870_not
g26283 not n2645 ; n2645_not
g26284 not n8720 ; n8720_not
g26285 not n8540 ; n8540_not
g26286 not n7280 ; n7280_not
g26287 not n7145 ; n7145_not
g26288 not n2654 ; n2654_not
g26289 not n2915 ; n2915_not
g26290 not n7208 ; n7208_not
g26291 not n7244 ; n7244_not
g26292 not n6830 ; n6830_not
g26293 not n4175 ; n4175_not
g26294 not n8234 ; n8234_not
g26295 not n8135 ; n8135_not
g26296 not n6236 ; n6236_not
g26297 not n9233 ; n9233_not
g26298 not n5427 ; n5427_not
g26299 not n4851 ; n4851_not
g26300 not n6345 ; n6345_not
g26301 not n5940 ; n5940_not
g26302 not n6129 ; n6129_not
g26303 not n9171 ; n9171_not
g26304 not n6390 ; n6390_not
g26305 not n9540 ; n9540_not
g26306 not n5904 ; n5904_not
g26307 not n6138 ; n6138_not
g26308 not n9054 ; n9054_not
g26309 not n7461 ; n7461_not
g26310 not n9162 ; n9162_not
g26311 not n7560 ; n7560_not
g26312 not n7191 ; n7191_not
g26313 not n6912 ; n6912_not
g26314 not n6471 ; n6471_not
g26315 not n7137 ; n7137_not
g26316 not n7146 ; n7146_not
g26317 not n9090 ; n9090_not
g26318 not n7128 ; n7128_not
g26319 not n6066 ; n6066_not
g26320 not n9270 ; n9270_not
g26321 not n6057 ; n6057_not
g26322 not n5832 ; n5832_not
g26323 not n7533 ; n7533_not
g26324 not n5463 ; n5463_not
g26325 not n6435 ; n6435_not
g26326 not n5760 ; n5760_not
g26327 not n6840 ; n6840_not
g26328 not n5094 ; n5094_not
g26329 not n5085 ; n5085_not
g26330 not n5157 ; n5157_not
g26331 not n6093 ; n6093_not
g26332 not n5724 ; n5724_not
g26333 not n7173 ; n7173_not
g26334 not n5166 ; n5166_not
g26335 not n6804 ; n6804_not
g26336 not n6507 ; n6507_not
g26337 not n6363 ; n6363_not
g26338 not n6318 ; n6318_not
g26339 not n9315 ; n9315_not
g26340 not n9612 ; n9612_not
g26341 not n9135 ; n9135_not
g26342 not n5319 ; n5319_not
g26343 not n7056 ; n7056_not
g26344 not n7245 ; n7245_not
g26345 not n5247 ; n5247_not
g26346 not n9126 ; n9126_not
g26347 not n6282 ; n6282_not
g26348 not n6273 ; n6273_not
g26349 not n5391 ; n5391_not
g26350 not n7317 ; n7317_not
g26351 not n5193 ; n5193_not
g26352 not n5355 ; n5355_not
g26353 not n6651 ; n6651_not
g26354 not n5571 ; n5571_not
g26355 not n9018 ; n9018_not
g26356 not n9063 ; n9063_not
g26357 not n6237 ; n6237_not
g26358 not n7281 ; n7281_not
g26359 not n6246 ; n6246_not
g26360 not n9027 ; n9027_not
g26361 not n7092 ; n7092_not
g26362 not n6615 ; n6615_not
g26363 not n9504 ; n9504_not
g26364 not n7209 ; n7209_not
g26365 not n5535 ; n5535_not
g26366 not n6543 ; n6543_not
g26367 not n9342 ; n9342_not
g26368 not n7425 ; n7425_not
g26369 not n5274 ; n5274_not
g26370 not n9720 ; n9720_not
g26371 not n5652 ; n5652_not
g26372 not n5256 ; n5256_not
g26373 not n9243 ; n9243_not
g26374 not n9234 ; n9234_not
g26375 not n5265 ; n5265_not
g26376 not n5049 ; n5049_not
g26377 not n5058 ; n5058_not
g26378 not n9432 ; n9432_not
g26379 not n6174 ; n6174_not
g26380 not n9207 ; n9207_not
g26381 not n6165 ; n6165_not
g26382 not n6741 ; n6741_not
g26383 not n6732 ; n6732_not
g26384 not n5625 ; n5625_not
g26385 not n7353 ; n7353_not
g26386 not n6723 ; n6723_not
g26387 not n9306 ; n9306_not
g26388 not n4950 ; n4950_not
g26389 not n6309 ; n6309_not
g26390 not n4752 ; n4752_not
g26391 not n8721 ; n8721_not
g26392 not n3078 ; n3078_not
g26393 not n2394 ; n2394_not
g26394 not n4716 ; n4716_not
g26395 not n2655 ; n2655_not
g26396 not n4680 ; n4680_not
g26397 not n2691 ; n2691_not
g26398 not n8505 ; n8505_not
g26399 not n2457 ; n2457_not
g26400 not n4644 ; n4644_not
g26401 not n2466 ; n2466_not
g26402 not n4608 ; n4608_not
g26403 not n2727 ; n2727_not
g26404 not n2493 ; n2493_not
g26405 not n2763 ; n2763_not
g26406 not n7623 ; n7623_not
g26407 not n7614 ; n7614_not
g26408 not n7551 ; n7551_not
g26409 not n2385 ; n2385_not
g26410 not n3384 ; n3384_not
g26411 not n4860 ; n4860_not
g26412 not n9360 ; n9360_not
g26413 not n2187 ; n2187_not
g26414 not n3357 ; n3357_not
g26415 not n3087 ; n3087_not
g26416 not n4824 ; n4824_not
g26417 not n7803 ; n7803_not
g26418 not n3375 ; n3375_not
g26419 not n2592 ; n2592_not
g26420 not n2583 ; n2583_not
g26421 not n4419 ; n4419_not
g26422 not n4086 ; n4086_not
g26423 not n2952 ; n2952_not
g26424 not n4077 ; n4077_not
g26425 not n4383 ; n4383_not
g26426 not n4347 ; n4347_not
g26427 not n4239 ; n4239_not
g26428 not n4248 ; n4248_not
g26429 not n8136 ; n8136_not
g26430 not n8541 ; n8541_not
g26431 not n2853 ; n2853_not
g26432 not n3096 ; n3096_not
g26433 not n4275 ; n4275_not
g26434 not n8172 ; n8172_not
g26435 not n7731 ; n7731_not
g26436 not n7722 ; n7722_not
g26437 not n4590 ; n4590_not
g26438 not n2529 ; n2529_not
g26439 not n2538 ; n2538_not
g26440 not n8064 ; n8064_not
g26441 not n4527 ; n4527_not
g26442 not n8208 ; n8208_not
g26443 not n4185 ; n4185_not
g26444 not n4194 ; n4194_not
g26445 not n4491 ; n4491_not
g26446 not n8613 ; n8613_not
g26447 not n7650 ; n7650_not
g26448 not n4158 ; n4158_not
g26449 not n4149 ; n4149_not
g26450 not n2880 ; n2880_not
g26451 not n4455 ; n4455_not
g26452 not n2916 ; n2916_not
g26453 not n1656 ; n1656_not
g26454 not n8280 ; n8280_not
g26455 not n1854 ; n1854_not
g26456 not n3294 ; n3294_not
g26457 not n1629 ; n1629_not
g26458 not n4941 ; n4941_not
g26459 not n1818 ; n1818_not
g26460 not n3285 ; n3285_not
g26461 not n3591 ; n3591_not
g26462 not n1593 ; n1593_not
g26463 not n1584 ; n1584_not
g26464 not n1278 ; n1278_not
g26465 not n1782 ; n1782_not
g26466 not n3780 ; n3780_not
g26467 not n3627 ; n3627_not
g26468 not n3636 ; n3636_not
g26469 not n3744 ; n3744_not
g26470 not n3708 ; n3708_not
g26471 not n3690 ; n3690_not
g26472 not n3645 ; n3645_not
g26473 not n1719 ; n1719_not
g26474 not n8451 ; n8451_not
g26475 not n1395 ; n1395_not
g26476 not n8316 ; n8316_not
g26477 not n1368 ; n1368_not
g26478 not n1467 ; n1467_not
g26479 not n7902 ; n7902_not
g26480 not n2268 ; n2268_not
g26481 not n3447 ; n3447_not
g26482 not n2196 ; n2196_not
g26483 not n3177 ; n3177_not
g26484 not n1935 ; n1935_not
g26485 not n8352 ; n8352_not
g26486 not n3186 ; n3186_not
g26487 not n2079 ; n2079_not
g26488 not n7911 ; n7911_not
g26489 not n1971 ; n1971_not
g26490 not n8019 ; n8019_not
g26491 not n3483 ; n3483_not
g26492 not n3852 ; n3852_not
g26493 not n1737 ; n1737_not
g26494 not n1665 ; n1665_not
g26495 not n1089 ; n1089_not
g26496 not n3555 ; n3555_not
g26497 not n1179 ; n1179_not
g26498 not n3672 ; n3672_not
g26499 not n7830 ; n7830_not
g26500 not n3816 ; n3816_not
g26501 not n3924 ; n3924_not
g26502 not n1890 ; n1890_not
g26503 not n8244 ; n8244_not
g26504 not n1908 ; n1908_not
g26505 not n3249 ; n3249_not
g26506 not n3519 ; n3519_not
g26507 not n2917 ; n2917_not
g26508 not n2926 ; n2926_not
g26509 not n3187 ; n3187_not
g26510 not n8353 ; n8353_not
g26511 not n3547 ; n3547_not
g26512 not n2881 ; n2881_not
g26513 not n9280 ; n9280_not
g26514 not n2890 ; n2890_not
g26515 not n6175 ; n6175_not
g26516 not n5806 ; n5806_not
g26517 not n5653 ; n5653_not
g26518 not n5662 ; n5662_not
g26519 not n3448 ; n3448_not
g26520 not n6067 ; n6067_not
g26521 not n3484 ; n3484_not
g26522 not n8470 ; n8470_not
g26523 not n3556 ; n3556_not
g26524 not n3079 ; n3079_not
g26525 not n3295 ; n3295_not
g26526 not n5734 ; n5734_not
g26527 not n5725 ; n5725_not
g26528 not n3259 ; n3259_not
g26529 not n2953 ; n2953_not
g26530 not n3592 ; n3592_not
g26531 not n3628 ; n3628_not
g26532 not n9505 ; n9505_not
g26533 not n2962 ; n2962_not
g26534 not n6139 ; n6139_not
g26535 not n5761 ; n5761_not
g26536 not n5770 ; n5770_not
g26537 not n9721 ; n9721_not
g26538 not n5590 ; n5590_not
g26539 not n5941 ; n5941_not
g26540 not n8803 ; n8803_not
g26541 not n3385 ; n3385_not
g26542 not n8515 ; n8515_not
g26543 not n1747 ; n1747_not
g26544 not n1549 ; n1549_not
g26545 not n1783 ; n1783_not
g26546 not n7057 ; n7057_not
g26547 not n6724 ; n6724_not
g26548 not n8650 ; n8650_not
g26549 not n1819 ; n1819_not
g26550 not n1855 ; n1855_not
g26551 not n9613 ; n9613_not
g26552 not n8902 ; n8902_not
g26553 not n9136 ; n9136_not
g26554 not n9910 ; n9910_not
g26555 not n1891 ; n1891_not
g26556 not n7093 ; n7093_not
g26557 not n6652 ; n6652_not
g26558 not n9541 ; n9541_not
g26559 not n1972 ; n1972_not
g26560 not n9172 ; n9172_not
g26561 not n6616 ; n6616_not
g26562 not n6580 ; n6580_not
g26563 not n9064 ; n9064_not
g26564 not n6913 ; n6913_not
g26565 not n9820 ; n9820_not
g26566 not n8614 ; n8614_not
g26567 not n9811 ; n9811_not
g26568 not n9028 ; n9028_not
g26569 not n8551 ; n8551_not
g26570 not n8542 ; n8542_not
g26571 not n1279 ; n1279_not
g26572 not n6841 ; n6841_not
g26573 not n1369 ; n1369_not
g26574 not n1378 ; n1378_not
g26575 not n8623 ; n8623_not
g26576 not n6805 ; n6805_not
g26577 not n8506 ; n8506_not
g26578 not n6364 ; n6364_not
g26579 not n1396 ; n1396_not
g26580 not n1594 ; n1594_not
g26581 not n1477 ; n1477_not
g26582 not n1468 ; n1468_not
g26583 not n1666 ; n1666_not
g26584 not n6373 ; n6373_not
g26585 not n2827 ; n2827_not
g26586 not n2854 ; n2854_not
g26587 not n2836 ; n2836_not
g26588 not n2863 ; n2863_not
g26589 not n5950 ; n5950_not
g26590 not n6319 ; n6319_not
g26591 not n5914 ; n5914_not
g26592 not n5905 ; n5905_not
g26593 not n6283 ; n6283_not
g26594 not n6247 ; n6247_not
g26595 not n3088 ; n3088_not
g26596 not n2818 ; n2818_not
g26597 not n5842 ; n5842_not
g26598 not n5833 ; n5833_not
g26599 not n9244 ; n9244_not
g26600 not n8731 ; n8731_not
g26601 not n8722 ; n8722_not
g26602 not n6544 ; n6544_not
g26603 not n2359 ; n2359_not
g26604 not n9532 ; n9532_not
g26605 not n2368 ; n2368_not
g26606 not n2395 ; n2395_not
g26607 not n2197 ; n2197_not
g26608 not n2467 ; n2467_not
g26609 not n6508 ; n6508_not
g26610 not n7129 ; n7129_not
g26611 not n2278 ; n2278_not
g26612 not n2269 ; n2269_not
g26613 not n2539 ; n2539_not
g26614 not n6472 ; n6472_not
g26615 not n2386 ; n2386_not
g26616 not n2656 ; n2656_not
g26617 not n9208 ; n9208_not
g26618 not n2692 ; n2692_not
g26619 not n6436 ; n6436_not
g26620 not n2728 ; n2728_not
g26621 not n2764 ; n2764_not
g26622 not n7462 ; n7462_not
g26623 not n7561 ; n7561_not
g26624 not n4915 ; n4915_not
g26625 not n9316 ; n9316_not
g26626 not n4087 ; n4087_not
g26627 not n3781 ; n3781_not
g26628 not n3790 ; n3790_not
g26629 not n7912 ; n7912_not
g26630 not n8245 ; n8245_not
g26631 not n7255 ; n7255_not
g26632 not n3826 ; n3826_not
g26633 not n3817 ; n3817_not
g26634 not n5635 ; n5635_not
g26635 not n4159 ; n4159_not
g26636 not n3853 ; n3853_not
g26637 not n5608 ; n5608_not
g26638 not n7840 ; n7840_not
g26639 not n4618 ; n4618_not
g26640 not n4951 ; n4951_not
g26641 not n7426 ; n7426_not
g26642 not n7435 ; n7435_not
g26643 not n8281 ; n8281_not
g26644 not n7552 ; n7552_not
g26645 not n4924 ; n4924_not
g26646 not n3709 ; n3709_not
g26647 not n3718 ; n3718_not
g26648 not n3754 ; n3754_not
g26649 not n3745 ; n3745_not
g26650 not n7534 ; n7534_not
g26651 not n7246 ; n7246_not
g26652 not n5266 ; n5266_not
g26653 not n7471 ; n7471_not
g26654 not n8137 ; n8137_not
g26655 not n5356 ; n5356_not
g26656 not n4348 ; n4348_not
g26657 not n4384 ; n4384_not
g26658 not n7624 ; n7624_not
g26659 not n9433 ; n9433_not
g26660 not n5536 ; n5536_not
g26661 not n4456 ; n4456_not
g26662 not n5392 ; n5392_not
g26663 not n4492 ; n4492_not
g26664 not n4528 ; n4528_not
g26665 not n8029 ; n8029_not
g26666 not n5428 ; n5428_not
g26667 not n4276 ; n4276_not
g26668 not n4609 ; n4609_not
g26669 not n8065 ; n8065_not
g26670 not n5464 ; n5464_not
g26671 not n5626 ; n5626_not
g26672 not n5284 ; n5284_not
g26673 not n8209 ; n8209_not
g26674 not n4195 ; n4195_not
g26675 not n4249 ; n4249_not
g26676 not n3943 ; n3943_not
g26677 not n7507 ; n7507_not
g26678 not n8173 ; n8173_not
g26679 not n7660 ; n7660_not
g26680 not n4942 ; n4942_not
g26681 not n4294 ; n4294_not
g26682 not n3970 ; n3970_not
g26683 not n7543 ; n7543_not
g26684 not n5572 ; n5572_not
g26685 not n9370 ; n9370_not
g26686 not n5095 ; n5095_not
g26687 not n7804 ; n7804_not
g26688 not n4645 ; n4645_not
g26689 not n4762 ; n4762_not
g26690 not n8911 ; n8911_not
g26691 not n7291 ; n7291_not
g26692 not n4870 ; n4870_not
g26693 not n4861 ; n4861_not
g26694 not n5167 ; n5167_not
g26695 not n7732 ; n7732_not
g26696 not n5059 ; n5059_not
g26697 not n7390 ; n7390_not
g26698 not n7363 ; n7363_not
g26699 not n3952 ; n3952_not
g26700 not n4681 ; n4681_not
g26701 not n4690 ; n4690_not
g26702 not n3961 ; n3961_not
g26703 not n4726 ; n4726_not
g26704 not n7318 ; n7318_not
g26705 not n4753 ; n4753_not
g26706 not n8317 ; n8317_not
g26707 not n7282 ; n7282_not
g26708 not n4654 ; n4654_not
g26709 not n8830 ; n8830_not
g26710 not n4717 ; n4717_not
g26711 not n4834 ; n4834_not
g26712 not n7327 ; n7327_not
g26713 not n4825 ; n4825_not
g26714 not n7354 ; n7354_not
g26715 not n8291 ; n8291_not
g26716 not n5096 ; n5096_not
g26717 not n5168 ; n5168_not
g26718 not n4493 ; n4493_not
g26719 not n9029 ; n9029_not
g26720 not n9650 ; n9650_not
g26721 not n2468 ; n2468_not
g26722 not n4835 ; n4835_not
g26723 not n9821 ; n9821_not
g26724 not n2396 ; n2396_not
g26725 not n7661 ; n7661_not
g26726 not n4529 ; n4529_not
g26727 not n8282 ; n8282_not
g26728 not n4538 ; n4538_not
g26729 not n4871 ; n4871_not
g26730 not n6554 ; n6554_not
g26731 not n6446 ; n6446_not
g26732 not n9551 ; n9551_not
g26733 not n2279 ; n2279_not
g26734 not n6437 ; n6437_not
g26735 not n9542 ; n9542_not
g26736 not n4349 ; n4349_not
g26737 not n6743 ; n6743_not
g26738 not n4358 ; n4358_not
g26739 not n6518 ; n6518_not
g26740 not n4655 ; n4655_not
g26741 not n6509 ; n6509_not
g26742 not n4619 ; n4619_not
g26743 not n9722 ; n9722_not
g26744 not n4592 ; n4592_not
g26745 not n4565 ; n4565_not
g26746 not n9731 ; n9731_not
g26747 not n8219 ; n8219_not
g26748 not n8660 ; n8660_not
g26749 not n9407 ; n9407_not
g26750 not n7157 ; n7157_not
g26751 not n7166 ; n7166_not
g26752 not n4466 ; n4466_not
g26753 not n7625 ; n7625_not
g26754 not n4457 ; n4457_not
g26755 not n8732 ; n8732_not
g26756 not n9209 ; n9209_not
g26757 not n9344 ; n9344_not
g26758 not n4763 ; n4763_not
g26759 not n6482 ; n6482_not
g26760 not n4727 ; n4727_not
g26761 not n8255 ; n8255_not
g26762 not n2369 ; n2369_not
g26763 not n4394 ; n4394_not
g26764 not n4385 ; n4385_not
g26765 not n6473 ; n6473_not
g26766 not n9065 ; n9065_not
g26767 not n4691 ; n4691_not
g26768 not n8246 ; n8246_not
g26769 not n1595 ; n1595_not
g26770 not n1928 ; n1928_not
g26771 not n9812 ; n9812_not
g26772 not n1667 ; n1667_not
g26773 not n1919 ; n1919_not
g26774 not n7913 ; n7913_not
g26775 not n6662 ; n6662_not
g26776 not n6653 ; n6653_not
g26777 not n8426 ; n8426_not
g26778 not n7841 ; n7841_not
g26779 not n8903 ; n8903_not
g26780 not n6761 ; n6761_not
g26781 not n6626 ; n6626_not
g26782 not n9137 ; n9137_not
g26783 not n6752 ; n6752_not
g26784 not n8471 ; n8471_not
g26785 not n9335 ; n9335_not
g26786 not n6347 ; n6347_not
g26787 not n9380 ; n9380_not
g26788 not n4952 ; n4952_not
g26789 not n6617 ; n6617_not
g26790 not n1748 ; n1748_not
g26791 not n8921 ; n8921_not
g26792 not n6338 ; n6338_not
g26793 not n6545 ; n6545_not
g26794 not n1982 ; n1982_not
g26795 not n1973 ; n1973_not
g26796 not n1937 ; n1937_not
g26797 not n9614 ; n9614_not
g26798 not n9623 ; n9623_not
g26799 not n8318 ; n8318_not
g26800 not n8327 ; n8327_not
g26801 not n1856 ; n1856_not
g26802 not n1865 ; n1865_not
g26803 not n1829 ; n1829_not
g26804 not n1784 ; n1784_not
g26805 not n1793 ; n1793_not
g26806 not n8804 ; n8804_not
g26807 not n8363 ; n8363_not
g26808 not n9371 ; n9371_not
g26809 not n8354 ; n8354_not
g26810 not n1757 ; n1757_not
g26811 not n9353 ; n9353_not
g26812 not n4925 ; n4925_not
g26813 not n1289 ; n1289_not
g26814 not n6581 ; n6581_not
g26815 not n6590 ; n6590_not
g26816 not n5285 ; n5285_not
g26817 not n8840 ; n8840_not
g26818 not n8390 ; n8390_not
g26819 not n9173 ; n9173_not
g26820 not n7733 ; n7733_not
g26821 not n1478 ; n1478_not
g26822 not n7805 ; n7805_not
g26823 not n1559 ; n1559_not
g26824 not n4088 ; n4088_not
g26825 not n7544 ; n7544_not
g26826 not n3674 ; n3674_not
g26827 not n8453 ; n8453_not
g26828 not n3980 ; n3980_not
g26829 not n7364 ; n7364_not
g26830 not n6950 ; n6950_not
g26831 not n9920 ; n9920_not
g26832 not n5357 ; n5357_not
g26833 not n5366 ; n5366_not
g26834 not n5735 ; n5735_not
g26835 not n3359 ; n3359_not
g26836 not n9317 ; n9317_not
g26837 not n3656 ; n3656_not
g26838 not n9803 ; n9803_not
g26839 not n3962 ; n3962_not
g26840 not n8444 ; n8444_not
g26841 not n5960 ; n5960_not
g26842 not n5627 ; n5627_not
g26843 not n8516 ; n8516_not
g26844 not n7148 ; n7148_not
g26845 not n9470 ; n9470_not
g26846 not n3296 ; n3296_not
g26847 not n7562 ; n7562_not
g26848 not n8039 ; n8039_not
g26849 not n7553 ; n7553_not
g26850 not n8480 ; n8480_not
g26851 not n7328 ; n7328_not
g26852 not n3386 ; n3386_not
g26853 not n3368 ; n3368_not
g26854 not n6923 ; n6923_not
g26855 not n6068 ; n6068_not
g26856 not n6914 ; n6914_not
g26857 not n5294 ; n5294_not
g26858 not n3395 ; n3395_not
g26859 not n5663 ; n5663_not
g26860 not n3485 ; n3485_not
g26861 not n3791 ; n3791_not
g26862 not n3647 ; n3647_not
g26863 not n3827 ; n3827_not
g26864 not n9434 ; n9434_not
g26865 not n7472 ; n7472_not
g26866 not n7067 ; n7067_not
g26867 not n7058 ; n7058_not
g26868 not n3593 ; n3593_not
g26869 not n5843 ; n5843_not
g26870 not n5465 ; n5465_not
g26871 not n5474 ; n5474_not
g26872 not n3566 ; n3566_not
g26873 not n3557 ; n3557_not
g26874 not n3863 ; n3863_not
g26875 not n7508 ; n7508_not
g26876 not n5429 ; n5429_not
g26877 not n5438 ; n5438_not
g26878 not n5807 ; n5807_not
g26879 not n9443 ; n9443_not
g26880 not n3665 ; n3665_not
g26881 not n5591 ; n5591_not
g26882 not n5951 ; n5951_not
g26883 not n5573 ; n5573_not
g26884 not n9281 ; n9281_not
g26885 not n5393 ; n5393_not
g26886 not n5771 ; n5771_not
g26887 not n7436 ; n7436_not
g26888 not n3719 ; n3719_not
g26889 not n5915 ; n5915_not
g26890 not n5537 ; n5537_not
g26891 not n5546 ; n5546_not
g26892 not n3449 ; n3449_not
g26893 not n3458 ; n3458_not
g26894 not n3755 ; n3755_not
g26895 not n7094 ; n7094_not
g26896 not n3494 ; n3494_not
g26897 not n8147 ; n8147_not
g26898 not n2891 ; n2891_not
g26899 not n2666 ; n2666_not
g26900 not n2657 ; n2657_not
g26901 not n2927 ; n2927_not
g26902 not n2963 ; n2963_not
g26903 not n2693 ; n2693_not
g26904 not n9245 ; n9245_not
g26905 not n9515 ; n9515_not
g26906 not n9506 ; n9506_not
g26907 not n6806 ; n6806_not
g26908 not n2738 ; n2738_not
g26909 not n6284 ; n6284_not
g26910 not n2729 ; n2729_not
g26911 not n6815 ; n6815_not
g26912 not n2765 ; n2765_not
g26913 not n2774 ; n2774_not
g26914 not n8552 ; n8552_not
g26915 not n2819 ; n2819_not
g26916 not n6383 ; n6383_not
g26917 not n2828 ; n2828_not
g26918 not n7175 ; n7175_not
g26919 not n6356 ; n6356_not
g26920 not n6374 ; n6374_not
g26921 not n8183 ; n8183_not
g26922 not n4583 ; n4583_not
g26923 not n8174 ; n8174_not
g26924 not n8624 ; n8624_not
g26925 not n6365 ; n6365_not
g26926 not n2855 ; n2855_not
g26927 not n7607 ; n7607_not
g26928 not n7652 ; n7652_not
g26929 not n6770 ; n6770_not
g26930 not n8138 ; n8138_not
g26931 not n8066 ; n8066_not
g26932 not n6851 ; n6851_not
g26933 not n7292 ; n7292_not
g26934 not n6176 ; n6176_not
g26935 not n8075 ; n8075_not
g26936 not n3188 ; n3188_not
g26937 not n7256 ; n7256_not
g26938 not n3089 ; n3089_not
g26939 not n6248 ; n6248_not
g26940 not n6842 ; n6842_not
g26941 not n4196 ; n4196_not
g26942 not n8364 ; n8364_not
g26943 not n8625 ; n8625_not
g26944 not n9345 ; n9345_not
g26945 not n8184 ; n8184_not
g26946 not n7626 ; n7626_not
g26947 not n6960 ; n6960_not
g26948 not n7635 ; n7635_not
g26949 not n7068 ; n7068_not
g26950 not n9552 ; n9552_not
g26951 not n7473 ; n7473_not
g26952 not n9075 ; n9075_not
g26953 not n7923 ; n7923_not
g26954 not n7293 ; n7293_not
g26955 not n9444 ; n9444_not
g26956 not n7509 ; n7509_not
g26957 not n7329 ; n7329_not
g26958 not n7914 ; n7914_not
g26959 not n9408 ; n9408_not
g26960 not n6924 ; n6924_not
g26961 not n9336 ; n9336_not
g26962 not n8517 ; n8517_not
g26963 not n8661 ; n8661_not
g26964 not n8841 ; n8841_not
g26965 not n7167 ; n7167_not
g26966 not n7770 ; n7770_not
g26967 not n8922 ; n8922_not
g26968 not n7707 ; n7707_not
g26969 not n7257 ; n7257_not
g26970 not n7842 ; n7842_not
g26971 not n8454 ; n8454_not
g26972 not n9318 ; n9318_not
g26973 not n9480 ; n9480_not
g26974 not n9039 ; n9039_not
g26975 not n7365 ; n7365_not
g26976 not n7851 ; n7851_not
g26977 not n8292 ; n8292_not
g26978 not n8256 ; n8256_not
g26979 not n7806 ; n7806_not
g26980 not n8931 ; n8931_not
g26981 not n8481 ; n8481_not
g26982 not n7815 ; n7815_not
g26983 not n7950 ; n7950_not
g26984 not n8328 ; n8328_not
g26985 not n9066 ; n9066_not
g26986 not n7734 ; n7734_not
g26987 not n8076 ; n8076_not
g26988 not n7185 ; n7185_not
g26989 not n8805 ; n8805_not
g26990 not n7743 ; n7743_not
g26991 not n9516 ; n9516_not
g26992 not n8553 ; n8553_not
g26993 not n8733 ; n8733_not
g26994 not n7671 ; n7671_not
g26995 not n7662 ; n7662_not
g26996 not n9372 ; n9372_not
g26997 not n7437 ; n7437_not
g26998 not n8148 ; n8148_not
g26999 not n7545 ; n7545_not
g27000 not n2964 ; n2964_not
g27001 not n4692 ; n4692_not
g27002 not n5295 ; n5295_not
g27003 not n9624 ; n9624_not
g27004 not n1794 ; n1794_not
g27005 not n4962 ; n4962_not
g27006 not n6375 ; n6375_not
g27007 not n4953 ; n4953_not
g27008 not n1596 ; n1596_not
g27009 not n2577 ; n2577_not
g27010 not n2856 ; n2856_not
g27011 not n9813 ; n9813_not
g27012 not n3666 ; n3666_not
g27013 not n1866 ; n1866_not
g27014 not n3567 ; n3567_not
g27015 not n1956 ; n1956_not
g27016 not n6555 ; n6555_not
g27017 not n6519 ; n6519_not
g27018 not n9219 ; n9219_not
g27019 not n6483 ; n6483_not
g27020 not n2397 ; n2397_not
g27021 not n6069 ; n6069_not
g27022 not n6078 ; n6078_not
g27023 not n9822 ; n9822_not
g27024 not n6447 ; n6447_not
g27025 not n1749 ; n1749_not
g27026 not n1758 ; n1758_not
g27027 not n5268 ; n5268_not
g27028 not n5736 ; n5736_not
g27029 not n9138 ; n9138_not
g27030 not n1569 ; n1569_not
g27031 not n9147 ; n9147_not
g27032 not n4728 ; n4728_not
g27033 not n2595 ; n2595_not
g27034 not n5664 ; n5664_not
g27035 not n5178 ; n5178_not
g27036 not n5646 ; n5646_not
g27037 not n1929 ; n1929_not
g27038 not n3297 ; n3297_not
g27039 not n5169 ; n5169_not
g27040 not n9327 ; n9327_not
g27041 not n5547 ; n5547_not
g27042 not n9660 ; n9660_not
g27043 not n3855 ; n3855_not
g27044 not n5592 ; n5592_not
g27045 not n5583 ; n5583_not
g27046 not n2379 ; n2379_not
g27047 not n4935 ; n4935_not
g27048 not n6348 ; n6348_not
g27049 not n9804 ; n9804_not
g27050 not n1947 ; n1947_not
g27051 not n6339 ; n6339_not
g27052 not n4872 ; n4872_not
g27053 not n1677 ; n1677_not
g27054 not n5628 ; n5628_not
g27055 not n5367 ; n5367_not
g27056 not n4656 ; n4656_not
g27057 not n5439 ; n5439_not
g27058 not n5097 ; n5097_not
g27059 not n1668 ; n1668_not
g27060 not n5475 ; n5475_not
g27061 not n4593 ; n4593_not
g27062 not n4278 ; n4278_not
g27063 not n5286 ; n5286_not
g27064 not n9183 ; n9183_not
g27065 not n9174 ; n9174_not
g27066 not n3198 ; n3198_not
g27067 not n4908 ; n4908_not
g27068 not n6816 ; n6816_not
g27069 not n4764 ; n4764_not
g27070 not n4089 ; n4089_not
g27071 not n3189 ; n3189_not
g27072 not n4926 ; n4926_not
g27073 not n3756 ; n3756_not
g27074 not n1389 ; n1389_not
g27075 not n6780 ; n6780_not
g27076 not n9246 ; n9246_not
g27077 not n2874 ; n2874_not
g27078 not n5844 ; n5844_not
g27079 not n2739 ; n2739_not
g27080 not n2469 ; n2469_not
g27081 not n1479 ; n1479_not
g27082 not n3459 ; n3459_not
g27083 not n2829 ; n2829_not
g27084 not n4359 ; n4359_not
g27085 not n3387 ; n3387_not
g27086 not n3792 ; n3792_not
g27087 not n2928 ; n2928_not
g27088 not n3990 ; n3990_not
g27089 not n3828 ; n3828_not
g27090 not n5880 ; n5880_not
g27091 not n4836 ; n4836_not
g27092 not n3864 ; n3864_not
g27093 not n9732 ; n9732_not
g27094 not n4395 ; n4395_not
g27095 not n6852 ; n6852_not
g27096 not n4098 ; n4098_not
g27097 not n5916 ; n5916_not
g27098 not n2775 ; n2775_not
g27099 not n2892 ; n2892_not
g27100 not n6663 ; n6663_not
g27101 not n5772 ; n5772_not
g27102 not n3981 ; n3981_not
g27103 not n6258 ; n6258_not
g27104 not n6249 ; n6249_not
g27105 not n9291 ; n9291_not
g27106 not n6627 ; n6627_not
g27107 not n9921 ; n9921_not
g27108 not n6591 ; n6591_not
g27109 not n4890 ; n4890_not
g27110 not n4197 ; n4197_not
g27111 not n5259 ; n5259_not
g27112 not n6186 ; n6186_not
g27113 not n6177 ; n6177_not
g27114 not n4539 ; n4539_not
g27115 not n3495 ; n3495_not
g27116 not n2478 ; n2478_not
g27117 not n6762 ; n6762_not
g27118 not n9255 ; n9255_not
g27119 not n5952 ; n5952_not
g27120 not n3684 ; n3684_not
g27121 not n2667 ; n2667_not
g27122 not n5808 ; n5808_not
g27123 not n4467 ; n4467_not
g27124 not n9282 ; n9282_not
g27125 not n4269 ; n4269_not
g27126 not n6294 ; n6294_not
g27127 not n6285 ; n6285_not
g27128 not n1983 ; n1983_not
g27129 not n8770 ; n8770_not
g27130 not n9445 ; n9445_not
g27131 not n5269 ; n5269_not
g27132 not n8077 ; n8077_not
g27133 not n4468 ; n4468_not
g27134 not n4396 ; n4396_not
g27135 not n9922 ; n9922_not
g27136 not n2938 ; n2938_not
g27137 not n2929 ; n2929_not
g27138 not n3199 ; n3199_not
g27139 not n2965 ; n2965_not
g27140 not n4882 ; n4882_not
g27141 not n4873 ; n4873_not
g27142 not n2668 ; n2668_not
g27143 not n4837 ; n4837_not
g27144 not n7294 ; n7294_not
g27145 not n4846 ; n4846_not
g27146 not n9346 ; n9346_not
g27147 not n5179 ; n5179_not
g27148 not n7744 ; n7744_not
g27149 not n9409 ; n9409_not
g27150 not n8743 ; n8743_not
g27151 not n7339 ; n7339_not
g27152 not n4765 ; n4765_not
g27153 not n4774 ; n4774_not
g27154 not n4738 ; n4738_not
g27155 not n7780 ; n7780_not
g27156 not n4729 ; n4729_not
g27157 not n4693 ; n4693_not
g27158 not n2776 ; n2776_not
g27159 not n7375 ; n7375_not
g27160 not n7366 ; n7366_not
g27161 not n7852 ; n7852_not
g27162 not n9373 ; n9373_not
g27163 not n7816 ; n7816_not
g27164 not n9391 ; n9391_not
g27165 not n4963 ; n4963_not
g27166 not n4666 ; n4666_not
g27167 not n4657 ; n4657_not
g27168 not n7564 ; n7564_not
g27169 not n4567 ; n4567_not
g27170 not n5584 ; n5584_not
g27171 not n2479 ; n2479_not
g27172 not n7573 ; n7573_not
g27173 not n4594 ; n4594_not
g27174 not n7582 ; n7582_not
g27175 not n5548 ; n5548_not
g27176 not n4576 ; n4576_not
g27177 not n9805 ; n9805_not
g27178 not n5476 ; n5476_not
g27179 not n2893 ; n2893_not
g27180 not n7195 ; n7195_not
g27181 not n5368 ; n5368_not
g27182 not n7591 ; n7591_not
g27183 not n7438 ; n7438_not
g27184 not n7636 ; n7636_not
g27185 not n7447 ; n7447_not
g27186 not n5296 ; n5296_not
g27187 not n7672 ; n7672_not
g27188 not n7258 ; n7258_not
g27189 not n7267 ; n7267_not
g27190 not n8923 ; n8923_not
g27191 not n9337 ; n9337_not
g27192 not n8734 ; n8734_not
g27193 not n7708 ; n7708_not
g27194 not n4891 ; n4891_not
g27195 not n8626 ; n8626_not
g27196 not n6664 ; n6664_not
g27197 not n3964 ; n3964_not
g27198 not n8806 ; n8806_not
g27199 not n6628 ; n6628_not
g27200 not n8482 ; n8482_not
g27201 not n8491 ; n8491_not
g27202 not n6592 ; n6592_not
g27203 not n8932 ; n8932_not
g27204 not n8293 ; n8293_not
g27205 not n6556 ; n6556_not
g27206 not n3991 ; n3991_not
g27207 not n6484 ; n6484_not
g27208 not n1759 ; n1759_not
g27209 not n6448 ; n6448_not
g27210 not n8842 ; n8842_not
g27211 not n9625 ; n9625_not
g27212 not n1795 ; n1795_not
g27213 not n8905 ; n8905_not
g27214 not n6394 ; n6394_not
g27215 not n3685 ; n3685_not
g27216 not n6367 ; n6367_not
g27217 not n8428 ; n8428_not
g27218 not n5971 ; n5971_not
g27219 not n1867 ; n1867_not
g27220 not n2695 ; n2695_not
g27221 not n7186 ; n7186_not
g27222 not n6349 ; n6349_not
g27223 not n8662 ; n8662_not
g27224 not n9661 ; n9661_not
g27225 not n7960 ; n7960_not
g27226 not n6925 ; n6925_not
g27227 not n9292 ; n9292_not
g27228 not n8590 ; n8590_not
g27229 not n9076 ; n9076_not
g27230 not n7519 ; n7519_not
g27231 not n8365 ; n8365_not
g27232 not n6961 ; n6961_not
g27233 not n6853 ; n6853_not
g27234 not n8554 ; n8554_not
g27235 not n8563 ; n8563_not
g27236 not n4558 ; n4558_not
g27237 not n6817 ; n6817_not
g27238 not n9553 ; n9553_not
g27239 not n3937 ; n3937_not
g27240 not n6376 ; n6376_not
g27241 not n6781 ; n6781_not
g27242 not n3955 ; n3955_not
g27243 not n8527 ; n8527_not
g27244 not n8329 ; n8329_not
g27245 not n8518 ; n8518_not
g27246 not n3388 ; n3388_not
g27247 not n8851 ; n8851_not
g27248 not n7924 ; n7924_not
g27249 not n8815 ; n8815_not
g27250 not n1489 ; n1489_not
g27251 not n8635 ; n8635_not
g27252 not n7069 ; n7069_not
g27253 not n1678 ; n1678_not
g27254 not n9148 ; n9148_not
g27255 not n5746 ; n5746_not
g27256 not n5737 ; n5737_not
g27257 not n6079 ; n6079_not
g27258 not n3874 ; n3874_not
g27259 not n1948 ; n1948_not
g27260 not n3865 ; n3865_not
g27261 not n5674 ; n5674_not
g27262 not n5665 ; n5665_not
g27263 not n8437 ; n8437_not
g27264 not n8464 ; n8464_not
g27265 not n8707 ; n8707_not
g27266 not n3568 ; n3568_not
g27267 not n1984 ; n1984_not
g27268 not n3496 ; n3496_not
g27269 not n5980 ; n5980_not
g27270 not n9481 ; n9481_not
g27271 not n8185 ; n8185_not
g27272 not n9733 ; n9733_not
g27273 not n4927 ; n4927_not
g27274 not n5575 ; n5575_not
g27275 not n4288 ; n4288_not
g27276 not n8149 ; n8149_not
g27277 not n3982 ; n3982_not
g27278 not n9931 ; n9931_not
g27279 not n9328 ; n9328_not
g27280 not n9184 ; n9184_not
g27281 not n4099 ; n4099_not
g27282 not n5845 ; n5845_not
g27283 not n7483 ; n7483_not
g27284 not n3766 ; n3766_not
g27285 not n8257 ; n8257_not
g27286 not n6259 ; n6259_not
g27287 not n5881 ; n5881_not
g27288 not n5890 ; n5890_not
g27289 not n3757 ; n3757_not
g27290 not n6295 ; n6295_not
g27291 not n5926 ; n5926_not
g27292 not n5917 ; n5917_not
g27293 not n9256 ; n9256_not
g27294 not n8671 ; n8671_not
g27295 not n3694 ; n3694_not
g27296 not n8419 ; n8419_not
g27297 not n5782 ; n5782_not
g27298 not n5773 ; n5773_not
g27299 not n8455 ; n8455_not
g27300 not n3838 ; n3838_not
g27301 not n9517 ; n9517_not
g27302 not n6187 ; n6187_not
g27303 not n5809 ; n5809_not
g27304 not n3829 ; n3829_not
g27305 not n7474 ; n7474_not
g27306 not n5818 ; n5818_not
g27307 not n3793 ; n3793_not
g27308 not n5854 ; n5854_not
g27309 not n8564 ; n8564_not
g27310 not n2786 ; n2786_not
g27311 not n2939 ; n2939_not
g27312 not n2975 ; n2975_not
g27313 not n2669 ; n2669_not
g27314 not n2678 ; n2678_not
g27315 not n4847 ; n4847_not
g27316 not n4469 ; n4469_not
g27317 not n4289 ; n4289_not
g27318 not n9257 ; n9257_not
g27319 not n8456 ; n8456_not
g27320 not n9446 ; n9446_not
g27321 not n3659 ; n3659_not
g27322 not n3668 ; n3668_not
g27323 not n3686 ; n3686_not
g27324 not n3992 ; n3992_not
g27325 not n8429 ; n8429_not
g27326 not n3695 ; n3695_not
g27327 not n9932 ; n9932_not
g27328 not n3875 ; n3875_not
g27329 not n3578 ; n3578_not
g27330 not n3569 ; n3569_not
g27331 not n3839 ; n3839_not
g27332 not n3767 ; n3767_not
g27333 not n9455 ; n9455_not
g27334 not n3497 ; n3497_not
g27335 not n9293 ; n9293_not
g27336 not n4478 ; n4478_not
g27337 not n2777 ; n2777_not
g27338 not n9491 ; n9491_not
g27339 not n9482 ; n9482_not
g27340 not n4775 ; n4775_not
g27341 not n2858 ; n2858_not
g27342 not n8087 ; n8087_not
g27343 not n8078 ; n8078_not
g27344 not n4739 ; n4739_not
g27345 not n4397 ; n4397_not
g27346 not n4667 ; n4667_not
g27347 not n8528 ; n8528_not
g27348 not n4298 ; n4298_not
g27349 not n4595 ; n4595_not
g27350 not n4568 ; n4568_not
g27351 not n4559 ; n4559_not
g27352 not n8492 ; n8492_not
g27353 not n9329 ; n9329_not
g27354 not n9419 ; n9419_not
g27355 not n3965 ; n3965_not
g27356 not n5990 ; n5990_not
g27357 not n6962 ; n6962_not
g27358 not n6971 ; n6971_not
g27359 not n7376 ; n7376_not
g27360 not n6935 ; n6935_not
g27361 not n6926 ; n6926_not
g27362 not n8852 ; n8852_not
g27363 not n1697 ; n1697_not
g27364 not n6890 ; n6890_not
g27365 not n6188 ; n6188_not
g27366 not n6863 ; n6863_not
g27367 not n6854 ; n6854_not
g27368 not n7268 ; n7268_not
g27369 not n9149 ; n9149_not
g27370 not n6818 ; n6818_not
g27371 not n6827 ; n6827_not
g27372 not n6296 ; n6296_not
g27373 not n7484 ; n7484_not
g27374 not n5855 ; n5855_not
g27375 not n8780 ; n8780_not
g27376 not n8339 ; n8339_not
g27377 not n1877 ; n1877_not
g27378 not n1868 ; n1868_not
g27379 not n5891 ; n5891_not
g27380 not n7448 ; n7448_not
g27381 not n1796 ; n1796_not
g27382 not n5549 ; n5549_not
g27383 not n5558 ; n5558_not
g27384 not n5927 ; n5927_not
g27385 not n8816 ; n8816_not
g27386 not n1769 ; n1769_not
g27387 not n8366 ; n8366_not
g27388 not n8375 ; n8375_not
g27389 not n9185 ; n9185_not
g27390 not n6593 ; n6593_not
g27391 not n9626 ; n9626_not
g27392 not n9635 ; n9635_not
g27393 not n9671 ; n9671_not
g27394 not n9662 ; n9662_not
g27395 not n6566 ; n6566_not
g27396 not n6557 ; n6557_not
g27397 not n9824 ; n9824_not
g27398 not n9707 ; n9707_not
g27399 not n6458 ; n6458_not
g27400 not n9851 ; n9851_not
g27401 not n6449 ; n6449_not
g27402 not n9743 ; n9743_not
g27403 not n9734 ; n9734_not
g27404 not n6485 ; n6485_not
g27405 not n6494 ; n6494_not
g27406 not n9077 ; n9077_not
g27407 not n6782 ; n6782_not
g27408 not n7196 ; n7196_not
g27409 not n7169 ; n7169_not
g27410 not n6737 ; n6737_not
g27411 not n8933 ; n8933_not
g27412 not n9590 ; n9590_not
g27413 not n6665 ; n6665_not
g27414 not n6674 ; n6674_not
g27415 not n6638 ; n6638_not
g27416 not n6629 ; n6629_not
g27417 not n9770 ; n9770_not
g27418 not n6755 ; n6755_not
g27419 not n1679 ; n1679_not
g27420 not n6764 ; n6764_not
g27421 not n8636 ; n8636_not
g27422 not n8195 ; n8195_not
g27423 not n8906 ; n8906_not
g27424 not n8186 ; n8186_not
g27425 not n7817 ; n7817_not
g27426 not n8672 ; n8672_not
g27427 not n7781 ; n7781_not
g27428 not n7745 ; n7745_not
g27429 not n7709 ; n7709_not
g27430 not n5279 ; n5279_not
g27431 not n4928 ; n4928_not
g27432 not n7673 ; n7673_not
g27433 not n8708 ; n8708_not
g27434 not n2579 ; n2579_not
g27435 not n8267 ; n8267_not
g27436 not n7637 ; n7637_not
g27437 not n7187 ; n7187_not
g27438 not n4883 ; n4883_not
g27439 not n7961 ; n7961_not
g27440 not n4892 ; n4892_not
g27441 not n8159 ; n8159_not
g27442 not n2849 ; n2849_not
g27443 not n7925 ; n7925_not
g27444 not n9527 ; n9527_not
g27445 not n9842 ; n9842_not
g27446 not n4946 ; n4946_not
g27447 not n9518 ; n9518_not
g27448 not n4964 ; n4964_not
g27449 not n7853 ; n7853_not
g27450 not n9833 ; n9833_not
g27451 not n1949 ; n1949_not
g27452 not n5675 ; n5675_not
g27453 not n5297 ; n5297_not
g27454 not n9554 ; n9554_not
g27455 not n1994 ; n1994_not
g27456 not n1985 ; n1985_not
g27457 not n5378 ; n5378_not
g27458 not n8294 ; n8294_not
g27459 not n8744 ; n8744_not
g27460 not n5369 ; n5369_not
g27461 not n5747 ; n5747_not
g27462 not n7583 ; n7583_not
g27463 not n5783 ; n5783_not
g27464 not n8258 ; n8258_not
g27465 not n5819 ; n5819_not
g27466 not n9563 ; n9563_not
g27467 not n2588 ; n2588_not
g27468 not n5486 ; n5486_not
g27469 not n5477 ; n5477_not
g27470 not n7079 ; n7079_not
g27471 not n8493 ; n8493_not
g27472 not n8565 ; n8565_not
g27473 not n8637 ; n8637_not
g27474 not n3768 ; n3768_not
g27475 not n7971 ; n7971_not
g27476 not n1995 ; n1995_not
g27477 not n2967 ; n2967_not
g27478 not n2868 ; n2868_not
g27479 not n7962 ; n7962_not
g27480 not n2976 ; n2976_not
g27481 not n8781 ; n8781_not
g27482 not n1698 ; n1698_not
g27483 not n1689 ; n1689_not
g27484 not n8880 ; n8880_not
g27485 not n1878 ; n1878_not
g27486 not n3579 ; n3579_not
g27487 not n8745 ; n8745_not
g27488 not n8853 ; n8853_not
g27489 not n8709 ; n8709_not
g27490 not n1959 ; n1959_not
g27491 not n8907 ; n8907_not
g27492 not n8916 ; n8916_not
g27493 not n2679 ; n2679_not
g27494 not n8529 ; n8529_not
g27495 not n8673 ; n8673_not
g27496 not n8457 ; n8457_not
g27497 not n2787 ; n2787_not
g27498 not n3696 ; n3696_not
g27499 not n8475 ; n8475_not
g27500 not n7980 ; n7980_not
g27501 not n8817 ; n8817_not
g27502 not n7197 ; n7197_not
g27503 not n6765 ; n6765_not
g27504 not n9636 ; n9636_not
g27505 not n9159 ; n9159_not
g27506 not n9348 ; n9348_not
g27507 not n4596 ; n4596_not
g27508 not n9843 ; n9843_not
g27509 not n9528 ; n9528_not
g27510 not n6459 ; n6459_not
g27511 not n6495 ; n6495_not
g27512 not n6567 ; n6567_not
g27513 not n9366 ; n9366_not
g27514 not n4884 ; n4884_not
g27515 not n9357 ; n9357_not
g27516 not n6198 ; n6198_not
g27517 not n4848 ; n4848_not
g27518 not n6189 ; n6189_not
g27519 not n6639 ; n6639_not
g27520 not n9861 ; n9861_not
g27521 not n9375 ; n9375_not
g27522 not n4776 ; n4776_not
g27523 not n8871 ; n8871_not
g27524 not n4668 ; n4668_not
g27525 not n6675 ; n6675_not
g27526 not n9708 ; n9708_not
g27527 not n9456 ; n9456_not
g27528 not n8970 ; n8970_not
g27529 not n7449 ; n7449_not
g27530 not n5928 ; n5928_not
g27531 not n5892 ; n5892_not
g27532 not n9672 ; n9672_not
g27533 not n7377 ; n7377_not
g27534 not n9258 ; n9258_not
g27535 not n9267 ; n9267_not
g27536 not n7485 ; n7485_not
g27537 not n9744 ; n9744_not
g27538 not n5856 ; n5856_not
g27539 not n9195 ; n9195_not
g27540 not n5784 ; n5784_not
g27541 not n9492 ; n9492_not
g27542 not n5748 ; n5748_not
g27543 not n9294 ; n9294_not
g27544 not n5676 ; n5676_not
g27545 not n9780 ; n9780_not
g27546 not n9186 ; n9186_not
g27547 not n5559 ; n5559_not
g27548 not n8934 ; n8934_not
g27549 not n8943 ; n8943_not
g27550 not n5487 ; n5487_not
g27551 not n5379 ; n5379_not
g27552 not n4974 ; n4974_not
g27553 not n4965 ; n4965_not
g27554 not n7269 ; n7269_not
g27555 not n7746 ; n7746_not
g27556 not n7755 ; n7755_not
g27557 not n8196 ; n8196_not
g27558 not n6378 ; n6378_not
g27559 not n6792 ; n6792_not
g27560 not n7791 ; n7791_not
g27561 not n7782 ; n7782_not
g27562 not n6972 ; n6972_not
g27563 not n6828 ; n6828_not
g27564 not n9087 ; n9087_not
g27565 not n7818 ; n7818_not
g27566 not n7827 ; n7827_not
g27567 not n6936 ; n6936_not
g27568 not n8268 ; n8268_not
g27569 not n3669 ; n3669_not
g27570 not n3975 ; n3975_not
g27571 not n7863 ; n7863_not
g27572 not n7854 ; n7854_not
g27573 not n3939 ; n3939_not
g27574 not n3948 ; n3948_not
g27575 not n3966 ; n3966_not
g27576 not n6864 ; n6864_not
g27577 not n9933 ; n9933_not
g27578 not n7890 ; n7890_not
g27579 not n3876 ; n3876_not
g27580 not n7935 ; n7935_not
g27581 not n7926 ; n7926_not
g27582 not n8376 ; n8376_not
g27583 not n9564 ; n9564_not
g27584 not n9078 ; n9078_not
g27585 not n7719 ; n7719_not
g27586 not n7674 ; n7674_not
g27587 not n7683 ; n7683_not
g27588 not n4479 ; n4479_not
g27589 not n8088 ; n8088_not
g27590 not n7638 ; n7638_not
g27591 not n7647 ; n7647_not
g27592 not n4299 ; n4299_not
g27593 not n3993 ; n3993_not
g27594 not n4569 ; n4569_not
g27595 not n6297 ; n6297_not
g27596 not n9907 ; n9907_not
g27597 not n8647 ; n8647_not
g27598 not n5677 ; n5677_not
g27599 not n8872 ; n8872_not
g27600 not n5686 ; n5686_not
g27601 not n5992 ; n5992_not
g27602 not n6865 ; n6865_not
g27603 not n8854 ; n8854_not
g27604 not n8638 ; n8638_not
g27605 not n8944 ; n8944_not
g27606 not n5965 ; n5965_not
g27607 not n1699 ; n1699_not
g27608 not n6739 ; n6739_not
g27609 not n9088 ; n9088_not
g27610 not n8980 ; n8980_not
g27611 not n6748 ; n6748_not
g27612 not n6766 ; n6766_not
g27613 not n6937 ; n6937_not
g27614 not n6676 ; n6676_not
g27615 not n9493 ; n9493_not
g27616 not n9709 ; n9709_not
g27617 not n5983 ; n5983_not
g27618 not n8494 ; n8494_not
g27619 not n6784 ; n6784_not
g27620 not n5938 ; n5938_not
g27621 not n6775 ; n6775_not
g27622 not n1879 ; n1879_not
g27623 not n8908 ; n8908_not
g27624 not n6829 ; n6829_not
g27625 not n6568 ; n6568_not
g27626 not n8539 ; n8539_not
g27627 not n9637 ; n9637_not
g27628 not n6496 ; n6496_not
g27629 not n9529 ; n9529_not
g27630 not n6793 ; n6793_not
g27631 not n6388 ; n6388_not
g27632 not n9565 ; n9565_not
g27633 not n9673 ; n9673_not
g27634 not n8566 ; n8566_not
g27635 not n8881 ; n8881_not
g27636 not n5758 ; n5758_not
g27637 not n9871 ; n9871_not
g27638 not n8674 ; n8674_not
g27639 not n6973 ; n6973_not
g27640 not n5749 ; n5749_not
g27641 not n5785 ; n5785_not
g27642 not n5794 ; n5794_not
g27643 not n6199 ; n6199_not
g27644 not n8683 ; n8683_not
g27645 not n5857 ; n5857_not
g27646 not n5866 ; n5866_not
g27647 not n5893 ; n5893_not
g27648 not n5929 ; n5929_not
g27649 not n8089 ; n8089_not
g27650 not n2878 ; n2878_not
g27651 not n7558 ; n7558_not
g27652 not n7990 ; n7990_not
g27653 not n7981 ; n7981_not
g27654 not n7972 ; n7972_not
g27655 not n9367 ; n9367_not
g27656 not n7936 ; n7936_not
g27657 not n9943 ; n9943_not
g27658 not n9862 ; n9862_not
g27659 not n2869 ; n2869_not
g27660 not n7486 ; n7486_not
g27661 not n7495 ; n7495_not
g27662 not n7459 ; n7459_not
g27663 not n7864 ; n7864_not
g27664 not n4975 ; n4975_not
g27665 not n7828 ; n7828_not
g27666 not n8827 ; n8827_not
g27667 not n8818 ; n8818_not
g27668 not n8377 ; n8377_not
g27669 not n3967 ; n3967_not
g27670 not n9268 ; n9268_not
g27671 not n3679 ; n3679_not
g27672 not n8269 ; n8269_not
g27673 not n3697 ; n3697_not
g27674 not n8791 ; n8791_not
g27675 not n3778 ; n3778_not
g27676 not n8782 ; n8782_not
g27677 not n3769 ; n3769_not
g27678 not n8863 ; n8863_not
g27679 not n3877 ; n3877_not
g27680 not n3886 ; n3886_not
g27681 not n8197 ; n8197_not
g27682 not n2977 ; n2977_not
g27683 not n2986 ; n2986_not
g27684 not n7576 ; n7576_not
g27685 not n9970 ; n9970_not
g27686 not n9196 ; n9196_not
g27687 not n7585 ; n7585_not
g27688 not n5488 ; n5488_not
g27689 not n9781 ; n9781_not
g27690 not n7198 ; n7198_not
g27691 not n7648 ; n7648_not
g27692 not n7684 ; n7684_not
g27693 not n7279 ; n7279_not
g27694 not n4849 ; n4849_not
g27695 not n1897 ; n1897_not
g27696 not n8719 ; n8719_not
g27697 not n9745 ; n9745_not
g27698 not n7387 ; n7387_not
g27699 not n8746 ; n8746_not
g27700 not n9934 ; n9934_not
g27701 not n8755 ; n8755_not
g27702 not n7378 ; n7378_not
g27703 not n2788 ; n2788_not
g27704 not n4678 ; n4678_not
g27705 not n1996 ; n1996_not
g27706 not n4669 ; n4669_not
g27707 not n7792 ; n7792_not
g27708 not n9385 ; n9385_not
g27709 not n4777 ; n4777_not
g27710 not n9457 ; n9457_not
g27711 not n7756 ; n7756_not
g27712 not n4786 ; n4786_not
g27713 not n9197 ; n9197_not
g27714 not n9269 ; n9269_not
g27715 not n9755 ; n9755_not
g27716 not n9863 ; n9863_not
g27717 not n9089 ; n9089_not
g27718 not n9719 ; n9719_not
g27719 not n9746 ; n9746_not
g27720 not n9683 ; n9683_not
g27721 not n9386 ; n9386_not
g27722 not n9818 ; n9818_not
g27723 not n9845 ; n9845_not
g27724 not n8909 ; n8909_not
g27725 not n9494 ; n9494_not
g27726 not n9836 ; n9836_not
g27727 not n9980 ; n9980_not
g27728 not n9872 ; n9872_not
g27729 not n9395 ; n9395_not
g27730 not n9467 ; n9467_not
g27731 not n9458 ; n9458_not
g27732 not n9944 ; n9944_not
g27733 not n9908 ; n9908_not
g27734 not n9566 ; n9566_not
g27735 not n9575 ; n9575_not
g27736 not n9647 ; n9647_not
g27737 not n9638 ; n9638_not
g27738 not n9674 ; n9674_not
g27739 not n7586 ; n7586_not
g27740 not n6839 ; n6839_not
g27741 not n6794 ; n6794_not
g27742 not n6686 ; n6686_not
g27743 not n6677 ; n6677_not
g27744 not n6569 ; n6569_not
g27745 not n6578 ; n6578_not
g27746 not n6497 ; n6497_not
g27747 not n3779 ; n3779_not
g27748 not n6398 ; n6398_not
g27749 not n6767 ; n6767_not
g27750 not n5993 ; n5993_not
g27751 not n6389 ; n6389_not
g27752 not n1898 ; n1898_not
g27753 not n8099 ; n8099_not
g27754 not n8576 ; n8576_not
g27755 not n3887 ; n3887_not
g27756 not n5597 ; n5597_not
g27757 not n3986 ; n3986_not
g27758 not n8648 ; n8648_not
g27759 not n8198 ; n8198_not
g27760 not n5939 ; n5939_not
g27761 not n7757 ; n7757_not
g27762 not n7685 ; n7685_not
g27763 not n7649 ; n7649_not
g27764 not n7793 ; n7793_not
g27765 not n7829 ; n7829_not
g27766 not n7865 ; n7865_not
g27767 not n7496 ; n7496_not
g27768 not n2789 ; n2789_not
g27769 not n7937 ; n7937_not
g27770 not n2798 ; n2798_not
g27771 not n7973 ; n7973_not
g27772 not n2987 ; n2987_not
g27773 not n6983 ; n6983_not
g27774 not n6974 ; n6974_not
g27775 not n7388 ; n7388_not
g27776 not n2879 ; n2879_not
g27777 not n1997 ; n1997_not
g27778 not n1889 ; n1889_not
g27779 not n6938 ; n6938_not
g27780 not n6947 ; n6947_not
g27781 not n6866 ; n6866_not
g27782 not n6875 ; n6875_not
g27783 not n8387 ; n8387_not
g27784 not n8378 ; n8378_not
g27785 not n5759 ; n5759_not
g27786 not n5687 ; n5687_not
g27787 not n8864 ; n8864_not
g27788 not n8873 ; n8873_not
g27789 not n8882 ; n8882_not
g27790 not n3968 ; n3968_not
g27791 not n4976 ; n4976_not
g27792 not n8927 ; n8927_not
g27793 not n8459 ; n8459_not
g27794 not n8945 ; n8945_not
g27795 not n4598 ; n4598_not
g27796 not n9791 ; n9791_not
g27797 not n9782 ; n9782_not
g27798 not n4859 ; n4859_not
g27799 not n8981 ; n8981_not
g27800 not n4787 ; n4787_not
g27801 not n4679 ; n4679_not
g27802 not n4589 ; n4589_not
g27803 not n8756 ; n8756_not
g27804 not n5498 ; n5498_not
g27805 not n8279 ; n8279_not
g27806 not n8792 ; n8792_not
g27807 not n8828 ; n8828_not
g27808 not n5489 ; n5489_not
g27809 not n5795 ; n5795_not
g27810 not n5867 ; n5867_not
g27811 not n8684 ; n8684_not
g27812 not n9684 ; n9684_not
g27813 not n9279 ; n9279_not
g27814 not n9468 ; n9468_not
g27815 not n9198 ; n9198_not
g27816 not n8982 ; n8982_not
g27817 not n5868 ; n5868_not
g27818 not n8991 ; n8991_not
g27819 not n5994 ; n5994_not
g27820 not n9981 ; n9981_not
g27821 not n7497 ; n7497_not
g27822 not n5967 ; n5967_not
g27823 not n8955 ; n8955_not
g27824 not n8946 ; n8946_not
g27825 not n9873 ; n9873_not
g27826 not n7587 ; n7587_not
g27827 not n4788 ; n4788_not
g27828 not n7569 ; n7569_not
g27829 not n7596 ; n7596_not
g27830 not n9387 ; n9387_not
g27831 not n6579 ; n6579_not
g27832 not n6687 ; n6687_not
g27833 not n9945 ; n9945_not
g27834 not n6399 ; n6399_not
g27835 not n5796 ; n5796_not
g27836 not n6876 ; n6876_not
g27837 not n3888 ; n3888_not
g27838 not n9576 ; n9576_not
g27839 not n9099 ; n9099_not
g27840 not n6948 ; n6948_not
g27841 not n9756 ; n9756_not
g27842 not n5688 ; n5688_not
g27843 not n6984 ; n6984_not
g27844 not n6768 ; n6768_not
g27845 not n5958 ; n5958_not
g27846 not n9648 ; n9648_not
g27847 not n9792 ; n9792_not
g27848 not n5499 ; n5499_not
g27849 not n4977 ; n4977_not
g27850 not n4986 ; n4986_not
g27851 not n9909 ; n9909_not
g27852 not n5976 ; n5976_not
g27853 not n7389 ; n7389_not
g27854 not n2799 ; n2799_not
g27855 not n7992 ; n7992_not
g27856 not n1899 ; n1899_not
g27857 not n8865 ; n8865_not
g27858 not n7695 ; n7695_not
g27859 not n7686 ; n7686_not
g27860 not n8829 ; n8829_not
g27861 not n8793 ; n8793_not
g27862 not n8757 ; n8757_not
g27863 not n8685 ; n8685_not
g27864 not n7767 ; n7767_not
g27865 not n7758 ; n7758_not
g27866 not n7794 ; n7794_not
g27867 not n8649 ; n8649_not
g27868 not n7839 ; n7839_not
g27869 not n7866 ; n7866_not
g27870 not n7875 ; n7875_not
g27871 not n8577 ; n8577_not
g27872 not n8469 ; n8469_not
g27873 not n7938 ; n7938_not
g27874 not n7947 ; n7947_not
g27875 not n8388 ; n8388_not
g27876 not n9846 ; n9846_not
g27877 not n2988 ; n2988_not
g27878 not n9369 ; n9369_not
g27879 not n9396 ; n9396_not
g27880 not n8568 ; n8568_not
g27881 not n8956 ; n8956_not
g27882 not n8758 ; n8758_not
g27883 not n5599 ; n5599_not
g27884 not n8767 ; n8767_not
g27885 not n5995 ; n5995_not
g27886 not n9856 ; n9856_not
g27887 not n4897 ; n4897_not
g27888 not n8992 ; n8992_not
g27889 not n9685 ; n9685_not
g27890 not n5689 ; n5689_not
g27891 not n5698 ; n5698_not
g27892 not n5797 ; n5797_not
g27893 not n5878 ; n5878_not
g27894 not n5869 ; n5869_not
g27895 not n5959 ; n5959_not
g27896 not n8587 ; n8587_not
g27897 not n8578 ; n8578_not
g27898 not n8794 ; n8794_not
g27899 not n9649 ; n9649_not
g27900 not n9991 ; n9991_not
g27901 not n9982 ; n9982_not
g27902 not n9883 ; n9883_not
g27903 not n9874 ; n9874_not
g27904 not n3889 ; n3889_not
g27905 not n8893 ; n8893_not
g27906 not n9793 ; n9793_not
g27907 not n8686 ; n8686_not
g27908 not n8695 ; n8695_not
g27909 not n8884 ; n8884_not
g27910 not n3898 ; n3898_not
g27911 not n4789 ; n4789_not
g27912 not n9955 ; n9955_not
g27913 not n4798 ; n4798_not
g27914 not n9757 ; n9757_not
g27915 not n4987 ; n4987_not
g27916 not n8659 ; n8659_not
g27917 not n8479 ; n8479_not
g27918 not n5968 ; n5968_not
g27919 not n9847 ; n9847_not
g27920 not n9829 ; n9829_not
g27921 not n7399 ; n7399_not
g27922 not n2998 ; n2998_not
g27923 not n2989 ; n2989_not
g27924 not n7498 ; n7498_not
g27925 not n9577 ; n9577_not
g27926 not n8839 ; n8839_not
g27927 not n7588 ; n7588_not
g27928 not n9397 ; n9397_not
g27929 not n7768 ; n7768_not
g27930 not n6877 ; n6877_not
g27931 not n9946 ; n9946_not
g27932 not n7948 ; n7948_not
g27933 not n6949 ; n6949_not
g27934 not n8389 ; n8389_not
g27935 not n7876 ; n7876_not
g27936 not n6688 ; n6688_not
g27937 not n9469 ; n9469_not
g27938 not n7696 ; n7696_not
g27939 not n9919 ; n9919_not
g27940 not n6985 ; n6985_not
g27941 not n9659 ; n9659_not
g27942 not n6959 ; n6959_not
g27943 not n6887 ; n6887_not
g27944 not n6878 ; n6878_not
g27945 not n5699 ; n5699_not
g27946 not n8399 ; n8399_not
g27947 not n9848 ; n9848_not
g27948 not n7589 ; n7589_not
g27949 not n9758 ; n9758_not
g27950 not n2999 ; n2999_not
g27951 not n9992 ; n9992_not
g27952 not n9794 ; n9794_not
g27953 not n4988 ; n4988_not
g27954 not a[2] ; a[2]_not
g27955 not n9695 ; n9695_not
g27956 not n9398 ; n9398_not
g27957 not n9686 ; n9686_not
g27958 not n6986 ; n6986_not
g27959 not n6995 ; n6995_not
g27960 not n7949 ; n7949_not
g27961 not n9884 ; n9884_not
g27962 not n9578 ; n9578_not
g27963 not n5996 ; n5996_not
g27964 not n9587 ; n9587_not
g27965 not n7697 ; n7697_not
g27966 not n9767 ; n9767_not
g27967 not n7769 ; n7769_not
g27968 not n8993 ; n8993_not
g27969 not n4799 ; n4799_not
g27970 not n3899 ; n3899_not
g27971 not n8588 ; n8588_not
g27972 not n7877 ; n7877_not
g27973 not n9479 ; n9479_not
g27974 not n9956 ; n9956_not
g27975 not n8768 ; n8768_not
g27976 not n6689 ; n6689_not
g27977 not n6698 ; n6698_not
g27978 not n8696 ; n8696_not
g27979 not n5879 ; n5879_not
g27980 not n8957 ; n8957_not
g27981 not n5969 ; n5969_not
g27982 not n9867 ; n9867_not
g27983 not n9993 ; n9993_not
g27984 not n9849 ; n9849_not
g27985 not n8958 ; n8958_not
g27986 not n4899 ; n4899_not
g27987 not n9885 ; n9885_not
g27988 not n8967 ; n8967_not
g27989 not n7986 ; n7986_not
g27990 not n7959 ; n7959_not
g27991 not n6699 ; n6699_not
g27992 not n6789 ; n6789_not
g27993 not n9588 ; n9588_not
g27994 not n7878 ; n7878_not
g27995 not n7887 ; n7887_not
g27996 not n8589 ; n8589_not
g27997 not n9957 ; n9957_not
g27998 not n9696 ; n9696_not
g27999 not n6888 ; n6888_not
g28000 not n7779 ; n7779_not
g28001 not n6996 ; n6996_not
g28002 not n7698 ; n7698_not
g28003 not n8697 ; n8697_not
g28004 not n8769 ; n8769_not
g28005 not n9768 ; n9768_not
g28006 not n8994 ; n8994_not
g28007 not n4998 ; n4998_not
g28008 not n4989 ; n4989_not
g28009 not n9886 ; n9886_not
g28010 not n9895 ; n9895_not
g28011 not a[4] ; a[4]_not
g28012 not n8878 ; n8878_not
g28013 not n7888 ; n7888_not
g28014 not n9967 ; n9967_not
g28015 not n8779 ; n8779_not
g28016 not n8698 ; n8698_not
g28017 not n6997 ; n6997_not
g28018 not n6889 ; n6889_not
g28019 not n9958 ; n9958_not
g28020 not n9589 ; n9589_not
g28021 not n8896 ; n8896_not
g28022 not n5998 ; n5998_not
g28023 not n8599 ; n8599_not
g28024 not n4999 ; n4999_not
g28025 not n8968 ; n8968_not
g28026 not n9994 ; n9994_not
g28027 not n9697 ; n9697_not
g28028 not n5989 ; n5989_not
g28029 not n9769 ; n9769_not
g28030 not n7997 ; n7997_not
g28031 not n7988 ; n7988_not
g28032 not n9698 ; n9698_not
g28033 not n9896 ; n9896_not
g28034 not n7889 ; n7889_not
g28035 not n7979 ; n7979_not
g28036 not n6998 ; n6998_not
g28037 not n9599 ; n9599_not
g28038 not n9968 ; n9968_not
g28039 not n6899 ; n6899_not
g28040 not n9779 ; n9779_not
g28041 not n8969 ; n8969_not
g28042 not n7899 ; n7899_not
g28043 not a[6] ; a[6]_not
g28044 not n8889 ; n8889_not
g28045 not n9969 ; n9969_not
g28046 not n9897 ; n9897_not
g28047 not n8979 ; n8979_not
g28048 not n7989 ; n7989_not
g28049 not n9898 ; n9898_not
g28050 not n9979 ; n9979_not
g28051 not a[8] ; a[8]_not
g28052 not n10100 ; n10100_not
g28053 not n10101 ; n10101_not
g28054 not n11100 ; n11100_not
g28055 not n20100 ; n20100_not
g28056 not n21010 ; n21010_not
g28057 not n12100 ; n12100_not
g28058 not n10300 ; n10300_not
g28059 not n20101 ; n20101_not
g28060 not n10210 ; n10210_not
g28061 not n10003 ; n10003_not
g28062 not n11101 ; n11101_not
g28063 not n10030 ; n10030_not
g28064 not n10111 ; n10111_not
g28065 not n10102 ; n10102_not
g28066 not n20003 ; n20003_not
g28067 not n10301 ; n10301_not
g28068 not n10220 ; n10220_not
g28069 not n13100 ; n13100_not
g28070 not n20102 ; n20102_not
g28071 not n20210 ; n20210_not
g28072 not n20030 ; n20030_not
g28073 not n11210 ; n11210_not
g28074 not n12101 ; n12101_not
g28075 not n10310 ; n10310_not
g28076 not n23000 ; n23000_not
g28077 not n11030 ; n11030_not
g28078 not n11111 ; n11111_not
g28079 not n20111 ; n20111_not
g28080 not n21020 ; n21020_not
g28081 not n11102 ; n11102_not
g28082 not n10040 ; n10040_not
g28083 not n10004 ; n10004_not
g28084 not n22100 ; n22100_not
g28085 not n10112 ; n10112_not
g28086 not n11003 ; n11003_not
g28087 not n21200 ; n21200_not
g28088 not n12102 ; n12102_not
g28089 not n13101 ; n13101_not
g28090 not n10221 ; n10221_not
g28091 not n23001 ; n23001_not
g28092 not n10041 ; n10041_not
g28093 not n11040 ; n11040_not
g28094 not n10032 ; n10032_not
g28095 not n20004 ; n20004_not
g28096 not n21021 ; n21021_not
g28097 not n10410 ; n10410_not
g28098 not n12030 ; n12030_not
g28099 not n22101 ; n22101_not
g28100 not n12210 ; n12210_not
g28101 not n10113 ; n10113_not
g28102 not n21201 ; n21201_not
g28103 not n11112 ; n11112_not
g28104 not n20220 ; n20220_not
g28105 not n14010 ; n14010_not
g28106 not n20400 ; n20400_not
g28107 not n10005 ; n10005_not
g28108 not n12003 ; n12003_not
g28109 not n11004 ; n11004_not
g28110 not n20112 ; n20112_not
g28111 not n12111 ; n12111_not
g28112 not n20040 ; n20040_not
g28113 not n11220 ; n11220_not
g28114 not n11113 ; n11113_not
g28115 not n10321 ; n10321_not
g28116 not n10330 ; n10330_not
g28117 not n10312 ; n10312_not
g28118 not n21310 ; n21310_not
g28119 not n13210 ; n13210_not
g28120 not n11311 ; n11311_not
g28121 not n23002 ; n23002_not
g28122 not n11320 ; n11320_not
g28123 not n10231 ; n10231_not
g28124 not n10222 ; n10222_not
g28125 not n20041 ; n20041_not
g28126 not n20221 ; n20221_not
g28127 not n10150 ; n10150_not
g28128 not n10114 ; n10114_not
g28129 not n10123 ; n10123_not
g28130 not n10600 ; n10600_not
g28131 not n11005 ; n11005_not
g28132 not n10042 ; n10042_not
g28133 not n10051 ; n10051_not
g28134 not n11041 ; n11041_not
g28135 not n10015 ; n10015_not
g28136 not n10006 ; n10006_not
g28137 not n15010 ; n15010_not
g28138 not n13003 ; n13003_not
g28139 not n13030 ; n13030_not
g28140 not n21202 ; n21202_not
g28141 not n10420 ; n10420_not
g28142 not n13111 ; n13111_not
g28143 not n13102 ; n13102_not
g28144 not n20401 ; n20401_not
g28145 not n12040 ; n12040_not
g28146 not n21103 ; n21103_not
g28147 not n23110 ; n23110_not
g28148 not n21022 ; n21022_not
g28149 not n21031 ; n21031_not
g28150 not n11221 ; n11221_not
g28151 not n12112 ; n12112_not
g28152 not n22030 ; n22030_not
g28153 not n22102 ; n22102_not
g28154 not n12004 ; n12004_not
g28155 not n20113 ; n20113_not
g28156 not n12220 ; n12220_not
g28157 not n22210 ; n22210_not
g28158 not n14101 ; n14101_not
g28159 not n14020 ; n14020_not
g28160 not n11410 ; n11410_not
g28161 not n20005 ; n20005_not
g28162 not n23111 ; n23111_not
g28163 not n15020 ; n15020_not
g28164 not n23120 ; n23120_not
g28165 not n22004 ; n22004_not
g28166 not n11600 ; n11600_not
g28167 not n11231 ; n11231_not
g28168 not n20123 ; n20123_not
g28169 not n20042 ; n20042_not
g28170 not n20303 ; n20303_not
g28171 not n22400 ; n22400_not
g28172 not n12221 ; n12221_not
g28173 not n11312 ; n11312_not
g28174 not n13400 ; n13400_not
g28175 not n15200 ; n15200_not
g28176 not n11150 ; n11150_not
g28177 not n11303 ; n11303_not
g28178 not n11006 ; n11006_not
g28179 not n21500 ; n21500_not
g28180 not n14111 ; n14111_not
g28181 not n20402 ; n20402_not
g28182 not n20411 ; n20411_not
g28183 not n11420 ; n11420_not
g28184 not n20600 ; n20600_not
g28185 not n22040 ; n22040_not
g28186 not n22031 ; n22031_not
g28187 not n20150 ; n20150_not
g28188 not n22220 ; n22220_not
g28189 not n21104 ; n21104_not
g28190 not n10331 ; n10331_not
g28191 not n13220 ; n13220_not
g28192 not n21320 ; n21320_not
g28193 not n21311 ; n21311_not
g28194 not n22211 ; n22211_not
g28195 not n11321 ; n11321_not
g28196 not n10601 ; n10601_not
g28197 not n11015 ; n11015_not
g28198 not n20114 ; n20114_not
g28199 not n16010 ; n16010_not
g28200 not n13112 ; n13112_not
g28201 not n10124 ; n10124_not
g28202 not n14102 ; n14102_not
g28203 not n11123 ; n11123_not
g28204 not n22112 ; n22112_not
g28205 not n12005 ; n12005_not
g28206 not n12041 ; n12041_not
g28207 not n10160 ; n10160_not
g28208 not n11051 ; n11051_not
g28209 not n23003 ; n23003_not
g28210 not n21032 ; n21032_not
g28211 not n11222 ; n11222_not
g28212 not n14021 ; n14021_not
g28213 not n20330 ; n20330_not
g28214 not n14210 ; n14210_not
g28215 not n24020 ; n24020_not
g28216 not n23012 ; n23012_not
g28217 not n10232 ; n10232_not
g28218 not n13040 ; n13040_not
g28219 not n17000 ; n17000_not
g28220 not n22103 ; n22103_not
g28221 not n20222 ; n20222_not
g28222 not n10016 ; n10016_not
g28223 not n10052 ; n10052_not
g28224 not n11114 ; n11114_not
g28225 not n12113 ; n12113_not
g28226 not n11042 ; n11042_not
g28227 not n20015 ; n20015_not
g28228 not n20231 ; n20231_not
g28229 not n10421 ; n10421_not
g28230 not n20006 ; n20006_not
g28231 not n21203 ; n21203_not
g28232 not n13004 ; n13004_not
g28233 not n21212 ; n21212_not
g28234 not n20051 ; n20051_not
g28235 not n12051 ; n12051_not
g28236 not n12600 ; n12600_not
g28237 not n14103 ; n14103_not
g28238 not n10431 ; n10431_not
g28239 not n10710 ; n10710_not
g28240 not n20124 ; n20124_not
g28241 not n20601 ; n20601_not
g28242 not n12042 ; n12042_not
g28243 not n12222 ; n12222_not
g28244 not n17100 ; n17100_not
g28245 not n23013 ; n23013_not
g28246 not n10800 ; n10800_not
g28247 not n13113 ; n13113_not
g28248 not n20016 ; n20016_not
g28249 not n12330 ; n12330_not
g28250 not n10611 ; n10611_not
g28251 not n12150 ; n12150_not
g28252 not n20412 ; n20412_not
g28253 not n12114 ; n12114_not
g28254 not n21105 ; n21105_not
g28255 not n11232 ; n11232_not
g28256 not n21321 ; n21321_not
g28257 not n10602 ; n10602_not
g28258 not n20232 ; n20232_not
g28259 not n12123 ; n12123_not
g28260 not n13221 ; n13221_not
g28261 not n12231 ; n12231_not
g28262 not n10422 ; n10422_not
g28263 not n22113 ; n22113_not
g28264 not n14400 ; n14400_not
g28265 not n15201 ; n15201_not
g28266 not n11304 ; n11304_not
g28267 not n10530 ; n10530_not
g28268 not n24021 ; n24021_not
g28269 not n14220 ; n14220_not
g28270 not n11052 ; n11052_not
g28271 not n10017 ; n10017_not
g28272 not n22221 ; n22221_not
g28273 not n12402 ; n12402_not
g28274 not n10053 ; n10053_not
g28275 not n21501 ; n21501_not
g28276 not n14112 ; n14112_not
g28277 not n11160 ; n11160_not
g28278 not n10125 ; n10125_not
g28279 not n21213 ; n21213_not
g28280 not n20160 ; n20160_not
g28281 not n10161 ; n10161_not
g28282 not n21033 ; n21033_not
g28283 not n20304 ; n20304_not
g28284 not n20340 ; n20340_not
g28285 not n13005 ; n13005_not
g28286 not n16200 ; n16200_not
g28287 not n10233 ; n10233_not
g28288 not n10350 ; n10350_not
g28289 not n17001 ; n17001_not
g28290 not n20052 ; n20052_not
g28291 not n11421 ; n11421_not
g28292 not n13041 ; n13041_not
g28293 not n13401 ; n13401_not
g28294 not n11124 ; n11124_not
g28295 not n16020 ; n16020_not
g28296 not n12411 ; n12411_not
g28297 not n14022 ; n14022_not
g28298 not n14031 ; n14031_not
g28299 not n12015 ; n12015_not
g28300 not n12006 ; n12006_not
g28301 not n24003 ; n24003_not
g28302 not n18000 ; n18000_not
g28303 not n11322 ; n11322_not
g28304 not n22005 ; n22005_not
g28305 not n11313 ; n11313_not
g28306 not n15021 ; n15021_not
g28307 not n10503 ; n10503_not
g28308 not n11016 ; n11016_not
g28309 not n22041 ; n22041_not
g28310 not n11601 ; n11601_not
g28311 not n22401 ; n22401_not
g28312 not n23121 ; n23121_not
g28313 not n12303 ; n12303_not
g28314 not n20341 ; n20341_not
g28315 not n10351 ; n10351_not
g28316 not n11503 ; n11503_not
g28317 not n12052 ; n12052_not
g28318 not n11530 ; n11530_not
g28319 not n11233 ; n11233_not
g28320 not n12016 ; n12016_not
g28321 not n23500 ; n23500_not
g28322 not n12124 ; n12124_not
g28323 not n11602 ; n11602_not
g28324 not n12160 ; n12160_not
g28325 not n12232 ; n12232_not
g28326 not n11710 ; n11710_not
g28327 not n11161 ; n11161_not
g28328 not n20440 ; n20440_not
g28329 not n24022 ; n24022_not
g28330 not n11422 ; n11422_not
g28331 not n12304 ; n12304_not
g28332 not n11431 ; n11431_not
g28333 not n11125 ; n11125_not
g28334 not n12340 ; n12340_not
g28335 not n11305 ; n11305_not
g28336 not n16201 ; n16201_not
g28337 not n12403 ; n12403_not
g28338 not n11053 ; n11053_not
g28339 not n12421 ; n12421_not
g28340 not n11017 ; n11017_not
g28341 not n23230 ; n23230_not
g28342 not n12601 ; n12601_not
g28343 not n16021 ; n16021_not
g28344 not n17101 ; n17101_not
g28345 not n20413 ; n20413_not
g28346 not n13330 ; n13330_not
g28347 not n15400 ; n15400_not
g28348 not n13303 ; n13303_not
g28349 not n20611 ; n20611_not
g28350 not n20602 ; n20602_not
g28351 not n21322 ; n21322_not
g28352 not n13222 ; n13222_not
g28353 not n10306 ; n10306_not
g28354 not n13231 ; n13231_not
g28355 not n10324 ; n10324_not
g28356 not n22510 ; n22510_not
g28357 not n13150 ; n13150_not
g28358 not n20530 ; n20530_not
g28359 not n10333 ; n10333_not
g28360 not n21250 ; n21250_not
g28361 not n13123 ; n13123_not
g28362 not n10360 ; n10360_not
g28363 not n13114 ; n13114_not
g28364 not n20503 ; n20503_not
g28365 not n21214 ; n21214_not
g28366 not n10432 ; n10432_not
g28367 not n13051 ; n13051_not
g28368 not n13042 ; n13042_not
g28369 not n13600 ; n13600_not
g28370 not n13006 ; n13006_not
g28371 not n13015 ; n13015_not
g28372 not n21142 ; n21142_not
g28373 not n21070 ; n21070_not
g28374 not n21043 ; n21043_not
g28375 not n21034 ; n21034_not
g28376 not n21106 ; n21106_not
g28377 not n21115 ; n21115_not
g28378 not n21007 ; n21007_not
g28379 not n17002 ; n17002_not
g28380 not n17011 ; n17011_not
g28381 not n20125 ; n20125_not
g28382 not n18001 ; n18001_not
g28383 not n22006 ; n22006_not
g28384 not n22042 ; n22042_not
g28385 not n22114 ; n22114_not
g28386 not n21610 ; n21610_not
g28387 not n14401 ; n14401_not
g28388 not n22150 ; n22150_not
g28389 not n22222 ; n22222_not
g28390 not n14221 ; n14221_not
g28391 not n20161 ; n20161_not
g28392 not n21502 ; n21502_not
g28393 not n14113 ; n14113_not
g28394 not n20710 ; n20710_not
g28395 not n21430 ; n21430_not
g28396 not n14032 ; n14032_not
g28397 not n22330 ; n22330_not
g28398 not n13411 ; n13411_not
g28399 not n13402 ; n13402_not
g28400 not n22402 ; n22402_not
g28401 not n10126 ; n10126_not
g28402 not n10135 ; n10135_not
g28403 not n15103 ; n15103_not
g28404 not n20053 ; n20053_not
g28405 not n20017 ; n20017_not
g28406 not n10171 ; n10171_not
g28407 not n20305 ; n20305_not
g28408 not n10162 ; n10162_not
g28409 not n15130 ; n15130_not
g28410 not n20233 ; n20233_not
g28411 not n10207 ; n10207_not
g28412 not n10720 ; n10720_not
g28413 not n10810 ; n10810_not
g28414 not n10243 ; n10243_not
g28415 not n10234 ; n10234_not
g28416 not n10801 ; n10801_not
g28417 not n15211 ; n15211_not
g28418 not n10270 ; n10270_not
g28419 not n17200 ; n17200_not
g28420 not n15202 ; n15202_not
g28421 not n23014 ; n23014_not
g28422 not n10504 ; n10504_not
g28423 not n15022 ; n15022_not
g28424 not n10027 ; n10027_not
g28425 not n10018 ; n10018_not
g28426 not n15031 ; n15031_not
g28427 not n13510 ; n13510_not
g28428 not n10540 ; n10540_not
g28429 not n23122 ; n23122_not
g28430 not n24004 ; n24004_not
g28431 not n13501 ; n13501_not
g28432 not n10054 ; n10054_not
g28433 not n10612 ; n10612_not
g28434 not n10090 ; n10090_not
g28435 not n23050 ; n23050_not
g28436 not n21151 ; n21151_not
g28437 not n21160 ; n21160_not
g28438 not n10063 ; n10063_not
g28439 not n11324 ; n11324_not
g28440 not n11027 ; n11027_not
g28441 not n20504 ; n20504_not
g28442 not n11063 ; n11063_not
g28443 not n23123 ; n23123_not
g28444 not n11054 ; n11054_not
g28445 not n11018 ; n11018_not
g28446 not n23132 ; n23132_not
g28447 not n11351 ; n11351_not
g28448 not n16031 ; n16031_not
g28449 not n11720 ; n11720_not
g28450 not n11207 ; n11207_not
g28451 not n16022 ; n16022_not
g28452 not n23051 ; n23051_not
g28453 not n20441 ; n20441_not
g28454 not n11171 ; n11171_not
g28455 not n23060 ; n23060_not
g28456 not n20414 ; n20414_not
g28457 not n11162 ; n11162_not
g28458 not n20432 ; n20432_not
g28459 not n11126 ; n11126_not
g28460 not n11234 ; n11234_not
g28461 not n11243 ; n11243_not
g28462 not n11135 ; n11135_not
g28463 not n11270 ; n11270_not
g28464 not n23024 ; n23024_not
g28465 not n23015 ; n23015_not
g28466 not n11090 ; n11090_not
g28467 not n11612 ; n11612_not
g28468 not n12017 ; n12017_not
g28469 not n14060 ; n14060_not
g28470 not n14033 ; n14033_not
g28471 not n21611 ; n21611_not
g28472 not n21620 ; n21620_not
g28473 not n15401 ; n15401_not
g28474 not n21800 ; n21800_not
g28475 not n22601 ; n22601_not
g28476 not n13601 ; n13601_not
g28477 not n22007 ; n22007_not
g28478 not n13511 ; n13511_not
g28479 not n22016 ; n22016_not
g28480 not n22052 ; n22052_not
g28481 not n22043 ; n22043_not
g28482 not n21161 ; n21161_not
g28483 not n13412 ; n13412_not
g28484 not n22124 ; n22124_not
g28485 not n22115 ; n22115_not
g28486 not n22151 ; n22151_not
g28487 not n13340 ; n13340_not
g28488 not n22160 ; n22160_not
g28489 not n13304 ; n13304_not
g28490 not n20423 ; n20423_not
g28491 not n12710 ; n12710_not
g28492 not n21116 ; n21116_not
g28493 not n14222 ; n14222_not
g28494 not n14231 ; n14231_not
g28495 not n14150 ; n14150_not
g28496 not n14114 ; n14114_not
g28497 not n14123 ; n14123_not
g28498 not n14303 ; n14303_not
g28499 not n14330 ; n14330_not
g28500 not n14051 ; n14051_not
g28501 not n21224 ; n21224_not
g28502 not n21215 ; n21215_not
g28503 not n21251 ; n21251_not
g28504 not n21260 ; n21260_not
g28505 not n14411 ; n14411_not
g28506 not n14402 ; n14402_not
g28507 not n21323 ; n21323_not
g28508 not n15032 ; n15032_not
g28509 not n21332 ; n21332_not
g28510 not n15104 ; n15104_not
g28511 not n14510 ; n14510_not
g28512 not n21404 ; n21404_not
g28513 not n15140 ; n15140_not
g28514 not n21440 ; n21440_not
g28515 not n21431 ; n21431_not
g28516 not n15212 ; n15212_not
g28517 not n21512 ; n21512_not
g28518 not n21503 ; n21503_not
g28519 not n20207 ; n20207_not
g28520 not n20900 ; n20900_not
g28521 not n20162 ; n20162_not
g28522 not n20171 ; n20171_not
g28523 not n22511 ; n22511_not
g28524 not n22520 ; n22520_not
g28525 not n20135 ; n20135_not
g28526 not n23303 ; n23303_not
g28527 not n20126 ; n20126_not
g28528 not n12422 ; n12422_not
g28529 not n20090 ; n20090_not
g28530 not n20063 ; n20063_not
g28531 not n23330 ; n23330_not
g28532 not n12341 ; n12341_not
g28533 not n20054 ; n20054_not
g28534 not n12305 ; n12305_not
g28535 not n20018 ; n20018_not
g28536 not n20027 ; n20027_not
g28537 not n20720 ; n20720_not
g28538 not n12233 ; n12233_not
g28539 not n12161 ; n12161_not
g28540 not n20612 ; n20612_not
g28541 not n22700 ; n22700_not
g28542 not n12125 ; n12125_not
g28543 not n20540 ; n20540_not
g28544 not n12053 ; n12053_not
g28545 not n23501 ; n23501_not
g28546 not n13232 ; n13232_not
g28547 not n22223 ; n22223_not
g28548 not n22232 ; n22232_not
g28549 not n12602 ; n12602_not
g28550 not n12611 ; n12611_not
g28551 not n13160 ; n13160_not
g28552 not n21080 ; n21080_not
g28553 not n13124 ; n13124_not
g28554 not n12530 ; n12530_not
g28555 not n12503 ; n12503_not
g28556 not n13052 ; n13052_not
g28557 not n20351 ; n20351_not
g28558 not n13016 ; n13016_not
g28559 not n20342 ; n20342_not
g28560 not n12431 ; n12431_not
g28561 not n22304 ; n22304_not
g28562 not n21044 ; n21044_not
g28563 not n22340 ; n22340_not
g28564 not n22331 ; n22331_not
g28565 not n20306 ; n20306_not
g28566 not n20315 ; n20315_not
g28567 not n21008 ; n21008_not
g28568 not n20270 ; n20270_not
g28569 not n22412 ; n22412_not
g28570 not n22403 ; n22403_not
g28571 not n20234 ; n20234_not
g28572 not n20243 ; n20243_not
g28573 not n12152 ; n12152_not
g28574 not n10208 ; n10208_not
g28575 not n16130 ; n16130_not
g28576 not n17201 ; n17201_not
g28577 not n24410 ; n24410_not
g28578 not n10433 ; n10433_not
g28579 not n10172 ; n10172_not
g28580 not n10334 ; n10334_not
g28581 not n18110 ; n18110_not
g28582 not n10910 ; n10910_not
g28583 not n24023 ; n24023_not
g28584 not n11432 ; n11432_not
g28585 not n11333 ; n11333_not
g28586 not n23204 ; n23204_not
g28587 not n11342 ; n11342_not
g28588 not n10028 ; n10028_not
g28589 not n16310 ; n16310_not
g28590 not n24050 ; n24050_not
g28591 not n16211 ; n16211_not
g28592 not n23231 ; n23231_not
g28593 not n23240 ; n23240_not
g28594 not n16202 ; n16202_not
g28595 not n10136 ; n10136_not
g28596 not n24005 ; n24005_not
g28597 not n17102 ; n17102_not
g28598 not n10064 ; n10064_not
g28599 not n10361 ; n10361_not
g28600 not n10613 ; n10613_not
g28601 not n24032 ; n24032_not
g28602 not n18011 ; n18011_not
g28603 not n10280 ; n10280_not
g28604 not n16103 ; n16103_not
g28605 not n18002 ; n18002_not
g28606 not n17012 ; n17012_not
g28607 not n10721 ; n10721_not
g28608 not n10505 ; n10505_not
g28609 not n24041 ; n24041_not
g28610 not n11504 ; n11504_not
g28611 not n11540 ; n11540_not
g28612 not n10244 ; n10244_not
g28613 not n10541 ; n10541_not
g28614 not n11604 ; n11604_not
g28615 not n22161 ; n22161_not
g28616 not n12720 ; n12720_not
g28617 not n10065 ; n10065_not
g28618 not n22233 ; n22233_not
g28619 not n10371 ; n10371_not
g28620 not n21144 ; n21144_not
g28621 not n12315 ; n12315_not
g28622 not n12306 ; n12306_not
g28623 not n12162 ; n12162_not
g28624 not n12171 ; n12171_not
g28625 not n14160 ; n14160_not
g28626 not n10407 ; n10407_not
g28627 not n10920 ; n10920_not
g28628 not n16320 ; n16320_not
g28629 not n15240 ; n15240_not
g28630 not n14124 ; n14124_not
g28631 not n14340 ; n14340_not
g28632 not n15213 ; n15213_not
g28633 not n21513 ; n21513_not
g28634 not n11244 ; n11244_not
g28635 not n12234 ; n12234_not
g28636 not n15303 ; n15303_not
g28637 not n20505 ; n20505_not
g28638 not n14232 ; n14232_not
g28639 not n12243 ; n12243_not
g28640 not n23610 ; n23610_not
g28641 not n10722 ; n10722_not
g28642 not n20541 ; n20541_not
g28643 not n10731 ; n10731_not
g28644 not n12270 ; n12270_not
g28645 not n10362 ; n10362_not
g28646 not n12207 ; n12207_not
g28647 not n10029 ; n10029_not
g28648 not n13611 ; n13611_not
g28649 not n13602 ; n13602_not
g28650 not n11208 ; n11208_not
g28651 not n24033 ; n24033_not
g28652 not n15330 ; n15330_not
g28653 not n20613 ; n20613_not
g28654 not n23133 ; n23133_not
g28655 not n11280 ; n11280_not
g28656 not n21225 ; n21225_not
g28657 not n13710 ; n13710_not
g28658 not n14304 ; n14304_not
g28659 not n10173 ; n10173_not
g28660 not n12018 ; n12018_not
g28661 not n12027 ; n12027_not
g28662 not n18300 ; n18300_not
g28663 not n15402 ; n15402_not
g28664 not n10308 ; n10308_not
g28665 not n23241 ; n23241_not
g28666 not n15411 ; n15411_not
g28667 not n17013 ; n17013_not
g28668 not n21405 ; n21405_not
g28669 not n10470 ; n10470_not
g28670 not n16032 ; n16032_not
g28671 not n10209 ; n10209_not
g28672 not n10245 ; n10245_not
g28673 not n16140 ; n16140_not
g28674 not n12540 ; n12540_not
g28675 not n10542 ; n10542_not
g28676 not n11064 ; n11064_not
g28677 not n22341 ; n22341_not
g28678 not n15510 ; n15510_not
g28679 not n12405 ; n12405_not
g28680 not n21333 ; n21333_not
g28681 not n12504 ; n12504_not
g28682 not n11028 ; n11028_not
g28683 not n23322 ; n23322_not
g28684 not n12432 ; n12432_not
g28685 not n10506 ; n10506_not
g28686 not n16104 ; n16104_not
g28687 not n10515 ; n10515_not
g28688 not n11910 ; n11910_not
g28689 not n10281 ; n10281_not
g28690 not n22413 ; n22413_not
g28691 not n12135 ; n12135_not
g28692 not n12126 ; n12126_not
g28693 not n20721 ; n20721_not
g28694 not n11172 ; n11172_not
g28695 not n10650 ; n10650_not
g28696 not n24042 ; n24042_not
g28697 not n20901 ; n20901_not
g28698 not n10344 ; n10344_not
g28699 not n10137 ; n10137_not
g28700 not n12090 ; n12090_not
g28701 not n23205 ; n23205_not
g28702 not n10443 ; n10443_not
g28703 not n21441 ; n21441_not
g28704 not n10434 ; n10434_not
g28705 not n14052 ; n14052_not
g28706 not n23340 ; n23340_not
g28707 not n10335 ; n10335_not
g28708 not n14034 ; n14034_not
g28709 not n10317 ; n10317_not
g28710 not n24051 ; n24051_not
g28711 not n16212 ; n16212_not
g28712 not n22521 ; n22521_not
g28713 not n14061 ; n14061_not
g28714 not n21261 ; n21261_not
g28715 not n12054 ; n12054_not
g28716 not n12063 ; n12063_not
g28717 not n22305 ; n22305_not
g28718 not n10614 ; n10614_not
g28719 not n10623 ; n10623_not
g28720 not n11136 ; n11136_not
g28721 not n12612 ; n12612_not
g28722 not n20208 ; n20208_not
g28723 not n13053 ; n13053_not
g28724 not n14043 ; n14043_not
g28725 not n20028 ; n20028_not
g28726 not n15231 ; n15231_not
g28727 not n24510 ; n24510_not
g28728 not n14007 ; n14007_not
g28729 not n23025 ; n23025_not
g28730 not n20244 ; n20244_not
g28731 not n13017 ; n13017_not
g28732 not n18012 ; n18012_not
g28733 not n13413 ; n13413_not
g28734 not n22017 ; n22017_not
g28735 not n10821 ; n10821_not
g28736 not n12423 ; n12423_not
g28737 not n20280 ; n20280_not
g28738 not n10830 ; n10830_not
g28739 not n14520 ; n14520_not
g28740 not n11361 ; n11361_not
g28741 not n15033 ; n15033_not
g28742 not n24411 ; n24411_not
g28743 not n23502 ; n23502_not
g28744 not n22053 ; n22053_not
g28745 not n11343 ; n11343_not
g28746 not n13233 ; n13233_not
g28747 not n11541 ; n11541_not
g28748 not n21117 ; n21117_not
g28749 not n21801 ; n21801_not
g28750 not n11505 ; n11505_not
g28751 not n20136 ; n20136_not
g28752 not n11613 ; n11613_not
g28753 not n24006 ; n24006_not
g28754 not n24015 ; n24015_not
g28755 not n13305 ; n13305_not
g28756 not n13161 ; n13161_not
g28757 not n21081 ; n21081_not
g28758 not n23331 ; n23331_not
g28759 not n17211 ; n17211_not
g28760 not n19110 ; n19110_not
g28761 not n17202 ; n17202_not
g28762 not n13125 ; n13125_not
g28763 not n13341 ; n13341_not
g28764 not n20172 ; n20172_not
g28765 not n23403 ; n23403_not
g28766 not n20064 ; n20064_not
g28767 not n21180 ; n21180_not
g28768 not n11721 ; n11721_not
g28769 not n17310 ; n17310_not
g28770 not n11433 ; n11433_not
g28771 not n23511 ; n23511_not
g28772 not n13530 ; n13530_not
g28773 not n23430 ; n23430_not
g28774 not n20424 ; n20424_not
g28775 not n12342 ; n12342_not
g28776 not n10812 ; n10812_not
g28777 not n12351 ; n12351_not
g28778 not n22701 ; n22701_not
g28779 not n20352 ; n20352_not
g28780 not n14412 ; n14412_not
g28781 not n12900 ; n12900_not
g28782 not n15105 ; n15105_not
g28783 not n21009 ; n21009_not
g28784 not n21045 ; n21045_not
g28785 not n18120 ; n18120_not
g28786 not n21621 ; n21621_not
g28787 not n20316 ; n20316_not
g28788 not n23061 ; n23061_not
g28789 not n20433 ; n20433_not
g28790 not n15141 ; n15141_not
g28791 not n20442 ; n20442_not
g28792 not n22125 ; n22125_not
g28793 not n21136 ; n21136_not
g28794 not n15007 ; n15007_not
g28795 not n18400 ; n18400_not
g28796 not n21118 ; n21118_not
g28797 not n12901 ; n12901_not
g28798 not n10309 ; n10309_not
g28799 not n21163 ; n21163_not
g28800 not n15214 ; n15214_not
g28801 not n16033 ; n16033_not
g28802 not n17113 ; n17113_not
g28803 not n10660 ; n10660_not
g28804 not n10291 ; n10291_not
g28805 not n10282 ; n10282_not
g28806 not n15106 ; n15106_not
g28807 not n23242 ; n23242_not
g28808 not n10336 ; n10336_not
g28809 not n15223 ; n15223_not
g28810 not n23134 ; n23134_not
g28811 not n13315 ; n13315_not
g28812 not n10219 ; n10219_not
g28813 not n13306 ; n13306_not
g28814 not n13540 ; n13540_not
g28815 not n15412 ; n15412_not
g28816 not n10732 ; n10732_not
g28817 not n15151 ; n15151_not
g28818 not n12505 ; n12505_not
g28819 not n13270 ; n13270_not
g28820 not n17212 ; n17212_not
g28821 not n22450 ; n22450_not
g28822 not n17122 ; n17122_not
g28823 not n15142 ; n15142_not
g28824 not n10183 ; n10183_not
g28825 not n10174 ; n10174_not
g28826 not n20614 ; n20614_not
g28827 not n20623 ; n20623_not
g28828 not n21334 ; n21334_not
g28829 not n13243 ; n13243_not
g28830 not n12541 ; n12541_not
g28831 not n22702 ; n22702_not
g28832 not n13234 ; n13234_not
g28833 not n13513 ; n13513_not
g28834 not n12712 ; n12712_not
g28835 not n10246 ; n10246_not
g28836 not n10255 ; n10255_not
g28837 not n17104 ; n17104_not
g28838 not n13126 ; n13126_not
g28839 not n10624 ; n10624_not
g28840 not n13135 ; n13135_not
g28841 not n10444 ; n10444_not
g28842 not n23206 ; n23206_not
g28843 not n15034 ; n15034_not
g28844 not n13063 ; n13063_not
g28845 not n23170 ; n23170_not
g28846 not n13054 ; n13054_not
g28847 not n10372 ; n10372_not
g28848 not n10066 ; n10066_not
g28849 not n10408 ; n10408_not
g28850 not n10831 ; n10831_not
g28851 not n10921 ; n10921_not
g28852 not n13090 ; n13090_not
g28853 not n22810 ; n22810_not
g28854 not n15070 ; n15070_not
g28855 not n12721 ; n12721_not
g28856 not n17320 ; n17320_not
g28857 not n12406 ; n12406_not
g28858 not n21154 ; n21154_not
g28859 not n23062 ; n23062_not
g28860 not n21226 ; n21226_not
g28861 not n20515 ; n20515_not
g28862 not n20506 ; n20506_not
g28863 not n22612 ; n22612_not
g28864 not n22522 ; n22522_not
g28865 not n13207 ; n13207_not
g28866 not n21190 ; n21190_not
g28867 not n10516 ; n10516_not
g28868 not n15115 ; n15115_not
g28869 not n21145 ; n21145_not
g28870 not n15232 ; n15232_not
g28871 not n12613 ; n12613_not
g28872 not n10138 ; n10138_not
g28873 not n23026 ; n23026_not
g28874 not n19120 ; n19120_not
g28875 not n10480 ; n10480_not
g28876 not n22630 ; n22630_not
g28877 not n10552 ; n10552_not
g28878 not n20542 ; n20542_not
g28879 not n13171 ; n13171_not
g28880 not n13162 ; n13162_not
g28881 not n20551 ; n20551_not
g28882 not n21262 ; n21262_not
g28883 not n13018 ; n13018_not
g28884 not n13027 ; n13027_not
g28885 not n15700 ; n15700_not
g28886 not n13504 ; n13504_not
g28887 not n13720 ; n13720_not
g28888 not n15043 ; n15043_not
g28889 not n10147 ; n10147_not
g28890 not n13612 ; n13612_not
g28891 not n15520 ; n15520_not
g28892 not n19300 ; n19300_not
g28893 not n10075 ; n10075_not
g28894 not n17500 ; n17500_not
g28895 not n12028 ; n12028_not
g28896 not n19111 ; n19111_not
g28897 not n24340 ; n24340_not
g28898 not n11470 ; n11470_not
g28899 not n11281 ; n11281_not
g28900 not n14305 ; n14305_not
g28901 not n21550 ; n21550_not
g28902 not n20830 ; n20830_not
g28903 not n23512 ; n23512_not
g28904 not n11443 ; n11443_not
g28905 not n11434 ; n11434_not
g28906 not n14341 ; n14341_not
g28907 not n22162 ; n22162_not
g28908 not n11407 ; n11407_not
g28909 not n24016 ; n24016_not
g28910 not n11920 ; n11920_not
g28911 not n20425 ; n20425_not
g28912 not n14413 ; n14413_not
g28913 not n22126 ; n22126_not
g28914 not n21514 ; n21514_not
g28915 not n11614 ; n11614_not
g28916 not n11623 ; n11623_not
g28917 not n12136 ; n12136_not
g28918 not n19030 ; n19030_not
g28919 not n15241 ; n15241_not
g28920 not n22234 ; n22234_not
g28921 not n11209 ; n11209_not
g28922 not n24034 ; n24034_not
g28923 not n20803 ; n20803_not
g28924 not n11245 ; n11245_not
g28925 not n11542 ; n11542_not
g28926 not n11551 ; n11551_not
g28927 not n14233 ; n14233_not
g28928 not n12064 ; n12064_not
g28929 not n24322 ; n24322_not
g28930 not n11515 ; n11515_not
g28931 not n11506 ; n11506_not
g28932 not n20065 ; n20065_not
g28933 not n17014 ; n17014_not
g28934 not n21910 ; n21910_not
g28935 not n17023 ; n17023_not
g28936 not n21730 ; n21730_not
g28937 not n20173 ; n20173_not
g28938 not n24700 ; n24700_not
g28939 not n21019 ; n21019_not
g28940 not n21127 ; n21127_not
g28941 not n17050 ; n17050_not
g28942 not n17131 ; n17131_not
g28943 not n21055 ; n21055_not
g28944 not n21046 ; n21046_not
g28945 not n21082 ; n21082_not
g28946 not n21802 ; n21802_not
g28947 not n20137 ; n20137_not
g28948 not n11371 ; n11371_not
g28949 not n23620 ; n23620_not
g28950 not n16510 ; n16510_not
g28951 not n21622 ; n21622_not
g28952 not n22090 ; n22090_not
g28953 not n20353 ; n20353_not
g28954 not n20911 ; n20911_not
g28955 not n20902 ; n20902_not
g28956 not n20317 ; n20317_not
g28957 not n18121 ; n18121_not
g28958 not n11362 ; n11362_not
g28959 not n14521 ; n14521_not
g28960 not n22054 ; n22054_not
g28961 not n20281 ; n20281_not
g28962 not n22018 ; n22018_not
g28963 not n18013 ; n18013_not
g28964 not n20245 ; n20245_not
g28965 not n20029 ; n20029_not
g28966 not n23800 ; n23800_not
g28967 not n20209 ; n20209_not
g28968 not n11731 ; n11731_not
g28969 not n21370 ; n21370_not
g28970 not n13351 ; n13351_not
g28971 not n12433 ; n12433_not
g28972 not n13342 ; n13342_not
g28973 not n20731 ; n20731_not
g28974 not n12280 ; n12280_not
g28975 not n20722 ; n20722_not
g28976 not n21442 ; n21442_not
g28977 not n20650 ; n20650_not
g28978 not n22306 ; n22306_not
g28979 not n14062 ; n14062_not
g28980 not n14053 ; n14053_not
g28981 not n12316 ; n12316_not
g28982 not n11137 ; n11137_not
g28983 not n15304 ; n15304_not
g28984 not n13423 ; n13423_not
g28985 not n23332 ; n23332_not
g28986 not n13414 ; n13414_not
g28987 not n22342 ; n22342_not
g28988 not n14710 ; n14710_not
g28989 not n14008 ; n14008_not
g28990 not n23305 ; n23305_not
g28991 not n13450 ; n13450_not
g28992 not n11065 ; n11065_not
g28993 not n12352 ; n12352_not
g28994 not n16213 ; n16213_not
g28995 not n19003 ; n19003_not
g28996 not n16141 ; n16141_not
g28997 not n15340 ; n15340_not
g28998 not n21406 ; n21406_not
g28999 not n11803 ; n11803_not
g29000 not n14044 ; n14044_not
g29001 not n12172 ; n12172_not
g29002 not n23440 ; n23440_not
g29003 not n16105 ; n16105_not
g29004 not n13900 ; n13900_not
g29005 not n14161 ; n14161_not
g29006 not n11650 ; n11650_not
g29007 not n16321 ; n16321_not
g29008 not n12208 ; n12208_not
g29009 not n13531 ; n13531_not
g29010 not n23404 ; n23404_not
g29011 not n14125 ; n14125_not
g29012 not n22414 ; n22414_not
g29013 not n18301 ; n18301_not
g29014 not n11029 ; n11029_not
g29015 not n11722 ; n11722_not
g29016 not n22270 ; n22270_not
g29017 not n12244 ; n12244_not
g29018 not n11173 ; n11173_not
g29019 not n14107 ; n14107_not
g29020 not n19040 ; n19040_not
g29021 not n14342 ; n14342_not
g29022 not n22136 ; n22136_not
g29023 not n14135 ; n14135_not
g29024 not n14351 ; n14351_not
g29025 not n21137 ; n21137_not
g29026 not n24530 ; n24530_not
g29027 not n22127 ; n22127_not
g29028 not n21632 ; n21632_not
g29029 not n12731 ; n12731_not
g29030 not n21227 ; n21227_not
g29031 not n21236 ; n21236_not
g29032 not n10256 ; n10256_not
g29033 not n10292 ; n10292_not
g29034 not n24512 ; n24512_not
g29035 not n18311 ; n18311_not
g29036 not n14243 ; n14243_not
g29037 not n18230 ; n18230_not
g29038 not n14270 ; n14270_not
g29039 not n18203 ; n18203_not
g29040 not n15341 ; n15341_not
g29041 not n12830 ; n12830_not
g29042 not n12722 ; n12722_not
g29043 not n21272 ; n21272_not
g29044 not n10625 ; n10625_not
g29045 not n21263 ; n21263_not
g29046 not n13901 ; n13901_not
g29047 not n15008 ; n15008_not
g29048 not n13316 ; n13316_not
g29049 not n13280 ; n13280_not
g29050 not n21731 ; n21731_not
g29051 not n22172 ; n22172_not
g29052 not n21740 ; n21740_not
g29053 not n24611 ; n24611_not
g29054 not n21128 ; n21128_not
g29055 not n14900 ; n14900_not
g29056 not n14315 ; n14315_not
g29057 not n14162 ; n14162_not
g29058 not n22163 ; n22163_not
g29059 not n21704 ; n21704_not
g29060 not n15413 ; n15413_not
g29061 not n14306 ; n14306_not
g29062 not n21164 ; n21164_not
g29063 not n18302 ; n18302_not
g29064 not n19004 ; n19004_not
g29065 not n14720 ; n14720_not
g29066 not n10661 ; n10661_not
g29067 not n14234 ; n14234_not
g29068 not n24053 ; n24053_not
g29069 not n14171 ; n14171_not
g29070 not n22208 ; n22208_not
g29071 not n13352 ; n13352_not
g29072 not n13244 ; n13244_not
g29073 not n14126 ; n14126_not
g29074 not n21623 ; n21623_not
g29075 not n12803 ; n12803_not
g29076 not n14207 ; n14207_not
g29077 not n21191 ; n21191_not
g29078 not n13514 ; n13514_not
g29079 not n14603 ; n14603_not
g29080 not n15521 ; n15521_not
g29081 not n21452 ; n21452_not
g29082 not n21911 ; n21911_not
g29083 not n21920 ; n21920_not
g29084 not n21560 ; n21560_not
g29085 not n21173 ; n21173_not
g29086 not n21443 ; n21443_not
g29087 not n21551 ; n21551_not
g29088 not n15305 ; n15305_not
g29089 not n15152 ; n15152_not
g29090 not n10148 ; n10148_not
g29091 not n14522 ; n14522_not
g29092 not n13541 ; n13541_not
g29093 not n14531 ; n14531_not
g29094 not n21407 ; n21407_not
g29095 not n21416 ; n21416_not
g29096 not n15242 ; n15242_not
g29097 not n21515 ; n21515_not
g29098 not n15233 ; n15233_not
g29099 not n21524 ; n21524_not
g29100 not n10409 ; n10409_not
g29101 not n10373 ; n10373_not
g29102 not n18401 ; n18401_not
g29103 not n24323 ; n24323_not
g29104 not n15224 ; n15224_not
g29105 not n10445 ; n10445_not
g29106 not n10355 ; n10355_not
g29107 not n10076 ; n10076_not
g29108 not n20471 ; n20471_not
g29109 not n13613 ; n13613_not
g29110 not n18500 ; n18500_not
g29111 not n13721 ; n13721_not
g29112 not n17501 ; n17501_not
g29113 not n10481 ; n10481_not
g29114 not n12902 ; n12902_not
g29115 not n13460 ; n13460_not
g29116 not n22064 ; n22064_not
g29117 not n15044 ; n15044_not
g29118 not n10184 ; n10184_not
g29119 not n21335 ; n21335_not
g29120 not n20444 ; n20444_not
g29121 not n21344 ; n21344_not
g29122 not n24305 ; n24305_not
g29123 not n21146 ; n21146_not
g29124 not n14009 ; n14009_not
g29125 not n17321 ; n17321_not
g29126 not n14423 ; n14423_not
g29127 not n13424 ; n13424_not
g29128 not n14414 ; n14414_not
g29129 not n22091 ; n22091_not
g29130 not n15701 ; n15701_not
g29131 not n21308 ; n21308_not
g29132 not n15116 ; n15116_not
g29133 not n10517 ; n10517_not
g29134 not n21803 ; n21803_not
g29135 not n18023 ; n18023_not
g29136 not n18014 ; n18014_not
g29137 not n10553 ; n10553_not
g29138 not n18050 ; n18050_not
g29139 not n22028 ; n22028_not
g29140 not n15080 ; n15080_not
g29141 not n22019 ; n22019_not
g29142 not n21380 ; n21380_not
g29143 not n21371 ; n21371_not
g29144 not n14045 ; n14045_not
g29145 not n14450 ; n14450_not
g29146 not n22055 ; n22055_not
g29147 not n12920 ; n12920_not
g29148 not n18122 ; n18122_not
g29149 not n18131 ; n18131_not
g29150 not n12911 ; n12911_not
g29151 not n22424 ; n22424_not
g29152 not n10922 ; n10922_not
g29153 not n12029 ; n12029_not
g29154 not n19301 ; n19301_not
g29155 not n20219 ; n20219_not
g29156 not n20912 ; n20912_not
g29157 not n11804 ; n11804_not
g29158 not n11372 ; n11372_not
g29159 not n11660 ; n11660_not
g29160 not n12065 ; n12065_not
g29161 not n22460 ; n22460_not
g29162 not n20516 ; n20516_not
g29163 not n11138 ; n11138_not
g29164 not n22451 ; n22451_not
g29165 not n23801 ; n23801_not
g29166 not n20552 ; n20552_not
g29167 not n16430 ; n16430_not
g29168 not n20183 ; n20183_not
g29169 not n11147 ; n11147_not
g29170 not n16043 ; n16043_not
g29171 not n16034 ; n16034_not
g29172 not n20174 ; n20174_not
g29173 not n22712 ; n22712_not
g29174 not n22703 ; n22703_not
g29175 not n12371 ; n12371_not
g29176 not n22811 ; n22811_not
g29177 not n23108 ; n23108_not
g29178 not n10337 ; n10337_not
g29179 not n22820 ; n22820_not
g29180 not n20453 ; n20453_not
g29181 not n20462 ; n20462_not
g29182 not n20282 ; n20282_not
g29183 not n23252 ; n23252_not
g29184 not n16151 ; n16151_not
g29185 not n20291 ; n20291_not
g29186 not n17123 ; n17123_not
g29187 not n16250 ; n16250_not
g29188 not n16142 ; n16142_not
g29189 not n11291 ; n11291_not
g29190 not n20255 ; n20255_not
g29191 not n20246 ; n20246_not
g29192 not n23513 ; n23513_not
g29193 not n11282 ; n11282_not
g29194 not n22415 ; n22415_not
g29195 not n10931 ; n10931_not
g29196 not n23306 ; n23306_not
g29197 not n22631 ; n22631_not
g29198 not n11255 ; n11255_not
g29199 not n12281 ; n12281_not
g29200 not n20732 ; n20732_not
g29201 not n16007 ; n16007_not
g29202 not n20039 ; n20039_not
g29203 not n12317 ; n12317_not
g29204 not n12416 ; n12416_not
g29205 not n23351 ; n23351_not
g29206 not n12380 ; n12380_not
g29207 not n12407 ; n12407_not
g29208 not n11732 ; n11732_not
g29209 not n10544 ; n10544_not
g29210 not n11219 ; n11219_not
g29211 not n12353 ; n12353_not
g29212 not n23333 ; n23333_not
g29213 not n20804 ; n20804_not
g29214 not n11408 ; n11408_not
g29215 not n20066 ; n20066_not
g29216 not n23207 ; n23207_not
g29217 not n23216 ; n23216_not
g29218 not n20075 ; n20075_not
g29219 not n12137 ; n12137_not
g29220 not n20624 ; n20624_not
g29221 not n23072 ; n23072_not
g29222 not n12173 ; n12173_not
g29223 not n11444 ; n11444_not
g29224 not n17060 ; n17060_not
g29225 not n23441 ; n23441_not
g29226 not n16403 ; n16403_not
g29227 not n23063 ; n23063_not
g29228 not n11183 ; n11183_not
g29229 not n20660 ; n20660_not
g29230 not n17024 ; n17024_not
g29231 not n12209 ; n12209_not
g29232 not n11174 ; n11174_not
g29233 not n22532 ; n22532_not
g29234 not n22523 ; n22523_not
g29235 not n23405 ; n23405_not
g29236 not n20138 ; n20138_not
g29237 not n12245 ; n12245_not
g29238 not n20147 ; n20147_not
g29239 not n11246 ; n11246_not
g29240 not n22640 ; n22640_not
g29241 not n16322 ; n16322_not
g29242 not n20840 ; n20840_not
g29243 not n16115 ; n16115_not
g29244 not n23027 ; n23027_not
g29245 not n12551 ; n12551_not
g29246 not n12542 ; n12542_not
g29247 not n22271 ; n22271_not
g29248 not n16214 ; n16214_not
g29249 not n11066 ; n11066_not
g29250 not n22280 ; n22280_not
g29251 not n20354 ; n20354_not
g29252 not n20363 ; n20363_not
g29253 not n12506 ; n12506_not
g29254 not n12515 ; n12515_not
g29255 not n16700 ; n16700_not
g29256 not n13064 ; n13064_not
g29257 not n19121 ; n19121_not
g29258 not n21056 ; n21056_not
g29259 not n16511 ; n16511_not
g29260 not n12470 ; n12470_not
g29261 not n16520 ; n16520_not
g29262 not n13028 ; n13028_not
g29263 not n11480 ; n11480_not
g29264 not n12434 ; n12434_not
g29265 not n23180 ; n23180_not
g29266 not n12443 ; n12443_not
g29267 not n11336 ; n11336_not
g29268 not n24017 ; n24017_not
g29269 not n23243 ; n23243_not
g29270 not n12650 ; n12650_not
g29271 not n11552 ; n11552_not
g29272 not n13208 ; n13208_not
g29273 not n11039 ; n11039_not
g29274 not n10733 ; n10733_not
g29275 not n23036 ; n23036_not
g29276 not n16070 ; n16070_not
g29277 not n22244 ; n22244_not
g29278 not n23135 ; n23135_not
g29279 not n11345 ; n11345_not
g29280 not n11516 ; n11516_not
g29281 not n20390 ; n20390_not
g29282 not n22235 ; n22235_not
g29283 not n21092 ; n21092_not
g29284 not n11318 ; n11318_not
g29285 not n12623 ; n12623_not
g29286 not n12614 ; n12614_not
g29287 not n13172 ; n13172_not
g29288 not n23144 ; n23144_not
g29289 not n17213 ; n17213_not
g29290 not n16223 ; n16223_not
g29291 not n13136 ; n13136_not
g29292 not n16106 ; n16106_not
g29293 not n11624 ; n11624_not
g29294 not n22307 ; n22307_not
g29295 not n10850 ; n10850_not
g29296 not n22343 ; n22343_not
g29297 not n11363 ; n11363_not
g29298 not n22352 ; n22352_not
g29299 not n11921 ; n11921_not
g29300 not n22316 ; n22316_not
g29301 not n20327 ; n20327_not
g29302 not n23171 ; n23171_not
g29303 not n23621 ; n23621_not
g29304 not n20318 ; n20318_not
g29305 not n17141 ; n17141_not
g29306 not n14073 ; n14073_not
g29307 not n10626 ; n10626_not
g29308 not n11292 ; n11292_not
g29309 not n14082 ; n14082_not
g29310 not n17511 ; n17511_not
g29311 not n20292 ; n20292_not
g29312 not n13902 ; n13902_not
g29313 not n10662 ; n10662_not
g29314 not n14604 ; n14604_not
g29315 not n17502 ; n17502_not
g29316 not n14064 ; n14064_not
g29317 not n11148 ; n11148_not
g29318 not n10770 ; n10770_not
g29319 not n22065 ; n22065_not
g29320 not n14019 ; n14019_not
g29321 not n21453 ; n21453_not
g29322 not n23622 ; n23622_not
g29323 not n23406 ; n23406_not
g29324 not n17610 ; n17610_not
g29325 not n20733 ; n20733_not
g29326 not n13911 ; n13911_not
g29327 not n15045 ; n15045_not
g29328 not n23415 ; n23415_not
g29329 not n15009 ; n15009_not
g29330 not n13803 ; n13803_not
g29331 not n12354 ; n12354_not
g29332 not n21633 ; n21633_not
g29333 not n11076 ; n11076_not
g29334 not n19311 ; n19311_not
g29335 not n19302 ; n19302_not
g29336 not n21417 ; n21417_not
g29337 not n12372 ; n12372_not
g29338 not n24360 ; n24360_not
g29339 not n17430 ; n17430_not
g29340 not n11373 ; n11373_not
g29341 not n24018 ; n24018_not
g29342 not n18024 ; n18024_not
g29343 not n10590 ; n10590_not
g29344 not n22137 ; n22137_not
g29345 not n11409 ; n11409_not
g29346 not n21561 ; n21561_not
g29347 not n19230 ; n19230_not
g29348 not n15603 ; n15603_not
g29349 not n20463 ; n20463_not
g29350 not n16224 ; n16224_not
g29351 not n18204 ; n18204_not
g29352 not n10635 ; n10635_not
g29353 not n14352 ; n14352_not
g29354 not n10149 ; n10149_not
g29355 not n24513 ; n24513_not
g29356 not n15630 ; n15630_not
g29357 not n16260 ; n16260_not
g29358 not n15153 ; n15153_not
g29359 not n22281 ; n22281_not
g29360 not n14424 ; n14424_not
g29361 not n18060 ; n18060_not
g29362 not n21525 ; n21525_not
g29363 not n19203 ; n19203_not
g29364 not n19122 ; n19122_not
g29365 not n14208 ; n14208_not
g29366 not n10806 ; n10806_not
g29367 not n20553 ; n20553_not
g29368 not n20364 ; n20364_not
g29369 not n18240 ; n18240_not
g29370 not n14460 ; n14460_not
g29371 not n16404 ; n16404_not
g29372 not n14280 ; n14280_not
g29373 not n16521 ; n16521_not
g29374 not n15225 ; n15225_not
g29375 not n20517 ; n20517_not
g29376 not n22173 ; n22173_not
g29377 not n11346 ; n11346_not
g29378 not n24342 ; n24342_not
g29379 not n13650 ; n13650_not
g29380 not n14244 ; n14244_not
g29381 not n22209 ; n22209_not
g29382 not n23550 ; n23550_not
g29383 not n10734 ; n10734_not
g29384 not n17403 ; n17403_not
g29385 not n10743 ; n10743_not
g29386 not n19131 ; n19131_not
g29387 not n15081 ; n15081_not
g29388 not n11256 ; n11256_not
g29389 not n14532 ; n14532_not
g29390 not n20256 ; n20256_not
g29391 not n10851 ; n10851_not
g29392 not n10671 ; n10671_not
g29393 not n23631 ; n23631_not
g29394 not n13551 ; n13551_not
g29395 not n13542 ; n13542_not
g29396 not n14136 ; n14136_not
g29397 not n22245 ; n22245_not
g29398 not n10077 ; n10077_not
g29399 not n20328 ; n20328_not
g29400 not n22029 ; n22029_not
g29401 not n15711 ; n15711_not
g29402 not n16440 ; n16440_not
g29403 not n14316 ; n14316_not
g29404 not n13731 ; n13731_not
g29405 not n15702 ; n15702_not
g29406 not n13722 ; n13722_not
g29407 not n16332 ; n16332_not
g29408 not n20661 ; n20661_not
g29409 not n15117 ; n15117_not
g29410 not n14172 ; n14172_not
g29411 not n11184 ; n11184_not
g29412 not n18132 ; n18132_not
g29413 not n15810 ; n15810_not
g29414 not n20625 ; n20625_not
g29415 not n13830 ; n13830_not
g29416 not n24441 ; n24441_not
g29417 not n20481 ; n20481_not
g29418 not n10707 ; n10707_not
g29419 not n11805 ; n11805_not
g29420 not n13623 ; n13623_not
g29421 not n13614 ; n13614_not
g29422 not n22641 ; n22641_not
g29423 not n11661 ; n11661_not
g29424 not n15900 ; n15900_not
g29425 not n14721 ; n14721_not
g29426 not n12291 ; n12291_not
g29427 not n12282 ; n12282_not
g29428 not n12840 ; n12840_not
g29429 not n17151 ; n17151_not
g29430 not n23514 ; n23514_not
g29431 not n12318 ; n12318_not
g29432 not n12327 ; n12327_not
g29433 not n22713 ; n22713_not
g29434 not n20076 ; n20076_not
g29435 not n23523 ; n23523_not
g29436 not n10860 ; n10860_not
g29437 not n13524 ; n13524_not
g29438 not n21165 ; n21165_not
g29439 not n23109 ; n23109_not
g29440 not n12363 ; n12363_not
g29441 not n13515 ; n13515_not
g29442 not n15342 ; n15342_not
g29443 not n15351 ; n15351_not
g29444 not n14091 ; n14091_not
g29445 not n12174 ; n12174_not
g29446 not n12183 ; n12183_not
g29447 not n12732 ; n12732_not
g29448 not n23181 ; n23181_not
g29449 not n24306 ; n24306_not
g29450 not n12219 ; n12219_not
g29451 not n14901 ; n14901_not
g29452 not n15315 ; n15315_not
g29453 not n10383 ; n10383_not
g29454 not n18501 ; n18501_not
g29455 not n15306 ; n15306_not
g29456 not n10374 ; n10374_not
g29457 not n23910 ; n23910_not
g29458 not n12246 ; n12246_not
g29459 not n23334 ; n23334_not
g29460 not n12255 ; n12255_not
g29461 not n12804 ; n12804_not
g29462 not n23145 ; n23145_not
g29463 not n10824 ; n10824_not
g29464 not n13029 ; n13029_not
g29465 not n13065 ; n13065_not
g29466 not n13353 ; n13353_not
g29467 not n23370 ; n23370_not
g29468 not n19410 ; n19410_not
g29469 not n21084 ; n21084_not
g29470 not n13137 ; n13137_not
g29471 not n19104 ; n19104_not
g29472 not n13317 ; n13317_not
g29473 not n11517 ; n11517_not
g29474 not n21129 ; n21129_not
g29475 not n19005 ; n19005_not
g29476 not n13173 ; n13173_not
g29477 not n21093 ; n21093_not
g29478 not n13281 ; n13281_not
g29479 not n19041 ; n19041_not
g29480 not n13209 ; n13209_not
g29481 not n13245 ; n13245_not
g29482 not n11553 ; n11553_not
g29483 not n12912 ; n12912_not
g29484 not n12921 ; n12921_not
g29485 not n11481 ; n11481_not
g29486 not n12930 ; n12930_not
g29487 not n16701 ; n16701_not
g29488 not n23442 ; n23442_not
g29489 not n20148 ; n20148_not
g29490 not n10833 ; n10833_not
g29491 not n23073 ; n23073_not
g29492 not n13461 ; n13461_not
g29493 not n21741 ; n21741_not
g29494 not n17142 ; n17142_not
g29495 not n22821 ; n22821_not
g29496 not n21813 ; n21813_not
g29497 not n15072 ; n15072_not
g29498 not n23037 ; n23037_not
g29499 not n23451 ; n23451_not
g29500 not n21057 ; n21057_not
g29501 not n13425 ; n13425_not
g29502 not n11625 ; n11625_not
g29503 not n12444 ; n12444_not
g29504 not n17025 ; n17025_not
g29505 not n17250 ; n17250_not
g29506 not n18312 ; n18312_not
g29507 not n23307 ; n23307_not
g29508 not n21345 ; n21345_not
g29509 not n11931 ; n11931_not
g29510 not n11922 ; n11922_not
g29511 not n12480 ; n12480_not
g29512 not n16080 ; n16080_not
g29513 not n15450 ; n15450_not
g29514 not n22425 ; n22425_not
g29515 not n11733 ; n11733_not
g29516 not n20184 ; n20184_not
g29517 not n17223 ; n17223_not
g29518 not n21705 ; n21705_not
g29519 not n10482 ; n10482_not
g29520 not n16044 ; n16044_not
g29521 not n12516 ; n12516_not
g29522 not n10185 ; n10185_not
g29523 not n22317 ; n22317_not
g29524 not n12381 ; n12381_not
g29525 not n10554 ; n10554_not
g29526 not n20805 ; n20805_not
g29527 not n17322 ; n17322_not
g29528 not n10563 ; n10563_not
g29529 not n16152 ; n16152_not
g29530 not n15531 ; n15531_not
g29531 not n15522 ; n15522_not
g29532 not n12408 ; n12408_not
g29533 not n22353 ; n22353_not
g29534 not n10527 ; n10527_not
g29535 not n17331 ; n17331_not
g29536 not n21381 ; n21381_not
g29537 not n10257 ; n10257_not
g29538 not n23703 ; n23703_not
g29539 not n16116 ; n16116_not
g29540 not n10518 ; n10518_not
g29541 not n20841 ; n20841_not
g29542 not n23802 ; n23802_not
g29543 not n10455 ; n10455_not
g29544 not n21273 ; n21273_not
g29545 not n22533 ; n22533_not
g29546 not n10446 ; n10446_not
g29547 not n23811 ; n23811_not
g29548 not n23730 ; n23730_not
g29549 not n12075 ; n12075_not
g29550 not n12066 ; n12066_not
g29551 not n12624 ; n12624_not
g29552 not n23217 ; n23217_not
g29553 not n16008 ; n16008_not
g29554 not n12660 ; n12660_not
g29555 not n10932 ; n10932_not
g29556 not n10419 ; n10419_not
g29557 not n17214 ; n17214_not
g29558 not n20913 ; n20913_not
g29559 not n12147 ; n12147_not
g29560 not n21237 ; n21237_not
g29561 not n12138 ; n12138_not
g29562 not n18402 ; n18402_not
g29563 not n10491 ; n10491_not
g29564 not n12552 ; n12552_not
g29565 not n11445 ; n11445_not
g29566 not n15423 ; n15423_not
g29567 not n21921 ; n21921_not
g29568 not n24612 ; n24612_not
g29569 not n10293 ; n10293_not
g29570 not n23253 ; n23253_not
g29571 not n22461 ; n22461_not
g29572 not n21309 ; n21309_not
g29573 not n15414 ; n15414_not
g29574 not n17061 ; n17061_not
g29575 not n12039 ; n12039_not
g29576 not n21634 ; n21634_not
g29577 not n21058 ; n21058_not
g29578 not n21706 ; n21706_not
g29579 not n17026 ; n17026_not
g29580 not n21742 ; n21742_not
g29581 not n17035 ; n17035_not
g29582 not n21670 ; n21670_not
g29583 not n20923 ; n20923_not
g29584 not n17143 ; n17143_not
g29585 not n18061 ; n18061_not
g29586 not n18025 ; n18025_not
g29587 not n20149 ; n20149_not
g29588 not n20257 ; n20257_not
g29589 not n20077 ; n20077_not
g29590 not n20185 ; n20185_not
g29591 not n20950 ; n20950_not
g29592 not n17062 ; n17062_not
g29593 not n17620 ; n17620_not
g29594 not n17071 ; n17071_not
g29595 not n20914 ; n20914_not
g29596 not n21166 ; n21166_not
g29597 not n15640 ; n15640_not
g29598 not n15019 ; n15019_not
g29599 not n21148 ; n21148_not
g29600 not n15901 ; n15901_not
g29601 not n15604 ; n15604_not
g29602 not n15271 ; n15271_not
g29603 not n21184 ; n21184_not
g29604 not n19204 ; n19204_not
g29605 not n17404 ; n17404_not
g29606 not n20491 ; n20491_not
g29607 not n17116 ; n17116_not
g29608 not n19240 ; n19240_not
g29609 not n21238 ; n21238_not
g29610 not n20527 ; n20527_not
g29611 not n20518 ; n20518_not
g29612 not n15532 ; n15532_not
g29613 not n18610 ; n18610_not
g29614 not n14911 ; n14911_not
g29615 not n16009 ; n16009_not
g29616 not n14902 ; n14902_not
g29617 not n21274 ; n21274_not
g29618 not n20554 ; n20554_not
g29619 not n20563 ; n20563_not
g29620 not n19312 ; n19312_not
g29621 not n20590 ; n20590_not
g29622 not n15460 ; n15460_not
g29623 not n17440 ; n17440_not
g29624 not n17224 ; n17224_not
g29625 not n19042 ; n19042_not
g29626 not n19060 ; n19060_not
g29627 not n16603 ; n16603_not
g29628 not n15154 ; n15154_not
g29629 not n15163 ; n15163_not
g29630 not n17260 ; n17260_not
g29631 not n15190 ; n15190_not
g29632 not n16630 ; n16630_not
g29633 not n15127 ; n15127_not
g29634 not n15820 ; n15820_not
g29635 not n15118 ; n15118_not
g29636 not n16522 ; n16522_not
g29637 not n16531 ; n16531_not
g29638 not n15712 ; n15712_not
g29639 not n15244 ; n15244_not
g29640 not n17152 ; n17152_not
g29641 not n15082 ; n15082_not
g29642 not n15091 ; n15091_not
g29643 not n19132 ; n19132_not
g29644 not n17125 ; n17125_not
g29645 not n18511 ; n18511_not
g29646 not n15055 ; n15055_not
g29647 not n15046 ; n15046_not
g29648 not n17332 ; n17332_not
g29649 not n16702 ; n16702_not
g29650 not n16711 ; n16711_not
g29651 not n18502 ; n18502_not
g29652 not n19015 ; n19015_not
g29653 not n15262 ; n15262_not
g29654 not n15253 ; n15253_not
g29655 not n19006 ; n19006_not
g29656 not n21490 ; n21490_not
g29657 not n20770 ; n20770_not
g29658 not n16333 ; n16333_not
g29659 not n19051 ; n19051_not
g29660 not n16405 ; n16405_not
g29661 not n18241 ; n18241_not
g29662 not n21526 ; n21526_not
g29663 not n20815 ; n20815_not
g29664 not n20806 ; n20806_not
g29665 not n16441 ; n16441_not
g29666 not n20482 ; n20482_not
g29667 not n21562 ; n21562_not
g29668 not n20842 ; n20842_not
g29669 not n20851 ; n20851_not
g29670 not n18205 ; n18205_not
g29671 not n17512 ; n17512_not
g29672 not n18133 ; n18133_not
g29673 not n16504 ; n16504_not
g29674 not n20365 ; n20365_not
g29675 not n20329 ; n20329_not
g29676 not n20293 ; n20293_not
g29677 not n19420 ; n19420_not
g29678 not n16045 ; n16045_not
g29679 not n14830 ; n14830_not
g29680 not n15424 ; n15424_not
g29681 not n21346 ; n21346_not
g29682 not n20626 ; n20626_not
g29683 not n20635 ; n20635_not
g29684 not n14803 ; n14803_not
g29685 not n16081 ; n16081_not
g29686 not n18313 ; n18313_not
g29687 not n16117 ; n16117_not
g29688 not n21382 ; n21382_not
g29689 not n20671 ; n20671_not
g29690 not n20662 ; n20662_not
g29691 not n15352 ; n15352_not
g29692 not n14722 ; n14722_not
g29693 not n14731 ; n14731_not
g29694 not n16153 ; n16153_not
g29695 not n21418 ; n21418_not
g29696 not n20707 ; n20707_not
g29697 not n16810 ; n16810_not
g29698 not n15316 ; n15316_not
g29699 not n19600 ; n19600_not
g29700 not n16225 ; n16225_not
g29701 not n16324 ; n16324_not
g29702 not n16261 ; n16261_not
g29703 not n21454 ; n21454_not
g29704 not n20743 ; n20743_not
g29705 not n20734 ; n20734_not
g29706 not n12661 ; n12661_not
g29707 not n12733 ; n12733_not
g29708 not n23182 ; n23182_not
g29709 not n12805 ; n12805_not
g29710 not n23146 ; n23146_not
g29711 not n12841 ; n12841_not
g29712 not n12913 ; n12913_not
g29713 not n23074 ; n23074_not
g29714 not n12409 ; n12409_not
g29715 not n23038 ; n23038_not
g29716 not n22930 ; n22930_not
g29717 not n22822 ; n22822_not
g29718 not n13480 ; n13480_not
g29719 not n13462 ; n13462_not
g29720 not n13516 ; n13516_not
g29721 not n22750 ; n22750_not
g29722 not n22714 ; n22714_not
g29723 not n13552 ; n13552_not
g29724 not n12292 ; n12292_not
g29725 not n11770 ; n11770_not
g29726 not n12328 ; n12328_not
g29727 not n11815 ; n11815_not
g29728 not n11806 ; n11806_not
g29729 not n12364 ; n12364_not
g29730 not n12373 ; n12373_not
g29731 not n12382 ; n12382_not
g29732 not n11842 ; n11842_not
g29733 not n12427 ; n12427_not
g29734 not n12445 ; n12445_not
g29735 not n23290 ; n23290_not
g29736 not n12481 ; n12481_not
g29737 not n12517 ; n12517_not
g29738 not n12553 ; n12553_not
g29739 not n23254 ; n23254_not
g29740 not n12625 ; n12625_not
g29741 not n23218 ; n23218_not
g29742 not n22462 ; n22462_not
g29743 not n13282 ; n13282_not
g29744 not n22426 ; n22426_not
g29745 not n13327 ; n13327_not
g29746 not n13318 ; n13318_not
g29747 not n13912 ; n13912_not
g29748 not n13354 ; n13354_not
g29749 not n13363 ; n13363_not
g29750 not n22390 ; n22390_not
g29751 not n22354 ; n22354_not
g29752 not n13390 ; n13390_not
g29753 not n13426 ; n13426_not
g29754 not n13435 ; n13435_not
g29755 not n22318 ; n22318_not
g29756 not n13471 ; n13471_not
g29757 not n14083 ; n14083_not
g29758 not n22282 ; n22282_not
g29759 not n22642 ; n22642_not
g29760 not n13039 ; n13039_not
g29761 not n13624 ; n13624_not
g29762 not n22606 ; n22606_not
g29763 not n13066 ; n13066_not
g29764 not n13075 ; n13075_not
g29765 not n13660 ; n13660_not
g29766 not n13138 ; n13138_not
g29767 not n13147 ; n13147_not
g29768 not n13732 ; n13732_not
g29769 not n13183 ; n13183_not
g29770 not n13174 ; n13174_not
g29771 not n21805 ; n21805_not
g29772 not n22534 ; n22534_not
g29773 not n13219 ; n13219_not
g29774 not n13804 ; n13804_not
g29775 not n13255 ; n13255_not
g29776 not n13246 ; n13246_not
g29777 not n13840 ; n13840_not
g29778 not n10708 ; n10708_not
g29779 not n10744 ; n10744_not
g29780 not n24262 ; n24262_not
g29781 not n10267 ; n10267_not
g29782 not n10258 ; n10258_not
g29783 not n10780 ; n10780_not
g29784 not n10861 ; n10861_not
g29785 not n10339 ; n10339_not
g29786 not n10933 ; n10933_not
g29787 not n11077 ; n11077_not
g29788 not n11149 ; n11149_not
g29789 not n11185 ; n11185_not
g29790 not n11257 ; n11257_not
g29791 not n23281 ; n23281_not
g29792 not n11293 ; n11293_not
g29793 not n11347 ; n11347_not
g29794 not n11329 ; n11329_not
g29795 not n11356 ; n11356_not
g29796 not n10834 ; n10834_not
g29797 not n24802 ; n24802_not
g29798 not n24730 ; n24730_not
g29799 not n24631 ; n24631_not
g29800 not n24442 ; n24442_not
g29801 not n24424 ; n24424_not
g29802 not n24343 ; n24343_not
g29803 not n24325 ; n24325_not
g29804 not n10384 ; n10384_not
g29805 not n10456 ; n10456_not
g29806 not n10492 ; n10492_not
g29807 not n10528 ; n10528_not
g29808 not n10564 ; n10564_not
g29809 not n10078 ; n10078_not
g29810 not n10087 ; n10087_not
g29811 not n10636 ; n10636_not
g29812 not n10159 ; n10159_not
g29813 not n10672 ; n10672_not
g29814 not n10195 ; n10195_not
g29815 not n10186 ; n10186_not
g29816 not n11527 ; n11527_not
g29817 not n11518 ; n11518_not
g29818 not n12076 ; n12076_not
g29819 not n11554 ; n11554_not
g29820 not n11563 ; n11563_not
g29821 not n23452 ; n23452_not
g29822 not n11590 ; n11590_not
g29823 not n12148 ; n12148_not
g29824 not n11626 ; n11626_not
g29825 not n11635 ; n11635_not
g29826 not n12184 ; n12184_not
g29827 not n23416 ; n23416_not
g29828 not n11671 ; n11671_not
g29829 not n11662 ; n11662_not
g29830 not n11707 ; n11707_not
g29831 not n12256 ; n12256_not
g29832 not n23380 ; n23380_not
g29833 not n11743 ; n11743_not
g29834 not n11734 ; n11734_not
g29835 not n23920 ; n23920_not
g29836 not n11068 ; n11068_not
g29837 not n23812 ; n23812_not
g29838 not n11860 ; n11860_not
g29839 not n23740 ; n23740_not
g29840 not n23704 ; n23704_not
g29841 not n23632 ; n23632_not
g29842 not n11383 ; n11383_not
g29843 not n11374 ; n11374_not
g29844 not n11932 ; n11932_not
g29845 not n11419 ; n11419_not
g29846 not n23560 ; n23560_not
g29847 not n23524 ; n23524_not
g29848 not n11455 ; n11455_not
g29849 not n11446 ; n11446_not
g29850 not n11482 ; n11482_not
g29851 not n11491 ; n11491_not
g29852 not n14245 ; n14245_not
g29853 not n21922 ; n21922_not
g29854 not n14209 ; n14209_not
g29855 not n21094 ; n21094_not
g29856 not n14425 ; n14425_not
g29857 not n22246 ; n22246_not
g29858 not n14173 ; n14173_not
g29859 not n14605 ; n14605_not
g29860 not n14461 ; n14461_not
g29861 not n14281 ; n14281_not
g29862 not n14353 ; n14353_not
g29863 not n22138 ; n22138_not
g29864 not n14137 ; n14137_not
g29865 not n14533 ; n14533_not
g29866 not n22174 ; n22174_not
g29867 not n22066 ; n22066_not
g29868 not n14317 ; n14317_not
g29869 not n21067 ; n21067_not
g29870 not n21814 ; n21814_not
g29871 not n20087 ; n20087_not
g29872 not n14318 ; n14318_not
g29873 not n23309 ; n23309_not
g29874 not n16271 ; n16271_not
g29875 not n16262 ; n16262_not
g29876 not n23327 ; n23327_not
g29877 not n16190 ; n16190_not
g29878 not n22652 ; n22652_not
g29879 not n22571 ; n22571_not
g29880 not n14912 ; n14912_not
g29881 not n22643 ; n22643_not
g29882 not n20816 ; n20816_not
g29883 not n11870 ; n11870_not
g29884 not n16307 ; n16307_not
g29885 not n23264 ; n23264_not
g29886 not n23255 ; n23255_not
g29887 not n14642 ; n14642_not
g29888 not n10088 ; n10088_not
g29889 not n24047 ; n24047_not
g29890 not n16343 ; n16343_not
g29891 not n14327 ; n14327_not
g29892 not n23381 ; n23381_not
g29893 not n22616 ; n22616_not
g29894 not n11348 ; n11348_not
g29895 not n20744 ; n20744_not
g29896 not n10808 ; n10808_not
g29897 not n12293 ; n12293_not
g29898 not n11294 ; n11294_not
g29899 not n16226 ; n16226_not
g29900 not n16235 ; n16235_not
g29901 not n21356 ; n21356_not
g29902 not n23345 ; n23345_not
g29903 not n12329 ; n12329_not
g29904 not n21347 ; n21347_not
g29905 not n15056 ; n15056_not
g29906 not n21167 ; n21167_not
g29907 not n12365 ; n12365_not
g29908 not n12257 ; n12257_not
g29909 not n14462 ; n14462_not
g29910 not n20780 ; n20780_not
g29911 not n20078 ; n20078_not
g29912 not n17072 ; n17072_not
g29913 not n16442 ; n16442_not
g29914 not n16451 ; n16451_not
g29915 not n17441 ; n17441_not
g29916 not n10385 ; n10385_not
g29917 not n19313 ; n19313_not
g29918 not n16460 ; n16460_not
g29919 not n20960 ; n20960_not
g29920 not n20267 ; n20267_not
g29921 not n21851 ; n21851_not
g29922 not n20258 ; n20258_not
g29923 not n22391 ; n22391_not
g29924 not n14840 ; n14840_not
g29925 not n20294 ; n20294_not
g29926 not n22355 ; n22355_not
g29927 not n22364 ; n22364_not
g29928 not n18413 ; n18413_not
g29929 not n17621 ; n17621_not
g29930 not n12941 ; n12941_not
g29931 not n19241 ; n19241_not
g29932 not n12950 ; n12950_not
g29933 not n21419 ; n21419_not
g29934 not n12932 ; n12932_not
g29935 not n22328 ; n22328_not
g29936 not n22319 ; n22319_not
g29937 not n20339 ; n20339_not
g29938 not n16334 ; n16334_not
g29939 not n22535 ; n22535_not
g29940 not n20852 ; n20852_not
g29941 not n10196 ; n10196_not
g29942 not n19601 ; n19601_not
g29943 not n20159 ; n20159_not
g29944 not n10268 ; n10268_not
g29945 not n15092 ; n15092_not
g29946 not n21392 ; n21392_not
g29947 not n16370 ; n16370_not
g29948 not n22508 ; n22508_not
g29949 not n14507 ; n14507_not
g29950 not n22472 ; n22472_not
g29951 not n21383 ; n21383_not
g29952 not n22463 ; n22463_not
g29953 not n20195 ; n20195_not
g29954 not n20186 ; n20186_not
g29955 not n17036 ; n17036_not
g29956 not n19421 ; n19421_not
g29957 not n24461 ; n24461_not
g29958 not n16415 ; n16415_not
g29959 not n16406 ; n16406_not
g29960 not n10349 ; n10349_not
g29961 not n20924 ; n20924_not
g29962 not n22427 ; n22427_not
g29963 not n22436 ; n22436_not
g29964 not n16532 ; n16532_not
g29965 not n22931 ; n22931_not
g29966 not n11672 ; n11672_not
g29967 not n14363 ; n14363_not
g29968 not n23075 ; n23075_not
g29969 not n16055 ; n16055_not
g29970 not n22940 ; n22940_not
g29971 not n16046 ; n16046_not
g29972 not n11636 ; n11636_not
g29973 not n22904 ; n22904_not
g29974 not n24326 ; n24326_not
g29975 not n14354 ; n14354_not
g29976 not n11078 ; n11078_not
g29977 not n11087 ; n11087_not
g29978 not n23633 ; n23633_not
g29979 not n11933 ; n11933_not
g29980 not n11564 ; n11564_not
g29981 not n22832 ; n22832_not
g29982 not n16712 ; n16712_not
g29983 not n22823 ; n22823_not
g29984 not n20438 ; n20438_not
g29985 not n20456 ; n20456_not
g29986 not n16082 ; n16082_not
g29987 not n16091 ; n16091_not
g29988 not n23561 ; n23561_not
g29989 not n23813 ; n23813_not
g29990 not n11744 ; n11744_not
g29991 not n11780 ; n11780_not
g29992 not n23048 ; n23048_not
g29993 not n11258 ; n11258_not
g29994 not n16604 ; n16604_not
g29995 not n11267 ; n11267_not
g29996 not n23039 ; n23039_not
g29997 not n14660 ; n14660_not
g29998 not n16640 ; n16640_not
g29999 not n11816 ; n11816_not
g30000 not n11195 ; n11195_not
g30001 not n16019 ; n16019_not
g30002 not n14804 ; n14804_not
g30003 not n11186 ; n11186_not
g30004 not n11708 ; n11708_not
g30005 not n23741 ; n23741_not
g30006 not n17513 ; n17513_not
g30007 not n23705 ; n23705_not
g30008 not n11159 ; n11159_not
g30009 not n15902 ; n15902_not
g30010 not n15911 ; n15911_not
g30011 not n23084 ; n23084_not
g30012 not n21239 ; n21239_not
g30013 not n23183 ; n23183_not
g30014 not n11456 ; n11456_not
g30015 not n20564 ; n20564_not
g30016 not n23192 ; n23192_not
g30017 not n21275 ; n21275_not
g30018 not n23453 ; n23453_not
g30019 not n21284 ; n21284_not
g30020 not n12149 ; n12149_not
g30021 not n16154 ; n16154_not
g30022 not n16163 ; n16163_not
g30023 not n20636 ; n20636_not
g30024 not n10907 ; n10907_not
g30025 not n23228 ; n23228_not
g30026 not n23219 ; n23219_not
g30027 not n12185 ; n12185_not
g30028 not n10862 ; n10862_not
g30029 not n10871 ; n10871_not
g30030 not n11384 ; n11384_not
g30031 not n23417 ; n23417_not
g30032 not n14435 ; n14435_not
g30033 not n16820 ; n16820_not
g30034 not n20672 ; n20672_not
g30035 not n14426 ; n14426_not
g30036 not n20708 ; n20708_not
g30037 not n24407 ; n24407_not
g30038 not n24425 ; n24425_not
g30039 not n11528 ; n11528_not
g30040 not n23156 ; n23156_not
g30041 not n23147 ; n23147_not
g30042 not n10970 ; n10970_not
g30043 not n20465 ; n20465_not
g30044 not n11492 ; n11492_not
g30045 not n23921 ; n23921_not
g30046 not n23525 ; n23525_not
g30047 not n16127 ; n16127_not
g30048 not n22760 ; n22760_not
g30049 not n22751 ; n22751_not
g30050 not n16118 ; n16118_not
g30051 not n20492 ; n20492_not
g30052 not n10934 ; n10934_not
g30053 not n14390 ; n14390_not
g30054 not n21248 ; n21248_not
g30055 not n12077 ; n12077_not
g30056 not n20528 ; n20528_not
g30057 not n22715 ; n22715_not
g30058 not n22724 ; n22724_not
g30059 not n10943 ; n10943_not
g30060 not n14732 ; n14732_not
g30061 not n22580 ; n22580_not
g30062 not n10745 ; n10745_not
g30063 not n15533 ; n15533_not
g30064 not n17225 ; n17225_not
g30065 not n24614 ; n24614_not
g30066 not n13733 ; n13733_not
g30067 not n18404 ; n18404_not
g30068 not n19070 ; n19070_not
g30069 not n14147 ; n14147_not
g30070 not n19061 ; n19061_not
g30071 not n21815 ; n21815_not
g30072 not n21824 ; n21824_not
g30073 not n14219 ; n14219_not
g30074 not n19052 ; n19052_not
g30075 not n21464 ; n21464_not
g30076 not n24632 ; n24632_not
g30077 not n10709 ; n10709_not
g30078 not n14138 ; n14138_not
g30079 not n21455 ; n21455_not
g30080 not n13805 ; n13805_not
g30081 not n17261 ; n17261_not
g30082 not n15461 ; n15461_not
g30083 not n21743 ; n21743_not
g30084 not n21752 ; n21752_not
g30085 not n13472 ; n13472_not
g30086 not n13481 ; n13481_not
g30087 not n13490 ; n13490_not
g30088 not n19133 ; n19133_not
g30089 not n15641 ; n15641_not
g30090 not n18431 ; n18431_not
g30091 not n13535 ; n13535_not
g30092 not n13553 ; n13553_not
g30093 not n21923 ; n21923_not
g30094 not n21932 ; n21932_not
g30095 not n19115 ; n19115_not
g30096 not n17810 ; n17810_not
g30097 not n15605 ; n15605_not
g30098 not n10781 ; n10781_not
g30099 not n17405 ; n17405_not
g30100 not n13625 ; n13625_not
g30101 not n20483 ; n20483_not
g30102 not n15164 ; n15164_not
g30103 not n14282 ; n14282_not
g30104 not n14291 ; n14291_not
g30105 not n14570 ; n14570_not
g30106 not n13661 ; n13661_not
g30107 not n22607 ; n22607_not
g30108 not n24560 ; n24560_not
g30109 not n18134 ; n18134_not
g30110 not n21608 ; n21608_not
g30111 not n18143 ; n18143_not
g30112 not n18800 ; n18800_not
g30113 not n10529 ; n10529_not
g30114 not n17126 ; n17126_not
g30115 not n15317 ; n15317_not
g30116 not n17333 ; n17333_not
g30117 not n14174 ; n14174_not
g30118 not n21572 ; n21572_not
g30119 not n21563 ; n21563_not
g30120 not n15281 ; n15281_not
g30121 not n24803 ; n24803_not
g30122 not n18107 ; n18107_not
g30123 not n18062 ; n18062_not
g30124 not n18071 ; n18071_not
g30125 not n23336 ; n23336_not
g30126 not n14183 ; n14183_not
g30127 not n21527 ; n21527_not
g30128 not n10565 ; n10565_not
g30129 not n18035 ; n18035_not
g30130 not n21536 ; n21536_not
g30131 not n15263 ; n15263_not
g30132 not n18026 ; n18026_not
g30133 not n13517 ; n13517_not
g30134 not n14255 ; n14255_not
g30135 not n18350 ; n18350_not
g30136 not n14606 ; n14606_not
g30137 not n14615 ; n14615_not
g30138 not n13841 ; n13841_not
g30139 not n19016 ; n19016_not
g30140 not n18512 ; n18512_not
g30141 not n21716 ; n21716_not
g30142 not n21707 ; n21707_not
g30143 not n15425 ; n15425_not
g30144 not n18620 ; n18620_not
g30145 not n18323 ; n18323_not
g30146 not n21491 ; n21491_not
g30147 not n18314 ; n18314_not
g30148 not n10673 ; n10673_not
g30149 not n13913 ; n13913_not
g30150 not n10493 ; n10493_not
g30151 not n14246 ; n14246_not
g30152 not n18251 ; n18251_not
g30153 not n18242 ; n18242_not
g30154 not n21671 ; n21671_not
g30155 not n21680 ; n21680_not
g30156 not n18206 ; n18206_not
g30157 not n24713 ; n24713_not
g30158 not n24731 ; n24731_not
g30159 not n18215 ; n18215_not
g30160 not n10637 ; n10637_not
g30161 not n18170 ; n18170_not
g30162 not n21644 ; n21644_not
g30163 not n15353 ; n15353_not
g30164 not n21635 ; n21635_not
g30165 not n17153 ; n17153_not
g30166 not n12527 ; n12527_not
g30167 not n10835 ; n10835_not
g30168 not n12563 ; n12563_not
g30169 not n12554 ; n12554_not
g30170 not n12662 ; n12662_not
g30171 not n10457 ; n10457_not
g30172 not n19205 ; n19205_not
g30173 not n12842 ; n12842_not
g30174 not n22256 ; n22256_not
g30175 not n15821 ; n15821_not
g30176 not n21068 ; n21068_not
g30177 not n12851 ; n12851_not
g30178 not n12626 ; n12626_not
g30179 not n13148 ; n13148_not
g30180 not n12590 ; n12590_not
g30181 not n10817 ; n10817_not
g30182 not n15713 ; n15713_not
g30183 not n12743 ; n12743_not
g30184 not n12815 ; n12815_not
g30185 not n12806 ; n12806_not
g30186 not n22247 ; n22247_not
g30187 not n13364 ; n13364_not
g30188 not n22148 ; n22148_not
g30189 not n20366 ; n20366_not
g30190 not n22139 ; n22139_not
g30191 not n12770 ; n12770_not
g30192 not n10844 ; n10844_not
g30193 not n13328 ; n13328_not
g30194 not n12635 ; n12635_not
g30195 not n13184 ; n13184_not
g30196 not n12455 ; n12455_not
g30197 not n22283 ; n22283_not
g30198 not n22292 ; n22292_not
g30199 not n12491 ; n12491_not
g30200 not n12482 ; n12482_not
g30201 not n12446 ; n12446_not
g30202 not n21428 ; n21428_not
g30203 not n12707 ; n12707_not
g30204 not n22184 ; n22184_not
g30205 not n22076 ; n22076_not
g30206 not n18422 ; n18422_not
g30207 not n22175 ; n22175_not
g30208 not n13076 ; n13076_not
g30209 not n21860 ; n21860_not
g30210 not n12518 ; n12518_not
g30211 not n13292 ; n13292_not
g30212 not n13256 ; n13256_not
g30213 not n22067 ; n22067_not
g30214 not n14543 ; n14543_not
g30215 not n24308 ; n24308_not
g30216 not n12671 ; n12671_not
g30217 not n14534 ; n14534_not
g30218 not n13436 ; n13436_not
g30219 not n15128 ; n15128_not
g30220 not n12734 ; n12734_not
g30221 not n17073 ; n17073_not
g30222 not n10467 ; n10467_not
g30223 not n11529 ; n11529_not
g30224 not n19431 ; n19431_not
g30225 not n17109 ; n17109_not
g30226 not n11565 ; n11565_not
g30227 not n17127 ; n17127_not
g30228 not n18360 ; n18360_not
g30229 not n24309 ; n24309_not
g30230 not n10458 ; n10458_not
g30231 not n18423 ; n18423_not
g30232 not n23643 ; n23643_not
g30233 not n11745 ; n11745_not
g30234 not n16641 ; n16641_not
g30235 not n20196 ; n20196_not
g30236 not n23562 ; n23562_not
g30237 not n10395 ; n10395_not
g30238 not n19503 ; n19503_not
g30239 not n10386 ; n10386_not
g30240 not n24291 ; n24291_not
g30241 not n23571 ; n23571_not
g30242 not n18801 ; n18801_not
g30243 not n11709 ; n11709_not
g30244 not n24273 ; n24273_not
g30245 not n10908 ; n10908_not
g30246 not n21753 ; n21753_not
g30247 not n23634 ; n23634_not
g30248 not n23715 ; n23715_not
g30249 not n11673 ; n11673_not
g30250 not n10944 ; n10944_not
g30251 not n11637 ; n11637_not
g30252 not n10872 ; n10872_not
g30253 not n10359 ; n10359_not
g30254 not n23706 ; n23706_not
g30255 not n23850 ; n23850_not
g30256 not n16713 ; n16713_not
g30257 not n14058 ; n14058_not
g30258 not n11385 ; n11385_not
g30259 not n18252 ; n18252_not
g30260 not n14733 ; n14733_not
g30261 not n23355 ; n23355_not
g30262 not n11367 ; n11367_not
g30263 not n11196 ; n11196_not
g30264 not n19314 ; n19314_not
g30265 not n19323 ; n19323_not
g30266 not n23382 ; n23382_not
g30267 not n21717 ; n21717_not
g30268 not n10719 ; n10719_not
g30269 not n14805 ; n14805_not
g30270 not n23391 ; n23391_not
g30271 not n19800 ; n19800_not
g30272 not n10755 ; n10755_not
g30273 not n10782 ; n10782_not
g30274 not n18441 ; n18441_not
g30275 not n10836 ; n10836_not
g30276 not n18216 ; n18216_not
g30277 not n19206 ; n19206_not
g30278 not n19170 ; n19170_not
g30279 not n19215 ; n19215_not
g30280 not n23418 ; n23418_not
g30281 not n19143 ; n19143_not
g30282 not n19251 ; n19251_not
g30283 not n19242 ; n19242_not
g30284 not n10791 ; n10791_not
g30285 not n19134 ; n19134_not
g30286 not n23427 ; n23427_not
g30287 not n11268 ; n11268_not
g30288 not n10809 ; n10809_not
g30289 not n10746 ; n10746_not
g30290 not n17136 ; n17136_not
g30291 not n23490 ; n23490_not
g30292 not n17550 ; n17550_not
g30293 not n18324 ; n18324_not
g30294 not n21825 ; n21825_not
g30295 not n20088 ; n20088_not
g30296 not n10539 ; n10539_not
g30297 not n11493 ; n11493_not
g30298 not n10494 ; n10494_not
g30299 not n23922 ; n23922_not
g30300 not n23931 ; n23931_not
g30301 not n17037 ; n17037_not
g30302 not n19017 ; n19017_not
g30303 not n17703 ; n17703_not
g30304 not n10980 ; n10980_not
g30305 not n18621 ; n18621_not
g30306 not n19422 ; n19422_not
g30307 not n10674 ; n10674_not
g30308 not n10089 ; n10089_not
g30309 not n10683 ; n10683_not
g30310 not n17622 ; n17622_not
g30311 not n16821 ; n16821_not
g30312 not n10647 ; n10647_not
g30313 not n10638 ; n10638_not
g30314 not n19350 ; n19350_not
g30315 not n10197 ; n10197_not
g30316 not n11088 ; n11088_not
g30317 not n10269 ; n10269_not
g30318 not n10575 ; n10575_not
g30319 not n11457 ; n11457_not
g30320 not n10566 ; n10566_not
g30321 not n18513 ; n18513_not
g30322 not n14913 ; n14913_not
g30323 not n19053 ; n19053_not
g30324 not n12294 ; n12294_not
g30325 not n12852 ; n12852_not
g30326 not n12339 ; n12339_not
g30327 not n14364 ; n14364_not
g30328 not n12384 ; n12384_not
g30329 not n23085 ; n23085_not
g30330 not n12951 ; n12951_not
g30331 not n23049 ; n23049_not
g30332 not n13770 ; n13770_not
g30333 not n21069 ; n21069_not
g30334 not n13077 ; n13077_not
g30335 not n15822 ; n15822_not
g30336 not n15840 ; n15840_not
g30337 not n13149 ; n13149_not
g30338 not n23607 ; n23607_not
g30339 not n13185 ; n13185_not
g30340 not n22941 ; n22941_not
g30341 not n13257 ; n13257_not
g30342 not n17343 ; n17343_not
g30343 not n13293 ; n13293_not
g30344 not n22905 ; n22905_not
g30345 not n13329 ; n13329_not
g30346 not n17334 ; n17334_not
g30347 not n13365 ; n13365_not
g30348 not n22833 ; n22833_not
g30349 not n13437 ; n13437_not
g30350 not n23670 ; n23670_not
g30351 not n13473 ; n13473_not
g30352 not n22149 ; n22149_not
g30353 not n22761 ; n22761_not
g30354 not n11970 ; n11970_not
g30355 not n12528 ; n12528_not
g30356 not n12564 ; n12564_not
g30357 not n23229 ; n23229_not
g30358 not n15390 ; n15390_not
g30359 not n12078 ; n12078_not
g30360 not n12087 ; n12087_not
g30361 not n12636 ; n12636_not
g30362 not n12672 ; n12672_not
g30363 not n15363 ; n15363_not
g30364 not n15354 ; n15354_not
g30365 not n23193 ; n23193_not
g30366 not n12708 ; n12708_not
g30367 not n12195 ; n12195_not
g30368 not n20925 ; n20925_not
g30369 not n12186 ; n12186_not
g30370 not n12744 ; n12744_not
g30371 not n13806 ; n13806_not
g30372 not n15318 ; n15318_not
g30373 not n15327 ; n15327_not
g30374 not n23157 ; n23157_not
g30375 not n12780 ; n12780_not
g30376 not n24462 ; n24462_not
g30377 not n13815 ; n13815_not
g30378 not n20961 ; n20961_not
g30379 not n12267 ; n12267_not
g30380 not n12258 ; n12258_not
g30381 not n15912 ; n15912_not
g30382 not n15291 ; n15291_not
g30383 not n12816 ; n12816_not
g30384 not n15129 ; n15129_not
g30385 not n14256 ; n14256_not
g30386 not n13662 ; n13662_not
g30387 not n22437 ; n22437_not
g30388 not n13671 ; n13671_not
g30389 not n13284 ; n13284_not
g30390 not n17154 ; n17154_not
g30391 not n13635 ; n13635_not
g30392 not n17163 ; n17163_not
g30393 not n24714 ; n24714_not
g30394 not n21357 ; n21357_not
g30395 not n13626 ; n13626_not
g30396 not n14184 ; n14184_not
g30397 not n13590 ; n13590_not
g30398 not n22365 ; n22365_not
g30399 not n21393 ; n21393_not
g30400 not n22329 ; n22329_not
g30401 not n14148 ; n14148_not
g30402 not n24750 ; n24750_not
g30403 not n13563 ; n13563_not
g30404 not n13554 ; n13554_not
g30405 not n22293 ; n22293_not
g30406 not n21429 ; n21429_not
g30407 not n14076 ; n14076_not
g30408 not n14670 ; n14670_not
g30409 not n15282 ; n15282_not
g30410 not n22257 ; n22257_not
g30411 not n14085 ; n14085_not
g30412 not n17091 ; n17091_not
g30413 not n21465 ; n21465_not
g30414 not n14328 ; n14328_not
g30415 not n22725 ; n22725_not
g30416 not n24543 ; n24543_not
g30417 not n13734 ; n13734_not
g30418 not n17307 ; n17307_not
g30419 not n15165 ; n15165_not
g30420 not n22653 ; n22653_not
g30421 not n20466 ; n20466_not
g30422 not n17271 ; n17271_not
g30423 not n17262 ; n17262_not
g30424 not n13743 ; n13743_not
g30425 not n22617 ; n22617_not
g30426 not n24561 ; n24561_not
g30427 not n17226 ; n17226_not
g30428 not n21537 ; n21537_not
g30429 not n17235 ; n17235_not
g30430 not n23751 ; n23751_not
g30431 not n23742 ; n23742_not
g30432 not n22545 ; n22545_not
g30433 not n24615 ; n24615_not
g30434 not n21249 ; n21249_not
g30435 not n14292 ; n14292_not
g30436 not n13707 ; n13707_not
g30437 not n23823 ; n23823_not
g30438 not n23814 ; n23814_not
g30439 not n17190 ; n17190_not
g30440 not n21285 ; n21285_not
g30441 not n22509 ; n22509_not
g30442 not n22473 ; n22473_not
g30443 not n22185 ; n22185_not
g30444 not n17820 ; n17820_not
g30445 not n17442 ; n17442_not
g30446 not n16470 ; n16470_not
g30447 not n16461 ; n16461_not
g30448 not n17451 ; n17451_not
g30449 not n16452 ; n16452_not
g30450 not n15831 ; n15831_not
g30451 not n20493 ; n20493_not
g30452 not n18072 ; n18072_not
g30453 not n16416 ; n16416_not
g30454 not n14616 ; n14616_not
g30455 not n20529 ; n20529_not
g30456 not n17415 ; n17415_not
g30457 not n16380 ; n16380_not
g30458 not n15750 ; n15750_not
g30459 not n20565 ; n20565_not
g30460 not n14580 ; n14580_not
g30461 not n14544 ; n14544_not
g30462 not n20637 ; n20637_not
g30463 not n16344 ; n16344_not
g30464 not n15723 ; n15723_not
g30465 not n15714 ; n15714_not
g30466 not n13950 ; n13950_not
g30467 not n14508 ; n14508_not
g30468 not n17406 ; n17406_not
g30469 not n13923 ; n13923_not
g30470 not n20673 ; n20673_not
g30471 not n16308 ; n16308_not
g30472 not n20709 ; n20709_not
g30473 not n11781 ; n11781_not
g30474 not n19530 ; n19530_not
g30475 not n16605 ; n16605_not
g30476 not n11817 ; n11817_not
g30477 not n20268 ; n20268_not
g30478 not n23463 ; n23463_not
g30479 not n11844 ; n11844_not
g30480 not n18180 ; n18180_not
g30481 not n19611 ; n19611_not
g30482 not n19602 ; n19602_not
g30483 not n21681 ; n21681_not
g30484 not n17514 ; n17514_not
g30485 not n17523 ; n17523_not
g30486 not n11871 ; n11871_not
g30487 not n11853 ; n11853_not
g30488 not n16533 ; n16533_not
g30489 not n11880 ; n11880_not
g30490 not n20376 ; n20376_not
g30491 not n16515 ; n16515_not
g30492 not n23454 ; n23454_not
g30493 not n11349 ; n11349_not
g30494 not n19710 ; n19710_not
g30495 not n18144 ; n18144_not
g30496 not n24390 ; n24390_not
g30497 not n24408 ; n24408_not
g30498 not n21933 ; n21933_not
g30499 not n21645 ; n21645_not
g30500 not n18108 ; n18108_not
g30501 not n16056 ; n16056_not
g30502 not n20817 ; n20817_not
g30503 not n16164 ; n16164_not
g30504 not n15534 ; n15534_not
g30505 not n15543 ; n15543_not
g30506 not n14436 ; n14436_not
g30507 not n23328 ; n23328_not
g30508 not n13851 ; n13851_not
g30509 not n12393 ; n12393_not
g30510 not n23319 ; n23319_not
g30511 not n23265 ; n23265_not
g30512 not n16128 ; n16128_not
g30513 not n15507 ; n15507_not
g30514 not n21573 ; n21573_not
g30515 not n18036 ; n18036_not
g30516 not n13842 ; n13842_not
g30517 not n12492 ; n12492_not
g30518 not n11943 ; n11943_not
g30519 not n11907 ; n11907_not
g30520 not n12456 ; n12456_not
g30521 not n15093 ; n15093_not
g30522 not n16092 ; n16092_not
g30523 not n15462 ; n15462_not
g30524 not n15471 ; n15471_not
g30525 not n11934 ; n11934_not
g30526 not n17370 ; n17370_not
g30527 not n20853 ; n20853_not
g30528 not n24444 ; n24444_not
g30529 not n13914 ; n13914_not
g30530 not n14841 ; n14841_not
g30531 not n16272 ; n16272_not
g30532 not n15651 ; n15651_not
g30533 not n15642 ; n15642_not
g30534 not n14472 ; n14472_not
g30535 not n20745 ; n20745_not
g30536 not n15057 ; n15057_not
g30537 not n22608 ; n22608_not
g30538 not n16236 ; n16236_not
g30539 not n15606 ; n15606_not
g30540 not n15615 ; n15615_not
g30541 not n23535 ; n23535_not
g30542 not n23346 ; n23346_not
g30543 not n22077 ; n22077_not
g30544 not n20781 ; n20781_not
g30545 not n15426 ; n15426_not
g30546 not n21609 ; n21609_not
g30547 not n15570 ; n15570_not
g30548 not n23526 ; n23526_not
g30549 not n15435 ; n15435_not
g30550 not n11835 ; n11835_not
g30551 not n18325 ; n18325_not
g30552 not n17092 ; n17092_not
g30553 not n24445 ; n24445_not
g30554 not n24805 ; n24805_not
g30555 not n24751 ; n24751_not
g30556 not n24373 ; n24373_not
g30557 not n21079 ; n21079_not
g30558 not n18361 ; n18361_not
g30559 not n18442 ; n18442_not
g30560 not n18073 ; n18073_not
g30561 not n24526 ; n24526_not
g30562 not n24544 ; n24544_not
g30563 not n24292 ; n24292_not
g30564 not n24580 ; n24580_not
g30565 not n18217 ; n18217_not
g30566 not n24427 ; n24427_not
g30567 not n18109 ; n18109_not
g30568 not n18253 ; n18253_not
g30569 not n18145 ; n18145_not
g30570 not n24391 ; n24391_not
g30571 not n17821 ; n17821_not
g30572 not n18181 ; n18181_not
g30573 not n24733 ; n24733_not
g30574 not n21790 ; n21790_not
g30575 not n18037 ; n18037_not
g30576 not n21178 ; n21178_not
g30577 not n22654 ; n22654_not
g30578 not n22690 ; n22690_not
g30579 not n22726 ; n22726_not
g30580 not n22762 ; n22762_not
g30581 not n22834 ; n22834_not
g30582 not n22870 ; n22870_not
g30583 not n22906 ; n22906_not
g30584 not n22942 ; n22942_not
g30585 not n20368 ; n20368_not
g30586 not n23086 ; n23086_not
g30587 not n23158 ; n23158_not
g30588 not n23194 ; n23194_not
g30589 not n21574 ; n21574_not
g30590 not n23266 ; n23266_not
g30591 not n20863 ; n20863_not
g30592 not n22537 ; n22537_not
g30593 not n20854 ; n20854_not
g30594 not n22573 ; n22573_not
g30595 not n20890 ; n20890_not
g30596 not n23356 ; n23356_not
g30597 not n22078 ; n22078_not
g30598 not n23392 ; n23392_not
g30599 not n23428 ; n23428_not
g30600 not n23464 ; n23464_not
g30601 not n21970 ; n21970_not
g30602 not n21646 ; n21646_not
g30603 not n20935 ; n20935_not
g30604 not n20476 ; n20476_not
g30605 not n20926 ; n20926_not
g30606 not n20755 ; n20755_not
g30607 not n20746 ; n20746_not
g30608 not n21466 ; n21466_not
g30609 not n22258 ; n22258_not
g30610 not n22294 ; n22294_not
g30611 not n20719 ; n20719_not
g30612 not n20791 ; n20791_not
g30613 not n20782 ; n20782_not
g30614 not n22366 ; n22366_not
g30615 not n20683 ; n20683_not
g30616 not n20674 ; n20674_not
g30617 not n21394 ; n21394_not
g30618 not n20638 ; n20638_not
g30619 not n20647 ; n20647_not
g30620 not n21358 ; n21358_not
g30621 not n22438 ; n22438_not
g30622 not n22474 ; n22474_not
g30623 not n20566 ; n20566_not
g30624 not n20575 ; n20575_not
g30625 not n21286 ; n21286_not
g30626 not n22186 ; n22186_not
g30627 not n22546 ; n22546_not
g30628 not n20539 ; n20539_not
g30629 not n21538 ; n21538_not
g30630 not n20818 ; n20818_not
g30631 not n21853 ; n21853_not
g30632 not n20827 ; n20827_not
g30633 not n22591 ; n22591_not
g30634 not n20494 ; n20494_not
g30635 not n22618 ; n22618_not
g30636 not n19540 ; n19540_not
g30637 not n19504 ; n19504_not
g30638 not n18811 ; n18811_not
g30639 not n18802 ; n18802_not
g30640 not n19432 ; n19432_not
g30641 not n18730 ; n18730_not
g30642 not n18703 ; n18703_not
g30643 not n19360 ; n19360_not
g30644 not n19324 ; n19324_not
g30645 not n18622 ; n18622_not
g30646 not n18631 ; n18631_not
g30647 not n19252 ; n19252_not
g30648 not n18550 ; n18550_not
g30649 not n19216 ; n19216_not
g30650 not n18523 ; n18523_not
g30651 not n18514 ; n18514_not
g30652 not n19180 ; n19180_not
g30653 not n19144 ; n19144_not
g30654 not n18451 ; n18451_not
g30655 not n23347 ; n23347_not
g30656 not n19072 ; n19072_not
g30657 not n19090 ; n19090_not
g30658 not n19081 ; n19081_not
g30659 not n24049 ; n24049_not
g30660 not n24265 ; n24265_not
g30661 not n24274 ; n24274_not
g30662 not n21826 ; n21826_not
g30663 not n21754 ; n21754_not
g30664 not n23536 ; n23536_not
g30665 not n20449 ; n20449_not
g30666 not n20467 ; n20467_not
g30667 not n23572 ; n23572_not
g30668 not n23608 ; n23608_not
g30669 not n21682 ; n21682_not
g30670 not n20962 ; n20962_not
g30671 not n23644 ; n23644_not
g30672 not n23680 ; n23680_not
g30673 not n20377 ; n20377_not
g30674 not n20971 ; n20971_not
g30675 not n23716 ; n23716_not
g30676 not n21934 ; n21934_not
g30677 not n23752 ; n23752_not
g30678 not n20269 ; n20269_not
g30679 not n20197 ; n20197_not
g30680 not n23824 ; n23824_not
g30681 not n23860 ; n23860_not
g30682 not n23932 ; n23932_not
g30683 not n20089 ; n20089_not
g30684 not n21718 ; n21718_not
g30685 not n21169 ; n21169_not
g30686 not n19801 ; n19801_not
g30687 not n19720 ; n19720_not
g30688 not n19027 ; n19027_not
g30689 not n19018 ; n19018_not
g30690 not n21871 ; n21871_not
g30691 not n19612 ; n19612_not
g30692 not n18910 ; n18910_not
g30693 not n14680 ; n14680_not
g30694 not n13672 ; n13672_not
g30695 not n12709 ; n12709_not
g30696 not n17272 ; n17272_not
g30697 not n13078 ; n13078_not
g30698 not n14086 ; n14086_not
g30699 not n11872 ; n11872_not
g30700 not n13087 ; n13087_not
g30701 not n12745 ; n12745_not
g30702 not n14950 ; n14950_not
g30703 not n15544 ; n15544_not
g30704 not n17524 ; n17524_not
g30705 not n14914 ; n14914_not
g30706 not n14923 ; n14923_not
g30707 not n12781 ; n12781_not
g30708 not n15508 ; n15508_not
g30709 not n12817 ; n12817_not
g30710 not n16615 ; n16615_not
g30711 not n10909 ; n10909_not
g30712 not n15472 ; n15472_not
g30713 not n16237 ; n16237_not
g30714 not n12853 ; n12853_not
g30715 not n17074 ; n17074_not
g30716 not n13636 ; n13636_not
g30717 not n16606 ; n16606_not
g30718 not n14842 ; n14842_not
g30719 not n10981 ; n10981_not
g30720 not n14545 ; n14545_not
g30721 not n12529 ; n12529_not
g30722 not n11386 ; n11386_not
g30723 not n11908 ; n11908_not
g30724 not n15058 ; n15058_not
g30725 not n15067 ; n15067_not
g30726 not n14581 ; n14581_not
g30727 not n15652 ; n15652_not
g30728 not n16930 ; n16930_not
g30729 not n16129 ; n16129_not
g30730 not n13708 ; n13708_not
g30731 not n12565 ; n12565_not
g30732 not n15616 ; n15616_not
g30733 not n16165 ; n16165_not
g30734 not n14617 ; n14617_not
g30735 not n12637 ; n12637_not
g30736 not n17380 ; n17380_not
g30737 not n17560 ; n17560_not
g30738 not n14644 ; n14644_not
g30739 not n12673 ; n12673_not
g30740 not n14671 ; n14671_not
g30741 not n16903 ; n16903_not
g30742 not n14653 ; n14653_not
g30743 not n15580 ; n15580_not
g30744 not n10945 ; n10945_not
g30745 not n10099 ; n10099_not
g30746 not n16570 ; n16570_not
g30747 not n14707 ; n14707_not
g30748 not n12970 ; n12970_not
g30749 not n10855 ; n10855_not
g30750 not n16309 ; n16309_not
g30751 not n10648 ; n10648_not
g30752 not n10684 ; n10684_not
g30753 not n16381 ; n16381_not
g30754 not n14464 ; n14464_not
g30755 not n15292 ; n15292_not
g30756 not n10792 ; n10792_not
g30757 not n15265 ; n15265_not
g30758 not n16345 ; n16345_not
g30759 not n15238 ; n15238_not
g30760 not n17164 ; n17164_not
g30761 not n10198 ; n10198_not
g30762 not n16534 ; n16534_not
g30763 not n10756 ; n10756_not
g30764 not n16543 ; n16543_not
g30765 not n14635 ; n14635_not
g30766 not n17416 ; n17416_not
g30767 not n10279 ; n10279_not
g30768 not n15256 ; n15256_not
g30769 not n11845 ; n11845_not
g30770 not n14851 ; n14851_not
g30771 not n11818 ; n11818_not
g30772 not n10396 ; n10396_not
g30773 not n15436 ; n15436_not
g30774 not n11836 ; n11836_not
g30775 not n10468 ; n10468_not
g30776 not n14815 ; n14815_not
g30777 not n14806 ; n14806_not
g30778 not n13492 ; n13492_not
g30779 not n16831 ; n16831_not
g30780 not n14770 ; n14770_not
g30781 not n10576 ; n10576_not
g30782 not n16822 ; n16822_not
g30783 not n16453 ; n16453_not
g30784 not n16273 ; n16273_not
g30785 not n17236 ; n17236_not
g30786 not n15364 ; n15364_not
g30787 not n13564 ; n13564_not
g30788 not n16750 ; n16750_not
g30789 not n10873 ; n10873_not
g30790 not n17452 ; n17452_not
g30791 not n14743 ; n14743_not
g30792 not n14734 ; n14734_not
g30793 not n15328 ; n15328_not
g30794 not n16417 ; n16417_not
g30795 not n17128 ; n17128_not
g30796 not n11638 ; n11638_not
g30797 not n17704 ; n17704_not
g30798 not n13186 ; n13186_not
g30799 not n13447 ; n13447_not
g30800 not n11647 ; n11647_not
g30801 not n13438 ; n13438_not
g30802 not n17047 ; n17047_not
g30803 not n17038 ; n17038_not
g30804 not n11782 ; n11782_not
g30805 not n11827 ; n11827_not
g30806 not n17344 ; n17344_not
g30807 not n13519 ; n13519_not
g30808 not n14149 ; n14149_not
g30809 not n11566 ; n11566_not
g30810 not n14185 ; n14185_not
g30811 not n13744 ; n13744_not
g30812 not n12457 ; n12457_not
g30813 not n11575 ; n11575_not
g30814 not n12088 ; n12088_not
g30815 not n14257 ; n14257_not
g30816 not n11539 ; n11539_not
g30817 not n15913 ; n15913_not
g30818 not n11269 ; n11269_not
g30819 not n15283 ; n15283_not
g30820 not n12268 ; n12268_not
g30821 not n13816 ; n13816_not
g30822 not n13258 ; n13258_not
g30823 not n13267 ; n13267_not
g30824 not n11719 ; n11719_not
g30825 not n17308 ; n17308_not
g30826 not n17083 ; n17083_not
g30827 not n13852 ; n13852_not
g30828 not n13294 ; n13294_not
g30829 not n11683 ; n11683_not
g30830 not n11674 ; n11674_not
g30831 not n12196 ; n12196_not
g30832 not n13339 ; n13339_not
g30833 not n13924 ; n13924_not
g30834 not n11197 ; n11197_not
g30835 not n11746 ; n11746_not
g30836 not n13375 ; n13375_not
g30837 not n13366 ; n13366_not
g30838 not n13780 ; n13780_not
g30839 not n11755 ; n11755_not
g30840 not n13960 ; n13960_not
g30841 not n11791 ; n11791_not
g30842 not n10837 ; n10837_not
g30843 not n13195 ; n13195_not
g30844 not n14365 ; n14365_not
g30845 not n13159 ; n13159_not
g30846 not n11980 ; n11980_not
g30847 not n14473 ; n14473_not
g30848 not n16723 ; n16723_not
g30849 not n11944 ; n11944_not
g30850 not n16057 ; n16057_not
g30851 not n11089 ; n11089_not
g30852 not n16714 ; n16714_not
g30853 not n16651 ; n16651_not
g30854 not n14437 ; n14437_not
g30855 not n15760 ; n15760_not
g30856 not n12493 ; n12493_not
g30857 not n15166 ; n15166_not
g30858 not n15175 ; n15175_not
g30859 not n16093 ; n16093_not
g30860 not n16642 ; n16642_not
g30861 not n17632 ; n17632_not
g30862 not n14509 ; n14509_not
g30863 not n15850 ; n15850_not
g30864 not n15094 ; n15094_not
g30865 not n15841 ; n15841_not
g30866 not n15724 ; n15724_not
g30867 not n14293 ; n14293_not
g30868 not n11494 ; n11494_not
g30869 not n11395 ; n11395_not
g30870 not n11467 ; n11467_not
g30871 not n14329 ; n14329_not
g30872 not n15832 ; n15832_not
g30873 not n15139 ; n15139_not
g30874 not n11458 ; n11458_not
g30875 not n18155 ; n18155_not
g30876 not n23195 ; n23195_not
g30877 not n10919 ; n10919_not
g30878 not n18146 ; n18146_not
g30879 not n12647 ; n12647_not
g30880 not n12638 ; n12638_not
g30881 not n18263 ; n18263_not
g30882 not n11099 ; n11099_not
g30883 not n12575 ; n12575_not
g30884 not n18920 ; n18920_not
g30885 not n23267 ; n23267_not
g30886 not n20648 ; n20648_not
g30887 not n18254 ; n18254_not
g30888 not n20684 ; n20684_not
g30889 not n18812 ; n18812_not
g30890 not n13196 ; n13196_not
g30891 not n11576 ; n11576_not
g30892 not n19091 ; n19091_not
g30893 not n23276 ; n23276_not
g30894 not n20828 ; n20828_not
g30895 not n22259 ; n22259_not
g30896 not n22268 ; n22268_not
g30897 not n18362 ; n18362_not
g30898 not n22196 ; n22196_not
g30899 not n20792 ; n20792_not
g30900 not n18191 ; n18191_not
g30901 not n18182 ; n18182_not
g30902 not n19028 ; n19028_not
g30903 not n22187 ; n22187_not
g30904 not n17309 ; n17309_not
g30905 not n10991 ; n10991_not
g30906 not n12674 ; n12674_not
g30907 not n20864 ; n20864_not
g30908 not n11396 ; n11396_not
g30909 not n20756 ; n20756_not
g30910 not n17273 ; n17273_not
g30911 not n12683 ; n12683_not
g30912 not n18335 ; n18335_not
g30913 not n18326 ; n18326_not
g30914 not n11468 ; n11468_not
g30915 not n18227 ; n18227_not
g30916 not n18218 ; n18218_not
g30917 not n10946 ; n10946_not
g30918 not n20936 ; n20936_not
g30919 not n10955 ; n10955_not
g30920 not n13268 ; n13268_not
g30921 not n23933 ; n23933_not
g30922 not n18290 ; n18290_not
g30923 not n17237 ; n17237_not
g30924 not n20099 ; n20099_not
g30925 not n10982 ; n10982_not
g30926 not n23168 ; n23168_not
g30927 not n23159 ; n23159_not
g30928 not n18371 ; n18371_not
g30929 not n10883 ; n10883_not
g30930 not n20198 ; n20198_not
g30931 not n10874 ; n10874_not
g30932 not n22547 ; n22547_not
g30933 not n22556 ; n22556_not
g30934 not n16139 ; n16139_not
g30935 not n16760 ; n16760_not
g30936 not n19613 ; n19613_not
g30937 not n16346 ; n16346_not
g30938 not n22808 ; n22808_not
g30939 not n16355 ; n16355_not
g30940 not n23573 ; n23573_not
g30941 not n16094 ; n16094_not
g30942 not n16724 ; n16724_not
g30943 not n11945 ; n11945_not
g30944 not n22844 ; n22844_not
g30945 not n22835 ; n22835_not
g30946 not n16067 ; n16067_not
g30947 not n23609 ; n23609_not
g30948 not n16058 ; n16058_not
g30949 not n19541 ; n19541_not
g30950 not n11909 ; n11909_not
g30951 not n22871 ; n22871_not
g30952 not n22880 ; n22880_not
g30953 not n23645 ; n23645_not
g30954 not n16652 ; n16652_not
g30955 not n19505 ; n19505_not
g30956 not n16616 ; n16616_not
g30957 not n11891 ; n11891_not
g30958 not n15950 ; n15950_not
g30959 not n22916 ; n22916_not
g30960 not n22907 ; n22907_not
g30961 not n22475 ; n22475_not
g30962 not n23681 ; n23681_not
g30963 not n22484 ; n22484_not
g30964 not n23393 ; n23393_not
g30965 not n16283 ; n16283_not
g30966 not n16274 ; n16274_not
g30967 not n12269 ; n12269_not
g30968 not n16904 ; n16904_not
g30969 not n22619 ; n22619_not
g30970 not n22628 ; n22628_not
g30971 not n22655 ; n22655_not
g30972 not n22664 ; n22664_not
g30973 not n23429 ; n23429_not
g30974 not n12197 ; n12197_not
g30975 not n23357 ; n23357_not
g30976 not n22592 ; n22592_not
g30977 not n16238 ; n16238_not
g30978 not n16247 ; n16247_not
g30979 not n22691 ; n22691_not
g30980 not n23465 ; n23465_not
g30981 not n16940 ; n16940_not
g30982 not n11873 ; n11873_not
g30983 not n19721 ; n19721_not
g30984 not n16319 ; n16319_not
g30985 not n12089 ; n12089_not
g30986 not n16832 ; n16832_not
g30987 not n22727 ; n22727_not
g30988 not n22736 ; n22736_not
g30989 not n22565 ; n22565_not
g30990 not n16166 ; n16166_not
g30991 not n16175 ; n16175_not
g30992 not n22772 ; n22772_not
g30993 not n22763 ; n22763_not
g30994 not n11981 ; n11981_not
g30995 not n23537 ; n23537_not
g30996 not n12926 ; n12926_not
g30997 not n11756 ; n11756_not
g30998 not n12944 ; n12944_not
g30999 not n11198 ; n11198_not
g31000 not n23825 ; n23825_not
g31001 not n19217 ; n19217_not
g31002 not n16472 ; n16472_not
g31003 not n19811 ; n19811_not
g31004 not n19802 ; n19802_not
g31005 not n11684 ; n11684_not
g31006 not n12953 ; n12953_not
g31007 not n19181 ; n19181_not
g31008 not n11648 ; n11648_not
g31009 not n12980 ; n12980_not
g31010 not n23087 ; n23087_not
g31011 not n23096 ; n23096_not
g31012 not n22295 ; n22295_not
g31013 not n17147 ; n17147_not
g31014 not n20576 ; n20576_not
g31015 not n12467 ; n12467_not
g31016 not n19145 ; n19145_not
g31017 not n23861 ; n23861_not
g31018 not n12458 ; n12458_not
g31019 not n18443 ; n18443_not
g31020 not n17165 ; n17165_not
g31021 not n12494 ; n12494_not
g31022 not n13088 ; n13088_not
g31023 not n19109 ; n19109_not
g31024 not n19910 ; n19910_not
g31025 not n12539 ; n12539_not
g31026 not n12566 ; n12566_not
g31027 not n16580 ; n16580_not
g31028 not n16391 ; n16391_not
g31029 not n19433 ; n19433_not
g31030 not n16382 ; n16382_not
g31031 not n15923 ; n15923_not
g31032 not n15914 ; n15914_not
g31033 not n16544 ; n16544_not
g31034 not n22943 ; n22943_not
g31035 not n22448 ; n22448_not
g31036 not n22952 ; n22952_not
g31037 not n22439 ; n22439_not
g31038 not n23717 ; n23717_not
g31039 not n17048 ; n17048_not
g31040 not n16418 ; n16418_not
g31041 not n19361 ; n19361_not
g31042 not n19253 ; n19253_not
g31043 not n20468 ; n20468_not
g31044 not n11792 ; n11792_not
g31045 not n22367 ; n22367_not
g31046 not n11279 ; n11279_not
g31047 not n22376 ; n22376_not
g31048 not n11828 ; n11828_not
g31049 not n16481 ; n16481_not
g31050 not n17093 ; n17093_not
g31051 not n11837 ; n11837_not
g31052 not n17084 ; n17084_not
g31053 not n19325 ; n19325_not
g31054 not n16490 ; n16490_not
g31055 not n16427 ; n16427_not
g31056 not n11846 ; n11846_not
g31057 not n23753 ; n23753_not
g31058 not n21908 ; n21908_not
g31059 not n14924 ; n14924_not
g31060 not n17624 ; n17624_not
g31061 not n14294 ; n14294_not
g31062 not n10577 ; n10577_not
g31063 not n13637 ; n13637_not
g31064 not n14258 ; n14258_not
g31065 not n10469 ; n10469_not
g31066 not n10397 ; n10397_not
g31067 not n14267 ; n14267_not
g31068 not n14852 ; n14852_not
g31069 not n14816 ; n14816_not
g31070 not n14186 ; n14186_not
g31071 not n14195 ; n14195_not
g31072 not n14780 ; n14780_not
g31073 not n14159 ; n14159_not
g31074 not n14744 ; n14744_not
g31075 not n24356 ; n24356_not
g31076 not n14708 ; n14708_not
g31077 not n21845 ; n21845_not
g31078 not n21827 ; n21827_not
g31079 not n21854 ; n21854_not
g31080 not n17525 ; n17525_not
g31081 not n24374 ; n24374_not
g31082 not n21872 ; n21872_not
g31083 not n21863 ; n21863_not
g31084 not n13673 ; n13673_not
g31085 not n21881 ; n21881_not
g31086 not n18416 ; n18416_not
g31087 not n10757 ; n10757_not
g31088 not n14636 ; n14636_not
g31089 not n14618 ; n14618_not
g31090 not n14627 ; n14627_not
g31091 not n14591 ; n14591_not
g31092 not n14582 ; n14582_not
g31093 not n15176 ; n15176_not
g31094 not n12971 ; n12971_not
g31095 not n14546 ; n14546_not
g31096 not n14555 ; n14555_not
g31097 not n14519 ; n14519_not
g31098 not n14474 ; n14474_not
g31099 not n21944 ; n21944_not
g31100 not n14483 ; n14483_not
g31101 not n21935 ; n21935_not
g31102 not n17453 ; n17453_not
g31103 not n10685 ; n10685_not
g31104 not n15068 ; n15068_not
g31105 not n14447 ; n14447_not
g31106 not n10649 ; n10649_not
g31107 not n14438 ; n14438_not
g31108 not n13565 ; n13565_not
g31109 not n14375 ; n14375_not
g31110 not n24275 ; n24275_not
g31111 not n14366 ; n14366_not
g31112 not n14960 ; n14960_not
g31113 not n14339 ; n14339_not
g31114 not n14096 ; n14096_not
g31115 not n14069 ; n14069_not
g31116 not n24662 ; n24662_not
g31117 not n14087 ; n14087_not
g31118 not n21539 ; n21539_not
g31119 not n21548 ; n21548_not
g31120 not n21584 ; n21584_not
g31121 not n21575 ; n21575_not
g31122 not n17705 ; n17705_not
g31123 not n24680 ; n24680_not
g31124 not n17129 ; n17129_not
g31125 not n21791 ; n21791_not
g31126 not n13781 ; n13781_not
g31127 not n24716 ; n24716_not
g31128 not n13961 ; n13961_not
g31129 not n21656 ; n21656_not
g31130 not n21647 ; n21647_not
g31131 not n13925 ; n13925_not
g31132 not n24734 ; n24734_not
g31133 not n21683 ; n21683_not
g31134 not n21692 ; n21692_not
g31135 not n21728 ; n21728_not
g31136 not n21719 ; n21719_not
g31137 not n13853 ; n13853_not
g31138 not n13817 ; n13817_not
g31139 not n21755 ; n21755_not
g31140 not n21764 ; n21764_not
g31141 not n24806 ; n24806_not
g31142 not n24428 ; n24428_not
g31143 not n14672 ; n14672_not
g31144 not n21188 ; n21188_not
g31145 not n17561 ; n17561_not
g31146 not n14645 ; n14645_not
g31147 not n22583 ; n22583_not
g31148 not n13709 ; n13709_not
g31149 not n22574 ; n22574_not
g31150 not n21296 ; n21296_not
g31151 not n21287 ; n21287_not
g31152 not n24509 ; n24509_not
g31153 not n17633 ; n17633_not
g31154 not n24527 ; n24527_not
g31155 not n21836 ; n21836_not
g31156 not n21368 ; n21368_not
g31157 not n21359 ; n21359_not
g31158 not n24563 ; n24563_not
g31159 not n21395 ; n21395_not
g31160 not n24581 ; n24581_not
g31161 not n13745 ; n13745_not
g31162 not n21467 ; n21467_not
g31163 not n21476 ; n21476_not
g31164 not n15725 ; n15725_not
g31165 not n12854 ; n12854_not
g31166 not n12863 ; n12863_not
g31167 not n18632 ; n18632_not
g31168 not n15653 ; n15653_not
g31169 not n15617 ; n15617_not
g31170 not n22088 ; n22088_not
g31171 not n21179 ; n21179_not
g31172 not n22079 ; n22079_not
g31173 not n17930 ; n17930_not
g31174 not n13448 ; n13448_not
g31175 not n15581 ; n15581_not
g31176 not n12890 ; n12890_not
g31177 not n15545 ; n15545_not
g31178 not n17903 ; n17903_not
g31179 not n18560 ; n18560_not
g31180 not n15509 ; n15509_not
g31181 not n15473 ; n15473_not
g31182 not n18524 ; n18524_not
g31183 not n15437 ; n15437_not
g31184 not n17345 ; n17345_not
g31185 not n18119 ; n18119_not
g31186 not n12755 ; n12755_not
g31187 not n20972 ; n20972_not
g31188 not n12746 ; n12746_not
g31189 not n20279 ; n20279_not
g31190 not n15266 ; n15266_not
g31191 not n12782 ; n12782_not
g31192 not n12791 ; n12791_not
g31193 not n18083 ; n18083_not
g31194 not n18074 ; n18074_not
g31195 not n18740 ; n18740_not
g31196 not n13376 ; n13376_not
g31197 not n18038 ; n18038_not
g31198 not n18047 ; n18047_not
g31199 not n18704 ; n18704_not
g31200 not n15833 ; n15833_not
g31201 not n20387 ; n20387_not
g31202 not n20378 ; n20378_not
g31203 not n12827 ; n12827_not
g31204 not n12818 ; n12818_not
g31205 not n17381 ; n17381_not
g31206 not n15761 ; n15761_not
g31207 not n15365 ; n15365_not
g31208 not n17417 ; n17417_not
g31209 not n15293 ; n15293_not
g31210 not n18425 ; n18425_not
g31211 not n15329 ; n15329_not
g31212 not n10793 ; n10793_not
g31213 not n17831 ; n17831_not
g31214 not n17822 ; n17822_not
g31215 not n21971 ; n21971_not
g31216 not n13529 ; n13529_not
g31217 not n18452 ; n18452_not
g31218 not n21980 ; n21980_not
g31219 not n13818 ; n13818_not
g31220 not n12468 ; n12468_not
g31221 not n13197 ; n13197_not
g31222 not n14376 ; n14376_not
g31223 not n13782 ; n13782_not
g31224 not n13791 ; n13791_not
g31225 not n19362 ; n19362_not
g31226 not n19371 ; n19371_not
g31227 not n20685 ; n20685_not
g31228 not n13755 ; n13755_not
g31229 not n13746 ; n13746_not
g31230 not n13719 ; n13719_not
g31231 not n13926 ; n13926_not
g31232 not n19335 ; n19335_not
g31233 not n19326 ; n19326_not
g31234 not n16833 ; n16833_not
g31235 not n21549 ; n21549_not
g31236 not n14268 ; n14268_not
g31237 not n13683 ; n13683_not
g31238 not n13674 ; n13674_not
g31239 not n15177 ; n15177_not
g31240 not n19443 ; n19443_not
g31241 not n20577 ; n20577_not
g31242 not n13890 ; n13890_not
g31243 not n16725 ; n16725_not
g31244 not n14673 ; n14673_not
g31245 not n16068 ; n16068_not
g31246 not n21585 ; n21585_not
g31247 not n22845 ; n22845_not
g31248 not n15438 ; n15438_not
g31249 not n23277 ; n23277_not
g31250 not n14484 ; n14484_not
g31251 not n15447 ; n15447_not
g31252 not n20865 ; n20865_not
g31253 not n22089 ; n22089_not
g31254 not n16761 ; n16761_not
g31255 not n14448 ; n14448_not
g31256 not n19434 ; n19434_not
g31257 not n19407 ; n19407_not
g31258 not n22557 ; n22557_not
g31259 not n11955 ; n11955_not
g31260 not n13935 ; n13935_not
g31261 not n13854 ; n13854_not
g31262 not n13863 ; n13863_not
g31263 not n13827 ; n13827_not
g31264 not n15276 ; n15276_not
g31265 not n13269 ; n13269_not
g31266 not n15960 ; n15960_not
g31267 not n15249 ; n15249_not
g31268 not n15339 ; n15339_not
g31269 not n19191 ; n19191_not
g31270 not n22917 ; n22917_not
g31271 not n19182 ; n19182_not
g31272 not n20937 ; n20937_not
g31273 not n22881 ; n22881_not
g31274 not n15852 ; n15852_not
g31275 not n19146 ; n19146_not
g31276 not n19155 ; n19155_not
g31277 not n22377 ; n22377_not
g31278 not n16356 ; n16356_not
g31279 not n15267 ; n15267_not
g31280 not n15924 ; n15924_not
g31281 not n15726 ; n15726_not
g31282 not n21477 ; n21477_not
g31283 not n16905 ; n16905_not
g31284 not n22449 ; n22449_not
g31285 not n15294 ; n15294_not
g31286 not n15735 ; n15735_not
g31287 not n20649 ; n20649_not
g31288 not n20973 ; n20973_not
g31289 not n22485 ; n22485_not
g31290 not n15690 ; n15690_not
g31291 not n22197 ; n22197_not
g31292 not n11919 ; n11919_not
g31293 not n13638 ; n13638_not
g31294 not n13647 ; n13647_not
g31295 not n14196 ; n14196_not
g31296 not n13566 ; n13566_not
g31297 not n13575 ; n13575_not
g31298 not n13539 ; n13539_not
g31299 not n19290 ; n19290_not
g31300 not n13377 ; n13377_not
g31301 not n15366 ; n15366_not
g31302 not n12378 ; n12378_not
g31303 not n12396 ; n12396_not
g31304 not n19263 ; n19263_not
g31305 not n19254 ; n19254_not
g31306 not n15375 ; n15375_not
g31307 not n15861 ; n15861_not
g31308 not n13089 ; n13089_not
g31309 not n22269 ; n22269_not
g31310 not n14088 ; n14088_not
g31311 not n15870 ; n15870_not
g31312 not n19920 ; n19920_not
g31313 not n19218 ; n19218_not
g31314 not n19227 ; n19227_not
g31315 not n15591 ; n15591_not
g31316 not n21657 ; n21657_not
g31317 not n15654 ; n15654_not
g31318 not n16491 ; n16491_not
g31319 not n14781 ; n14781_not
g31320 not n19740 ; n19740_not
g31321 not n20793 ; n20793_not
g31322 not n16392 ; n16392_not
g31323 not n12828 ; n12828_not
g31324 not n12279 ; n12279_not
g31325 not n22665 ; n22665_not
g31326 not n19722 ; n19722_not
g31327 not n19731 ; n19731_not
g31328 not n14745 ; n14745_not
g31329 not n16284 ; n16284_not
g31330 not n16176 ; n16176_not
g31331 not n21189 ; n21189_not
g31332 not n12792 ; n12792_not
g31333 not n21837 ; n21837_not
g31334 not n14709 ; n14709_not
g31335 not n20388 ; n20388_not
g31336 not n16509 ; n16509_not
g31337 not n12756 ; n12756_not
g31338 not n12198 ; n12198_not
g31339 not n23169 ; n23169_not
g31340 not n21693 ; n21693_not
g31341 not n15627 ; n15627_not
g31342 not n16428 ; n16428_not
g31343 not n15618 ; n15618_not
g31344 not n20487 ; n20487_not
g31345 not n22737 ; n22737_not
g31346 not n14961 ; n14961_not
g31347 not n14925 ; n14925_not
g31348 not n20757 ; n20757_not
g31349 not n23097 ; n23097_not
g31350 not n22629 ; n22629_not
g31351 not n15807 ; n15807_not
g31352 not n21729 ; n21729_not
g31353 not n16248 ; n16248_not
g31354 not n21297 ; n21297_not
g31355 not n12864 ; n12864_not
g31356 not n22773 ; n22773_not
g31357 not n15582 ; n15582_not
g31358 not n14853 ; n14853_not
g31359 not n21765 ; n21765_not
g31360 not n15663 ; n15663_not
g31361 not n14817 ; n14817_not
g31362 not n13449 ; n13449_not
g31363 not n14628 ; n14628_not
g31364 not n21945 ; n21945_not
g31365 not n20829 ; n20829_not
g31366 not n14592 ; n14592_not
g31367 not n19551 ; n19551_not
g31368 not n19542 ; n19542_not
g31369 not n16617 ; n16617_not
g31370 not n22953 ; n22953_not
g31371 not n12576 ; n12576_not
g31372 not n19506 ; n19506_not
g31373 not n15483 ; n15483_not
g31374 not n19515 ; n19515_not
g31375 not n16653 ; n16653_not
g31376 not n21981 ; n21981_not
g31377 not n22575 ; n22575_not
g31378 not n22566 ; n22566_not
g31379 not n12954 ; n12954_not
g31380 not n11991 ; n11991_not
g31381 not n19470 ; n19470_not
g31382 not n15474 ; n15474_not
g31383 not n14556 ; n14556_not
g31384 not n13971 ; n13971_not
g31385 not n11982 ; n11982_not
g31386 not n13962 ; n13962_not
g31387 not n11946 ; n11946_not
g31388 not n20469 ; n20469_not
g31389 not n21369 ; n21369_not
g31390 not n21846 ; n21846_not
g31391 not n15555 ; n15555_not
g31392 not n21855 ; n21855_not
g31393 not n19650 ; n19650_not
g31394 not n15546 ; n15546_not
g31395 not n22809 ; n22809_not
g31396 not n14691 ; n14691_not
g31397 not n16545 ; n16545_not
g31398 not n15771 ; n15771_not
g31399 not n21873 ; n21873_not
g31400 not n15762 ; n15762_not
g31401 not n22593 ; n22593_not
g31402 not n15069 ; n15069_not
g31403 not n19623 ; n19623_not
g31404 not n19614 ; n19614_not
g31405 not n12981 ; n12981_not
g31406 not n12684 ; n12684_not
g31407 not n16581 ; n16581_not
g31408 not n15519 ; n15519_not
g31409 not n12648 ; n12648_not
g31410 not n21909 ; n21909_not
g31411 not n12099 ; n12099_not
g31412 not n14646 ; n14646_not
g31413 not n14637 ; n14637_not
g31414 not n23826 ; n23826_not
g31415 not n23835 ; n23835_not
g31416 not n18633 ; n18633_not
g31417 not n23754 ; n23754_not
g31418 not n23763 ; n23763_not
g31419 not n10956 ; n10956_not
g31420 not n23682 ; n23682_not
g31421 not n23691 ; n23691_not
g31422 not n18561 ; n18561_not
g31423 not n10398 ; n10398_not
g31424 not n23619 ; n23619_not
g31425 not n18525 ; n18525_not
g31426 not n10884 ; n10884_not
g31427 not n23538 ; n23538_not
g31428 not n23547 ; n23547_not
g31429 not n23466 ; n23466_not
g31430 not n23475 ; n23475_not
g31431 not n10299 ; n10299_not
g31432 not n23394 ; n23394_not
g31433 not n18453 ; n18453_not
g31434 not n17742 ; n17742_not
g31435 not n18372 ; n18372_not
g31436 not n17706 ; n17706_not
g31437 not n17715 ; n17715_not
g31438 not n18336 ; n18336_not
g31439 not n17670 ; n17670_not
g31440 not n17634 ; n17634_not
g31441 not n17049 ; n17049_not
g31442 not n17085 ; n17085_not
g31443 not n11829 ; n11829_not
g31444 not n11793 ; n11793_not
g31445 not n11757 ; n11757_not
g31446 not n11685 ; n11685_not
g31447 not n11649 ; n11649_not
g31448 not n18426 ; n18426_not
g31449 not n11577 ; n11577_not
g31450 not n19029 ; n19029_not
g31451 not n11469 ; n11469_not
g31452 not n18921 ; n18921_not
g31453 not n11397 ; n11397_not
g31454 not n10839 ; n10839_not
g31455 not n18813 ; n18813_not
g31456 not n10767 ; n10767_not
g31457 not n10758 ; n10758_not
g31458 not n10695 ; n10695_not
g31459 not n10686 ; n10686_not
g31460 not n10659 ; n10659_not
g31461 not n18741 ; n18741_not
g31462 not n10578 ; n10578_not
g31463 not n10587 ; n10587_not
g31464 not n18705 ; n18705_not
g31465 not n10992 ; n10992_not
g31466 not n23970 ; n23970_not
g31467 not n10479 ; n10479_not
g31468 not n23907 ; n23907_not
g31469 not n17355 ; n17355_not
g31470 not n23655 ; n23655_not
g31471 not n23646 ; n23646_not
g31472 not n24546 ; n24546_not
g31473 not n17319 ; n17319_not
g31474 not n23727 ; n23727_not
g31475 not n23718 ; n23718_not
g31476 not n24564 ; n24564_not
g31477 not n17940 ; n17940_not
g31478 not n17274 ; n17274_not
g31479 not n17283 ; n17283_not
g31480 not n17904 ; n17904_not
g31481 not n17247 ; n17247_not
g31482 not n17238 ; n17238_not
g31483 not n23790 ; n23790_not
g31484 not n24645 ; n24645_not
g31485 not n24663 ; n24663_not
g31486 not n23871 ; n23871_not
g31487 not n23862 ; n23862_not
g31488 not n17832 ; n17832_not
g31489 not n17175 ; n17175_not
g31490 not n17166 ; n17166_not
g31491 not n23943 ; n23943_not
g31492 not n23934 ; n23934_not
g31493 not n24717 ; n24717_not
g31494 not n17760 ; n17760_not
g31495 not n17643 ; n17643_not
g31496 not n18264 ; n18264_not
g31497 not n17607 ; n17607_not
g31498 not n23367 ; n23367_not
g31499 not n18228 ; n18228_not
g31500 not n17562 ; n17562_not
g31501 not n17571 ; n17571_not
g31502 not n23358 ; n23358_not
g31503 not n24339 ; n24339_not
g31504 not n24357 ; n24357_not
g31505 not n23439 ; n23439_not
g31506 not n18192 ; n18192_not
g31507 not n17535 ; n17535_not
g31508 not n17526 ; n17526_not
g31509 not n18156 ; n18156_not
g31510 not n17490 ; n17490_not
g31511 not n24393 ; n24393_not
g31512 not n17463 ; n17463_not
g31513 not n17454 ; n17454_not
g31514 not n18084 ; n18084_not
g31515 not n17418 ; n17418_not
g31516 not n17427 ; n17427_not
g31517 not n23583 ; n23583_not
g31518 not n23574 ; n23574_not
g31519 not n18048 ; n18048_not
g31520 not n17391 ; n17391_not
g31521 not n17382 ; n17382_not
g31522 not n24492 ; n24492_not
g31523 not n17346 ; n17346_not
g31524 not n19812 ; n19812_not
g31525 not n19119 ; n19119_not
g31526 not n16941 ; n16941_not
g31527 not n23944 ; n23944_not
g31528 not n20974 ; n20974_not
g31529 not n17464 ; n17464_not
g31530 not n22954 ; n22954_not
g31531 not n13576 ; n13576_not
g31532 not n16177 ; n16177_not
g31533 not n18292 ; n18292_not
g31534 not n11875 ; n11875_not
g31535 not n17284 ; n17284_not
g31536 not n23908 ; n23908_not
g31537 not n16618 ; n16618_not
g31538 not n16627 ; n16627_not
g31539 not n18265 ; n18265_not
g31540 not n11848 ; n11848_not
g31541 not n21766 ; n21766_not
g31542 not n16843 ; n16843_not
g31543 not n16834 ; n16834_not
g31544 not n20866 ; n20866_not
g31545 not n20875 ; n20875_not
g31546 not n12469 ; n12469_not
g31547 not n18373 ; n18373_not
g31548 not n23278 ; n23278_not
g31549 not n19039 ; n19039_not
g31550 not n18337 ; n18337_not
g31551 not n12991 ; n12991_not
g31552 not n22666 ; n22666_not
g31553 not n16654 ; n16654_not
g31554 not n23980 ; n23980_not
g31555 not n21658 ; n21658_not
g31556 not n16069 ; n16069_not
g31557 not n20938 ; n20938_not
g31558 not n20947 ; n20947_not
g31559 not n16807 ; n16807_not
g31560 not n10588 ; n10588_not
g31561 not n12982 ; n12982_not
g31562 not n21694 ; n21694_not
g31563 not n20983 ; n20983_not
g31564 not n16546 ; n16546_not
g31565 not n14089 ; n14089_not
g31566 not n24376 ; n24376_not
g31567 not n16555 ; n16555_not
g31568 not n19750 ; n19750_not
g31569 not n18157 ; n18157_not
g31570 not n21874 ; n21874_not
g31571 not n16357 ; n16357_not
g31572 not n13099 ; n13099_not
g31573 not n24394 ; n24394_not
g31574 not n19066 ; n19066_not
g31575 not n19093 ; n19093_not
g31576 not n17536 ; n17536_not
g31577 not n17176 ; n17176_not
g31578 not n21892 ; n21892_not
g31579 not n22594 ; n22594_not
g31580 not n16519 ; n16519_not
g31581 not n16915 ; n16915_not
g31582 not n23584 ; n23584_not
g31583 not n16249 ; n16249_not
g31584 not n17248 ; n17248_not
g31585 not n18229 ; n18229_not
g31586 not n16285 ; n16285_not
g31587 not n16591 ; n16591_not
g31588 not n16582 ; n16582_not
g31589 not n18391 ; n18391_not
g31590 not n13648 ; n13648_not
g31591 not n19732 ; n19732_not
g31592 not n21838 ; n21838_not
g31593 not n11398 ; n11398_not
g31594 not n11578 ; n11578_not
g31595 not n19741 ; n19741_not
g31596 not n18193 ; n18193_not
g31597 not n19084 ; n19084_not
g31598 not n23872 ; n23872_not
g31599 not n22990 ; n22990_not
g31600 not n16870 ; n16870_not
g31601 not n15448 ; n15448_not
g31602 not n14818 ; n14818_not
g31603 not n16735 ; n16735_not
g31604 not n11992 ; n11992_not
g31605 not n14827 ; n14827_not
g31606 not n15628 ; n15628_not
g31607 not n14791 ; n14791_not
g31608 not n15664 ; n15664_not
g31609 not n14782 ; n14782_not
g31610 not n11479 ; n11479_not
g31611 not n15376 ; n15376_not
g31612 not n22846 ; n22846_not
g31613 not n20659 ; n20659_not
g31614 not n17392 ; n17392_not
g31615 not n22738 ; n22738_not
g31616 not n13486 ; n13486_not
g31617 not n15736 ; n15736_not
g31618 not n10993 ; n10993_not
g31619 not n14746 ; n14746_not
g31620 not n14755 ; n14755_not
g31621 not n14890 ; n14890_not
g31622 not n19660 ; n19660_not
g31623 not n14926 ; n14926_not
g31624 not n14935 ; n14935_not
g31625 not n12928 ; n12928_not
g31626 not n12919 ; n12919_not
g31627 not n15556 ; n15556_not
g31628 not n22774 ; n22774_not
g31629 not n15484 ; n15484_not
g31630 not n14971 ; n14971_not
g31631 not n14962 ; n14962_not
g31632 not n10957 ; n10957_not
g31633 not n14863 ; n14863_not
g31634 not n21298 ; n21298_not
g31635 not n20578 ; n20578_not
g31636 not n20587 ; n20587_not
g31637 not n15592 ; n15592_not
g31638 not n14854 ; n14854_not
g31639 not n18427 ; n18427_not
g31640 not n21478 ; n21478_not
g31641 not n15871 ; n15871_not
g31642 not n20767 ; n20767_not
g31643 not n20758 ; n20758_not
g31644 not n10768 ; n10768_not
g31645 not n20794 ; n20794_not
g31646 not n10696 ; n10696_not
g31647 not n16690 ; n16690_not
g31648 not n18931 ; n18931_not
g31649 not n17428 ; n17428_not
g31650 not n18922 ; n18922_not
g31651 not n20839 ; n20839_not
g31652 not n23548 ; n23548_not
g31653 not n15925 ; n15925_not
g31654 not n22918 ; n22918_not
g31655 not n21586 ; n21586_not
g31656 not n15961 ; n15961_not
g31657 not n11956 ; n11956_not
g31658 not n16663 ; n16663_not
g31659 not n10885 ; n10885_not
g31660 not n10849 ; n10849_not
g31661 not n15772 ; n15772_not
g31662 not n20695 ; n20695_not
g31663 not n20686 ; n20686_not
g31664 not n16726 ; n16726_not
g31665 not n14719 ; n14719_not
g31666 not n19624 ; n19624_not
g31667 not n15187 ; n15187_not
g31668 not n15178 ; n15178_not
g31669 not n23476 ; n23476_not
g31670 not n15808 ; n15808_not
g31671 not n17770 ; n17770_not
g31672 not n17356 ; n17356_not
g31673 not n18436 ; n18436_not
g31674 not n16771 ; n16771_not
g31675 not n16762 ; n16762_not
g31676 not n22882 ; n22882_not
g31677 not n15268 ; n15268_not
g31678 not n18409 ; n18409_not
g31679 not n13378 ; n13378_not
g31680 not n12793 ; n12793_not
g31681 not n14269 ; n14269_not
g31682 not n17716 ; n17716_not
g31683 not n23368 ; n23368_not
g31684 not n17905 ; n17905_not
g31685 not n23728 ; n23728_not
g31686 not n11857 ; n11857_not
g31687 not n22198 ; n22198_not
g31688 not n19336 ; n19336_not
g31689 not n22378 ; n22378_not
g31690 not n12829 ; n12829_not
g31691 not n17644 ; n17644_not
g31692 not n17941 ; n17941_not
g31693 not n18643 ; n18643_not
g31694 not n18634 ; n18634_not
g31695 not n14377 ; n14377_not
g31696 not n11767 ; n11767_not
g31697 not n23764 ; n23764_not
g31698 not n12865 ; n12865_not
g31699 not n19480 ; n19480_not
g31700 not n19813 ; n19813_not
g31701 not n18607 ; n18607_not
g31702 not n11758 ; n11758_not
g31703 not n14449 ; n14449_not
g31704 not n24547 ; n24547_not
g31705 not n24529 ; n24529_not
g31706 not n19264 ; n19264_not
g31707 not n13936 ; n13936_not
g31708 not n22558 ; n22558_not
g31709 not n14485 ; n14485_not
g31710 not n18751 ; n18751_not
g31711 not n13756 ; n13756_not
g31712 not n11695 ; n11695_not
g31713 not n18742 ; n18742_not
g31714 not n19408 ; n19408_not
g31715 not n23692 ; n23692_not
g31716 not n11659 ; n11659_not
g31717 not n18715 ; n18715_not
g31718 not n11686 ; n11686_not
g31719 not n18706 ; n18706_not
g31720 not n17833 ; n17833_not
g31721 not n13459 ; n13459_not
g31722 not n17680 ; n17680_not
g31723 not n18670 ; n18670_not
g31724 not n13387 ; n13387_not
g31725 not n23656 ; n23656_not
g31726 not n13198 ; n13198_not
g31727 not n13972 ; n13972_not
g31728 not n24628 ; n24628_not
g31729 not n12649 ; n12649_not
g31730 not n20389 ; n20389_not
g31731 not n24646 ; n24646_not
g31732 not n14197 ; n14197_not
g31733 not n19372 ; n19372_not
g31734 not n19444 ; n19444_not
g31735 not n12757 ; n12757_not
g31736 not n24682 ; n24682_not
g31737 not n17059 ; n17059_not
g31738 not n12685 ; n12685_not
g31739 not n11866 ; n11866_not
g31740 not n18049 ; n18049_not
g31741 not n19156 ; n19156_not
g31742 not n12577 ; n12577_not
g31743 not n18526 ; n18526_not
g31744 not n18814 ; n18814_not
g31745 not n16429 ; n16429_not
g31746 not n23836 ; n23836_not
g31747 not n12955 ; n12955_not
g31748 not n12937 ; n12937_not
g31749 not n18535 ; n18535_not
g31750 not n13279 ; n13279_not
g31751 not n24475 ; n24475_not
g31752 not n11794 ; n11794_not
g31753 not n14593 ; n14593_not
g31754 not n19516 ; n19516_not
g31755 not n17572 ; n17572_not
g31756 not n21982 ; n21982_not
g31757 not n19921 ; n19921_not
g31758 not n19192 ; n19192_not
g31759 not n16393 ; n16393_not
g31760 not n14629 ; n14629_not
g31761 not n18490 ; n18490_not
g31762 not n12964 ; n12964_not
g31763 not n11587 ; n11587_not
g31764 not n18085 ; n18085_not
g31765 not n13828 ; n13828_not
g31766 not n24781 ; n24781_not
g31767 not n19552 ; n19552_not
g31768 not n22486 ; n22486_not
g31769 not n18463 ; n18463_not
g31770 not n13792 ; n13792_not
g31771 not n17608 ; n17608_not
g31772 not n18571 ; n18571_not
g31773 not n13684 ; n13684_not
g31774 not n18454 ; n18454_not
g31775 not n18562 ; n18562_not
g31776 not n16906 ; n16906_not
g31777 not n23098 ; n23098_not
g31778 not n24493 ; n24493_not
g31779 not n19228 ; n19228_not
g31780 not n13864 ; n13864_not
g31781 not n16942 ; n16942_not
g31782 not n18823 ; n18823_not
g31783 not n18850 ; n18850_not
g31784 not n14557 ; n14557_not
g31785 not n21946 ; n21946_not
g31786 not n16951 ; n16951_not
g31787 not n21596 ; n21596_not
g31788 not n17807 ; n17807_not
g31789 not n13829 ; n13829_not
g31790 not n16844 ; n16844_not
g31791 not n18464 ; n18464_not
g31792 not n14675 ; n14675_not
g31793 not n16808 ; n16808_not
g31794 not n21992 ; n21992_not
g31795 not n24782 ; n24782_not
g31796 not n21587 ; n21587_not
g31797 not n17870 ; n17870_not
g31798 not n21983 ; n21983_not
g31799 not n13937 ; n13937_not
g31800 not n15449 ; n15449_not
g31801 not n17753 ; n17753_not
g31802 not n17771 ; n17771_not
g31803 not n21668 ; n21668_not
g31804 not n21767 ; n21767_not
g31805 not n21659 ; n21659_not
g31806 not n13793 ; n13793_not
g31807 not n16178 ; n16178_not
g31808 not n17393 ; n17393_not
g31809 not n17843 ; n17843_not
g31810 not n18536 ; n18536_not
g31811 not n17744 ; n17744_not
g31812 not n21776 ; n21776_not
g31813 not n21695 ; n21695_not
g31814 not n17834 ; n17834_not
g31815 not n16187 ; n16187_not
g31816 not n17780 ; n17780_not
g31817 not n13865 ; n13865_not
g31818 not n16916 ; n16916_not
g31819 not n15485 ; n15485_not
g31820 not n15377 ; n15377_not
g31821 not n13973 ; n13973_not
g31822 not n22739 ; n22739_not
g31823 not n24683 ; n24683_not
g31824 not n17717 ; n17717_not
g31825 not n24764 ; n24764_not
g31826 not n22748 ; n22748_not
g31827 not n14792 ; n14792_not
g31828 not n14198 ; n14198_not
g31829 not n21299 ; n21299_not
g31830 not n14828 ; n14828_not
g31831 not n17609 ; n17609_not
g31832 not n14864 ; n14864_not
g31833 not n21875 ; n21875_not
g31834 not n14279 ; n14279_not
g31835 not n12389 ; n12389_not
g31836 not n24287 ; n24287_not
g31837 not n16259 ; n16259_not
g31838 not n14936 ; n14936_not
g31839 not n22667 ; n22667_not
g31840 not n13577 ; n13577_not
g31841 not n22595 ; n22595_not
g31842 not n17645 ; n17645_not
g31843 not n10589 ; n10589_not
g31844 not n17465 ; n17465_not
g31845 not n14666 ; n14666_not
g31846 not n13685 ; n13685_not
g31847 not n16286 ; n16286_not
g31848 not n14648 ; n14648_not
g31849 not n14657 ; n14657_not
g31850 not n22577 ; n22577_not
g31851 not n17573 ; n17573_not
g31852 not n24458 ; n24458_not
g31853 not n21857 ; n21857_not
g31854 not n24377 ; n24377_not
g31855 not n17537 ; n17537_not
g31856 not n24476 ; n24476_not
g31857 not n16880 ; n16880_not
g31858 not n24359 ; n24359_not
g31859 not n14756 ; n14756_not
g31860 not n13649 ; n13649_not
g31861 not n16295 ; n16295_not
g31862 not n19733 ; n19733_not
g31863 not n24269 ; n24269_not
g31864 not n22676 ; n22676_not
g31865 not n17735 ; n17735_not
g31866 not n17681 ; n17681_not
g31867 not n15188 ; n15188_not
g31868 not n14594 ; n14594_not
g31869 not n10769 ; n10769_not
g31870 not n23477 ; n23477_not
g31871 not n17429 ; n17429_not
g31872 not n18428 ; n18428_not
g31873 not n24665 ; n24665_not
g31874 not n19094 ; n19094_not
g31875 not n13757 ; n13757_not
g31876 not n15287 ; n15287_not
g31877 not n23369 ; n23369_not
g31878 not n14972 ; n14972_not
g31879 not n14387 ; n14387_not
g31880 not n14378 ; n14378_not
g31881 not n14459 ; n14459_not
g31882 not n16952 ; n16952_not
g31883 not n21956 ; n21956_not
g31884 not n21488 ; n21488_not
g31885 not n21479 ; n21479_not
g31886 not n24629 ; n24629_not
g31887 not n14486 ; n14486_not
g31888 not n14495 ; n14495_not
g31889 not n21947 ; n21947_not
g31890 not n18392 ; n18392_not
g31891 not n10697 ; n10697_not
g31892 not n18374 ; n18374_not
g31893 not n14558 ; n14558_not
g31894 not n14567 ; n14567_not
g31895 not n11867 ; n11867_not
g31896 not n12686 ; n12686_not
g31897 not n20876 ; n20876_not
g31898 not n23981 ; n23981_not
g31899 not n10895 ; n10895_not
g31900 not n10886 ; n10886_not
g31901 not n18239 ; n18239_not
g31902 not n19373 ; n19373_not
g31903 not n16736 ; n16736_not
g31904 not n16493 ; n16493_not
g31905 not n16466 ; n16466_not
g31906 not n23729 ; n23729_not
g31907 not n22991 ; n22991_not
g31908 not n18932 ; n18932_not
g31909 not n18266 ; n18266_not
g31910 not n18275 ; n18275_not
g31911 not n11957 ; n11957_not
g31912 not n23945 ; n23945_not
g31913 not n10967 ; n10967_not
g31914 not n10958 ; n10958_not
g31915 not n23765 ; n23765_not
g31916 not n17285 ; n17285_not
g31917 not n23297 ; n23297_not
g31918 not n12758 ; n12758_not
g31919 not n20984 ; n20984_not
g31920 not n23549 ; n23549_not
g31921 not n15935 ; n15935_not
g31922 not n16556 ; n16556_not
g31923 not n15269 ; n15269_not
g31924 not n23279 ; n23279_not
g31925 not n16394 ; n16394_not
g31926 not n20948 ; n20948_not
g31927 not n18824 ; n18824_not
g31928 not n18167 ; n18167_not
g31929 not n18158 ; n18158_not
g31930 not n10859 ; n10859_not
g31931 not n22847 ; n22847_not
g31932 not n19409 ; n19409_not
g31933 not n18860 ; n18860_not
g31934 not n22964 ; n22964_not
g31935 not n18194 ; n18194_not
g31936 not n12695 ; n12695_not
g31937 not n22955 ; n22955_not
g31938 not n22199 ; n22199_not
g31939 not n23873 ; n23873_not
g31940 not n11768 ; n11768_not
g31941 not n19922 ; n19922_not
g31942 not n19931 ; n19931_not
g31943 not n23099 ; n23099_not
g31944 not n23585 ; n23585_not
g31945 not n17177 ; n17177_not
g31946 not n16079 ; n16079_not
g31947 not n19229 ; n19229_not
g31948 not n12956 ; n12956_not
g31949 not n11696 ; n11696_not
g31950 not n12479 ; n12479_not
g31951 not n20588 ; n20588_not
g31952 not n12992 ; n12992_not
g31953 not n19157 ; n19157_not
g31954 not n19814 ; n19814_not
g31955 not n19823 ; n19823_not
g31956 not n19850 ; n19850_not
g31957 not n19193 ; n19193_not
g31958 not n23837 ; n23837_not
g31959 not n12659 ; n12659_not
g31960 not n20768 ; n20768_not
g31961 not n18338 ; n18338_not
g31962 not n19337 ; n19337_not
g31963 not n16439 ; n16439_not
g31964 not n18347 ; n18347_not
g31965 not n23909 ; n23909_not
g31966 not n18383 ; n18383_not
g31967 not n17249 ; n17249_not
g31968 not n22379 ; n22379_not
g31969 not n10994 ; n10994_not
g31970 not n22388 ; n22388_not
g31971 not n16484 ; n16484_not
g31972 not n20696 ; n20696_not
g31973 not n12929 ; n12929_not
g31974 not n19265 ; n19265_not
g31975 not n12578 ; n12578_not
g31976 not n12587 ; n12587_not
g31977 not n15692 ; n15692_not
g31978 not n11588 ; n11588_not
g31979 not n22496 ; n22496_not
g31980 not n15773 ; n15773_not
g31981 not n22487 ; n22487_not
g31982 not n20399 ; n20399_not
g31983 not n18680 ; n18680_not
g31984 not n19517 ; n19517_not
g31985 not n11885 ; n11885_not
g31986 not n16772 ; n16772_not
g31987 not n23657 ; n23657_not
g31988 not n15809 ; n15809_not
g31989 not n15971 ; n15971_not
g31990 not n15962 ; n15962_not
g31991 not n22784 ; n22784_not
g31992 not n15593 ; n15593_not
g31993 not n18716 ; n18716_not
g31994 not n16592 ; n16592_not
g31995 not n18059 ; n18059_not
g31996 not n12875 ; n12875_not
g31997 not n12866 ; n12866_not
g31998 not n11993 ; n11993_not
g31999 not n22775 ; n22775_not
g32000 not n15665 ; n15665_not
g32001 not n16358 ; n16358_not
g32002 not n15629 ; n15629_not
g32003 not n18644 ; n18644_not
g32004 not n17942 ; n17942_not
g32005 not n12839 ; n12839_not
g32006 not n22892 ; n22892_not
g32007 not n17951 ; n17951_not
g32008 not n18608 ; n18608_not
g32009 not n15737 ; n15737_not
g32010 not n16628 ; n16628_not
g32011 not n13388 ; n13388_not
g32012 not n22883 ; n22883_not
g32013 not n16367 ; n16367_not
g32014 not n18095 ; n18095_not
g32015 not n18572 ; n18572_not
g32016 not n15557 ; n15557_not
g32017 not n18086 ; n18086_not
g32018 not n22856 ; n22856_not
g32019 not n18752 ; n18752_not
g32020 not n23693 ; n23693_not
g32021 not n19553 ; n19553_not
g32022 not n22928 ; n22928_not
g32023 not n12794 ; n12794_not
g32024 not n17357 ; n17357_not
g32025 not n19625 ; n19625_not
g32026 not n19661 ; n19661_not
g32027 not n19445 ; n19445_not
g32028 not n19481 ; n19481_not
g32029 not n15926 ; n15926_not
g32030 not n12767 ; n12767_not
g32031 not n17906 ; n17906_not
g32032 not n15890 ; n15890_not
g32033 not n16664 ; n16664_not
g32034 not n22919 ; n22919_not
g32035 not n17915 ; n17915_not
g32036 not n14496 ; n14496_not
g32037 not n23991 ; n23991_not
g32038 not n19194 ; n19194_not
g32039 not n17745 ; n17745_not
g32040 not n11967 ; n11967_not
g32041 not n24747 ; n24747_not
g32042 not n11958 ; n11958_not
g32043 not n15783 ; n15783_not
g32044 not n19761 ; n19761_not
g32045 not n16494 ; n16494_not
g32046 not n13866 ; n13866_not
g32047 not n19446 ; n19446_not
g32048 not n19752 ; n19752_not
g32049 not n22497 ; n22497_not
g32050 not n23694 ; n23694_not
g32051 not n11769 ; n11769_not
g32052 not n19491 ; n19491_not
g32053 not n19482 ; n19482_not
g32054 not n24765 ; n24765_not
g32055 not n16665 ; n16665_not
g32056 not n24495 ; n24495_not
g32057 not n17736 ; n17736_not
g32058 not n13983 ; n13983_not
g32059 not n13974 ; n13974_not
g32060 not n14568 ; n14568_not
g32061 not n15819 ; n15819_not
g32062 not n21993 ; n21993_not
g32063 not n19068 ; n19068_not
g32064 not n13947 ; n13947_not
g32065 not n13938 ; n13938_not
g32066 not n11994 ; n11994_not
g32067 not n17367 ; n17367_not
g32068 not n23982 ; n23982_not
g32069 not n17358 ; n17358_not
g32070 not n17394 ; n17394_not
g32071 not n15846 ; n15846_not
g32072 not n17718 ; n17718_not
g32073 not n11697 ; n11697_not
g32074 not n15774 ; n15774_not
g32075 not n19824 ; n19824_not
g32076 not n12768 ; n12768_not
g32077 not n13659 ; n13659_not
g32078 not n19563 ; n19563_not
g32079 not n19554 ; n19554_not
g32080 not n17880 ; n17880_not
g32081 not n24648 ; n24648_not
g32082 not n23919 ; n23919_not
g32083 not n13587 ; n13587_not
g32084 not n13578 ; n13578_not
g32085 not n23847 ; n23847_not
g32086 not n16593 ; n16593_not
g32087 not n23838 ; n23838_not
g32088 not n19662 ; n19662_not
g32089 not n15891 ; n15891_not
g32090 not n17844 ; n17844_not
g32091 not n17178 ; n17178_not
g32092 not n17187 ; n17187_not
g32093 not n11886 ; n11886_not
g32094 not n12696 ; n12696_not
g32095 not n16557 ; n16557_not
g32096 not n19590 ; n19590_not
g32097 not n13488 ; n13488_not
g32098 not n19626 ; n19626_not
g32099 not n19635 ; n19635_not
g32100 not n17808 ; n17808_not
g32101 not n24666 ; n24666_not
g32102 not n13479 ; n13479_not
g32103 not n12876 ; n12876_not
g32104 not n13839 ; n13839_not
g32105 not n17772 ; n17772_not
g32106 not n17952 ; n17952_not
g32107 not n17295 ; n17295_not
g32108 not n14388 ; n14388_not
g32109 not n13794 ; n13794_not
g32110 not n19518 ; n19518_not
g32111 not n17286 ; n17286_not
g32112 not n19455 ; n19455_not
g32113 not n19770 ; n19770_not
g32114 not n19527 ; n19527_not
g32115 not n16629 ; n16629_not
g32116 not n13758 ; n13758_not
g32117 not n13767 ; n13767_not
g32118 not n24594 ; n24594_not
g32119 not n23775 ; n23775_not
g32120 not n17916 ; n17916_not
g32121 not n17259 ; n17259_not
g32122 not n22389 ; n22389_not
g32123 not n13686 ; n13686_not
g32124 not n13695 ; n13695_not
g32125 not n23766 ; n23766_not
g32126 not n12588 ; n12588_not
g32127 not n19860 ; n19860_not
g32128 not n19167 ; n19167_not
g32129 not n19158 ; n19158_not
g32130 not n16917 ; n16917_not
g32131 not n19707 ; n19707_not
g32132 not n17727 ; n17727_not
g32133 not n10779 ; n10779_not
g32134 not n15936 ; n15936_not
g32135 not n20949 ; n20949_not
g32136 not n18825 ; n18825_not
g32137 not n18384 ; n18384_not
g32138 not n19419 ; n19419_not
g32139 not n18393 ; n18393_not
g32140 not n15189 ; n15189_not
g32141 not n10698 ; n10698_not
g32142 not n20985 ; n20985_not
g32143 not n23298 ; n23298_not
g32144 not n15873 ; n15873_not
g32145 not n22893 ; n22893_not
g32146 not n12957 ; n12957_not
g32147 not n21489 ; n21489_not
g32148 not n16773 ; n16773_not
g32149 not n18933 ; n18933_not
g32150 not n17646 ; n17646_not
g32151 not n17655 ; n17655_not
g32152 not n14973 ; n14973_not
g32153 not n21669 ; n21669_not
g32154 not n15459 ; n15459_not
g32155 not n20877 ; n20877_not
g32156 not n15387 ; n15387_not
g32157 not n15378 ; n15378_not
g32158 not n17691 ; n17691_not
g32159 not n17682 ; n17682_not
g32160 not n18348 ; n18348_not
g32161 not n22929 ; n22929_not
g32162 not n11895 ; n11895_not
g32163 not n21597 ; n21597_not
g32164 not n18861 ; n18861_not
g32165 not n22677 ; n22677_not
g32166 not n15972 ; n15972_not
g32167 not n18645 ; n18645_not
g32168 not n13497 ; n13497_not
g32169 not n10968 ; n10968_not
g32170 not n22749 ; n22749_not
g32171 not n23595 ; n23595_not
g32172 not n18537 ; n18537_not
g32173 not n23586 ; n23586_not
g32174 not n19347 ; n19347_not
g32175 not n18609 ; n18609_not
g32176 not n16809 ; n16809_not
g32177 not n23289 ; n23289_not
g32178 not n23739 ; n23739_not
g32179 not n10896 ; n10896_not
g32180 not n22785 ; n22785_not
g32181 not n19338 ; n19338_not
g32182 not n18573 ; n18573_not
g32183 not n23667 ; n23667_not
g32184 not n23658 ; n23658_not
g32185 not n18753 ; n18753_not
g32186 not n15864 ; n15864_not
g32187 not n10599 ; n10599_not
g32188 not n23379 ; n23379_not
g32189 not n18447 ; n18447_not
g32190 not n18717 ; n18717_not
g32191 not n16845 ; n16845_not
g32192 not n18465 ; n18465_not
g32193 not n13389 ; n13389_not
g32194 not n22857 ; n22857_not
g32195 not n19383 ; n19383_not
g32196 not n18681 ; n18681_not
g32197 not n23946 ; n23946_not
g32198 not n23955 ; n23955_not
g32199 not n19374 ; n19374_not
g32200 not n23874 ; n23874_not
g32201 not n23883 ; n23883_not
g32202 not n23487 ; n23487_not
g32203 not n19077 ; n19077_not
g32204 not n19095 ; n19095_not
g32205 not n19932 ; n19932_not
g32206 not n19059 ; n19059_not
g32207 not n14685 ; n14685_not
g32208 not n11589 ; n11589_not
g32209 not n18168 ; n18168_not
g32210 not n16881 ; n16881_not
g32211 not n20697 ; n20697_not
g32212 not n22965 ; n22965_not
g32213 not n17547 ; n17547_not
g32214 not n17538 ; n17538_not
g32215 not n14757 ; n14757_not
g32216 not n16296 ; n16296_not
g32217 not n15675 ; n15675_not
g32218 not n21957 ; n21957_not
g32219 not n12975 ; n12975_not
g32220 not n12993 ; n12993_not
g32221 not n17439 ; n17439_not
g32222 not n18096 ; n18096_not
g32223 not n20589 ; n20589_not
g32224 not n14667 ; n14667_not
g32225 not n16368 ; n16368_not
g32226 not n24459 ; n24459_not
g32227 not n15747 ; n15747_not
g32228 not n19239 ; n19239_not
g32229 not n23559 ; n23559_not
g32230 not n15738 ; n15738_not
g32231 not n18429 ; n18429_not
g32232 not n17475 ; n17475_not
g32233 not n17466 ; n17466_not
g32234 not n23478 ; n23478_not
g32235 not n15495 ; n15495_not
g32236 not n15486 ; n15486_not
g32237 not n16953 ; n16953_not
g32238 not n14937 ; n14937_not
g32239 not n18276 ; n18276_not
g32240 not n17619 ; n17619_not
g32241 not n15567 ; n15567_not
g32242 not n15558 ; n15558_not
g32243 not n16188 ; n16188_not
g32244 not n14865 ; n14865_not
g32245 not n15594 ; n15594_not
g32246 not n20769 ; n20769_not
g32247 not n17583 ; n17583_not
g32248 not n17574 ; n17574_not
g32249 not n14829 ; n14829_not
g32250 not n21777 ; n21777_not
g32251 not n14793 ; n14793_not
g32252 not n15639 ; n15639_not
g32253 not n19275 ; n19275_not
g32254 not n15666 ; n15666_not
g32255 not n19266 ; n19266_not
g32256 not n16737 ; n16737_not
g32257 not n10897 ; n10897_not
g32258 not n12769 ; n12769_not
g32259 not n22498 ; n22498_not
g32260 not n13588 ; n13588_not
g32261 not n11599 ; n11599_not
g32262 not n23956 ; n23956_not
g32263 not n22966 ; n22966_not
g32264 not n23776 ; n23776_not
g32265 not n12697 ; n12697_not
g32266 not n24478 ; n24478_not
g32267 not n24289 ; n24289_not
g32268 not n24784 ; n24784_not
g32269 not n11698 ; n11698_not
g32270 not n13489 ; n13489_not
g32271 not n23848 ; n23848_not
g32272 not n11896 ; n11896_not
g32273 not n23596 ; n23596_not
g32274 not n13696 ; n13696_not
g32275 not n22786 ; n22786_not
g32276 not n12994 ; n12994_not
g32277 not n23668 ; n23668_not
g32278 not n11779 ; n11779_not
g32279 not n24496 ; n24496_not
g32280 not n11968 ; n11968_not
g32281 not n21877 ; n21877_not
g32282 not n24577 ; n24577_not
g32283 not n23992 ; n23992_not
g32284 not n24649 ; n24649_not
g32285 not n12877 ; n12877_not
g32286 not n23488 ; n23488_not
g32287 not n13768 ; n13768_not
g32288 not n22894 ; n22894_not
g32289 not n22858 ; n22858_not
g32290 not n23884 ; n23884_not
g32291 not n11869 ; n11869_not
g32292 not n24595 ; n24595_not
g32293 not n22678 ; n22678_not
g32294 not n11887 ; n11887_not
g32295 not n24748 ; n24748_not
g32296 not n22588 ; n22588_not
g32297 not n22597 ; n22597_not
g32298 not n12589 ; n12589_not
g32299 not n10969 ; n10969_not
g32300 not n19069 ; n19069_not
g32301 not n16567 ; n16567_not
g32302 not n15676 ; n15676_not
g32303 not n16558 ; n16558_not
g32304 not n17188 ; n17188_not
g32305 not n19096 ; n19096_not
g32306 not n15748 ; n15748_not
g32307 not n15784 ; n15784_not
g32308 not n18466 ; n18466_not
g32309 not n18475 ; n18475_not
g32310 not n15199 ; n15199_not
g32311 not n19168 ; n19168_not
g32312 not n17098 ; n17098_not
g32313 not n16468 ; n16468_not
g32314 not n18538 ; n18538_not
g32315 not n18547 ; n18547_not
g32316 not n18583 ; n18583_not
g32317 not n18574 ; n18574_not
g32318 not n19276 ; n19276_not
g32319 not n14695 ; n14695_not
g32320 not n16666 ; n16666_not
g32321 not n20698 ; n20698_not
g32322 not n14758 ; n14758_not
g32323 not n14767 ; n14767_not
g32324 not n16675 ; n16675_not
g32325 not n15388 ; n15388_not
g32326 not n14794 ; n14794_not
g32327 not n14839 ; n14839_not
g32328 not n20599 ; n20599_not
g32329 not n14875 ; n14875_not
g32330 not n14866 ; n14866_not
g32331 not n17296 ; n17296_not
g32332 not n15496 ; n15496_not
g32333 not n14947 ; n14947_not
g32334 not n14938 ; n14938_not
g32335 not n15568 ; n15568_not
g32336 not n14974 ; n14974_not
g32337 not n16639 ; n16639_not
g32338 not n14983 ; n14983_not
g32339 not n16594 ; n16594_not
g32340 not n19528 ; n19528_not
g32341 not n16369 ; n16369_not
g32342 not n18871 ; n18871_not
g32343 not n18862 ; n18862_not
g32344 not n19564 ; n19564_not
g32345 not n18907 ; n18907_not
g32346 not n18943 ; n18943_not
g32347 not n18934 ; n18934_not
g32348 not n19636 ; n19636_not
g32349 not n18970 ; n18970_not
g32350 not n19672 ; n19672_not
g32351 not n19708 ; n19708_not
g32352 not n19771 ; n19771_not
g32353 not n19825 ; n19825_not
g32354 not n19861 ; n19861_not
g32355 not n19933 ; n19933_not
g32356 not n16495 ; n16495_not
g32357 not n16477 ; n16477_not
g32358 not n15874 ; n15874_not
g32359 not n16459 ; n16459_not
g32360 not n15937 ; n15937_not
g32361 not n18619 ; n18619_not
g32362 not n18655 ; n18655_not
g32363 not n18646 ; n18646_not
g32364 not n15973 ; n15973_not
g32365 not n19348 ; n19348_not
g32366 not n18682 ; n18682_not
g32367 not n18691 ; n18691_not
g32368 not n19384 ; n19384_not
g32369 not n16189 ; n16189_not
g32370 not n18727 ; n18727_not
g32371 not n16297 ; n16297_not
g32372 not n18718 ; n18718_not
g32373 not n18754 ; n18754_not
g32374 not n18763 ; n18763_not
g32375 not n19456 ; n19456_not
g32376 not n18790 ; n18790_not
g32377 not n19492 ; n19492_not
g32378 not n18826 ; n18826_not
g32379 not n18835 ; n18835_not
g32380 not n16891 ; n16891_not
g32381 not n14686 ; n14686_not
g32382 not n21868 ; n21868_not
g32383 not n16855 ; n16855_not
g32384 not n16846 ; n16846_not
g32385 not n17476 ; n17476_not
g32386 not n18277 ; n18277_not
g32387 not n17692 ; n17692_not
g32388 not n16819 ; n16819_not
g32389 not n21778 ; n21778_not
g32390 not n17809 ; n17809_not
g32391 not n18349 ; n18349_not
g32392 not n18385 ; n18385_not
g32393 not n16783 ; n16783_not
g32394 not n16774 ; n16774_not
g32395 not n17791 ; n17791_not
g32396 not n17773 ; n17773_not
g32397 not n16738 ; n16738_not
g32398 not n13984 ; n13984_not
g32399 not n16990 ; n16990_not
g32400 not n17953 ; n17953_not
g32401 not n17917 ; n17917_not
g32402 not n14389 ; n14389_not
g32403 not n14497 ; n14497_not
g32404 not n16954 ; n16954_not
g32405 not n14569 ; n14569_not
g32406 not n16963 ; n16963_not
g32407 not n17656 ; n17656_not
g32408 not n21994 ; n21994_not
g32409 not n17584 ; n17584_not
g32410 not n17881 ; n17881_not
g32411 not n21958 ; n21958_not
g32412 not n16927 ; n16927_not
g32413 not n16918 ; n16918_not
g32414 not n17845 ; n17845_not
g32415 not n18097 ; n18097_not
g32416 not n17548 ; n17548_not
g32417 not n16882 ; n16882_not
g32418 not n21886 ; n21886_not
g32419 not n18169 ; n18169_not
g32420 not n17728 ; n17728_not
g32421 not n20779 ; n20779_not
g32422 not n13876 ; n13876_not
g32423 not n17368 ; n17368_not
g32424 not n17737 ; n17737_not
g32425 not n21598 ; n21598_not
g32426 not n20887 ; n20887_not
g32427 not n20878 ; n20878_not
g32428 not n17746 ; n17746_not
g32429 not n13948 ; n13948_not
g32430 not n13399 ; n13399_not
g32431 not n16747 ; n16747_not
g32432 not n20995 ; n20995_not
g32433 not n20959 ; n20959_not
g32434 not n20986 ; n20986_not
g32435 not n23597 ; n23597_not
g32436 not n16964 ; n16964_not
g32437 not n22499 ; n22499_not
g32438 not n19565 ; n19565_not
g32439 not n15974 ; n15974_not
g32440 not n15983 ; n15983_not
g32441 not n15947 ; n15947_not
g32442 not n15938 ; n15938_not
g32443 not n23489 ; n23489_not
g32444 not n24785 ; n24785_not
g32445 not n17657 ; n17657_not
g32446 not n16568 ; n16568_not
g32447 not n19673 ; n19673_not
g32448 not n22868 ; n22868_not
g32449 not n22859 ; n22859_not
g32450 not n19529 ; n19529_not
g32451 not n19664 ; n19664_not
g32452 not n22688 ; n22688_not
g32453 not n22679 ; n22679_not
g32454 not n16928 ; n16928_not
g32455 not n19790 ; n19790_not
g32456 not n19097 ; n19097_not
g32457 not n19637 ; n19637_not
g32458 not n17729 ; n17729_not
g32459 not n16892 ; n16892_not
g32460 not n22796 ; n22796_not
g32461 not n16298 ; n16298_not
g32462 not n22787 ; n22787_not
g32463 not n16856 ; n16856_not
g32464 not n16199 ; n16199_not
g32465 not n16784 ; n16784_not
g32466 not n11969 ; n11969_not
g32467 not n24767 ; n24767_not
g32468 not n16748 ; n16748_not
g32469 not n19709 ; n19709_not
g32470 not n16676 ; n16676_not
g32471 not n17693 ; n17693_not
g32472 not n18548 ; n18548_not
g32473 not n18278 ; n18278_not
g32474 not n18287 ; n18287_not
g32475 not n17882 ; n17882_not
g32476 not n18944 ; n18944_not
g32477 not n23957 ; n23957_not
g32478 not n10898 ; n10898_not
g32479 not n17891 ; n17891_not
g32480 not n18584 ; n18584_not
g32481 not n17297 ; n17297_not
g32482 not n17927 ; n17927_not
g32483 not n18908 ; n18908_not
g32484 not n17918 ; n17918_not
g32485 not n23993 ; n23993_not
g32486 not n18872 ; n18872_not
g32487 not n17954 ; n17954_not
g32488 not n18179 ; n18179_not
g32489 not n17963 ; n17963_not
g32490 not n18656 ; n18656_not
g32491 not n18836 ; n18836_not
g32492 not n10799 ; n10799_not
g32493 not n17990 ; n17990_not
g32494 not n18692 ; n18692_not
g32495 not n17369 ; n17369_not
g32496 not n18728 ; n18728_not
g32497 not n18098 ; n18098_not
g32498 not n18764 ; n18764_not
g32499 not n11897 ; n11897_not
g32500 not n16379 ; n16379_not
g32501 not n19493 ; n19493_not
g32502 not n24578 ; n24578_not
g32503 not n22895 ; n22895_not
g32504 not n23669 ; n23669_not
g32505 not n19457 ; n19457_not
g32506 not n24479 ; n24479_not
g32507 not n17585 ; n17585_not
g32508 not n19385 ; n19385_not
g32509 not n22967 ; n22967_not
g32510 not n22976 ; n22976_not
g32511 not n19349 ; n19349_not
g32512 not n17549 ; n17549_not
g32513 not n23777 ; n23777_not
g32514 not n19277 ; n19277_not
g32515 not n17477 ; n17477_not
g32516 not n23849 ; n23849_not
g32517 not n19169 ; n19169_not
g32518 not n17189 ; n17189_not
g32519 not n18476 ; n18476_not
g32520 not n17819 ; n17819_not
g32521 not n23885 ; n23885_not
g32522 not n17855 ; n17855_not
g32523 not n18359 ; n18359_not
g32524 not n10979 ; n10979_not
g32525 not n18980 ; n18980_not
g32526 not n17846 ; n17846_not
g32527 not n21887 ; n21887_not
g32528 not n15875 ; n15875_not
g32529 not n15857 ; n15857_not
g32530 not n15848 ; n15848_not
g32531 not n12779 ; n12779_not
g32532 not n15884 ; n15884_not
g32533 not n20996 ; n20996_not
g32534 not n12698 ; n12698_not
g32535 not n20888 ; n20888_not
g32536 not n22589 ; n22589_not
g32537 not n13697 ; n13697_not
g32538 not n19970 ; n19970_not
g32539 not n12599 ; n12599_not
g32540 not n19943 ; n19943_not
g32541 not n19934 ; n19934_not
g32542 not n19907 ; n19907_not
g32543 not n19871 ; n19871_not
g32544 not n19862 ; n19862_not
g32545 not n19826 ; n19826_not
g32546 not n19835 ; n19835_not
g32547 not n13868 ; n13868_not
g32548 not n16469 ; n16469_not
g32549 not n15839 ; n15839_not
g32550 not n13769 ; n13769_not
g32551 not n21599 ; n21599_not
g32552 not n13589 ; n13589_not
g32553 not n14948 ; n14948_not
g32554 not n21896 ; n21896_not
g32555 not n14984 ; n14984_not
g32556 not n14399 ; n14399_not
g32557 not n14498 ; n14498_not
g32558 not n14579 ; n14579_not
g32559 not n21959 ; n21959_not
g32560 not n21968 ; n21968_not
g32561 not n12959 ; n12959_not
g32562 not n14876 ; n14876_not
g32563 not n14687 ; n14687_not
g32564 not n15389 ; n15389_not
g32565 not n21995 ; n21995_not
g32566 not n14768 ; n14768_not
g32567 not n15497 ; n15497_not
g32568 not n14696 ; n14696_not
g32569 not n15569 ; n15569_not
g32570 not n12887 ; n12887_not
g32571 not n12878 ; n12878_not
g32572 not n15677 ; n15677_not
g32573 not n21869 ; n21869_not
g32574 not n15749 ; n15749_not
g32575 not n15785 ; n15785_not
g32576 not n14669 ; n14669_not
g32577 not n13949 ; n13949_not
g32578 not n21779 ; n21779_not
g32579 not n21788 ; n21788_not
g32580 not n13877 ; n13877_not
g32581 not n13985 ; n13985_not
g32582 not n16496 ; n16496_not
g32583 not n17964 ; n17964_not
g32584 not n18288 ; n18288_not
g32585 not n23679 ; n23679_not
g32586 not n14769 ; n14769_not
g32587 not n18909 ; n18909_not
g32588 not n13959 ; n13959_not
g32589 not n19395 ; n19395_not
g32590 not n13986 ; n13986_not
g32591 not n24768 ; n24768_not
g32592 not n17379 ; n17379_not
g32593 not n19386 ; n19386_not
g32594 not n18945 ; n18945_not
g32595 not n17586 ; n17586_not
g32596 not n22797 ; n22797_not
g32597 not n18873 ; n18873_not
g32598 not n17298 ; n17298_not
g32599 not n21789 ; n21789_not
g32600 not n16785 ; n16785_not
g32601 not n17667 ; n17667_not
g32602 not n17658 ; n17658_not
g32603 not n15759 ; n15759_not
g32604 not n12969 ; n12969_not
g32605 not n18837 ; n18837_not
g32606 not n19719 ; n19719_not
g32607 not n13878 ; n13878_not
g32608 not n17928 ; n17928_not
g32609 not n14877 ; n14877_not
g32610 not n17694 ; n17694_not
g32611 not n18972 ; n18972_not
g32612 not n16569 ; n16569_not
g32613 not n15399 ; n15399_not
g32614 not n20889 ; n20889_not
g32615 not n19467 ; n19467_not
g32616 not n19458 ; n19458_not
g32617 not n15849 ; n15849_not
g32618 not n15984 ; n15984_not
g32619 not n21897 ; n21897_not
g32620 not n22869 ; n22869_not
g32621 not n17478 ; n17478_not
g32622 not n15948 ; n15948_not
g32623 not n15876 ; n15876_not
g32624 not n17487 ; n17487_not
g32625 not n19746 ; n19746_not
g32626 not n19494 ; n19494_not
g32627 not n16677 ; n16677_not
g32628 not n20997 ; n20997_not
g32629 not n11979 ; n11979_not
g32630 not n17595 ; n17595_not
g32631 not n13995 ; n13995_not
g32632 not n23598 ; n23598_not
g32633 not n17757 ; n17757_not
g32634 not n15678 ; n15678_not
g32635 not n22977 ; n22977_not
g32636 not n18981 ; n18981_not
g32637 not n19575 ; n19575_not
g32638 not n16749 ; n16749_not
g32639 not n21969 ; n21969_not
g32640 not n17559 ; n17559_not
g32641 not n19566 ; n19566_not
g32642 not n15687 ; n15687_not
g32643 not n14697 ; n14697_not
g32644 not n15579 ; n15579_not
g32645 not n19539 ; n19539_not
g32646 not n15498 ; n15498_not
g32647 not n16497 ; n16497_not
g32648 not n17748 ; n17748_not
g32649 not n22689 ; n22689_not
g32650 not n21888 ; n21888_not
g32651 not n18657 ; n18657_not
g32652 not n23859 ; n23859_not
g32653 not n14949 ; n14949_not
g32654 not n19773 ; n19773_not
g32655 not n17856 ; n17856_not
g32656 not n17199 ; n17199_not
g32657 not n16929 ; n16929_not
g32658 not n23778 ; n23778_not
g32659 not n16857 ; n16857_not
g32660 not n12888 ; n12888_not
g32661 not n23787 ; n23787_not
g32662 not n19836 ; n19836_not
g32663 not n24696 ; n24696_not
g32664 not n17766 ; n17766_not
g32665 not n19944 ; n19944_not
g32666 not n18585 ; n18585_not
g32667 not n18549 ; n18549_not
g32668 not n19908 ; n19908_not
g32669 not n19179 ; n19179_not
g32670 not n17775 ; n17775_not
g32671 not n19872 ; n19872_not
g32672 not n19683 ; n19683_not
g32673 not n16893 ; n16893_not
g32674 not n23895 ; n23895_not
g32675 not n23886 ; n23886_not
g32676 not n14985 ; n14985_not
g32677 not n19674 ; n19674_not
g32678 not n19638 ; n19638_not
g32679 not n15786 ; n15786_not
g32680 not n18765 ; n18765_not
g32681 not n13887 ; n13887_not
g32682 not n24597 ; n24597_not
g32683 not n18477 ; n18477_not
g32684 not n23958 ; n23958_not
g32685 not n23967 ; n23967_not
g32686 not n15795 ; n15795_not
g32687 not n19647 ; n19647_not
g32688 not n18729 ; n18729_not
g32689 not n19359 ; n19359_not
g32690 not n16965 ; n16965_not
g32691 not n19791 ; n19791_not
g32692 not n19980 ; n19980_not
g32693 not n17892 ; n17892_not
g32694 not n13779 ; n13779_not
g32695 not n13698 ; n13698_not
g32696 not n11898 ; n11898_not
g32697 not n23994 ; n23994_not
g32698 not n13599 ; n13599_not
g32699 not n24795 ; n24795_not
g32700 not n23499 ; n23499_not
g32701 not n19764 ; n19764_not
g32702 not n18693 ; n18693_not
g32703 not n19287 ; n19287_not
g32704 not n19278 ; n19278_not
g32705 not n23788 ; n23788_not
g32706 not n20998 ; n20998_not
g32707 not n15796 ; n15796_not
g32708 not n16858 ; n16858_not
g32709 not n16867 ; n16867_not
g32710 not n24796 ; n24796_not
g32711 not n18487 ; n18487_not
g32712 not n18478 ; n18478_not
g32713 not n18559 ; n18559_not
g32714 not n16786 ; n16786_not
g32715 not n16687 ; n16687_not
g32716 not n16678 ; n16678_not
g32717 not n14698 ; n14698_not
g32718 not n16795 ; n16795_not
g32719 not n14779 ; n14779_not
g32720 not n13888 ; n13888_not
g32721 not n18289 ; n18289_not
g32722 not n14878 ; n14878_not
g32723 not n23968 ; n23968_not
g32724 not n14887 ; n14887_not
g32725 not n15877 ; n15877_not
g32726 not n22798 ; n22798_not
g32727 not n14959 ; n14959_not
g32728 not n12979 ; n12979_not
g32729 not n20899 ; n20899_not
g32730 not n17488 ; n17488_not
g32731 not n16759 ; n16759_not
g32732 not n14995 ; n14995_not
g32733 not n14986 ; n14986_not
g32734 not n23896 ; n23896_not
g32735 not a[10] ; a[10]_not
g32736 not n16579 ; n16579_not
g32737 not n15688 ; n15688_not
g32738 not n18982 ; n18982_not
g32739 not n18991 ; n18991_not
g32740 not n17767 ; n17767_not
g32741 not n19648 ; n19648_not
g32742 not n18955 ; n18955_not
g32743 not n18946 ; n18946_not
g32744 not n17965 ; n17965_not
g32745 not n18919 ; n18919_not
g32746 not n19576 ; n19576_not
g32747 not n16966 ; n16966_not
g32748 not n18883 ; n18883_not
g32749 not n18874 ; n18874_not
g32750 not n17596 ; n17596_not
g32751 not n18838 ; n18838_not
g32752 not n18847 ; n18847_not
g32753 not n16939 ; n16939_not
g32754 not n19468 ; n19468_not
g32755 not n22978 ; n22978_not
g32756 not n19981 ; n19981_not
g32757 not n17785 ; n17785_not
g32758 not n19945 ; n19945_not
g32759 not n19909 ; n19909_not
g32760 not n24697 ; n24697_not
g32761 not n24679 ; n24679_not
g32762 not n19873 ; n19873_not
g32763 not n13996 ; n13996_not
g32764 not n17857 ; n17857_not
g32765 not n19837 ; n19837_not
g32766 not n19099 ; n19099_not
g32767 not n12889 ; n12889_not
g32768 not n19774 ; n19774_not
g32769 not n17668 ; n17668_not
g32770 not n17893 ; n17893_not
g32771 not n24598 ; n24598_not
g32772 not n17929 ; n17929_not
g32773 not n19684 ; n19684_not
g32774 not n16894 ; n16894_not
g32775 not n18667 ; n18667_not
g32776 not n18694 ; n18694_not
g32777 not n18658 ; n18658_not
g32778 not n15985 ; n15985_not
g32779 not n19396 ; n19396_not
g32780 not n15949 ; n15949_not
g32781 not n19288 ; n19288_not
g32782 not n18739 ; n18739_not
g32783 not n15895 ; n15895_not
g32784 not n21898 ; n21898_not
g32785 not n18766 ; n18766_not
g32786 not n18586 ; n18586_not
g32787 not n18595 ; n18595_not
g32788 not n18775 ; n18775_not
g32789 not n19748 ; n19748_not
g32790 not n18398 ; n18398_not
g32791 not n19757 ; n19757_not
g32792 not n19775 ; n19775_not
g32793 not n14888 ; n14888_not
g32794 not n18668 ; n18668_not
g32795 not n17795 ; n17795_not
g32796 not n17669 ; n17669_not
g32797 not n16868 ; n16868_not
g32798 not n22979 ; n22979_not
g32799 not n22988 ; n22988_not
g32800 not n15986 ; n15986_not
g32801 not n19685 ; n19685_not
g32802 not n17867 ; n17867_not
g32803 not n23789 ; n23789_not
g32804 not a[20] ; a[20]_not
g32805 not n19289 ; n19289_not
g32806 not n17858 ; n17858_not
g32807 not n17894 ; n17894_not
g32808 not n13889 ; n13889_not
g32809 not n21899 ; n21899_not
g32810 not n17786 ; n17786_not
g32811 not n14996 ; n14996_not
g32812 not n18488 ; n18488_not
g32813 not n18596 ; n18596_not
g32814 not n17939 ; n17939_not
g32815 not n13997 ; n13997_not
g32816 not n15995 ; n15995_not
g32817 not n24788 ; n24788_not
g32818 not n17975 ; n17975_not
g32819 not n17966 ; n17966_not
g32820 not n19784 ; n19784_not
g32821 not n23897 ; n23897_not
g32822 not n19739 ; n19739_not
g32823 not n15959 ; n15959_not
g32824 not n19577 ; n19577_not
g32825 not n18884 ; n18884_not
g32826 not n19874 ; n19874_not
g32827 not n17489 ; n17489_not
g32828 not n15689 ; n15689_not
g32829 not n23969 ; n23969_not
g32830 not n19919 ; n19919_not
g32831 not n17597 ; n17597_not
g32832 not n19991 ; n19991_not
g32833 not n19955 ; n19955_not
g32834 not n19946 ; n19946_not
g32835 not n12899 ; n12899_not
g32836 not n18956 ; n18956_not
g32837 not n19469 ; n19469_not
g32838 not n16796 ; n16796_not
g32839 not n18776 ; n18776_not
g32840 not n15797 ; n15797_not
g32841 not n16499 ; n16499_not
g32842 not n16688 ; n16688_not
g32843 not n19649 ; n19649_not
g32844 not n19838 ; n19838_not
g32845 not n19397 ; n19397_not
g32846 not n19847 ; n19847_not
g32847 not n16976 ; n16976_not
g32848 not n18992 ; n18992_not
g32849 not n19982 ; n19982_not
g32850 not n22799 ; n22799_not
g32851 not n18848 ; n18848_not
g32852 not n19883 ; n19883_not
g32853 not n24699 ; n24699_not
g32854 not n13998 ; n13998_not
g32855 not n17787 ; n17787_not
g32856 not n17769 ; n17769_not
g32857 not n17796 ; n17796_not
g32858 not a[30] ; a[30]_not
g32859 not n17598 ; n17598_not
g32860 not n17499 ; n17499_not
g32861 not n16968 ; n16968_not
g32862 not n17976 ; n17976_not
g32863 not n17868 ; n17868_not
g32864 not n14889 ; n14889_not
g32865 not n13899 ; n13899_not
g32866 not n23799 ; n23799_not
g32867 not n17679 ; n17679_not
g32868 not n19398 ; n19398_not
g32869 not n16797 ; n16797_not
g32870 not n16869 ; n16869_not
g32871 not n19992 ; n19992_not
g32872 not n18849 ; n18849_not
g32873 not n19299 ; n19299_not
g32874 not n18885 ; n18885_not
g32875 not n19956 ; n19956_not
g32876 not n22989 ; n22989_not
g32877 not n18957 ; n18957_not
g32878 not n19884 ; n19884_not
g32879 not n18993 ; n18993_not
g32880 not a[12] ; a[12]_not
g32881 not n19848 ; n19848_not
g32882 not n19776 ; n19776_not
g32883 not n15798 ; n15798_not
g32884 not n19749 ; n19749_not
g32885 not n16977 ; n16977_not
g32886 not n19695 ; n19695_not
g32887 not n19686 ; n19686_not
g32888 not n15879 ; n15879_not
g32889 not n18489 ; n18489_not
g32890 not n14997 ; n14997_not
g32891 not n18597 ; n18597_not
g32892 not n19659 ; n19659_not
g32893 not n19578 ; n19578_not
g32894 not n19587 ; n19587_not
g32895 not n23898 ; n23898_not
g32896 not n15996 ; n15996_not
g32897 not n18777 ; n18777_not
g32898 not n18669 ; n18669_not
g32899 not n19479 ; n19479_not
g32900 not n23979 ; n23979_not
g32901 not n16689 ; n16689_not
g32902 not n16879 ; n16879_not
g32903 not a[22] ; a[22]_not
g32904 not n18958 ; n18958_not
g32905 not n18967 ; n18967_not
g32906 not n19588 ; n19588_not
g32907 not n15997 ; n15997_not
g32908 not n17977 ; n17977_not
g32909 not n18778 ; n18778_not
g32910 not n18598 ; n18598_not
g32911 not n15889 ; n15889_not
g32912 not a[40] ; a[40]_not
g32913 not n16978 ; n16978_not
g32914 not n18886 ; n18886_not
g32915 not n16987 ; n16987_not
g32916 not n18679 ; n18679_not
g32917 not n18895 ; n18895_not
g32918 not n18859 ; n18859_not
g32919 not n18787 ; n18787_not
g32920 not n16798 ; n16798_not
g32921 not n16699 ; n16699_not
g32922 not n19993 ; n19993_not
g32923 not n19957 ; n19957_not
g32924 not n14899 ; n14899_not
g32925 not n17797 ; n17797_not
g32926 not n19885 ; n19885_not
g32927 not n19849 ; n19849_not
g32928 not n19795 ; n19795_not
g32929 not n17869 ; n17869_not
g32930 not n18994 ; n18994_not
g32931 not n14998 ; n14998_not
g32932 not n18499 ; n18499_not
g32933 not n19696 ; n19696_not
g32934 not n19777 ; n19777_not
g32935 not n15899 ; n15899_not
g32936 not n15998 ; n15998_not
g32937 not n19994 ; n19994_not
g32938 not n19697 ; n19697_not
g32939 not n19967 ; n19967_not
g32940 not n19859 ; n19859_not
g32941 not n19958 ; n19958_not
g32942 not n16988 ; n16988_not
g32943 not n19895 ; n19895_not
g32944 not n19886 ; n19886_not
g32945 not a[14] ; a[14]_not
g32946 not a[32] ; a[32]_not
g32947 not n19589 ; n19589_not
g32948 not n17798 ; n17798_not
g32949 not a[50] ; a[50]_not
g32950 not n18968 ; n18968_not
g32951 not n18896 ; n18896_not
g32952 not n18788 ; n18788_not
g32953 not n17987 ; n17987_not
g32954 not n17879 ; n17879_not
g32955 not n17978 ; n17978_not
g32956 not n16989 ; n16989_not
g32957 not a[60] ; a[60]_not
g32958 not n19779 ; n19779_not
g32959 not n19599 ; n19599_not
g32960 not a[24] ; a[24]_not
g32961 not n18969 ; n18969_not
g32962 not n19896 ; n19896_not
g32963 not n19698 ; n19698_not
g32964 not n18897 ; n18897_not
g32965 not n19968 ; n19968_not
g32966 not a[42] ; a[42]_not
g32967 not n18789 ; n18789_not
g32968 not n17988 ; n17988_not
g32969 not n18799 ; n18799_not
g32970 not a[34] ; a[34]_not
g32971 not n19969 ; n19969_not
g32972 not n19897 ; n19897_not
g32973 not n19789 ; n19789_not
g32974 not a[52] ; a[52]_not
g32975 not a[70] ; a[70]_not
g32976 not a[16] ; a[16]_not
g32977 not n16999 ; n16999_not
g32978 not n18898 ; n18898_not
g32979 not n17989 ; n17989_not
g32980 not n19979 ; n19979_not
g32981 not n19799 ; n19799_not
g32982 not a[26] ; a[26]_not
g32983 not n19898 ; n19898_not
g32984 not n17999 ; n17999_not
g32985 not a[44] ; a[44]_not
g32986 not a[62] ; a[62]_not
g32987 not a[80] ; a[80]_not
g32988 not a[54] ; a[54]_not
g32989 not a[36] ; a[36]_not
g32990 not a[72] ; a[72]_not
g32991 not a[90] ; a[90]_not
g32992 not a[18] ; a[18]_not
g32993 not a[28] ; a[28]_not
g32994 not a[46] ; a[46]_not
g32995 not a[82] ; a[82]_not
g32996 not a[64] ; a[64]_not
g32997 not a[38] ; a[38]_not
g32998 not a[74] ; a[74]_not
g32999 not a[92] ; a[92]_not
g33000 not a[56] ; a[56]_not
g33001 not a[84] ; a[84]_not
g33002 not a[66] ; a[66]_not
g33003 not a[48] ; a[48]_not
g33004 not a[94] ; a[94]_not
g33005 not a[58] ; a[58]_not
g33006 not a[76] ; a[76]_not
g33007 not a[86] ; a[86]_not
g33008 not a[68] ; a[68]_not
g33009 not a[78] ; a[78]_not
g33010 not a[96] ; a[96]_not
g33011 not a[88] ; a[88]_not
g33012 not a[98] ; a[98]_not
g33013 not a[100] ; a[100]_not
g33014 not a[110] ; a[110]_not
g33015 not a[120] ; a[120]_not
g33016 not a[102] ; a[102]_not
g33017 not a[112] ; a[112]_not
g33018 not a[122] ; a[122]_not
g33019 not a[104] ; a[104]_not
g33020 not a[114] ; a[114]_not
g33021 not a[124] ; a[124]_not
g33022 not a[106] ; a[106]_not
g33023 not a[116] ; a[116]_not
g33024 not a[108] ; a[108]_not
g33025 not a[118] ; a[118]_not
