name div
i a[0]
i a[1]
i a[2]
i a[3]
i a[4]
i a[5]
i a[6]
i a[7]
i a[8]
i a[9]
i a[10]
i a[11]
i a[12]
i a[13]
i a[14]
i a[15]
i a[16]
i a[17]
i a[18]
i a[19]
i a[20]
i a[21]
i a[22]
i a[23]
i a[24]
i a[25]
i a[26]
i a[27]
i a[28]
i a[29]
i a[30]
i a[31]
i a[32]
i a[33]
i a[34]
i a[35]
i a[36]
i a[37]
i a[38]
i a[39]
i a[40]
i a[41]
i a[42]
i a[43]
i a[44]
i a[45]
i a[46]
i a[47]
i a[48]
i a[49]
i a[50]
i a[51]
i a[52]
i a[53]
i a[54]
i a[55]
i a[56]
i a[57]
i a[58]
i a[59]
i a[60]
i a[61]
i a[62]
i a[63]
i b[0]
i b[1]
i b[2]
i b[3]
i b[4]
i b[5]
i b[6]
i b[7]
i b[8]
i b[9]
i b[10]
i b[11]
i b[12]
i b[13]
i b[14]
i b[15]
i b[16]
i b[17]
i b[18]
i b[19]
i b[20]
i b[21]
i b[22]
i b[23]
i b[24]
i b[25]
i b[26]
i b[27]
i b[28]
i b[29]
i b[30]
i b[31]
i b[32]
i b[33]
i b[34]
i b[35]
i b[36]
i b[37]
i b[38]
i b[39]
i b[40]
i b[41]
i b[42]
i b[43]
i b[44]
i b[45]
i b[46]
i b[47]
i b[48]
i b[49]
i b[50]
i b[51]
i b[52]
i b[53]
i b[54]
i b[55]
i b[56]
i b[57]
i b[58]
i b[59]
i b[60]
i b[61]
i b[62]
i b[63]

g1 and a[63]_not b[0] ; n257
g2 and b[0] b[1]_not ; n258
g3 and b[2]_not b[3]_not ; n259
g4 and n258 n259 ; n260
g5 and n257_not n260 ; n261
g6 and b[8]_not b[9]_not ; n262
g7 and b[10]_not b[11]_not ; n263
g8 and n262 n263 ; n264
g9 and b[4]_not b[5]_not ; n265
g10 and b[6]_not b[7]_not ; n266
g11 and n265 n266 ; n267
g12 and n264 n267 ; n268
g13 and b[16]_not b[17]_not ; n269
g14 and b[18]_not b[19]_not ; n270
g15 and n269 n270 ; n271
g16 and b[12]_not b[13]_not ; n272
g17 and b[14]_not b[15]_not ; n273
g18 and n272 n273 ; n274
g19 and n271 n274 ; n275
g20 and n268 n275 ; n276
g21 and n261 n276 ; n277
g22 and b[60]_not b[61]_not ; n278
g23 and b[62]_not b[63]_not ; n279
g24 and n278 n279 ; n280
g25 and b[56]_not b[57]_not ; n281
g26 and b[58]_not b[59]_not ; n282
g27 and n281 n282 ; n283
g28 and b[52]_not b[53]_not ; n284
g29 and b[54]_not b[55]_not ; n285
g30 and n284 n285 ; n286
g31 and n283 n286 ; n287
g32 and n280 n287 ; n288
g33 and b[40]_not b[41]_not ; n289
g34 and b[42]_not b[43]_not ; n290
g35 and n289 n290 ; n291
g36 and b[36]_not b[37]_not ; n292
g37 and b[38]_not b[39]_not ; n293
g38 and n292 n293 ; n294
g39 and n291 n294 ; n295
g40 and b[48]_not b[49]_not ; n296
g41 and b[50]_not b[51]_not ; n297
g42 and n296 n297 ; n298
g43 and b[44]_not b[45]_not ; n299
g44 and b[46]_not b[47]_not ; n300
g45 and n299 n300 ; n301
g46 and n298 n301 ; n302
g47 and n295 n302 ; n303
g48 and b[24]_not b[25]_not ; n304
g49 and b[26]_not b[27]_not ; n305
g50 and n304 n305 ; n306
g51 and b[20]_not b[21]_not ; n307
g52 and b[22]_not b[23]_not ; n308
g53 and n307 n308 ; n309
g54 and n306 n309 ; n310
g55 and b[32]_not b[33]_not ; n311
g56 and b[34]_not b[35]_not ; n312
g57 and n311 n312 ; n313
g58 and b[28]_not b[29]_not ; n314
g59 and b[30]_not b[31]_not ; n315
g60 and n314 n315 ; n316
g61 and n313 n316 ; n317
g62 and n310 n317 ; n318
g63 and n303 n318 ; n319
g64 and n288 n319 ; n320
g65 and n277 n320 ; n321
g66 and a[62]_not b[0] ; n322
g67 and b[1] n322 ; n323
g68 and a[63] n323_not ; n324
g69 and n321_not n324 ; n325
g70 and b[1]_not n322_not ; n326
g71 and n325_not n326_not ; n327
g72 and a[63] n321_not ; n328
g73 and b[1] n322_not ; n329
g74 and b[1]_not n322 ; n330
g75 and n329_not n330_not ; n331
g76 and n259 n267 ; n332
g77 and n264 n274 ; n333
g78 and n332 n333 ; n334
g79 and n331_not n334 ; n335
g80 and n286 n298 ; n336
g81 and n280 n283 ; n337
g82 and n336 n337 ; n338
g83 and n294 n313 ; n339
g84 and n291 n301 ; n340
g85 and n339 n340 ; n341
g86 and n271 n309 ; n342
g87 and n306 n316 ; n343
g88 and n342 n343 ; n344
g89 and n341 n344 ; n345
g90 and n338 n345 ; n346
g91 and n335 n346 ; n347
g92 and n328_not n347 ; n348
g93 and n327_not n348 ; n349
g94 and n333 n342 ; n350
g95 and n332 n350 ; n351
g96 and n323_not n326_not ; n352
g97 and n337 n352 ; n353
g98 and n336 n340 ; n354
g99 and n339 n343 ; n355
g100 and n354 n355 ; n356
g101 and n353 n356 ; n357
g102 and n351 n357 ; n358
g103 and n327_not n358 ; n359
g104 and n328 n359_not ; n360
g105 and n349_not n360_not ; n361
g106 and a[61]_not b[0] ; n362
g107 and b[1] n362 ; n363
g108 and b[21]_not b[22]_not ; n364
g109 and b[23]_not b[24]_not ; n365
g110 and n364 n365 ; n366
g111 and b[17]_not b[18]_not ; n367
g112 and b[19]_not b[20]_not ; n368
g113 and n367 n368 ; n369
g114 and n366 n369 ; n370
g115 and b[29]_not b[30]_not ; n371
g116 and b[31]_not b[32]_not ; n372
g117 and n371 n372 ; n373
g118 and b[25]_not b[26]_not ; n374
g119 and b[27]_not b[28]_not ; n375
g120 and n374 n375 ; n376
g121 and n373 n376 ; n377
g122 and n370 n377 ; n378
g123 and b[5]_not b[6]_not ; n379
g124 and b[7]_not b[8]_not ; n380
g125 and n379 n380 ; n381
g126 and b[0] b[2]_not ; n382
g127 and b[3]_not b[4]_not ; n383
g128 and n382 n383 ; n384
g129 and n381 n384 ; n385
g130 and b[13]_not b[14]_not ; n386
g131 and b[15]_not b[16]_not ; n387
g132 and n386 n387 ; n388
g133 and b[9]_not b[10]_not ; n389
g134 and b[11]_not b[12]_not ; n390
g135 and n389 n390 ; n391
g136 and n388 n391 ; n392
g137 and n385 n392 ; n393
g138 and n378 n393 ; n394
g139 and b[53]_not b[54]_not ; n395
g140 and b[55]_not b[56]_not ; n396
g141 and n395 n396 ; n397
g142 and b[49]_not b[50]_not ; n398
g143 and b[51]_not b[52]_not ; n399
g144 and n398 n399 ; n400
g145 and n397 n400 ; n401
g146 and b[61]_not b[62]_not ; n402
g147 and b[63]_not n402 ; n403
g148 and b[57]_not b[58]_not ; n404
g149 and b[59]_not b[60]_not ; n405
g150 and n404 n405 ; n406
g151 and n403 n406 ; n407
g152 and n401 n407 ; n408
g153 and b[37]_not b[38]_not ; n409
g154 and b[39]_not b[40]_not ; n410
g155 and n409 n410 ; n411
g156 and b[33]_not b[34]_not ; n412
g157 and b[35]_not b[36]_not ; n413
g158 and n412 n413 ; n414
g159 and n411 n414 ; n415
g160 and b[45]_not b[46]_not ; n416
g161 and b[47]_not b[48]_not ; n417
g162 and n416 n417 ; n418
g163 and b[41]_not b[42]_not ; n419
g164 and b[43]_not b[44]_not ; n420
g165 and n419 n420 ; n421
g166 and n418 n421 ; n422
g167 and n415 n422 ; n423
g168 and n408 n423 ; n424
g169 and n394 n424 ; n425
g170 and n327_not n425 ; n426
g171 and a[62] n426_not ; n427
g172 and n259 n322 ; n428
g173 and n267 n428 ; n429
g174 and n333 n429 ; n430
g175 and n344 n430 ; n431
g176 and n338 n341 ; n432
g177 and n431 n432 ; n433
g178 and n327_not n433 ; n434
g179 and n427_not n434_not ; n435
g180 and n363_not n435_not ; n436
g181 and b[1]_not n362_not ; n437
g182 and n436_not n437_not ; n438
g183 and b[2] n349_not ; n439
g184 and n360_not n439 ; n440
g185 and b[2]_not n361_not ; n441
g186 and n440_not n441_not ; n442
g187 and n438 n442_not ; n443
g188 and b[2]_not n443_not ; n444
g189 and n438_not n440_not ; n445
g190 and n441_not n445_not ; n446
g191 and n381 n383 ; n447
g192 and n392 n447 ; n448
g193 and n378 n448 ; n449
g194 and n424 n449 ; n450
g195 and n446_not n450 ; quotient[61]
g196 and n444_not quotient[61] ; n452
g197 and n361_not n452_not ; n453
g198 and n445_not n450 ; n454
g199 and n443_not n454 ; n455
g200 and n446_not n455 ; n456
g201 and b[3] n456_not ; n457
g202 and n453_not n457 ; n458
g203 and n370 n392 ; n459
g204 and n447 n459 ; n460
g205 and n363_not n437_not ; n461
g206 and n407 n461 ; n462
g207 and n401 n422 ; n463
g208 and n377 n415 ; n464
g209 and n463 n464 ; n465
g210 and n462 n465 ; n466
g211 and n460 n466 ; n467
g212 and n446_not n467 ; n468
g213 and n435_not n468_not ; n469
g214 and b[1] n362_not ; n470
g215 and b[1]_not n362 ; n471
g216 and n470_not n471_not ; n472
g217 and n448 n472_not ; n473
g218 and n378 n423 ; n474
g219 and n408 n474 ; n475
g220 and n473 n475 ; n476
g221 and n434_not n476 ; n477
g222 and n427_not n477 ; n478
g223 and n446_not n478 ; n479
g224 and n469_not n479_not ; n480
g225 and b[2]_not n480_not ; n481
g226 and b[2] n479_not ; n482
g227 and n469_not n482 ; n483
g228 and b[0] b[3]_not ; n484
g229 and n267 n484 ; n485
g230 and n333 n485 ; n486
g231 and n344 n486 ; n487
g232 and n432 n487 ; n488
g233 and n446_not n488 ; n489
g234 and a[61] n489_not ; n490
g235 and n362 n383 ; n491
g236 and n381 n491 ; n492
g237 and n392 n492 ; n493
g238 and n378 n493 ; n494
g239 and n424 n494 ; n495
g240 and n446_not n495 ; n496
g241 and n490_not n496_not ; n497
g242 and a[60]_not b[0] ; n498
g243 and b[1] n498 ; n499
g244 and n497_not n499_not ; n500
g245 and b[1]_not n498_not ; n501
g246 and n500_not n501_not ; n502
g247 and n483_not n502_not ; n503
g248 and n481_not n503_not ; n504
g249 and n458_not n504_not ; n505
g250 and n453_not n456_not ; n506
g251 and b[3]_not n506_not ; n507
g252 and n505_not n507_not ; n508
g253 and n458_not n507_not ; n509
g254 and n504_not n509 ; n510
g255 and n276 n318 ; n511
g256 and n288 n303 ; n512
g257 and n511 n512 ; n513
g258 and n504 n509_not ; n514
g259 and n513 n514_not ; n515
g260 and n510_not n515 ; n516
g261 and n508_not n516 ; n517
g262 and n508_not n513 ; quotient[60]
g263 and n506_not quotient[60]_not ; n519
g264 and b[4] n519_not ; n520
g265 and n517_not n520 ; n521
g266 and n481_not n483_not ; n522
g267 and n502 n522_not ; n523
g268 and n503_not n513 ; n524
g269 and n523_not n524 ; n525
g270 and n508_not n525 ; n526
g271 and b[2]_not n523_not ; n527
g272 and n513 n527_not ; n528
g273 and n508_not n528 ; n529
g274 and n480_not n529_not ; n530
g275 and n526_not n530_not ; n531
g276 and b[3]_not n531_not ; n532
g277 and b[3] n526_not ; n533
g278 and n530_not n533 ; n534
g279 and n275 n310 ; n535
g280 and n268 n535 ; n536
g281 and n280 n499_not ; n537
g282 and n501_not n537 ; n538
g283 and n287 n302 ; n539
g284 and n295 n317 ; n540
g285 and n539 n540 ; n541
g286 and n538 n541 ; n542
g287 and n536 n542 ; n543
g288 and n508_not n543 ; n544
g289 and n497_not n544_not ; n545
g290 and b[1] n498_not ; n546
g291 and b[1]_not n498 ; n547
g292 and n546_not n547_not ; n548
g293 and n276 n548_not ; n549
g294 and n320 n549 ; n550
g295 and n496_not n550 ; n551
g296 and n490_not n551 ; n552
g297 and n508_not n552 ; n553
g298 and n545_not n553_not ; n554
g299 and b[2]_not n554_not ; n555
g300 and b[2] n553_not ; n556
g301 and n545_not n556 ; n557
g302 and a[59]_not b[0] ; n558
g303 and b[1] n558 ; n559
g304 and b[0] b[4]_not ; n560
g305 and n381 n560 ; n561
g306 and n392 n561 ; n562
g307 and n378 n562 ; n563
g308 and n424 n563 ; n564
g309 and n508_not n564 ; n565
g310 and a[60] n565_not ; n566
g311 and n267 n498 ; n567
g312 and n333 n567 ; n568
g313 and n344 n568 ; n569
g314 and n432 n569 ; n570
g315 and n508_not n570 ; n571
g316 and n566_not n571_not ; n572
g317 and n559_not n572_not ; n573
g318 and b[1]_not n558_not ; n574
g319 and n573_not n574_not ; n575
g320 and n557_not n575_not ; n576
g321 and n555_not n576_not ; n577
g322 and n534_not n577_not ; n578
g323 and n532_not n578_not ; n579
g324 and n521_not n579_not ; n580
g325 and n517_not n519_not ; n581
g326 and b[4]_not n581_not ; n582
g327 and n580_not n582_not ; n583
g328 and n532_not n534_not ; n584
g329 and n555_not n584_not ; n585
g330 and n576_not n585 ; n586
g331 and n366 n376 ; n587
g332 and n373 n414 ; n588
g333 and n587 n588 ; n589
g334 and n381 n391 ; n590
g335 and n369 n388 ; n591
g336 and n590 n591 ; n592
g337 and n589 n592 ; n593
g338 and n397 n406 ; n594
g339 and n403 n594 ; n595
g340 and n411 n421 ; n596
g341 and n400 n418 ; n597
g342 and n596 n597 ; n598
g343 and n595 n598 ; n599
g344 and n593 n599 ; n600
g345 and n586_not n600 ; n601
g346 and n578_not n601 ; n602
g347 and n583_not n602 ; n603
g348 and b[3]_not n586_not ; n604
g349 and n600 n604_not ; n605
g350 and n583_not n605 ; n606
g351 and n531_not n606_not ; n607
g352 and n603_not n607_not ; n608
g353 and b[4] n608_not ; n609
g354 and b[4]_not n603_not ; n610
g355 and n607_not n610 ; n611
g356 and n609_not n611_not ; n612
g357 and n555_not n557_not ; n613
g358 and n575 n613_not ; n614
g359 and n576_not n600 ; n615
g360 and n614_not n615 ; n616
g361 and n583_not n616 ; n617
g362 and b[2]_not n614_not ; n618
g363 and n600 n618_not ; n619
g364 and n583_not n619 ; n620
g365 and n554_not n620_not ; n621
g366 and n617_not n621_not ; n622
g367 and b[3] n622_not ; n623
g368 and b[3]_not n617_not ; n624
g369 and n621_not n624 ; n625
g370 and n623_not n625_not ; n626
g371 and n587 n591 ; n627
g372 and n590 n627 ; n628
g373 and n403 n559_not ; n629
g374 and n574_not n629 ; n630
g375 and n594 n597 ; n631
g376 and n588 n596 ; n632
g377 and n631 n632 ; n633
g378 and n630 n633 ; n634
g379 and n628 n634 ; n635
g380 and n583_not n635 ; n636
g381 and n572_not n636_not ; n637
g382 and b[1] n558_not ; n638
g383 and b[1]_not n558 ; n639
g384 and n638_not n639_not ; n640
g385 and n592 n640_not ; n641
g386 and n589 n598 ; n642
g387 and n595 n642 ; n643
g388 and n641 n643 ; n644
g389 and n571_not n644 ; n645
g390 and n566_not n645 ; n646
g391 and n583_not n646 ; n647
g392 and n637_not n647_not ; n648
g393 and b[2]_not n648_not ; n649
g394 and b[0] b[5]_not ; n650
g395 and n266 n650 ; n651
g396 and n264 n651 ; n652
g397 and n275 n652 ; n653
g398 and n318 n653 ; n654
g399 and n512 n654 ; n655
g400 and n583_not n655 ; n656
g401 and a[59] n656_not ; n657
g402 and n381 n558 ; n658
g403 and n392 n658 ; n659
g404 and n378 n659 ; n660
g405 and n424 n660 ; n661
g406 and n583_not n661 ; n662
g407 and n657_not n662_not ; n663
g408 and b[1] n663_not ; n664
g409 and b[1]_not n662_not ; n665
g410 and n657_not n665 ; n666
g411 and n664_not n666_not ; n667
g412 and a[58]_not b[0] ; n668
g413 and n667_not n668_not ; n669
g414 and b[1]_not n663_not ; n670
g415 and n669_not n670_not ; n671
g416 and b[2] n647_not ; n672
g417 and n637_not n672 ; n673
g418 and n649_not n673_not ; n674
g419 and n671_not n674 ; n675
g420 and n649_not n675_not ; n676
g421 and n626_not n676_not ; n677
g422 and b[3]_not n622_not ; n678
g423 and n677_not n678_not ; n679
g424 and n612_not n679_not ; n680
g425 and b[4]_not n608_not ; n681
g426 and n680_not n681_not ; n682
g427 and n521_not n582_not ; n683
g428 and n532_not n683_not ; n684
g429 and n578_not n684 ; n685
g430 and n600 n685_not ; n686
g431 and n580_not n686 ; n687
g432 and n583_not n687 ; n688
g433 and b[4]_not n685_not ; n689
g434 and n600 n689_not ; n690
g435 and n583_not n690 ; n691
g436 and n581_not n691_not ; n692
g437 and n688_not n692_not ; n693
g438 and b[5] n693_not ; n694
g439 and b[5]_not n688_not ; n695
g440 and n692_not n695 ; n696
g441 and n694_not n696_not ; n697
g442 and n264 n266 ; n698
g443 and n275 n698 ; n699
g444 and n318 n699 ; n700
g445 and n512 n700 ; n701
g446 and n697_not n701 ; n702
g447 and n682_not n702 ; n703
g448 and n600 n693_not ; n704
g449 and n703_not n704_not ; quotient[58]
g450 and n612 n678_not ; n706
g451 and n677_not n706 ; n707
g452 and n680_not n707_not ; n708
g453 and quotient[58] n708 ; n709
g454 and n608_not n704_not ; n710
g455 and n703_not n710 ; n711
g456 and n709_not n711_not ; n712
g457 and n682_not n697_not ; n713
g458 and n681_not n697 ; n714
g459 and n680_not n714 ; n715
g460 and n713_not n715_not ; n716
g461 and quotient[58] n716 ; n717
g462 and n693_not n704_not ; n718
g463 and n703_not n718 ; n719
g464 and n717_not n719_not ; n720
g465 and b[6]_not n720_not ; n721
g466 and b[5]_not n712_not ; n722
g467 and n626 n649_not ; n723
g468 and n675_not n723 ; n724
g469 and n677_not n724_not ; n725
g470 and quotient[58] n725 ; n726
g471 and n622_not n704_not ; n727
g472 and n703_not n727 ; n728
g473 and n726_not n728_not ; n729
g474 and b[4]_not n729_not ; n730
g475 and n670_not n674 ; n731
g476 and n669_not n731 ; n732
g477 and n671_not n674_not ; n733
g478 and n732_not n733_not ; n734
g479 and quotient[58] n734_not ; n735
g480 and n648_not n704_not ; n736
g481 and n703_not n736 ; n737
g482 and n735_not n737_not ; n738
g483 and b[3]_not n738_not ; n739
g484 and n666_not n668 ; n740
g485 and n664_not n740 ; n741
g486 and n669_not n741_not ; n742
g487 and quotient[58] n742 ; n743
g488 and n663_not n704_not ; n744
g489 and n703_not n744 ; n745
g490 and n743_not n745_not ; n746
g491 and b[2]_not n746_not ; n747
g492 and b[0] quotient[58] ; n748
g493 and a[58] n748_not ; n749
g494 and n668 quotient[58] ; n750
g495 and n749_not n750_not ; n751
g496 and b[1] n751_not ; n752
g497 and b[1]_not n750_not ; n753
g498 and n749_not n753 ; n754
g499 and n752_not n754_not ; n755
g500 and a[57]_not b[0] ; n756
g501 and n755_not n756_not ; n757
g502 and b[1]_not n751_not ; n758
g503 and n757_not n758_not ; n759
g504 and b[2] n745_not ; n760
g505 and n743_not n760 ; n761
g506 and n747_not n761_not ; n762
g507 and n759_not n762 ; n763
g508 and n747_not n763_not ; n764
g509 and b[3] n737_not ; n765
g510 and n735_not n765 ; n766
g511 and n739_not n766_not ; n767
g512 and n764_not n767 ; n768
g513 and n739_not n768_not ; n769
g514 and b[4] n728_not ; n770
g515 and n726_not n770 ; n771
g516 and n730_not n771_not ; n772
g517 and n769_not n772 ; n773
g518 and n730_not n773_not ; n774
g519 and b[5] n711_not ; n775
g520 and n709_not n775 ; n776
g521 and n722_not n776_not ; n777
g522 and n774_not n777 ; n778
g523 and n722_not n778_not ; n779
g524 and b[6] n719_not ; n780
g525 and n717_not n780 ; n781
g526 and n721_not n781_not ; n782
g527 and n779_not n782 ; n783
g528 and n721_not n783_not ; n784
g529 and n380 n391 ; n785
g530 and n591 n785 ; n786
g531 and n589 n786 ; n787
g532 and n599 n787 ; n788
g533 and n784_not n788 ; quotient[57]
g534 and n712_not quotient[57]_not ; n790
g535 and n730_not n777 ; n791
g536 and n773_not n791 ; n792
g537 and n774_not n777_not ; n793
g538 and n792_not n793_not ; n794
g539 and n788 n794_not ; n795
g540 and n784_not n795 ; n796
g541 and n790_not n796_not ; n797
g542 and n720_not quotient[57]_not ; n798
g543 and n722_not n782 ; n799
g544 and n778_not n799 ; n800
g545 and n779_not n782_not ; n801
g546 and n800_not n801_not ; n802
g547 and quotient[57] n802_not ; n803
g548 and n798_not n803_not ; n804
g549 and b[7]_not n804_not ; n805
g550 and b[6]_not n797_not ; n806
g551 and n729_not quotient[57]_not ; n807
g552 and n739_not n772 ; n808
g553 and n768_not n808 ; n809
g554 and n769_not n772_not ; n810
g555 and n809_not n810_not ; n811
g556 and n788 n811_not ; n812
g557 and n784_not n812 ; n813
g558 and n807_not n813_not ; n814
g559 and b[5]_not n814_not ; n815
g560 and n738_not quotient[57]_not ; n816
g561 and n747_not n767 ; n817
g562 and n763_not n817 ; n818
g563 and n764_not n767_not ; n819
g564 and n818_not n819_not ; n820
g565 and n788 n820_not ; n821
g566 and n784_not n821 ; n822
g567 and n816_not n822_not ; n823
g568 and b[4]_not n823_not ; n824
g569 and n746_not quotient[57]_not ; n825
g570 and n758_not n762 ; n826
g571 and n757_not n826 ; n827
g572 and n759_not n762_not ; n828
g573 and n827_not n828_not ; n829
g574 and n788 n829_not ; n830
g575 and n784_not n830 ; n831
g576 and n825_not n831_not ; n832
g577 and b[3]_not n832_not ; n833
g578 and n751_not quotient[57]_not ; n834
g579 and n754_not n756 ; n835
g580 and n752_not n835 ; n836
g581 and n788 n836_not ; n837
g582 and n757_not n837 ; n838
g583 and n784_not n838 ; n839
g584 and n834_not n839_not ; n840
g585 and b[2]_not n840_not ; n841
g586 and b[0] b[7]_not ; n842
g587 and n264 n842 ; n843
g588 and n275 n843 ; n844
g589 and n318 n844 ; n845
g590 and n512 n845 ; n846
g591 and n784_not n846 ; n847
g592 and a[57] n847_not ; n848
g593 and n380 n756 ; n849
g594 and n391 n849 ; n850
g595 and n591 n850 ; n851
g596 and n589 n851 ; n852
g597 and n599 n852 ; n853
g598 and n784_not n853 ; n854
g599 and n848_not n854_not ; n855
g600 and b[1] n855_not ; n856
g601 and b[1]_not n854_not ; n857
g602 and n848_not n857 ; n858
g603 and n856_not n858_not ; n859
g604 and a[56]_not b[0] ; n860
g605 and n859_not n860_not ; n861
g606 and b[1]_not n855_not ; n862
g607 and n861_not n862_not ; n863
g608 and b[2] n839_not ; n864
g609 and n834_not n864 ; n865
g610 and n841_not n865_not ; n866
g611 and n863_not n866 ; n867
g612 and n841_not n867_not ; n868
g613 and b[3] n831_not ; n869
g614 and n825_not n869 ; n870
g615 and n833_not n870_not ; n871
g616 and n868_not n871 ; n872
g617 and n833_not n872_not ; n873
g618 and b[4] n822_not ; n874
g619 and n816_not n874 ; n875
g620 and n824_not n875_not ; n876
g621 and n873_not n876 ; n877
g622 and n824_not n877_not ; n878
g623 and b[5] n813_not ; n879
g624 and n807_not n879 ; n880
g625 and n815_not n880_not ; n881
g626 and n878_not n881 ; n882
g627 and n815_not n882_not ; n883
g628 and b[6] n796_not ; n884
g629 and n790_not n884 ; n885
g630 and n806_not n885_not ; n886
g631 and n883_not n886 ; n887
g632 and n806_not n887_not ; n888
g633 and b[7] n798_not ; n889
g634 and n803_not n889 ; n890
g635 and n805_not n890_not ; n891
g636 and n888_not n891 ; n892
g637 and n805_not n892_not ; n893
g638 and n333 n344 ; n894
g639 and n432 n894 ; n895
g640 and n893_not n895 ; quotient[56]
g641 and n797_not quotient[56]_not ; n897
g642 and n815_not n886 ; n898
g643 and n882_not n898 ; n899
g644 and n883_not n886_not ; n900
g645 and n899_not n900_not ; n901
g646 and n895 n901_not ; n902
g647 and n893_not n902 ; n903
g648 and n897_not n903_not ; n904
g649 and b[7]_not n904_not ; n905
g650 and n814_not quotient[56]_not ; n906
g651 and n824_not n881 ; n907
g652 and n877_not n907 ; n908
g653 and n878_not n881_not ; n909
g654 and n908_not n909_not ; n910
g655 and n895 n910_not ; n911
g656 and n893_not n911 ; n912
g657 and n906_not n912_not ; n913
g658 and b[6]_not n913_not ; n914
g659 and n823_not quotient[56]_not ; n915
g660 and n833_not n876 ; n916
g661 and n872_not n916 ; n917
g662 and n873_not n876_not ; n918
g663 and n917_not n918_not ; n919
g664 and n895 n919_not ; n920
g665 and n893_not n920 ; n921
g666 and n915_not n921_not ; n922
g667 and b[5]_not n922_not ; n923
g668 and n832_not quotient[56]_not ; n924
g669 and n841_not n871 ; n925
g670 and n867_not n925 ; n926
g671 and n868_not n871_not ; n927
g672 and n926_not n927_not ; n928
g673 and n895 n928_not ; n929
g674 and n893_not n929 ; n930
g675 and n924_not n930_not ; n931
g676 and b[4]_not n931_not ; n932
g677 and n840_not quotient[56]_not ; n933
g678 and n862_not n866 ; n934
g679 and n861_not n934 ; n935
g680 and n863_not n866_not ; n936
g681 and n935_not n936_not ; n937
g682 and n895 n937_not ; n938
g683 and n893_not n938 ; n939
g684 and n933_not n939_not ; n940
g685 and b[3]_not n940_not ; n941
g686 and n855_not quotient[56]_not ; n942
g687 and n858_not n860 ; n943
g688 and n856_not n943 ; n944
g689 and n895 n944_not ; n945
g690 and n861_not n945 ; n946
g691 and n893_not n946 ; n947
g692 and n942_not n947_not ; n948
g693 and b[2]_not n948_not ; n949
g694 and b[0] b[8]_not ; n950
g695 and n391 n950 ; n951
g696 and n591 n951 ; n952
g697 and n589 n952 ; n953
g698 and n599 n953 ; n954
g699 and n893_not n954 ; n955
g700 and a[56] n955_not ; n956
g701 and n264 n860 ; n957
g702 and n275 n957 ; n958
g703 and n318 n958 ; n959
g704 and n512 n959 ; n960
g705 and n893_not n960 ; n961
g706 and n956_not n961_not ; n962
g707 and b[1] n962_not ; n963
g708 and b[1]_not n961_not ; n964
g709 and n956_not n964 ; n965
g710 and n963_not n965_not ; n966
g711 and a[55]_not b[0] ; n967
g712 and n966_not n967_not ; n968
g713 and b[1]_not n962_not ; n969
g714 and n968_not n969_not ; n970
g715 and b[2] n947_not ; n971
g716 and n942_not n971 ; n972
g717 and n949_not n972_not ; n973
g718 and n970_not n973 ; n974
g719 and n949_not n974_not ; n975
g720 and b[3] n939_not ; n976
g721 and n933_not n976 ; n977
g722 and n941_not n977_not ; n978
g723 and n975_not n978 ; n979
g724 and n941_not n979_not ; n980
g725 and b[4] n930_not ; n981
g726 and n924_not n981 ; n982
g727 and n932_not n982_not ; n983
g728 and n980_not n983 ; n984
g729 and n932_not n984_not ; n985
g730 and b[5] n921_not ; n986
g731 and n915_not n986 ; n987
g732 and n923_not n987_not ; n988
g733 and n985_not n988 ; n989
g734 and n923_not n989_not ; n990
g735 and b[6] n912_not ; n991
g736 and n906_not n991 ; n992
g737 and n914_not n992_not ; n993
g738 and n990_not n993 ; n994
g739 and n914_not n994_not ; n995
g740 and b[7] n903_not ; n996
g741 and n897_not n996 ; n997
g742 and n905_not n997_not ; n998
g743 and n995_not n998 ; n999
g744 and n905_not n999_not ; n1000
g745 and n804_not quotient[56]_not ; n1001
g746 and n806_not n891 ; n1002
g747 and n887_not n1002 ; n1003
g748 and n888_not n891_not ; n1004
g749 and n1003_not n1004_not ; n1005
g750 and quotient[56] n1005_not ; n1006
g751 and n1001_not n1006_not ; n1007
g752 and b[8]_not n1007_not ; n1008
g753 and b[8] n1001_not ; n1009
g754 and n1006_not n1009 ; n1010
g755 and n378 n392 ; n1011
g756 and n424 n1011 ; n1012
g757 and n1010_not n1012 ; n1013
g758 and n1008_not n1013 ; n1014
g759 and n1000_not n1014 ; n1015
g760 and n895 n1007_not ; n1016
g761 and n1015_not n1016_not ; quotient[55]
g762 and n914_not n998 ; n1018
g763 and n994_not n1018 ; n1019
g764 and n995_not n998_not ; n1020
g765 and n1019_not n1020_not ; n1021
g766 and quotient[55] n1021_not ; n1022
g767 and n904_not n1016_not ; n1023
g768 and n1015_not n1023 ; n1024
g769 and n1022_not n1024_not ; n1025
g770 and n905_not n1010_not ; n1026
g771 and n1008_not n1026 ; n1027
g772 and n999_not n1027 ; n1028
g773 and n1008_not n1010_not ; n1029
g774 and n1000_not n1029_not ; n1030
g775 and n1028_not n1030_not ; n1031
g776 and quotient[55] n1031_not ; n1032
g777 and n1007_not n1016_not ; n1033
g778 and n1015_not n1033 ; n1034
g779 and n1032_not n1034_not ; n1035
g780 and b[9]_not n1035_not ; n1036
g781 and b[8]_not n1025_not ; n1037
g782 and n923_not n993 ; n1038
g783 and n989_not n1038 ; n1039
g784 and n990_not n993_not ; n1040
g785 and n1039_not n1040_not ; n1041
g786 and quotient[55] n1041_not ; n1042
g787 and n913_not n1016_not ; n1043
g788 and n1015_not n1043 ; n1044
g789 and n1042_not n1044_not ; n1045
g790 and b[7]_not n1045_not ; n1046
g791 and n932_not n988 ; n1047
g792 and n984_not n1047 ; n1048
g793 and n985_not n988_not ; n1049
g794 and n1048_not n1049_not ; n1050
g795 and quotient[55] n1050_not ; n1051
g796 and n922_not n1016_not ; n1052
g797 and n1015_not n1052 ; n1053
g798 and n1051_not n1053_not ; n1054
g799 and b[6]_not n1054_not ; n1055
g800 and n941_not n983 ; n1056
g801 and n979_not n1056 ; n1057
g802 and n980_not n983_not ; n1058
g803 and n1057_not n1058_not ; n1059
g804 and quotient[55] n1059_not ; n1060
g805 and n931_not n1016_not ; n1061
g806 and n1015_not n1061 ; n1062
g807 and n1060_not n1062_not ; n1063
g808 and b[5]_not n1063_not ; n1064
g809 and n949_not n978 ; n1065
g810 and n974_not n1065 ; n1066
g811 and n975_not n978_not ; n1067
g812 and n1066_not n1067_not ; n1068
g813 and quotient[55] n1068_not ; n1069
g814 and n940_not n1016_not ; n1070
g815 and n1015_not n1070 ; n1071
g816 and n1069_not n1071_not ; n1072
g817 and b[4]_not n1072_not ; n1073
g818 and n969_not n973 ; n1074
g819 and n968_not n1074 ; n1075
g820 and n970_not n973_not ; n1076
g821 and n1075_not n1076_not ; n1077
g822 and quotient[55] n1077_not ; n1078
g823 and n948_not n1016_not ; n1079
g824 and n1015_not n1079 ; n1080
g825 and n1078_not n1080_not ; n1081
g826 and b[3]_not n1081_not ; n1082
g827 and n965_not n967 ; n1083
g828 and n963_not n1083 ; n1084
g829 and n968_not n1084_not ; n1085
g830 and quotient[55] n1085 ; n1086
g831 and n962_not n1016_not ; n1087
g832 and n1015_not n1087 ; n1088
g833 and n1086_not n1088_not ; n1089
g834 and b[2]_not n1089_not ; n1090
g835 and b[0] quotient[55] ; n1091
g836 and a[55] n1091_not ; n1092
g837 and n967 quotient[55] ; n1093
g838 and n1092_not n1093_not ; n1094
g839 and b[1] n1094_not ; n1095
g840 and b[1]_not n1093_not ; n1096
g841 and n1092_not n1096 ; n1097
g842 and n1095_not n1097_not ; n1098
g843 and a[54]_not b[0] ; n1099
g844 and n1098_not n1099_not ; n1100
g845 and b[1]_not n1094_not ; n1101
g846 and n1100_not n1101_not ; n1102
g847 and b[2] n1088_not ; n1103
g848 and n1086_not n1103 ; n1104
g849 and n1090_not n1104_not ; n1105
g850 and n1102_not n1105 ; n1106
g851 and n1090_not n1106_not ; n1107
g852 and b[3] n1080_not ; n1108
g853 and n1078_not n1108 ; n1109
g854 and n1082_not n1109_not ; n1110
g855 and n1107_not n1110 ; n1111
g856 and n1082_not n1111_not ; n1112
g857 and b[4] n1071_not ; n1113
g858 and n1069_not n1113 ; n1114
g859 and n1073_not n1114_not ; n1115
g860 and n1112_not n1115 ; n1116
g861 and n1073_not n1116_not ; n1117
g862 and b[5] n1062_not ; n1118
g863 and n1060_not n1118 ; n1119
g864 and n1064_not n1119_not ; n1120
g865 and n1117_not n1120 ; n1121
g866 and n1064_not n1121_not ; n1122
g867 and b[6] n1053_not ; n1123
g868 and n1051_not n1123 ; n1124
g869 and n1055_not n1124_not ; n1125
g870 and n1122_not n1125 ; n1126
g871 and n1055_not n1126_not ; n1127
g872 and b[7] n1044_not ; n1128
g873 and n1042_not n1128 ; n1129
g874 and n1046_not n1129_not ; n1130
g875 and n1127_not n1130 ; n1131
g876 and n1046_not n1131_not ; n1132
g877 and b[8] n1024_not ; n1133
g878 and n1022_not n1133 ; n1134
g879 and n1037_not n1134_not ; n1135
g880 and n1132_not n1135 ; n1136
g881 and n1037_not n1136_not ; n1137
g882 and b[9] n1034_not ; n1138
g883 and n1032_not n1138 ; n1139
g884 and n1036_not n1139_not ; n1140
g885 and n1137_not n1140 ; n1141
g886 and n1036_not n1141_not ; n1142
g887 and n263 n274 ; n1143
g888 and n344 n1143 ; n1144
g889 and n432 n1144 ; n1145
g890 and n1142_not n1145 ; quotient[54]
g891 and n1025_not quotient[54]_not ; n1147
g892 and n1046_not n1135 ; n1148
g893 and n1131_not n1148 ; n1149
g894 and n1132_not n1135_not ; n1150
g895 and n1149_not n1150_not ; n1151
g896 and n1145 n1151_not ; n1152
g897 and n1142_not n1152 ; n1153
g898 and n1147_not n1153_not ; n1154
g899 and n1035_not quotient[54]_not ; n1155
g900 and n1037_not n1140 ; n1156
g901 and n1136_not n1156 ; n1157
g902 and n1137_not n1140_not ; n1158
g903 and n1157_not n1158_not ; n1159
g904 and quotient[54] n1159_not ; n1160
g905 and n1155_not n1160_not ; n1161
g906 and b[10]_not n1161_not ; n1162
g907 and b[9]_not n1154_not ; n1163
g908 and n1045_not quotient[54]_not ; n1164
g909 and n1055_not n1130 ; n1165
g910 and n1126_not n1165 ; n1166
g911 and n1127_not n1130_not ; n1167
g912 and n1166_not n1167_not ; n1168
g913 and n1145 n1168_not ; n1169
g914 and n1142_not n1169 ; n1170
g915 and n1164_not n1170_not ; n1171
g916 and b[8]_not n1171_not ; n1172
g917 and n1054_not quotient[54]_not ; n1173
g918 and n1064_not n1125 ; n1174
g919 and n1121_not n1174 ; n1175
g920 and n1122_not n1125_not ; n1176
g921 and n1175_not n1176_not ; n1177
g922 and n1145 n1177_not ; n1178
g923 and n1142_not n1178 ; n1179
g924 and n1173_not n1179_not ; n1180
g925 and b[7]_not n1180_not ; n1181
g926 and n1063_not quotient[54]_not ; n1182
g927 and n1073_not n1120 ; n1183
g928 and n1116_not n1183 ; n1184
g929 and n1117_not n1120_not ; n1185
g930 and n1184_not n1185_not ; n1186
g931 and n1145 n1186_not ; n1187
g932 and n1142_not n1187 ; n1188
g933 and n1182_not n1188_not ; n1189
g934 and b[6]_not n1189_not ; n1190
g935 and n1072_not quotient[54]_not ; n1191
g936 and n1082_not n1115 ; n1192
g937 and n1111_not n1192 ; n1193
g938 and n1112_not n1115_not ; n1194
g939 and n1193_not n1194_not ; n1195
g940 and n1145 n1195_not ; n1196
g941 and n1142_not n1196 ; n1197
g942 and n1191_not n1197_not ; n1198
g943 and b[5]_not n1198_not ; n1199
g944 and n1081_not quotient[54]_not ; n1200
g945 and n1090_not n1110 ; n1201
g946 and n1106_not n1201 ; n1202
g947 and n1107_not n1110_not ; n1203
g948 and n1202_not n1203_not ; n1204
g949 and n1145 n1204_not ; n1205
g950 and n1142_not n1205 ; n1206
g951 and n1200_not n1206_not ; n1207
g952 and b[4]_not n1207_not ; n1208
g953 and n1089_not quotient[54]_not ; n1209
g954 and n1101_not n1105 ; n1210
g955 and n1100_not n1210 ; n1211
g956 and n1102_not n1105_not ; n1212
g957 and n1211_not n1212_not ; n1213
g958 and n1145 n1213_not ; n1214
g959 and n1142_not n1214 ; n1215
g960 and n1209_not n1215_not ; n1216
g961 and b[3]_not n1216_not ; n1217
g962 and n1094_not quotient[54]_not ; n1218
g963 and n1097_not n1099 ; n1219
g964 and n1095_not n1219 ; n1220
g965 and n1145 n1220_not ; n1221
g966 and n1100_not n1221 ; n1222
g967 and n1142_not n1222 ; n1223
g968 and n1218_not n1223_not ; n1224
g969 and b[2]_not n1224_not ; n1225
g970 and b[0] b[10]_not ; n1226
g971 and n390 n1226 ; n1227
g972 and n388 n1227 ; n1228
g973 and n378 n1228 ; n1229
g974 and n424 n1229 ; n1230
g975 and n1142_not n1230 ; n1231
g976 and a[54] n1231_not ; n1232
g977 and n263 n1099 ; n1233
g978 and n274 n1233 ; n1234
g979 and n344 n1234 ; n1235
g980 and n432 n1235 ; n1236
g981 and n1142_not n1236 ; n1237
g982 and n1232_not n1237_not ; n1238
g983 and b[1] n1238_not ; n1239
g984 and b[1]_not n1237_not ; n1240
g985 and n1232_not n1240 ; n1241
g986 and n1239_not n1241_not ; n1242
g987 and a[53]_not b[0] ; n1243
g988 and n1242_not n1243_not ; n1244
g989 and b[1]_not n1238_not ; n1245
g990 and n1244_not n1245_not ; n1246
g991 and b[2] n1223_not ; n1247
g992 and n1218_not n1247 ; n1248
g993 and n1225_not n1248_not ; n1249
g994 and n1246_not n1249 ; n1250
g995 and n1225_not n1250_not ; n1251
g996 and b[3] n1215_not ; n1252
g997 and n1209_not n1252 ; n1253
g998 and n1217_not n1253_not ; n1254
g999 and n1251_not n1254 ; n1255
g1000 and n1217_not n1255_not ; n1256
g1001 and b[4] n1206_not ; n1257
g1002 and n1200_not n1257 ; n1258
g1003 and n1208_not n1258_not ; n1259
g1004 and n1256_not n1259 ; n1260
g1005 and n1208_not n1260_not ; n1261
g1006 and b[5] n1197_not ; n1262
g1007 and n1191_not n1262 ; n1263
g1008 and n1199_not n1263_not ; n1264
g1009 and n1261_not n1264 ; n1265
g1010 and n1199_not n1265_not ; n1266
g1011 and b[6] n1188_not ; n1267
g1012 and n1182_not n1267 ; n1268
g1013 and n1190_not n1268_not ; n1269
g1014 and n1266_not n1269 ; n1270
g1015 and n1190_not n1270_not ; n1271
g1016 and b[7] n1179_not ; n1272
g1017 and n1173_not n1272 ; n1273
g1018 and n1181_not n1273_not ; n1274
g1019 and n1271_not n1274 ; n1275
g1020 and n1181_not n1275_not ; n1276
g1021 and b[8] n1170_not ; n1277
g1022 and n1164_not n1277 ; n1278
g1023 and n1172_not n1278_not ; n1279
g1024 and n1276_not n1279 ; n1280
g1025 and n1172_not n1280_not ; n1281
g1026 and b[9] n1153_not ; n1282
g1027 and n1147_not n1282 ; n1283
g1028 and n1163_not n1283_not ; n1284
g1029 and n1281_not n1284 ; n1285
g1030 and n1163_not n1285_not ; n1286
g1031 and b[10] n1155_not ; n1287
g1032 and n1160_not n1287 ; n1288
g1033 and n1162_not n1288_not ; n1289
g1034 and n1286_not n1289 ; n1290
g1035 and n1162_not n1290_not ; n1291
g1036 and n388 n390 ; n1292
g1037 and n378 n1292 ; n1293
g1038 and n424 n1293 ; n1294
g1039 and n1291_not n1294 ; quotient[53]
g1040 and n1154_not quotient[53]_not ; n1296
g1041 and n1172_not n1284 ; n1297
g1042 and n1280_not n1297 ; n1298
g1043 and n1281_not n1284_not ; n1299
g1044 and n1298_not n1299_not ; n1300
g1045 and n1294 n1300_not ; n1301
g1046 and n1291_not n1301 ; n1302
g1047 and n1296_not n1302_not ; n1303
g1048 and b[10]_not n1303_not ; n1304
g1049 and n1171_not quotient[53]_not ; n1305
g1050 and n1181_not n1279 ; n1306
g1051 and n1275_not n1306 ; n1307
g1052 and n1276_not n1279_not ; n1308
g1053 and n1307_not n1308_not ; n1309
g1054 and n1294 n1309_not ; n1310
g1055 and n1291_not n1310 ; n1311
g1056 and n1305_not n1311_not ; n1312
g1057 and b[9]_not n1312_not ; n1313
g1058 and n1180_not quotient[53]_not ; n1314
g1059 and n1190_not n1274 ; n1315
g1060 and n1270_not n1315 ; n1316
g1061 and n1271_not n1274_not ; n1317
g1062 and n1316_not n1317_not ; n1318
g1063 and n1294 n1318_not ; n1319
g1064 and n1291_not n1319 ; n1320
g1065 and n1314_not n1320_not ; n1321
g1066 and b[8]_not n1321_not ; n1322
g1067 and n1189_not quotient[53]_not ; n1323
g1068 and n1199_not n1269 ; n1324
g1069 and n1265_not n1324 ; n1325
g1070 and n1266_not n1269_not ; n1326
g1071 and n1325_not n1326_not ; n1327
g1072 and n1294 n1327_not ; n1328
g1073 and n1291_not n1328 ; n1329
g1074 and n1323_not n1329_not ; n1330
g1075 and b[7]_not n1330_not ; n1331
g1076 and n1198_not quotient[53]_not ; n1332
g1077 and n1208_not n1264 ; n1333
g1078 and n1260_not n1333 ; n1334
g1079 and n1261_not n1264_not ; n1335
g1080 and n1334_not n1335_not ; n1336
g1081 and n1294 n1336_not ; n1337
g1082 and n1291_not n1337 ; n1338
g1083 and n1332_not n1338_not ; n1339
g1084 and b[6]_not n1339_not ; n1340
g1085 and n1207_not quotient[53]_not ; n1341
g1086 and n1217_not n1259 ; n1342
g1087 and n1255_not n1342 ; n1343
g1088 and n1256_not n1259_not ; n1344
g1089 and n1343_not n1344_not ; n1345
g1090 and n1294 n1345_not ; n1346
g1091 and n1291_not n1346 ; n1347
g1092 and n1341_not n1347_not ; n1348
g1093 and b[5]_not n1348_not ; n1349
g1094 and n1216_not quotient[53]_not ; n1350
g1095 and n1225_not n1254 ; n1351
g1096 and n1250_not n1351 ; n1352
g1097 and n1251_not n1254_not ; n1353
g1098 and n1352_not n1353_not ; n1354
g1099 and n1294 n1354_not ; n1355
g1100 and n1291_not n1355 ; n1356
g1101 and n1350_not n1356_not ; n1357
g1102 and b[4]_not n1357_not ; n1358
g1103 and n1224_not quotient[53]_not ; n1359
g1104 and n1245_not n1249 ; n1360
g1105 and n1244_not n1360 ; n1361
g1106 and n1246_not n1249_not ; n1362
g1107 and n1361_not n1362_not ; n1363
g1108 and n1294 n1363_not ; n1364
g1109 and n1291_not n1364 ; n1365
g1110 and n1359_not n1365_not ; n1366
g1111 and b[3]_not n1366_not ; n1367
g1112 and n1238_not quotient[53]_not ; n1368
g1113 and n1241_not n1243 ; n1369
g1114 and n1239_not n1369 ; n1370
g1115 and n1294 n1370_not ; n1371
g1116 and n1244_not n1371 ; n1372
g1117 and n1291_not n1372 ; n1373
g1118 and n1368_not n1373_not ; n1374
g1119 and b[2]_not n1374_not ; n1375
g1120 and b[0] b[11]_not ; n1376
g1121 and n274 n1376 ; n1377
g1122 and n344 n1377 ; n1378
g1123 and n432 n1378 ; n1379
g1124 and n1291_not n1379 ; n1380
g1125 and a[53] n1380_not ; n1381
g1126 and n390 n1243 ; n1382
g1127 and n388 n1382 ; n1383
g1128 and n378 n1383 ; n1384
g1129 and n424 n1384 ; n1385
g1130 and n1291_not n1385 ; n1386
g1131 and n1381_not n1386_not ; n1387
g1132 and b[1] n1387_not ; n1388
g1133 and b[1]_not n1386_not ; n1389
g1134 and n1381_not n1389 ; n1390
g1135 and n1388_not n1390_not ; n1391
g1136 and a[52]_not b[0] ; n1392
g1137 and n1391_not n1392_not ; n1393
g1138 and b[1]_not n1387_not ; n1394
g1139 and n1393_not n1394_not ; n1395
g1140 and b[2] n1373_not ; n1396
g1141 and n1368_not n1396 ; n1397
g1142 and n1375_not n1397_not ; n1398
g1143 and n1395_not n1398 ; n1399
g1144 and n1375_not n1399_not ; n1400
g1145 and b[3] n1365_not ; n1401
g1146 and n1359_not n1401 ; n1402
g1147 and n1367_not n1402_not ; n1403
g1148 and n1400_not n1403 ; n1404
g1149 and n1367_not n1404_not ; n1405
g1150 and b[4] n1356_not ; n1406
g1151 and n1350_not n1406 ; n1407
g1152 and n1358_not n1407_not ; n1408
g1153 and n1405_not n1408 ; n1409
g1154 and n1358_not n1409_not ; n1410
g1155 and b[5] n1347_not ; n1411
g1156 and n1341_not n1411 ; n1412
g1157 and n1349_not n1412_not ; n1413
g1158 and n1410_not n1413 ; n1414
g1159 and n1349_not n1414_not ; n1415
g1160 and b[6] n1338_not ; n1416
g1161 and n1332_not n1416 ; n1417
g1162 and n1340_not n1417_not ; n1418
g1163 and n1415_not n1418 ; n1419
g1164 and n1340_not n1419_not ; n1420
g1165 and b[7] n1329_not ; n1421
g1166 and n1323_not n1421 ; n1422
g1167 and n1331_not n1422_not ; n1423
g1168 and n1420_not n1423 ; n1424
g1169 and n1331_not n1424_not ; n1425
g1170 and b[8] n1320_not ; n1426
g1171 and n1314_not n1426 ; n1427
g1172 and n1322_not n1427_not ; n1428
g1173 and n1425_not n1428 ; n1429
g1174 and n1322_not n1429_not ; n1430
g1175 and b[9] n1311_not ; n1431
g1176 and n1305_not n1431 ; n1432
g1177 and n1313_not n1432_not ; n1433
g1178 and n1430_not n1433 ; n1434
g1179 and n1313_not n1434_not ; n1435
g1180 and b[10] n1302_not ; n1436
g1181 and n1296_not n1436 ; n1437
g1182 and n1304_not n1437_not ; n1438
g1183 and n1435_not n1438 ; n1439
g1184 and n1304_not n1439_not ; n1440
g1185 and n1161_not quotient[53]_not ; n1441
g1186 and n1163_not n1289 ; n1442
g1187 and n1285_not n1442 ; n1443
g1188 and n1286_not n1289_not ; n1444
g1189 and n1443_not n1444_not ; n1445
g1190 and quotient[53] n1445_not ; n1446
g1191 and n1441_not n1446_not ; n1447
g1192 and b[11]_not n1447_not ; n1448
g1193 and b[11] n1441_not ; n1449
g1194 and n1446_not n1449 ; n1450
g1195 and n275 n318 ; n1451
g1196 and n512 n1451 ; n1452
g1197 and n1450_not n1452 ; n1453
g1198 and n1448_not n1453 ; n1454
g1199 and n1440_not n1454 ; n1455
g1200 and n1294 n1447_not ; n1456
g1201 and n1455_not n1456_not ; quotient[52]
g1202 and n1313_not n1438 ; n1458
g1203 and n1434_not n1458 ; n1459
g1204 and n1435_not n1438_not ; n1460
g1205 and n1459_not n1460_not ; n1461
g1206 and quotient[52] n1461_not ; n1462
g1207 and n1303_not n1456_not ; n1463
g1208 and n1455_not n1463 ; n1464
g1209 and n1462_not n1464_not ; n1465
g1210 and n1304_not n1450_not ; n1466
g1211 and n1448_not n1466 ; n1467
g1212 and n1439_not n1467 ; n1468
g1213 and n1448_not n1450_not ; n1469
g1214 and n1440_not n1469_not ; n1470
g1215 and n1468_not n1470_not ; n1471
g1216 and quotient[52] n1471_not ; n1472
g1217 and n1447_not n1456_not ; n1473
g1218 and n1455_not n1473 ; n1474
g1219 and n1472_not n1474_not ; n1475
g1220 and b[12]_not n1475_not ; n1476
g1221 and b[11]_not n1465_not ; n1477
g1222 and n1322_not n1433 ; n1478
g1223 and n1429_not n1478 ; n1479
g1224 and n1430_not n1433_not ; n1480
g1225 and n1479_not n1480_not ; n1481
g1226 and quotient[52] n1481_not ; n1482
g1227 and n1312_not n1456_not ; n1483
g1228 and n1455_not n1483 ; n1484
g1229 and n1482_not n1484_not ; n1485
g1230 and b[10]_not n1485_not ; n1486
g1231 and n1331_not n1428 ; n1487
g1232 and n1424_not n1487 ; n1488
g1233 and n1425_not n1428_not ; n1489
g1234 and n1488_not n1489_not ; n1490
g1235 and quotient[52] n1490_not ; n1491
g1236 and n1321_not n1456_not ; n1492
g1237 and n1455_not n1492 ; n1493
g1238 and n1491_not n1493_not ; n1494
g1239 and b[9]_not n1494_not ; n1495
g1240 and n1340_not n1423 ; n1496
g1241 and n1419_not n1496 ; n1497
g1242 and n1420_not n1423_not ; n1498
g1243 and n1497_not n1498_not ; n1499
g1244 and quotient[52] n1499_not ; n1500
g1245 and n1330_not n1456_not ; n1501
g1246 and n1455_not n1501 ; n1502
g1247 and n1500_not n1502_not ; n1503
g1248 and b[8]_not n1503_not ; n1504
g1249 and n1349_not n1418 ; n1505
g1250 and n1414_not n1505 ; n1506
g1251 and n1415_not n1418_not ; n1507
g1252 and n1506_not n1507_not ; n1508
g1253 and quotient[52] n1508_not ; n1509
g1254 and n1339_not n1456_not ; n1510
g1255 and n1455_not n1510 ; n1511
g1256 and n1509_not n1511_not ; n1512
g1257 and b[7]_not n1512_not ; n1513
g1258 and n1358_not n1413 ; n1514
g1259 and n1409_not n1514 ; n1515
g1260 and n1410_not n1413_not ; n1516
g1261 and n1515_not n1516_not ; n1517
g1262 and quotient[52] n1517_not ; n1518
g1263 and n1348_not n1456_not ; n1519
g1264 and n1455_not n1519 ; n1520
g1265 and n1518_not n1520_not ; n1521
g1266 and b[6]_not n1521_not ; n1522
g1267 and n1367_not n1408 ; n1523
g1268 and n1404_not n1523 ; n1524
g1269 and n1405_not n1408_not ; n1525
g1270 and n1524_not n1525_not ; n1526
g1271 and quotient[52] n1526_not ; n1527
g1272 and n1357_not n1456_not ; n1528
g1273 and n1455_not n1528 ; n1529
g1274 and n1527_not n1529_not ; n1530
g1275 and b[5]_not n1530_not ; n1531
g1276 and n1375_not n1403 ; n1532
g1277 and n1399_not n1532 ; n1533
g1278 and n1400_not n1403_not ; n1534
g1279 and n1533_not n1534_not ; n1535
g1280 and quotient[52] n1535_not ; n1536
g1281 and n1366_not n1456_not ; n1537
g1282 and n1455_not n1537 ; n1538
g1283 and n1536_not n1538_not ; n1539
g1284 and b[4]_not n1539_not ; n1540
g1285 and n1394_not n1398 ; n1541
g1286 and n1393_not n1541 ; n1542
g1287 and n1395_not n1398_not ; n1543
g1288 and n1542_not n1543_not ; n1544
g1289 and quotient[52] n1544_not ; n1545
g1290 and n1374_not n1456_not ; n1546
g1291 and n1455_not n1546 ; n1547
g1292 and n1545_not n1547_not ; n1548
g1293 and b[3]_not n1548_not ; n1549
g1294 and n1390_not n1392 ; n1550
g1295 and n1388_not n1550 ; n1551
g1296 and n1393_not n1551_not ; n1552
g1297 and quotient[52] n1552 ; n1553
g1298 and n1387_not n1456_not ; n1554
g1299 and n1455_not n1554 ; n1555
g1300 and n1553_not n1555_not ; n1556
g1301 and b[2]_not n1556_not ; n1557
g1302 and b[0] quotient[52] ; n1558
g1303 and a[52] n1558_not ; n1559
g1304 and n1392 quotient[52] ; n1560
g1305 and n1559_not n1560_not ; n1561
g1306 and b[1] n1561_not ; n1562
g1307 and b[1]_not n1560_not ; n1563
g1308 and n1559_not n1563 ; n1564
g1309 and n1562_not n1564_not ; n1565
g1310 and a[51]_not b[0] ; n1566
g1311 and n1565_not n1566_not ; n1567
g1312 and b[1]_not n1561_not ; n1568
g1313 and n1567_not n1568_not ; n1569
g1314 and b[2] n1555_not ; n1570
g1315 and n1553_not n1570 ; n1571
g1316 and n1557_not n1571_not ; n1572
g1317 and n1569_not n1572 ; n1573
g1318 and n1557_not n1573_not ; n1574
g1319 and b[3] n1547_not ; n1575
g1320 and n1545_not n1575 ; n1576
g1321 and n1549_not n1576_not ; n1577
g1322 and n1574_not n1577 ; n1578
g1323 and n1549_not n1578_not ; n1579
g1324 and b[4] n1538_not ; n1580
g1325 and n1536_not n1580 ; n1581
g1326 and n1540_not n1581_not ; n1582
g1327 and n1579_not n1582 ; n1583
g1328 and n1540_not n1583_not ; n1584
g1329 and b[5] n1529_not ; n1585
g1330 and n1527_not n1585 ; n1586
g1331 and n1531_not n1586_not ; n1587
g1332 and n1584_not n1587 ; n1588
g1333 and n1531_not n1588_not ; n1589
g1334 and b[6] n1520_not ; n1590
g1335 and n1518_not n1590 ; n1591
g1336 and n1522_not n1591_not ; n1592
g1337 and n1589_not n1592 ; n1593
g1338 and n1522_not n1593_not ; n1594
g1339 and b[7] n1511_not ; n1595
g1340 and n1509_not n1595 ; n1596
g1341 and n1513_not n1596_not ; n1597
g1342 and n1594_not n1597 ; n1598
g1343 and n1513_not n1598_not ; n1599
g1344 and b[8] n1502_not ; n1600
g1345 and n1500_not n1600 ; n1601
g1346 and n1504_not n1601_not ; n1602
g1347 and n1599_not n1602 ; n1603
g1348 and n1504_not n1603_not ; n1604
g1349 and b[9] n1493_not ; n1605
g1350 and n1491_not n1605 ; n1606
g1351 and n1495_not n1606_not ; n1607
g1352 and n1604_not n1607 ; n1608
g1353 and n1495_not n1608_not ; n1609
g1354 and b[10] n1484_not ; n1610
g1355 and n1482_not n1610 ; n1611
g1356 and n1486_not n1611_not ; n1612
g1357 and n1609_not n1612 ; n1613
g1358 and n1486_not n1613_not ; n1614
g1359 and b[11] n1464_not ; n1615
g1360 and n1462_not n1615 ; n1616
g1361 and n1477_not n1616_not ; n1617
g1362 and n1614_not n1617 ; n1618
g1363 and n1477_not n1618_not ; n1619
g1364 and b[12] n1474_not ; n1620
g1365 and n1472_not n1620 ; n1621
g1366 and n1476_not n1621_not ; n1622
g1367 and n1619_not n1622 ; n1623
g1368 and n1476_not n1623_not ; n1624
g1369 and n589 n591 ; n1625
g1370 and n599 n1625 ; n1626
g1371 and n1624_not n1626 ; quotient[51]
g1372 and n1465_not quotient[51]_not ; n1628
g1373 and n1486_not n1617 ; n1629
g1374 and n1613_not n1629 ; n1630
g1375 and n1614_not n1617_not ; n1631
g1376 and n1630_not n1631_not ; n1632
g1377 and n1626 n1632_not ; n1633
g1378 and n1624_not n1633 ; n1634
g1379 and n1628_not n1634_not ; n1635
g1380 and n1475_not quotient[51]_not ; n1636
g1381 and n1477_not n1622 ; n1637
g1382 and n1618_not n1637 ; n1638
g1383 and n1619_not n1622_not ; n1639
g1384 and n1638_not n1639_not ; n1640
g1385 and quotient[51] n1640_not ; n1641
g1386 and n1636_not n1641_not ; n1642
g1387 and b[13]_not n1642_not ; n1643
g1388 and b[12]_not n1635_not ; n1644
g1389 and n1485_not quotient[51]_not ; n1645
g1390 and n1495_not n1612 ; n1646
g1391 and n1608_not n1646 ; n1647
g1392 and n1609_not n1612_not ; n1648
g1393 and n1647_not n1648_not ; n1649
g1394 and n1626 n1649_not ; n1650
g1395 and n1624_not n1650 ; n1651
g1396 and n1645_not n1651_not ; n1652
g1397 and b[11]_not n1652_not ; n1653
g1398 and n1494_not quotient[51]_not ; n1654
g1399 and n1504_not n1607 ; n1655
g1400 and n1603_not n1655 ; n1656
g1401 and n1604_not n1607_not ; n1657
g1402 and n1656_not n1657_not ; n1658
g1403 and n1626 n1658_not ; n1659
g1404 and n1624_not n1659 ; n1660
g1405 and n1654_not n1660_not ; n1661
g1406 and b[10]_not n1661_not ; n1662
g1407 and n1503_not quotient[51]_not ; n1663
g1408 and n1513_not n1602 ; n1664
g1409 and n1598_not n1664 ; n1665
g1410 and n1599_not n1602_not ; n1666
g1411 and n1665_not n1666_not ; n1667
g1412 and n1626 n1667_not ; n1668
g1413 and n1624_not n1668 ; n1669
g1414 and n1663_not n1669_not ; n1670
g1415 and b[9]_not n1670_not ; n1671
g1416 and n1512_not quotient[51]_not ; n1672
g1417 and n1522_not n1597 ; n1673
g1418 and n1593_not n1673 ; n1674
g1419 and n1594_not n1597_not ; n1675
g1420 and n1674_not n1675_not ; n1676
g1421 and n1626 n1676_not ; n1677
g1422 and n1624_not n1677 ; n1678
g1423 and n1672_not n1678_not ; n1679
g1424 and b[8]_not n1679_not ; n1680
g1425 and n1521_not quotient[51]_not ; n1681
g1426 and n1531_not n1592 ; n1682
g1427 and n1588_not n1682 ; n1683
g1428 and n1589_not n1592_not ; n1684
g1429 and n1683_not n1684_not ; n1685
g1430 and n1626 n1685_not ; n1686
g1431 and n1624_not n1686 ; n1687
g1432 and n1681_not n1687_not ; n1688
g1433 and b[7]_not n1688_not ; n1689
g1434 and n1530_not quotient[51]_not ; n1690
g1435 and n1540_not n1587 ; n1691
g1436 and n1583_not n1691 ; n1692
g1437 and n1584_not n1587_not ; n1693
g1438 and n1692_not n1693_not ; n1694
g1439 and n1626 n1694_not ; n1695
g1440 and n1624_not n1695 ; n1696
g1441 and n1690_not n1696_not ; n1697
g1442 and b[6]_not n1697_not ; n1698
g1443 and n1539_not quotient[51]_not ; n1699
g1444 and n1549_not n1582 ; n1700
g1445 and n1578_not n1700 ; n1701
g1446 and n1579_not n1582_not ; n1702
g1447 and n1701_not n1702_not ; n1703
g1448 and n1626 n1703_not ; n1704
g1449 and n1624_not n1704 ; n1705
g1450 and n1699_not n1705_not ; n1706
g1451 and b[5]_not n1706_not ; n1707
g1452 and n1548_not quotient[51]_not ; n1708
g1453 and n1557_not n1577 ; n1709
g1454 and n1573_not n1709 ; n1710
g1455 and n1574_not n1577_not ; n1711
g1456 and n1710_not n1711_not ; n1712
g1457 and n1626 n1712_not ; n1713
g1458 and n1624_not n1713 ; n1714
g1459 and n1708_not n1714_not ; n1715
g1460 and b[4]_not n1715_not ; n1716
g1461 and n1556_not quotient[51]_not ; n1717
g1462 and n1568_not n1572 ; n1718
g1463 and n1567_not n1718 ; n1719
g1464 and n1569_not n1572_not ; n1720
g1465 and n1719_not n1720_not ; n1721
g1466 and n1626 n1721_not ; n1722
g1467 and n1624_not n1722 ; n1723
g1468 and n1717_not n1723_not ; n1724
g1469 and b[3]_not n1724_not ; n1725
g1470 and n1561_not quotient[51]_not ; n1726
g1471 and n1564_not n1566 ; n1727
g1472 and n1562_not n1727 ; n1728
g1473 and n1626 n1728_not ; n1729
g1474 and n1567_not n1729 ; n1730
g1475 and n1624_not n1730 ; n1731
g1476 and n1726_not n1731_not ; n1732
g1477 and b[2]_not n1732_not ; n1733
g1478 and b[0] b[13]_not ; n1734
g1479 and n273 n1734 ; n1735
g1480 and n271 n1735 ; n1736
g1481 and n318 n1736 ; n1737
g1482 and n512 n1737 ; n1738
g1483 and n1624_not n1738 ; n1739
g1484 and a[51] n1739_not ; n1740
g1485 and n388 n1566 ; n1741
g1486 and n378 n1741 ; n1742
g1487 and n424 n1742 ; n1743
g1488 and n1624_not n1743 ; n1744
g1489 and n1740_not n1744_not ; n1745
g1490 and b[1] n1745_not ; n1746
g1491 and b[1]_not n1744_not ; n1747
g1492 and n1740_not n1747 ; n1748
g1493 and n1746_not n1748_not ; n1749
g1494 and a[50]_not b[0] ; n1750
g1495 and n1749_not n1750_not ; n1751
g1496 and b[1]_not n1745_not ; n1752
g1497 and n1751_not n1752_not ; n1753
g1498 and b[2] n1731_not ; n1754
g1499 and n1726_not n1754 ; n1755
g1500 and n1733_not n1755_not ; n1756
g1501 and n1753_not n1756 ; n1757
g1502 and n1733_not n1757_not ; n1758
g1503 and b[3] n1723_not ; n1759
g1504 and n1717_not n1759 ; n1760
g1505 and n1725_not n1760_not ; n1761
g1506 and n1758_not n1761 ; n1762
g1507 and n1725_not n1762_not ; n1763
g1508 and b[4] n1714_not ; n1764
g1509 and n1708_not n1764 ; n1765
g1510 and n1716_not n1765_not ; n1766
g1511 and n1763_not n1766 ; n1767
g1512 and n1716_not n1767_not ; n1768
g1513 and b[5] n1705_not ; n1769
g1514 and n1699_not n1769 ; n1770
g1515 and n1707_not n1770_not ; n1771
g1516 and n1768_not n1771 ; n1772
g1517 and n1707_not n1772_not ; n1773
g1518 and b[6] n1696_not ; n1774
g1519 and n1690_not n1774 ; n1775
g1520 and n1698_not n1775_not ; n1776
g1521 and n1773_not n1776 ; n1777
g1522 and n1698_not n1777_not ; n1778
g1523 and b[7] n1687_not ; n1779
g1524 and n1681_not n1779 ; n1780
g1525 and n1689_not n1780_not ; n1781
g1526 and n1778_not n1781 ; n1782
g1527 and n1689_not n1782_not ; n1783
g1528 and b[8] n1678_not ; n1784
g1529 and n1672_not n1784 ; n1785
g1530 and n1680_not n1785_not ; n1786
g1531 and n1783_not n1786 ; n1787
g1532 and n1680_not n1787_not ; n1788
g1533 and b[9] n1669_not ; n1789
g1534 and n1663_not n1789 ; n1790
g1535 and n1671_not n1790_not ; n1791
g1536 and n1788_not n1791 ; n1792
g1537 and n1671_not n1792_not ; n1793
g1538 and b[10] n1660_not ; n1794
g1539 and n1654_not n1794 ; n1795
g1540 and n1662_not n1795_not ; n1796
g1541 and n1793_not n1796 ; n1797
g1542 and n1662_not n1797_not ; n1798
g1543 and b[11] n1651_not ; n1799
g1544 and n1645_not n1799 ; n1800
g1545 and n1653_not n1800_not ; n1801
g1546 and n1798_not n1801 ; n1802
g1547 and n1653_not n1802_not ; n1803
g1548 and b[12] n1634_not ; n1804
g1549 and n1628_not n1804 ; n1805
g1550 and n1644_not n1805_not ; n1806
g1551 and n1803_not n1806 ; n1807
g1552 and n1644_not n1807_not ; n1808
g1553 and b[13] n1636_not ; n1809
g1554 and n1641_not n1809 ; n1810
g1555 and n1643_not n1810_not ; n1811
g1556 and n1808_not n1811 ; n1812
g1557 and n1643_not n1812_not ; n1813
g1558 and n271 n273 ; n1814
g1559 and n318 n1814 ; n1815
g1560 and n512 n1815 ; n1816
g1561 and n1813_not n1816 ; quotient[50]
g1562 and n1635_not quotient[50]_not ; n1818
g1563 and n1653_not n1806 ; n1819
g1564 and n1802_not n1819 ; n1820
g1565 and n1803_not n1806_not ; n1821
g1566 and n1820_not n1821_not ; n1822
g1567 and n1816 n1822_not ; n1823
g1568 and n1813_not n1823 ; n1824
g1569 and n1818_not n1824_not ; n1825
g1570 and b[13]_not n1825_not ; n1826
g1571 and n1652_not quotient[50]_not ; n1827
g1572 and n1662_not n1801 ; n1828
g1573 and n1797_not n1828 ; n1829
g1574 and n1798_not n1801_not ; n1830
g1575 and n1829_not n1830_not ; n1831
g1576 and n1816 n1831_not ; n1832
g1577 and n1813_not n1832 ; n1833
g1578 and n1827_not n1833_not ; n1834
g1579 and b[12]_not n1834_not ; n1835
g1580 and n1661_not quotient[50]_not ; n1836
g1581 and n1671_not n1796 ; n1837
g1582 and n1792_not n1837 ; n1838
g1583 and n1793_not n1796_not ; n1839
g1584 and n1838_not n1839_not ; n1840
g1585 and n1816 n1840_not ; n1841
g1586 and n1813_not n1841 ; n1842
g1587 and n1836_not n1842_not ; n1843
g1588 and b[11]_not n1843_not ; n1844
g1589 and n1670_not quotient[50]_not ; n1845
g1590 and n1680_not n1791 ; n1846
g1591 and n1787_not n1846 ; n1847
g1592 and n1788_not n1791_not ; n1848
g1593 and n1847_not n1848_not ; n1849
g1594 and n1816 n1849_not ; n1850
g1595 and n1813_not n1850 ; n1851
g1596 and n1845_not n1851_not ; n1852
g1597 and b[10]_not n1852_not ; n1853
g1598 and n1679_not quotient[50]_not ; n1854
g1599 and n1689_not n1786 ; n1855
g1600 and n1782_not n1855 ; n1856
g1601 and n1783_not n1786_not ; n1857
g1602 and n1856_not n1857_not ; n1858
g1603 and n1816 n1858_not ; n1859
g1604 and n1813_not n1859 ; n1860
g1605 and n1854_not n1860_not ; n1861
g1606 and b[9]_not n1861_not ; n1862
g1607 and n1688_not quotient[50]_not ; n1863
g1608 and n1698_not n1781 ; n1864
g1609 and n1777_not n1864 ; n1865
g1610 and n1778_not n1781_not ; n1866
g1611 and n1865_not n1866_not ; n1867
g1612 and n1816 n1867_not ; n1868
g1613 and n1813_not n1868 ; n1869
g1614 and n1863_not n1869_not ; n1870
g1615 and b[8]_not n1870_not ; n1871
g1616 and n1697_not quotient[50]_not ; n1872
g1617 and n1707_not n1776 ; n1873
g1618 and n1772_not n1873 ; n1874
g1619 and n1773_not n1776_not ; n1875
g1620 and n1874_not n1875_not ; n1876
g1621 and n1816 n1876_not ; n1877
g1622 and n1813_not n1877 ; n1878
g1623 and n1872_not n1878_not ; n1879
g1624 and b[7]_not n1879_not ; n1880
g1625 and n1706_not quotient[50]_not ; n1881
g1626 and n1716_not n1771 ; n1882
g1627 and n1767_not n1882 ; n1883
g1628 and n1768_not n1771_not ; n1884
g1629 and n1883_not n1884_not ; n1885
g1630 and n1816 n1885_not ; n1886
g1631 and n1813_not n1886 ; n1887
g1632 and n1881_not n1887_not ; n1888
g1633 and b[6]_not n1888_not ; n1889
g1634 and n1715_not quotient[50]_not ; n1890
g1635 and n1725_not n1766 ; n1891
g1636 and n1762_not n1891 ; n1892
g1637 and n1763_not n1766_not ; n1893
g1638 and n1892_not n1893_not ; n1894
g1639 and n1816 n1894_not ; n1895
g1640 and n1813_not n1895 ; n1896
g1641 and n1890_not n1896_not ; n1897
g1642 and b[5]_not n1897_not ; n1898
g1643 and n1724_not quotient[50]_not ; n1899
g1644 and n1733_not n1761 ; n1900
g1645 and n1757_not n1900 ; n1901
g1646 and n1758_not n1761_not ; n1902
g1647 and n1901_not n1902_not ; n1903
g1648 and n1816 n1903_not ; n1904
g1649 and n1813_not n1904 ; n1905
g1650 and n1899_not n1905_not ; n1906
g1651 and b[4]_not n1906_not ; n1907
g1652 and n1732_not quotient[50]_not ; n1908
g1653 and n1752_not n1756 ; n1909
g1654 and n1751_not n1909 ; n1910
g1655 and n1753_not n1756_not ; n1911
g1656 and n1910_not n1911_not ; n1912
g1657 and n1816 n1912_not ; n1913
g1658 and n1813_not n1913 ; n1914
g1659 and n1908_not n1914_not ; n1915
g1660 and b[3]_not n1915_not ; n1916
g1661 and n1745_not quotient[50]_not ; n1917
g1662 and n1748_not n1750 ; n1918
g1663 and n1746_not n1918 ; n1919
g1664 and n1816 n1919_not ; n1920
g1665 and n1751_not n1920 ; n1921
g1666 and n1813_not n1921 ; n1922
g1667 and n1917_not n1922_not ; n1923
g1668 and b[2]_not n1923_not ; n1924
g1669 and b[0] b[14]_not ; n1925
g1670 and n387 n1925 ; n1926
g1671 and n369 n1926 ; n1927
g1672 and n589 n1927 ; n1928
g1673 and n599 n1928 ; n1929
g1674 and n1813_not n1929 ; n1930
g1675 and a[50] n1930_not ; n1931
g1676 and n273 n1750 ; n1932
g1677 and n271 n1932 ; n1933
g1678 and n318 n1933 ; n1934
g1679 and n512 n1934 ; n1935
g1680 and n1813_not n1935 ; n1936
g1681 and n1931_not n1936_not ; n1937
g1682 and b[1] n1937_not ; n1938
g1683 and b[1]_not n1936_not ; n1939
g1684 and n1931_not n1939 ; n1940
g1685 and n1938_not n1940_not ; n1941
g1686 and a[49]_not b[0] ; n1942
g1687 and n1941_not n1942_not ; n1943
g1688 and b[1]_not n1937_not ; n1944
g1689 and n1943_not n1944_not ; n1945
g1690 and b[2] n1922_not ; n1946
g1691 and n1917_not n1946 ; n1947
g1692 and n1924_not n1947_not ; n1948
g1693 and n1945_not n1948 ; n1949
g1694 and n1924_not n1949_not ; n1950
g1695 and b[3] n1914_not ; n1951
g1696 and n1908_not n1951 ; n1952
g1697 and n1916_not n1952_not ; n1953
g1698 and n1950_not n1953 ; n1954
g1699 and n1916_not n1954_not ; n1955
g1700 and b[4] n1905_not ; n1956
g1701 and n1899_not n1956 ; n1957
g1702 and n1907_not n1957_not ; n1958
g1703 and n1955_not n1958 ; n1959
g1704 and n1907_not n1959_not ; n1960
g1705 and b[5] n1896_not ; n1961
g1706 and n1890_not n1961 ; n1962
g1707 and n1898_not n1962_not ; n1963
g1708 and n1960_not n1963 ; n1964
g1709 and n1898_not n1964_not ; n1965
g1710 and b[6] n1887_not ; n1966
g1711 and n1881_not n1966 ; n1967
g1712 and n1889_not n1967_not ; n1968
g1713 and n1965_not n1968 ; n1969
g1714 and n1889_not n1969_not ; n1970
g1715 and b[7] n1878_not ; n1971
g1716 and n1872_not n1971 ; n1972
g1717 and n1880_not n1972_not ; n1973
g1718 and n1970_not n1973 ; n1974
g1719 and n1880_not n1974_not ; n1975
g1720 and b[8] n1869_not ; n1976
g1721 and n1863_not n1976 ; n1977
g1722 and n1871_not n1977_not ; n1978
g1723 and n1975_not n1978 ; n1979
g1724 and n1871_not n1979_not ; n1980
g1725 and b[9] n1860_not ; n1981
g1726 and n1854_not n1981 ; n1982
g1727 and n1862_not n1982_not ; n1983
g1728 and n1980_not n1983 ; n1984
g1729 and n1862_not n1984_not ; n1985
g1730 and b[10] n1851_not ; n1986
g1731 and n1845_not n1986 ; n1987
g1732 and n1853_not n1987_not ; n1988
g1733 and n1985_not n1988 ; n1989
g1734 and n1853_not n1989_not ; n1990
g1735 and b[11] n1842_not ; n1991
g1736 and n1836_not n1991 ; n1992
g1737 and n1844_not n1992_not ; n1993
g1738 and n1990_not n1993 ; n1994
g1739 and n1844_not n1994_not ; n1995
g1740 and b[12] n1833_not ; n1996
g1741 and n1827_not n1996 ; n1997
g1742 and n1835_not n1997_not ; n1998
g1743 and n1995_not n1998 ; n1999
g1744 and n1835_not n1999_not ; n2000
g1745 and b[13] n1824_not ; n2001
g1746 and n1818_not n2001 ; n2002
g1747 and n1826_not n2002_not ; n2003
g1748 and n2000_not n2003 ; n2004
g1749 and n1826_not n2004_not ; n2005
g1750 and n1642_not quotient[50]_not ; n2006
g1751 and n1644_not n1811 ; n2007
g1752 and n1807_not n2007 ; n2008
g1753 and n1808_not n1811_not ; n2009
g1754 and n2008_not n2009_not ; n2010
g1755 and quotient[50] n2010_not ; n2011
g1756 and n2006_not n2011_not ; n2012
g1757 and b[14]_not n2012_not ; n2013
g1758 and b[14] n2006_not ; n2014
g1759 and n2011_not n2014 ; n2015
g1760 and n369 n387 ; n2016
g1761 and n589 n2016 ; n2017
g1762 and n599 n2017 ; n2018
g1763 and n2015_not n2018 ; n2019
g1764 and n2013_not n2019 ; n2020
g1765 and n2005_not n2020 ; n2021
g1766 and n1816 n2012_not ; n2022
g1767 and n2021_not n2022_not ; quotient[49]
g1768 and n1835_not n2003 ; n2024
g1769 and n1999_not n2024 ; n2025
g1770 and n2000_not n2003_not ; n2026
g1771 and n2025_not n2026_not ; n2027
g1772 and quotient[49] n2027_not ; n2028
g1773 and n1825_not n2022_not ; n2029
g1774 and n2021_not n2029 ; n2030
g1775 and n2028_not n2030_not ; n2031
g1776 and n1826_not n2015_not ; n2032
g1777 and n2013_not n2032 ; n2033
g1778 and n2004_not n2033 ; n2034
g1779 and n2013_not n2015_not ; n2035
g1780 and n2005_not n2035_not ; n2036
g1781 and n2034_not n2036_not ; n2037
g1782 and quotient[49] n2037_not ; n2038
g1783 and n2012_not n2022_not ; n2039
g1784 and n2021_not n2039 ; n2040
g1785 and n2038_not n2040_not ; n2041
g1786 and b[15]_not n2041_not ; n2042
g1787 and b[14]_not n2031_not ; n2043
g1788 and n1844_not n1998 ; n2044
g1789 and n1994_not n2044 ; n2045
g1790 and n1995_not n1998_not ; n2046
g1791 and n2045_not n2046_not ; n2047
g1792 and quotient[49] n2047_not ; n2048
g1793 and n1834_not n2022_not ; n2049
g1794 and n2021_not n2049 ; n2050
g1795 and n2048_not n2050_not ; n2051
g1796 and b[13]_not n2051_not ; n2052
g1797 and n1853_not n1993 ; n2053
g1798 and n1989_not n2053 ; n2054
g1799 and n1990_not n1993_not ; n2055
g1800 and n2054_not n2055_not ; n2056
g1801 and quotient[49] n2056_not ; n2057
g1802 and n1843_not n2022_not ; n2058
g1803 and n2021_not n2058 ; n2059
g1804 and n2057_not n2059_not ; n2060
g1805 and b[12]_not n2060_not ; n2061
g1806 and n1862_not n1988 ; n2062
g1807 and n1984_not n2062 ; n2063
g1808 and n1985_not n1988_not ; n2064
g1809 and n2063_not n2064_not ; n2065
g1810 and quotient[49] n2065_not ; n2066
g1811 and n1852_not n2022_not ; n2067
g1812 and n2021_not n2067 ; n2068
g1813 and n2066_not n2068_not ; n2069
g1814 and b[11]_not n2069_not ; n2070
g1815 and n1871_not n1983 ; n2071
g1816 and n1979_not n2071 ; n2072
g1817 and n1980_not n1983_not ; n2073
g1818 and n2072_not n2073_not ; n2074
g1819 and quotient[49] n2074_not ; n2075
g1820 and n1861_not n2022_not ; n2076
g1821 and n2021_not n2076 ; n2077
g1822 and n2075_not n2077_not ; n2078
g1823 and b[10]_not n2078_not ; n2079
g1824 and n1880_not n1978 ; n2080
g1825 and n1974_not n2080 ; n2081
g1826 and n1975_not n1978_not ; n2082
g1827 and n2081_not n2082_not ; n2083
g1828 and quotient[49] n2083_not ; n2084
g1829 and n1870_not n2022_not ; n2085
g1830 and n2021_not n2085 ; n2086
g1831 and n2084_not n2086_not ; n2087
g1832 and b[9]_not n2087_not ; n2088
g1833 and n1889_not n1973 ; n2089
g1834 and n1969_not n2089 ; n2090
g1835 and n1970_not n1973_not ; n2091
g1836 and n2090_not n2091_not ; n2092
g1837 and quotient[49] n2092_not ; n2093
g1838 and n1879_not n2022_not ; n2094
g1839 and n2021_not n2094 ; n2095
g1840 and n2093_not n2095_not ; n2096
g1841 and b[8]_not n2096_not ; n2097
g1842 and n1898_not n1968 ; n2098
g1843 and n1964_not n2098 ; n2099
g1844 and n1965_not n1968_not ; n2100
g1845 and n2099_not n2100_not ; n2101
g1846 and quotient[49] n2101_not ; n2102
g1847 and n1888_not n2022_not ; n2103
g1848 and n2021_not n2103 ; n2104
g1849 and n2102_not n2104_not ; n2105
g1850 and b[7]_not n2105_not ; n2106
g1851 and n1907_not n1963 ; n2107
g1852 and n1959_not n2107 ; n2108
g1853 and n1960_not n1963_not ; n2109
g1854 and n2108_not n2109_not ; n2110
g1855 and quotient[49] n2110_not ; n2111
g1856 and n1897_not n2022_not ; n2112
g1857 and n2021_not n2112 ; n2113
g1858 and n2111_not n2113_not ; n2114
g1859 and b[6]_not n2114_not ; n2115
g1860 and n1916_not n1958 ; n2116
g1861 and n1954_not n2116 ; n2117
g1862 and n1955_not n1958_not ; n2118
g1863 and n2117_not n2118_not ; n2119
g1864 and quotient[49] n2119_not ; n2120
g1865 and n1906_not n2022_not ; n2121
g1866 and n2021_not n2121 ; n2122
g1867 and n2120_not n2122_not ; n2123
g1868 and b[5]_not n2123_not ; n2124
g1869 and n1924_not n1953 ; n2125
g1870 and n1949_not n2125 ; n2126
g1871 and n1950_not n1953_not ; n2127
g1872 and n2126_not n2127_not ; n2128
g1873 and quotient[49] n2128_not ; n2129
g1874 and n1915_not n2022_not ; n2130
g1875 and n2021_not n2130 ; n2131
g1876 and n2129_not n2131_not ; n2132
g1877 and b[4]_not n2132_not ; n2133
g1878 and n1944_not n1948 ; n2134
g1879 and n1943_not n2134 ; n2135
g1880 and n1945_not n1948_not ; n2136
g1881 and n2135_not n2136_not ; n2137
g1882 and quotient[49] n2137_not ; n2138
g1883 and n1923_not n2022_not ; n2139
g1884 and n2021_not n2139 ; n2140
g1885 and n2138_not n2140_not ; n2141
g1886 and b[3]_not n2141_not ; n2142
g1887 and n1940_not n1942 ; n2143
g1888 and n1938_not n2143 ; n2144
g1889 and n1943_not n2144_not ; n2145
g1890 and quotient[49] n2145 ; n2146
g1891 and n1937_not n2022_not ; n2147
g1892 and n2021_not n2147 ; n2148
g1893 and n2146_not n2148_not ; n2149
g1894 and b[2]_not n2149_not ; n2150
g1895 and b[0] quotient[49] ; n2151
g1896 and a[49] n2151_not ; n2152
g1897 and n1942 quotient[49] ; n2153
g1898 and n2152_not n2153_not ; n2154
g1899 and b[1] n2154_not ; n2155
g1900 and b[1]_not n2153_not ; n2156
g1901 and n2152_not n2156 ; n2157
g1902 and n2155_not n2157_not ; n2158
g1903 and a[48]_not b[0] ; n2159
g1904 and n2158_not n2159_not ; n2160
g1905 and b[1]_not n2154_not ; n2161
g1906 and n2160_not n2161_not ; n2162
g1907 and b[2] n2148_not ; n2163
g1908 and n2146_not n2163 ; n2164
g1909 and n2150_not n2164_not ; n2165
g1910 and n2162_not n2165 ; n2166
g1911 and n2150_not n2166_not ; n2167
g1912 and b[3] n2140_not ; n2168
g1913 and n2138_not n2168 ; n2169
g1914 and n2142_not n2169_not ; n2170
g1915 and n2167_not n2170 ; n2171
g1916 and n2142_not n2171_not ; n2172
g1917 and b[4] n2131_not ; n2173
g1918 and n2129_not n2173 ; n2174
g1919 and n2133_not n2174_not ; n2175
g1920 and n2172_not n2175 ; n2176
g1921 and n2133_not n2176_not ; n2177
g1922 and b[5] n2122_not ; n2178
g1923 and n2120_not n2178 ; n2179
g1924 and n2124_not n2179_not ; n2180
g1925 and n2177_not n2180 ; n2181
g1926 and n2124_not n2181_not ; n2182
g1927 and b[6] n2113_not ; n2183
g1928 and n2111_not n2183 ; n2184
g1929 and n2115_not n2184_not ; n2185
g1930 and n2182_not n2185 ; n2186
g1931 and n2115_not n2186_not ; n2187
g1932 and b[7] n2104_not ; n2188
g1933 and n2102_not n2188 ; n2189
g1934 and n2106_not n2189_not ; n2190
g1935 and n2187_not n2190 ; n2191
g1936 and n2106_not n2191_not ; n2192
g1937 and b[8] n2095_not ; n2193
g1938 and n2093_not n2193 ; n2194
g1939 and n2097_not n2194_not ; n2195
g1940 and n2192_not n2195 ; n2196
g1941 and n2097_not n2196_not ; n2197
g1942 and b[9] n2086_not ; n2198
g1943 and n2084_not n2198 ; n2199
g1944 and n2088_not n2199_not ; n2200
g1945 and n2197_not n2200 ; n2201
g1946 and n2088_not n2201_not ; n2202
g1947 and b[10] n2077_not ; n2203
g1948 and n2075_not n2203 ; n2204
g1949 and n2079_not n2204_not ; n2205
g1950 and n2202_not n2205 ; n2206
g1951 and n2079_not n2206_not ; n2207
g1952 and b[11] n2068_not ; n2208
g1953 and n2066_not n2208 ; n2209
g1954 and n2070_not n2209_not ; n2210
g1955 and n2207_not n2210 ; n2211
g1956 and n2070_not n2211_not ; n2212
g1957 and b[12] n2059_not ; n2213
g1958 and n2057_not n2213 ; n2214
g1959 and n2061_not n2214_not ; n2215
g1960 and n2212_not n2215 ; n2216
g1961 and n2061_not n2216_not ; n2217
g1962 and b[13] n2050_not ; n2218
g1963 and n2048_not n2218 ; n2219
g1964 and n2052_not n2219_not ; n2220
g1965 and n2217_not n2220 ; n2221
g1966 and n2052_not n2221_not ; n2222
g1967 and b[14] n2030_not ; n2223
g1968 and n2028_not n2223 ; n2224
g1969 and n2043_not n2224_not ; n2225
g1970 and n2222_not n2225 ; n2226
g1971 and n2043_not n2226_not ; n2227
g1972 and b[15] n2040_not ; n2228
g1973 and n2038_not n2228 ; n2229
g1974 and n2042_not n2229_not ; n2230
g1975 and n2227_not n2230 ; n2231
g1976 and n2042_not n2231_not ; n2232
g1977 and n346 n2232_not ; quotient[48]
g1978 and n2031_not quotient[48]_not ; n2234
g1979 and n2052_not n2225 ; n2235
g1980 and n2221_not n2235 ; n2236
g1981 and n2222_not n2225_not ; n2237
g1982 and n2236_not n2237_not ; n2238
g1983 and n346 n2238_not ; n2239
g1984 and n2232_not n2239 ; n2240
g1985 and n2234_not n2240_not ; n2241
g1986 and n2041_not quotient[48]_not ; n2242
g1987 and n2043_not n2230 ; n2243
g1988 and n2226_not n2243 ; n2244
g1989 and n2227_not n2230_not ; n2245
g1990 and n2244_not n2245_not ; n2246
g1991 and quotient[48] n2246_not ; n2247
g1992 and n2242_not n2247_not ; n2248
g1993 and b[16]_not n2248_not ; n2249
g1994 and b[15]_not n2241_not ; n2250
g1995 and n2051_not quotient[48]_not ; n2251
g1996 and n2061_not n2220 ; n2252
g1997 and n2216_not n2252 ; n2253
g1998 and n2217_not n2220_not ; n2254
g1999 and n2253_not n2254_not ; n2255
g2000 and n346 n2255_not ; n2256
g2001 and n2232_not n2256 ; n2257
g2002 and n2251_not n2257_not ; n2258
g2003 and b[14]_not n2258_not ; n2259
g2004 and n2060_not quotient[48]_not ; n2260
g2005 and n2070_not n2215 ; n2261
g2006 and n2211_not n2261 ; n2262
g2007 and n2212_not n2215_not ; n2263
g2008 and n2262_not n2263_not ; n2264
g2009 and n346 n2264_not ; n2265
g2010 and n2232_not n2265 ; n2266
g2011 and n2260_not n2266_not ; n2267
g2012 and b[13]_not n2267_not ; n2268
g2013 and n2069_not quotient[48]_not ; n2269
g2014 and n2079_not n2210 ; n2270
g2015 and n2206_not n2270 ; n2271
g2016 and n2207_not n2210_not ; n2272
g2017 and n2271_not n2272_not ; n2273
g2018 and n346 n2273_not ; n2274
g2019 and n2232_not n2274 ; n2275
g2020 and n2269_not n2275_not ; n2276
g2021 and b[12]_not n2276_not ; n2277
g2022 and n2078_not quotient[48]_not ; n2278
g2023 and n2088_not n2205 ; n2279
g2024 and n2201_not n2279 ; n2280
g2025 and n2202_not n2205_not ; n2281
g2026 and n2280_not n2281_not ; n2282
g2027 and n346 n2282_not ; n2283
g2028 and n2232_not n2283 ; n2284
g2029 and n2278_not n2284_not ; n2285
g2030 and b[11]_not n2285_not ; n2286
g2031 and n2087_not quotient[48]_not ; n2287
g2032 and n2097_not n2200 ; n2288
g2033 and n2196_not n2288 ; n2289
g2034 and n2197_not n2200_not ; n2290
g2035 and n2289_not n2290_not ; n2291
g2036 and n346 n2291_not ; n2292
g2037 and n2232_not n2292 ; n2293
g2038 and n2287_not n2293_not ; n2294
g2039 and b[10]_not n2294_not ; n2295
g2040 and n2096_not quotient[48]_not ; n2296
g2041 and n2106_not n2195 ; n2297
g2042 and n2191_not n2297 ; n2298
g2043 and n2192_not n2195_not ; n2299
g2044 and n2298_not n2299_not ; n2300
g2045 and n346 n2300_not ; n2301
g2046 and n2232_not n2301 ; n2302
g2047 and n2296_not n2302_not ; n2303
g2048 and b[9]_not n2303_not ; n2304
g2049 and n2105_not quotient[48]_not ; n2305
g2050 and n2115_not n2190 ; n2306
g2051 and n2186_not n2306 ; n2307
g2052 and n2187_not n2190_not ; n2308
g2053 and n2307_not n2308_not ; n2309
g2054 and n346 n2309_not ; n2310
g2055 and n2232_not n2310 ; n2311
g2056 and n2305_not n2311_not ; n2312
g2057 and b[8]_not n2312_not ; n2313
g2058 and n2114_not quotient[48]_not ; n2314
g2059 and n2124_not n2185 ; n2315
g2060 and n2181_not n2315 ; n2316
g2061 and n2182_not n2185_not ; n2317
g2062 and n2316_not n2317_not ; n2318
g2063 and n346 n2318_not ; n2319
g2064 and n2232_not n2319 ; n2320
g2065 and n2314_not n2320_not ; n2321
g2066 and b[7]_not n2321_not ; n2322
g2067 and n2123_not quotient[48]_not ; n2323
g2068 and n2133_not n2180 ; n2324
g2069 and n2176_not n2324 ; n2325
g2070 and n2177_not n2180_not ; n2326
g2071 and n2325_not n2326_not ; n2327
g2072 and n346 n2327_not ; n2328
g2073 and n2232_not n2328 ; n2329
g2074 and n2323_not n2329_not ; n2330
g2075 and b[6]_not n2330_not ; n2331
g2076 and n2132_not quotient[48]_not ; n2332
g2077 and n2142_not n2175 ; n2333
g2078 and n2171_not n2333 ; n2334
g2079 and n2172_not n2175_not ; n2335
g2080 and n2334_not n2335_not ; n2336
g2081 and n346 n2336_not ; n2337
g2082 and n2232_not n2337 ; n2338
g2083 and n2332_not n2338_not ; n2339
g2084 and b[5]_not n2339_not ; n2340
g2085 and n2141_not quotient[48]_not ; n2341
g2086 and n2150_not n2170 ; n2342
g2087 and n2166_not n2342 ; n2343
g2088 and n2167_not n2170_not ; n2344
g2089 and n2343_not n2344_not ; n2345
g2090 and n346 n2345_not ; n2346
g2091 and n2232_not n2346 ; n2347
g2092 and n2341_not n2347_not ; n2348
g2093 and b[4]_not n2348_not ; n2349
g2094 and n2149_not quotient[48]_not ; n2350
g2095 and n2161_not n2165 ; n2351
g2096 and n2160_not n2351 ; n2352
g2097 and n2162_not n2165_not ; n2353
g2098 and n2352_not n2353_not ; n2354
g2099 and n346 n2354_not ; n2355
g2100 and n2232_not n2355 ; n2356
g2101 and n2350_not n2356_not ; n2357
g2102 and b[3]_not n2357_not ; n2358
g2103 and n2154_not quotient[48]_not ; n2359
g2104 and n2157_not n2159 ; n2360
g2105 and n2155_not n2360 ; n2361
g2106 and n346 n2361_not ; n2362
g2107 and n2160_not n2362 ; n2363
g2108 and n2232_not n2363 ; n2364
g2109 and n2359_not n2364_not ; n2365
g2110 and b[2]_not n2365_not ; n2366
g2111 and b[0] b[16]_not ; n2367
g2112 and n369 n2367 ; n2368
g2113 and n589 n2368 ; n2369
g2114 and n599 n2369 ; n2370
g2115 and n2232_not n2370 ; n2371
g2116 and a[48] n2371_not ; n2372
g2117 and n271 n2159 ; n2373
g2118 and n318 n2373 ; n2374
g2119 and n512 n2374 ; n2375
g2120 and n2232_not n2375 ; n2376
g2121 and n2372_not n2376_not ; n2377
g2122 and b[1] n2377_not ; n2378
g2123 and b[1]_not n2376_not ; n2379
g2124 and n2372_not n2379 ; n2380
g2125 and n2378_not n2380_not ; n2381
g2126 and a[47]_not b[0] ; n2382
g2127 and n2381_not n2382_not ; n2383
g2128 and b[1]_not n2377_not ; n2384
g2129 and n2383_not n2384_not ; n2385
g2130 and b[2] n2364_not ; n2386
g2131 and n2359_not n2386 ; n2387
g2132 and n2366_not n2387_not ; n2388
g2133 and n2385_not n2388 ; n2389
g2134 and n2366_not n2389_not ; n2390
g2135 and b[3] n2356_not ; n2391
g2136 and n2350_not n2391 ; n2392
g2137 and n2358_not n2392_not ; n2393
g2138 and n2390_not n2393 ; n2394
g2139 and n2358_not n2394_not ; n2395
g2140 and b[4] n2347_not ; n2396
g2141 and n2341_not n2396 ; n2397
g2142 and n2349_not n2397_not ; n2398
g2143 and n2395_not n2398 ; n2399
g2144 and n2349_not n2399_not ; n2400
g2145 and b[5] n2338_not ; n2401
g2146 and n2332_not n2401 ; n2402
g2147 and n2340_not n2402_not ; n2403
g2148 and n2400_not n2403 ; n2404
g2149 and n2340_not n2404_not ; n2405
g2150 and b[6] n2329_not ; n2406
g2151 and n2323_not n2406 ; n2407
g2152 and n2331_not n2407_not ; n2408
g2153 and n2405_not n2408 ; n2409
g2154 and n2331_not n2409_not ; n2410
g2155 and b[7] n2320_not ; n2411
g2156 and n2314_not n2411 ; n2412
g2157 and n2322_not n2412_not ; n2413
g2158 and n2410_not n2413 ; n2414
g2159 and n2322_not n2414_not ; n2415
g2160 and b[8] n2311_not ; n2416
g2161 and n2305_not n2416 ; n2417
g2162 and n2313_not n2417_not ; n2418
g2163 and n2415_not n2418 ; n2419
g2164 and n2313_not n2419_not ; n2420
g2165 and b[9] n2302_not ; n2421
g2166 and n2296_not n2421 ; n2422
g2167 and n2304_not n2422_not ; n2423
g2168 and n2420_not n2423 ; n2424
g2169 and n2304_not n2424_not ; n2425
g2170 and b[10] n2293_not ; n2426
g2171 and n2287_not n2426 ; n2427
g2172 and n2295_not n2427_not ; n2428
g2173 and n2425_not n2428 ; n2429
g2174 and n2295_not n2429_not ; n2430
g2175 and b[11] n2284_not ; n2431
g2176 and n2278_not n2431 ; n2432
g2177 and n2286_not n2432_not ; n2433
g2178 and n2430_not n2433 ; n2434
g2179 and n2286_not n2434_not ; n2435
g2180 and b[12] n2275_not ; n2436
g2181 and n2269_not n2436 ; n2437
g2182 and n2277_not n2437_not ; n2438
g2183 and n2435_not n2438 ; n2439
g2184 and n2277_not n2439_not ; n2440
g2185 and b[13] n2266_not ; n2441
g2186 and n2260_not n2441 ; n2442
g2187 and n2268_not n2442_not ; n2443
g2188 and n2440_not n2443 ; n2444
g2189 and n2268_not n2444_not ; n2445
g2190 and b[14] n2257_not ; n2446
g2191 and n2251_not n2446 ; n2447
g2192 and n2259_not n2447_not ; n2448
g2193 and n2445_not n2448 ; n2449
g2194 and n2259_not n2449_not ; n2450
g2195 and b[15] n2240_not ; n2451
g2196 and n2234_not n2451 ; n2452
g2197 and n2250_not n2452_not ; n2453
g2198 and n2450_not n2453 ; n2454
g2199 and n2250_not n2454_not ; n2455
g2200 and b[16] n2242_not ; n2456
g2201 and n2247_not n2456 ; n2457
g2202 and n2249_not n2457_not ; n2458
g2203 and n2455_not n2458 ; n2459
g2204 and n2249_not n2459_not ; n2460
g2205 and n475 n2460_not ; quotient[47]
g2206 and n2241_not quotient[47]_not ; n2462
g2207 and n2259_not n2453 ; n2463
g2208 and n2449_not n2463 ; n2464
g2209 and n2450_not n2453_not ; n2465
g2210 and n2464_not n2465_not ; n2466
g2211 and n475 n2466_not ; n2467
g2212 and n2460_not n2467 ; n2468
g2213 and n2462_not n2468_not ; n2469
g2214 and b[16]_not n2469_not ; n2470
g2215 and n2258_not quotient[47]_not ; n2471
g2216 and n2268_not n2448 ; n2472
g2217 and n2444_not n2472 ; n2473
g2218 and n2445_not n2448_not ; n2474
g2219 and n2473_not n2474_not ; n2475
g2220 and n475 n2475_not ; n2476
g2221 and n2460_not n2476 ; n2477
g2222 and n2471_not n2477_not ; n2478
g2223 and b[15]_not n2478_not ; n2479
g2224 and n2267_not quotient[47]_not ; n2480
g2225 and n2277_not n2443 ; n2481
g2226 and n2439_not n2481 ; n2482
g2227 and n2440_not n2443_not ; n2483
g2228 and n2482_not n2483_not ; n2484
g2229 and n475 n2484_not ; n2485
g2230 and n2460_not n2485 ; n2486
g2231 and n2480_not n2486_not ; n2487
g2232 and b[14]_not n2487_not ; n2488
g2233 and n2276_not quotient[47]_not ; n2489
g2234 and n2286_not n2438 ; n2490
g2235 and n2434_not n2490 ; n2491
g2236 and n2435_not n2438_not ; n2492
g2237 and n2491_not n2492_not ; n2493
g2238 and n475 n2493_not ; n2494
g2239 and n2460_not n2494 ; n2495
g2240 and n2489_not n2495_not ; n2496
g2241 and b[13]_not n2496_not ; n2497
g2242 and n2285_not quotient[47]_not ; n2498
g2243 and n2295_not n2433 ; n2499
g2244 and n2429_not n2499 ; n2500
g2245 and n2430_not n2433_not ; n2501
g2246 and n2500_not n2501_not ; n2502
g2247 and n475 n2502_not ; n2503
g2248 and n2460_not n2503 ; n2504
g2249 and n2498_not n2504_not ; n2505
g2250 and b[12]_not n2505_not ; n2506
g2251 and n2294_not quotient[47]_not ; n2507
g2252 and n2304_not n2428 ; n2508
g2253 and n2424_not n2508 ; n2509
g2254 and n2425_not n2428_not ; n2510
g2255 and n2509_not n2510_not ; n2511
g2256 and n475 n2511_not ; n2512
g2257 and n2460_not n2512 ; n2513
g2258 and n2507_not n2513_not ; n2514
g2259 and b[11]_not n2514_not ; n2515
g2260 and n2303_not quotient[47]_not ; n2516
g2261 and n2313_not n2423 ; n2517
g2262 and n2419_not n2517 ; n2518
g2263 and n2420_not n2423_not ; n2519
g2264 and n2518_not n2519_not ; n2520
g2265 and n475 n2520_not ; n2521
g2266 and n2460_not n2521 ; n2522
g2267 and n2516_not n2522_not ; n2523
g2268 and b[10]_not n2523_not ; n2524
g2269 and n2312_not quotient[47]_not ; n2525
g2270 and n2322_not n2418 ; n2526
g2271 and n2414_not n2526 ; n2527
g2272 and n2415_not n2418_not ; n2528
g2273 and n2527_not n2528_not ; n2529
g2274 and n475 n2529_not ; n2530
g2275 and n2460_not n2530 ; n2531
g2276 and n2525_not n2531_not ; n2532
g2277 and b[9]_not n2532_not ; n2533
g2278 and n2321_not quotient[47]_not ; n2534
g2279 and n2331_not n2413 ; n2535
g2280 and n2409_not n2535 ; n2536
g2281 and n2410_not n2413_not ; n2537
g2282 and n2536_not n2537_not ; n2538
g2283 and n475 n2538_not ; n2539
g2284 and n2460_not n2539 ; n2540
g2285 and n2534_not n2540_not ; n2541
g2286 and b[8]_not n2541_not ; n2542
g2287 and n2330_not quotient[47]_not ; n2543
g2288 and n2340_not n2408 ; n2544
g2289 and n2404_not n2544 ; n2545
g2290 and n2405_not n2408_not ; n2546
g2291 and n2545_not n2546_not ; n2547
g2292 and n475 n2547_not ; n2548
g2293 and n2460_not n2548 ; n2549
g2294 and n2543_not n2549_not ; n2550
g2295 and b[7]_not n2550_not ; n2551
g2296 and n2339_not quotient[47]_not ; n2552
g2297 and n2349_not n2403 ; n2553
g2298 and n2399_not n2553 ; n2554
g2299 and n2400_not n2403_not ; n2555
g2300 and n2554_not n2555_not ; n2556
g2301 and n475 n2556_not ; n2557
g2302 and n2460_not n2557 ; n2558
g2303 and n2552_not n2558_not ; n2559
g2304 and b[6]_not n2559_not ; n2560
g2305 and n2348_not quotient[47]_not ; n2561
g2306 and n2358_not n2398 ; n2562
g2307 and n2394_not n2562 ; n2563
g2308 and n2395_not n2398_not ; n2564
g2309 and n2563_not n2564_not ; n2565
g2310 and n475 n2565_not ; n2566
g2311 and n2460_not n2566 ; n2567
g2312 and n2561_not n2567_not ; n2568
g2313 and b[5]_not n2568_not ; n2569
g2314 and n2357_not quotient[47]_not ; n2570
g2315 and n2366_not n2393 ; n2571
g2316 and n2389_not n2571 ; n2572
g2317 and n2390_not n2393_not ; n2573
g2318 and n2572_not n2573_not ; n2574
g2319 and n475 n2574_not ; n2575
g2320 and n2460_not n2575 ; n2576
g2321 and n2570_not n2576_not ; n2577
g2322 and b[4]_not n2577_not ; n2578
g2323 and n2365_not quotient[47]_not ; n2579
g2324 and n2384_not n2388 ; n2580
g2325 and n2383_not n2580 ; n2581
g2326 and n2385_not n2388_not ; n2582
g2327 and n2581_not n2582_not ; n2583
g2328 and n475 n2583_not ; n2584
g2329 and n2460_not n2584 ; n2585
g2330 and n2579_not n2585_not ; n2586
g2331 and b[3]_not n2586_not ; n2587
g2332 and n2377_not quotient[47]_not ; n2588
g2333 and n2380_not n2382 ; n2589
g2334 and n2378_not n2589 ; n2590
g2335 and n475 n2590_not ; n2591
g2336 and n2383_not n2591 ; n2592
g2337 and n2460_not n2592 ; n2593
g2338 and n2588_not n2593_not ; n2594
g2339 and b[2]_not n2594_not ; n2595
g2340 and b[0] b[17]_not ; n2596
g2341 and n270 n2596 ; n2597
g2342 and n309 n2597 ; n2598
g2343 and n343 n2598 ; n2599
g2344 and n341 n2599 ; n2600
g2345 and n338 n2600 ; n2601
g2346 and n2460_not n2601 ; n2602
g2347 and a[47] n2602_not ; n2603
g2348 and n369 n2382 ; n2604
g2349 and n589 n2604 ; n2605
g2350 and n599 n2605 ; n2606
g2351 and n2460_not n2606 ; n2607
g2352 and n2603_not n2607_not ; n2608
g2353 and b[1] n2608_not ; n2609
g2354 and b[1]_not n2607_not ; n2610
g2355 and n2603_not n2610 ; n2611
g2356 and n2609_not n2611_not ; n2612
g2357 and a[46]_not b[0] ; n2613
g2358 and n2612_not n2613_not ; n2614
g2359 and b[1]_not n2608_not ; n2615
g2360 and n2614_not n2615_not ; n2616
g2361 and b[2] n2593_not ; n2617
g2362 and n2588_not n2617 ; n2618
g2363 and n2595_not n2618_not ; n2619
g2364 and n2616_not n2619 ; n2620
g2365 and n2595_not n2620_not ; n2621
g2366 and b[3] n2585_not ; n2622
g2367 and n2579_not n2622 ; n2623
g2368 and n2587_not n2623_not ; n2624
g2369 and n2621_not n2624 ; n2625
g2370 and n2587_not n2625_not ; n2626
g2371 and b[4] n2576_not ; n2627
g2372 and n2570_not n2627 ; n2628
g2373 and n2578_not n2628_not ; n2629
g2374 and n2626_not n2629 ; n2630
g2375 and n2578_not n2630_not ; n2631
g2376 and b[5] n2567_not ; n2632
g2377 and n2561_not n2632 ; n2633
g2378 and n2569_not n2633_not ; n2634
g2379 and n2631_not n2634 ; n2635
g2380 and n2569_not n2635_not ; n2636
g2381 and b[6] n2558_not ; n2637
g2382 and n2552_not n2637 ; n2638
g2383 and n2560_not n2638_not ; n2639
g2384 and n2636_not n2639 ; n2640
g2385 and n2560_not n2640_not ; n2641
g2386 and b[7] n2549_not ; n2642
g2387 and n2543_not n2642 ; n2643
g2388 and n2551_not n2643_not ; n2644
g2389 and n2641_not n2644 ; n2645
g2390 and n2551_not n2645_not ; n2646
g2391 and b[8] n2540_not ; n2647
g2392 and n2534_not n2647 ; n2648
g2393 and n2542_not n2648_not ; n2649
g2394 and n2646_not n2649 ; n2650
g2395 and n2542_not n2650_not ; n2651
g2396 and b[9] n2531_not ; n2652
g2397 and n2525_not n2652 ; n2653
g2398 and n2533_not n2653_not ; n2654
g2399 and n2651_not n2654 ; n2655
g2400 and n2533_not n2655_not ; n2656
g2401 and b[10] n2522_not ; n2657
g2402 and n2516_not n2657 ; n2658
g2403 and n2524_not n2658_not ; n2659
g2404 and n2656_not n2659 ; n2660
g2405 and n2524_not n2660_not ; n2661
g2406 and b[11] n2513_not ; n2662
g2407 and n2507_not n2662 ; n2663
g2408 and n2515_not n2663_not ; n2664
g2409 and n2661_not n2664 ; n2665
g2410 and n2515_not n2665_not ; n2666
g2411 and b[12] n2504_not ; n2667
g2412 and n2498_not n2667 ; n2668
g2413 and n2506_not n2668_not ; n2669
g2414 and n2666_not n2669 ; n2670
g2415 and n2506_not n2670_not ; n2671
g2416 and b[13] n2495_not ; n2672
g2417 and n2489_not n2672 ; n2673
g2418 and n2497_not n2673_not ; n2674
g2419 and n2671_not n2674 ; n2675
g2420 and n2497_not n2675_not ; n2676
g2421 and b[14] n2486_not ; n2677
g2422 and n2480_not n2677 ; n2678
g2423 and n2488_not n2678_not ; n2679
g2424 and n2676_not n2679 ; n2680
g2425 and n2488_not n2680_not ; n2681
g2426 and b[15] n2477_not ; n2682
g2427 and n2471_not n2682 ; n2683
g2428 and n2479_not n2683_not ; n2684
g2429 and n2681_not n2684 ; n2685
g2430 and n2479_not n2685_not ; n2686
g2431 and b[16] n2468_not ; n2687
g2432 and n2462_not n2687 ; n2688
g2433 and n2470_not n2688_not ; n2689
g2434 and n2686_not n2689 ; n2690
g2435 and n2470_not n2690_not ; n2691
g2436 and n2248_not quotient[47]_not ; n2692
g2437 and n2250_not n2458 ; n2693
g2438 and n2454_not n2693 ; n2694
g2439 and n2455_not n2458_not ; n2695
g2440 and n2694_not n2695_not ; n2696
g2441 and quotient[47] n2696_not ; n2697
g2442 and n2692_not n2697_not ; n2698
g2443 and b[17]_not n2698_not ; n2699
g2444 and b[17] n2692_not ; n2700
g2445 and n2697_not n2700 ; n2701
g2446 and n270 n309 ; n2702
g2447 and n343 n2702 ; n2703
g2448 and n341 n2703 ; n2704
g2449 and n338 n2704 ; n2705
g2450 and n2701_not n2705 ; n2706
g2451 and n2699_not n2706 ; n2707
g2452 and n2691_not n2707 ; n2708
g2453 and n475 n2698_not ; n2709
g2454 and n2708_not n2709_not ; quotient[46]
g2455 and n2479_not n2689 ; n2711
g2456 and n2685_not n2711 ; n2712
g2457 and n2686_not n2689_not ; n2713
g2458 and n2712_not n2713_not ; n2714
g2459 and quotient[46] n2714_not ; n2715
g2460 and n2469_not n2709_not ; n2716
g2461 and n2708_not n2716 ; n2717
g2462 and n2715_not n2717_not ; n2718
g2463 and n2470_not n2701_not ; n2719
g2464 and n2699_not n2719 ; n2720
g2465 and n2690_not n2720 ; n2721
g2466 and n2699_not n2701_not ; n2722
g2467 and n2691_not n2722_not ; n2723
g2468 and n2721_not n2723_not ; n2724
g2469 and quotient[46] n2724_not ; n2725
g2470 and n2698_not n2709_not ; n2726
g2471 and n2708_not n2726 ; n2727
g2472 and n2725_not n2727_not ; n2728
g2473 and b[18]_not n2728_not ; n2729
g2474 and b[17]_not n2718_not ; n2730
g2475 and n2488_not n2684 ; n2731
g2476 and n2680_not n2731 ; n2732
g2477 and n2681_not n2684_not ; n2733
g2478 and n2732_not n2733_not ; n2734
g2479 and quotient[46] n2734_not ; n2735
g2480 and n2478_not n2709_not ; n2736
g2481 and n2708_not n2736 ; n2737
g2482 and n2735_not n2737_not ; n2738
g2483 and b[16]_not n2738_not ; n2739
g2484 and n2497_not n2679 ; n2740
g2485 and n2675_not n2740 ; n2741
g2486 and n2676_not n2679_not ; n2742
g2487 and n2741_not n2742_not ; n2743
g2488 and quotient[46] n2743_not ; n2744
g2489 and n2487_not n2709_not ; n2745
g2490 and n2708_not n2745 ; n2746
g2491 and n2744_not n2746_not ; n2747
g2492 and b[15]_not n2747_not ; n2748
g2493 and n2506_not n2674 ; n2749
g2494 and n2670_not n2749 ; n2750
g2495 and n2671_not n2674_not ; n2751
g2496 and n2750_not n2751_not ; n2752
g2497 and quotient[46] n2752_not ; n2753
g2498 and n2496_not n2709_not ; n2754
g2499 and n2708_not n2754 ; n2755
g2500 and n2753_not n2755_not ; n2756
g2501 and b[14]_not n2756_not ; n2757
g2502 and n2515_not n2669 ; n2758
g2503 and n2665_not n2758 ; n2759
g2504 and n2666_not n2669_not ; n2760
g2505 and n2759_not n2760_not ; n2761
g2506 and quotient[46] n2761_not ; n2762
g2507 and n2505_not n2709_not ; n2763
g2508 and n2708_not n2763 ; n2764
g2509 and n2762_not n2764_not ; n2765
g2510 and b[13]_not n2765_not ; n2766
g2511 and n2524_not n2664 ; n2767
g2512 and n2660_not n2767 ; n2768
g2513 and n2661_not n2664_not ; n2769
g2514 and n2768_not n2769_not ; n2770
g2515 and quotient[46] n2770_not ; n2771
g2516 and n2514_not n2709_not ; n2772
g2517 and n2708_not n2772 ; n2773
g2518 and n2771_not n2773_not ; n2774
g2519 and b[12]_not n2774_not ; n2775
g2520 and n2533_not n2659 ; n2776
g2521 and n2655_not n2776 ; n2777
g2522 and n2656_not n2659_not ; n2778
g2523 and n2777_not n2778_not ; n2779
g2524 and quotient[46] n2779_not ; n2780
g2525 and n2523_not n2709_not ; n2781
g2526 and n2708_not n2781 ; n2782
g2527 and n2780_not n2782_not ; n2783
g2528 and b[11]_not n2783_not ; n2784
g2529 and n2542_not n2654 ; n2785
g2530 and n2650_not n2785 ; n2786
g2531 and n2651_not n2654_not ; n2787
g2532 and n2786_not n2787_not ; n2788
g2533 and quotient[46] n2788_not ; n2789
g2534 and n2532_not n2709_not ; n2790
g2535 and n2708_not n2790 ; n2791
g2536 and n2789_not n2791_not ; n2792
g2537 and b[10]_not n2792_not ; n2793
g2538 and n2551_not n2649 ; n2794
g2539 and n2645_not n2794 ; n2795
g2540 and n2646_not n2649_not ; n2796
g2541 and n2795_not n2796_not ; n2797
g2542 and quotient[46] n2797_not ; n2798
g2543 and n2541_not n2709_not ; n2799
g2544 and n2708_not n2799 ; n2800
g2545 and n2798_not n2800_not ; n2801
g2546 and b[9]_not n2801_not ; n2802
g2547 and n2560_not n2644 ; n2803
g2548 and n2640_not n2803 ; n2804
g2549 and n2641_not n2644_not ; n2805
g2550 and n2804_not n2805_not ; n2806
g2551 and quotient[46] n2806_not ; n2807
g2552 and n2550_not n2709_not ; n2808
g2553 and n2708_not n2808 ; n2809
g2554 and n2807_not n2809_not ; n2810
g2555 and b[8]_not n2810_not ; n2811
g2556 and n2569_not n2639 ; n2812
g2557 and n2635_not n2812 ; n2813
g2558 and n2636_not n2639_not ; n2814
g2559 and n2813_not n2814_not ; n2815
g2560 and quotient[46] n2815_not ; n2816
g2561 and n2559_not n2709_not ; n2817
g2562 and n2708_not n2817 ; n2818
g2563 and n2816_not n2818_not ; n2819
g2564 and b[7]_not n2819_not ; n2820
g2565 and n2578_not n2634 ; n2821
g2566 and n2630_not n2821 ; n2822
g2567 and n2631_not n2634_not ; n2823
g2568 and n2822_not n2823_not ; n2824
g2569 and quotient[46] n2824_not ; n2825
g2570 and n2568_not n2709_not ; n2826
g2571 and n2708_not n2826 ; n2827
g2572 and n2825_not n2827_not ; n2828
g2573 and b[6]_not n2828_not ; n2829
g2574 and n2587_not n2629 ; n2830
g2575 and n2625_not n2830 ; n2831
g2576 and n2626_not n2629_not ; n2832
g2577 and n2831_not n2832_not ; n2833
g2578 and quotient[46] n2833_not ; n2834
g2579 and n2577_not n2709_not ; n2835
g2580 and n2708_not n2835 ; n2836
g2581 and n2834_not n2836_not ; n2837
g2582 and b[5]_not n2837_not ; n2838
g2583 and n2595_not n2624 ; n2839
g2584 and n2620_not n2839 ; n2840
g2585 and n2621_not n2624_not ; n2841
g2586 and n2840_not n2841_not ; n2842
g2587 and quotient[46] n2842_not ; n2843
g2588 and n2586_not n2709_not ; n2844
g2589 and n2708_not n2844 ; n2845
g2590 and n2843_not n2845_not ; n2846
g2591 and b[4]_not n2846_not ; n2847
g2592 and n2615_not n2619 ; n2848
g2593 and n2614_not n2848 ; n2849
g2594 and n2616_not n2619_not ; n2850
g2595 and n2849_not n2850_not ; n2851
g2596 and quotient[46] n2851_not ; n2852
g2597 and n2594_not n2709_not ; n2853
g2598 and n2708_not n2853 ; n2854
g2599 and n2852_not n2854_not ; n2855
g2600 and b[3]_not n2855_not ; n2856
g2601 and n2611_not n2613 ; n2857
g2602 and n2609_not n2857 ; n2858
g2603 and n2614_not n2858_not ; n2859
g2604 and quotient[46] n2859 ; n2860
g2605 and n2608_not n2709_not ; n2861
g2606 and n2708_not n2861 ; n2862
g2607 and n2860_not n2862_not ; n2863
g2608 and b[2]_not n2863_not ; n2864
g2609 and b[0] quotient[46] ; n2865
g2610 and a[46] n2865_not ; n2866
g2611 and n2613 quotient[46] ; n2867
g2612 and n2866_not n2867_not ; n2868
g2613 and b[1] n2868_not ; n2869
g2614 and b[1]_not n2867_not ; n2870
g2615 and n2866_not n2870 ; n2871
g2616 and n2869_not n2871_not ; n2872
g2617 and a[45]_not b[0] ; n2873
g2618 and n2872_not n2873_not ; n2874
g2619 and b[1]_not n2868_not ; n2875
g2620 and n2874_not n2875_not ; n2876
g2621 and b[2] n2862_not ; n2877
g2622 and n2860_not n2877 ; n2878
g2623 and n2864_not n2878_not ; n2879
g2624 and n2876_not n2879 ; n2880
g2625 and n2864_not n2880_not ; n2881
g2626 and b[3] n2854_not ; n2882
g2627 and n2852_not n2882 ; n2883
g2628 and n2856_not n2883_not ; n2884
g2629 and n2881_not n2884 ; n2885
g2630 and n2856_not n2885_not ; n2886
g2631 and b[4] n2845_not ; n2887
g2632 and n2843_not n2887 ; n2888
g2633 and n2847_not n2888_not ; n2889
g2634 and n2886_not n2889 ; n2890
g2635 and n2847_not n2890_not ; n2891
g2636 and b[5] n2836_not ; n2892
g2637 and n2834_not n2892 ; n2893
g2638 and n2838_not n2893_not ; n2894
g2639 and n2891_not n2894 ; n2895
g2640 and n2838_not n2895_not ; n2896
g2641 and b[6] n2827_not ; n2897
g2642 and n2825_not n2897 ; n2898
g2643 and n2829_not n2898_not ; n2899
g2644 and n2896_not n2899 ; n2900
g2645 and n2829_not n2900_not ; n2901
g2646 and b[7] n2818_not ; n2902
g2647 and n2816_not n2902 ; n2903
g2648 and n2820_not n2903_not ; n2904
g2649 and n2901_not n2904 ; n2905
g2650 and n2820_not n2905_not ; n2906
g2651 and b[8] n2809_not ; n2907
g2652 and n2807_not n2907 ; n2908
g2653 and n2811_not n2908_not ; n2909
g2654 and n2906_not n2909 ; n2910
g2655 and n2811_not n2910_not ; n2911
g2656 and b[9] n2800_not ; n2912
g2657 and n2798_not n2912 ; n2913
g2658 and n2802_not n2913_not ; n2914
g2659 and n2911_not n2914 ; n2915
g2660 and n2802_not n2915_not ; n2916
g2661 and b[10] n2791_not ; n2917
g2662 and n2789_not n2917 ; n2918
g2663 and n2793_not n2918_not ; n2919
g2664 and n2916_not n2919 ; n2920
g2665 and n2793_not n2920_not ; n2921
g2666 and b[11] n2782_not ; n2922
g2667 and n2780_not n2922 ; n2923
g2668 and n2784_not n2923_not ; n2924
g2669 and n2921_not n2924 ; n2925
g2670 and n2784_not n2925_not ; n2926
g2671 and b[12] n2773_not ; n2927
g2672 and n2771_not n2927 ; n2928
g2673 and n2775_not n2928_not ; n2929
g2674 and n2926_not n2929 ; n2930
g2675 and n2775_not n2930_not ; n2931
g2676 and b[13] n2764_not ; n2932
g2677 and n2762_not n2932 ; n2933
g2678 and n2766_not n2933_not ; n2934
g2679 and n2931_not n2934 ; n2935
g2680 and n2766_not n2935_not ; n2936
g2681 and b[14] n2755_not ; n2937
g2682 and n2753_not n2937 ; n2938
g2683 and n2757_not n2938_not ; n2939
g2684 and n2936_not n2939 ; n2940
g2685 and n2757_not n2940_not ; n2941
g2686 and b[15] n2746_not ; n2942
g2687 and n2744_not n2942 ; n2943
g2688 and n2748_not n2943_not ; n2944
g2689 and n2941_not n2944 ; n2945
g2690 and n2748_not n2945_not ; n2946
g2691 and b[16] n2737_not ; n2947
g2692 and n2735_not n2947 ; n2948
g2693 and n2739_not n2948_not ; n2949
g2694 and n2946_not n2949 ; n2950
g2695 and n2739_not n2950_not ; n2951
g2696 and b[17] n2717_not ; n2952
g2697 and n2715_not n2952 ; n2953
g2698 and n2730_not n2953_not ; n2954
g2699 and n2951_not n2954 ; n2955
g2700 and n2730_not n2955_not ; n2956
g2701 and b[18] n2727_not ; n2957
g2702 and n2725_not n2957 ; n2958
g2703 and n2729_not n2958_not ; n2959
g2704 and n2956_not n2959 ; n2960
g2705 and n2729_not n2960_not ; n2961
g2706 and n366 n368 ; n2962
g2707 and n377 n2962 ; n2963
g2708 and n423 n2963 ; n2964
g2709 and n408 n2964 ; n2965
g2710 and n2961_not n2965 ; quotient[45]
g2711 and n2718_not quotient[45]_not ; n2967
g2712 and n2739_not n2954 ; n2968
g2713 and n2950_not n2968 ; n2969
g2714 and n2951_not n2954_not ; n2970
g2715 and n2969_not n2970_not ; n2971
g2716 and n2965 n2971_not ; n2972
g2717 and n2961_not n2972 ; n2973
g2718 and n2967_not n2973_not ; n2974
g2719 and n2728_not quotient[45]_not ; n2975
g2720 and n2730_not n2959 ; n2976
g2721 and n2955_not n2976 ; n2977
g2722 and n2956_not n2959_not ; n2978
g2723 and n2977_not n2978_not ; n2979
g2724 and quotient[45] n2979_not ; n2980
g2725 and n2975_not n2980_not ; n2981
g2726 and b[19]_not n2981_not ; n2982
g2727 and b[18]_not n2974_not ; n2983
g2728 and n2738_not quotient[45]_not ; n2984
g2729 and n2748_not n2949 ; n2985
g2730 and n2945_not n2985 ; n2986
g2731 and n2946_not n2949_not ; n2987
g2732 and n2986_not n2987_not ; n2988
g2733 and n2965 n2988_not ; n2989
g2734 and n2961_not n2989 ; n2990
g2735 and n2984_not n2990_not ; n2991
g2736 and b[17]_not n2991_not ; n2992
g2737 and n2747_not quotient[45]_not ; n2993
g2738 and n2757_not n2944 ; n2994
g2739 and n2940_not n2994 ; n2995
g2740 and n2941_not n2944_not ; n2996
g2741 and n2995_not n2996_not ; n2997
g2742 and n2965 n2997_not ; n2998
g2743 and n2961_not n2998 ; n2999
g2744 and n2993_not n2999_not ; n3000
g2745 and b[16]_not n3000_not ; n3001
g2746 and n2756_not quotient[45]_not ; n3002
g2747 and n2766_not n2939 ; n3003
g2748 and n2935_not n3003 ; n3004
g2749 and n2936_not n2939_not ; n3005
g2750 and n3004_not n3005_not ; n3006
g2751 and n2965 n3006_not ; n3007
g2752 and n2961_not n3007 ; n3008
g2753 and n3002_not n3008_not ; n3009
g2754 and b[15]_not n3009_not ; n3010
g2755 and n2765_not quotient[45]_not ; n3011
g2756 and n2775_not n2934 ; n3012
g2757 and n2930_not n3012 ; n3013
g2758 and n2931_not n2934_not ; n3014
g2759 and n3013_not n3014_not ; n3015
g2760 and n2965 n3015_not ; n3016
g2761 and n2961_not n3016 ; n3017
g2762 and n3011_not n3017_not ; n3018
g2763 and b[14]_not n3018_not ; n3019
g2764 and n2774_not quotient[45]_not ; n3020
g2765 and n2784_not n2929 ; n3021
g2766 and n2925_not n3021 ; n3022
g2767 and n2926_not n2929_not ; n3023
g2768 and n3022_not n3023_not ; n3024
g2769 and n2965 n3024_not ; n3025
g2770 and n2961_not n3025 ; n3026
g2771 and n3020_not n3026_not ; n3027
g2772 and b[13]_not n3027_not ; n3028
g2773 and n2783_not quotient[45]_not ; n3029
g2774 and n2793_not n2924 ; n3030
g2775 and n2920_not n3030 ; n3031
g2776 and n2921_not n2924_not ; n3032
g2777 and n3031_not n3032_not ; n3033
g2778 and n2965 n3033_not ; n3034
g2779 and n2961_not n3034 ; n3035
g2780 and n3029_not n3035_not ; n3036
g2781 and b[12]_not n3036_not ; n3037
g2782 and n2792_not quotient[45]_not ; n3038
g2783 and n2802_not n2919 ; n3039
g2784 and n2915_not n3039 ; n3040
g2785 and n2916_not n2919_not ; n3041
g2786 and n3040_not n3041_not ; n3042
g2787 and n2965 n3042_not ; n3043
g2788 and n2961_not n3043 ; n3044
g2789 and n3038_not n3044_not ; n3045
g2790 and b[11]_not n3045_not ; n3046
g2791 and n2801_not quotient[45]_not ; n3047
g2792 and n2811_not n2914 ; n3048
g2793 and n2910_not n3048 ; n3049
g2794 and n2911_not n2914_not ; n3050
g2795 and n3049_not n3050_not ; n3051
g2796 and n2965 n3051_not ; n3052
g2797 and n2961_not n3052 ; n3053
g2798 and n3047_not n3053_not ; n3054
g2799 and b[10]_not n3054_not ; n3055
g2800 and n2810_not quotient[45]_not ; n3056
g2801 and n2820_not n2909 ; n3057
g2802 and n2905_not n3057 ; n3058
g2803 and n2906_not n2909_not ; n3059
g2804 and n3058_not n3059_not ; n3060
g2805 and n2965 n3060_not ; n3061
g2806 and n2961_not n3061 ; n3062
g2807 and n3056_not n3062_not ; n3063
g2808 and b[9]_not n3063_not ; n3064
g2809 and n2819_not quotient[45]_not ; n3065
g2810 and n2829_not n2904 ; n3066
g2811 and n2900_not n3066 ; n3067
g2812 and n2901_not n2904_not ; n3068
g2813 and n3067_not n3068_not ; n3069
g2814 and n2965 n3069_not ; n3070
g2815 and n2961_not n3070 ; n3071
g2816 and n3065_not n3071_not ; n3072
g2817 and b[8]_not n3072_not ; n3073
g2818 and n2828_not quotient[45]_not ; n3074
g2819 and n2838_not n2899 ; n3075
g2820 and n2895_not n3075 ; n3076
g2821 and n2896_not n2899_not ; n3077
g2822 and n3076_not n3077_not ; n3078
g2823 and n2965 n3078_not ; n3079
g2824 and n2961_not n3079 ; n3080
g2825 and n3074_not n3080_not ; n3081
g2826 and b[7]_not n3081_not ; n3082
g2827 and n2837_not quotient[45]_not ; n3083
g2828 and n2847_not n2894 ; n3084
g2829 and n2890_not n3084 ; n3085
g2830 and n2891_not n2894_not ; n3086
g2831 and n3085_not n3086_not ; n3087
g2832 and n2965 n3087_not ; n3088
g2833 and n2961_not n3088 ; n3089
g2834 and n3083_not n3089_not ; n3090
g2835 and b[6]_not n3090_not ; n3091
g2836 and n2846_not quotient[45]_not ; n3092
g2837 and n2856_not n2889 ; n3093
g2838 and n2885_not n3093 ; n3094
g2839 and n2886_not n2889_not ; n3095
g2840 and n3094_not n3095_not ; n3096
g2841 and n2965 n3096_not ; n3097
g2842 and n2961_not n3097 ; n3098
g2843 and n3092_not n3098_not ; n3099
g2844 and b[5]_not n3099_not ; n3100
g2845 and n2855_not quotient[45]_not ; n3101
g2846 and n2864_not n2884 ; n3102
g2847 and n2880_not n3102 ; n3103
g2848 and n2881_not n2884_not ; n3104
g2849 and n3103_not n3104_not ; n3105
g2850 and n2965 n3105_not ; n3106
g2851 and n2961_not n3106 ; n3107
g2852 and n3101_not n3107_not ; n3108
g2853 and b[4]_not n3108_not ; n3109
g2854 and n2863_not quotient[45]_not ; n3110
g2855 and n2875_not n2879 ; n3111
g2856 and n2874_not n3111 ; n3112
g2857 and n2876_not n2879_not ; n3113
g2858 and n3112_not n3113_not ; n3114
g2859 and n2965 n3114_not ; n3115
g2860 and n2961_not n3115 ; n3116
g2861 and n3110_not n3116_not ; n3117
g2862 and b[3]_not n3117_not ; n3118
g2863 and n2868_not quotient[45]_not ; n3119
g2864 and n2871_not n2873 ; n3120
g2865 and n2869_not n3120 ; n3121
g2866 and n2965 n3121_not ; n3122
g2867 and n2874_not n3122 ; n3123
g2868 and n2961_not n3123 ; n3124
g2869 and n3119_not n3124_not ; n3125
g2870 and b[2]_not n3125_not ; n3126
g2871 and b[0] b[19]_not ; n3127
g2872 and n309 n3127 ; n3128
g2873 and n343 n3128 ; n3129
g2874 and n341 n3129 ; n3130
g2875 and n338 n3130 ; n3131
g2876 and n2961_not n3131 ; n3132
g2877 and a[45] n3132_not ; n3133
g2878 and n368 n2873 ; n3134
g2879 and n366 n3134 ; n3135
g2880 and n377 n3135 ; n3136
g2881 and n423 n3136 ; n3137
g2882 and n408 n3137 ; n3138
g2883 and n2961_not n3138 ; n3139
g2884 and n3133_not n3139_not ; n3140
g2885 and b[1] n3140_not ; n3141
g2886 and b[1]_not n3139_not ; n3142
g2887 and n3133_not n3142 ; n3143
g2888 and n3141_not n3143_not ; n3144
g2889 and a[44]_not b[0] ; n3145
g2890 and n3144_not n3145_not ; n3146
g2891 and b[1]_not n3140_not ; n3147
g2892 and n3146_not n3147_not ; n3148
g2893 and b[2] n3124_not ; n3149
g2894 and n3119_not n3149 ; n3150
g2895 and n3126_not n3150_not ; n3151
g2896 and n3148_not n3151 ; n3152
g2897 and n3126_not n3152_not ; n3153
g2898 and b[3] n3116_not ; n3154
g2899 and n3110_not n3154 ; n3155
g2900 and n3118_not n3155_not ; n3156
g2901 and n3153_not n3156 ; n3157
g2902 and n3118_not n3157_not ; n3158
g2903 and b[4] n3107_not ; n3159
g2904 and n3101_not n3159 ; n3160
g2905 and n3109_not n3160_not ; n3161
g2906 and n3158_not n3161 ; n3162
g2907 and n3109_not n3162_not ; n3163
g2908 and b[5] n3098_not ; n3164
g2909 and n3092_not n3164 ; n3165
g2910 and n3100_not n3165_not ; n3166
g2911 and n3163_not n3166 ; n3167
g2912 and n3100_not n3167_not ; n3168
g2913 and b[6] n3089_not ; n3169
g2914 and n3083_not n3169 ; n3170
g2915 and n3091_not n3170_not ; n3171
g2916 and n3168_not n3171 ; n3172
g2917 and n3091_not n3172_not ; n3173
g2918 and b[7] n3080_not ; n3174
g2919 and n3074_not n3174 ; n3175
g2920 and n3082_not n3175_not ; n3176
g2921 and n3173_not n3176 ; n3177
g2922 and n3082_not n3177_not ; n3178
g2923 and b[8] n3071_not ; n3179
g2924 and n3065_not n3179 ; n3180
g2925 and n3073_not n3180_not ; n3181
g2926 and n3178_not n3181 ; n3182
g2927 and n3073_not n3182_not ; n3183
g2928 and b[9] n3062_not ; n3184
g2929 and n3056_not n3184 ; n3185
g2930 and n3064_not n3185_not ; n3186
g2931 and n3183_not n3186 ; n3187
g2932 and n3064_not n3187_not ; n3188
g2933 and b[10] n3053_not ; n3189
g2934 and n3047_not n3189 ; n3190
g2935 and n3055_not n3190_not ; n3191
g2936 and n3188_not n3191 ; n3192
g2937 and n3055_not n3192_not ; n3193
g2938 and b[11] n3044_not ; n3194
g2939 and n3038_not n3194 ; n3195
g2940 and n3046_not n3195_not ; n3196
g2941 and n3193_not n3196 ; n3197
g2942 and n3046_not n3197_not ; n3198
g2943 and b[12] n3035_not ; n3199
g2944 and n3029_not n3199 ; n3200
g2945 and n3037_not n3200_not ; n3201
g2946 and n3198_not n3201 ; n3202
g2947 and n3037_not n3202_not ; n3203
g2948 and b[13] n3026_not ; n3204
g2949 and n3020_not n3204 ; n3205
g2950 and n3028_not n3205_not ; n3206
g2951 and n3203_not n3206 ; n3207
g2952 and n3028_not n3207_not ; n3208
g2953 and b[14] n3017_not ; n3209
g2954 and n3011_not n3209 ; n3210
g2955 and n3019_not n3210_not ; n3211
g2956 and n3208_not n3211 ; n3212
g2957 and n3019_not n3212_not ; n3213
g2958 and b[15] n3008_not ; n3214
g2959 and n3002_not n3214 ; n3215
g2960 and n3010_not n3215_not ; n3216
g2961 and n3213_not n3216 ; n3217
g2962 and n3010_not n3217_not ; n3218
g2963 and b[16] n2999_not ; n3219
g2964 and n2993_not n3219 ; n3220
g2965 and n3001_not n3220_not ; n3221
g2966 and n3218_not n3221 ; n3222
g2967 and n3001_not n3222_not ; n3223
g2968 and b[17] n2990_not ; n3224
g2969 and n2984_not n3224 ; n3225
g2970 and n2992_not n3225_not ; n3226
g2971 and n3223_not n3226 ; n3227
g2972 and n2992_not n3227_not ; n3228
g2973 and b[18] n2973_not ; n3229
g2974 and n2967_not n3229 ; n3230
g2975 and n2983_not n3230_not ; n3231
g2976 and n3228_not n3231 ; n3232
g2977 and n2983_not n3232_not ; n3233
g2978 and b[19] n2975_not ; n3234
g2979 and n2980_not n3234 ; n3235
g2980 and n2982_not n3235_not ; n3236
g2981 and n3233_not n3236 ; n3237
g2982 and n2982_not n3237_not ; n3238
g2983 and n320 n3238_not ; quotient[44]
g2984 and n2974_not quotient[44]_not ; n3240
g2985 and n2992_not n3231 ; n3241
g2986 and n3227_not n3241 ; n3242
g2987 and n3228_not n3231_not ; n3243
g2988 and n3242_not n3243_not ; n3244
g2989 and n320 n3244_not ; n3245
g2990 and n3238_not n3245 ; n3246
g2991 and n3240_not n3246_not ; n3247
g2992 and b[19]_not n3247_not ; n3248
g2993 and n2991_not quotient[44]_not ; n3249
g2994 and n3001_not n3226 ; n3250
g2995 and n3222_not n3250 ; n3251
g2996 and n3223_not n3226_not ; n3252
g2997 and n3251_not n3252_not ; n3253
g2998 and n320 n3253_not ; n3254
g2999 and n3238_not n3254 ; n3255
g3000 and n3249_not n3255_not ; n3256
g3001 and b[18]_not n3256_not ; n3257
g3002 and n3000_not quotient[44]_not ; n3258
g3003 and n3010_not n3221 ; n3259
g3004 and n3217_not n3259 ; n3260
g3005 and n3218_not n3221_not ; n3261
g3006 and n3260_not n3261_not ; n3262
g3007 and n320 n3262_not ; n3263
g3008 and n3238_not n3263 ; n3264
g3009 and n3258_not n3264_not ; n3265
g3010 and b[17]_not n3265_not ; n3266
g3011 and n3009_not quotient[44]_not ; n3267
g3012 and n3019_not n3216 ; n3268
g3013 and n3212_not n3268 ; n3269
g3014 and n3213_not n3216_not ; n3270
g3015 and n3269_not n3270_not ; n3271
g3016 and n320 n3271_not ; n3272
g3017 and n3238_not n3272 ; n3273
g3018 and n3267_not n3273_not ; n3274
g3019 and b[16]_not n3274_not ; n3275
g3020 and n3018_not quotient[44]_not ; n3276
g3021 and n3028_not n3211 ; n3277
g3022 and n3207_not n3277 ; n3278
g3023 and n3208_not n3211_not ; n3279
g3024 and n3278_not n3279_not ; n3280
g3025 and n320 n3280_not ; n3281
g3026 and n3238_not n3281 ; n3282
g3027 and n3276_not n3282_not ; n3283
g3028 and b[15]_not n3283_not ; n3284
g3029 and n3027_not quotient[44]_not ; n3285
g3030 and n3037_not n3206 ; n3286
g3031 and n3202_not n3286 ; n3287
g3032 and n3203_not n3206_not ; n3288
g3033 and n3287_not n3288_not ; n3289
g3034 and n320 n3289_not ; n3290
g3035 and n3238_not n3290 ; n3291
g3036 and n3285_not n3291_not ; n3292
g3037 and b[14]_not n3292_not ; n3293
g3038 and n3036_not quotient[44]_not ; n3294
g3039 and n3046_not n3201 ; n3295
g3040 and n3197_not n3295 ; n3296
g3041 and n3198_not n3201_not ; n3297
g3042 and n3296_not n3297_not ; n3298
g3043 and n320 n3298_not ; n3299
g3044 and n3238_not n3299 ; n3300
g3045 and n3294_not n3300_not ; n3301
g3046 and b[13]_not n3301_not ; n3302
g3047 and n3045_not quotient[44]_not ; n3303
g3048 and n3055_not n3196 ; n3304
g3049 and n3192_not n3304 ; n3305
g3050 and n3193_not n3196_not ; n3306
g3051 and n3305_not n3306_not ; n3307
g3052 and n320 n3307_not ; n3308
g3053 and n3238_not n3308 ; n3309
g3054 and n3303_not n3309_not ; n3310
g3055 and b[12]_not n3310_not ; n3311
g3056 and n3054_not quotient[44]_not ; n3312
g3057 and n3064_not n3191 ; n3313
g3058 and n3187_not n3313 ; n3314
g3059 and n3188_not n3191_not ; n3315
g3060 and n3314_not n3315_not ; n3316
g3061 and n320 n3316_not ; n3317
g3062 and n3238_not n3317 ; n3318
g3063 and n3312_not n3318_not ; n3319
g3064 and b[11]_not n3319_not ; n3320
g3065 and n3063_not quotient[44]_not ; n3321
g3066 and n3073_not n3186 ; n3322
g3067 and n3182_not n3322 ; n3323
g3068 and n3183_not n3186_not ; n3324
g3069 and n3323_not n3324_not ; n3325
g3070 and n320 n3325_not ; n3326
g3071 and n3238_not n3326 ; n3327
g3072 and n3321_not n3327_not ; n3328
g3073 and b[10]_not n3328_not ; n3329
g3074 and n3072_not quotient[44]_not ; n3330
g3075 and n3082_not n3181 ; n3331
g3076 and n3177_not n3331 ; n3332
g3077 and n3178_not n3181_not ; n3333
g3078 and n3332_not n3333_not ; n3334
g3079 and n320 n3334_not ; n3335
g3080 and n3238_not n3335 ; n3336
g3081 and n3330_not n3336_not ; n3337
g3082 and b[9]_not n3337_not ; n3338
g3083 and n3081_not quotient[44]_not ; n3339
g3084 and n3091_not n3176 ; n3340
g3085 and n3172_not n3340 ; n3341
g3086 and n3173_not n3176_not ; n3342
g3087 and n3341_not n3342_not ; n3343
g3088 and n320 n3343_not ; n3344
g3089 and n3238_not n3344 ; n3345
g3090 and n3339_not n3345_not ; n3346
g3091 and b[8]_not n3346_not ; n3347
g3092 and n3090_not quotient[44]_not ; n3348
g3093 and n3100_not n3171 ; n3349
g3094 and n3167_not n3349 ; n3350
g3095 and n3168_not n3171_not ; n3351
g3096 and n3350_not n3351_not ; n3352
g3097 and n320 n3352_not ; n3353
g3098 and n3238_not n3353 ; n3354
g3099 and n3348_not n3354_not ; n3355
g3100 and b[7]_not n3355_not ; n3356
g3101 and n3099_not quotient[44]_not ; n3357
g3102 and n3109_not n3166 ; n3358
g3103 and n3162_not n3358 ; n3359
g3104 and n3163_not n3166_not ; n3360
g3105 and n3359_not n3360_not ; n3361
g3106 and n320 n3361_not ; n3362
g3107 and n3238_not n3362 ; n3363
g3108 and n3357_not n3363_not ; n3364
g3109 and b[6]_not n3364_not ; n3365
g3110 and n3108_not quotient[44]_not ; n3366
g3111 and n3118_not n3161 ; n3367
g3112 and n3157_not n3367 ; n3368
g3113 and n3158_not n3161_not ; n3369
g3114 and n3368_not n3369_not ; n3370
g3115 and n320 n3370_not ; n3371
g3116 and n3238_not n3371 ; n3372
g3117 and n3366_not n3372_not ; n3373
g3118 and b[5]_not n3373_not ; n3374
g3119 and n3117_not quotient[44]_not ; n3375
g3120 and n3126_not n3156 ; n3376
g3121 and n3152_not n3376 ; n3377
g3122 and n3153_not n3156_not ; n3378
g3123 and n3377_not n3378_not ; n3379
g3124 and n320 n3379_not ; n3380
g3125 and n3238_not n3380 ; n3381
g3126 and n3375_not n3381_not ; n3382
g3127 and b[4]_not n3382_not ; n3383
g3128 and n3125_not quotient[44]_not ; n3384
g3129 and n3147_not n3151 ; n3385
g3130 and n3146_not n3385 ; n3386
g3131 and n3148_not n3151_not ; n3387
g3132 and n3386_not n3387_not ; n3388
g3133 and n320 n3388_not ; n3389
g3134 and n3238_not n3389 ; n3390
g3135 and n3384_not n3390_not ; n3391
g3136 and b[3]_not n3391_not ; n3392
g3137 and n3140_not quotient[44]_not ; n3393
g3138 and n3143_not n3145 ; n3394
g3139 and n3141_not n3394 ; n3395
g3140 and n320 n3395_not ; n3396
g3141 and n3146_not n3396 ; n3397
g3142 and n3238_not n3397 ; n3398
g3143 and n3393_not n3398_not ; n3399
g3144 and b[2]_not n3399_not ; n3400
g3145 and b[0] b[20]_not ; n3401
g3146 and n366 n3401 ; n3402
g3147 and n377 n3402 ; n3403
g3148 and n423 n3403 ; n3404
g3149 and n408 n3404 ; n3405
g3150 and n3238_not n3405 ; n3406
g3151 and a[44] n3406_not ; n3407
g3152 and n309 n3145 ; n3408
g3153 and n343 n3408 ; n3409
g3154 and n341 n3409 ; n3410
g3155 and n338 n3410 ; n3411
g3156 and n3238_not n3411 ; n3412
g3157 and n3407_not n3412_not ; n3413
g3158 and b[1] n3413_not ; n3414
g3159 and b[1]_not n3412_not ; n3415
g3160 and n3407_not n3415 ; n3416
g3161 and n3414_not n3416_not ; n3417
g3162 and a[43]_not b[0] ; n3418
g3163 and n3417_not n3418_not ; n3419
g3164 and b[1]_not n3413_not ; n3420
g3165 and n3419_not n3420_not ; n3421
g3166 and b[2] n3398_not ; n3422
g3167 and n3393_not n3422 ; n3423
g3168 and n3400_not n3423_not ; n3424
g3169 and n3421_not n3424 ; n3425
g3170 and n3400_not n3425_not ; n3426
g3171 and b[3] n3390_not ; n3427
g3172 and n3384_not n3427 ; n3428
g3173 and n3392_not n3428_not ; n3429
g3174 and n3426_not n3429 ; n3430
g3175 and n3392_not n3430_not ; n3431
g3176 and b[4] n3381_not ; n3432
g3177 and n3375_not n3432 ; n3433
g3178 and n3383_not n3433_not ; n3434
g3179 and n3431_not n3434 ; n3435
g3180 and n3383_not n3435_not ; n3436
g3181 and b[5] n3372_not ; n3437
g3182 and n3366_not n3437 ; n3438
g3183 and n3374_not n3438_not ; n3439
g3184 and n3436_not n3439 ; n3440
g3185 and n3374_not n3440_not ; n3441
g3186 and b[6] n3363_not ; n3442
g3187 and n3357_not n3442 ; n3443
g3188 and n3365_not n3443_not ; n3444
g3189 and n3441_not n3444 ; n3445
g3190 and n3365_not n3445_not ; n3446
g3191 and b[7] n3354_not ; n3447
g3192 and n3348_not n3447 ; n3448
g3193 and n3356_not n3448_not ; n3449
g3194 and n3446_not n3449 ; n3450
g3195 and n3356_not n3450_not ; n3451
g3196 and b[8] n3345_not ; n3452
g3197 and n3339_not n3452 ; n3453
g3198 and n3347_not n3453_not ; n3454
g3199 and n3451_not n3454 ; n3455
g3200 and n3347_not n3455_not ; n3456
g3201 and b[9] n3336_not ; n3457
g3202 and n3330_not n3457 ; n3458
g3203 and n3338_not n3458_not ; n3459
g3204 and n3456_not n3459 ; n3460
g3205 and n3338_not n3460_not ; n3461
g3206 and b[10] n3327_not ; n3462
g3207 and n3321_not n3462 ; n3463
g3208 and n3329_not n3463_not ; n3464
g3209 and n3461_not n3464 ; n3465
g3210 and n3329_not n3465_not ; n3466
g3211 and b[11] n3318_not ; n3467
g3212 and n3312_not n3467 ; n3468
g3213 and n3320_not n3468_not ; n3469
g3214 and n3466_not n3469 ; n3470
g3215 and n3320_not n3470_not ; n3471
g3216 and b[12] n3309_not ; n3472
g3217 and n3303_not n3472 ; n3473
g3218 and n3311_not n3473_not ; n3474
g3219 and n3471_not n3474 ; n3475
g3220 and n3311_not n3475_not ; n3476
g3221 and b[13] n3300_not ; n3477
g3222 and n3294_not n3477 ; n3478
g3223 and n3302_not n3478_not ; n3479
g3224 and n3476_not n3479 ; n3480
g3225 and n3302_not n3480_not ; n3481
g3226 and b[14] n3291_not ; n3482
g3227 and n3285_not n3482 ; n3483
g3228 and n3293_not n3483_not ; n3484
g3229 and n3481_not n3484 ; n3485
g3230 and n3293_not n3485_not ; n3486
g3231 and b[15] n3282_not ; n3487
g3232 and n3276_not n3487 ; n3488
g3233 and n3284_not n3488_not ; n3489
g3234 and n3486_not n3489 ; n3490
g3235 and n3284_not n3490_not ; n3491
g3236 and b[16] n3273_not ; n3492
g3237 and n3267_not n3492 ; n3493
g3238 and n3275_not n3493_not ; n3494
g3239 and n3491_not n3494 ; n3495
g3240 and n3275_not n3495_not ; n3496
g3241 and b[17] n3264_not ; n3497
g3242 and n3258_not n3497 ; n3498
g3243 and n3266_not n3498_not ; n3499
g3244 and n3496_not n3499 ; n3500
g3245 and n3266_not n3500_not ; n3501
g3246 and b[18] n3255_not ; n3502
g3247 and n3249_not n3502 ; n3503
g3248 and n3257_not n3503_not ; n3504
g3249 and n3501_not n3504 ; n3505
g3250 and n3257_not n3505_not ; n3506
g3251 and b[19] n3246_not ; n3507
g3252 and n3240_not n3507 ; n3508
g3253 and n3248_not n3508_not ; n3509
g3254 and n3506_not n3509 ; n3510
g3255 and n3248_not n3510_not ; n3511
g3256 and n2981_not quotient[44]_not ; n3512
g3257 and n2983_not n3236 ; n3513
g3258 and n3232_not n3513 ; n3514
g3259 and n3233_not n3236_not ; n3515
g3260 and n3514_not n3515_not ; n3516
g3261 and quotient[44] n3516_not ; n3517
g3262 and n3512_not n3517_not ; n3518
g3263 and b[20]_not n3518_not ; n3519
g3264 and b[20] n3512_not ; n3520
g3265 and n3517_not n3520 ; n3521
g3266 and n643 n3521_not ; n3522
g3267 and n3519_not n3522 ; n3523
g3268 and n3511_not n3523 ; n3524
g3269 and n320 n3518_not ; n3525
g3270 and n3524_not n3525_not ; quotient[43]
g3271 and n3257_not n3509 ; n3527
g3272 and n3505_not n3527 ; n3528
g3273 and n3506_not n3509_not ; n3529
g3274 and n3528_not n3529_not ; n3530
g3275 and quotient[43] n3530_not ; n3531
g3276 and n3247_not n3525_not ; n3532
g3277 and n3524_not n3532 ; n3533
g3278 and n3531_not n3533_not ; n3534
g3279 and n3248_not n3521_not ; n3535
g3280 and n3519_not n3535 ; n3536
g3281 and n3510_not n3536 ; n3537
g3282 and n3519_not n3521_not ; n3538
g3283 and n3511_not n3538_not ; n3539
g3284 and n3537_not n3539_not ; n3540
g3285 and quotient[43] n3540_not ; n3541
g3286 and n3518_not n3525_not ; n3542
g3287 and n3524_not n3542 ; n3543
g3288 and n3541_not n3543_not ; n3544
g3289 and b[21]_not n3544_not ; n3545
g3290 and b[20]_not n3534_not ; n3546
g3291 and n3266_not n3504 ; n3547
g3292 and n3500_not n3547 ; n3548
g3293 and n3501_not n3504_not ; n3549
g3294 and n3548_not n3549_not ; n3550
g3295 and quotient[43] n3550_not ; n3551
g3296 and n3256_not n3525_not ; n3552
g3297 and n3524_not n3552 ; n3553
g3298 and n3551_not n3553_not ; n3554
g3299 and b[19]_not n3554_not ; n3555
g3300 and n3275_not n3499 ; n3556
g3301 and n3495_not n3556 ; n3557
g3302 and n3496_not n3499_not ; n3558
g3303 and n3557_not n3558_not ; n3559
g3304 and quotient[43] n3559_not ; n3560
g3305 and n3265_not n3525_not ; n3561
g3306 and n3524_not n3561 ; n3562
g3307 and n3560_not n3562_not ; n3563
g3308 and b[18]_not n3563_not ; n3564
g3309 and n3284_not n3494 ; n3565
g3310 and n3490_not n3565 ; n3566
g3311 and n3491_not n3494_not ; n3567
g3312 and n3566_not n3567_not ; n3568
g3313 and quotient[43] n3568_not ; n3569
g3314 and n3274_not n3525_not ; n3570
g3315 and n3524_not n3570 ; n3571
g3316 and n3569_not n3571_not ; n3572
g3317 and b[17]_not n3572_not ; n3573
g3318 and n3293_not n3489 ; n3574
g3319 and n3485_not n3574 ; n3575
g3320 and n3486_not n3489_not ; n3576
g3321 and n3575_not n3576_not ; n3577
g3322 and quotient[43] n3577_not ; n3578
g3323 and n3283_not n3525_not ; n3579
g3324 and n3524_not n3579 ; n3580
g3325 and n3578_not n3580_not ; n3581
g3326 and b[16]_not n3581_not ; n3582
g3327 and n3302_not n3484 ; n3583
g3328 and n3480_not n3583 ; n3584
g3329 and n3481_not n3484_not ; n3585
g3330 and n3584_not n3585_not ; n3586
g3331 and quotient[43] n3586_not ; n3587
g3332 and n3292_not n3525_not ; n3588
g3333 and n3524_not n3588 ; n3589
g3334 and n3587_not n3589_not ; n3590
g3335 and b[15]_not n3590_not ; n3591
g3336 and n3311_not n3479 ; n3592
g3337 and n3475_not n3592 ; n3593
g3338 and n3476_not n3479_not ; n3594
g3339 and n3593_not n3594_not ; n3595
g3340 and quotient[43] n3595_not ; n3596
g3341 and n3301_not n3525_not ; n3597
g3342 and n3524_not n3597 ; n3598
g3343 and n3596_not n3598_not ; n3599
g3344 and b[14]_not n3599_not ; n3600
g3345 and n3320_not n3474 ; n3601
g3346 and n3470_not n3601 ; n3602
g3347 and n3471_not n3474_not ; n3603
g3348 and n3602_not n3603_not ; n3604
g3349 and quotient[43] n3604_not ; n3605
g3350 and n3310_not n3525_not ; n3606
g3351 and n3524_not n3606 ; n3607
g3352 and n3605_not n3607_not ; n3608
g3353 and b[13]_not n3608_not ; n3609
g3354 and n3329_not n3469 ; n3610
g3355 and n3465_not n3610 ; n3611
g3356 and n3466_not n3469_not ; n3612
g3357 and n3611_not n3612_not ; n3613
g3358 and quotient[43] n3613_not ; n3614
g3359 and n3319_not n3525_not ; n3615
g3360 and n3524_not n3615 ; n3616
g3361 and n3614_not n3616_not ; n3617
g3362 and b[12]_not n3617_not ; n3618
g3363 and n3338_not n3464 ; n3619
g3364 and n3460_not n3619 ; n3620
g3365 and n3461_not n3464_not ; n3621
g3366 and n3620_not n3621_not ; n3622
g3367 and quotient[43] n3622_not ; n3623
g3368 and n3328_not n3525_not ; n3624
g3369 and n3524_not n3624 ; n3625
g3370 and n3623_not n3625_not ; n3626
g3371 and b[11]_not n3626_not ; n3627
g3372 and n3347_not n3459 ; n3628
g3373 and n3455_not n3628 ; n3629
g3374 and n3456_not n3459_not ; n3630
g3375 and n3629_not n3630_not ; n3631
g3376 and quotient[43] n3631_not ; n3632
g3377 and n3337_not n3525_not ; n3633
g3378 and n3524_not n3633 ; n3634
g3379 and n3632_not n3634_not ; n3635
g3380 and b[10]_not n3635_not ; n3636
g3381 and n3356_not n3454 ; n3637
g3382 and n3450_not n3637 ; n3638
g3383 and n3451_not n3454_not ; n3639
g3384 and n3638_not n3639_not ; n3640
g3385 and quotient[43] n3640_not ; n3641
g3386 and n3346_not n3525_not ; n3642
g3387 and n3524_not n3642 ; n3643
g3388 and n3641_not n3643_not ; n3644
g3389 and b[9]_not n3644_not ; n3645
g3390 and n3365_not n3449 ; n3646
g3391 and n3445_not n3646 ; n3647
g3392 and n3446_not n3449_not ; n3648
g3393 and n3647_not n3648_not ; n3649
g3394 and quotient[43] n3649_not ; n3650
g3395 and n3355_not n3525_not ; n3651
g3396 and n3524_not n3651 ; n3652
g3397 and n3650_not n3652_not ; n3653
g3398 and b[8]_not n3653_not ; n3654
g3399 and n3374_not n3444 ; n3655
g3400 and n3440_not n3655 ; n3656
g3401 and n3441_not n3444_not ; n3657
g3402 and n3656_not n3657_not ; n3658
g3403 and quotient[43] n3658_not ; n3659
g3404 and n3364_not n3525_not ; n3660
g3405 and n3524_not n3660 ; n3661
g3406 and n3659_not n3661_not ; n3662
g3407 and b[7]_not n3662_not ; n3663
g3408 and n3383_not n3439 ; n3664
g3409 and n3435_not n3664 ; n3665
g3410 and n3436_not n3439_not ; n3666
g3411 and n3665_not n3666_not ; n3667
g3412 and quotient[43] n3667_not ; n3668
g3413 and n3373_not n3525_not ; n3669
g3414 and n3524_not n3669 ; n3670
g3415 and n3668_not n3670_not ; n3671
g3416 and b[6]_not n3671_not ; n3672
g3417 and n3392_not n3434 ; n3673
g3418 and n3430_not n3673 ; n3674
g3419 and n3431_not n3434_not ; n3675
g3420 and n3674_not n3675_not ; n3676
g3421 and quotient[43] n3676_not ; n3677
g3422 and n3382_not n3525_not ; n3678
g3423 and n3524_not n3678 ; n3679
g3424 and n3677_not n3679_not ; n3680
g3425 and b[5]_not n3680_not ; n3681
g3426 and n3400_not n3429 ; n3682
g3427 and n3425_not n3682 ; n3683
g3428 and n3426_not n3429_not ; n3684
g3429 and n3683_not n3684_not ; n3685
g3430 and quotient[43] n3685_not ; n3686
g3431 and n3391_not n3525_not ; n3687
g3432 and n3524_not n3687 ; n3688
g3433 and n3686_not n3688_not ; n3689
g3434 and b[4]_not n3689_not ; n3690
g3435 and n3420_not n3424 ; n3691
g3436 and n3419_not n3691 ; n3692
g3437 and n3421_not n3424_not ; n3693
g3438 and n3692_not n3693_not ; n3694
g3439 and quotient[43] n3694_not ; n3695
g3440 and n3399_not n3525_not ; n3696
g3441 and n3524_not n3696 ; n3697
g3442 and n3695_not n3697_not ; n3698
g3443 and b[3]_not n3698_not ; n3699
g3444 and n3416_not n3418 ; n3700
g3445 and n3414_not n3700 ; n3701
g3446 and n3419_not n3701_not ; n3702
g3447 and quotient[43] n3702 ; n3703
g3448 and n3413_not n3525_not ; n3704
g3449 and n3524_not n3704 ; n3705
g3450 and n3703_not n3705_not ; n3706
g3451 and b[2]_not n3706_not ; n3707
g3452 and b[0] quotient[43] ; n3708
g3453 and a[43] n3708_not ; n3709
g3454 and n3418 quotient[43] ; n3710
g3455 and n3709_not n3710_not ; n3711
g3456 and b[1] n3711_not ; n3712
g3457 and b[1]_not n3710_not ; n3713
g3458 and n3709_not n3713 ; n3714
g3459 and n3712_not n3714_not ; n3715
g3460 and a[42]_not b[0] ; n3716
g3461 and n3715_not n3716_not ; n3717
g3462 and b[1]_not n3711_not ; n3718
g3463 and n3717_not n3718_not ; n3719
g3464 and b[2] n3705_not ; n3720
g3465 and n3703_not n3720 ; n3721
g3466 and n3707_not n3721_not ; n3722
g3467 and n3719_not n3722 ; n3723
g3468 and n3707_not n3723_not ; n3724
g3469 and b[3] n3697_not ; n3725
g3470 and n3695_not n3725 ; n3726
g3471 and n3699_not n3726_not ; n3727
g3472 and n3724_not n3727 ; n3728
g3473 and n3699_not n3728_not ; n3729
g3474 and b[4] n3688_not ; n3730
g3475 and n3686_not n3730 ; n3731
g3476 and n3690_not n3731_not ; n3732
g3477 and n3729_not n3732 ; n3733
g3478 and n3690_not n3733_not ; n3734
g3479 and b[5] n3679_not ; n3735
g3480 and n3677_not n3735 ; n3736
g3481 and n3681_not n3736_not ; n3737
g3482 and n3734_not n3737 ; n3738
g3483 and n3681_not n3738_not ; n3739
g3484 and b[6] n3670_not ; n3740
g3485 and n3668_not n3740 ; n3741
g3486 and n3672_not n3741_not ; n3742
g3487 and n3739_not n3742 ; n3743
g3488 and n3672_not n3743_not ; n3744
g3489 and b[7] n3661_not ; n3745
g3490 and n3659_not n3745 ; n3746
g3491 and n3663_not n3746_not ; n3747
g3492 and n3744_not n3747 ; n3748
g3493 and n3663_not n3748_not ; n3749
g3494 and b[8] n3652_not ; n3750
g3495 and n3650_not n3750 ; n3751
g3496 and n3654_not n3751_not ; n3752
g3497 and n3749_not n3752 ; n3753
g3498 and n3654_not n3753_not ; n3754
g3499 and b[9] n3643_not ; n3755
g3500 and n3641_not n3755 ; n3756
g3501 and n3645_not n3756_not ; n3757
g3502 and n3754_not n3757 ; n3758
g3503 and n3645_not n3758_not ; n3759
g3504 and b[10] n3634_not ; n3760
g3505 and n3632_not n3760 ; n3761
g3506 and n3636_not n3761_not ; n3762
g3507 and n3759_not n3762 ; n3763
g3508 and n3636_not n3763_not ; n3764
g3509 and b[11] n3625_not ; n3765
g3510 and n3623_not n3765 ; n3766
g3511 and n3627_not n3766_not ; n3767
g3512 and n3764_not n3767 ; n3768
g3513 and n3627_not n3768_not ; n3769
g3514 and b[12] n3616_not ; n3770
g3515 and n3614_not n3770 ; n3771
g3516 and n3618_not n3771_not ; n3772
g3517 and n3769_not n3772 ; n3773
g3518 and n3618_not n3773_not ; n3774
g3519 and b[13] n3607_not ; n3775
g3520 and n3605_not n3775 ; n3776
g3521 and n3609_not n3776_not ; n3777
g3522 and n3774_not n3777 ; n3778
g3523 and n3609_not n3778_not ; n3779
g3524 and b[14] n3598_not ; n3780
g3525 and n3596_not n3780 ; n3781
g3526 and n3600_not n3781_not ; n3782
g3527 and n3779_not n3782 ; n3783
g3528 and n3600_not n3783_not ; n3784
g3529 and b[15] n3589_not ; n3785
g3530 and n3587_not n3785 ; n3786
g3531 and n3591_not n3786_not ; n3787
g3532 and n3784_not n3787 ; n3788
g3533 and n3591_not n3788_not ; n3789
g3534 and b[16] n3580_not ; n3790
g3535 and n3578_not n3790 ; n3791
g3536 and n3582_not n3791_not ; n3792
g3537 and n3789_not n3792 ; n3793
g3538 and n3582_not n3793_not ; n3794
g3539 and b[17] n3571_not ; n3795
g3540 and n3569_not n3795 ; n3796
g3541 and n3573_not n3796_not ; n3797
g3542 and n3794_not n3797 ; n3798
g3543 and n3573_not n3798_not ; n3799
g3544 and b[18] n3562_not ; n3800
g3545 and n3560_not n3800 ; n3801
g3546 and n3564_not n3801_not ; n3802
g3547 and n3799_not n3802 ; n3803
g3548 and n3564_not n3803_not ; n3804
g3549 and b[19] n3553_not ; n3805
g3550 and n3551_not n3805 ; n3806
g3551 and n3555_not n3806_not ; n3807
g3552 and n3804_not n3807 ; n3808
g3553 and n3555_not n3808_not ; n3809
g3554 and b[20] n3533_not ; n3810
g3555 and n3531_not n3810 ; n3811
g3556 and n3546_not n3811_not ; n3812
g3557 and n3809_not n3812 ; n3813
g3558 and n3546_not n3813_not ; n3814
g3559 and b[21] n3543_not ; n3815
g3560 and n3541_not n3815 ; n3816
g3561 and n3545_not n3816_not ; n3817
g3562 and n3814_not n3817 ; n3818
g3563 and n3545_not n3818_not ; n3819
g3564 and n306 n308 ; n3820
g3565 and n317 n3820 ; n3821
g3566 and n303 n3821 ; n3822
g3567 and n288 n3822 ; n3823
g3568 and n3819_not n3823 ; quotient[42]
g3569 and n3534_not quotient[42]_not ; n3825
g3570 and n3555_not n3812 ; n3826
g3571 and n3808_not n3826 ; n3827
g3572 and n3809_not n3812_not ; n3828
g3573 and n3827_not n3828_not ; n3829
g3574 and n3823 n3829_not ; n3830
g3575 and n3819_not n3830 ; n3831
g3576 and n3825_not n3831_not ; n3832
g3577 and n3544_not quotient[42]_not ; n3833
g3578 and n3546_not n3817 ; n3834
g3579 and n3813_not n3834 ; n3835
g3580 and n3814_not n3817_not ; n3836
g3581 and n3835_not n3836_not ; n3837
g3582 and quotient[42] n3837_not ; n3838
g3583 and n3833_not n3838_not ; n3839
g3584 and b[22]_not n3839_not ; n3840
g3585 and b[21]_not n3832_not ; n3841
g3586 and n3554_not quotient[42]_not ; n3842
g3587 and n3564_not n3807 ; n3843
g3588 and n3803_not n3843 ; n3844
g3589 and n3804_not n3807_not ; n3845
g3590 and n3844_not n3845_not ; n3846
g3591 and n3823 n3846_not ; n3847
g3592 and n3819_not n3847 ; n3848
g3593 and n3842_not n3848_not ; n3849
g3594 and b[20]_not n3849_not ; n3850
g3595 and n3563_not quotient[42]_not ; n3851
g3596 and n3573_not n3802 ; n3852
g3597 and n3798_not n3852 ; n3853
g3598 and n3799_not n3802_not ; n3854
g3599 and n3853_not n3854_not ; n3855
g3600 and n3823 n3855_not ; n3856
g3601 and n3819_not n3856 ; n3857
g3602 and n3851_not n3857_not ; n3858
g3603 and b[19]_not n3858_not ; n3859
g3604 and n3572_not quotient[42]_not ; n3860
g3605 and n3582_not n3797 ; n3861
g3606 and n3793_not n3861 ; n3862
g3607 and n3794_not n3797_not ; n3863
g3608 and n3862_not n3863_not ; n3864
g3609 and n3823 n3864_not ; n3865
g3610 and n3819_not n3865 ; n3866
g3611 and n3860_not n3866_not ; n3867
g3612 and b[18]_not n3867_not ; n3868
g3613 and n3581_not quotient[42]_not ; n3869
g3614 and n3591_not n3792 ; n3870
g3615 and n3788_not n3870 ; n3871
g3616 and n3789_not n3792_not ; n3872
g3617 and n3871_not n3872_not ; n3873
g3618 and n3823 n3873_not ; n3874
g3619 and n3819_not n3874 ; n3875
g3620 and n3869_not n3875_not ; n3876
g3621 and b[17]_not n3876_not ; n3877
g3622 and n3590_not quotient[42]_not ; n3878
g3623 and n3600_not n3787 ; n3879
g3624 and n3783_not n3879 ; n3880
g3625 and n3784_not n3787_not ; n3881
g3626 and n3880_not n3881_not ; n3882
g3627 and n3823 n3882_not ; n3883
g3628 and n3819_not n3883 ; n3884
g3629 and n3878_not n3884_not ; n3885
g3630 and b[16]_not n3885_not ; n3886
g3631 and n3599_not quotient[42]_not ; n3887
g3632 and n3609_not n3782 ; n3888
g3633 and n3778_not n3888 ; n3889
g3634 and n3779_not n3782_not ; n3890
g3635 and n3889_not n3890_not ; n3891
g3636 and n3823 n3891_not ; n3892
g3637 and n3819_not n3892 ; n3893
g3638 and n3887_not n3893_not ; n3894
g3639 and b[15]_not n3894_not ; n3895
g3640 and n3608_not quotient[42]_not ; n3896
g3641 and n3618_not n3777 ; n3897
g3642 and n3773_not n3897 ; n3898
g3643 and n3774_not n3777_not ; n3899
g3644 and n3898_not n3899_not ; n3900
g3645 and n3823 n3900_not ; n3901
g3646 and n3819_not n3901 ; n3902
g3647 and n3896_not n3902_not ; n3903
g3648 and b[14]_not n3903_not ; n3904
g3649 and n3617_not quotient[42]_not ; n3905
g3650 and n3627_not n3772 ; n3906
g3651 and n3768_not n3906 ; n3907
g3652 and n3769_not n3772_not ; n3908
g3653 and n3907_not n3908_not ; n3909
g3654 and n3823 n3909_not ; n3910
g3655 and n3819_not n3910 ; n3911
g3656 and n3905_not n3911_not ; n3912
g3657 and b[13]_not n3912_not ; n3913
g3658 and n3626_not quotient[42]_not ; n3914
g3659 and n3636_not n3767 ; n3915
g3660 and n3763_not n3915 ; n3916
g3661 and n3764_not n3767_not ; n3917
g3662 and n3916_not n3917_not ; n3918
g3663 and n3823 n3918_not ; n3919
g3664 and n3819_not n3919 ; n3920
g3665 and n3914_not n3920_not ; n3921
g3666 and b[12]_not n3921_not ; n3922
g3667 and n3635_not quotient[42]_not ; n3923
g3668 and n3645_not n3762 ; n3924
g3669 and n3758_not n3924 ; n3925
g3670 and n3759_not n3762_not ; n3926
g3671 and n3925_not n3926_not ; n3927
g3672 and n3823 n3927_not ; n3928
g3673 and n3819_not n3928 ; n3929
g3674 and n3923_not n3929_not ; n3930
g3675 and b[11]_not n3930_not ; n3931
g3676 and n3644_not quotient[42]_not ; n3932
g3677 and n3654_not n3757 ; n3933
g3678 and n3753_not n3933 ; n3934
g3679 and n3754_not n3757_not ; n3935
g3680 and n3934_not n3935_not ; n3936
g3681 and n3823 n3936_not ; n3937
g3682 and n3819_not n3937 ; n3938
g3683 and n3932_not n3938_not ; n3939
g3684 and b[10]_not n3939_not ; n3940
g3685 and n3653_not quotient[42]_not ; n3941
g3686 and n3663_not n3752 ; n3942
g3687 and n3748_not n3942 ; n3943
g3688 and n3749_not n3752_not ; n3944
g3689 and n3943_not n3944_not ; n3945
g3690 and n3823 n3945_not ; n3946
g3691 and n3819_not n3946 ; n3947
g3692 and n3941_not n3947_not ; n3948
g3693 and b[9]_not n3948_not ; n3949
g3694 and n3662_not quotient[42]_not ; n3950
g3695 and n3672_not n3747 ; n3951
g3696 and n3743_not n3951 ; n3952
g3697 and n3744_not n3747_not ; n3953
g3698 and n3952_not n3953_not ; n3954
g3699 and n3823 n3954_not ; n3955
g3700 and n3819_not n3955 ; n3956
g3701 and n3950_not n3956_not ; n3957
g3702 and b[8]_not n3957_not ; n3958
g3703 and n3671_not quotient[42]_not ; n3959
g3704 and n3681_not n3742 ; n3960
g3705 and n3738_not n3960 ; n3961
g3706 and n3739_not n3742_not ; n3962
g3707 and n3961_not n3962_not ; n3963
g3708 and n3823 n3963_not ; n3964
g3709 and n3819_not n3964 ; n3965
g3710 and n3959_not n3965_not ; n3966
g3711 and b[7]_not n3966_not ; n3967
g3712 and n3680_not quotient[42]_not ; n3968
g3713 and n3690_not n3737 ; n3969
g3714 and n3733_not n3969 ; n3970
g3715 and n3734_not n3737_not ; n3971
g3716 and n3970_not n3971_not ; n3972
g3717 and n3823 n3972_not ; n3973
g3718 and n3819_not n3973 ; n3974
g3719 and n3968_not n3974_not ; n3975
g3720 and b[6]_not n3975_not ; n3976
g3721 and n3689_not quotient[42]_not ; n3977
g3722 and n3699_not n3732 ; n3978
g3723 and n3728_not n3978 ; n3979
g3724 and n3729_not n3732_not ; n3980
g3725 and n3979_not n3980_not ; n3981
g3726 and n3823 n3981_not ; n3982
g3727 and n3819_not n3982 ; n3983
g3728 and n3977_not n3983_not ; n3984
g3729 and b[5]_not n3984_not ; n3985
g3730 and n3698_not quotient[42]_not ; n3986
g3731 and n3707_not n3727 ; n3987
g3732 and n3723_not n3987 ; n3988
g3733 and n3724_not n3727_not ; n3989
g3734 and n3988_not n3989_not ; n3990
g3735 and n3823 n3990_not ; n3991
g3736 and n3819_not n3991 ; n3992
g3737 and n3986_not n3992_not ; n3993
g3738 and b[4]_not n3993_not ; n3994
g3739 and n3706_not quotient[42]_not ; n3995
g3740 and n3718_not n3722 ; n3996
g3741 and n3717_not n3996 ; n3997
g3742 and n3719_not n3722_not ; n3998
g3743 and n3997_not n3998_not ; n3999
g3744 and n3823 n3999_not ; n4000
g3745 and n3819_not n4000 ; n4001
g3746 and n3995_not n4001_not ; n4002
g3747 and b[3]_not n4002_not ; n4003
g3748 and n3711_not quotient[42]_not ; n4004
g3749 and n3714_not n3716 ; n4005
g3750 and n3712_not n4005 ; n4006
g3751 and n3823 n4006_not ; n4007
g3752 and n3717_not n4007 ; n4008
g3753 and n3819_not n4008 ; n4009
g3754 and n4004_not n4009_not ; n4010
g3755 and b[2]_not n4010_not ; n4011
g3756 and b[0] b[22]_not ; n4012
g3757 and n365 n4012 ; n4013
g3758 and n376 n4013 ; n4014
g3759 and n588 n4014 ; n4015
g3760 and n598 n4015 ; n4016
g3761 and n595 n4016 ; n4017
g3762 and n3819_not n4017 ; n4018
g3763 and a[42] n4018_not ; n4019
g3764 and n308 n3716 ; n4020
g3765 and n306 n4020 ; n4021
g3766 and n317 n4021 ; n4022
g3767 and n303 n4022 ; n4023
g3768 and n288 n4023 ; n4024
g3769 and n3819_not n4024 ; n4025
g3770 and n4019_not n4025_not ; n4026
g3771 and b[1] n4026_not ; n4027
g3772 and b[1]_not n4025_not ; n4028
g3773 and n4019_not n4028 ; n4029
g3774 and n4027_not n4029_not ; n4030
g3775 and a[41]_not b[0] ; n4031
g3776 and n4030_not n4031_not ; n4032
g3777 and b[1]_not n4026_not ; n4033
g3778 and n4032_not n4033_not ; n4034
g3779 and b[2] n4009_not ; n4035
g3780 and n4004_not n4035 ; n4036
g3781 and n4011_not n4036_not ; n4037
g3782 and n4034_not n4037 ; n4038
g3783 and n4011_not n4038_not ; n4039
g3784 and b[3] n4001_not ; n4040
g3785 and n3995_not n4040 ; n4041
g3786 and n4003_not n4041_not ; n4042
g3787 and n4039_not n4042 ; n4043
g3788 and n4003_not n4043_not ; n4044
g3789 and b[4] n3992_not ; n4045
g3790 and n3986_not n4045 ; n4046
g3791 and n3994_not n4046_not ; n4047
g3792 and n4044_not n4047 ; n4048
g3793 and n3994_not n4048_not ; n4049
g3794 and b[5] n3983_not ; n4050
g3795 and n3977_not n4050 ; n4051
g3796 and n3985_not n4051_not ; n4052
g3797 and n4049_not n4052 ; n4053
g3798 and n3985_not n4053_not ; n4054
g3799 and b[6] n3974_not ; n4055
g3800 and n3968_not n4055 ; n4056
g3801 and n3976_not n4056_not ; n4057
g3802 and n4054_not n4057 ; n4058
g3803 and n3976_not n4058_not ; n4059
g3804 and b[7] n3965_not ; n4060
g3805 and n3959_not n4060 ; n4061
g3806 and n3967_not n4061_not ; n4062
g3807 and n4059_not n4062 ; n4063
g3808 and n3967_not n4063_not ; n4064
g3809 and b[8] n3956_not ; n4065
g3810 and n3950_not n4065 ; n4066
g3811 and n3958_not n4066_not ; n4067
g3812 and n4064_not n4067 ; n4068
g3813 and n3958_not n4068_not ; n4069
g3814 and b[9] n3947_not ; n4070
g3815 and n3941_not n4070 ; n4071
g3816 and n3949_not n4071_not ; n4072
g3817 and n4069_not n4072 ; n4073
g3818 and n3949_not n4073_not ; n4074
g3819 and b[10] n3938_not ; n4075
g3820 and n3932_not n4075 ; n4076
g3821 and n3940_not n4076_not ; n4077
g3822 and n4074_not n4077 ; n4078
g3823 and n3940_not n4078_not ; n4079
g3824 and b[11] n3929_not ; n4080
g3825 and n3923_not n4080 ; n4081
g3826 and n3931_not n4081_not ; n4082
g3827 and n4079_not n4082 ; n4083
g3828 and n3931_not n4083_not ; n4084
g3829 and b[12] n3920_not ; n4085
g3830 and n3914_not n4085 ; n4086
g3831 and n3922_not n4086_not ; n4087
g3832 and n4084_not n4087 ; n4088
g3833 and n3922_not n4088_not ; n4089
g3834 and b[13] n3911_not ; n4090
g3835 and n3905_not n4090 ; n4091
g3836 and n3913_not n4091_not ; n4092
g3837 and n4089_not n4092 ; n4093
g3838 and n3913_not n4093_not ; n4094
g3839 and b[14] n3902_not ; n4095
g3840 and n3896_not n4095 ; n4096
g3841 and n3904_not n4096_not ; n4097
g3842 and n4094_not n4097 ; n4098
g3843 and n3904_not n4098_not ; n4099
g3844 and b[15] n3893_not ; n4100
g3845 and n3887_not n4100 ; n4101
g3846 and n3895_not n4101_not ; n4102
g3847 and n4099_not n4102 ; n4103
g3848 and n3895_not n4103_not ; n4104
g3849 and b[16] n3884_not ; n4105
g3850 and n3878_not n4105 ; n4106
g3851 and n3886_not n4106_not ; n4107
g3852 and n4104_not n4107 ; n4108
g3853 and n3886_not n4108_not ; n4109
g3854 and b[17] n3875_not ; n4110
g3855 and n3869_not n4110 ; n4111
g3856 and n3877_not n4111_not ; n4112
g3857 and n4109_not n4112 ; n4113
g3858 and n3877_not n4113_not ; n4114
g3859 and b[18] n3866_not ; n4115
g3860 and n3860_not n4115 ; n4116
g3861 and n3868_not n4116_not ; n4117
g3862 and n4114_not n4117 ; n4118
g3863 and n3868_not n4118_not ; n4119
g3864 and b[19] n3857_not ; n4120
g3865 and n3851_not n4120 ; n4121
g3866 and n3859_not n4121_not ; n4122
g3867 and n4119_not n4122 ; n4123
g3868 and n3859_not n4123_not ; n4124
g3869 and b[20] n3848_not ; n4125
g3870 and n3842_not n4125 ; n4126
g3871 and n3850_not n4126_not ; n4127
g3872 and n4124_not n4127 ; n4128
g3873 and n3850_not n4128_not ; n4129
g3874 and b[21] n3831_not ; n4130
g3875 and n3825_not n4130 ; n4131
g3876 and n3841_not n4131_not ; n4132
g3877 and n4129_not n4132 ; n4133
g3878 and n3841_not n4133_not ; n4134
g3879 and b[22] n3833_not ; n4135
g3880 and n3838_not n4135 ; n4136
g3881 and n3840_not n4136_not ; n4137
g3882 and n4134_not n4137 ; n4138
g3883 and n3840_not n4138_not ; n4139
g3884 and n365 n376 ; n4140
g3885 and n588 n4140 ; n4141
g3886 and n598 n4141 ; n4142
g3887 and n595 n4142 ; n4143
g3888 and n4139_not n4143 ; quotient[41]
g3889 and n3832_not quotient[41]_not ; n4145
g3890 and n3850_not n4132 ; n4146
g3891 and n4128_not n4146 ; n4147
g3892 and n4129_not n4132_not ; n4148
g3893 and n4147_not n4148_not ; n4149
g3894 and n4143 n4149_not ; n4150
g3895 and n4139_not n4150 ; n4151
g3896 and n4145_not n4151_not ; n4152
g3897 and b[22]_not n4152_not ; n4153
g3898 and n3849_not quotient[41]_not ; n4154
g3899 and n3859_not n4127 ; n4155
g3900 and n4123_not n4155 ; n4156
g3901 and n4124_not n4127_not ; n4157
g3902 and n4156_not n4157_not ; n4158
g3903 and n4143 n4158_not ; n4159
g3904 and n4139_not n4159 ; n4160
g3905 and n4154_not n4160_not ; n4161
g3906 and b[21]_not n4161_not ; n4162
g3907 and n3858_not quotient[41]_not ; n4163
g3908 and n3868_not n4122 ; n4164
g3909 and n4118_not n4164 ; n4165
g3910 and n4119_not n4122_not ; n4166
g3911 and n4165_not n4166_not ; n4167
g3912 and n4143 n4167_not ; n4168
g3913 and n4139_not n4168 ; n4169
g3914 and n4163_not n4169_not ; n4170
g3915 and b[20]_not n4170_not ; n4171
g3916 and n3867_not quotient[41]_not ; n4172
g3917 and n3877_not n4117 ; n4173
g3918 and n4113_not n4173 ; n4174
g3919 and n4114_not n4117_not ; n4175
g3920 and n4174_not n4175_not ; n4176
g3921 and n4143 n4176_not ; n4177
g3922 and n4139_not n4177 ; n4178
g3923 and n4172_not n4178_not ; n4179
g3924 and b[19]_not n4179_not ; n4180
g3925 and n3876_not quotient[41]_not ; n4181
g3926 and n3886_not n4112 ; n4182
g3927 and n4108_not n4182 ; n4183
g3928 and n4109_not n4112_not ; n4184
g3929 and n4183_not n4184_not ; n4185
g3930 and n4143 n4185_not ; n4186
g3931 and n4139_not n4186 ; n4187
g3932 and n4181_not n4187_not ; n4188
g3933 and b[18]_not n4188_not ; n4189
g3934 and n3885_not quotient[41]_not ; n4190
g3935 and n3895_not n4107 ; n4191
g3936 and n4103_not n4191 ; n4192
g3937 and n4104_not n4107_not ; n4193
g3938 and n4192_not n4193_not ; n4194
g3939 and n4143 n4194_not ; n4195
g3940 and n4139_not n4195 ; n4196
g3941 and n4190_not n4196_not ; n4197
g3942 and b[17]_not n4197_not ; n4198
g3943 and n3894_not quotient[41]_not ; n4199
g3944 and n3904_not n4102 ; n4200
g3945 and n4098_not n4200 ; n4201
g3946 and n4099_not n4102_not ; n4202
g3947 and n4201_not n4202_not ; n4203
g3948 and n4143 n4203_not ; n4204
g3949 and n4139_not n4204 ; n4205
g3950 and n4199_not n4205_not ; n4206
g3951 and b[16]_not n4206_not ; n4207
g3952 and n3903_not quotient[41]_not ; n4208
g3953 and n3913_not n4097 ; n4209
g3954 and n4093_not n4209 ; n4210
g3955 and n4094_not n4097_not ; n4211
g3956 and n4210_not n4211_not ; n4212
g3957 and n4143 n4212_not ; n4213
g3958 and n4139_not n4213 ; n4214
g3959 and n4208_not n4214_not ; n4215
g3960 and b[15]_not n4215_not ; n4216
g3961 and n3912_not quotient[41]_not ; n4217
g3962 and n3922_not n4092 ; n4218
g3963 and n4088_not n4218 ; n4219
g3964 and n4089_not n4092_not ; n4220
g3965 and n4219_not n4220_not ; n4221
g3966 and n4143 n4221_not ; n4222
g3967 and n4139_not n4222 ; n4223
g3968 and n4217_not n4223_not ; n4224
g3969 and b[14]_not n4224_not ; n4225
g3970 and n3921_not quotient[41]_not ; n4226
g3971 and n3931_not n4087 ; n4227
g3972 and n4083_not n4227 ; n4228
g3973 and n4084_not n4087_not ; n4229
g3974 and n4228_not n4229_not ; n4230
g3975 and n4143 n4230_not ; n4231
g3976 and n4139_not n4231 ; n4232
g3977 and n4226_not n4232_not ; n4233
g3978 and b[13]_not n4233_not ; n4234
g3979 and n3930_not quotient[41]_not ; n4235
g3980 and n3940_not n4082 ; n4236
g3981 and n4078_not n4236 ; n4237
g3982 and n4079_not n4082_not ; n4238
g3983 and n4237_not n4238_not ; n4239
g3984 and n4143 n4239_not ; n4240
g3985 and n4139_not n4240 ; n4241
g3986 and n4235_not n4241_not ; n4242
g3987 and b[12]_not n4242_not ; n4243
g3988 and n3939_not quotient[41]_not ; n4244
g3989 and n3949_not n4077 ; n4245
g3990 and n4073_not n4245 ; n4246
g3991 and n4074_not n4077_not ; n4247
g3992 and n4246_not n4247_not ; n4248
g3993 and n4143 n4248_not ; n4249
g3994 and n4139_not n4249 ; n4250
g3995 and n4244_not n4250_not ; n4251
g3996 and b[11]_not n4251_not ; n4252
g3997 and n3948_not quotient[41]_not ; n4253
g3998 and n3958_not n4072 ; n4254
g3999 and n4068_not n4254 ; n4255
g4000 and n4069_not n4072_not ; n4256
g4001 and n4255_not n4256_not ; n4257
g4002 and n4143 n4257_not ; n4258
g4003 and n4139_not n4258 ; n4259
g4004 and n4253_not n4259_not ; n4260
g4005 and b[10]_not n4260_not ; n4261
g4006 and n3957_not quotient[41]_not ; n4262
g4007 and n3967_not n4067 ; n4263
g4008 and n4063_not n4263 ; n4264
g4009 and n4064_not n4067_not ; n4265
g4010 and n4264_not n4265_not ; n4266
g4011 and n4143 n4266_not ; n4267
g4012 and n4139_not n4267 ; n4268
g4013 and n4262_not n4268_not ; n4269
g4014 and b[9]_not n4269_not ; n4270
g4015 and n3966_not quotient[41]_not ; n4271
g4016 and n3976_not n4062 ; n4272
g4017 and n4058_not n4272 ; n4273
g4018 and n4059_not n4062_not ; n4274
g4019 and n4273_not n4274_not ; n4275
g4020 and n4143 n4275_not ; n4276
g4021 and n4139_not n4276 ; n4277
g4022 and n4271_not n4277_not ; n4278
g4023 and b[8]_not n4278_not ; n4279
g4024 and n3975_not quotient[41]_not ; n4280
g4025 and n3985_not n4057 ; n4281
g4026 and n4053_not n4281 ; n4282
g4027 and n4054_not n4057_not ; n4283
g4028 and n4282_not n4283_not ; n4284
g4029 and n4143 n4284_not ; n4285
g4030 and n4139_not n4285 ; n4286
g4031 and n4280_not n4286_not ; n4287
g4032 and b[7]_not n4287_not ; n4288
g4033 and n3984_not quotient[41]_not ; n4289
g4034 and n3994_not n4052 ; n4290
g4035 and n4048_not n4290 ; n4291
g4036 and n4049_not n4052_not ; n4292
g4037 and n4291_not n4292_not ; n4293
g4038 and n4143 n4293_not ; n4294
g4039 and n4139_not n4294 ; n4295
g4040 and n4289_not n4295_not ; n4296
g4041 and b[6]_not n4296_not ; n4297
g4042 and n3993_not quotient[41]_not ; n4298
g4043 and n4003_not n4047 ; n4299
g4044 and n4043_not n4299 ; n4300
g4045 and n4044_not n4047_not ; n4301
g4046 and n4300_not n4301_not ; n4302
g4047 and n4143 n4302_not ; n4303
g4048 and n4139_not n4303 ; n4304
g4049 and n4298_not n4304_not ; n4305
g4050 and b[5]_not n4305_not ; n4306
g4051 and n4002_not quotient[41]_not ; n4307
g4052 and n4011_not n4042 ; n4308
g4053 and n4038_not n4308 ; n4309
g4054 and n4039_not n4042_not ; n4310
g4055 and n4309_not n4310_not ; n4311
g4056 and n4143 n4311_not ; n4312
g4057 and n4139_not n4312 ; n4313
g4058 and n4307_not n4313_not ; n4314
g4059 and b[4]_not n4314_not ; n4315
g4060 and n4010_not quotient[41]_not ; n4316
g4061 and n4033_not n4037 ; n4317
g4062 and n4032_not n4317 ; n4318
g4063 and n4034_not n4037_not ; n4319
g4064 and n4318_not n4319_not ; n4320
g4065 and n4143 n4320_not ; n4321
g4066 and n4139_not n4321 ; n4322
g4067 and n4316_not n4322_not ; n4323
g4068 and b[3]_not n4323_not ; n4324
g4069 and n4026_not quotient[41]_not ; n4325
g4070 and n4029_not n4031 ; n4326
g4071 and n4027_not n4326 ; n4327
g4072 and n4143 n4327_not ; n4328
g4073 and n4032_not n4328 ; n4329
g4074 and n4139_not n4329 ; n4330
g4075 and n4325_not n4330_not ; n4331
g4076 and b[2]_not n4331_not ; n4332
g4077 and b[0] b[23]_not ; n4333
g4078 and n306 n4333 ; n4334
g4079 and n317 n4334 ; n4335
g4080 and n303 n4335 ; n4336
g4081 and n288 n4336 ; n4337
g4082 and n4139_not n4337 ; n4338
g4083 and a[41] n4338_not ; n4339
g4084 and n365 n4031 ; n4340
g4085 and n376 n4340 ; n4341
g4086 and n588 n4341 ; n4342
g4087 and n598 n4342 ; n4343
g4088 and n595 n4343 ; n4344
g4089 and n4139_not n4344 ; n4345
g4090 and n4339_not n4345_not ; n4346
g4091 and b[1] n4346_not ; n4347
g4092 and b[1]_not n4345_not ; n4348
g4093 and n4339_not n4348 ; n4349
g4094 and n4347_not n4349_not ; n4350
g4095 and a[40]_not b[0] ; n4351
g4096 and n4350_not n4351_not ; n4352
g4097 and b[1]_not n4346_not ; n4353
g4098 and n4352_not n4353_not ; n4354
g4099 and b[2] n4330_not ; n4355
g4100 and n4325_not n4355 ; n4356
g4101 and n4332_not n4356_not ; n4357
g4102 and n4354_not n4357 ; n4358
g4103 and n4332_not n4358_not ; n4359
g4104 and b[3] n4322_not ; n4360
g4105 and n4316_not n4360 ; n4361
g4106 and n4324_not n4361_not ; n4362
g4107 and n4359_not n4362 ; n4363
g4108 and n4324_not n4363_not ; n4364
g4109 and b[4] n4313_not ; n4365
g4110 and n4307_not n4365 ; n4366
g4111 and n4315_not n4366_not ; n4367
g4112 and n4364_not n4367 ; n4368
g4113 and n4315_not n4368_not ; n4369
g4114 and b[5] n4304_not ; n4370
g4115 and n4298_not n4370 ; n4371
g4116 and n4306_not n4371_not ; n4372
g4117 and n4369_not n4372 ; n4373
g4118 and n4306_not n4373_not ; n4374
g4119 and b[6] n4295_not ; n4375
g4120 and n4289_not n4375 ; n4376
g4121 and n4297_not n4376_not ; n4377
g4122 and n4374_not n4377 ; n4378
g4123 and n4297_not n4378_not ; n4379
g4124 and b[7] n4286_not ; n4380
g4125 and n4280_not n4380 ; n4381
g4126 and n4288_not n4381_not ; n4382
g4127 and n4379_not n4382 ; n4383
g4128 and n4288_not n4383_not ; n4384
g4129 and b[8] n4277_not ; n4385
g4130 and n4271_not n4385 ; n4386
g4131 and n4279_not n4386_not ; n4387
g4132 and n4384_not n4387 ; n4388
g4133 and n4279_not n4388_not ; n4389
g4134 and b[9] n4268_not ; n4390
g4135 and n4262_not n4390 ; n4391
g4136 and n4270_not n4391_not ; n4392
g4137 and n4389_not n4392 ; n4393
g4138 and n4270_not n4393_not ; n4394
g4139 and b[10] n4259_not ; n4395
g4140 and n4253_not n4395 ; n4396
g4141 and n4261_not n4396_not ; n4397
g4142 and n4394_not n4397 ; n4398
g4143 and n4261_not n4398_not ; n4399
g4144 and b[11] n4250_not ; n4400
g4145 and n4244_not n4400 ; n4401
g4146 and n4252_not n4401_not ; n4402
g4147 and n4399_not n4402 ; n4403
g4148 and n4252_not n4403_not ; n4404
g4149 and b[12] n4241_not ; n4405
g4150 and n4235_not n4405 ; n4406
g4151 and n4243_not n4406_not ; n4407
g4152 and n4404_not n4407 ; n4408
g4153 and n4243_not n4408_not ; n4409
g4154 and b[13] n4232_not ; n4410
g4155 and n4226_not n4410 ; n4411
g4156 and n4234_not n4411_not ; n4412
g4157 and n4409_not n4412 ; n4413
g4158 and n4234_not n4413_not ; n4414
g4159 and b[14] n4223_not ; n4415
g4160 and n4217_not n4415 ; n4416
g4161 and n4225_not n4416_not ; n4417
g4162 and n4414_not n4417 ; n4418
g4163 and n4225_not n4418_not ; n4419
g4164 and b[15] n4214_not ; n4420
g4165 and n4208_not n4420 ; n4421
g4166 and n4216_not n4421_not ; n4422
g4167 and n4419_not n4422 ; n4423
g4168 and n4216_not n4423_not ; n4424
g4169 and b[16] n4205_not ; n4425
g4170 and n4199_not n4425 ; n4426
g4171 and n4207_not n4426_not ; n4427
g4172 and n4424_not n4427 ; n4428
g4173 and n4207_not n4428_not ; n4429
g4174 and b[17] n4196_not ; n4430
g4175 and n4190_not n4430 ; n4431
g4176 and n4198_not n4431_not ; n4432
g4177 and n4429_not n4432 ; n4433
g4178 and n4198_not n4433_not ; n4434
g4179 and b[18] n4187_not ; n4435
g4180 and n4181_not n4435 ; n4436
g4181 and n4189_not n4436_not ; n4437
g4182 and n4434_not n4437 ; n4438
g4183 and n4189_not n4438_not ; n4439
g4184 and b[19] n4178_not ; n4440
g4185 and n4172_not n4440 ; n4441
g4186 and n4180_not n4441_not ; n4442
g4187 and n4439_not n4442 ; n4443
g4188 and n4180_not n4443_not ; n4444
g4189 and b[20] n4169_not ; n4445
g4190 and n4163_not n4445 ; n4446
g4191 and n4171_not n4446_not ; n4447
g4192 and n4444_not n4447 ; n4448
g4193 and n4171_not n4448_not ; n4449
g4194 and b[21] n4160_not ; n4450
g4195 and n4154_not n4450 ; n4451
g4196 and n4162_not n4451_not ; n4452
g4197 and n4449_not n4452 ; n4453
g4198 and n4162_not n4453_not ; n4454
g4199 and b[22] n4151_not ; n4455
g4200 and n4145_not n4455 ; n4456
g4201 and n4153_not n4456_not ; n4457
g4202 and n4454_not n4457 ; n4458
g4203 and n4153_not n4458_not ; n4459
g4204 and n3839_not quotient[41]_not ; n4460
g4205 and n3841_not n4137 ; n4461
g4206 and n4133_not n4461 ; n4462
g4207 and n4134_not n4137_not ; n4463
g4208 and n4462_not n4463_not ; n4464
g4209 and quotient[41] n4464_not ; n4465
g4210 and n4460_not n4465_not ; n4466
g4211 and b[23]_not n4466_not ; n4467
g4212 and b[23] n4460_not ; n4468
g4213 and n4465_not n4468 ; n4469
g4214 and n341 n343 ; n4470
g4215 and n338 n4470 ; n4471
g4216 and n4469_not n4471 ; n4472
g4217 and n4467_not n4472 ; n4473
g4218 and n4459_not n4473 ; n4474
g4219 and n4143 n4466_not ; n4475
g4220 and n4474_not n4475_not ; quotient[40]
g4221 and n4162_not n4457 ; n4477
g4222 and n4453_not n4477 ; n4478
g4223 and n4454_not n4457_not ; n4479
g4224 and n4478_not n4479_not ; n4480
g4225 and quotient[40] n4480_not ; n4481
g4226 and n4152_not n4475_not ; n4482
g4227 and n4474_not n4482 ; n4483
g4228 and n4481_not n4483_not ; n4484
g4229 and n4153_not n4469_not ; n4485
g4230 and n4467_not n4485 ; n4486
g4231 and n4458_not n4486 ; n4487
g4232 and n4467_not n4469_not ; n4488
g4233 and n4459_not n4488_not ; n4489
g4234 and n4487_not n4489_not ; n4490
g4235 and quotient[40] n4490_not ; n4491
g4236 and n4466_not n4475_not ; n4492
g4237 and n4474_not n4492 ; n4493
g4238 and n4491_not n4493_not ; n4494
g4239 and b[24]_not n4494_not ; n4495
g4240 and b[23]_not n4484_not ; n4496
g4241 and n4171_not n4452 ; n4497
g4242 and n4448_not n4497 ; n4498
g4243 and n4449_not n4452_not ; n4499
g4244 and n4498_not n4499_not ; n4500
g4245 and quotient[40] n4500_not ; n4501
g4246 and n4161_not n4475_not ; n4502
g4247 and n4474_not n4502 ; n4503
g4248 and n4501_not n4503_not ; n4504
g4249 and b[22]_not n4504_not ; n4505
g4250 and n4180_not n4447 ; n4506
g4251 and n4443_not n4506 ; n4507
g4252 and n4444_not n4447_not ; n4508
g4253 and n4507_not n4508_not ; n4509
g4254 and quotient[40] n4509_not ; n4510
g4255 and n4170_not n4475_not ; n4511
g4256 and n4474_not n4511 ; n4512
g4257 and n4510_not n4512_not ; n4513
g4258 and b[21]_not n4513_not ; n4514
g4259 and n4189_not n4442 ; n4515
g4260 and n4438_not n4515 ; n4516
g4261 and n4439_not n4442_not ; n4517
g4262 and n4516_not n4517_not ; n4518
g4263 and quotient[40] n4518_not ; n4519
g4264 and n4179_not n4475_not ; n4520
g4265 and n4474_not n4520 ; n4521
g4266 and n4519_not n4521_not ; n4522
g4267 and b[20]_not n4522_not ; n4523
g4268 and n4198_not n4437 ; n4524
g4269 and n4433_not n4524 ; n4525
g4270 and n4434_not n4437_not ; n4526
g4271 and n4525_not n4526_not ; n4527
g4272 and quotient[40] n4527_not ; n4528
g4273 and n4188_not n4475_not ; n4529
g4274 and n4474_not n4529 ; n4530
g4275 and n4528_not n4530_not ; n4531
g4276 and b[19]_not n4531_not ; n4532
g4277 and n4207_not n4432 ; n4533
g4278 and n4428_not n4533 ; n4534
g4279 and n4429_not n4432_not ; n4535
g4280 and n4534_not n4535_not ; n4536
g4281 and quotient[40] n4536_not ; n4537
g4282 and n4197_not n4475_not ; n4538
g4283 and n4474_not n4538 ; n4539
g4284 and n4537_not n4539_not ; n4540
g4285 and b[18]_not n4540_not ; n4541
g4286 and n4216_not n4427 ; n4542
g4287 and n4423_not n4542 ; n4543
g4288 and n4424_not n4427_not ; n4544
g4289 and n4543_not n4544_not ; n4545
g4290 and quotient[40] n4545_not ; n4546
g4291 and n4206_not n4475_not ; n4547
g4292 and n4474_not n4547 ; n4548
g4293 and n4546_not n4548_not ; n4549
g4294 and b[17]_not n4549_not ; n4550
g4295 and n4225_not n4422 ; n4551
g4296 and n4418_not n4551 ; n4552
g4297 and n4419_not n4422_not ; n4553
g4298 and n4552_not n4553_not ; n4554
g4299 and quotient[40] n4554_not ; n4555
g4300 and n4215_not n4475_not ; n4556
g4301 and n4474_not n4556 ; n4557
g4302 and n4555_not n4557_not ; n4558
g4303 and b[16]_not n4558_not ; n4559
g4304 and n4234_not n4417 ; n4560
g4305 and n4413_not n4560 ; n4561
g4306 and n4414_not n4417_not ; n4562
g4307 and n4561_not n4562_not ; n4563
g4308 and quotient[40] n4563_not ; n4564
g4309 and n4224_not n4475_not ; n4565
g4310 and n4474_not n4565 ; n4566
g4311 and n4564_not n4566_not ; n4567
g4312 and b[15]_not n4567_not ; n4568
g4313 and n4243_not n4412 ; n4569
g4314 and n4408_not n4569 ; n4570
g4315 and n4409_not n4412_not ; n4571
g4316 and n4570_not n4571_not ; n4572
g4317 and quotient[40] n4572_not ; n4573
g4318 and n4233_not n4475_not ; n4574
g4319 and n4474_not n4574 ; n4575
g4320 and n4573_not n4575_not ; n4576
g4321 and b[14]_not n4576_not ; n4577
g4322 and n4252_not n4407 ; n4578
g4323 and n4403_not n4578 ; n4579
g4324 and n4404_not n4407_not ; n4580
g4325 and n4579_not n4580_not ; n4581
g4326 and quotient[40] n4581_not ; n4582
g4327 and n4242_not n4475_not ; n4583
g4328 and n4474_not n4583 ; n4584
g4329 and n4582_not n4584_not ; n4585
g4330 and b[13]_not n4585_not ; n4586
g4331 and n4261_not n4402 ; n4587
g4332 and n4398_not n4587 ; n4588
g4333 and n4399_not n4402_not ; n4589
g4334 and n4588_not n4589_not ; n4590
g4335 and quotient[40] n4590_not ; n4591
g4336 and n4251_not n4475_not ; n4592
g4337 and n4474_not n4592 ; n4593
g4338 and n4591_not n4593_not ; n4594
g4339 and b[12]_not n4594_not ; n4595
g4340 and n4270_not n4397 ; n4596
g4341 and n4393_not n4596 ; n4597
g4342 and n4394_not n4397_not ; n4598
g4343 and n4597_not n4598_not ; n4599
g4344 and quotient[40] n4599_not ; n4600
g4345 and n4260_not n4475_not ; n4601
g4346 and n4474_not n4601 ; n4602
g4347 and n4600_not n4602_not ; n4603
g4348 and b[11]_not n4603_not ; n4604
g4349 and n4279_not n4392 ; n4605
g4350 and n4388_not n4605 ; n4606
g4351 and n4389_not n4392_not ; n4607
g4352 and n4606_not n4607_not ; n4608
g4353 and quotient[40] n4608_not ; n4609
g4354 and n4269_not n4475_not ; n4610
g4355 and n4474_not n4610 ; n4611
g4356 and n4609_not n4611_not ; n4612
g4357 and b[10]_not n4612_not ; n4613
g4358 and n4288_not n4387 ; n4614
g4359 and n4383_not n4614 ; n4615
g4360 and n4384_not n4387_not ; n4616
g4361 and n4615_not n4616_not ; n4617
g4362 and quotient[40] n4617_not ; n4618
g4363 and n4278_not n4475_not ; n4619
g4364 and n4474_not n4619 ; n4620
g4365 and n4618_not n4620_not ; n4621
g4366 and b[9]_not n4621_not ; n4622
g4367 and n4297_not n4382 ; n4623
g4368 and n4378_not n4623 ; n4624
g4369 and n4379_not n4382_not ; n4625
g4370 and n4624_not n4625_not ; n4626
g4371 and quotient[40] n4626_not ; n4627
g4372 and n4287_not n4475_not ; n4628
g4373 and n4474_not n4628 ; n4629
g4374 and n4627_not n4629_not ; n4630
g4375 and b[8]_not n4630_not ; n4631
g4376 and n4306_not n4377 ; n4632
g4377 and n4373_not n4632 ; n4633
g4378 and n4374_not n4377_not ; n4634
g4379 and n4633_not n4634_not ; n4635
g4380 and quotient[40] n4635_not ; n4636
g4381 and n4296_not n4475_not ; n4637
g4382 and n4474_not n4637 ; n4638
g4383 and n4636_not n4638_not ; n4639
g4384 and b[7]_not n4639_not ; n4640
g4385 and n4315_not n4372 ; n4641
g4386 and n4368_not n4641 ; n4642
g4387 and n4369_not n4372_not ; n4643
g4388 and n4642_not n4643_not ; n4644
g4389 and quotient[40] n4644_not ; n4645
g4390 and n4305_not n4475_not ; n4646
g4391 and n4474_not n4646 ; n4647
g4392 and n4645_not n4647_not ; n4648
g4393 and b[6]_not n4648_not ; n4649
g4394 and n4324_not n4367 ; n4650
g4395 and n4363_not n4650 ; n4651
g4396 and n4364_not n4367_not ; n4652
g4397 and n4651_not n4652_not ; n4653
g4398 and quotient[40] n4653_not ; n4654
g4399 and n4314_not n4475_not ; n4655
g4400 and n4474_not n4655 ; n4656
g4401 and n4654_not n4656_not ; n4657
g4402 and b[5]_not n4657_not ; n4658
g4403 and n4332_not n4362 ; n4659
g4404 and n4358_not n4659 ; n4660
g4405 and n4359_not n4362_not ; n4661
g4406 and n4660_not n4661_not ; n4662
g4407 and quotient[40] n4662_not ; n4663
g4408 and n4323_not n4475_not ; n4664
g4409 and n4474_not n4664 ; n4665
g4410 and n4663_not n4665_not ; n4666
g4411 and b[4]_not n4666_not ; n4667
g4412 and n4353_not n4357 ; n4668
g4413 and n4352_not n4668 ; n4669
g4414 and n4354_not n4357_not ; n4670
g4415 and n4669_not n4670_not ; n4671
g4416 and quotient[40] n4671_not ; n4672
g4417 and n4331_not n4475_not ; n4673
g4418 and n4474_not n4673 ; n4674
g4419 and n4672_not n4674_not ; n4675
g4420 and b[3]_not n4675_not ; n4676
g4421 and n4349_not n4351 ; n4677
g4422 and n4347_not n4677 ; n4678
g4423 and n4352_not n4678_not ; n4679
g4424 and quotient[40] n4679 ; n4680
g4425 and n4346_not n4475_not ; n4681
g4426 and n4474_not n4681 ; n4682
g4427 and n4680_not n4682_not ; n4683
g4428 and b[2]_not n4683_not ; n4684
g4429 and b[0] quotient[40] ; n4685
g4430 and a[40] n4685_not ; n4686
g4431 and n4351 quotient[40] ; n4687
g4432 and n4686_not n4687_not ; n4688
g4433 and b[1] n4688_not ; n4689
g4434 and b[1]_not n4687_not ; n4690
g4435 and n4686_not n4690 ; n4691
g4436 and n4689_not n4691_not ; n4692
g4437 and a[39]_not b[0] ; n4693
g4438 and n4692_not n4693_not ; n4694
g4439 and b[1]_not n4688_not ; n4695
g4440 and n4694_not n4695_not ; n4696
g4441 and b[2] n4682_not ; n4697
g4442 and n4680_not n4697 ; n4698
g4443 and n4684_not n4698_not ; n4699
g4444 and n4696_not n4699 ; n4700
g4445 and n4684_not n4700_not ; n4701
g4446 and b[3] n4674_not ; n4702
g4447 and n4672_not n4702 ; n4703
g4448 and n4676_not n4703_not ; n4704
g4449 and n4701_not n4704 ; n4705
g4450 and n4676_not n4705_not ; n4706
g4451 and b[4] n4665_not ; n4707
g4452 and n4663_not n4707 ; n4708
g4453 and n4667_not n4708_not ; n4709
g4454 and n4706_not n4709 ; n4710
g4455 and n4667_not n4710_not ; n4711
g4456 and b[5] n4656_not ; n4712
g4457 and n4654_not n4712 ; n4713
g4458 and n4658_not n4713_not ; n4714
g4459 and n4711_not n4714 ; n4715
g4460 and n4658_not n4715_not ; n4716
g4461 and b[6] n4647_not ; n4717
g4462 and n4645_not n4717 ; n4718
g4463 and n4649_not n4718_not ; n4719
g4464 and n4716_not n4719 ; n4720
g4465 and n4649_not n4720_not ; n4721
g4466 and b[7] n4638_not ; n4722
g4467 and n4636_not n4722 ; n4723
g4468 and n4640_not n4723_not ; n4724
g4469 and n4721_not n4724 ; n4725
g4470 and n4640_not n4725_not ; n4726
g4471 and b[8] n4629_not ; n4727
g4472 and n4627_not n4727 ; n4728
g4473 and n4631_not n4728_not ; n4729
g4474 and n4726_not n4729 ; n4730
g4475 and n4631_not n4730_not ; n4731
g4476 and b[9] n4620_not ; n4732
g4477 and n4618_not n4732 ; n4733
g4478 and n4622_not n4733_not ; n4734
g4479 and n4731_not n4734 ; n4735
g4480 and n4622_not n4735_not ; n4736
g4481 and b[10] n4611_not ; n4737
g4482 and n4609_not n4737 ; n4738
g4483 and n4613_not n4738_not ; n4739
g4484 and n4736_not n4739 ; n4740
g4485 and n4613_not n4740_not ; n4741
g4486 and b[11] n4602_not ; n4742
g4487 and n4600_not n4742 ; n4743
g4488 and n4604_not n4743_not ; n4744
g4489 and n4741_not n4744 ; n4745
g4490 and n4604_not n4745_not ; n4746
g4491 and b[12] n4593_not ; n4747
g4492 and n4591_not n4747 ; n4748
g4493 and n4595_not n4748_not ; n4749
g4494 and n4746_not n4749 ; n4750
g4495 and n4595_not n4750_not ; n4751
g4496 and b[13] n4584_not ; n4752
g4497 and n4582_not n4752 ; n4753
g4498 and n4586_not n4753_not ; n4754
g4499 and n4751_not n4754 ; n4755
g4500 and n4586_not n4755_not ; n4756
g4501 and b[14] n4575_not ; n4757
g4502 and n4573_not n4757 ; n4758
g4503 and n4577_not n4758_not ; n4759
g4504 and n4756_not n4759 ; n4760
g4505 and n4577_not n4760_not ; n4761
g4506 and b[15] n4566_not ; n4762
g4507 and n4564_not n4762 ; n4763
g4508 and n4568_not n4763_not ; n4764
g4509 and n4761_not n4764 ; n4765
g4510 and n4568_not n4765_not ; n4766
g4511 and b[16] n4557_not ; n4767
g4512 and n4555_not n4767 ; n4768
g4513 and n4559_not n4768_not ; n4769
g4514 and n4766_not n4769 ; n4770
g4515 and n4559_not n4770_not ; n4771
g4516 and b[17] n4548_not ; n4772
g4517 and n4546_not n4772 ; n4773
g4518 and n4550_not n4773_not ; n4774
g4519 and n4771_not n4774 ; n4775
g4520 and n4550_not n4775_not ; n4776
g4521 and b[18] n4539_not ; n4777
g4522 and n4537_not n4777 ; n4778
g4523 and n4541_not n4778_not ; n4779
g4524 and n4776_not n4779 ; n4780
g4525 and n4541_not n4780_not ; n4781
g4526 and b[19] n4530_not ; n4782
g4527 and n4528_not n4782 ; n4783
g4528 and n4532_not n4783_not ; n4784
g4529 and n4781_not n4784 ; n4785
g4530 and n4532_not n4785_not ; n4786
g4531 and b[20] n4521_not ; n4787
g4532 and n4519_not n4787 ; n4788
g4533 and n4523_not n4788_not ; n4789
g4534 and n4786_not n4789 ; n4790
g4535 and n4523_not n4790_not ; n4791
g4536 and b[21] n4512_not ; n4792
g4537 and n4510_not n4792 ; n4793
g4538 and n4514_not n4793_not ; n4794
g4539 and n4791_not n4794 ; n4795
g4540 and n4514_not n4795_not ; n4796
g4541 and b[22] n4503_not ; n4797
g4542 and n4501_not n4797 ; n4798
g4543 and n4505_not n4798_not ; n4799
g4544 and n4796_not n4799 ; n4800
g4545 and n4505_not n4800_not ; n4801
g4546 and b[23] n4483_not ; n4802
g4547 and n4481_not n4802 ; n4803
g4548 and n4496_not n4803_not ; n4804
g4549 and n4801_not n4804 ; n4805
g4550 and n4496_not n4805_not ; n4806
g4551 and b[24] n4493_not ; n4807
g4552 and n4491_not n4807 ; n4808
g4553 and n4495_not n4808_not ; n4809
g4554 and n4806_not n4809 ; n4810
g4555 and n4495_not n4810_not ; n4811
g4556 and n377 n423 ; n4812
g4557 and n408 n4812 ; n4813
g4558 and n4811_not n4813 ; quotient[39]
g4559 and n4484_not quotient[39]_not ; n4815
g4560 and n4505_not n4804 ; n4816
g4561 and n4800_not n4816 ; n4817
g4562 and n4801_not n4804_not ; n4818
g4563 and n4817_not n4818_not ; n4819
g4564 and n4813 n4819_not ; n4820
g4565 and n4811_not n4820 ; n4821
g4566 and n4815_not n4821_not ; n4822
g4567 and n4494_not quotient[39]_not ; n4823
g4568 and n4496_not n4809 ; n4824
g4569 and n4805_not n4824 ; n4825
g4570 and n4806_not n4809_not ; n4826
g4571 and n4825_not n4826_not ; n4827
g4572 and quotient[39] n4827_not ; n4828
g4573 and n4823_not n4828_not ; n4829
g4574 and b[25]_not n4829_not ; n4830
g4575 and b[24]_not n4822_not ; n4831
g4576 and n4504_not quotient[39]_not ; n4832
g4577 and n4514_not n4799 ; n4833
g4578 and n4795_not n4833 ; n4834
g4579 and n4796_not n4799_not ; n4835
g4580 and n4834_not n4835_not ; n4836
g4581 and n4813 n4836_not ; n4837
g4582 and n4811_not n4837 ; n4838
g4583 and n4832_not n4838_not ; n4839
g4584 and b[23]_not n4839_not ; n4840
g4585 and n4513_not quotient[39]_not ; n4841
g4586 and n4523_not n4794 ; n4842
g4587 and n4790_not n4842 ; n4843
g4588 and n4791_not n4794_not ; n4844
g4589 and n4843_not n4844_not ; n4845
g4590 and n4813 n4845_not ; n4846
g4591 and n4811_not n4846 ; n4847
g4592 and n4841_not n4847_not ; n4848
g4593 and b[22]_not n4848_not ; n4849
g4594 and n4522_not quotient[39]_not ; n4850
g4595 and n4532_not n4789 ; n4851
g4596 and n4785_not n4851 ; n4852
g4597 and n4786_not n4789_not ; n4853
g4598 and n4852_not n4853_not ; n4854
g4599 and n4813 n4854_not ; n4855
g4600 and n4811_not n4855 ; n4856
g4601 and n4850_not n4856_not ; n4857
g4602 and b[21]_not n4857_not ; n4858
g4603 and n4531_not quotient[39]_not ; n4859
g4604 and n4541_not n4784 ; n4860
g4605 and n4780_not n4860 ; n4861
g4606 and n4781_not n4784_not ; n4862
g4607 and n4861_not n4862_not ; n4863
g4608 and n4813 n4863_not ; n4864
g4609 and n4811_not n4864 ; n4865
g4610 and n4859_not n4865_not ; n4866
g4611 and b[20]_not n4866_not ; n4867
g4612 and n4540_not quotient[39]_not ; n4868
g4613 and n4550_not n4779 ; n4869
g4614 and n4775_not n4869 ; n4870
g4615 and n4776_not n4779_not ; n4871
g4616 and n4870_not n4871_not ; n4872
g4617 and n4813 n4872_not ; n4873
g4618 and n4811_not n4873 ; n4874
g4619 and n4868_not n4874_not ; n4875
g4620 and b[19]_not n4875_not ; n4876
g4621 and n4549_not quotient[39]_not ; n4877
g4622 and n4559_not n4774 ; n4878
g4623 and n4770_not n4878 ; n4879
g4624 and n4771_not n4774_not ; n4880
g4625 and n4879_not n4880_not ; n4881
g4626 and n4813 n4881_not ; n4882
g4627 and n4811_not n4882 ; n4883
g4628 and n4877_not n4883_not ; n4884
g4629 and b[18]_not n4884_not ; n4885
g4630 and n4558_not quotient[39]_not ; n4886
g4631 and n4568_not n4769 ; n4887
g4632 and n4765_not n4887 ; n4888
g4633 and n4766_not n4769_not ; n4889
g4634 and n4888_not n4889_not ; n4890
g4635 and n4813 n4890_not ; n4891
g4636 and n4811_not n4891 ; n4892
g4637 and n4886_not n4892_not ; n4893
g4638 and b[17]_not n4893_not ; n4894
g4639 and n4567_not quotient[39]_not ; n4895
g4640 and n4577_not n4764 ; n4896
g4641 and n4760_not n4896 ; n4897
g4642 and n4761_not n4764_not ; n4898
g4643 and n4897_not n4898_not ; n4899
g4644 and n4813 n4899_not ; n4900
g4645 and n4811_not n4900 ; n4901
g4646 and n4895_not n4901_not ; n4902
g4647 and b[16]_not n4902_not ; n4903
g4648 and n4576_not quotient[39]_not ; n4904
g4649 and n4586_not n4759 ; n4905
g4650 and n4755_not n4905 ; n4906
g4651 and n4756_not n4759_not ; n4907
g4652 and n4906_not n4907_not ; n4908
g4653 and n4813 n4908_not ; n4909
g4654 and n4811_not n4909 ; n4910
g4655 and n4904_not n4910_not ; n4911
g4656 and b[15]_not n4911_not ; n4912
g4657 and n4585_not quotient[39]_not ; n4913
g4658 and n4595_not n4754 ; n4914
g4659 and n4750_not n4914 ; n4915
g4660 and n4751_not n4754_not ; n4916
g4661 and n4915_not n4916_not ; n4917
g4662 and n4813 n4917_not ; n4918
g4663 and n4811_not n4918 ; n4919
g4664 and n4913_not n4919_not ; n4920
g4665 and b[14]_not n4920_not ; n4921
g4666 and n4594_not quotient[39]_not ; n4922
g4667 and n4604_not n4749 ; n4923
g4668 and n4745_not n4923 ; n4924
g4669 and n4746_not n4749_not ; n4925
g4670 and n4924_not n4925_not ; n4926
g4671 and n4813 n4926_not ; n4927
g4672 and n4811_not n4927 ; n4928
g4673 and n4922_not n4928_not ; n4929
g4674 and b[13]_not n4929_not ; n4930
g4675 and n4603_not quotient[39]_not ; n4931
g4676 and n4613_not n4744 ; n4932
g4677 and n4740_not n4932 ; n4933
g4678 and n4741_not n4744_not ; n4934
g4679 and n4933_not n4934_not ; n4935
g4680 and n4813 n4935_not ; n4936
g4681 and n4811_not n4936 ; n4937
g4682 and n4931_not n4937_not ; n4938
g4683 and b[12]_not n4938_not ; n4939
g4684 and n4612_not quotient[39]_not ; n4940
g4685 and n4622_not n4739 ; n4941
g4686 and n4735_not n4941 ; n4942
g4687 and n4736_not n4739_not ; n4943
g4688 and n4942_not n4943_not ; n4944
g4689 and n4813 n4944_not ; n4945
g4690 and n4811_not n4945 ; n4946
g4691 and n4940_not n4946_not ; n4947
g4692 and b[11]_not n4947_not ; n4948
g4693 and n4621_not quotient[39]_not ; n4949
g4694 and n4631_not n4734 ; n4950
g4695 and n4730_not n4950 ; n4951
g4696 and n4731_not n4734_not ; n4952
g4697 and n4951_not n4952_not ; n4953
g4698 and n4813 n4953_not ; n4954
g4699 and n4811_not n4954 ; n4955
g4700 and n4949_not n4955_not ; n4956
g4701 and b[10]_not n4956_not ; n4957
g4702 and n4630_not quotient[39]_not ; n4958
g4703 and n4640_not n4729 ; n4959
g4704 and n4725_not n4959 ; n4960
g4705 and n4726_not n4729_not ; n4961
g4706 and n4960_not n4961_not ; n4962
g4707 and n4813 n4962_not ; n4963
g4708 and n4811_not n4963 ; n4964
g4709 and n4958_not n4964_not ; n4965
g4710 and b[9]_not n4965_not ; n4966
g4711 and n4639_not quotient[39]_not ; n4967
g4712 and n4649_not n4724 ; n4968
g4713 and n4720_not n4968 ; n4969
g4714 and n4721_not n4724_not ; n4970
g4715 and n4969_not n4970_not ; n4971
g4716 and n4813 n4971_not ; n4972
g4717 and n4811_not n4972 ; n4973
g4718 and n4967_not n4973_not ; n4974
g4719 and b[8]_not n4974_not ; n4975
g4720 and n4648_not quotient[39]_not ; n4976
g4721 and n4658_not n4719 ; n4977
g4722 and n4715_not n4977 ; n4978
g4723 and n4716_not n4719_not ; n4979
g4724 and n4978_not n4979_not ; n4980
g4725 and n4813 n4980_not ; n4981
g4726 and n4811_not n4981 ; n4982
g4727 and n4976_not n4982_not ; n4983
g4728 and b[7]_not n4983_not ; n4984
g4729 and n4657_not quotient[39]_not ; n4985
g4730 and n4667_not n4714 ; n4986
g4731 and n4710_not n4986 ; n4987
g4732 and n4711_not n4714_not ; n4988
g4733 and n4987_not n4988_not ; n4989
g4734 and n4813 n4989_not ; n4990
g4735 and n4811_not n4990 ; n4991
g4736 and n4985_not n4991_not ; n4992
g4737 and b[6]_not n4992_not ; n4993
g4738 and n4666_not quotient[39]_not ; n4994
g4739 and n4676_not n4709 ; n4995
g4740 and n4705_not n4995 ; n4996
g4741 and n4706_not n4709_not ; n4997
g4742 and n4996_not n4997_not ; n4998
g4743 and n4813 n4998_not ; n4999
g4744 and n4811_not n4999 ; n5000
g4745 and n4994_not n5000_not ; n5001
g4746 and b[5]_not n5001_not ; n5002
g4747 and n4675_not quotient[39]_not ; n5003
g4748 and n4684_not n4704 ; n5004
g4749 and n4700_not n5004 ; n5005
g4750 and n4701_not n4704_not ; n5006
g4751 and n5005_not n5006_not ; n5007
g4752 and n4813 n5007_not ; n5008
g4753 and n4811_not n5008 ; n5009
g4754 and n5003_not n5009_not ; n5010
g4755 and b[4]_not n5010_not ; n5011
g4756 and n4683_not quotient[39]_not ; n5012
g4757 and n4695_not n4699 ; n5013
g4758 and n4694_not n5013 ; n5014
g4759 and n4696_not n4699_not ; n5015
g4760 and n5014_not n5015_not ; n5016
g4761 and n4813 n5016_not ; n5017
g4762 and n4811_not n5017 ; n5018
g4763 and n5012_not n5018_not ; n5019
g4764 and b[3]_not n5019_not ; n5020
g4765 and n4688_not quotient[39]_not ; n5021
g4766 and n4691_not n4693 ; n5022
g4767 and n4689_not n5022 ; n5023
g4768 and n4813 n5023_not ; n5024
g4769 and n4694_not n5024 ; n5025
g4770 and n4811_not n5025 ; n5026
g4771 and n5021_not n5026_not ; n5027
g4772 and b[2]_not n5027_not ; n5028
g4773 and b[0] b[25]_not ; n5029
g4774 and n305 n5029 ; n5030
g4775 and n316 n5030 ; n5031
g4776 and n341 n5031 ; n5032
g4777 and n338 n5032 ; n5033
g4778 and n4811_not n5033 ; n5034
g4779 and a[39] n5034_not ; n5035
g4780 and n376 n4693 ; n5036
g4781 and n588 n5036 ; n5037
g4782 and n598 n5037 ; n5038
g4783 and n595 n5038 ; n5039
g4784 and n4811_not n5039 ; n5040
g4785 and n5035_not n5040_not ; n5041
g4786 and b[1] n5041_not ; n5042
g4787 and b[1]_not n5040_not ; n5043
g4788 and n5035_not n5043 ; n5044
g4789 and n5042_not n5044_not ; n5045
g4790 and a[38]_not b[0] ; n5046
g4791 and n5045_not n5046_not ; n5047
g4792 and b[1]_not n5041_not ; n5048
g4793 and n5047_not n5048_not ; n5049
g4794 and b[2] n5026_not ; n5050
g4795 and n5021_not n5050 ; n5051
g4796 and n5028_not n5051_not ; n5052
g4797 and n5049_not n5052 ; n5053
g4798 and n5028_not n5053_not ; n5054
g4799 and b[3] n5018_not ; n5055
g4800 and n5012_not n5055 ; n5056
g4801 and n5020_not n5056_not ; n5057
g4802 and n5054_not n5057 ; n5058
g4803 and n5020_not n5058_not ; n5059
g4804 and b[4] n5009_not ; n5060
g4805 and n5003_not n5060 ; n5061
g4806 and n5011_not n5061_not ; n5062
g4807 and n5059_not n5062 ; n5063
g4808 and n5011_not n5063_not ; n5064
g4809 and b[5] n5000_not ; n5065
g4810 and n4994_not n5065 ; n5066
g4811 and n5002_not n5066_not ; n5067
g4812 and n5064_not n5067 ; n5068
g4813 and n5002_not n5068_not ; n5069
g4814 and b[6] n4991_not ; n5070
g4815 and n4985_not n5070 ; n5071
g4816 and n4993_not n5071_not ; n5072
g4817 and n5069_not n5072 ; n5073
g4818 and n4993_not n5073_not ; n5074
g4819 and b[7] n4982_not ; n5075
g4820 and n4976_not n5075 ; n5076
g4821 and n4984_not n5076_not ; n5077
g4822 and n5074_not n5077 ; n5078
g4823 and n4984_not n5078_not ; n5079
g4824 and b[8] n4973_not ; n5080
g4825 and n4967_not n5080 ; n5081
g4826 and n4975_not n5081_not ; n5082
g4827 and n5079_not n5082 ; n5083
g4828 and n4975_not n5083_not ; n5084
g4829 and b[9] n4964_not ; n5085
g4830 and n4958_not n5085 ; n5086
g4831 and n4966_not n5086_not ; n5087
g4832 and n5084_not n5087 ; n5088
g4833 and n4966_not n5088_not ; n5089
g4834 and b[10] n4955_not ; n5090
g4835 and n4949_not n5090 ; n5091
g4836 and n4957_not n5091_not ; n5092
g4837 and n5089_not n5092 ; n5093
g4838 and n4957_not n5093_not ; n5094
g4839 and b[11] n4946_not ; n5095
g4840 and n4940_not n5095 ; n5096
g4841 and n4948_not n5096_not ; n5097
g4842 and n5094_not n5097 ; n5098
g4843 and n4948_not n5098_not ; n5099
g4844 and b[12] n4937_not ; n5100
g4845 and n4931_not n5100 ; n5101
g4846 and n4939_not n5101_not ; n5102
g4847 and n5099_not n5102 ; n5103
g4848 and n4939_not n5103_not ; n5104
g4849 and b[13] n4928_not ; n5105
g4850 and n4922_not n5105 ; n5106
g4851 and n4930_not n5106_not ; n5107
g4852 and n5104_not n5107 ; n5108
g4853 and n4930_not n5108_not ; n5109
g4854 and b[14] n4919_not ; n5110
g4855 and n4913_not n5110 ; n5111
g4856 and n4921_not n5111_not ; n5112
g4857 and n5109_not n5112 ; n5113
g4858 and n4921_not n5113_not ; n5114
g4859 and b[15] n4910_not ; n5115
g4860 and n4904_not n5115 ; n5116
g4861 and n4912_not n5116_not ; n5117
g4862 and n5114_not n5117 ; n5118
g4863 and n4912_not n5118_not ; n5119
g4864 and b[16] n4901_not ; n5120
g4865 and n4895_not n5120 ; n5121
g4866 and n4903_not n5121_not ; n5122
g4867 and n5119_not n5122 ; n5123
g4868 and n4903_not n5123_not ; n5124
g4869 and b[17] n4892_not ; n5125
g4870 and n4886_not n5125 ; n5126
g4871 and n4894_not n5126_not ; n5127
g4872 and n5124_not n5127 ; n5128
g4873 and n4894_not n5128_not ; n5129
g4874 and b[18] n4883_not ; n5130
g4875 and n4877_not n5130 ; n5131
g4876 and n4885_not n5131_not ; n5132
g4877 and n5129_not n5132 ; n5133
g4878 and n4885_not n5133_not ; n5134
g4879 and b[19] n4874_not ; n5135
g4880 and n4868_not n5135 ; n5136
g4881 and n4876_not n5136_not ; n5137
g4882 and n5134_not n5137 ; n5138
g4883 and n4876_not n5138_not ; n5139
g4884 and b[20] n4865_not ; n5140
g4885 and n4859_not n5140 ; n5141
g4886 and n4867_not n5141_not ; n5142
g4887 and n5139_not n5142 ; n5143
g4888 and n4867_not n5143_not ; n5144
g4889 and b[21] n4856_not ; n5145
g4890 and n4850_not n5145 ; n5146
g4891 and n4858_not n5146_not ; n5147
g4892 and n5144_not n5147 ; n5148
g4893 and n4858_not n5148_not ; n5149
g4894 and b[22] n4847_not ; n5150
g4895 and n4841_not n5150 ; n5151
g4896 and n4849_not n5151_not ; n5152
g4897 and n5149_not n5152 ; n5153
g4898 and n4849_not n5153_not ; n5154
g4899 and b[23] n4838_not ; n5155
g4900 and n4832_not n5155 ; n5156
g4901 and n4840_not n5156_not ; n5157
g4902 and n5154_not n5157 ; n5158
g4903 and n4840_not n5158_not ; n5159
g4904 and b[24] n4821_not ; n5160
g4905 and n4815_not n5160 ; n5161
g4906 and n4831_not n5161_not ; n5162
g4907 and n5159_not n5162 ; n5163
g4908 and n4831_not n5163_not ; n5164
g4909 and b[25] n4823_not ; n5165
g4910 and n4828_not n5165 ; n5166
g4911 and n4830_not n5166_not ; n5167
g4912 and n5164_not n5167 ; n5168
g4913 and n4830_not n5168_not ; n5169
g4914 and n305 n316 ; n5170
g4915 and n341 n5170 ; n5171
g4916 and n338 n5171 ; n5172
g4917 and n5169_not n5172 ; quotient[38]
g4918 and n4822_not quotient[38]_not ; n5174
g4919 and n4840_not n5162 ; n5175
g4920 and n5158_not n5175 ; n5176
g4921 and n5159_not n5162_not ; n5177
g4922 and n5176_not n5177_not ; n5178
g4923 and n5172 n5178_not ; n5179
g4924 and n5169_not n5179 ; n5180
g4925 and n5174_not n5180_not ; n5181
g4926 and b[25]_not n5181_not ; n5182
g4927 and n4839_not quotient[38]_not ; n5183
g4928 and n4849_not n5157 ; n5184
g4929 and n5153_not n5184 ; n5185
g4930 and n5154_not n5157_not ; n5186
g4931 and n5185_not n5186_not ; n5187
g4932 and n5172 n5187_not ; n5188
g4933 and n5169_not n5188 ; n5189
g4934 and n5183_not n5189_not ; n5190
g4935 and b[24]_not n5190_not ; n5191
g4936 and n4848_not quotient[38]_not ; n5192
g4937 and n4858_not n5152 ; n5193
g4938 and n5148_not n5193 ; n5194
g4939 and n5149_not n5152_not ; n5195
g4940 and n5194_not n5195_not ; n5196
g4941 and n5172 n5196_not ; n5197
g4942 and n5169_not n5197 ; n5198
g4943 and n5192_not n5198_not ; n5199
g4944 and b[23]_not n5199_not ; n5200
g4945 and n4857_not quotient[38]_not ; n5201
g4946 and n4867_not n5147 ; n5202
g4947 and n5143_not n5202 ; n5203
g4948 and n5144_not n5147_not ; n5204
g4949 and n5203_not n5204_not ; n5205
g4950 and n5172 n5205_not ; n5206
g4951 and n5169_not n5206 ; n5207
g4952 and n5201_not n5207_not ; n5208
g4953 and b[22]_not n5208_not ; n5209
g4954 and n4866_not quotient[38]_not ; n5210
g4955 and n4876_not n5142 ; n5211
g4956 and n5138_not n5211 ; n5212
g4957 and n5139_not n5142_not ; n5213
g4958 and n5212_not n5213_not ; n5214
g4959 and n5172 n5214_not ; n5215
g4960 and n5169_not n5215 ; n5216
g4961 and n5210_not n5216_not ; n5217
g4962 and b[21]_not n5217_not ; n5218
g4963 and n4875_not quotient[38]_not ; n5219
g4964 and n4885_not n5137 ; n5220
g4965 and n5133_not n5220 ; n5221
g4966 and n5134_not n5137_not ; n5222
g4967 and n5221_not n5222_not ; n5223
g4968 and n5172 n5223_not ; n5224
g4969 and n5169_not n5224 ; n5225
g4970 and n5219_not n5225_not ; n5226
g4971 and b[20]_not n5226_not ; n5227
g4972 and n4884_not quotient[38]_not ; n5228
g4973 and n4894_not n5132 ; n5229
g4974 and n5128_not n5229 ; n5230
g4975 and n5129_not n5132_not ; n5231
g4976 and n5230_not n5231_not ; n5232
g4977 and n5172 n5232_not ; n5233
g4978 and n5169_not n5233 ; n5234
g4979 and n5228_not n5234_not ; n5235
g4980 and b[19]_not n5235_not ; n5236
g4981 and n4893_not quotient[38]_not ; n5237
g4982 and n4903_not n5127 ; n5238
g4983 and n5123_not n5238 ; n5239
g4984 and n5124_not n5127_not ; n5240
g4985 and n5239_not n5240_not ; n5241
g4986 and n5172 n5241_not ; n5242
g4987 and n5169_not n5242 ; n5243
g4988 and n5237_not n5243_not ; n5244
g4989 and b[18]_not n5244_not ; n5245
g4990 and n4902_not quotient[38]_not ; n5246
g4991 and n4912_not n5122 ; n5247
g4992 and n5118_not n5247 ; n5248
g4993 and n5119_not n5122_not ; n5249
g4994 and n5248_not n5249_not ; n5250
g4995 and n5172 n5250_not ; n5251
g4996 and n5169_not n5251 ; n5252
g4997 and n5246_not n5252_not ; n5253
g4998 and b[17]_not n5253_not ; n5254
g4999 and n4911_not quotient[38]_not ; n5255
g5000 and n4921_not n5117 ; n5256
g5001 and n5113_not n5256 ; n5257
g5002 and n5114_not n5117_not ; n5258
g5003 and n5257_not n5258_not ; n5259
g5004 and n5172 n5259_not ; n5260
g5005 and n5169_not n5260 ; n5261
g5006 and n5255_not n5261_not ; n5262
g5007 and b[16]_not n5262_not ; n5263
g5008 and n4920_not quotient[38]_not ; n5264
g5009 and n4930_not n5112 ; n5265
g5010 and n5108_not n5265 ; n5266
g5011 and n5109_not n5112_not ; n5267
g5012 and n5266_not n5267_not ; n5268
g5013 and n5172 n5268_not ; n5269
g5014 and n5169_not n5269 ; n5270
g5015 and n5264_not n5270_not ; n5271
g5016 and b[15]_not n5271_not ; n5272
g5017 and n4929_not quotient[38]_not ; n5273
g5018 and n4939_not n5107 ; n5274
g5019 and n5103_not n5274 ; n5275
g5020 and n5104_not n5107_not ; n5276
g5021 and n5275_not n5276_not ; n5277
g5022 and n5172 n5277_not ; n5278
g5023 and n5169_not n5278 ; n5279
g5024 and n5273_not n5279_not ; n5280
g5025 and b[14]_not n5280_not ; n5281
g5026 and n4938_not quotient[38]_not ; n5282
g5027 and n4948_not n5102 ; n5283
g5028 and n5098_not n5283 ; n5284
g5029 and n5099_not n5102_not ; n5285
g5030 and n5284_not n5285_not ; n5286
g5031 and n5172 n5286_not ; n5287
g5032 and n5169_not n5287 ; n5288
g5033 and n5282_not n5288_not ; n5289
g5034 and b[13]_not n5289_not ; n5290
g5035 and n4947_not quotient[38]_not ; n5291
g5036 and n4957_not n5097 ; n5292
g5037 and n5093_not n5292 ; n5293
g5038 and n5094_not n5097_not ; n5294
g5039 and n5293_not n5294_not ; n5295
g5040 and n5172 n5295_not ; n5296
g5041 and n5169_not n5296 ; n5297
g5042 and n5291_not n5297_not ; n5298
g5043 and b[12]_not n5298_not ; n5299
g5044 and n4956_not quotient[38]_not ; n5300
g5045 and n4966_not n5092 ; n5301
g5046 and n5088_not n5301 ; n5302
g5047 and n5089_not n5092_not ; n5303
g5048 and n5302_not n5303_not ; n5304
g5049 and n5172 n5304_not ; n5305
g5050 and n5169_not n5305 ; n5306
g5051 and n5300_not n5306_not ; n5307
g5052 and b[11]_not n5307_not ; n5308
g5053 and n4965_not quotient[38]_not ; n5309
g5054 and n4975_not n5087 ; n5310
g5055 and n5083_not n5310 ; n5311
g5056 and n5084_not n5087_not ; n5312
g5057 and n5311_not n5312_not ; n5313
g5058 and n5172 n5313_not ; n5314
g5059 and n5169_not n5314 ; n5315
g5060 and n5309_not n5315_not ; n5316
g5061 and b[10]_not n5316_not ; n5317
g5062 and n4974_not quotient[38]_not ; n5318
g5063 and n4984_not n5082 ; n5319
g5064 and n5078_not n5319 ; n5320
g5065 and n5079_not n5082_not ; n5321
g5066 and n5320_not n5321_not ; n5322
g5067 and n5172 n5322_not ; n5323
g5068 and n5169_not n5323 ; n5324
g5069 and n5318_not n5324_not ; n5325
g5070 and b[9]_not n5325_not ; n5326
g5071 and n4983_not quotient[38]_not ; n5327
g5072 and n4993_not n5077 ; n5328
g5073 and n5073_not n5328 ; n5329
g5074 and n5074_not n5077_not ; n5330
g5075 and n5329_not n5330_not ; n5331
g5076 and n5172 n5331_not ; n5332
g5077 and n5169_not n5332 ; n5333
g5078 and n5327_not n5333_not ; n5334
g5079 and b[8]_not n5334_not ; n5335
g5080 and n4992_not quotient[38]_not ; n5336
g5081 and n5002_not n5072 ; n5337
g5082 and n5068_not n5337 ; n5338
g5083 and n5069_not n5072_not ; n5339
g5084 and n5338_not n5339_not ; n5340
g5085 and n5172 n5340_not ; n5341
g5086 and n5169_not n5341 ; n5342
g5087 and n5336_not n5342_not ; n5343
g5088 and b[7]_not n5343_not ; n5344
g5089 and n5001_not quotient[38]_not ; n5345
g5090 and n5011_not n5067 ; n5346
g5091 and n5063_not n5346 ; n5347
g5092 and n5064_not n5067_not ; n5348
g5093 and n5347_not n5348_not ; n5349
g5094 and n5172 n5349_not ; n5350
g5095 and n5169_not n5350 ; n5351
g5096 and n5345_not n5351_not ; n5352
g5097 and b[6]_not n5352_not ; n5353
g5098 and n5010_not quotient[38]_not ; n5354
g5099 and n5020_not n5062 ; n5355
g5100 and n5058_not n5355 ; n5356
g5101 and n5059_not n5062_not ; n5357
g5102 and n5356_not n5357_not ; n5358
g5103 and n5172 n5358_not ; n5359
g5104 and n5169_not n5359 ; n5360
g5105 and n5354_not n5360_not ; n5361
g5106 and b[5]_not n5361_not ; n5362
g5107 and n5019_not quotient[38]_not ; n5363
g5108 and n5028_not n5057 ; n5364
g5109 and n5053_not n5364 ; n5365
g5110 and n5054_not n5057_not ; n5366
g5111 and n5365_not n5366_not ; n5367
g5112 and n5172 n5367_not ; n5368
g5113 and n5169_not n5368 ; n5369
g5114 and n5363_not n5369_not ; n5370
g5115 and b[4]_not n5370_not ; n5371
g5116 and n5027_not quotient[38]_not ; n5372
g5117 and n5048_not n5052 ; n5373
g5118 and n5047_not n5373 ; n5374
g5119 and n5049_not n5052_not ; n5375
g5120 and n5374_not n5375_not ; n5376
g5121 and n5172 n5376_not ; n5377
g5122 and n5169_not n5377 ; n5378
g5123 and n5372_not n5378_not ; n5379
g5124 and b[3]_not n5379_not ; n5380
g5125 and n5041_not quotient[38]_not ; n5381
g5126 and n5044_not n5046 ; n5382
g5127 and n5042_not n5382 ; n5383
g5128 and n5172 n5383_not ; n5384
g5129 and n5047_not n5384 ; n5385
g5130 and n5169_not n5385 ; n5386
g5131 and n5381_not n5386_not ; n5387
g5132 and b[2]_not n5387_not ; n5388
g5133 and b[0] b[26]_not ; n5389
g5134 and n375 n5389 ; n5390
g5135 and n373 n5390 ; n5391
g5136 and n423 n5391 ; n5392
g5137 and n408 n5392 ; n5393
g5138 and n5169_not n5393 ; n5394
g5139 and a[38] n5394_not ; n5395
g5140 and n305 n5046 ; n5396
g5141 and n316 n5396 ; n5397
g5142 and n341 n5397 ; n5398
g5143 and n338 n5398 ; n5399
g5144 and n5169_not n5399 ; n5400
g5145 and n5395_not n5400_not ; n5401
g5146 and b[1] n5401_not ; n5402
g5147 and b[1]_not n5400_not ; n5403
g5148 and n5395_not n5403 ; n5404
g5149 and n5402_not n5404_not ; n5405
g5150 and a[37]_not b[0] ; n5406
g5151 and n5405_not n5406_not ; n5407
g5152 and b[1]_not n5401_not ; n5408
g5153 and n5407_not n5408_not ; n5409
g5154 and b[2] n5386_not ; n5410
g5155 and n5381_not n5410 ; n5411
g5156 and n5388_not n5411_not ; n5412
g5157 and n5409_not n5412 ; n5413
g5158 and n5388_not n5413_not ; n5414
g5159 and b[3] n5378_not ; n5415
g5160 and n5372_not n5415 ; n5416
g5161 and n5380_not n5416_not ; n5417
g5162 and n5414_not n5417 ; n5418
g5163 and n5380_not n5418_not ; n5419
g5164 and b[4] n5369_not ; n5420
g5165 and n5363_not n5420 ; n5421
g5166 and n5371_not n5421_not ; n5422
g5167 and n5419_not n5422 ; n5423
g5168 and n5371_not n5423_not ; n5424
g5169 and b[5] n5360_not ; n5425
g5170 and n5354_not n5425 ; n5426
g5171 and n5362_not n5426_not ; n5427
g5172 and n5424_not n5427 ; n5428
g5173 and n5362_not n5428_not ; n5429
g5174 and b[6] n5351_not ; n5430
g5175 and n5345_not n5430 ; n5431
g5176 and n5353_not n5431_not ; n5432
g5177 and n5429_not n5432 ; n5433
g5178 and n5353_not n5433_not ; n5434
g5179 and b[7] n5342_not ; n5435
g5180 and n5336_not n5435 ; n5436
g5181 and n5344_not n5436_not ; n5437
g5182 and n5434_not n5437 ; n5438
g5183 and n5344_not n5438_not ; n5439
g5184 and b[8] n5333_not ; n5440
g5185 and n5327_not n5440 ; n5441
g5186 and n5335_not n5441_not ; n5442
g5187 and n5439_not n5442 ; n5443
g5188 and n5335_not n5443_not ; n5444
g5189 and b[9] n5324_not ; n5445
g5190 and n5318_not n5445 ; n5446
g5191 and n5326_not n5446_not ; n5447
g5192 and n5444_not n5447 ; n5448
g5193 and n5326_not n5448_not ; n5449
g5194 and b[10] n5315_not ; n5450
g5195 and n5309_not n5450 ; n5451
g5196 and n5317_not n5451_not ; n5452
g5197 and n5449_not n5452 ; n5453
g5198 and n5317_not n5453_not ; n5454
g5199 and b[11] n5306_not ; n5455
g5200 and n5300_not n5455 ; n5456
g5201 and n5308_not n5456_not ; n5457
g5202 and n5454_not n5457 ; n5458
g5203 and n5308_not n5458_not ; n5459
g5204 and b[12] n5297_not ; n5460
g5205 and n5291_not n5460 ; n5461
g5206 and n5299_not n5461_not ; n5462
g5207 and n5459_not n5462 ; n5463
g5208 and n5299_not n5463_not ; n5464
g5209 and b[13] n5288_not ; n5465
g5210 and n5282_not n5465 ; n5466
g5211 and n5290_not n5466_not ; n5467
g5212 and n5464_not n5467 ; n5468
g5213 and n5290_not n5468_not ; n5469
g5214 and b[14] n5279_not ; n5470
g5215 and n5273_not n5470 ; n5471
g5216 and n5281_not n5471_not ; n5472
g5217 and n5469_not n5472 ; n5473
g5218 and n5281_not n5473_not ; n5474
g5219 and b[15] n5270_not ; n5475
g5220 and n5264_not n5475 ; n5476
g5221 and n5272_not n5476_not ; n5477
g5222 and n5474_not n5477 ; n5478
g5223 and n5272_not n5478_not ; n5479
g5224 and b[16] n5261_not ; n5480
g5225 and n5255_not n5480 ; n5481
g5226 and n5263_not n5481_not ; n5482
g5227 and n5479_not n5482 ; n5483
g5228 and n5263_not n5483_not ; n5484
g5229 and b[17] n5252_not ; n5485
g5230 and n5246_not n5485 ; n5486
g5231 and n5254_not n5486_not ; n5487
g5232 and n5484_not n5487 ; n5488
g5233 and n5254_not n5488_not ; n5489
g5234 and b[18] n5243_not ; n5490
g5235 and n5237_not n5490 ; n5491
g5236 and n5245_not n5491_not ; n5492
g5237 and n5489_not n5492 ; n5493
g5238 and n5245_not n5493_not ; n5494
g5239 and b[19] n5234_not ; n5495
g5240 and n5228_not n5495 ; n5496
g5241 and n5236_not n5496_not ; n5497
g5242 and n5494_not n5497 ; n5498
g5243 and n5236_not n5498_not ; n5499
g5244 and b[20] n5225_not ; n5500
g5245 and n5219_not n5500 ; n5501
g5246 and n5227_not n5501_not ; n5502
g5247 and n5499_not n5502 ; n5503
g5248 and n5227_not n5503_not ; n5504
g5249 and b[21] n5216_not ; n5505
g5250 and n5210_not n5505 ; n5506
g5251 and n5218_not n5506_not ; n5507
g5252 and n5504_not n5507 ; n5508
g5253 and n5218_not n5508_not ; n5509
g5254 and b[22] n5207_not ; n5510
g5255 and n5201_not n5510 ; n5511
g5256 and n5209_not n5511_not ; n5512
g5257 and n5509_not n5512 ; n5513
g5258 and n5209_not n5513_not ; n5514
g5259 and b[23] n5198_not ; n5515
g5260 and n5192_not n5515 ; n5516
g5261 and n5200_not n5516_not ; n5517
g5262 and n5514_not n5517 ; n5518
g5263 and n5200_not n5518_not ; n5519
g5264 and b[24] n5189_not ; n5520
g5265 and n5183_not n5520 ; n5521
g5266 and n5191_not n5521_not ; n5522
g5267 and n5519_not n5522 ; n5523
g5268 and n5191_not n5523_not ; n5524
g5269 and b[25] n5180_not ; n5525
g5270 and n5174_not n5525 ; n5526
g5271 and n5182_not n5526_not ; n5527
g5272 and n5524_not n5527 ; n5528
g5273 and n5182_not n5528_not ; n5529
g5274 and n4829_not quotient[38]_not ; n5530
g5275 and n4831_not n5167 ; n5531
g5276 and n5163_not n5531 ; n5532
g5277 and n5164_not n5167_not ; n5533
g5278 and n5532_not n5533_not ; n5534
g5279 and quotient[38] n5534_not ; n5535
g5280 and n5530_not n5535_not ; n5536
g5281 and b[26]_not n5536_not ; n5537
g5282 and b[26] n5530_not ; n5538
g5283 and n5535_not n5538 ; n5539
g5284 and n373 n375 ; n5540
g5285 and n423 n5540 ; n5541
g5286 and n408 n5541 ; n5542
g5287 and n5539_not n5542 ; n5543
g5288 and n5537_not n5543 ; n5544
g5289 and n5529_not n5544 ; n5545
g5290 and n5172 n5536_not ; n5546
g5291 and n5545_not n5546_not ; quotient[37]
g5292 and n5191_not n5527 ; n5548
g5293 and n5523_not n5548 ; n5549
g5294 and n5524_not n5527_not ; n5550
g5295 and n5549_not n5550_not ; n5551
g5296 and quotient[37] n5551_not ; n5552
g5297 and n5181_not n5546_not ; n5553
g5298 and n5545_not n5553 ; n5554
g5299 and n5552_not n5554_not ; n5555
g5300 and n5182_not n5539_not ; n5556
g5301 and n5537_not n5556 ; n5557
g5302 and n5528_not n5557 ; n5558
g5303 and n5537_not n5539_not ; n5559
g5304 and n5529_not n5559_not ; n5560
g5305 and n5558_not n5560_not ; n5561
g5306 and quotient[37] n5561_not ; n5562
g5307 and n5536_not n5546_not ; n5563
g5308 and n5545_not n5563 ; n5564
g5309 and n5562_not n5564_not ; n5565
g5310 and b[27]_not n5565_not ; n5566
g5311 and b[26]_not n5555_not ; n5567
g5312 and n5200_not n5522 ; n5568
g5313 and n5518_not n5568 ; n5569
g5314 and n5519_not n5522_not ; n5570
g5315 and n5569_not n5570_not ; n5571
g5316 and quotient[37] n5571_not ; n5572
g5317 and n5190_not n5546_not ; n5573
g5318 and n5545_not n5573 ; n5574
g5319 and n5572_not n5574_not ; n5575
g5320 and b[25]_not n5575_not ; n5576
g5321 and n5209_not n5517 ; n5577
g5322 and n5513_not n5577 ; n5578
g5323 and n5514_not n5517_not ; n5579
g5324 and n5578_not n5579_not ; n5580
g5325 and quotient[37] n5580_not ; n5581
g5326 and n5199_not n5546_not ; n5582
g5327 and n5545_not n5582 ; n5583
g5328 and n5581_not n5583_not ; n5584
g5329 and b[24]_not n5584_not ; n5585
g5330 and n5218_not n5512 ; n5586
g5331 and n5508_not n5586 ; n5587
g5332 and n5509_not n5512_not ; n5588
g5333 and n5587_not n5588_not ; n5589
g5334 and quotient[37] n5589_not ; n5590
g5335 and n5208_not n5546_not ; n5591
g5336 and n5545_not n5591 ; n5592
g5337 and n5590_not n5592_not ; n5593
g5338 and b[23]_not n5593_not ; n5594
g5339 and n5227_not n5507 ; n5595
g5340 and n5503_not n5595 ; n5596
g5341 and n5504_not n5507_not ; n5597
g5342 and n5596_not n5597_not ; n5598
g5343 and quotient[37] n5598_not ; n5599
g5344 and n5217_not n5546_not ; n5600
g5345 and n5545_not n5600 ; n5601
g5346 and n5599_not n5601_not ; n5602
g5347 and b[22]_not n5602_not ; n5603
g5348 and n5236_not n5502 ; n5604
g5349 and n5498_not n5604 ; n5605
g5350 and n5499_not n5502_not ; n5606
g5351 and n5605_not n5606_not ; n5607
g5352 and quotient[37] n5607_not ; n5608
g5353 and n5226_not n5546_not ; n5609
g5354 and n5545_not n5609 ; n5610
g5355 and n5608_not n5610_not ; n5611
g5356 and b[21]_not n5611_not ; n5612
g5357 and n5245_not n5497 ; n5613
g5358 and n5493_not n5613 ; n5614
g5359 and n5494_not n5497_not ; n5615
g5360 and n5614_not n5615_not ; n5616
g5361 and quotient[37] n5616_not ; n5617
g5362 and n5235_not n5546_not ; n5618
g5363 and n5545_not n5618 ; n5619
g5364 and n5617_not n5619_not ; n5620
g5365 and b[20]_not n5620_not ; n5621
g5366 and n5254_not n5492 ; n5622
g5367 and n5488_not n5622 ; n5623
g5368 and n5489_not n5492_not ; n5624
g5369 and n5623_not n5624_not ; n5625
g5370 and quotient[37] n5625_not ; n5626
g5371 and n5244_not n5546_not ; n5627
g5372 and n5545_not n5627 ; n5628
g5373 and n5626_not n5628_not ; n5629
g5374 and b[19]_not n5629_not ; n5630
g5375 and n5263_not n5487 ; n5631
g5376 and n5483_not n5631 ; n5632
g5377 and n5484_not n5487_not ; n5633
g5378 and n5632_not n5633_not ; n5634
g5379 and quotient[37] n5634_not ; n5635
g5380 and n5253_not n5546_not ; n5636
g5381 and n5545_not n5636 ; n5637
g5382 and n5635_not n5637_not ; n5638
g5383 and b[18]_not n5638_not ; n5639
g5384 and n5272_not n5482 ; n5640
g5385 and n5478_not n5640 ; n5641
g5386 and n5479_not n5482_not ; n5642
g5387 and n5641_not n5642_not ; n5643
g5388 and quotient[37] n5643_not ; n5644
g5389 and n5262_not n5546_not ; n5645
g5390 and n5545_not n5645 ; n5646
g5391 and n5644_not n5646_not ; n5647
g5392 and b[17]_not n5647_not ; n5648
g5393 and n5281_not n5477 ; n5649
g5394 and n5473_not n5649 ; n5650
g5395 and n5474_not n5477_not ; n5651
g5396 and n5650_not n5651_not ; n5652
g5397 and quotient[37] n5652_not ; n5653
g5398 and n5271_not n5546_not ; n5654
g5399 and n5545_not n5654 ; n5655
g5400 and n5653_not n5655_not ; n5656
g5401 and b[16]_not n5656_not ; n5657
g5402 and n5290_not n5472 ; n5658
g5403 and n5468_not n5658 ; n5659
g5404 and n5469_not n5472_not ; n5660
g5405 and n5659_not n5660_not ; n5661
g5406 and quotient[37] n5661_not ; n5662
g5407 and n5280_not n5546_not ; n5663
g5408 and n5545_not n5663 ; n5664
g5409 and n5662_not n5664_not ; n5665
g5410 and b[15]_not n5665_not ; n5666
g5411 and n5299_not n5467 ; n5667
g5412 and n5463_not n5667 ; n5668
g5413 and n5464_not n5467_not ; n5669
g5414 and n5668_not n5669_not ; n5670
g5415 and quotient[37] n5670_not ; n5671
g5416 and n5289_not n5546_not ; n5672
g5417 and n5545_not n5672 ; n5673
g5418 and n5671_not n5673_not ; n5674
g5419 and b[14]_not n5674_not ; n5675
g5420 and n5308_not n5462 ; n5676
g5421 and n5458_not n5676 ; n5677
g5422 and n5459_not n5462_not ; n5678
g5423 and n5677_not n5678_not ; n5679
g5424 and quotient[37] n5679_not ; n5680
g5425 and n5298_not n5546_not ; n5681
g5426 and n5545_not n5681 ; n5682
g5427 and n5680_not n5682_not ; n5683
g5428 and b[13]_not n5683_not ; n5684
g5429 and n5317_not n5457 ; n5685
g5430 and n5453_not n5685 ; n5686
g5431 and n5454_not n5457_not ; n5687
g5432 and n5686_not n5687_not ; n5688
g5433 and quotient[37] n5688_not ; n5689
g5434 and n5307_not n5546_not ; n5690
g5435 and n5545_not n5690 ; n5691
g5436 and n5689_not n5691_not ; n5692
g5437 and b[12]_not n5692_not ; n5693
g5438 and n5326_not n5452 ; n5694
g5439 and n5448_not n5694 ; n5695
g5440 and n5449_not n5452_not ; n5696
g5441 and n5695_not n5696_not ; n5697
g5442 and quotient[37] n5697_not ; n5698
g5443 and n5316_not n5546_not ; n5699
g5444 and n5545_not n5699 ; n5700
g5445 and n5698_not n5700_not ; n5701
g5446 and b[11]_not n5701_not ; n5702
g5447 and n5335_not n5447 ; n5703
g5448 and n5443_not n5703 ; n5704
g5449 and n5444_not n5447_not ; n5705
g5450 and n5704_not n5705_not ; n5706
g5451 and quotient[37] n5706_not ; n5707
g5452 and n5325_not n5546_not ; n5708
g5453 and n5545_not n5708 ; n5709
g5454 and n5707_not n5709_not ; n5710
g5455 and b[10]_not n5710_not ; n5711
g5456 and n5344_not n5442 ; n5712
g5457 and n5438_not n5712 ; n5713
g5458 and n5439_not n5442_not ; n5714
g5459 and n5713_not n5714_not ; n5715
g5460 and quotient[37] n5715_not ; n5716
g5461 and n5334_not n5546_not ; n5717
g5462 and n5545_not n5717 ; n5718
g5463 and n5716_not n5718_not ; n5719
g5464 and b[9]_not n5719_not ; n5720
g5465 and n5353_not n5437 ; n5721
g5466 and n5433_not n5721 ; n5722
g5467 and n5434_not n5437_not ; n5723
g5468 and n5722_not n5723_not ; n5724
g5469 and quotient[37] n5724_not ; n5725
g5470 and n5343_not n5546_not ; n5726
g5471 and n5545_not n5726 ; n5727
g5472 and n5725_not n5727_not ; n5728
g5473 and b[8]_not n5728_not ; n5729
g5474 and n5362_not n5432 ; n5730
g5475 and n5428_not n5730 ; n5731
g5476 and n5429_not n5432_not ; n5732
g5477 and n5731_not n5732_not ; n5733
g5478 and quotient[37] n5733_not ; n5734
g5479 and n5352_not n5546_not ; n5735
g5480 and n5545_not n5735 ; n5736
g5481 and n5734_not n5736_not ; n5737
g5482 and b[7]_not n5737_not ; n5738
g5483 and n5371_not n5427 ; n5739
g5484 and n5423_not n5739 ; n5740
g5485 and n5424_not n5427_not ; n5741
g5486 and n5740_not n5741_not ; n5742
g5487 and quotient[37] n5742_not ; n5743
g5488 and n5361_not n5546_not ; n5744
g5489 and n5545_not n5744 ; n5745
g5490 and n5743_not n5745_not ; n5746
g5491 and b[6]_not n5746_not ; n5747
g5492 and n5380_not n5422 ; n5748
g5493 and n5418_not n5748 ; n5749
g5494 and n5419_not n5422_not ; n5750
g5495 and n5749_not n5750_not ; n5751
g5496 and quotient[37] n5751_not ; n5752
g5497 and n5370_not n5546_not ; n5753
g5498 and n5545_not n5753 ; n5754
g5499 and n5752_not n5754_not ; n5755
g5500 and b[5]_not n5755_not ; n5756
g5501 and n5388_not n5417 ; n5757
g5502 and n5413_not n5757 ; n5758
g5503 and n5414_not n5417_not ; n5759
g5504 and n5758_not n5759_not ; n5760
g5505 and quotient[37] n5760_not ; n5761
g5506 and n5379_not n5546_not ; n5762
g5507 and n5545_not n5762 ; n5763
g5508 and n5761_not n5763_not ; n5764
g5509 and b[4]_not n5764_not ; n5765
g5510 and n5408_not n5412 ; n5766
g5511 and n5407_not n5766 ; n5767
g5512 and n5409_not n5412_not ; n5768
g5513 and n5767_not n5768_not ; n5769
g5514 and quotient[37] n5769_not ; n5770
g5515 and n5387_not n5546_not ; n5771
g5516 and n5545_not n5771 ; n5772
g5517 and n5770_not n5772_not ; n5773
g5518 and b[3]_not n5773_not ; n5774
g5519 and n5404_not n5406 ; n5775
g5520 and n5402_not n5775 ; n5776
g5521 and n5407_not n5776_not ; n5777
g5522 and quotient[37] n5777 ; n5778
g5523 and n5401_not n5546_not ; n5779
g5524 and n5545_not n5779 ; n5780
g5525 and n5778_not n5780_not ; n5781
g5526 and b[2]_not n5781_not ; n5782
g5527 and b[0] quotient[37] ; n5783
g5528 and a[37] n5783_not ; n5784
g5529 and n5406 quotient[37] ; n5785
g5530 and n5784_not n5785_not ; n5786
g5531 and b[1] n5786_not ; n5787
g5532 and b[1]_not n5785_not ; n5788
g5533 and n5784_not n5788 ; n5789
g5534 and n5787_not n5789_not ; n5790
g5535 and a[36]_not b[0] ; n5791
g5536 and n5790_not n5791_not ; n5792
g5537 and b[1]_not n5786_not ; n5793
g5538 and n5792_not n5793_not ; n5794
g5539 and b[2] n5780_not ; n5795
g5540 and n5778_not n5795 ; n5796
g5541 and n5782_not n5796_not ; n5797
g5542 and n5794_not n5797 ; n5798
g5543 and n5782_not n5798_not ; n5799
g5544 and b[3] n5772_not ; n5800
g5545 and n5770_not n5800 ; n5801
g5546 and n5774_not n5801_not ; n5802
g5547 and n5799_not n5802 ; n5803
g5548 and n5774_not n5803_not ; n5804
g5549 and b[4] n5763_not ; n5805
g5550 and n5761_not n5805 ; n5806
g5551 and n5765_not n5806_not ; n5807
g5552 and n5804_not n5807 ; n5808
g5553 and n5765_not n5808_not ; n5809
g5554 and b[5] n5754_not ; n5810
g5555 and n5752_not n5810 ; n5811
g5556 and n5756_not n5811_not ; n5812
g5557 and n5809_not n5812 ; n5813
g5558 and n5756_not n5813_not ; n5814
g5559 and b[6] n5745_not ; n5815
g5560 and n5743_not n5815 ; n5816
g5561 and n5747_not n5816_not ; n5817
g5562 and n5814_not n5817 ; n5818
g5563 and n5747_not n5818_not ; n5819
g5564 and b[7] n5736_not ; n5820
g5565 and n5734_not n5820 ; n5821
g5566 and n5738_not n5821_not ; n5822
g5567 and n5819_not n5822 ; n5823
g5568 and n5738_not n5823_not ; n5824
g5569 and b[8] n5727_not ; n5825
g5570 and n5725_not n5825 ; n5826
g5571 and n5729_not n5826_not ; n5827
g5572 and n5824_not n5827 ; n5828
g5573 and n5729_not n5828_not ; n5829
g5574 and b[9] n5718_not ; n5830
g5575 and n5716_not n5830 ; n5831
g5576 and n5720_not n5831_not ; n5832
g5577 and n5829_not n5832 ; n5833
g5578 and n5720_not n5833_not ; n5834
g5579 and b[10] n5709_not ; n5835
g5580 and n5707_not n5835 ; n5836
g5581 and n5711_not n5836_not ; n5837
g5582 and n5834_not n5837 ; n5838
g5583 and n5711_not n5838_not ; n5839
g5584 and b[11] n5700_not ; n5840
g5585 and n5698_not n5840 ; n5841
g5586 and n5702_not n5841_not ; n5842
g5587 and n5839_not n5842 ; n5843
g5588 and n5702_not n5843_not ; n5844
g5589 and b[12] n5691_not ; n5845
g5590 and n5689_not n5845 ; n5846
g5591 and n5693_not n5846_not ; n5847
g5592 and n5844_not n5847 ; n5848
g5593 and n5693_not n5848_not ; n5849
g5594 and b[13] n5682_not ; n5850
g5595 and n5680_not n5850 ; n5851
g5596 and n5684_not n5851_not ; n5852
g5597 and n5849_not n5852 ; n5853
g5598 and n5684_not n5853_not ; n5854
g5599 and b[14] n5673_not ; n5855
g5600 and n5671_not n5855 ; n5856
g5601 and n5675_not n5856_not ; n5857
g5602 and n5854_not n5857 ; n5858
g5603 and n5675_not n5858_not ; n5859
g5604 and b[15] n5664_not ; n5860
g5605 and n5662_not n5860 ; n5861
g5606 and n5666_not n5861_not ; n5862
g5607 and n5859_not n5862 ; n5863
g5608 and n5666_not n5863_not ; n5864
g5609 and b[16] n5655_not ; n5865
g5610 and n5653_not n5865 ; n5866
g5611 and n5657_not n5866_not ; n5867
g5612 and n5864_not n5867 ; n5868
g5613 and n5657_not n5868_not ; n5869
g5614 and b[17] n5646_not ; n5870
g5615 and n5644_not n5870 ; n5871
g5616 and n5648_not n5871_not ; n5872
g5617 and n5869_not n5872 ; n5873
g5618 and n5648_not n5873_not ; n5874
g5619 and b[18] n5637_not ; n5875
g5620 and n5635_not n5875 ; n5876
g5621 and n5639_not n5876_not ; n5877
g5622 and n5874_not n5877 ; n5878
g5623 and n5639_not n5878_not ; n5879
g5624 and b[19] n5628_not ; n5880
g5625 and n5626_not n5880 ; n5881
g5626 and n5630_not n5881_not ; n5882
g5627 and n5879_not n5882 ; n5883
g5628 and n5630_not n5883_not ; n5884
g5629 and b[20] n5619_not ; n5885
g5630 and n5617_not n5885 ; n5886
g5631 and n5621_not n5886_not ; n5887
g5632 and n5884_not n5887 ; n5888
g5633 and n5621_not n5888_not ; n5889
g5634 and b[21] n5610_not ; n5890
g5635 and n5608_not n5890 ; n5891
g5636 and n5612_not n5891_not ; n5892
g5637 and n5889_not n5892 ; n5893
g5638 and n5612_not n5893_not ; n5894
g5639 and b[22] n5601_not ; n5895
g5640 and n5599_not n5895 ; n5896
g5641 and n5603_not n5896_not ; n5897
g5642 and n5894_not n5897 ; n5898
g5643 and n5603_not n5898_not ; n5899
g5644 and b[23] n5592_not ; n5900
g5645 and n5590_not n5900 ; n5901
g5646 and n5594_not n5901_not ; n5902
g5647 and n5899_not n5902 ; n5903
g5648 and n5594_not n5903_not ; n5904
g5649 and b[24] n5583_not ; n5905
g5650 and n5581_not n5905 ; n5906
g5651 and n5585_not n5906_not ; n5907
g5652 and n5904_not n5907 ; n5908
g5653 and n5585_not n5908_not ; n5909
g5654 and b[25] n5574_not ; n5910
g5655 and n5572_not n5910 ; n5911
g5656 and n5576_not n5911_not ; n5912
g5657 and n5909_not n5912 ; n5913
g5658 and n5576_not n5913_not ; n5914
g5659 and b[26] n5554_not ; n5915
g5660 and n5552_not n5915 ; n5916
g5661 and n5567_not n5916_not ; n5917
g5662 and n5914_not n5917 ; n5918
g5663 and n5567_not n5918_not ; n5919
g5664 and b[27] n5564_not ; n5920
g5665 and n5562_not n5920 ; n5921
g5666 and n5566_not n5921_not ; n5922
g5667 and n5919_not n5922 ; n5923
g5668 and n5566_not n5923_not ; n5924
g5669 and n303 n317 ; n5925
g5670 and n288 n5925 ; n5926
g5671 and n5924_not n5926 ; quotient[36]
g5672 and n5555_not quotient[36]_not ; n5928
g5673 and n5576_not n5917 ; n5929
g5674 and n5913_not n5929 ; n5930
g5675 and n5914_not n5917_not ; n5931
g5676 and n5930_not n5931_not ; n5932
g5677 and n5926 n5932_not ; n5933
g5678 and n5924_not n5933 ; n5934
g5679 and n5928_not n5934_not ; n5935
g5680 and n5565_not quotient[36]_not ; n5936
g5681 and n5567_not n5922 ; n5937
g5682 and n5918_not n5937 ; n5938
g5683 and n5919_not n5922_not ; n5939
g5684 and n5938_not n5939_not ; n5940
g5685 and quotient[36] n5940_not ; n5941
g5686 and n5936_not n5941_not ; n5942
g5687 and b[28]_not n5942_not ; n5943
g5688 and b[27]_not n5935_not ; n5944
g5689 and n5575_not quotient[36]_not ; n5945
g5690 and n5585_not n5912 ; n5946
g5691 and n5908_not n5946 ; n5947
g5692 and n5909_not n5912_not ; n5948
g5693 and n5947_not n5948_not ; n5949
g5694 and n5926 n5949_not ; n5950
g5695 and n5924_not n5950 ; n5951
g5696 and n5945_not n5951_not ; n5952
g5697 and b[26]_not n5952_not ; n5953
g5698 and n5584_not quotient[36]_not ; n5954
g5699 and n5594_not n5907 ; n5955
g5700 and n5903_not n5955 ; n5956
g5701 and n5904_not n5907_not ; n5957
g5702 and n5956_not n5957_not ; n5958
g5703 and n5926 n5958_not ; n5959
g5704 and n5924_not n5959 ; n5960
g5705 and n5954_not n5960_not ; n5961
g5706 and b[25]_not n5961_not ; n5962
g5707 and n5593_not quotient[36]_not ; n5963
g5708 and n5603_not n5902 ; n5964
g5709 and n5898_not n5964 ; n5965
g5710 and n5899_not n5902_not ; n5966
g5711 and n5965_not n5966_not ; n5967
g5712 and n5926 n5967_not ; n5968
g5713 and n5924_not n5968 ; n5969
g5714 and n5963_not n5969_not ; n5970
g5715 and b[24]_not n5970_not ; n5971
g5716 and n5602_not quotient[36]_not ; n5972
g5717 and n5612_not n5897 ; n5973
g5718 and n5893_not n5973 ; n5974
g5719 and n5894_not n5897_not ; n5975
g5720 and n5974_not n5975_not ; n5976
g5721 and n5926 n5976_not ; n5977
g5722 and n5924_not n5977 ; n5978
g5723 and n5972_not n5978_not ; n5979
g5724 and b[23]_not n5979_not ; n5980
g5725 and n5611_not quotient[36]_not ; n5981
g5726 and n5621_not n5892 ; n5982
g5727 and n5888_not n5982 ; n5983
g5728 and n5889_not n5892_not ; n5984
g5729 and n5983_not n5984_not ; n5985
g5730 and n5926 n5985_not ; n5986
g5731 and n5924_not n5986 ; n5987
g5732 and n5981_not n5987_not ; n5988
g5733 and b[22]_not n5988_not ; n5989
g5734 and n5620_not quotient[36]_not ; n5990
g5735 and n5630_not n5887 ; n5991
g5736 and n5883_not n5991 ; n5992
g5737 and n5884_not n5887_not ; n5993
g5738 and n5992_not n5993_not ; n5994
g5739 and n5926 n5994_not ; n5995
g5740 and n5924_not n5995 ; n5996
g5741 and n5990_not n5996_not ; n5997
g5742 and b[21]_not n5997_not ; n5998
g5743 and n5629_not quotient[36]_not ; n5999
g5744 and n5639_not n5882 ; n6000
g5745 and n5878_not n6000 ; n6001
g5746 and n5879_not n5882_not ; n6002
g5747 and n6001_not n6002_not ; n6003
g5748 and n5926 n6003_not ; n6004
g5749 and n5924_not n6004 ; n6005
g5750 and n5999_not n6005_not ; n6006
g5751 and b[20]_not n6006_not ; n6007
g5752 and n5638_not quotient[36]_not ; n6008
g5753 and n5648_not n5877 ; n6009
g5754 and n5873_not n6009 ; n6010
g5755 and n5874_not n5877_not ; n6011
g5756 and n6010_not n6011_not ; n6012
g5757 and n5926 n6012_not ; n6013
g5758 and n5924_not n6013 ; n6014
g5759 and n6008_not n6014_not ; n6015
g5760 and b[19]_not n6015_not ; n6016
g5761 and n5647_not quotient[36]_not ; n6017
g5762 and n5657_not n5872 ; n6018
g5763 and n5868_not n6018 ; n6019
g5764 and n5869_not n5872_not ; n6020
g5765 and n6019_not n6020_not ; n6021
g5766 and n5926 n6021_not ; n6022
g5767 and n5924_not n6022 ; n6023
g5768 and n6017_not n6023_not ; n6024
g5769 and b[18]_not n6024_not ; n6025
g5770 and n5656_not quotient[36]_not ; n6026
g5771 and n5666_not n5867 ; n6027
g5772 and n5863_not n6027 ; n6028
g5773 and n5864_not n5867_not ; n6029
g5774 and n6028_not n6029_not ; n6030
g5775 and n5926 n6030_not ; n6031
g5776 and n5924_not n6031 ; n6032
g5777 and n6026_not n6032_not ; n6033
g5778 and b[17]_not n6033_not ; n6034
g5779 and n5665_not quotient[36]_not ; n6035
g5780 and n5675_not n5862 ; n6036
g5781 and n5858_not n6036 ; n6037
g5782 and n5859_not n5862_not ; n6038
g5783 and n6037_not n6038_not ; n6039
g5784 and n5926 n6039_not ; n6040
g5785 and n5924_not n6040 ; n6041
g5786 and n6035_not n6041_not ; n6042
g5787 and b[16]_not n6042_not ; n6043
g5788 and n5674_not quotient[36]_not ; n6044
g5789 and n5684_not n5857 ; n6045
g5790 and n5853_not n6045 ; n6046
g5791 and n5854_not n5857_not ; n6047
g5792 and n6046_not n6047_not ; n6048
g5793 and n5926 n6048_not ; n6049
g5794 and n5924_not n6049 ; n6050
g5795 and n6044_not n6050_not ; n6051
g5796 and b[15]_not n6051_not ; n6052
g5797 and n5683_not quotient[36]_not ; n6053
g5798 and n5693_not n5852 ; n6054
g5799 and n5848_not n6054 ; n6055
g5800 and n5849_not n5852_not ; n6056
g5801 and n6055_not n6056_not ; n6057
g5802 and n5926 n6057_not ; n6058
g5803 and n5924_not n6058 ; n6059
g5804 and n6053_not n6059_not ; n6060
g5805 and b[14]_not n6060_not ; n6061
g5806 and n5692_not quotient[36]_not ; n6062
g5807 and n5702_not n5847 ; n6063
g5808 and n5843_not n6063 ; n6064
g5809 and n5844_not n5847_not ; n6065
g5810 and n6064_not n6065_not ; n6066
g5811 and n5926 n6066_not ; n6067
g5812 and n5924_not n6067 ; n6068
g5813 and n6062_not n6068_not ; n6069
g5814 and b[13]_not n6069_not ; n6070
g5815 and n5701_not quotient[36]_not ; n6071
g5816 and n5711_not n5842 ; n6072
g5817 and n5838_not n6072 ; n6073
g5818 and n5839_not n5842_not ; n6074
g5819 and n6073_not n6074_not ; n6075
g5820 and n5926 n6075_not ; n6076
g5821 and n5924_not n6076 ; n6077
g5822 and n6071_not n6077_not ; n6078
g5823 and b[12]_not n6078_not ; n6079
g5824 and n5710_not quotient[36]_not ; n6080
g5825 and n5720_not n5837 ; n6081
g5826 and n5833_not n6081 ; n6082
g5827 and n5834_not n5837_not ; n6083
g5828 and n6082_not n6083_not ; n6084
g5829 and n5926 n6084_not ; n6085
g5830 and n5924_not n6085 ; n6086
g5831 and n6080_not n6086_not ; n6087
g5832 and b[11]_not n6087_not ; n6088
g5833 and n5719_not quotient[36]_not ; n6089
g5834 and n5729_not n5832 ; n6090
g5835 and n5828_not n6090 ; n6091
g5836 and n5829_not n5832_not ; n6092
g5837 and n6091_not n6092_not ; n6093
g5838 and n5926 n6093_not ; n6094
g5839 and n5924_not n6094 ; n6095
g5840 and n6089_not n6095_not ; n6096
g5841 and b[10]_not n6096_not ; n6097
g5842 and n5728_not quotient[36]_not ; n6098
g5843 and n5738_not n5827 ; n6099
g5844 and n5823_not n6099 ; n6100
g5845 and n5824_not n5827_not ; n6101
g5846 and n6100_not n6101_not ; n6102
g5847 and n5926 n6102_not ; n6103
g5848 and n5924_not n6103 ; n6104
g5849 and n6098_not n6104_not ; n6105
g5850 and b[9]_not n6105_not ; n6106
g5851 and n5737_not quotient[36]_not ; n6107
g5852 and n5747_not n5822 ; n6108
g5853 and n5818_not n6108 ; n6109
g5854 and n5819_not n5822_not ; n6110
g5855 and n6109_not n6110_not ; n6111
g5856 and n5926 n6111_not ; n6112
g5857 and n5924_not n6112 ; n6113
g5858 and n6107_not n6113_not ; n6114
g5859 and b[8]_not n6114_not ; n6115
g5860 and n5746_not quotient[36]_not ; n6116
g5861 and n5756_not n5817 ; n6117
g5862 and n5813_not n6117 ; n6118
g5863 and n5814_not n5817_not ; n6119
g5864 and n6118_not n6119_not ; n6120
g5865 and n5926 n6120_not ; n6121
g5866 and n5924_not n6121 ; n6122
g5867 and n6116_not n6122_not ; n6123
g5868 and b[7]_not n6123_not ; n6124
g5869 and n5755_not quotient[36]_not ; n6125
g5870 and n5765_not n5812 ; n6126
g5871 and n5808_not n6126 ; n6127
g5872 and n5809_not n5812_not ; n6128
g5873 and n6127_not n6128_not ; n6129
g5874 and n5926 n6129_not ; n6130
g5875 and n5924_not n6130 ; n6131
g5876 and n6125_not n6131_not ; n6132
g5877 and b[6]_not n6132_not ; n6133
g5878 and n5764_not quotient[36]_not ; n6134
g5879 and n5774_not n5807 ; n6135
g5880 and n5803_not n6135 ; n6136
g5881 and n5804_not n5807_not ; n6137
g5882 and n6136_not n6137_not ; n6138
g5883 and n5926 n6138_not ; n6139
g5884 and n5924_not n6139 ; n6140
g5885 and n6134_not n6140_not ; n6141
g5886 and b[5]_not n6141_not ; n6142
g5887 and n5773_not quotient[36]_not ; n6143
g5888 and n5782_not n5802 ; n6144
g5889 and n5798_not n6144 ; n6145
g5890 and n5799_not n5802_not ; n6146
g5891 and n6145_not n6146_not ; n6147
g5892 and n5926 n6147_not ; n6148
g5893 and n5924_not n6148 ; n6149
g5894 and n6143_not n6149_not ; n6150
g5895 and b[4]_not n6150_not ; n6151
g5896 and n5781_not quotient[36]_not ; n6152
g5897 and n5793_not n5797 ; n6153
g5898 and n5792_not n6153 ; n6154
g5899 and n5794_not n5797_not ; n6155
g5900 and n6154_not n6155_not ; n6156
g5901 and n5926 n6156_not ; n6157
g5902 and n5924_not n6157 ; n6158
g5903 and n6152_not n6158_not ; n6159
g5904 and b[3]_not n6159_not ; n6160
g5905 and n5786_not quotient[36]_not ; n6161
g5906 and n5789_not n5791 ; n6162
g5907 and n5787_not n6162 ; n6163
g5908 and n5926 n6163_not ; n6164
g5909 and n5792_not n6164 ; n6165
g5910 and n5924_not n6165 ; n6166
g5911 and n6161_not n6166_not ; n6167
g5912 and b[2]_not n6167_not ; n6168
g5913 and b[0] b[28]_not ; n6169
g5914 and n373 n6169 ; n6170
g5915 and n423 n6170 ; n6171
g5916 and n408 n6171 ; n6172
g5917 and n5924_not n6172 ; n6173
g5918 and a[36] n6173_not ; n6174
g5919 and n316 n5791 ; n6175
g5920 and n341 n6175 ; n6176
g5921 and n338 n6176 ; n6177
g5922 and n5924_not n6177 ; n6178
g5923 and n6174_not n6178_not ; n6179
g5924 and b[1] n6179_not ; n6180
g5925 and b[1]_not n6178_not ; n6181
g5926 and n6174_not n6181 ; n6182
g5927 and n6180_not n6182_not ; n6183
g5928 and a[35]_not b[0] ; n6184
g5929 and n6183_not n6184_not ; n6185
g5930 and b[1]_not n6179_not ; n6186
g5931 and n6185_not n6186_not ; n6187
g5932 and b[2] n6166_not ; n6188
g5933 and n6161_not n6188 ; n6189
g5934 and n6168_not n6189_not ; n6190
g5935 and n6187_not n6190 ; n6191
g5936 and n6168_not n6191_not ; n6192
g5937 and b[3] n6158_not ; n6193
g5938 and n6152_not n6193 ; n6194
g5939 and n6160_not n6194_not ; n6195
g5940 and n6192_not n6195 ; n6196
g5941 and n6160_not n6196_not ; n6197
g5942 and b[4] n6149_not ; n6198
g5943 and n6143_not n6198 ; n6199
g5944 and n6151_not n6199_not ; n6200
g5945 and n6197_not n6200 ; n6201
g5946 and n6151_not n6201_not ; n6202
g5947 and b[5] n6140_not ; n6203
g5948 and n6134_not n6203 ; n6204
g5949 and n6142_not n6204_not ; n6205
g5950 and n6202_not n6205 ; n6206
g5951 and n6142_not n6206_not ; n6207
g5952 and b[6] n6131_not ; n6208
g5953 and n6125_not n6208 ; n6209
g5954 and n6133_not n6209_not ; n6210
g5955 and n6207_not n6210 ; n6211
g5956 and n6133_not n6211_not ; n6212
g5957 and b[7] n6122_not ; n6213
g5958 and n6116_not n6213 ; n6214
g5959 and n6124_not n6214_not ; n6215
g5960 and n6212_not n6215 ; n6216
g5961 and n6124_not n6216_not ; n6217
g5962 and b[8] n6113_not ; n6218
g5963 and n6107_not n6218 ; n6219
g5964 and n6115_not n6219_not ; n6220
g5965 and n6217_not n6220 ; n6221
g5966 and n6115_not n6221_not ; n6222
g5967 and b[9] n6104_not ; n6223
g5968 and n6098_not n6223 ; n6224
g5969 and n6106_not n6224_not ; n6225
g5970 and n6222_not n6225 ; n6226
g5971 and n6106_not n6226_not ; n6227
g5972 and b[10] n6095_not ; n6228
g5973 and n6089_not n6228 ; n6229
g5974 and n6097_not n6229_not ; n6230
g5975 and n6227_not n6230 ; n6231
g5976 and n6097_not n6231_not ; n6232
g5977 and b[11] n6086_not ; n6233
g5978 and n6080_not n6233 ; n6234
g5979 and n6088_not n6234_not ; n6235
g5980 and n6232_not n6235 ; n6236
g5981 and n6088_not n6236_not ; n6237
g5982 and b[12] n6077_not ; n6238
g5983 and n6071_not n6238 ; n6239
g5984 and n6079_not n6239_not ; n6240
g5985 and n6237_not n6240 ; n6241
g5986 and n6079_not n6241_not ; n6242
g5987 and b[13] n6068_not ; n6243
g5988 and n6062_not n6243 ; n6244
g5989 and n6070_not n6244_not ; n6245
g5990 and n6242_not n6245 ; n6246
g5991 and n6070_not n6246_not ; n6247
g5992 and b[14] n6059_not ; n6248
g5993 and n6053_not n6248 ; n6249
g5994 and n6061_not n6249_not ; n6250
g5995 and n6247_not n6250 ; n6251
g5996 and n6061_not n6251_not ; n6252
g5997 and b[15] n6050_not ; n6253
g5998 and n6044_not n6253 ; n6254
g5999 and n6052_not n6254_not ; n6255
g6000 and n6252_not n6255 ; n6256
g6001 and n6052_not n6256_not ; n6257
g6002 and b[16] n6041_not ; n6258
g6003 and n6035_not n6258 ; n6259
g6004 and n6043_not n6259_not ; n6260
g6005 and n6257_not n6260 ; n6261
g6006 and n6043_not n6261_not ; n6262
g6007 and b[17] n6032_not ; n6263
g6008 and n6026_not n6263 ; n6264
g6009 and n6034_not n6264_not ; n6265
g6010 and n6262_not n6265 ; n6266
g6011 and n6034_not n6266_not ; n6267
g6012 and b[18] n6023_not ; n6268
g6013 and n6017_not n6268 ; n6269
g6014 and n6025_not n6269_not ; n6270
g6015 and n6267_not n6270 ; n6271
g6016 and n6025_not n6271_not ; n6272
g6017 and b[19] n6014_not ; n6273
g6018 and n6008_not n6273 ; n6274
g6019 and n6016_not n6274_not ; n6275
g6020 and n6272_not n6275 ; n6276
g6021 and n6016_not n6276_not ; n6277
g6022 and b[20] n6005_not ; n6278
g6023 and n5999_not n6278 ; n6279
g6024 and n6007_not n6279_not ; n6280
g6025 and n6277_not n6280 ; n6281
g6026 and n6007_not n6281_not ; n6282
g6027 and b[21] n5996_not ; n6283
g6028 and n5990_not n6283 ; n6284
g6029 and n5998_not n6284_not ; n6285
g6030 and n6282_not n6285 ; n6286
g6031 and n5998_not n6286_not ; n6287
g6032 and b[22] n5987_not ; n6288
g6033 and n5981_not n6288 ; n6289
g6034 and n5989_not n6289_not ; n6290
g6035 and n6287_not n6290 ; n6291
g6036 and n5989_not n6291_not ; n6292
g6037 and b[23] n5978_not ; n6293
g6038 and n5972_not n6293 ; n6294
g6039 and n5980_not n6294_not ; n6295
g6040 and n6292_not n6295 ; n6296
g6041 and n5980_not n6296_not ; n6297
g6042 and b[24] n5969_not ; n6298
g6043 and n5963_not n6298 ; n6299
g6044 and n5971_not n6299_not ; n6300
g6045 and n6297_not n6300 ; n6301
g6046 and n5971_not n6301_not ; n6302
g6047 and b[25] n5960_not ; n6303
g6048 and n5954_not n6303 ; n6304
g6049 and n5962_not n6304_not ; n6305
g6050 and n6302_not n6305 ; n6306
g6051 and n5962_not n6306_not ; n6307
g6052 and b[26] n5951_not ; n6308
g6053 and n5945_not n6308 ; n6309
g6054 and n5953_not n6309_not ; n6310
g6055 and n6307_not n6310 ; n6311
g6056 and n5953_not n6311_not ; n6312
g6057 and b[27] n5934_not ; n6313
g6058 and n5928_not n6313 ; n6314
g6059 and n5944_not n6314_not ; n6315
g6060 and n6312_not n6315 ; n6316
g6061 and n5944_not n6316_not ; n6317
g6062 and b[28] n5936_not ; n6318
g6063 and n5941_not n6318 ; n6319
g6064 and n5943_not n6319_not ; n6320
g6065 and n6317_not n6320 ; n6321
g6066 and n5943_not n6321_not ; n6322
g6067 and n588 n598 ; n6323
g6068 and n595 n6323 ; n6324
g6069 and n6322_not n6324 ; quotient[35]
g6070 and n5935_not quotient[35]_not ; n6326
g6071 and n5953_not n6315 ; n6327
g6072 and n6311_not n6327 ; n6328
g6073 and n6312_not n6315_not ; n6329
g6074 and n6328_not n6329_not ; n6330
g6075 and n6324 n6330_not ; n6331
g6076 and n6322_not n6331 ; n6332
g6077 and n6326_not n6332_not ; n6333
g6078 and b[28]_not n6333_not ; n6334
g6079 and n5952_not quotient[35]_not ; n6335
g6080 and n5962_not n6310 ; n6336
g6081 and n6306_not n6336 ; n6337
g6082 and n6307_not n6310_not ; n6338
g6083 and n6337_not n6338_not ; n6339
g6084 and n6324 n6339_not ; n6340
g6085 and n6322_not n6340 ; n6341
g6086 and n6335_not n6341_not ; n6342
g6087 and b[27]_not n6342_not ; n6343
g6088 and n5961_not quotient[35]_not ; n6344
g6089 and n5971_not n6305 ; n6345
g6090 and n6301_not n6345 ; n6346
g6091 and n6302_not n6305_not ; n6347
g6092 and n6346_not n6347_not ; n6348
g6093 and n6324 n6348_not ; n6349
g6094 and n6322_not n6349 ; n6350
g6095 and n6344_not n6350_not ; n6351
g6096 and b[26]_not n6351_not ; n6352
g6097 and n5970_not quotient[35]_not ; n6353
g6098 and n5980_not n6300 ; n6354
g6099 and n6296_not n6354 ; n6355
g6100 and n6297_not n6300_not ; n6356
g6101 and n6355_not n6356_not ; n6357
g6102 and n6324 n6357_not ; n6358
g6103 and n6322_not n6358 ; n6359
g6104 and n6353_not n6359_not ; n6360
g6105 and b[25]_not n6360_not ; n6361
g6106 and n5979_not quotient[35]_not ; n6362
g6107 and n5989_not n6295 ; n6363
g6108 and n6291_not n6363 ; n6364
g6109 and n6292_not n6295_not ; n6365
g6110 and n6364_not n6365_not ; n6366
g6111 and n6324 n6366_not ; n6367
g6112 and n6322_not n6367 ; n6368
g6113 and n6362_not n6368_not ; n6369
g6114 and b[24]_not n6369_not ; n6370
g6115 and n5988_not quotient[35]_not ; n6371
g6116 and n5998_not n6290 ; n6372
g6117 and n6286_not n6372 ; n6373
g6118 and n6287_not n6290_not ; n6374
g6119 and n6373_not n6374_not ; n6375
g6120 and n6324 n6375_not ; n6376
g6121 and n6322_not n6376 ; n6377
g6122 and n6371_not n6377_not ; n6378
g6123 and b[23]_not n6378_not ; n6379
g6124 and n5997_not quotient[35]_not ; n6380
g6125 and n6007_not n6285 ; n6381
g6126 and n6281_not n6381 ; n6382
g6127 and n6282_not n6285_not ; n6383
g6128 and n6382_not n6383_not ; n6384
g6129 and n6324 n6384_not ; n6385
g6130 and n6322_not n6385 ; n6386
g6131 and n6380_not n6386_not ; n6387
g6132 and b[22]_not n6387_not ; n6388
g6133 and n6006_not quotient[35]_not ; n6389
g6134 and n6016_not n6280 ; n6390
g6135 and n6276_not n6390 ; n6391
g6136 and n6277_not n6280_not ; n6392
g6137 and n6391_not n6392_not ; n6393
g6138 and n6324 n6393_not ; n6394
g6139 and n6322_not n6394 ; n6395
g6140 and n6389_not n6395_not ; n6396
g6141 and b[21]_not n6396_not ; n6397
g6142 and n6015_not quotient[35]_not ; n6398
g6143 and n6025_not n6275 ; n6399
g6144 and n6271_not n6399 ; n6400
g6145 and n6272_not n6275_not ; n6401
g6146 and n6400_not n6401_not ; n6402
g6147 and n6324 n6402_not ; n6403
g6148 and n6322_not n6403 ; n6404
g6149 and n6398_not n6404_not ; n6405
g6150 and b[20]_not n6405_not ; n6406
g6151 and n6024_not quotient[35]_not ; n6407
g6152 and n6034_not n6270 ; n6408
g6153 and n6266_not n6408 ; n6409
g6154 and n6267_not n6270_not ; n6410
g6155 and n6409_not n6410_not ; n6411
g6156 and n6324 n6411_not ; n6412
g6157 and n6322_not n6412 ; n6413
g6158 and n6407_not n6413_not ; n6414
g6159 and b[19]_not n6414_not ; n6415
g6160 and n6033_not quotient[35]_not ; n6416
g6161 and n6043_not n6265 ; n6417
g6162 and n6261_not n6417 ; n6418
g6163 and n6262_not n6265_not ; n6419
g6164 and n6418_not n6419_not ; n6420
g6165 and n6324 n6420_not ; n6421
g6166 and n6322_not n6421 ; n6422
g6167 and n6416_not n6422_not ; n6423
g6168 and b[18]_not n6423_not ; n6424
g6169 and n6042_not quotient[35]_not ; n6425
g6170 and n6052_not n6260 ; n6426
g6171 and n6256_not n6426 ; n6427
g6172 and n6257_not n6260_not ; n6428
g6173 and n6427_not n6428_not ; n6429
g6174 and n6324 n6429_not ; n6430
g6175 and n6322_not n6430 ; n6431
g6176 and n6425_not n6431_not ; n6432
g6177 and b[17]_not n6432_not ; n6433
g6178 and n6051_not quotient[35]_not ; n6434
g6179 and n6061_not n6255 ; n6435
g6180 and n6251_not n6435 ; n6436
g6181 and n6252_not n6255_not ; n6437
g6182 and n6436_not n6437_not ; n6438
g6183 and n6324 n6438_not ; n6439
g6184 and n6322_not n6439 ; n6440
g6185 and n6434_not n6440_not ; n6441
g6186 and b[16]_not n6441_not ; n6442
g6187 and n6060_not quotient[35]_not ; n6443
g6188 and n6070_not n6250 ; n6444
g6189 and n6246_not n6444 ; n6445
g6190 and n6247_not n6250_not ; n6446
g6191 and n6445_not n6446_not ; n6447
g6192 and n6324 n6447_not ; n6448
g6193 and n6322_not n6448 ; n6449
g6194 and n6443_not n6449_not ; n6450
g6195 and b[15]_not n6450_not ; n6451
g6196 and n6069_not quotient[35]_not ; n6452
g6197 and n6079_not n6245 ; n6453
g6198 and n6241_not n6453 ; n6454
g6199 and n6242_not n6245_not ; n6455
g6200 and n6454_not n6455_not ; n6456
g6201 and n6324 n6456_not ; n6457
g6202 and n6322_not n6457 ; n6458
g6203 and n6452_not n6458_not ; n6459
g6204 and b[14]_not n6459_not ; n6460
g6205 and n6078_not quotient[35]_not ; n6461
g6206 and n6088_not n6240 ; n6462
g6207 and n6236_not n6462 ; n6463
g6208 and n6237_not n6240_not ; n6464
g6209 and n6463_not n6464_not ; n6465
g6210 and n6324 n6465_not ; n6466
g6211 and n6322_not n6466 ; n6467
g6212 and n6461_not n6467_not ; n6468
g6213 and b[13]_not n6468_not ; n6469
g6214 and n6087_not quotient[35]_not ; n6470
g6215 and n6097_not n6235 ; n6471
g6216 and n6231_not n6471 ; n6472
g6217 and n6232_not n6235_not ; n6473
g6218 and n6472_not n6473_not ; n6474
g6219 and n6324 n6474_not ; n6475
g6220 and n6322_not n6475 ; n6476
g6221 and n6470_not n6476_not ; n6477
g6222 and b[12]_not n6477_not ; n6478
g6223 and n6096_not quotient[35]_not ; n6479
g6224 and n6106_not n6230 ; n6480
g6225 and n6226_not n6480 ; n6481
g6226 and n6227_not n6230_not ; n6482
g6227 and n6481_not n6482_not ; n6483
g6228 and n6324 n6483_not ; n6484
g6229 and n6322_not n6484 ; n6485
g6230 and n6479_not n6485_not ; n6486
g6231 and b[11]_not n6486_not ; n6487
g6232 and n6105_not quotient[35]_not ; n6488
g6233 and n6115_not n6225 ; n6489
g6234 and n6221_not n6489 ; n6490
g6235 and n6222_not n6225_not ; n6491
g6236 and n6490_not n6491_not ; n6492
g6237 and n6324 n6492_not ; n6493
g6238 and n6322_not n6493 ; n6494
g6239 and n6488_not n6494_not ; n6495
g6240 and b[10]_not n6495_not ; n6496
g6241 and n6114_not quotient[35]_not ; n6497
g6242 and n6124_not n6220 ; n6498
g6243 and n6216_not n6498 ; n6499
g6244 and n6217_not n6220_not ; n6500
g6245 and n6499_not n6500_not ; n6501
g6246 and n6324 n6501_not ; n6502
g6247 and n6322_not n6502 ; n6503
g6248 and n6497_not n6503_not ; n6504
g6249 and b[9]_not n6504_not ; n6505
g6250 and n6123_not quotient[35]_not ; n6506
g6251 and n6133_not n6215 ; n6507
g6252 and n6211_not n6507 ; n6508
g6253 and n6212_not n6215_not ; n6509
g6254 and n6508_not n6509_not ; n6510
g6255 and n6324 n6510_not ; n6511
g6256 and n6322_not n6511 ; n6512
g6257 and n6506_not n6512_not ; n6513
g6258 and b[8]_not n6513_not ; n6514
g6259 and n6132_not quotient[35]_not ; n6515
g6260 and n6142_not n6210 ; n6516
g6261 and n6206_not n6516 ; n6517
g6262 and n6207_not n6210_not ; n6518
g6263 and n6517_not n6518_not ; n6519
g6264 and n6324 n6519_not ; n6520
g6265 and n6322_not n6520 ; n6521
g6266 and n6515_not n6521_not ; n6522
g6267 and b[7]_not n6522_not ; n6523
g6268 and n6141_not quotient[35]_not ; n6524
g6269 and n6151_not n6205 ; n6525
g6270 and n6201_not n6525 ; n6526
g6271 and n6202_not n6205_not ; n6527
g6272 and n6526_not n6527_not ; n6528
g6273 and n6324 n6528_not ; n6529
g6274 and n6322_not n6529 ; n6530
g6275 and n6524_not n6530_not ; n6531
g6276 and b[6]_not n6531_not ; n6532
g6277 and n6150_not quotient[35]_not ; n6533
g6278 and n6160_not n6200 ; n6534
g6279 and n6196_not n6534 ; n6535
g6280 and n6197_not n6200_not ; n6536
g6281 and n6535_not n6536_not ; n6537
g6282 and n6324 n6537_not ; n6538
g6283 and n6322_not n6538 ; n6539
g6284 and n6533_not n6539_not ; n6540
g6285 and b[5]_not n6540_not ; n6541
g6286 and n6159_not quotient[35]_not ; n6542
g6287 and n6168_not n6195 ; n6543
g6288 and n6191_not n6543 ; n6544
g6289 and n6192_not n6195_not ; n6545
g6290 and n6544_not n6545_not ; n6546
g6291 and n6324 n6546_not ; n6547
g6292 and n6322_not n6547 ; n6548
g6293 and n6542_not n6548_not ; n6549
g6294 and b[4]_not n6549_not ; n6550
g6295 and n6167_not quotient[35]_not ; n6551
g6296 and n6186_not n6190 ; n6552
g6297 and n6185_not n6552 ; n6553
g6298 and n6187_not n6190_not ; n6554
g6299 and n6553_not n6554_not ; n6555
g6300 and n6324 n6555_not ; n6556
g6301 and n6322_not n6556 ; n6557
g6302 and n6551_not n6557_not ; n6558
g6303 and b[3]_not n6558_not ; n6559
g6304 and n6179_not quotient[35]_not ; n6560
g6305 and n6182_not n6184 ; n6561
g6306 and n6180_not n6561 ; n6562
g6307 and n6324 n6562_not ; n6563
g6308 and n6185_not n6563 ; n6564
g6309 and n6322_not n6564 ; n6565
g6310 and n6560_not n6565_not ; n6566
g6311 and b[2]_not n6566_not ; n6567
g6312 and b[0] b[29]_not ; n6568
g6313 and n315 n6568 ; n6569
g6314 and n313 n6569 ; n6570
g6315 and n303 n6570 ; n6571
g6316 and n288 n6571 ; n6572
g6317 and n6322_not n6572 ; n6573
g6318 and a[35] n6573_not ; n6574
g6319 and n373 n6184 ; n6575
g6320 and n423 n6575 ; n6576
g6321 and n408 n6576 ; n6577
g6322 and n6322_not n6577 ; n6578
g6323 and n6574_not n6578_not ; n6579
g6324 and b[1] n6579_not ; n6580
g6325 and b[1]_not n6578_not ; n6581
g6326 and n6574_not n6581 ; n6582
g6327 and n6580_not n6582_not ; n6583
g6328 and a[34]_not b[0] ; n6584
g6329 and n6583_not n6584_not ; n6585
g6330 and b[1]_not n6579_not ; n6586
g6331 and n6585_not n6586_not ; n6587
g6332 and b[2] n6565_not ; n6588
g6333 and n6560_not n6588 ; n6589
g6334 and n6567_not n6589_not ; n6590
g6335 and n6587_not n6590 ; n6591
g6336 and n6567_not n6591_not ; n6592
g6337 and b[3] n6557_not ; n6593
g6338 and n6551_not n6593 ; n6594
g6339 and n6559_not n6594_not ; n6595
g6340 and n6592_not n6595 ; n6596
g6341 and n6559_not n6596_not ; n6597
g6342 and b[4] n6548_not ; n6598
g6343 and n6542_not n6598 ; n6599
g6344 and n6550_not n6599_not ; n6600
g6345 and n6597_not n6600 ; n6601
g6346 and n6550_not n6601_not ; n6602
g6347 and b[5] n6539_not ; n6603
g6348 and n6533_not n6603 ; n6604
g6349 and n6541_not n6604_not ; n6605
g6350 and n6602_not n6605 ; n6606
g6351 and n6541_not n6606_not ; n6607
g6352 and b[6] n6530_not ; n6608
g6353 and n6524_not n6608 ; n6609
g6354 and n6532_not n6609_not ; n6610
g6355 and n6607_not n6610 ; n6611
g6356 and n6532_not n6611_not ; n6612
g6357 and b[7] n6521_not ; n6613
g6358 and n6515_not n6613 ; n6614
g6359 and n6523_not n6614_not ; n6615
g6360 and n6612_not n6615 ; n6616
g6361 and n6523_not n6616_not ; n6617
g6362 and b[8] n6512_not ; n6618
g6363 and n6506_not n6618 ; n6619
g6364 and n6514_not n6619_not ; n6620
g6365 and n6617_not n6620 ; n6621
g6366 and n6514_not n6621_not ; n6622
g6367 and b[9] n6503_not ; n6623
g6368 and n6497_not n6623 ; n6624
g6369 and n6505_not n6624_not ; n6625
g6370 and n6622_not n6625 ; n6626
g6371 and n6505_not n6626_not ; n6627
g6372 and b[10] n6494_not ; n6628
g6373 and n6488_not n6628 ; n6629
g6374 and n6496_not n6629_not ; n6630
g6375 and n6627_not n6630 ; n6631
g6376 and n6496_not n6631_not ; n6632
g6377 and b[11] n6485_not ; n6633
g6378 and n6479_not n6633 ; n6634
g6379 and n6487_not n6634_not ; n6635
g6380 and n6632_not n6635 ; n6636
g6381 and n6487_not n6636_not ; n6637
g6382 and b[12] n6476_not ; n6638
g6383 and n6470_not n6638 ; n6639
g6384 and n6478_not n6639_not ; n6640
g6385 and n6637_not n6640 ; n6641
g6386 and n6478_not n6641_not ; n6642
g6387 and b[13] n6467_not ; n6643
g6388 and n6461_not n6643 ; n6644
g6389 and n6469_not n6644_not ; n6645
g6390 and n6642_not n6645 ; n6646
g6391 and n6469_not n6646_not ; n6647
g6392 and b[14] n6458_not ; n6648
g6393 and n6452_not n6648 ; n6649
g6394 and n6460_not n6649_not ; n6650
g6395 and n6647_not n6650 ; n6651
g6396 and n6460_not n6651_not ; n6652
g6397 and b[15] n6449_not ; n6653
g6398 and n6443_not n6653 ; n6654
g6399 and n6451_not n6654_not ; n6655
g6400 and n6652_not n6655 ; n6656
g6401 and n6451_not n6656_not ; n6657
g6402 and b[16] n6440_not ; n6658
g6403 and n6434_not n6658 ; n6659
g6404 and n6442_not n6659_not ; n6660
g6405 and n6657_not n6660 ; n6661
g6406 and n6442_not n6661_not ; n6662
g6407 and b[17] n6431_not ; n6663
g6408 and n6425_not n6663 ; n6664
g6409 and n6433_not n6664_not ; n6665
g6410 and n6662_not n6665 ; n6666
g6411 and n6433_not n6666_not ; n6667
g6412 and b[18] n6422_not ; n6668
g6413 and n6416_not n6668 ; n6669
g6414 and n6424_not n6669_not ; n6670
g6415 and n6667_not n6670 ; n6671
g6416 and n6424_not n6671_not ; n6672
g6417 and b[19] n6413_not ; n6673
g6418 and n6407_not n6673 ; n6674
g6419 and n6415_not n6674_not ; n6675
g6420 and n6672_not n6675 ; n6676
g6421 and n6415_not n6676_not ; n6677
g6422 and b[20] n6404_not ; n6678
g6423 and n6398_not n6678 ; n6679
g6424 and n6406_not n6679_not ; n6680
g6425 and n6677_not n6680 ; n6681
g6426 and n6406_not n6681_not ; n6682
g6427 and b[21] n6395_not ; n6683
g6428 and n6389_not n6683 ; n6684
g6429 and n6397_not n6684_not ; n6685
g6430 and n6682_not n6685 ; n6686
g6431 and n6397_not n6686_not ; n6687
g6432 and b[22] n6386_not ; n6688
g6433 and n6380_not n6688 ; n6689
g6434 and n6388_not n6689_not ; n6690
g6435 and n6687_not n6690 ; n6691
g6436 and n6388_not n6691_not ; n6692
g6437 and b[23] n6377_not ; n6693
g6438 and n6371_not n6693 ; n6694
g6439 and n6379_not n6694_not ; n6695
g6440 and n6692_not n6695 ; n6696
g6441 and n6379_not n6696_not ; n6697
g6442 and b[24] n6368_not ; n6698
g6443 and n6362_not n6698 ; n6699
g6444 and n6370_not n6699_not ; n6700
g6445 and n6697_not n6700 ; n6701
g6446 and n6370_not n6701_not ; n6702
g6447 and b[25] n6359_not ; n6703
g6448 and n6353_not n6703 ; n6704
g6449 and n6361_not n6704_not ; n6705
g6450 and n6702_not n6705 ; n6706
g6451 and n6361_not n6706_not ; n6707
g6452 and b[26] n6350_not ; n6708
g6453 and n6344_not n6708 ; n6709
g6454 and n6352_not n6709_not ; n6710
g6455 and n6707_not n6710 ; n6711
g6456 and n6352_not n6711_not ; n6712
g6457 and b[27] n6341_not ; n6713
g6458 and n6335_not n6713 ; n6714
g6459 and n6343_not n6714_not ; n6715
g6460 and n6712_not n6715 ; n6716
g6461 and n6343_not n6716_not ; n6717
g6462 and b[28] n6332_not ; n6718
g6463 and n6326_not n6718 ; n6719
g6464 and n6334_not n6719_not ; n6720
g6465 and n6717_not n6720 ; n6721
g6466 and n6334_not n6721_not ; n6722
g6467 and n5942_not quotient[35]_not ; n6723
g6468 and n5944_not n6320 ; n6724
g6469 and n6316_not n6724 ; n6725
g6470 and n6317_not n6320_not ; n6726
g6471 and n6725_not n6726_not ; n6727
g6472 and quotient[35] n6727_not ; n6728
g6473 and n6723_not n6728_not ; n6729
g6474 and b[29]_not n6729_not ; n6730
g6475 and b[29] n6723_not ; n6731
g6476 and n6728_not n6731 ; n6732
g6477 and n313 n315 ; n6733
g6478 and n303 n6733 ; n6734
g6479 and n288 n6734 ; n6735
g6480 and n6732_not n6735 ; n6736
g6481 and n6730_not n6736 ; n6737
g6482 and n6722_not n6737 ; n6738
g6483 and n6324 n6729_not ; n6739
g6484 and n6738_not n6739_not ; quotient[34]
g6485 and n6343_not n6720 ; n6741
g6486 and n6716_not n6741 ; n6742
g6487 and n6717_not n6720_not ; n6743
g6488 and n6742_not n6743_not ; n6744
g6489 and quotient[34] n6744_not ; n6745
g6490 and n6333_not n6739_not ; n6746
g6491 and n6738_not n6746 ; n6747
g6492 and n6745_not n6747_not ; n6748
g6493 and n6334_not n6732_not ; n6749
g6494 and n6730_not n6749 ; n6750
g6495 and n6721_not n6750 ; n6751
g6496 and n6730_not n6732_not ; n6752
g6497 and n6722_not n6752_not ; n6753
g6498 and n6751_not n6753_not ; n6754
g6499 and quotient[34] n6754_not ; n6755
g6500 and n6729_not n6739_not ; n6756
g6501 and n6738_not n6756 ; n6757
g6502 and n6755_not n6757_not ; n6758
g6503 and b[30]_not n6758_not ; n6759
g6504 and b[29]_not n6748_not ; n6760
g6505 and n6352_not n6715 ; n6761
g6506 and n6711_not n6761 ; n6762
g6507 and n6712_not n6715_not ; n6763
g6508 and n6762_not n6763_not ; n6764
g6509 and quotient[34] n6764_not ; n6765
g6510 and n6342_not n6739_not ; n6766
g6511 and n6738_not n6766 ; n6767
g6512 and n6765_not n6767_not ; n6768
g6513 and b[28]_not n6768_not ; n6769
g6514 and n6361_not n6710 ; n6770
g6515 and n6706_not n6770 ; n6771
g6516 and n6707_not n6710_not ; n6772
g6517 and n6771_not n6772_not ; n6773
g6518 and quotient[34] n6773_not ; n6774
g6519 and n6351_not n6739_not ; n6775
g6520 and n6738_not n6775 ; n6776
g6521 and n6774_not n6776_not ; n6777
g6522 and b[27]_not n6777_not ; n6778
g6523 and n6370_not n6705 ; n6779
g6524 and n6701_not n6779 ; n6780
g6525 and n6702_not n6705_not ; n6781
g6526 and n6780_not n6781_not ; n6782
g6527 and quotient[34] n6782_not ; n6783
g6528 and n6360_not n6739_not ; n6784
g6529 and n6738_not n6784 ; n6785
g6530 and n6783_not n6785_not ; n6786
g6531 and b[26]_not n6786_not ; n6787
g6532 and n6379_not n6700 ; n6788
g6533 and n6696_not n6788 ; n6789
g6534 and n6697_not n6700_not ; n6790
g6535 and n6789_not n6790_not ; n6791
g6536 and quotient[34] n6791_not ; n6792
g6537 and n6369_not n6739_not ; n6793
g6538 and n6738_not n6793 ; n6794
g6539 and n6792_not n6794_not ; n6795
g6540 and b[25]_not n6795_not ; n6796
g6541 and n6388_not n6695 ; n6797
g6542 and n6691_not n6797 ; n6798
g6543 and n6692_not n6695_not ; n6799
g6544 and n6798_not n6799_not ; n6800
g6545 and quotient[34] n6800_not ; n6801
g6546 and n6378_not n6739_not ; n6802
g6547 and n6738_not n6802 ; n6803
g6548 and n6801_not n6803_not ; n6804
g6549 and b[24]_not n6804_not ; n6805
g6550 and n6397_not n6690 ; n6806
g6551 and n6686_not n6806 ; n6807
g6552 and n6687_not n6690_not ; n6808
g6553 and n6807_not n6808_not ; n6809
g6554 and quotient[34] n6809_not ; n6810
g6555 and n6387_not n6739_not ; n6811
g6556 and n6738_not n6811 ; n6812
g6557 and n6810_not n6812_not ; n6813
g6558 and b[23]_not n6813_not ; n6814
g6559 and n6406_not n6685 ; n6815
g6560 and n6681_not n6815 ; n6816
g6561 and n6682_not n6685_not ; n6817
g6562 and n6816_not n6817_not ; n6818
g6563 and quotient[34] n6818_not ; n6819
g6564 and n6396_not n6739_not ; n6820
g6565 and n6738_not n6820 ; n6821
g6566 and n6819_not n6821_not ; n6822
g6567 and b[22]_not n6822_not ; n6823
g6568 and n6415_not n6680 ; n6824
g6569 and n6676_not n6824 ; n6825
g6570 and n6677_not n6680_not ; n6826
g6571 and n6825_not n6826_not ; n6827
g6572 and quotient[34] n6827_not ; n6828
g6573 and n6405_not n6739_not ; n6829
g6574 and n6738_not n6829 ; n6830
g6575 and n6828_not n6830_not ; n6831
g6576 and b[21]_not n6831_not ; n6832
g6577 and n6424_not n6675 ; n6833
g6578 and n6671_not n6833 ; n6834
g6579 and n6672_not n6675_not ; n6835
g6580 and n6834_not n6835_not ; n6836
g6581 and quotient[34] n6836_not ; n6837
g6582 and n6414_not n6739_not ; n6838
g6583 and n6738_not n6838 ; n6839
g6584 and n6837_not n6839_not ; n6840
g6585 and b[20]_not n6840_not ; n6841
g6586 and n6433_not n6670 ; n6842
g6587 and n6666_not n6842 ; n6843
g6588 and n6667_not n6670_not ; n6844
g6589 and n6843_not n6844_not ; n6845
g6590 and quotient[34] n6845_not ; n6846
g6591 and n6423_not n6739_not ; n6847
g6592 and n6738_not n6847 ; n6848
g6593 and n6846_not n6848_not ; n6849
g6594 and b[19]_not n6849_not ; n6850
g6595 and n6442_not n6665 ; n6851
g6596 and n6661_not n6851 ; n6852
g6597 and n6662_not n6665_not ; n6853
g6598 and n6852_not n6853_not ; n6854
g6599 and quotient[34] n6854_not ; n6855
g6600 and n6432_not n6739_not ; n6856
g6601 and n6738_not n6856 ; n6857
g6602 and n6855_not n6857_not ; n6858
g6603 and b[18]_not n6858_not ; n6859
g6604 and n6451_not n6660 ; n6860
g6605 and n6656_not n6860 ; n6861
g6606 and n6657_not n6660_not ; n6862
g6607 and n6861_not n6862_not ; n6863
g6608 and quotient[34] n6863_not ; n6864
g6609 and n6441_not n6739_not ; n6865
g6610 and n6738_not n6865 ; n6866
g6611 and n6864_not n6866_not ; n6867
g6612 and b[17]_not n6867_not ; n6868
g6613 and n6460_not n6655 ; n6869
g6614 and n6651_not n6869 ; n6870
g6615 and n6652_not n6655_not ; n6871
g6616 and n6870_not n6871_not ; n6872
g6617 and quotient[34] n6872_not ; n6873
g6618 and n6450_not n6739_not ; n6874
g6619 and n6738_not n6874 ; n6875
g6620 and n6873_not n6875_not ; n6876
g6621 and b[16]_not n6876_not ; n6877
g6622 and n6469_not n6650 ; n6878
g6623 and n6646_not n6878 ; n6879
g6624 and n6647_not n6650_not ; n6880
g6625 and n6879_not n6880_not ; n6881
g6626 and quotient[34] n6881_not ; n6882
g6627 and n6459_not n6739_not ; n6883
g6628 and n6738_not n6883 ; n6884
g6629 and n6882_not n6884_not ; n6885
g6630 and b[15]_not n6885_not ; n6886
g6631 and n6478_not n6645 ; n6887
g6632 and n6641_not n6887 ; n6888
g6633 and n6642_not n6645_not ; n6889
g6634 and n6888_not n6889_not ; n6890
g6635 and quotient[34] n6890_not ; n6891
g6636 and n6468_not n6739_not ; n6892
g6637 and n6738_not n6892 ; n6893
g6638 and n6891_not n6893_not ; n6894
g6639 and b[14]_not n6894_not ; n6895
g6640 and n6487_not n6640 ; n6896
g6641 and n6636_not n6896 ; n6897
g6642 and n6637_not n6640_not ; n6898
g6643 and n6897_not n6898_not ; n6899
g6644 and quotient[34] n6899_not ; n6900
g6645 and n6477_not n6739_not ; n6901
g6646 and n6738_not n6901 ; n6902
g6647 and n6900_not n6902_not ; n6903
g6648 and b[13]_not n6903_not ; n6904
g6649 and n6496_not n6635 ; n6905
g6650 and n6631_not n6905 ; n6906
g6651 and n6632_not n6635_not ; n6907
g6652 and n6906_not n6907_not ; n6908
g6653 and quotient[34] n6908_not ; n6909
g6654 and n6486_not n6739_not ; n6910
g6655 and n6738_not n6910 ; n6911
g6656 and n6909_not n6911_not ; n6912
g6657 and b[12]_not n6912_not ; n6913
g6658 and n6505_not n6630 ; n6914
g6659 and n6626_not n6914 ; n6915
g6660 and n6627_not n6630_not ; n6916
g6661 and n6915_not n6916_not ; n6917
g6662 and quotient[34] n6917_not ; n6918
g6663 and n6495_not n6739_not ; n6919
g6664 and n6738_not n6919 ; n6920
g6665 and n6918_not n6920_not ; n6921
g6666 and b[11]_not n6921_not ; n6922
g6667 and n6514_not n6625 ; n6923
g6668 and n6621_not n6923 ; n6924
g6669 and n6622_not n6625_not ; n6925
g6670 and n6924_not n6925_not ; n6926
g6671 and quotient[34] n6926_not ; n6927
g6672 and n6504_not n6739_not ; n6928
g6673 and n6738_not n6928 ; n6929
g6674 and n6927_not n6929_not ; n6930
g6675 and b[10]_not n6930_not ; n6931
g6676 and n6523_not n6620 ; n6932
g6677 and n6616_not n6932 ; n6933
g6678 and n6617_not n6620_not ; n6934
g6679 and n6933_not n6934_not ; n6935
g6680 and quotient[34] n6935_not ; n6936
g6681 and n6513_not n6739_not ; n6937
g6682 and n6738_not n6937 ; n6938
g6683 and n6936_not n6938_not ; n6939
g6684 and b[9]_not n6939_not ; n6940
g6685 and n6532_not n6615 ; n6941
g6686 and n6611_not n6941 ; n6942
g6687 and n6612_not n6615_not ; n6943
g6688 and n6942_not n6943_not ; n6944
g6689 and quotient[34] n6944_not ; n6945
g6690 and n6522_not n6739_not ; n6946
g6691 and n6738_not n6946 ; n6947
g6692 and n6945_not n6947_not ; n6948
g6693 and b[8]_not n6948_not ; n6949
g6694 and n6541_not n6610 ; n6950
g6695 and n6606_not n6950 ; n6951
g6696 and n6607_not n6610_not ; n6952
g6697 and n6951_not n6952_not ; n6953
g6698 and quotient[34] n6953_not ; n6954
g6699 and n6531_not n6739_not ; n6955
g6700 and n6738_not n6955 ; n6956
g6701 and n6954_not n6956_not ; n6957
g6702 and b[7]_not n6957_not ; n6958
g6703 and n6550_not n6605 ; n6959
g6704 and n6601_not n6959 ; n6960
g6705 and n6602_not n6605_not ; n6961
g6706 and n6960_not n6961_not ; n6962
g6707 and quotient[34] n6962_not ; n6963
g6708 and n6540_not n6739_not ; n6964
g6709 and n6738_not n6964 ; n6965
g6710 and n6963_not n6965_not ; n6966
g6711 and b[6]_not n6966_not ; n6967
g6712 and n6559_not n6600 ; n6968
g6713 and n6596_not n6968 ; n6969
g6714 and n6597_not n6600_not ; n6970
g6715 and n6969_not n6970_not ; n6971
g6716 and quotient[34] n6971_not ; n6972
g6717 and n6549_not n6739_not ; n6973
g6718 and n6738_not n6973 ; n6974
g6719 and n6972_not n6974_not ; n6975
g6720 and b[5]_not n6975_not ; n6976
g6721 and n6567_not n6595 ; n6977
g6722 and n6591_not n6977 ; n6978
g6723 and n6592_not n6595_not ; n6979
g6724 and n6978_not n6979_not ; n6980
g6725 and quotient[34] n6980_not ; n6981
g6726 and n6558_not n6739_not ; n6982
g6727 and n6738_not n6982 ; n6983
g6728 and n6981_not n6983_not ; n6984
g6729 and b[4]_not n6984_not ; n6985
g6730 and n6586_not n6590 ; n6986
g6731 and n6585_not n6986 ; n6987
g6732 and n6587_not n6590_not ; n6988
g6733 and n6987_not n6988_not ; n6989
g6734 and quotient[34] n6989_not ; n6990
g6735 and n6566_not n6739_not ; n6991
g6736 and n6738_not n6991 ; n6992
g6737 and n6990_not n6992_not ; n6993
g6738 and b[3]_not n6993_not ; n6994
g6739 and n6582_not n6584 ; n6995
g6740 and n6580_not n6995 ; n6996
g6741 and n6585_not n6996_not ; n6997
g6742 and quotient[34] n6997 ; n6998
g6743 and n6579_not n6739_not ; n6999
g6744 and n6738_not n6999 ; n7000
g6745 and n6998_not n7000_not ; n7001
g6746 and b[2]_not n7001_not ; n7002
g6747 and b[0] quotient[34] ; n7003
g6748 and a[34] n7003_not ; n7004
g6749 and n6584 quotient[34] ; n7005
g6750 and n7004_not n7005_not ; n7006
g6751 and b[1] n7006_not ; n7007
g6752 and b[1]_not n7005_not ; n7008
g6753 and n7004_not n7008 ; n7009
g6754 and n7007_not n7009_not ; n7010
g6755 and a[33]_not b[0] ; n7011
g6756 and n7010_not n7011_not ; n7012
g6757 and b[1]_not n7006_not ; n7013
g6758 and n7012_not n7013_not ; n7014
g6759 and b[2] n7000_not ; n7015
g6760 and n6998_not n7015 ; n7016
g6761 and n7002_not n7016_not ; n7017
g6762 and n7014_not n7017 ; n7018
g6763 and n7002_not n7018_not ; n7019
g6764 and b[3] n6992_not ; n7020
g6765 and n6990_not n7020 ; n7021
g6766 and n6994_not n7021_not ; n7022
g6767 and n7019_not n7022 ; n7023
g6768 and n6994_not n7023_not ; n7024
g6769 and b[4] n6983_not ; n7025
g6770 and n6981_not n7025 ; n7026
g6771 and n6985_not n7026_not ; n7027
g6772 and n7024_not n7027 ; n7028
g6773 and n6985_not n7028_not ; n7029
g6774 and b[5] n6974_not ; n7030
g6775 and n6972_not n7030 ; n7031
g6776 and n6976_not n7031_not ; n7032
g6777 and n7029_not n7032 ; n7033
g6778 and n6976_not n7033_not ; n7034
g6779 and b[6] n6965_not ; n7035
g6780 and n6963_not n7035 ; n7036
g6781 and n6967_not n7036_not ; n7037
g6782 and n7034_not n7037 ; n7038
g6783 and n6967_not n7038_not ; n7039
g6784 and b[7] n6956_not ; n7040
g6785 and n6954_not n7040 ; n7041
g6786 and n6958_not n7041_not ; n7042
g6787 and n7039_not n7042 ; n7043
g6788 and n6958_not n7043_not ; n7044
g6789 and b[8] n6947_not ; n7045
g6790 and n6945_not n7045 ; n7046
g6791 and n6949_not n7046_not ; n7047
g6792 and n7044_not n7047 ; n7048
g6793 and n6949_not n7048_not ; n7049
g6794 and b[9] n6938_not ; n7050
g6795 and n6936_not n7050 ; n7051
g6796 and n6940_not n7051_not ; n7052
g6797 and n7049_not n7052 ; n7053
g6798 and n6940_not n7053_not ; n7054
g6799 and b[10] n6929_not ; n7055
g6800 and n6927_not n7055 ; n7056
g6801 and n6931_not n7056_not ; n7057
g6802 and n7054_not n7057 ; n7058
g6803 and n6931_not n7058_not ; n7059
g6804 and b[11] n6920_not ; n7060
g6805 and n6918_not n7060 ; n7061
g6806 and n6922_not n7061_not ; n7062
g6807 and n7059_not n7062 ; n7063
g6808 and n6922_not n7063_not ; n7064
g6809 and b[12] n6911_not ; n7065
g6810 and n6909_not n7065 ; n7066
g6811 and n6913_not n7066_not ; n7067
g6812 and n7064_not n7067 ; n7068
g6813 and n6913_not n7068_not ; n7069
g6814 and b[13] n6902_not ; n7070
g6815 and n6900_not n7070 ; n7071
g6816 and n6904_not n7071_not ; n7072
g6817 and n7069_not n7072 ; n7073
g6818 and n6904_not n7073_not ; n7074
g6819 and b[14] n6893_not ; n7075
g6820 and n6891_not n7075 ; n7076
g6821 and n6895_not n7076_not ; n7077
g6822 and n7074_not n7077 ; n7078
g6823 and n6895_not n7078_not ; n7079
g6824 and b[15] n6884_not ; n7080
g6825 and n6882_not n7080 ; n7081
g6826 and n6886_not n7081_not ; n7082
g6827 and n7079_not n7082 ; n7083
g6828 and n6886_not n7083_not ; n7084
g6829 and b[16] n6875_not ; n7085
g6830 and n6873_not n7085 ; n7086
g6831 and n6877_not n7086_not ; n7087
g6832 and n7084_not n7087 ; n7088
g6833 and n6877_not n7088_not ; n7089
g6834 and b[17] n6866_not ; n7090
g6835 and n6864_not n7090 ; n7091
g6836 and n6868_not n7091_not ; n7092
g6837 and n7089_not n7092 ; n7093
g6838 and n6868_not n7093_not ; n7094
g6839 and b[18] n6857_not ; n7095
g6840 and n6855_not n7095 ; n7096
g6841 and n6859_not n7096_not ; n7097
g6842 and n7094_not n7097 ; n7098
g6843 and n6859_not n7098_not ; n7099
g6844 and b[19] n6848_not ; n7100
g6845 and n6846_not n7100 ; n7101
g6846 and n6850_not n7101_not ; n7102
g6847 and n7099_not n7102 ; n7103
g6848 and n6850_not n7103_not ; n7104
g6849 and b[20] n6839_not ; n7105
g6850 and n6837_not n7105 ; n7106
g6851 and n6841_not n7106_not ; n7107
g6852 and n7104_not n7107 ; n7108
g6853 and n6841_not n7108_not ; n7109
g6854 and b[21] n6830_not ; n7110
g6855 and n6828_not n7110 ; n7111
g6856 and n6832_not n7111_not ; n7112
g6857 and n7109_not n7112 ; n7113
g6858 and n6832_not n7113_not ; n7114
g6859 and b[22] n6821_not ; n7115
g6860 and n6819_not n7115 ; n7116
g6861 and n6823_not n7116_not ; n7117
g6862 and n7114_not n7117 ; n7118
g6863 and n6823_not n7118_not ; n7119
g6864 and b[23] n6812_not ; n7120
g6865 and n6810_not n7120 ; n7121
g6866 and n6814_not n7121_not ; n7122
g6867 and n7119_not n7122 ; n7123
g6868 and n6814_not n7123_not ; n7124
g6869 and b[24] n6803_not ; n7125
g6870 and n6801_not n7125 ; n7126
g6871 and n6805_not n7126_not ; n7127
g6872 and n7124_not n7127 ; n7128
g6873 and n6805_not n7128_not ; n7129
g6874 and b[25] n6794_not ; n7130
g6875 and n6792_not n7130 ; n7131
g6876 and n6796_not n7131_not ; n7132
g6877 and n7129_not n7132 ; n7133
g6878 and n6796_not n7133_not ; n7134
g6879 and b[26] n6785_not ; n7135
g6880 and n6783_not n7135 ; n7136
g6881 and n6787_not n7136_not ; n7137
g6882 and n7134_not n7137 ; n7138
g6883 and n6787_not n7138_not ; n7139
g6884 and b[27] n6776_not ; n7140
g6885 and n6774_not n7140 ; n7141
g6886 and n6778_not n7141_not ; n7142
g6887 and n7139_not n7142 ; n7143
g6888 and n6778_not n7143_not ; n7144
g6889 and b[28] n6767_not ; n7145
g6890 and n6765_not n7145 ; n7146
g6891 and n6769_not n7146_not ; n7147
g6892 and n7144_not n7147 ; n7148
g6893 and n6769_not n7148_not ; n7149
g6894 and b[29] n6747_not ; n7150
g6895 and n6745_not n7150 ; n7151
g6896 and n6760_not n7151_not ; n7152
g6897 and n7149_not n7152 ; n7153
g6898 and n6760_not n7153_not ; n7154
g6899 and b[30] n6757_not ; n7155
g6900 and n6755_not n7155 ; n7156
g6901 and n6759_not n7156_not ; n7157
g6902 and n7154_not n7157 ; n7158
g6903 and n6759_not n7158_not ; n7159
g6904 and n372 n414 ; n7160
g6905 and n598 n7160 ; n7161
g6906 and n595 n7161 ; n7162
g6907 and n7159_not n7162 ; quotient[33]
g6908 and n6748_not quotient[33]_not ; n7164
g6909 and n6769_not n7152 ; n7165
g6910 and n7148_not n7165 ; n7166
g6911 and n7149_not n7152_not ; n7167
g6912 and n7166_not n7167_not ; n7168
g6913 and n7162 n7168_not ; n7169
g6914 and n7159_not n7169 ; n7170
g6915 and n7164_not n7170_not ; n7171
g6916 and n6758_not quotient[33]_not ; n7172
g6917 and n6760_not n7157 ; n7173
g6918 and n7153_not n7173 ; n7174
g6919 and n7154_not n7157_not ; n7175
g6920 and n7174_not n7175_not ; n7176
g6921 and quotient[33] n7176_not ; n7177
g6922 and n7172_not n7177_not ; n7178
g6923 and b[31]_not n7178_not ; n7179
g6924 and b[30]_not n7171_not ; n7180
g6925 and n6768_not quotient[33]_not ; n7181
g6926 and n6778_not n7147 ; n7182
g6927 and n7143_not n7182 ; n7183
g6928 and n7144_not n7147_not ; n7184
g6929 and n7183_not n7184_not ; n7185
g6930 and n7162 n7185_not ; n7186
g6931 and n7159_not n7186 ; n7187
g6932 and n7181_not n7187_not ; n7188
g6933 and b[29]_not n7188_not ; n7189
g6934 and n6777_not quotient[33]_not ; n7190
g6935 and n6787_not n7142 ; n7191
g6936 and n7138_not n7191 ; n7192
g6937 and n7139_not n7142_not ; n7193
g6938 and n7192_not n7193_not ; n7194
g6939 and n7162 n7194_not ; n7195
g6940 and n7159_not n7195 ; n7196
g6941 and n7190_not n7196_not ; n7197
g6942 and b[28]_not n7197_not ; n7198
g6943 and n6786_not quotient[33]_not ; n7199
g6944 and n6796_not n7137 ; n7200
g6945 and n7133_not n7200 ; n7201
g6946 and n7134_not n7137_not ; n7202
g6947 and n7201_not n7202_not ; n7203
g6948 and n7162 n7203_not ; n7204
g6949 and n7159_not n7204 ; n7205
g6950 and n7199_not n7205_not ; n7206
g6951 and b[27]_not n7206_not ; n7207
g6952 and n6795_not quotient[33]_not ; n7208
g6953 and n6805_not n7132 ; n7209
g6954 and n7128_not n7209 ; n7210
g6955 and n7129_not n7132_not ; n7211
g6956 and n7210_not n7211_not ; n7212
g6957 and n7162 n7212_not ; n7213
g6958 and n7159_not n7213 ; n7214
g6959 and n7208_not n7214_not ; n7215
g6960 and b[26]_not n7215_not ; n7216
g6961 and n6804_not quotient[33]_not ; n7217
g6962 and n6814_not n7127 ; n7218
g6963 and n7123_not n7218 ; n7219
g6964 and n7124_not n7127_not ; n7220
g6965 and n7219_not n7220_not ; n7221
g6966 and n7162 n7221_not ; n7222
g6967 and n7159_not n7222 ; n7223
g6968 and n7217_not n7223_not ; n7224
g6969 and b[25]_not n7224_not ; n7225
g6970 and n6813_not quotient[33]_not ; n7226
g6971 and n6823_not n7122 ; n7227
g6972 and n7118_not n7227 ; n7228
g6973 and n7119_not n7122_not ; n7229
g6974 and n7228_not n7229_not ; n7230
g6975 and n7162 n7230_not ; n7231
g6976 and n7159_not n7231 ; n7232
g6977 and n7226_not n7232_not ; n7233
g6978 and b[24]_not n7233_not ; n7234
g6979 and n6822_not quotient[33]_not ; n7235
g6980 and n6832_not n7117 ; n7236
g6981 and n7113_not n7236 ; n7237
g6982 and n7114_not n7117_not ; n7238
g6983 and n7237_not n7238_not ; n7239
g6984 and n7162 n7239_not ; n7240
g6985 and n7159_not n7240 ; n7241
g6986 and n7235_not n7241_not ; n7242
g6987 and b[23]_not n7242_not ; n7243
g6988 and n6831_not quotient[33]_not ; n7244
g6989 and n6841_not n7112 ; n7245
g6990 and n7108_not n7245 ; n7246
g6991 and n7109_not n7112_not ; n7247
g6992 and n7246_not n7247_not ; n7248
g6993 and n7162 n7248_not ; n7249
g6994 and n7159_not n7249 ; n7250
g6995 and n7244_not n7250_not ; n7251
g6996 and b[22]_not n7251_not ; n7252
g6997 and n6840_not quotient[33]_not ; n7253
g6998 and n6850_not n7107 ; n7254
g6999 and n7103_not n7254 ; n7255
g7000 and n7104_not n7107_not ; n7256
g7001 and n7255_not n7256_not ; n7257
g7002 and n7162 n7257_not ; n7258
g7003 and n7159_not n7258 ; n7259
g7004 and n7253_not n7259_not ; n7260
g7005 and b[21]_not n7260_not ; n7261
g7006 and n6849_not quotient[33]_not ; n7262
g7007 and n6859_not n7102 ; n7263
g7008 and n7098_not n7263 ; n7264
g7009 and n7099_not n7102_not ; n7265
g7010 and n7264_not n7265_not ; n7266
g7011 and n7162 n7266_not ; n7267
g7012 and n7159_not n7267 ; n7268
g7013 and n7262_not n7268_not ; n7269
g7014 and b[20]_not n7269_not ; n7270
g7015 and n6858_not quotient[33]_not ; n7271
g7016 and n6868_not n7097 ; n7272
g7017 and n7093_not n7272 ; n7273
g7018 and n7094_not n7097_not ; n7274
g7019 and n7273_not n7274_not ; n7275
g7020 and n7162 n7275_not ; n7276
g7021 and n7159_not n7276 ; n7277
g7022 and n7271_not n7277_not ; n7278
g7023 and b[19]_not n7278_not ; n7279
g7024 and n6867_not quotient[33]_not ; n7280
g7025 and n6877_not n7092 ; n7281
g7026 and n7088_not n7281 ; n7282
g7027 and n7089_not n7092_not ; n7283
g7028 and n7282_not n7283_not ; n7284
g7029 and n7162 n7284_not ; n7285
g7030 and n7159_not n7285 ; n7286
g7031 and n7280_not n7286_not ; n7287
g7032 and b[18]_not n7287_not ; n7288
g7033 and n6876_not quotient[33]_not ; n7289
g7034 and n6886_not n7087 ; n7290
g7035 and n7083_not n7290 ; n7291
g7036 and n7084_not n7087_not ; n7292
g7037 and n7291_not n7292_not ; n7293
g7038 and n7162 n7293_not ; n7294
g7039 and n7159_not n7294 ; n7295
g7040 and n7289_not n7295_not ; n7296
g7041 and b[17]_not n7296_not ; n7297
g7042 and n6885_not quotient[33]_not ; n7298
g7043 and n6895_not n7082 ; n7299
g7044 and n7078_not n7299 ; n7300
g7045 and n7079_not n7082_not ; n7301
g7046 and n7300_not n7301_not ; n7302
g7047 and n7162 n7302_not ; n7303
g7048 and n7159_not n7303 ; n7304
g7049 and n7298_not n7304_not ; n7305
g7050 and b[16]_not n7305_not ; n7306
g7051 and n6894_not quotient[33]_not ; n7307
g7052 and n6904_not n7077 ; n7308
g7053 and n7073_not n7308 ; n7309
g7054 and n7074_not n7077_not ; n7310
g7055 and n7309_not n7310_not ; n7311
g7056 and n7162 n7311_not ; n7312
g7057 and n7159_not n7312 ; n7313
g7058 and n7307_not n7313_not ; n7314
g7059 and b[15]_not n7314_not ; n7315
g7060 and n6903_not quotient[33]_not ; n7316
g7061 and n6913_not n7072 ; n7317
g7062 and n7068_not n7317 ; n7318
g7063 and n7069_not n7072_not ; n7319
g7064 and n7318_not n7319_not ; n7320
g7065 and n7162 n7320_not ; n7321
g7066 and n7159_not n7321 ; n7322
g7067 and n7316_not n7322_not ; n7323
g7068 and b[14]_not n7323_not ; n7324
g7069 and n6912_not quotient[33]_not ; n7325
g7070 and n6922_not n7067 ; n7326
g7071 and n7063_not n7326 ; n7327
g7072 and n7064_not n7067_not ; n7328
g7073 and n7327_not n7328_not ; n7329
g7074 and n7162 n7329_not ; n7330
g7075 and n7159_not n7330 ; n7331
g7076 and n7325_not n7331_not ; n7332
g7077 and b[13]_not n7332_not ; n7333
g7078 and n6921_not quotient[33]_not ; n7334
g7079 and n6931_not n7062 ; n7335
g7080 and n7058_not n7335 ; n7336
g7081 and n7059_not n7062_not ; n7337
g7082 and n7336_not n7337_not ; n7338
g7083 and n7162 n7338_not ; n7339
g7084 and n7159_not n7339 ; n7340
g7085 and n7334_not n7340_not ; n7341
g7086 and b[12]_not n7341_not ; n7342
g7087 and n6930_not quotient[33]_not ; n7343
g7088 and n6940_not n7057 ; n7344
g7089 and n7053_not n7344 ; n7345
g7090 and n7054_not n7057_not ; n7346
g7091 and n7345_not n7346_not ; n7347
g7092 and n7162 n7347_not ; n7348
g7093 and n7159_not n7348 ; n7349
g7094 and n7343_not n7349_not ; n7350
g7095 and b[11]_not n7350_not ; n7351
g7096 and n6939_not quotient[33]_not ; n7352
g7097 and n6949_not n7052 ; n7353
g7098 and n7048_not n7353 ; n7354
g7099 and n7049_not n7052_not ; n7355
g7100 and n7354_not n7355_not ; n7356
g7101 and n7162 n7356_not ; n7357
g7102 and n7159_not n7357 ; n7358
g7103 and n7352_not n7358_not ; n7359
g7104 and b[10]_not n7359_not ; n7360
g7105 and n6948_not quotient[33]_not ; n7361
g7106 and n6958_not n7047 ; n7362
g7107 and n7043_not n7362 ; n7363
g7108 and n7044_not n7047_not ; n7364
g7109 and n7363_not n7364_not ; n7365
g7110 and n7162 n7365_not ; n7366
g7111 and n7159_not n7366 ; n7367
g7112 and n7361_not n7367_not ; n7368
g7113 and b[9]_not n7368_not ; n7369
g7114 and n6957_not quotient[33]_not ; n7370
g7115 and n6967_not n7042 ; n7371
g7116 and n7038_not n7371 ; n7372
g7117 and n7039_not n7042_not ; n7373
g7118 and n7372_not n7373_not ; n7374
g7119 and n7162 n7374_not ; n7375
g7120 and n7159_not n7375 ; n7376
g7121 and n7370_not n7376_not ; n7377
g7122 and b[8]_not n7377_not ; n7378
g7123 and n6966_not quotient[33]_not ; n7379
g7124 and n6976_not n7037 ; n7380
g7125 and n7033_not n7380 ; n7381
g7126 and n7034_not n7037_not ; n7382
g7127 and n7381_not n7382_not ; n7383
g7128 and n7162 n7383_not ; n7384
g7129 and n7159_not n7384 ; n7385
g7130 and n7379_not n7385_not ; n7386
g7131 and b[7]_not n7386_not ; n7387
g7132 and n6975_not quotient[33]_not ; n7388
g7133 and n6985_not n7032 ; n7389
g7134 and n7028_not n7389 ; n7390
g7135 and n7029_not n7032_not ; n7391
g7136 and n7390_not n7391_not ; n7392
g7137 and n7162 n7392_not ; n7393
g7138 and n7159_not n7393 ; n7394
g7139 and n7388_not n7394_not ; n7395
g7140 and b[6]_not n7395_not ; n7396
g7141 and n6984_not quotient[33]_not ; n7397
g7142 and n6994_not n7027 ; n7398
g7143 and n7023_not n7398 ; n7399
g7144 and n7024_not n7027_not ; n7400
g7145 and n7399_not n7400_not ; n7401
g7146 and n7162 n7401_not ; n7402
g7147 and n7159_not n7402 ; n7403
g7148 and n7397_not n7403_not ; n7404
g7149 and b[5]_not n7404_not ; n7405
g7150 and n6993_not quotient[33]_not ; n7406
g7151 and n7002_not n7022 ; n7407
g7152 and n7018_not n7407 ; n7408
g7153 and n7019_not n7022_not ; n7409
g7154 and n7408_not n7409_not ; n7410
g7155 and n7162 n7410_not ; n7411
g7156 and n7159_not n7411 ; n7412
g7157 and n7406_not n7412_not ; n7413
g7158 and b[4]_not n7413_not ; n7414
g7159 and n7001_not quotient[33]_not ; n7415
g7160 and n7013_not n7017 ; n7416
g7161 and n7012_not n7416 ; n7417
g7162 and n7014_not n7017_not ; n7418
g7163 and n7417_not n7418_not ; n7419
g7164 and n7162 n7419_not ; n7420
g7165 and n7159_not n7420 ; n7421
g7166 and n7415_not n7421_not ; n7422
g7167 and b[3]_not n7422_not ; n7423
g7168 and n7006_not quotient[33]_not ; n7424
g7169 and n7009_not n7011 ; n7425
g7170 and n7007_not n7425 ; n7426
g7171 and n7162 n7426_not ; n7427
g7172 and n7012_not n7427 ; n7428
g7173 and n7159_not n7428 ; n7429
g7174 and n7424_not n7429_not ; n7430
g7175 and b[2]_not n7430_not ; n7431
g7176 and b[0] b[31]_not ; n7432
g7177 and n313 n7432 ; n7433
g7178 and n303 n7433 ; n7434
g7179 and n288 n7434 ; n7435
g7180 and n7159_not n7435 ; n7436
g7181 and a[33] n7436_not ; n7437
g7182 and n372 n7011 ; n7438
g7183 and n414 n7438 ; n7439
g7184 and n598 n7439 ; n7440
g7185 and n595 n7440 ; n7441
g7186 and n7159_not n7441 ; n7442
g7187 and n7437_not n7442_not ; n7443
g7188 and b[1] n7443_not ; n7444
g7189 and b[1]_not n7442_not ; n7445
g7190 and n7437_not n7445 ; n7446
g7191 and n7444_not n7446_not ; n7447
g7192 and a[32]_not b[0] ; n7448
g7193 and n7447_not n7448_not ; n7449
g7194 and b[1]_not n7443_not ; n7450
g7195 and n7449_not n7450_not ; n7451
g7196 and b[2] n7429_not ; n7452
g7197 and n7424_not n7452 ; n7453
g7198 and n7431_not n7453_not ; n7454
g7199 and n7451_not n7454 ; n7455
g7200 and n7431_not n7455_not ; n7456
g7201 and b[3] n7421_not ; n7457
g7202 and n7415_not n7457 ; n7458
g7203 and n7423_not n7458_not ; n7459
g7204 and n7456_not n7459 ; n7460
g7205 and n7423_not n7460_not ; n7461
g7206 and b[4] n7412_not ; n7462
g7207 and n7406_not n7462 ; n7463
g7208 and n7414_not n7463_not ; n7464
g7209 and n7461_not n7464 ; n7465
g7210 and n7414_not n7465_not ; n7466
g7211 and b[5] n7403_not ; n7467
g7212 and n7397_not n7467 ; n7468
g7213 and n7405_not n7468_not ; n7469
g7214 and n7466_not n7469 ; n7470
g7215 and n7405_not n7470_not ; n7471
g7216 and b[6] n7394_not ; n7472
g7217 and n7388_not n7472 ; n7473
g7218 and n7396_not n7473_not ; n7474
g7219 and n7471_not n7474 ; n7475
g7220 and n7396_not n7475_not ; n7476
g7221 and b[7] n7385_not ; n7477
g7222 and n7379_not n7477 ; n7478
g7223 and n7387_not n7478_not ; n7479
g7224 and n7476_not n7479 ; n7480
g7225 and n7387_not n7480_not ; n7481
g7226 and b[8] n7376_not ; n7482
g7227 and n7370_not n7482 ; n7483
g7228 and n7378_not n7483_not ; n7484
g7229 and n7481_not n7484 ; n7485
g7230 and n7378_not n7485_not ; n7486
g7231 and b[9] n7367_not ; n7487
g7232 and n7361_not n7487 ; n7488
g7233 and n7369_not n7488_not ; n7489
g7234 and n7486_not n7489 ; n7490
g7235 and n7369_not n7490_not ; n7491
g7236 and b[10] n7358_not ; n7492
g7237 and n7352_not n7492 ; n7493
g7238 and n7360_not n7493_not ; n7494
g7239 and n7491_not n7494 ; n7495
g7240 and n7360_not n7495_not ; n7496
g7241 and b[11] n7349_not ; n7497
g7242 and n7343_not n7497 ; n7498
g7243 and n7351_not n7498_not ; n7499
g7244 and n7496_not n7499 ; n7500
g7245 and n7351_not n7500_not ; n7501
g7246 and b[12] n7340_not ; n7502
g7247 and n7334_not n7502 ; n7503
g7248 and n7342_not n7503_not ; n7504
g7249 and n7501_not n7504 ; n7505
g7250 and n7342_not n7505_not ; n7506
g7251 and b[13] n7331_not ; n7507
g7252 and n7325_not n7507 ; n7508
g7253 and n7333_not n7508_not ; n7509
g7254 and n7506_not n7509 ; n7510
g7255 and n7333_not n7510_not ; n7511
g7256 and b[14] n7322_not ; n7512
g7257 and n7316_not n7512 ; n7513
g7258 and n7324_not n7513_not ; n7514
g7259 and n7511_not n7514 ; n7515
g7260 and n7324_not n7515_not ; n7516
g7261 and b[15] n7313_not ; n7517
g7262 and n7307_not n7517 ; n7518
g7263 and n7315_not n7518_not ; n7519
g7264 and n7516_not n7519 ; n7520
g7265 and n7315_not n7520_not ; n7521
g7266 and b[16] n7304_not ; n7522
g7267 and n7298_not n7522 ; n7523
g7268 and n7306_not n7523_not ; n7524
g7269 and n7521_not n7524 ; n7525
g7270 and n7306_not n7525_not ; n7526
g7271 and b[17] n7295_not ; n7527
g7272 and n7289_not n7527 ; n7528
g7273 and n7297_not n7528_not ; n7529
g7274 and n7526_not n7529 ; n7530
g7275 and n7297_not n7530_not ; n7531
g7276 and b[18] n7286_not ; n7532
g7277 and n7280_not n7532 ; n7533
g7278 and n7288_not n7533_not ; n7534
g7279 and n7531_not n7534 ; n7535
g7280 and n7288_not n7535_not ; n7536
g7281 and b[19] n7277_not ; n7537
g7282 and n7271_not n7537 ; n7538
g7283 and n7279_not n7538_not ; n7539
g7284 and n7536_not n7539 ; n7540
g7285 and n7279_not n7540_not ; n7541
g7286 and b[20] n7268_not ; n7542
g7287 and n7262_not n7542 ; n7543
g7288 and n7270_not n7543_not ; n7544
g7289 and n7541_not n7544 ; n7545
g7290 and n7270_not n7545_not ; n7546
g7291 and b[21] n7259_not ; n7547
g7292 and n7253_not n7547 ; n7548
g7293 and n7261_not n7548_not ; n7549
g7294 and n7546_not n7549 ; n7550
g7295 and n7261_not n7550_not ; n7551
g7296 and b[22] n7250_not ; n7552
g7297 and n7244_not n7552 ; n7553
g7298 and n7252_not n7553_not ; n7554
g7299 and n7551_not n7554 ; n7555
g7300 and n7252_not n7555_not ; n7556
g7301 and b[23] n7241_not ; n7557
g7302 and n7235_not n7557 ; n7558
g7303 and n7243_not n7558_not ; n7559
g7304 and n7556_not n7559 ; n7560
g7305 and n7243_not n7560_not ; n7561
g7306 and b[24] n7232_not ; n7562
g7307 and n7226_not n7562 ; n7563
g7308 and n7234_not n7563_not ; n7564
g7309 and n7561_not n7564 ; n7565
g7310 and n7234_not n7565_not ; n7566
g7311 and b[25] n7223_not ; n7567
g7312 and n7217_not n7567 ; n7568
g7313 and n7225_not n7568_not ; n7569
g7314 and n7566_not n7569 ; n7570
g7315 and n7225_not n7570_not ; n7571
g7316 and b[26] n7214_not ; n7572
g7317 and n7208_not n7572 ; n7573
g7318 and n7216_not n7573_not ; n7574
g7319 and n7571_not n7574 ; n7575
g7320 and n7216_not n7575_not ; n7576
g7321 and b[27] n7205_not ; n7577
g7322 and n7199_not n7577 ; n7578
g7323 and n7207_not n7578_not ; n7579
g7324 and n7576_not n7579 ; n7580
g7325 and n7207_not n7580_not ; n7581
g7326 and b[28] n7196_not ; n7582
g7327 and n7190_not n7582 ; n7583
g7328 and n7198_not n7583_not ; n7584
g7329 and n7581_not n7584 ; n7585
g7330 and n7198_not n7585_not ; n7586
g7331 and b[29] n7187_not ; n7587
g7332 and n7181_not n7587 ; n7588
g7333 and n7189_not n7588_not ; n7589
g7334 and n7586_not n7589 ; n7590
g7335 and n7189_not n7590_not ; n7591
g7336 and b[30] n7170_not ; n7592
g7337 and n7164_not n7592 ; n7593
g7338 and n7180_not n7593_not ; n7594
g7339 and n7591_not n7594 ; n7595
g7340 and n7180_not n7595_not ; n7596
g7341 and b[31] n7172_not ; n7597
g7342 and n7177_not n7597 ; n7598
g7343 and n7179_not n7598_not ; n7599
g7344 and n7596_not n7599 ; n7600
g7345 and n7179_not n7600_not ; n7601
g7346 and n432 n7601_not ; quotient[32]
g7347 and n7171_not quotient[32]_not ; n7603
g7348 and n7189_not n7594 ; n7604
g7349 and n7590_not n7604 ; n7605
g7350 and n7591_not n7594_not ; n7606
g7351 and n7605_not n7606_not ; n7607
g7352 and n432 n7607_not ; n7608
g7353 and n7601_not n7608 ; n7609
g7354 and n7603_not n7609_not ; n7610
g7355 and b[31]_not n7610_not ; n7611
g7356 and n7188_not quotient[32]_not ; n7612
g7357 and n7198_not n7589 ; n7613
g7358 and n7585_not n7613 ; n7614
g7359 and n7586_not n7589_not ; n7615
g7360 and n7614_not n7615_not ; n7616
g7361 and n432 n7616_not ; n7617
g7362 and n7601_not n7617 ; n7618
g7363 and n7612_not n7618_not ; n7619
g7364 and b[30]_not n7619_not ; n7620
g7365 and n7197_not quotient[32]_not ; n7621
g7366 and n7207_not n7584 ; n7622
g7367 and n7580_not n7622 ; n7623
g7368 and n7581_not n7584_not ; n7624
g7369 and n7623_not n7624_not ; n7625
g7370 and n432 n7625_not ; n7626
g7371 and n7601_not n7626 ; n7627
g7372 and n7621_not n7627_not ; n7628
g7373 and b[29]_not n7628_not ; n7629
g7374 and n7206_not quotient[32]_not ; n7630
g7375 and n7216_not n7579 ; n7631
g7376 and n7575_not n7631 ; n7632
g7377 and n7576_not n7579_not ; n7633
g7378 and n7632_not n7633_not ; n7634
g7379 and n432 n7634_not ; n7635
g7380 and n7601_not n7635 ; n7636
g7381 and n7630_not n7636_not ; n7637
g7382 and b[28]_not n7637_not ; n7638
g7383 and n7215_not quotient[32]_not ; n7639
g7384 and n7225_not n7574 ; n7640
g7385 and n7570_not n7640 ; n7641
g7386 and n7571_not n7574_not ; n7642
g7387 and n7641_not n7642_not ; n7643
g7388 and n432 n7643_not ; n7644
g7389 and n7601_not n7644 ; n7645
g7390 and n7639_not n7645_not ; n7646
g7391 and b[27]_not n7646_not ; n7647
g7392 and n7224_not quotient[32]_not ; n7648
g7393 and n7234_not n7569 ; n7649
g7394 and n7565_not n7649 ; n7650
g7395 and n7566_not n7569_not ; n7651
g7396 and n7650_not n7651_not ; n7652
g7397 and n432 n7652_not ; n7653
g7398 and n7601_not n7653 ; n7654
g7399 and n7648_not n7654_not ; n7655
g7400 and b[26]_not n7655_not ; n7656
g7401 and n7233_not quotient[32]_not ; n7657
g7402 and n7243_not n7564 ; n7658
g7403 and n7560_not n7658 ; n7659
g7404 and n7561_not n7564_not ; n7660
g7405 and n7659_not n7660_not ; n7661
g7406 and n432 n7661_not ; n7662
g7407 and n7601_not n7662 ; n7663
g7408 and n7657_not n7663_not ; n7664
g7409 and b[25]_not n7664_not ; n7665
g7410 and n7242_not quotient[32]_not ; n7666
g7411 and n7252_not n7559 ; n7667
g7412 and n7555_not n7667 ; n7668
g7413 and n7556_not n7559_not ; n7669
g7414 and n7668_not n7669_not ; n7670
g7415 and n432 n7670_not ; n7671
g7416 and n7601_not n7671 ; n7672
g7417 and n7666_not n7672_not ; n7673
g7418 and b[24]_not n7673_not ; n7674
g7419 and n7251_not quotient[32]_not ; n7675
g7420 and n7261_not n7554 ; n7676
g7421 and n7550_not n7676 ; n7677
g7422 and n7551_not n7554_not ; n7678
g7423 and n7677_not n7678_not ; n7679
g7424 and n432 n7679_not ; n7680
g7425 and n7601_not n7680 ; n7681
g7426 and n7675_not n7681_not ; n7682
g7427 and b[23]_not n7682_not ; n7683
g7428 and n7260_not quotient[32]_not ; n7684
g7429 and n7270_not n7549 ; n7685
g7430 and n7545_not n7685 ; n7686
g7431 and n7546_not n7549_not ; n7687
g7432 and n7686_not n7687_not ; n7688
g7433 and n432 n7688_not ; n7689
g7434 and n7601_not n7689 ; n7690
g7435 and n7684_not n7690_not ; n7691
g7436 and b[22]_not n7691_not ; n7692
g7437 and n7269_not quotient[32]_not ; n7693
g7438 and n7279_not n7544 ; n7694
g7439 and n7540_not n7694 ; n7695
g7440 and n7541_not n7544_not ; n7696
g7441 and n7695_not n7696_not ; n7697
g7442 and n432 n7697_not ; n7698
g7443 and n7601_not n7698 ; n7699
g7444 and n7693_not n7699_not ; n7700
g7445 and b[21]_not n7700_not ; n7701
g7446 and n7278_not quotient[32]_not ; n7702
g7447 and n7288_not n7539 ; n7703
g7448 and n7535_not n7703 ; n7704
g7449 and n7536_not n7539_not ; n7705
g7450 and n7704_not n7705_not ; n7706
g7451 and n432 n7706_not ; n7707
g7452 and n7601_not n7707 ; n7708
g7453 and n7702_not n7708_not ; n7709
g7454 and b[20]_not n7709_not ; n7710
g7455 and n7287_not quotient[32]_not ; n7711
g7456 and n7297_not n7534 ; n7712
g7457 and n7530_not n7712 ; n7713
g7458 and n7531_not n7534_not ; n7714
g7459 and n7713_not n7714_not ; n7715
g7460 and n432 n7715_not ; n7716
g7461 and n7601_not n7716 ; n7717
g7462 and n7711_not n7717_not ; n7718
g7463 and b[19]_not n7718_not ; n7719
g7464 and n7296_not quotient[32]_not ; n7720
g7465 and n7306_not n7529 ; n7721
g7466 and n7525_not n7721 ; n7722
g7467 and n7526_not n7529_not ; n7723
g7468 and n7722_not n7723_not ; n7724
g7469 and n432 n7724_not ; n7725
g7470 and n7601_not n7725 ; n7726
g7471 and n7720_not n7726_not ; n7727
g7472 and b[18]_not n7727_not ; n7728
g7473 and n7305_not quotient[32]_not ; n7729
g7474 and n7315_not n7524 ; n7730
g7475 and n7520_not n7730 ; n7731
g7476 and n7521_not n7524_not ; n7732
g7477 and n7731_not n7732_not ; n7733
g7478 and n432 n7733_not ; n7734
g7479 and n7601_not n7734 ; n7735
g7480 and n7729_not n7735_not ; n7736
g7481 and b[17]_not n7736_not ; n7737
g7482 and n7314_not quotient[32]_not ; n7738
g7483 and n7324_not n7519 ; n7739
g7484 and n7515_not n7739 ; n7740
g7485 and n7516_not n7519_not ; n7741
g7486 and n7740_not n7741_not ; n7742
g7487 and n432 n7742_not ; n7743
g7488 and n7601_not n7743 ; n7744
g7489 and n7738_not n7744_not ; n7745
g7490 and b[16]_not n7745_not ; n7746
g7491 and n7323_not quotient[32]_not ; n7747
g7492 and n7333_not n7514 ; n7748
g7493 and n7510_not n7748 ; n7749
g7494 and n7511_not n7514_not ; n7750
g7495 and n7749_not n7750_not ; n7751
g7496 and n432 n7751_not ; n7752
g7497 and n7601_not n7752 ; n7753
g7498 and n7747_not n7753_not ; n7754
g7499 and b[15]_not n7754_not ; n7755
g7500 and n7332_not quotient[32]_not ; n7756
g7501 and n7342_not n7509 ; n7757
g7502 and n7505_not n7757 ; n7758
g7503 and n7506_not n7509_not ; n7759
g7504 and n7758_not n7759_not ; n7760
g7505 and n432 n7760_not ; n7761
g7506 and n7601_not n7761 ; n7762
g7507 and n7756_not n7762_not ; n7763
g7508 and b[14]_not n7763_not ; n7764
g7509 and n7341_not quotient[32]_not ; n7765
g7510 and n7351_not n7504 ; n7766
g7511 and n7500_not n7766 ; n7767
g7512 and n7501_not n7504_not ; n7768
g7513 and n7767_not n7768_not ; n7769
g7514 and n432 n7769_not ; n7770
g7515 and n7601_not n7770 ; n7771
g7516 and n7765_not n7771_not ; n7772
g7517 and b[13]_not n7772_not ; n7773
g7518 and n7350_not quotient[32]_not ; n7774
g7519 and n7360_not n7499 ; n7775
g7520 and n7495_not n7775 ; n7776
g7521 and n7496_not n7499_not ; n7777
g7522 and n7776_not n7777_not ; n7778
g7523 and n432 n7778_not ; n7779
g7524 and n7601_not n7779 ; n7780
g7525 and n7774_not n7780_not ; n7781
g7526 and b[12]_not n7781_not ; n7782
g7527 and n7359_not quotient[32]_not ; n7783
g7528 and n7369_not n7494 ; n7784
g7529 and n7490_not n7784 ; n7785
g7530 and n7491_not n7494_not ; n7786
g7531 and n7785_not n7786_not ; n7787
g7532 and n432 n7787_not ; n7788
g7533 and n7601_not n7788 ; n7789
g7534 and n7783_not n7789_not ; n7790
g7535 and b[11]_not n7790_not ; n7791
g7536 and n7368_not quotient[32]_not ; n7792
g7537 and n7378_not n7489 ; n7793
g7538 and n7485_not n7793 ; n7794
g7539 and n7486_not n7489_not ; n7795
g7540 and n7794_not n7795_not ; n7796
g7541 and n432 n7796_not ; n7797
g7542 and n7601_not n7797 ; n7798
g7543 and n7792_not n7798_not ; n7799
g7544 and b[10]_not n7799_not ; n7800
g7545 and n7377_not quotient[32]_not ; n7801
g7546 and n7387_not n7484 ; n7802
g7547 and n7480_not n7802 ; n7803
g7548 and n7481_not n7484_not ; n7804
g7549 and n7803_not n7804_not ; n7805
g7550 and n432 n7805_not ; n7806
g7551 and n7601_not n7806 ; n7807
g7552 and n7801_not n7807_not ; n7808
g7553 and b[9]_not n7808_not ; n7809
g7554 and n7386_not quotient[32]_not ; n7810
g7555 and n7396_not n7479 ; n7811
g7556 and n7475_not n7811 ; n7812
g7557 and n7476_not n7479_not ; n7813
g7558 and n7812_not n7813_not ; n7814
g7559 and n432 n7814_not ; n7815
g7560 and n7601_not n7815 ; n7816
g7561 and n7810_not n7816_not ; n7817
g7562 and b[8]_not n7817_not ; n7818
g7563 and n7395_not quotient[32]_not ; n7819
g7564 and n7405_not n7474 ; n7820
g7565 and n7470_not n7820 ; n7821
g7566 and n7471_not n7474_not ; n7822
g7567 and n7821_not n7822_not ; n7823
g7568 and n432 n7823_not ; n7824
g7569 and n7601_not n7824 ; n7825
g7570 and n7819_not n7825_not ; n7826
g7571 and b[7]_not n7826_not ; n7827
g7572 and n7404_not quotient[32]_not ; n7828
g7573 and n7414_not n7469 ; n7829
g7574 and n7465_not n7829 ; n7830
g7575 and n7466_not n7469_not ; n7831
g7576 and n7830_not n7831_not ; n7832
g7577 and n432 n7832_not ; n7833
g7578 and n7601_not n7833 ; n7834
g7579 and n7828_not n7834_not ; n7835
g7580 and b[6]_not n7835_not ; n7836
g7581 and n7413_not quotient[32]_not ; n7837
g7582 and n7423_not n7464 ; n7838
g7583 and n7460_not n7838 ; n7839
g7584 and n7461_not n7464_not ; n7840
g7585 and n7839_not n7840_not ; n7841
g7586 and n432 n7841_not ; n7842
g7587 and n7601_not n7842 ; n7843
g7588 and n7837_not n7843_not ; n7844
g7589 and b[5]_not n7844_not ; n7845
g7590 and n7422_not quotient[32]_not ; n7846
g7591 and n7431_not n7459 ; n7847
g7592 and n7455_not n7847 ; n7848
g7593 and n7456_not n7459_not ; n7849
g7594 and n7848_not n7849_not ; n7850
g7595 and n432 n7850_not ; n7851
g7596 and n7601_not n7851 ; n7852
g7597 and n7846_not n7852_not ; n7853
g7598 and b[4]_not n7853_not ; n7854
g7599 and n7430_not quotient[32]_not ; n7855
g7600 and n7450_not n7454 ; n7856
g7601 and n7449_not n7856 ; n7857
g7602 and n7451_not n7454_not ; n7858
g7603 and n7857_not n7858_not ; n7859
g7604 and n432 n7859_not ; n7860
g7605 and n7601_not n7860 ; n7861
g7606 and n7855_not n7861_not ; n7862
g7607 and b[3]_not n7862_not ; n7863
g7608 and n7443_not quotient[32]_not ; n7864
g7609 and n7446_not n7448 ; n7865
g7610 and n7444_not n7865 ; n7866
g7611 and n432 n7866_not ; n7867
g7612 and n7449_not n7867 ; n7868
g7613 and n7601_not n7868 ; n7869
g7614 and n7864_not n7869_not ; n7870
g7615 and b[2]_not n7870_not ; n7871
g7616 and b[0] b[32]_not ; n7872
g7617 and n414 n7872 ; n7873
g7618 and n598 n7873 ; n7874
g7619 and n595 n7874 ; n7875
g7620 and n7601_not n7875 ; n7876
g7621 and a[32] n7876_not ; n7877
g7622 and n313 n7448 ; n7878
g7623 and n303 n7878 ; n7879
g7624 and n288 n7879 ; n7880
g7625 and n7601_not n7880 ; n7881
g7626 and n7877_not n7881_not ; n7882
g7627 and b[1] n7882_not ; n7883
g7628 and b[1]_not n7881_not ; n7884
g7629 and n7877_not n7884 ; n7885
g7630 and n7883_not n7885_not ; n7886
g7631 and a[31]_not b[0] ; n7887
g7632 and n7886_not n7887_not ; n7888
g7633 and b[1]_not n7882_not ; n7889
g7634 and n7888_not n7889_not ; n7890
g7635 and b[2] n7869_not ; n7891
g7636 and n7864_not n7891 ; n7892
g7637 and n7871_not n7892_not ; n7893
g7638 and n7890_not n7893 ; n7894
g7639 and n7871_not n7894_not ; n7895
g7640 and b[3] n7861_not ; n7896
g7641 and n7855_not n7896 ; n7897
g7642 and n7863_not n7897_not ; n7898
g7643 and n7895_not n7898 ; n7899
g7644 and n7863_not n7899_not ; n7900
g7645 and b[4] n7852_not ; n7901
g7646 and n7846_not n7901 ; n7902
g7647 and n7854_not n7902_not ; n7903
g7648 and n7900_not n7903 ; n7904
g7649 and n7854_not n7904_not ; n7905
g7650 and b[5] n7843_not ; n7906
g7651 and n7837_not n7906 ; n7907
g7652 and n7845_not n7907_not ; n7908
g7653 and n7905_not n7908 ; n7909
g7654 and n7845_not n7909_not ; n7910
g7655 and b[6] n7834_not ; n7911
g7656 and n7828_not n7911 ; n7912
g7657 and n7836_not n7912_not ; n7913
g7658 and n7910_not n7913 ; n7914
g7659 and n7836_not n7914_not ; n7915
g7660 and b[7] n7825_not ; n7916
g7661 and n7819_not n7916 ; n7917
g7662 and n7827_not n7917_not ; n7918
g7663 and n7915_not n7918 ; n7919
g7664 and n7827_not n7919_not ; n7920
g7665 and b[8] n7816_not ; n7921
g7666 and n7810_not n7921 ; n7922
g7667 and n7818_not n7922_not ; n7923
g7668 and n7920_not n7923 ; n7924
g7669 and n7818_not n7924_not ; n7925
g7670 and b[9] n7807_not ; n7926
g7671 and n7801_not n7926 ; n7927
g7672 and n7809_not n7927_not ; n7928
g7673 and n7925_not n7928 ; n7929
g7674 and n7809_not n7929_not ; n7930
g7675 and b[10] n7798_not ; n7931
g7676 and n7792_not n7931 ; n7932
g7677 and n7800_not n7932_not ; n7933
g7678 and n7930_not n7933 ; n7934
g7679 and n7800_not n7934_not ; n7935
g7680 and b[11] n7789_not ; n7936
g7681 and n7783_not n7936 ; n7937
g7682 and n7791_not n7937_not ; n7938
g7683 and n7935_not n7938 ; n7939
g7684 and n7791_not n7939_not ; n7940
g7685 and b[12] n7780_not ; n7941
g7686 and n7774_not n7941 ; n7942
g7687 and n7782_not n7942_not ; n7943
g7688 and n7940_not n7943 ; n7944
g7689 and n7782_not n7944_not ; n7945
g7690 and b[13] n7771_not ; n7946
g7691 and n7765_not n7946 ; n7947
g7692 and n7773_not n7947_not ; n7948
g7693 and n7945_not n7948 ; n7949
g7694 and n7773_not n7949_not ; n7950
g7695 and b[14] n7762_not ; n7951
g7696 and n7756_not n7951 ; n7952
g7697 and n7764_not n7952_not ; n7953
g7698 and n7950_not n7953 ; n7954
g7699 and n7764_not n7954_not ; n7955
g7700 and b[15] n7753_not ; n7956
g7701 and n7747_not n7956 ; n7957
g7702 and n7755_not n7957_not ; n7958
g7703 and n7955_not n7958 ; n7959
g7704 and n7755_not n7959_not ; n7960
g7705 and b[16] n7744_not ; n7961
g7706 and n7738_not n7961 ; n7962
g7707 and n7746_not n7962_not ; n7963
g7708 and n7960_not n7963 ; n7964
g7709 and n7746_not n7964_not ; n7965
g7710 and b[17] n7735_not ; n7966
g7711 and n7729_not n7966 ; n7967
g7712 and n7737_not n7967_not ; n7968
g7713 and n7965_not n7968 ; n7969
g7714 and n7737_not n7969_not ; n7970
g7715 and b[18] n7726_not ; n7971
g7716 and n7720_not n7971 ; n7972
g7717 and n7728_not n7972_not ; n7973
g7718 and n7970_not n7973 ; n7974
g7719 and n7728_not n7974_not ; n7975
g7720 and b[19] n7717_not ; n7976
g7721 and n7711_not n7976 ; n7977
g7722 and n7719_not n7977_not ; n7978
g7723 and n7975_not n7978 ; n7979
g7724 and n7719_not n7979_not ; n7980
g7725 and b[20] n7708_not ; n7981
g7726 and n7702_not n7981 ; n7982
g7727 and n7710_not n7982_not ; n7983
g7728 and n7980_not n7983 ; n7984
g7729 and n7710_not n7984_not ; n7985
g7730 and b[21] n7699_not ; n7986
g7731 and n7693_not n7986 ; n7987
g7732 and n7701_not n7987_not ; n7988
g7733 and n7985_not n7988 ; n7989
g7734 and n7701_not n7989_not ; n7990
g7735 and b[22] n7690_not ; n7991
g7736 and n7684_not n7991 ; n7992
g7737 and n7692_not n7992_not ; n7993
g7738 and n7990_not n7993 ; n7994
g7739 and n7692_not n7994_not ; n7995
g7740 and b[23] n7681_not ; n7996
g7741 and n7675_not n7996 ; n7997
g7742 and n7683_not n7997_not ; n7998
g7743 and n7995_not n7998 ; n7999
g7744 and n7683_not n7999_not ; n8000
g7745 and b[24] n7672_not ; n8001
g7746 and n7666_not n8001 ; n8002
g7747 and n7674_not n8002_not ; n8003
g7748 and n8000_not n8003 ; n8004
g7749 and n7674_not n8004_not ; n8005
g7750 and b[25] n7663_not ; n8006
g7751 and n7657_not n8006 ; n8007
g7752 and n7665_not n8007_not ; n8008
g7753 and n8005_not n8008 ; n8009
g7754 and n7665_not n8009_not ; n8010
g7755 and b[26] n7654_not ; n8011
g7756 and n7648_not n8011 ; n8012
g7757 and n7656_not n8012_not ; n8013
g7758 and n8010_not n8013 ; n8014
g7759 and n7656_not n8014_not ; n8015
g7760 and b[27] n7645_not ; n8016
g7761 and n7639_not n8016 ; n8017
g7762 and n7647_not n8017_not ; n8018
g7763 and n8015_not n8018 ; n8019
g7764 and n7647_not n8019_not ; n8020
g7765 and b[28] n7636_not ; n8021
g7766 and n7630_not n8021 ; n8022
g7767 and n7638_not n8022_not ; n8023
g7768 and n8020_not n8023 ; n8024
g7769 and n7638_not n8024_not ; n8025
g7770 and b[29] n7627_not ; n8026
g7771 and n7621_not n8026 ; n8027
g7772 and n7629_not n8027_not ; n8028
g7773 and n8025_not n8028 ; n8029
g7774 and n7629_not n8029_not ; n8030
g7775 and b[30] n7618_not ; n8031
g7776 and n7612_not n8031 ; n8032
g7777 and n7620_not n8032_not ; n8033
g7778 and n8030_not n8033 ; n8034
g7779 and n7620_not n8034_not ; n8035
g7780 and b[31] n7609_not ; n8036
g7781 and n7603_not n8036 ; n8037
g7782 and n7611_not n8037_not ; n8038
g7783 and n8035_not n8038 ; n8039
g7784 and n7611_not n8039_not ; n8040
g7785 and n7178_not quotient[32]_not ; n8041
g7786 and n7180_not n7599 ; n8042
g7787 and n7595_not n8042 ; n8043
g7788 and n7596_not n7599_not ; n8044
g7789 and n8043_not n8044_not ; n8045
g7790 and quotient[32] n8045_not ; n8046
g7791 and n8041_not n8046_not ; n8047
g7792 and b[32]_not n8047_not ; n8048
g7793 and b[32] n8041_not ; n8049
g7794 and n8046_not n8049 ; n8050
g7795 and n424 n8050_not ; n8051
g7796 and n8048_not n8051 ; n8052
g7797 and n8040_not n8052 ; n8053
g7798 and n432 n8047_not ; n8054
g7799 and n8053_not n8054_not ; quotient[31]
g7800 and n7620_not n8038 ; n8056
g7801 and n8034_not n8056 ; n8057
g7802 and n8035_not n8038_not ; n8058
g7803 and n8057_not n8058_not ; n8059
g7804 and quotient[31] n8059_not ; n8060
g7805 and n7610_not n8054_not ; n8061
g7806 and n8053_not n8061 ; n8062
g7807 and n8060_not n8062_not ; n8063
g7808 and n7611_not n8050_not ; n8064
g7809 and n8048_not n8064 ; n8065
g7810 and n8039_not n8065 ; n8066
g7811 and n8048_not n8050_not ; n8067
g7812 and n8040_not n8067_not ; n8068
g7813 and n8066_not n8068_not ; n8069
g7814 and quotient[31] n8069_not ; n8070
g7815 and n8047_not n8054_not ; n8071
g7816 and n8053_not n8071 ; n8072
g7817 and n8070_not n8072_not ; n8073
g7818 and b[33]_not n8073_not ; n8074
g7819 and b[32]_not n8063_not ; n8075
g7820 and n7629_not n8033 ; n8076
g7821 and n8029_not n8076 ; n8077
g7822 and n8030_not n8033_not ; n8078
g7823 and n8077_not n8078_not ; n8079
g7824 and quotient[31] n8079_not ; n8080
g7825 and n7619_not n8054_not ; n8081
g7826 and n8053_not n8081 ; n8082
g7827 and n8080_not n8082_not ; n8083
g7828 and b[31]_not n8083_not ; n8084
g7829 and n7638_not n8028 ; n8085
g7830 and n8024_not n8085 ; n8086
g7831 and n8025_not n8028_not ; n8087
g7832 and n8086_not n8087_not ; n8088
g7833 and quotient[31] n8088_not ; n8089
g7834 and n7628_not n8054_not ; n8090
g7835 and n8053_not n8090 ; n8091
g7836 and n8089_not n8091_not ; n8092
g7837 and b[30]_not n8092_not ; n8093
g7838 and n7647_not n8023 ; n8094
g7839 and n8019_not n8094 ; n8095
g7840 and n8020_not n8023_not ; n8096
g7841 and n8095_not n8096_not ; n8097
g7842 and quotient[31] n8097_not ; n8098
g7843 and n7637_not n8054_not ; n8099
g7844 and n8053_not n8099 ; n8100
g7845 and n8098_not n8100_not ; n8101
g7846 and b[29]_not n8101_not ; n8102
g7847 and n7656_not n8018 ; n8103
g7848 and n8014_not n8103 ; n8104
g7849 and n8015_not n8018_not ; n8105
g7850 and n8104_not n8105_not ; n8106
g7851 and quotient[31] n8106_not ; n8107
g7852 and n7646_not n8054_not ; n8108
g7853 and n8053_not n8108 ; n8109
g7854 and n8107_not n8109_not ; n8110
g7855 and b[28]_not n8110_not ; n8111
g7856 and n7665_not n8013 ; n8112
g7857 and n8009_not n8112 ; n8113
g7858 and n8010_not n8013_not ; n8114
g7859 and n8113_not n8114_not ; n8115
g7860 and quotient[31] n8115_not ; n8116
g7861 and n7655_not n8054_not ; n8117
g7862 and n8053_not n8117 ; n8118
g7863 and n8116_not n8118_not ; n8119
g7864 and b[27]_not n8119_not ; n8120
g7865 and n7674_not n8008 ; n8121
g7866 and n8004_not n8121 ; n8122
g7867 and n8005_not n8008_not ; n8123
g7868 and n8122_not n8123_not ; n8124
g7869 and quotient[31] n8124_not ; n8125
g7870 and n7664_not n8054_not ; n8126
g7871 and n8053_not n8126 ; n8127
g7872 and n8125_not n8127_not ; n8128
g7873 and b[26]_not n8128_not ; n8129
g7874 and n7683_not n8003 ; n8130
g7875 and n7999_not n8130 ; n8131
g7876 and n8000_not n8003_not ; n8132
g7877 and n8131_not n8132_not ; n8133
g7878 and quotient[31] n8133_not ; n8134
g7879 and n7673_not n8054_not ; n8135
g7880 and n8053_not n8135 ; n8136
g7881 and n8134_not n8136_not ; n8137
g7882 and b[25]_not n8137_not ; n8138
g7883 and n7692_not n7998 ; n8139
g7884 and n7994_not n8139 ; n8140
g7885 and n7995_not n7998_not ; n8141
g7886 and n8140_not n8141_not ; n8142
g7887 and quotient[31] n8142_not ; n8143
g7888 and n7682_not n8054_not ; n8144
g7889 and n8053_not n8144 ; n8145
g7890 and n8143_not n8145_not ; n8146
g7891 and b[24]_not n8146_not ; n8147
g7892 and n7701_not n7993 ; n8148
g7893 and n7989_not n8148 ; n8149
g7894 and n7990_not n7993_not ; n8150
g7895 and n8149_not n8150_not ; n8151
g7896 and quotient[31] n8151_not ; n8152
g7897 and n7691_not n8054_not ; n8153
g7898 and n8053_not n8153 ; n8154
g7899 and n8152_not n8154_not ; n8155
g7900 and b[23]_not n8155_not ; n8156
g7901 and n7710_not n7988 ; n8157
g7902 and n7984_not n8157 ; n8158
g7903 and n7985_not n7988_not ; n8159
g7904 and n8158_not n8159_not ; n8160
g7905 and quotient[31] n8160_not ; n8161
g7906 and n7700_not n8054_not ; n8162
g7907 and n8053_not n8162 ; n8163
g7908 and n8161_not n8163_not ; n8164
g7909 and b[22]_not n8164_not ; n8165
g7910 and n7719_not n7983 ; n8166
g7911 and n7979_not n8166 ; n8167
g7912 and n7980_not n7983_not ; n8168
g7913 and n8167_not n8168_not ; n8169
g7914 and quotient[31] n8169_not ; n8170
g7915 and n7709_not n8054_not ; n8171
g7916 and n8053_not n8171 ; n8172
g7917 and n8170_not n8172_not ; n8173
g7918 and b[21]_not n8173_not ; n8174
g7919 and n7728_not n7978 ; n8175
g7920 and n7974_not n8175 ; n8176
g7921 and n7975_not n7978_not ; n8177
g7922 and n8176_not n8177_not ; n8178
g7923 and quotient[31] n8178_not ; n8179
g7924 and n7718_not n8054_not ; n8180
g7925 and n8053_not n8180 ; n8181
g7926 and n8179_not n8181_not ; n8182
g7927 and b[20]_not n8182_not ; n8183
g7928 and n7737_not n7973 ; n8184
g7929 and n7969_not n8184 ; n8185
g7930 and n7970_not n7973_not ; n8186
g7931 and n8185_not n8186_not ; n8187
g7932 and quotient[31] n8187_not ; n8188
g7933 and n7727_not n8054_not ; n8189
g7934 and n8053_not n8189 ; n8190
g7935 and n8188_not n8190_not ; n8191
g7936 and b[19]_not n8191_not ; n8192
g7937 and n7746_not n7968 ; n8193
g7938 and n7964_not n8193 ; n8194
g7939 and n7965_not n7968_not ; n8195
g7940 and n8194_not n8195_not ; n8196
g7941 and quotient[31] n8196_not ; n8197
g7942 and n7736_not n8054_not ; n8198
g7943 and n8053_not n8198 ; n8199
g7944 and n8197_not n8199_not ; n8200
g7945 and b[18]_not n8200_not ; n8201
g7946 and n7755_not n7963 ; n8202
g7947 and n7959_not n8202 ; n8203
g7948 and n7960_not n7963_not ; n8204
g7949 and n8203_not n8204_not ; n8205
g7950 and quotient[31] n8205_not ; n8206
g7951 and n7745_not n8054_not ; n8207
g7952 and n8053_not n8207 ; n8208
g7953 and n8206_not n8208_not ; n8209
g7954 and b[17]_not n8209_not ; n8210
g7955 and n7764_not n7958 ; n8211
g7956 and n7954_not n8211 ; n8212
g7957 and n7955_not n7958_not ; n8213
g7958 and n8212_not n8213_not ; n8214
g7959 and quotient[31] n8214_not ; n8215
g7960 and n7754_not n8054_not ; n8216
g7961 and n8053_not n8216 ; n8217
g7962 and n8215_not n8217_not ; n8218
g7963 and b[16]_not n8218_not ; n8219
g7964 and n7773_not n7953 ; n8220
g7965 and n7949_not n8220 ; n8221
g7966 and n7950_not n7953_not ; n8222
g7967 and n8221_not n8222_not ; n8223
g7968 and quotient[31] n8223_not ; n8224
g7969 and n7763_not n8054_not ; n8225
g7970 and n8053_not n8225 ; n8226
g7971 and n8224_not n8226_not ; n8227
g7972 and b[15]_not n8227_not ; n8228
g7973 and n7782_not n7948 ; n8229
g7974 and n7944_not n8229 ; n8230
g7975 and n7945_not n7948_not ; n8231
g7976 and n8230_not n8231_not ; n8232
g7977 and quotient[31] n8232_not ; n8233
g7978 and n7772_not n8054_not ; n8234
g7979 and n8053_not n8234 ; n8235
g7980 and n8233_not n8235_not ; n8236
g7981 and b[14]_not n8236_not ; n8237
g7982 and n7791_not n7943 ; n8238
g7983 and n7939_not n8238 ; n8239
g7984 and n7940_not n7943_not ; n8240
g7985 and n8239_not n8240_not ; n8241
g7986 and quotient[31] n8241_not ; n8242
g7987 and n7781_not n8054_not ; n8243
g7988 and n8053_not n8243 ; n8244
g7989 and n8242_not n8244_not ; n8245
g7990 and b[13]_not n8245_not ; n8246
g7991 and n7800_not n7938 ; n8247
g7992 and n7934_not n8247 ; n8248
g7993 and n7935_not n7938_not ; n8249
g7994 and n8248_not n8249_not ; n8250
g7995 and quotient[31] n8250_not ; n8251
g7996 and n7790_not n8054_not ; n8252
g7997 and n8053_not n8252 ; n8253
g7998 and n8251_not n8253_not ; n8254
g7999 and b[12]_not n8254_not ; n8255
g8000 and n7809_not n7933 ; n8256
g8001 and n7929_not n8256 ; n8257
g8002 and n7930_not n7933_not ; n8258
g8003 and n8257_not n8258_not ; n8259
g8004 and quotient[31] n8259_not ; n8260
g8005 and n7799_not n8054_not ; n8261
g8006 and n8053_not n8261 ; n8262
g8007 and n8260_not n8262_not ; n8263
g8008 and b[11]_not n8263_not ; n8264
g8009 and n7818_not n7928 ; n8265
g8010 and n7924_not n8265 ; n8266
g8011 and n7925_not n7928_not ; n8267
g8012 and n8266_not n8267_not ; n8268
g8013 and quotient[31] n8268_not ; n8269
g8014 and n7808_not n8054_not ; n8270
g8015 and n8053_not n8270 ; n8271
g8016 and n8269_not n8271_not ; n8272
g8017 and b[10]_not n8272_not ; n8273
g8018 and n7827_not n7923 ; n8274
g8019 and n7919_not n8274 ; n8275
g8020 and n7920_not n7923_not ; n8276
g8021 and n8275_not n8276_not ; n8277
g8022 and quotient[31] n8277_not ; n8278
g8023 and n7817_not n8054_not ; n8279
g8024 and n8053_not n8279 ; n8280
g8025 and n8278_not n8280_not ; n8281
g8026 and b[9]_not n8281_not ; n8282
g8027 and n7836_not n7918 ; n8283
g8028 and n7914_not n8283 ; n8284
g8029 and n7915_not n7918_not ; n8285
g8030 and n8284_not n8285_not ; n8286
g8031 and quotient[31] n8286_not ; n8287
g8032 and n7826_not n8054_not ; n8288
g8033 and n8053_not n8288 ; n8289
g8034 and n8287_not n8289_not ; n8290
g8035 and b[8]_not n8290_not ; n8291
g8036 and n7845_not n7913 ; n8292
g8037 and n7909_not n8292 ; n8293
g8038 and n7910_not n7913_not ; n8294
g8039 and n8293_not n8294_not ; n8295
g8040 and quotient[31] n8295_not ; n8296
g8041 and n7835_not n8054_not ; n8297
g8042 and n8053_not n8297 ; n8298
g8043 and n8296_not n8298_not ; n8299
g8044 and b[7]_not n8299_not ; n8300
g8045 and n7854_not n7908 ; n8301
g8046 and n7904_not n8301 ; n8302
g8047 and n7905_not n7908_not ; n8303
g8048 and n8302_not n8303_not ; n8304
g8049 and quotient[31] n8304_not ; n8305
g8050 and n7844_not n8054_not ; n8306
g8051 and n8053_not n8306 ; n8307
g8052 and n8305_not n8307_not ; n8308
g8053 and b[6]_not n8308_not ; n8309
g8054 and n7863_not n7903 ; n8310
g8055 and n7899_not n8310 ; n8311
g8056 and n7900_not n7903_not ; n8312
g8057 and n8311_not n8312_not ; n8313
g8058 and quotient[31] n8313_not ; n8314
g8059 and n7853_not n8054_not ; n8315
g8060 and n8053_not n8315 ; n8316
g8061 and n8314_not n8316_not ; n8317
g8062 and b[5]_not n8317_not ; n8318
g8063 and n7871_not n7898 ; n8319
g8064 and n7894_not n8319 ; n8320
g8065 and n7895_not n7898_not ; n8321
g8066 and n8320_not n8321_not ; n8322
g8067 and quotient[31] n8322_not ; n8323
g8068 and n7862_not n8054_not ; n8324
g8069 and n8053_not n8324 ; n8325
g8070 and n8323_not n8325_not ; n8326
g8071 and b[4]_not n8326_not ; n8327
g8072 and n7889_not n7893 ; n8328
g8073 and n7888_not n8328 ; n8329
g8074 and n7890_not n7893_not ; n8330
g8075 and n8329_not n8330_not ; n8331
g8076 and quotient[31] n8331_not ; n8332
g8077 and n7870_not n8054_not ; n8333
g8078 and n8053_not n8333 ; n8334
g8079 and n8332_not n8334_not ; n8335
g8080 and b[3]_not n8335_not ; n8336
g8081 and n7885_not n7887 ; n8337
g8082 and n7883_not n8337 ; n8338
g8083 and n7888_not n8338_not ; n8339
g8084 and quotient[31] n8339 ; n8340
g8085 and n7882_not n8054_not ; n8341
g8086 and n8053_not n8341 ; n8342
g8087 and n8340_not n8342_not ; n8343
g8088 and b[2]_not n8343_not ; n8344
g8089 and b[0] quotient[31] ; n8345
g8090 and a[31] n8345_not ; n8346
g8091 and n7887 quotient[31] ; n8347
g8092 and n8346_not n8347_not ; n8348
g8093 and b[1] n8348_not ; n8349
g8094 and b[1]_not n8347_not ; n8350
g8095 and n8346_not n8350 ; n8351
g8096 and n8349_not n8351_not ; n8352
g8097 and a[30]_not b[0] ; n8353
g8098 and n8352_not n8353_not ; n8354
g8099 and b[1]_not n8348_not ; n8355
g8100 and n8354_not n8355_not ; n8356
g8101 and b[2] n8342_not ; n8357
g8102 and n8340_not n8357 ; n8358
g8103 and n8344_not n8358_not ; n8359
g8104 and n8356_not n8359 ; n8360
g8105 and n8344_not n8360_not ; n8361
g8106 and b[3] n8334_not ; n8362
g8107 and n8332_not n8362 ; n8363
g8108 and n8336_not n8363_not ; n8364
g8109 and n8361_not n8364 ; n8365
g8110 and n8336_not n8365_not ; n8366
g8111 and b[4] n8325_not ; n8367
g8112 and n8323_not n8367 ; n8368
g8113 and n8327_not n8368_not ; n8369
g8114 and n8366_not n8369 ; n8370
g8115 and n8327_not n8370_not ; n8371
g8116 and b[5] n8316_not ; n8372
g8117 and n8314_not n8372 ; n8373
g8118 and n8318_not n8373_not ; n8374
g8119 and n8371_not n8374 ; n8375
g8120 and n8318_not n8375_not ; n8376
g8121 and b[6] n8307_not ; n8377
g8122 and n8305_not n8377 ; n8378
g8123 and n8309_not n8378_not ; n8379
g8124 and n8376_not n8379 ; n8380
g8125 and n8309_not n8380_not ; n8381
g8126 and b[7] n8298_not ; n8382
g8127 and n8296_not n8382 ; n8383
g8128 and n8300_not n8383_not ; n8384
g8129 and n8381_not n8384 ; n8385
g8130 and n8300_not n8385_not ; n8386
g8131 and b[8] n8289_not ; n8387
g8132 and n8287_not n8387 ; n8388
g8133 and n8291_not n8388_not ; n8389
g8134 and n8386_not n8389 ; n8390
g8135 and n8291_not n8390_not ; n8391
g8136 and b[9] n8280_not ; n8392
g8137 and n8278_not n8392 ; n8393
g8138 and n8282_not n8393_not ; n8394
g8139 and n8391_not n8394 ; n8395
g8140 and n8282_not n8395_not ; n8396
g8141 and b[10] n8271_not ; n8397
g8142 and n8269_not n8397 ; n8398
g8143 and n8273_not n8398_not ; n8399
g8144 and n8396_not n8399 ; n8400
g8145 and n8273_not n8400_not ; n8401
g8146 and b[11] n8262_not ; n8402
g8147 and n8260_not n8402 ; n8403
g8148 and n8264_not n8403_not ; n8404
g8149 and n8401_not n8404 ; n8405
g8150 and n8264_not n8405_not ; n8406
g8151 and b[12] n8253_not ; n8407
g8152 and n8251_not n8407 ; n8408
g8153 and n8255_not n8408_not ; n8409
g8154 and n8406_not n8409 ; n8410
g8155 and n8255_not n8410_not ; n8411
g8156 and b[13] n8244_not ; n8412
g8157 and n8242_not n8412 ; n8413
g8158 and n8246_not n8413_not ; n8414
g8159 and n8411_not n8414 ; n8415
g8160 and n8246_not n8415_not ; n8416
g8161 and b[14] n8235_not ; n8417
g8162 and n8233_not n8417 ; n8418
g8163 and n8237_not n8418_not ; n8419
g8164 and n8416_not n8419 ; n8420
g8165 and n8237_not n8420_not ; n8421
g8166 and b[15] n8226_not ; n8422
g8167 and n8224_not n8422 ; n8423
g8168 and n8228_not n8423_not ; n8424
g8169 and n8421_not n8424 ; n8425
g8170 and n8228_not n8425_not ; n8426
g8171 and b[16] n8217_not ; n8427
g8172 and n8215_not n8427 ; n8428
g8173 and n8219_not n8428_not ; n8429
g8174 and n8426_not n8429 ; n8430
g8175 and n8219_not n8430_not ; n8431
g8176 and b[17] n8208_not ; n8432
g8177 and n8206_not n8432 ; n8433
g8178 and n8210_not n8433_not ; n8434
g8179 and n8431_not n8434 ; n8435
g8180 and n8210_not n8435_not ; n8436
g8181 and b[18] n8199_not ; n8437
g8182 and n8197_not n8437 ; n8438
g8183 and n8201_not n8438_not ; n8439
g8184 and n8436_not n8439 ; n8440
g8185 and n8201_not n8440_not ; n8441
g8186 and b[19] n8190_not ; n8442
g8187 and n8188_not n8442 ; n8443
g8188 and n8192_not n8443_not ; n8444
g8189 and n8441_not n8444 ; n8445
g8190 and n8192_not n8445_not ; n8446
g8191 and b[20] n8181_not ; n8447
g8192 and n8179_not n8447 ; n8448
g8193 and n8183_not n8448_not ; n8449
g8194 and n8446_not n8449 ; n8450
g8195 and n8183_not n8450_not ; n8451
g8196 and b[21] n8172_not ; n8452
g8197 and n8170_not n8452 ; n8453
g8198 and n8174_not n8453_not ; n8454
g8199 and n8451_not n8454 ; n8455
g8200 and n8174_not n8455_not ; n8456
g8201 and b[22] n8163_not ; n8457
g8202 and n8161_not n8457 ; n8458
g8203 and n8165_not n8458_not ; n8459
g8204 and n8456_not n8459 ; n8460
g8205 and n8165_not n8460_not ; n8461
g8206 and b[23] n8154_not ; n8462
g8207 and n8152_not n8462 ; n8463
g8208 and n8156_not n8463_not ; n8464
g8209 and n8461_not n8464 ; n8465
g8210 and n8156_not n8465_not ; n8466
g8211 and b[24] n8145_not ; n8467
g8212 and n8143_not n8467 ; n8468
g8213 and n8147_not n8468_not ; n8469
g8214 and n8466_not n8469 ; n8470
g8215 and n8147_not n8470_not ; n8471
g8216 and b[25] n8136_not ; n8472
g8217 and n8134_not n8472 ; n8473
g8218 and n8138_not n8473_not ; n8474
g8219 and n8471_not n8474 ; n8475
g8220 and n8138_not n8475_not ; n8476
g8221 and b[26] n8127_not ; n8477
g8222 and n8125_not n8477 ; n8478
g8223 and n8129_not n8478_not ; n8479
g8224 and n8476_not n8479 ; n8480
g8225 and n8129_not n8480_not ; n8481
g8226 and b[27] n8118_not ; n8482
g8227 and n8116_not n8482 ; n8483
g8228 and n8120_not n8483_not ; n8484
g8229 and n8481_not n8484 ; n8485
g8230 and n8120_not n8485_not ; n8486
g8231 and b[28] n8109_not ; n8487
g8232 and n8107_not n8487 ; n8488
g8233 and n8111_not n8488_not ; n8489
g8234 and n8486_not n8489 ; n8490
g8235 and n8111_not n8490_not ; n8491
g8236 and b[29] n8100_not ; n8492
g8237 and n8098_not n8492 ; n8493
g8238 and n8102_not n8493_not ; n8494
g8239 and n8491_not n8494 ; n8495
g8240 and n8102_not n8495_not ; n8496
g8241 and b[30] n8091_not ; n8497
g8242 and n8089_not n8497 ; n8498
g8243 and n8093_not n8498_not ; n8499
g8244 and n8496_not n8499 ; n8500
g8245 and n8093_not n8500_not ; n8501
g8246 and b[31] n8082_not ; n8502
g8247 and n8080_not n8502 ; n8503
g8248 and n8084_not n8503_not ; n8504
g8249 and n8501_not n8504 ; n8505
g8250 and n8084_not n8505_not ; n8506
g8251 and b[32] n8062_not ; n8507
g8252 and n8060_not n8507 ; n8508
g8253 and n8075_not n8508_not ; n8509
g8254 and n8506_not n8509 ; n8510
g8255 and n8075_not n8510_not ; n8511
g8256 and b[33] n8072_not ; n8512
g8257 and n8070_not n8512 ; n8513
g8258 and n8074_not n8513_not ; n8514
g8259 and n8511_not n8514 ; n8515
g8260 and n8074_not n8515_not ; n8516
g8261 and n294 n312 ; n8517
g8262 and n340 n8517 ; n8518
g8263 and n338 n8518 ; n8519
g8264 and n8516_not n8519 ; quotient[30]
g8265 and n8063_not quotient[30]_not ; n8521
g8266 and n8084_not n8509 ; n8522
g8267 and n8505_not n8522 ; n8523
g8268 and n8506_not n8509_not ; n8524
g8269 and n8523_not n8524_not ; n8525
g8270 and n8519 n8525_not ; n8526
g8271 and n8516_not n8526 ; n8527
g8272 and n8521_not n8527_not ; n8528
g8273 and n8073_not quotient[30]_not ; n8529
g8274 and n8075_not n8514 ; n8530
g8275 and n8510_not n8530 ; n8531
g8276 and n8511_not n8514_not ; n8532
g8277 and n8531_not n8532_not ; n8533
g8278 and quotient[30] n8533_not ; n8534
g8279 and n8529_not n8534_not ; n8535
g8280 and b[34]_not n8535_not ; n8536
g8281 and b[33]_not n8528_not ; n8537
g8282 and n8083_not quotient[30]_not ; n8538
g8283 and n8093_not n8504 ; n8539
g8284 and n8500_not n8539 ; n8540
g8285 and n8501_not n8504_not ; n8541
g8286 and n8540_not n8541_not ; n8542
g8287 and n8519 n8542_not ; n8543
g8288 and n8516_not n8543 ; n8544
g8289 and n8538_not n8544_not ; n8545
g8290 and b[32]_not n8545_not ; n8546
g8291 and n8092_not quotient[30]_not ; n8547
g8292 and n8102_not n8499 ; n8548
g8293 and n8495_not n8548 ; n8549
g8294 and n8496_not n8499_not ; n8550
g8295 and n8549_not n8550_not ; n8551
g8296 and n8519 n8551_not ; n8552
g8297 and n8516_not n8552 ; n8553
g8298 and n8547_not n8553_not ; n8554
g8299 and b[31]_not n8554_not ; n8555
g8300 and n8101_not quotient[30]_not ; n8556
g8301 and n8111_not n8494 ; n8557
g8302 and n8490_not n8557 ; n8558
g8303 and n8491_not n8494_not ; n8559
g8304 and n8558_not n8559_not ; n8560
g8305 and n8519 n8560_not ; n8561
g8306 and n8516_not n8561 ; n8562
g8307 and n8556_not n8562_not ; n8563
g8308 and b[30]_not n8563_not ; n8564
g8309 and n8110_not quotient[30]_not ; n8565
g8310 and n8120_not n8489 ; n8566
g8311 and n8485_not n8566 ; n8567
g8312 and n8486_not n8489_not ; n8568
g8313 and n8567_not n8568_not ; n8569
g8314 and n8519 n8569_not ; n8570
g8315 and n8516_not n8570 ; n8571
g8316 and n8565_not n8571_not ; n8572
g8317 and b[29]_not n8572_not ; n8573
g8318 and n8119_not quotient[30]_not ; n8574
g8319 and n8129_not n8484 ; n8575
g8320 and n8480_not n8575 ; n8576
g8321 and n8481_not n8484_not ; n8577
g8322 and n8576_not n8577_not ; n8578
g8323 and n8519 n8578_not ; n8579
g8324 and n8516_not n8579 ; n8580
g8325 and n8574_not n8580_not ; n8581
g8326 and b[28]_not n8581_not ; n8582
g8327 and n8128_not quotient[30]_not ; n8583
g8328 and n8138_not n8479 ; n8584
g8329 and n8475_not n8584 ; n8585
g8330 and n8476_not n8479_not ; n8586
g8331 and n8585_not n8586_not ; n8587
g8332 and n8519 n8587_not ; n8588
g8333 and n8516_not n8588 ; n8589
g8334 and n8583_not n8589_not ; n8590
g8335 and b[27]_not n8590_not ; n8591
g8336 and n8137_not quotient[30]_not ; n8592
g8337 and n8147_not n8474 ; n8593
g8338 and n8470_not n8593 ; n8594
g8339 and n8471_not n8474_not ; n8595
g8340 and n8594_not n8595_not ; n8596
g8341 and n8519 n8596_not ; n8597
g8342 and n8516_not n8597 ; n8598
g8343 and n8592_not n8598_not ; n8599
g8344 and b[26]_not n8599_not ; n8600
g8345 and n8146_not quotient[30]_not ; n8601
g8346 and n8156_not n8469 ; n8602
g8347 and n8465_not n8602 ; n8603
g8348 and n8466_not n8469_not ; n8604
g8349 and n8603_not n8604_not ; n8605
g8350 and n8519 n8605_not ; n8606
g8351 and n8516_not n8606 ; n8607
g8352 and n8601_not n8607_not ; n8608
g8353 and b[25]_not n8608_not ; n8609
g8354 and n8155_not quotient[30]_not ; n8610
g8355 and n8165_not n8464 ; n8611
g8356 and n8460_not n8611 ; n8612
g8357 and n8461_not n8464_not ; n8613
g8358 and n8612_not n8613_not ; n8614
g8359 and n8519 n8614_not ; n8615
g8360 and n8516_not n8615 ; n8616
g8361 and n8610_not n8616_not ; n8617
g8362 and b[24]_not n8617_not ; n8618
g8363 and n8164_not quotient[30]_not ; n8619
g8364 and n8174_not n8459 ; n8620
g8365 and n8455_not n8620 ; n8621
g8366 and n8456_not n8459_not ; n8622
g8367 and n8621_not n8622_not ; n8623
g8368 and n8519 n8623_not ; n8624
g8369 and n8516_not n8624 ; n8625
g8370 and n8619_not n8625_not ; n8626
g8371 and b[23]_not n8626_not ; n8627
g8372 and n8173_not quotient[30]_not ; n8628
g8373 and n8183_not n8454 ; n8629
g8374 and n8450_not n8629 ; n8630
g8375 and n8451_not n8454_not ; n8631
g8376 and n8630_not n8631_not ; n8632
g8377 and n8519 n8632_not ; n8633
g8378 and n8516_not n8633 ; n8634
g8379 and n8628_not n8634_not ; n8635
g8380 and b[22]_not n8635_not ; n8636
g8381 and n8182_not quotient[30]_not ; n8637
g8382 and n8192_not n8449 ; n8638
g8383 and n8445_not n8638 ; n8639
g8384 and n8446_not n8449_not ; n8640
g8385 and n8639_not n8640_not ; n8641
g8386 and n8519 n8641_not ; n8642
g8387 and n8516_not n8642 ; n8643
g8388 and n8637_not n8643_not ; n8644
g8389 and b[21]_not n8644_not ; n8645
g8390 and n8191_not quotient[30]_not ; n8646
g8391 and n8201_not n8444 ; n8647
g8392 and n8440_not n8647 ; n8648
g8393 and n8441_not n8444_not ; n8649
g8394 and n8648_not n8649_not ; n8650
g8395 and n8519 n8650_not ; n8651
g8396 and n8516_not n8651 ; n8652
g8397 and n8646_not n8652_not ; n8653
g8398 and b[20]_not n8653_not ; n8654
g8399 and n8200_not quotient[30]_not ; n8655
g8400 and n8210_not n8439 ; n8656
g8401 and n8435_not n8656 ; n8657
g8402 and n8436_not n8439_not ; n8658
g8403 and n8657_not n8658_not ; n8659
g8404 and n8519 n8659_not ; n8660
g8405 and n8516_not n8660 ; n8661
g8406 and n8655_not n8661_not ; n8662
g8407 and b[19]_not n8662_not ; n8663
g8408 and n8209_not quotient[30]_not ; n8664
g8409 and n8219_not n8434 ; n8665
g8410 and n8430_not n8665 ; n8666
g8411 and n8431_not n8434_not ; n8667
g8412 and n8666_not n8667_not ; n8668
g8413 and n8519 n8668_not ; n8669
g8414 and n8516_not n8669 ; n8670
g8415 and n8664_not n8670_not ; n8671
g8416 and b[18]_not n8671_not ; n8672
g8417 and n8218_not quotient[30]_not ; n8673
g8418 and n8228_not n8429 ; n8674
g8419 and n8425_not n8674 ; n8675
g8420 and n8426_not n8429_not ; n8676
g8421 and n8675_not n8676_not ; n8677
g8422 and n8519 n8677_not ; n8678
g8423 and n8516_not n8678 ; n8679
g8424 and n8673_not n8679_not ; n8680
g8425 and b[17]_not n8680_not ; n8681
g8426 and n8227_not quotient[30]_not ; n8682
g8427 and n8237_not n8424 ; n8683
g8428 and n8420_not n8683 ; n8684
g8429 and n8421_not n8424_not ; n8685
g8430 and n8684_not n8685_not ; n8686
g8431 and n8519 n8686_not ; n8687
g8432 and n8516_not n8687 ; n8688
g8433 and n8682_not n8688_not ; n8689
g8434 and b[16]_not n8689_not ; n8690
g8435 and n8236_not quotient[30]_not ; n8691
g8436 and n8246_not n8419 ; n8692
g8437 and n8415_not n8692 ; n8693
g8438 and n8416_not n8419_not ; n8694
g8439 and n8693_not n8694_not ; n8695
g8440 and n8519 n8695_not ; n8696
g8441 and n8516_not n8696 ; n8697
g8442 and n8691_not n8697_not ; n8698
g8443 and b[15]_not n8698_not ; n8699
g8444 and n8245_not quotient[30]_not ; n8700
g8445 and n8255_not n8414 ; n8701
g8446 and n8410_not n8701 ; n8702
g8447 and n8411_not n8414_not ; n8703
g8448 and n8702_not n8703_not ; n8704
g8449 and n8519 n8704_not ; n8705
g8450 and n8516_not n8705 ; n8706
g8451 and n8700_not n8706_not ; n8707
g8452 and b[14]_not n8707_not ; n8708
g8453 and n8254_not quotient[30]_not ; n8709
g8454 and n8264_not n8409 ; n8710
g8455 and n8405_not n8710 ; n8711
g8456 and n8406_not n8409_not ; n8712
g8457 and n8711_not n8712_not ; n8713
g8458 and n8519 n8713_not ; n8714
g8459 and n8516_not n8714 ; n8715
g8460 and n8709_not n8715_not ; n8716
g8461 and b[13]_not n8716_not ; n8717
g8462 and n8263_not quotient[30]_not ; n8718
g8463 and n8273_not n8404 ; n8719
g8464 and n8400_not n8719 ; n8720
g8465 and n8401_not n8404_not ; n8721
g8466 and n8720_not n8721_not ; n8722
g8467 and n8519 n8722_not ; n8723
g8468 and n8516_not n8723 ; n8724
g8469 and n8718_not n8724_not ; n8725
g8470 and b[12]_not n8725_not ; n8726
g8471 and n8272_not quotient[30]_not ; n8727
g8472 and n8282_not n8399 ; n8728
g8473 and n8395_not n8728 ; n8729
g8474 and n8396_not n8399_not ; n8730
g8475 and n8729_not n8730_not ; n8731
g8476 and n8519 n8731_not ; n8732
g8477 and n8516_not n8732 ; n8733
g8478 and n8727_not n8733_not ; n8734
g8479 and b[11]_not n8734_not ; n8735
g8480 and n8281_not quotient[30]_not ; n8736
g8481 and n8291_not n8394 ; n8737
g8482 and n8390_not n8737 ; n8738
g8483 and n8391_not n8394_not ; n8739
g8484 and n8738_not n8739_not ; n8740
g8485 and n8519 n8740_not ; n8741
g8486 and n8516_not n8741 ; n8742
g8487 and n8736_not n8742_not ; n8743
g8488 and b[10]_not n8743_not ; n8744
g8489 and n8290_not quotient[30]_not ; n8745
g8490 and n8300_not n8389 ; n8746
g8491 and n8385_not n8746 ; n8747
g8492 and n8386_not n8389_not ; n8748
g8493 and n8747_not n8748_not ; n8749
g8494 and n8519 n8749_not ; n8750
g8495 and n8516_not n8750 ; n8751
g8496 and n8745_not n8751_not ; n8752
g8497 and b[9]_not n8752_not ; n8753
g8498 and n8299_not quotient[30]_not ; n8754
g8499 and n8309_not n8384 ; n8755
g8500 and n8380_not n8755 ; n8756
g8501 and n8381_not n8384_not ; n8757
g8502 and n8756_not n8757_not ; n8758
g8503 and n8519 n8758_not ; n8759
g8504 and n8516_not n8759 ; n8760
g8505 and n8754_not n8760_not ; n8761
g8506 and b[8]_not n8761_not ; n8762
g8507 and n8308_not quotient[30]_not ; n8763
g8508 and n8318_not n8379 ; n8764
g8509 and n8375_not n8764 ; n8765
g8510 and n8376_not n8379_not ; n8766
g8511 and n8765_not n8766_not ; n8767
g8512 and n8519 n8767_not ; n8768
g8513 and n8516_not n8768 ; n8769
g8514 and n8763_not n8769_not ; n8770
g8515 and b[7]_not n8770_not ; n8771
g8516 and n8317_not quotient[30]_not ; n8772
g8517 and n8327_not n8374 ; n8773
g8518 and n8370_not n8773 ; n8774
g8519 and n8371_not n8374_not ; n8775
g8520 and n8774_not n8775_not ; n8776
g8521 and n8519 n8776_not ; n8777
g8522 and n8516_not n8777 ; n8778
g8523 and n8772_not n8778_not ; n8779
g8524 and b[6]_not n8779_not ; n8780
g8525 and n8326_not quotient[30]_not ; n8781
g8526 and n8336_not n8369 ; n8782
g8527 and n8365_not n8782 ; n8783
g8528 and n8366_not n8369_not ; n8784
g8529 and n8783_not n8784_not ; n8785
g8530 and n8519 n8785_not ; n8786
g8531 and n8516_not n8786 ; n8787
g8532 and n8781_not n8787_not ; n8788
g8533 and b[5]_not n8788_not ; n8789
g8534 and n8335_not quotient[30]_not ; n8790
g8535 and n8344_not n8364 ; n8791
g8536 and n8360_not n8791 ; n8792
g8537 and n8361_not n8364_not ; n8793
g8538 and n8792_not n8793_not ; n8794
g8539 and n8519 n8794_not ; n8795
g8540 and n8516_not n8795 ; n8796
g8541 and n8790_not n8796_not ; n8797
g8542 and b[4]_not n8797_not ; n8798
g8543 and n8343_not quotient[30]_not ; n8799
g8544 and n8355_not n8359 ; n8800
g8545 and n8354_not n8800 ; n8801
g8546 and n8356_not n8359_not ; n8802
g8547 and n8801_not n8802_not ; n8803
g8548 and n8519 n8803_not ; n8804
g8549 and n8516_not n8804 ; n8805
g8550 and n8799_not n8805_not ; n8806
g8551 and b[3]_not n8806_not ; n8807
g8552 and n8348_not quotient[30]_not ; n8808
g8553 and n8351_not n8353 ; n8809
g8554 and n8349_not n8809 ; n8810
g8555 and n8519 n8810_not ; n8811
g8556 and n8354_not n8811 ; n8812
g8557 and n8516_not n8812 ; n8813
g8558 and n8808_not n8813_not ; n8814
g8559 and b[2]_not n8814_not ; n8815
g8560 and b[0] b[34]_not ; n8816
g8561 and n413 n8816 ; n8817
g8562 and n411 n8817 ; n8818
g8563 and n422 n8818 ; n8819
g8564 and n408 n8819 ; n8820
g8565 and n8516_not n8820 ; n8821
g8566 and a[30] n8821_not ; n8822
g8567 and n312 n8353 ; n8823
g8568 and n294 n8823 ; n8824
g8569 and n340 n8824 ; n8825
g8570 and n338 n8825 ; n8826
g8571 and n8516_not n8826 ; n8827
g8572 and n8822_not n8827_not ; n8828
g8573 and b[1] n8828_not ; n8829
g8574 and b[1]_not n8827_not ; n8830
g8575 and n8822_not n8830 ; n8831
g8576 and n8829_not n8831_not ; n8832
g8577 and a[29]_not b[0] ; n8833
g8578 and n8832_not n8833_not ; n8834
g8579 and b[1]_not n8828_not ; n8835
g8580 and n8834_not n8835_not ; n8836
g8581 and b[2] n8813_not ; n8837
g8582 and n8808_not n8837 ; n8838
g8583 and n8815_not n8838_not ; n8839
g8584 and n8836_not n8839 ; n8840
g8585 and n8815_not n8840_not ; n8841
g8586 and b[3] n8805_not ; n8842
g8587 and n8799_not n8842 ; n8843
g8588 and n8807_not n8843_not ; n8844
g8589 and n8841_not n8844 ; n8845
g8590 and n8807_not n8845_not ; n8846
g8591 and b[4] n8796_not ; n8847
g8592 and n8790_not n8847 ; n8848
g8593 and n8798_not n8848_not ; n8849
g8594 and n8846_not n8849 ; n8850
g8595 and n8798_not n8850_not ; n8851
g8596 and b[5] n8787_not ; n8852
g8597 and n8781_not n8852 ; n8853
g8598 and n8789_not n8853_not ; n8854
g8599 and n8851_not n8854 ; n8855
g8600 and n8789_not n8855_not ; n8856
g8601 and b[6] n8778_not ; n8857
g8602 and n8772_not n8857 ; n8858
g8603 and n8780_not n8858_not ; n8859
g8604 and n8856_not n8859 ; n8860
g8605 and n8780_not n8860_not ; n8861
g8606 and b[7] n8769_not ; n8862
g8607 and n8763_not n8862 ; n8863
g8608 and n8771_not n8863_not ; n8864
g8609 and n8861_not n8864 ; n8865
g8610 and n8771_not n8865_not ; n8866
g8611 and b[8] n8760_not ; n8867
g8612 and n8754_not n8867 ; n8868
g8613 and n8762_not n8868_not ; n8869
g8614 and n8866_not n8869 ; n8870
g8615 and n8762_not n8870_not ; n8871
g8616 and b[9] n8751_not ; n8872
g8617 and n8745_not n8872 ; n8873
g8618 and n8753_not n8873_not ; n8874
g8619 and n8871_not n8874 ; n8875
g8620 and n8753_not n8875_not ; n8876
g8621 and b[10] n8742_not ; n8877
g8622 and n8736_not n8877 ; n8878
g8623 and n8744_not n8878_not ; n8879
g8624 and n8876_not n8879 ; n8880
g8625 and n8744_not n8880_not ; n8881
g8626 and b[11] n8733_not ; n8882
g8627 and n8727_not n8882 ; n8883
g8628 and n8735_not n8883_not ; n8884
g8629 and n8881_not n8884 ; n8885
g8630 and n8735_not n8885_not ; n8886
g8631 and b[12] n8724_not ; n8887
g8632 and n8718_not n8887 ; n8888
g8633 and n8726_not n8888_not ; n8889
g8634 and n8886_not n8889 ; n8890
g8635 and n8726_not n8890_not ; n8891
g8636 and b[13] n8715_not ; n8892
g8637 and n8709_not n8892 ; n8893
g8638 and n8717_not n8893_not ; n8894
g8639 and n8891_not n8894 ; n8895
g8640 and n8717_not n8895_not ; n8896
g8641 and b[14] n8706_not ; n8897
g8642 and n8700_not n8897 ; n8898
g8643 and n8708_not n8898_not ; n8899
g8644 and n8896_not n8899 ; n8900
g8645 and n8708_not n8900_not ; n8901
g8646 and b[15] n8697_not ; n8902
g8647 and n8691_not n8902 ; n8903
g8648 and n8699_not n8903_not ; n8904
g8649 and n8901_not n8904 ; n8905
g8650 and n8699_not n8905_not ; n8906
g8651 and b[16] n8688_not ; n8907
g8652 and n8682_not n8907 ; n8908
g8653 and n8690_not n8908_not ; n8909
g8654 and n8906_not n8909 ; n8910
g8655 and n8690_not n8910_not ; n8911
g8656 and b[17] n8679_not ; n8912
g8657 and n8673_not n8912 ; n8913
g8658 and n8681_not n8913_not ; n8914
g8659 and n8911_not n8914 ; n8915
g8660 and n8681_not n8915_not ; n8916
g8661 and b[18] n8670_not ; n8917
g8662 and n8664_not n8917 ; n8918
g8663 and n8672_not n8918_not ; n8919
g8664 and n8916_not n8919 ; n8920
g8665 and n8672_not n8920_not ; n8921
g8666 and b[19] n8661_not ; n8922
g8667 and n8655_not n8922 ; n8923
g8668 and n8663_not n8923_not ; n8924
g8669 and n8921_not n8924 ; n8925
g8670 and n8663_not n8925_not ; n8926
g8671 and b[20] n8652_not ; n8927
g8672 and n8646_not n8927 ; n8928
g8673 and n8654_not n8928_not ; n8929
g8674 and n8926_not n8929 ; n8930
g8675 and n8654_not n8930_not ; n8931
g8676 and b[21] n8643_not ; n8932
g8677 and n8637_not n8932 ; n8933
g8678 and n8645_not n8933_not ; n8934
g8679 and n8931_not n8934 ; n8935
g8680 and n8645_not n8935_not ; n8936
g8681 and b[22] n8634_not ; n8937
g8682 and n8628_not n8937 ; n8938
g8683 and n8636_not n8938_not ; n8939
g8684 and n8936_not n8939 ; n8940
g8685 and n8636_not n8940_not ; n8941
g8686 and b[23] n8625_not ; n8942
g8687 and n8619_not n8942 ; n8943
g8688 and n8627_not n8943_not ; n8944
g8689 and n8941_not n8944 ; n8945
g8690 and n8627_not n8945_not ; n8946
g8691 and b[24] n8616_not ; n8947
g8692 and n8610_not n8947 ; n8948
g8693 and n8618_not n8948_not ; n8949
g8694 and n8946_not n8949 ; n8950
g8695 and n8618_not n8950_not ; n8951
g8696 and b[25] n8607_not ; n8952
g8697 and n8601_not n8952 ; n8953
g8698 and n8609_not n8953_not ; n8954
g8699 and n8951_not n8954 ; n8955
g8700 and n8609_not n8955_not ; n8956
g8701 and b[26] n8598_not ; n8957
g8702 and n8592_not n8957 ; n8958
g8703 and n8600_not n8958_not ; n8959
g8704 and n8956_not n8959 ; n8960
g8705 and n8600_not n8960_not ; n8961
g8706 and b[27] n8589_not ; n8962
g8707 and n8583_not n8962 ; n8963
g8708 and n8591_not n8963_not ; n8964
g8709 and n8961_not n8964 ; n8965
g8710 and n8591_not n8965_not ; n8966
g8711 and b[28] n8580_not ; n8967
g8712 and n8574_not n8967 ; n8968
g8713 and n8582_not n8968_not ; n8969
g8714 and n8966_not n8969 ; n8970
g8715 and n8582_not n8970_not ; n8971
g8716 and b[29] n8571_not ; n8972
g8717 and n8565_not n8972 ; n8973
g8718 and n8573_not n8973_not ; n8974
g8719 and n8971_not n8974 ; n8975
g8720 and n8573_not n8975_not ; n8976
g8721 and b[30] n8562_not ; n8977
g8722 and n8556_not n8977 ; n8978
g8723 and n8564_not n8978_not ; n8979
g8724 and n8976_not n8979 ; n8980
g8725 and n8564_not n8980_not ; n8981
g8726 and b[31] n8553_not ; n8982
g8727 and n8547_not n8982 ; n8983
g8728 and n8555_not n8983_not ; n8984
g8729 and n8981_not n8984 ; n8985
g8730 and n8555_not n8985_not ; n8986
g8731 and b[32] n8544_not ; n8987
g8732 and n8538_not n8987 ; n8988
g8733 and n8546_not n8988_not ; n8989
g8734 and n8986_not n8989 ; n8990
g8735 and n8546_not n8990_not ; n8991
g8736 and b[33] n8527_not ; n8992
g8737 and n8521_not n8992 ; n8993
g8738 and n8537_not n8993_not ; n8994
g8739 and n8991_not n8994 ; n8995
g8740 and n8537_not n8995_not ; n8996
g8741 and b[34] n8529_not ; n8997
g8742 and n8534_not n8997 ; n8998
g8743 and n8536_not n8998_not ; n8999
g8744 and n8996_not n8999 ; n9000
g8745 and n8536_not n9000_not ; n9001
g8746 and n411 n413 ; n9002
g8747 and n422 n9002 ; n9003
g8748 and n408 n9003 ; n9004
g8749 and n9001_not n9004 ; quotient[29]
g8750 and n8528_not quotient[29]_not ; n9006
g8751 and n8546_not n8994 ; n9007
g8752 and n8990_not n9007 ; n9008
g8753 and n8991_not n8994_not ; n9009
g8754 and n9008_not n9009_not ; n9010
g8755 and n9004 n9010_not ; n9011
g8756 and n9001_not n9011 ; n9012
g8757 and n9006_not n9012_not ; n9013
g8758 and b[34]_not n9013_not ; n9014
g8759 and n8545_not quotient[29]_not ; n9015
g8760 and n8555_not n8989 ; n9016
g8761 and n8985_not n9016 ; n9017
g8762 and n8986_not n8989_not ; n9018
g8763 and n9017_not n9018_not ; n9019
g8764 and n9004 n9019_not ; n9020
g8765 and n9001_not n9020 ; n9021
g8766 and n9015_not n9021_not ; n9022
g8767 and b[33]_not n9022_not ; n9023
g8768 and n8554_not quotient[29]_not ; n9024
g8769 and n8564_not n8984 ; n9025
g8770 and n8980_not n9025 ; n9026
g8771 and n8981_not n8984_not ; n9027
g8772 and n9026_not n9027_not ; n9028
g8773 and n9004 n9028_not ; n9029
g8774 and n9001_not n9029 ; n9030
g8775 and n9024_not n9030_not ; n9031
g8776 and b[32]_not n9031_not ; n9032
g8777 and n8563_not quotient[29]_not ; n9033
g8778 and n8573_not n8979 ; n9034
g8779 and n8975_not n9034 ; n9035
g8780 and n8976_not n8979_not ; n9036
g8781 and n9035_not n9036_not ; n9037
g8782 and n9004 n9037_not ; n9038
g8783 and n9001_not n9038 ; n9039
g8784 and n9033_not n9039_not ; n9040
g8785 and b[31]_not n9040_not ; n9041
g8786 and n8572_not quotient[29]_not ; n9042
g8787 and n8582_not n8974 ; n9043
g8788 and n8970_not n9043 ; n9044
g8789 and n8971_not n8974_not ; n9045
g8790 and n9044_not n9045_not ; n9046
g8791 and n9004 n9046_not ; n9047
g8792 and n9001_not n9047 ; n9048
g8793 and n9042_not n9048_not ; n9049
g8794 and b[30]_not n9049_not ; n9050
g8795 and n8581_not quotient[29]_not ; n9051
g8796 and n8591_not n8969 ; n9052
g8797 and n8965_not n9052 ; n9053
g8798 and n8966_not n8969_not ; n9054
g8799 and n9053_not n9054_not ; n9055
g8800 and n9004 n9055_not ; n9056
g8801 and n9001_not n9056 ; n9057
g8802 and n9051_not n9057_not ; n9058
g8803 and b[29]_not n9058_not ; n9059
g8804 and n8590_not quotient[29]_not ; n9060
g8805 and n8600_not n8964 ; n9061
g8806 and n8960_not n9061 ; n9062
g8807 and n8961_not n8964_not ; n9063
g8808 and n9062_not n9063_not ; n9064
g8809 and n9004 n9064_not ; n9065
g8810 and n9001_not n9065 ; n9066
g8811 and n9060_not n9066_not ; n9067
g8812 and b[28]_not n9067_not ; n9068
g8813 and n8599_not quotient[29]_not ; n9069
g8814 and n8609_not n8959 ; n9070
g8815 and n8955_not n9070 ; n9071
g8816 and n8956_not n8959_not ; n9072
g8817 and n9071_not n9072_not ; n9073
g8818 and n9004 n9073_not ; n9074
g8819 and n9001_not n9074 ; n9075
g8820 and n9069_not n9075_not ; n9076
g8821 and b[27]_not n9076_not ; n9077
g8822 and n8608_not quotient[29]_not ; n9078
g8823 and n8618_not n8954 ; n9079
g8824 and n8950_not n9079 ; n9080
g8825 and n8951_not n8954_not ; n9081
g8826 and n9080_not n9081_not ; n9082
g8827 and n9004 n9082_not ; n9083
g8828 and n9001_not n9083 ; n9084
g8829 and n9078_not n9084_not ; n9085
g8830 and b[26]_not n9085_not ; n9086
g8831 and n8617_not quotient[29]_not ; n9087
g8832 and n8627_not n8949 ; n9088
g8833 and n8945_not n9088 ; n9089
g8834 and n8946_not n8949_not ; n9090
g8835 and n9089_not n9090_not ; n9091
g8836 and n9004 n9091_not ; n9092
g8837 and n9001_not n9092 ; n9093
g8838 and n9087_not n9093_not ; n9094
g8839 and b[25]_not n9094_not ; n9095
g8840 and n8626_not quotient[29]_not ; n9096
g8841 and n8636_not n8944 ; n9097
g8842 and n8940_not n9097 ; n9098
g8843 and n8941_not n8944_not ; n9099
g8844 and n9098_not n9099_not ; n9100
g8845 and n9004 n9100_not ; n9101
g8846 and n9001_not n9101 ; n9102
g8847 and n9096_not n9102_not ; n9103
g8848 and b[24]_not n9103_not ; n9104
g8849 and n8635_not quotient[29]_not ; n9105
g8850 and n8645_not n8939 ; n9106
g8851 and n8935_not n9106 ; n9107
g8852 and n8936_not n8939_not ; n9108
g8853 and n9107_not n9108_not ; n9109
g8854 and n9004 n9109_not ; n9110
g8855 and n9001_not n9110 ; n9111
g8856 and n9105_not n9111_not ; n9112
g8857 and b[23]_not n9112_not ; n9113
g8858 and n8644_not quotient[29]_not ; n9114
g8859 and n8654_not n8934 ; n9115
g8860 and n8930_not n9115 ; n9116
g8861 and n8931_not n8934_not ; n9117
g8862 and n9116_not n9117_not ; n9118
g8863 and n9004 n9118_not ; n9119
g8864 and n9001_not n9119 ; n9120
g8865 and n9114_not n9120_not ; n9121
g8866 and b[22]_not n9121_not ; n9122
g8867 and n8653_not quotient[29]_not ; n9123
g8868 and n8663_not n8929 ; n9124
g8869 and n8925_not n9124 ; n9125
g8870 and n8926_not n8929_not ; n9126
g8871 and n9125_not n9126_not ; n9127
g8872 and n9004 n9127_not ; n9128
g8873 and n9001_not n9128 ; n9129
g8874 and n9123_not n9129_not ; n9130
g8875 and b[21]_not n9130_not ; n9131
g8876 and n8662_not quotient[29]_not ; n9132
g8877 and n8672_not n8924 ; n9133
g8878 and n8920_not n9133 ; n9134
g8879 and n8921_not n8924_not ; n9135
g8880 and n9134_not n9135_not ; n9136
g8881 and n9004 n9136_not ; n9137
g8882 and n9001_not n9137 ; n9138
g8883 and n9132_not n9138_not ; n9139
g8884 and b[20]_not n9139_not ; n9140
g8885 and n8671_not quotient[29]_not ; n9141
g8886 and n8681_not n8919 ; n9142
g8887 and n8915_not n9142 ; n9143
g8888 and n8916_not n8919_not ; n9144
g8889 and n9143_not n9144_not ; n9145
g8890 and n9004 n9145_not ; n9146
g8891 and n9001_not n9146 ; n9147
g8892 and n9141_not n9147_not ; n9148
g8893 and b[19]_not n9148_not ; n9149
g8894 and n8680_not quotient[29]_not ; n9150
g8895 and n8690_not n8914 ; n9151
g8896 and n8910_not n9151 ; n9152
g8897 and n8911_not n8914_not ; n9153
g8898 and n9152_not n9153_not ; n9154
g8899 and n9004 n9154_not ; n9155
g8900 and n9001_not n9155 ; n9156
g8901 and n9150_not n9156_not ; n9157
g8902 and b[18]_not n9157_not ; n9158
g8903 and n8689_not quotient[29]_not ; n9159
g8904 and n8699_not n8909 ; n9160
g8905 and n8905_not n9160 ; n9161
g8906 and n8906_not n8909_not ; n9162
g8907 and n9161_not n9162_not ; n9163
g8908 and n9004 n9163_not ; n9164
g8909 and n9001_not n9164 ; n9165
g8910 and n9159_not n9165_not ; n9166
g8911 and b[17]_not n9166_not ; n9167
g8912 and n8698_not quotient[29]_not ; n9168
g8913 and n8708_not n8904 ; n9169
g8914 and n8900_not n9169 ; n9170
g8915 and n8901_not n8904_not ; n9171
g8916 and n9170_not n9171_not ; n9172
g8917 and n9004 n9172_not ; n9173
g8918 and n9001_not n9173 ; n9174
g8919 and n9168_not n9174_not ; n9175
g8920 and b[16]_not n9175_not ; n9176
g8921 and n8707_not quotient[29]_not ; n9177
g8922 and n8717_not n8899 ; n9178
g8923 and n8895_not n9178 ; n9179
g8924 and n8896_not n8899_not ; n9180
g8925 and n9179_not n9180_not ; n9181
g8926 and n9004 n9181_not ; n9182
g8927 and n9001_not n9182 ; n9183
g8928 and n9177_not n9183_not ; n9184
g8929 and b[15]_not n9184_not ; n9185
g8930 and n8716_not quotient[29]_not ; n9186
g8931 and n8726_not n8894 ; n9187
g8932 and n8890_not n9187 ; n9188
g8933 and n8891_not n8894_not ; n9189
g8934 and n9188_not n9189_not ; n9190
g8935 and n9004 n9190_not ; n9191
g8936 and n9001_not n9191 ; n9192
g8937 and n9186_not n9192_not ; n9193
g8938 and b[14]_not n9193_not ; n9194
g8939 and n8725_not quotient[29]_not ; n9195
g8940 and n8735_not n8889 ; n9196
g8941 and n8885_not n9196 ; n9197
g8942 and n8886_not n8889_not ; n9198
g8943 and n9197_not n9198_not ; n9199
g8944 and n9004 n9199_not ; n9200
g8945 and n9001_not n9200 ; n9201
g8946 and n9195_not n9201_not ; n9202
g8947 and b[13]_not n9202_not ; n9203
g8948 and n8734_not quotient[29]_not ; n9204
g8949 and n8744_not n8884 ; n9205
g8950 and n8880_not n9205 ; n9206
g8951 and n8881_not n8884_not ; n9207
g8952 and n9206_not n9207_not ; n9208
g8953 and n9004 n9208_not ; n9209
g8954 and n9001_not n9209 ; n9210
g8955 and n9204_not n9210_not ; n9211
g8956 and b[12]_not n9211_not ; n9212
g8957 and n8743_not quotient[29]_not ; n9213
g8958 and n8753_not n8879 ; n9214
g8959 and n8875_not n9214 ; n9215
g8960 and n8876_not n8879_not ; n9216
g8961 and n9215_not n9216_not ; n9217
g8962 and n9004 n9217_not ; n9218
g8963 and n9001_not n9218 ; n9219
g8964 and n9213_not n9219_not ; n9220
g8965 and b[11]_not n9220_not ; n9221
g8966 and n8752_not quotient[29]_not ; n9222
g8967 and n8762_not n8874 ; n9223
g8968 and n8870_not n9223 ; n9224
g8969 and n8871_not n8874_not ; n9225
g8970 and n9224_not n9225_not ; n9226
g8971 and n9004 n9226_not ; n9227
g8972 and n9001_not n9227 ; n9228
g8973 and n9222_not n9228_not ; n9229
g8974 and b[10]_not n9229_not ; n9230
g8975 and n8761_not quotient[29]_not ; n9231
g8976 and n8771_not n8869 ; n9232
g8977 and n8865_not n9232 ; n9233
g8978 and n8866_not n8869_not ; n9234
g8979 and n9233_not n9234_not ; n9235
g8980 and n9004 n9235_not ; n9236
g8981 and n9001_not n9236 ; n9237
g8982 and n9231_not n9237_not ; n9238
g8983 and b[9]_not n9238_not ; n9239
g8984 and n8770_not quotient[29]_not ; n9240
g8985 and n8780_not n8864 ; n9241
g8986 and n8860_not n9241 ; n9242
g8987 and n8861_not n8864_not ; n9243
g8988 and n9242_not n9243_not ; n9244
g8989 and n9004 n9244_not ; n9245
g8990 and n9001_not n9245 ; n9246
g8991 and n9240_not n9246_not ; n9247
g8992 and b[8]_not n9247_not ; n9248
g8993 and n8779_not quotient[29]_not ; n9249
g8994 and n8789_not n8859 ; n9250
g8995 and n8855_not n9250 ; n9251
g8996 and n8856_not n8859_not ; n9252
g8997 and n9251_not n9252_not ; n9253
g8998 and n9004 n9253_not ; n9254
g8999 and n9001_not n9254 ; n9255
g9000 and n9249_not n9255_not ; n9256
g9001 and b[7]_not n9256_not ; n9257
g9002 and n8788_not quotient[29]_not ; n9258
g9003 and n8798_not n8854 ; n9259
g9004 and n8850_not n9259 ; n9260
g9005 and n8851_not n8854_not ; n9261
g9006 and n9260_not n9261_not ; n9262
g9007 and n9004 n9262_not ; n9263
g9008 and n9001_not n9263 ; n9264
g9009 and n9258_not n9264_not ; n9265
g9010 and b[6]_not n9265_not ; n9266
g9011 and n8797_not quotient[29]_not ; n9267
g9012 and n8807_not n8849 ; n9268
g9013 and n8845_not n9268 ; n9269
g9014 and n8846_not n8849_not ; n9270
g9015 and n9269_not n9270_not ; n9271
g9016 and n9004 n9271_not ; n9272
g9017 and n9001_not n9272 ; n9273
g9018 and n9267_not n9273_not ; n9274
g9019 and b[5]_not n9274_not ; n9275
g9020 and n8806_not quotient[29]_not ; n9276
g9021 and n8815_not n8844 ; n9277
g9022 and n8840_not n9277 ; n9278
g9023 and n8841_not n8844_not ; n9279
g9024 and n9278_not n9279_not ; n9280
g9025 and n9004 n9280_not ; n9281
g9026 and n9001_not n9281 ; n9282
g9027 and n9276_not n9282_not ; n9283
g9028 and b[4]_not n9283_not ; n9284
g9029 and n8814_not quotient[29]_not ; n9285
g9030 and n8835_not n8839 ; n9286
g9031 and n8834_not n9286 ; n9287
g9032 and n8836_not n8839_not ; n9288
g9033 and n9287_not n9288_not ; n9289
g9034 and n9004 n9289_not ; n9290
g9035 and n9001_not n9290 ; n9291
g9036 and n9285_not n9291_not ; n9292
g9037 and b[3]_not n9292_not ; n9293
g9038 and n8828_not quotient[29]_not ; n9294
g9039 and n8831_not n8833 ; n9295
g9040 and n8829_not n9295 ; n9296
g9041 and n9004 n9296_not ; n9297
g9042 and n8834_not n9297 ; n9298
g9043 and n9001_not n9298 ; n9299
g9044 and n9294_not n9299_not ; n9300
g9045 and b[2]_not n9300_not ; n9301
g9046 and b[0] b[35]_not ; n9302
g9047 and n294 n9302 ; n9303
g9048 and n340 n9303 ; n9304
g9049 and n338 n9304 ; n9305
g9050 and n9001_not n9305 ; n9306
g9051 and a[29] n9306_not ; n9307
g9052 and n413 n8833 ; n9308
g9053 and n411 n9308 ; n9309
g9054 and n422 n9309 ; n9310
g9055 and n408 n9310 ; n9311
g9056 and n9001_not n9311 ; n9312
g9057 and n9307_not n9312_not ; n9313
g9058 and b[1] n9313_not ; n9314
g9059 and b[1]_not n9312_not ; n9315
g9060 and n9307_not n9315 ; n9316
g9061 and n9314_not n9316_not ; n9317
g9062 and a[28]_not b[0] ; n9318
g9063 and n9317_not n9318_not ; n9319
g9064 and b[1]_not n9313_not ; n9320
g9065 and n9319_not n9320_not ; n9321
g9066 and b[2] n9299_not ; n9322
g9067 and n9294_not n9322 ; n9323
g9068 and n9301_not n9323_not ; n9324
g9069 and n9321_not n9324 ; n9325
g9070 and n9301_not n9325_not ; n9326
g9071 and b[3] n9291_not ; n9327
g9072 and n9285_not n9327 ; n9328
g9073 and n9293_not n9328_not ; n9329
g9074 and n9326_not n9329 ; n9330
g9075 and n9293_not n9330_not ; n9331
g9076 and b[4] n9282_not ; n9332
g9077 and n9276_not n9332 ; n9333
g9078 and n9284_not n9333_not ; n9334
g9079 and n9331_not n9334 ; n9335
g9080 and n9284_not n9335_not ; n9336
g9081 and b[5] n9273_not ; n9337
g9082 and n9267_not n9337 ; n9338
g9083 and n9275_not n9338_not ; n9339
g9084 and n9336_not n9339 ; n9340
g9085 and n9275_not n9340_not ; n9341
g9086 and b[6] n9264_not ; n9342
g9087 and n9258_not n9342 ; n9343
g9088 and n9266_not n9343_not ; n9344
g9089 and n9341_not n9344 ; n9345
g9090 and n9266_not n9345_not ; n9346
g9091 and b[7] n9255_not ; n9347
g9092 and n9249_not n9347 ; n9348
g9093 and n9257_not n9348_not ; n9349
g9094 and n9346_not n9349 ; n9350
g9095 and n9257_not n9350_not ; n9351
g9096 and b[8] n9246_not ; n9352
g9097 and n9240_not n9352 ; n9353
g9098 and n9248_not n9353_not ; n9354
g9099 and n9351_not n9354 ; n9355
g9100 and n9248_not n9355_not ; n9356
g9101 and b[9] n9237_not ; n9357
g9102 and n9231_not n9357 ; n9358
g9103 and n9239_not n9358_not ; n9359
g9104 and n9356_not n9359 ; n9360
g9105 and n9239_not n9360_not ; n9361
g9106 and b[10] n9228_not ; n9362
g9107 and n9222_not n9362 ; n9363
g9108 and n9230_not n9363_not ; n9364
g9109 and n9361_not n9364 ; n9365
g9110 and n9230_not n9365_not ; n9366
g9111 and b[11] n9219_not ; n9367
g9112 and n9213_not n9367 ; n9368
g9113 and n9221_not n9368_not ; n9369
g9114 and n9366_not n9369 ; n9370
g9115 and n9221_not n9370_not ; n9371
g9116 and b[12] n9210_not ; n9372
g9117 and n9204_not n9372 ; n9373
g9118 and n9212_not n9373_not ; n9374
g9119 and n9371_not n9374 ; n9375
g9120 and n9212_not n9375_not ; n9376
g9121 and b[13] n9201_not ; n9377
g9122 and n9195_not n9377 ; n9378
g9123 and n9203_not n9378_not ; n9379
g9124 and n9376_not n9379 ; n9380
g9125 and n9203_not n9380_not ; n9381
g9126 and b[14] n9192_not ; n9382
g9127 and n9186_not n9382 ; n9383
g9128 and n9194_not n9383_not ; n9384
g9129 and n9381_not n9384 ; n9385
g9130 and n9194_not n9385_not ; n9386
g9131 and b[15] n9183_not ; n9387
g9132 and n9177_not n9387 ; n9388
g9133 and n9185_not n9388_not ; n9389
g9134 and n9386_not n9389 ; n9390
g9135 and n9185_not n9390_not ; n9391
g9136 and b[16] n9174_not ; n9392
g9137 and n9168_not n9392 ; n9393
g9138 and n9176_not n9393_not ; n9394
g9139 and n9391_not n9394 ; n9395
g9140 and n9176_not n9395_not ; n9396
g9141 and b[17] n9165_not ; n9397
g9142 and n9159_not n9397 ; n9398
g9143 and n9167_not n9398_not ; n9399
g9144 and n9396_not n9399 ; n9400
g9145 and n9167_not n9400_not ; n9401
g9146 and b[18] n9156_not ; n9402
g9147 and n9150_not n9402 ; n9403
g9148 and n9158_not n9403_not ; n9404
g9149 and n9401_not n9404 ; n9405
g9150 and n9158_not n9405_not ; n9406
g9151 and b[19] n9147_not ; n9407
g9152 and n9141_not n9407 ; n9408
g9153 and n9149_not n9408_not ; n9409
g9154 and n9406_not n9409 ; n9410
g9155 and n9149_not n9410_not ; n9411
g9156 and b[20] n9138_not ; n9412
g9157 and n9132_not n9412 ; n9413
g9158 and n9140_not n9413_not ; n9414
g9159 and n9411_not n9414 ; n9415
g9160 and n9140_not n9415_not ; n9416
g9161 and b[21] n9129_not ; n9417
g9162 and n9123_not n9417 ; n9418
g9163 and n9131_not n9418_not ; n9419
g9164 and n9416_not n9419 ; n9420
g9165 and n9131_not n9420_not ; n9421
g9166 and b[22] n9120_not ; n9422
g9167 and n9114_not n9422 ; n9423
g9168 and n9122_not n9423_not ; n9424
g9169 and n9421_not n9424 ; n9425
g9170 and n9122_not n9425_not ; n9426
g9171 and b[23] n9111_not ; n9427
g9172 and n9105_not n9427 ; n9428
g9173 and n9113_not n9428_not ; n9429
g9174 and n9426_not n9429 ; n9430
g9175 and n9113_not n9430_not ; n9431
g9176 and b[24] n9102_not ; n9432
g9177 and n9096_not n9432 ; n9433
g9178 and n9104_not n9433_not ; n9434
g9179 and n9431_not n9434 ; n9435
g9180 and n9104_not n9435_not ; n9436
g9181 and b[25] n9093_not ; n9437
g9182 and n9087_not n9437 ; n9438
g9183 and n9095_not n9438_not ; n9439
g9184 and n9436_not n9439 ; n9440
g9185 and n9095_not n9440_not ; n9441
g9186 and b[26] n9084_not ; n9442
g9187 and n9078_not n9442 ; n9443
g9188 and n9086_not n9443_not ; n9444
g9189 and n9441_not n9444 ; n9445
g9190 and n9086_not n9445_not ; n9446
g9191 and b[27] n9075_not ; n9447
g9192 and n9069_not n9447 ; n9448
g9193 and n9077_not n9448_not ; n9449
g9194 and n9446_not n9449 ; n9450
g9195 and n9077_not n9450_not ; n9451
g9196 and b[28] n9066_not ; n9452
g9197 and n9060_not n9452 ; n9453
g9198 and n9068_not n9453_not ; n9454
g9199 and n9451_not n9454 ; n9455
g9200 and n9068_not n9455_not ; n9456
g9201 and b[29] n9057_not ; n9457
g9202 and n9051_not n9457 ; n9458
g9203 and n9059_not n9458_not ; n9459
g9204 and n9456_not n9459 ; n9460
g9205 and n9059_not n9460_not ; n9461
g9206 and b[30] n9048_not ; n9462
g9207 and n9042_not n9462 ; n9463
g9208 and n9050_not n9463_not ; n9464
g9209 and n9461_not n9464 ; n9465
g9210 and n9050_not n9465_not ; n9466
g9211 and b[31] n9039_not ; n9467
g9212 and n9033_not n9467 ; n9468
g9213 and n9041_not n9468_not ; n9469
g9214 and n9466_not n9469 ; n9470
g9215 and n9041_not n9470_not ; n9471
g9216 and b[32] n9030_not ; n9472
g9217 and n9024_not n9472 ; n9473
g9218 and n9032_not n9473_not ; n9474
g9219 and n9471_not n9474 ; n9475
g9220 and n9032_not n9475_not ; n9476
g9221 and b[33] n9021_not ; n9477
g9222 and n9015_not n9477 ; n9478
g9223 and n9023_not n9478_not ; n9479
g9224 and n9476_not n9479 ; n9480
g9225 and n9023_not n9480_not ; n9481
g9226 and b[34] n9012_not ; n9482
g9227 and n9006_not n9482 ; n9483
g9228 and n9014_not n9483_not ; n9484
g9229 and n9481_not n9484 ; n9485
g9230 and n9014_not n9485_not ; n9486
g9231 and n8535_not quotient[29]_not ; n9487
g9232 and n8537_not n8999 ; n9488
g9233 and n8995_not n9488 ; n9489
g9234 and n8996_not n8999_not ; n9490
g9235 and n9489_not n9490_not ; n9491
g9236 and quotient[29] n9491_not ; n9492
g9237 and n9487_not n9492_not ; n9493
g9238 and b[35]_not n9493_not ; n9494
g9239 and b[35] n9487_not ; n9495
g9240 and n9492_not n9495 ; n9496
g9241 and n512 n9496_not ; n9497
g9242 and n9494_not n9497 ; n9498
g9243 and n9486_not n9498 ; n9499
g9244 and n9004 n9493_not ; n9500
g9245 and n9499_not n9500_not ; quotient[28]
g9246 and n9023_not n9484 ; n9502
g9247 and n9480_not n9502 ; n9503
g9248 and n9481_not n9484_not ; n9504
g9249 and n9503_not n9504_not ; n9505
g9250 and quotient[28] n9505_not ; n9506
g9251 and n9013_not n9500_not ; n9507
g9252 and n9499_not n9507 ; n9508
g9253 and n9506_not n9508_not ; n9509
g9254 and n9014_not n9496_not ; n9510
g9255 and n9494_not n9510 ; n9511
g9256 and n9485_not n9511 ; n9512
g9257 and n9494_not n9496_not ; n9513
g9258 and n9486_not n9513_not ; n9514
g9259 and n9512_not n9514_not ; n9515
g9260 and quotient[28] n9515_not ; n9516
g9261 and n9493_not n9500_not ; n9517
g9262 and n9499_not n9517 ; n9518
g9263 and n9516_not n9518_not ; n9519
g9264 and b[36]_not n9519_not ; n9520
g9265 and b[35]_not n9509_not ; n9521
g9266 and n9032_not n9479 ; n9522
g9267 and n9475_not n9522 ; n9523
g9268 and n9476_not n9479_not ; n9524
g9269 and n9523_not n9524_not ; n9525
g9270 and quotient[28] n9525_not ; n9526
g9271 and n9022_not n9500_not ; n9527
g9272 and n9499_not n9527 ; n9528
g9273 and n9526_not n9528_not ; n9529
g9274 and b[34]_not n9529_not ; n9530
g9275 and n9041_not n9474 ; n9531
g9276 and n9470_not n9531 ; n9532
g9277 and n9471_not n9474_not ; n9533
g9278 and n9532_not n9533_not ; n9534
g9279 and quotient[28] n9534_not ; n9535
g9280 and n9031_not n9500_not ; n9536
g9281 and n9499_not n9536 ; n9537
g9282 and n9535_not n9537_not ; n9538
g9283 and b[33]_not n9538_not ; n9539
g9284 and n9050_not n9469 ; n9540
g9285 and n9465_not n9540 ; n9541
g9286 and n9466_not n9469_not ; n9542
g9287 and n9541_not n9542_not ; n9543
g9288 and quotient[28] n9543_not ; n9544
g9289 and n9040_not n9500_not ; n9545
g9290 and n9499_not n9545 ; n9546
g9291 and n9544_not n9546_not ; n9547
g9292 and b[32]_not n9547_not ; n9548
g9293 and n9059_not n9464 ; n9549
g9294 and n9460_not n9549 ; n9550
g9295 and n9461_not n9464_not ; n9551
g9296 and n9550_not n9551_not ; n9552
g9297 and quotient[28] n9552_not ; n9553
g9298 and n9049_not n9500_not ; n9554
g9299 and n9499_not n9554 ; n9555
g9300 and n9553_not n9555_not ; n9556
g9301 and b[31]_not n9556_not ; n9557
g9302 and n9068_not n9459 ; n9558
g9303 and n9455_not n9558 ; n9559
g9304 and n9456_not n9459_not ; n9560
g9305 and n9559_not n9560_not ; n9561
g9306 and quotient[28] n9561_not ; n9562
g9307 and n9058_not n9500_not ; n9563
g9308 and n9499_not n9563 ; n9564
g9309 and n9562_not n9564_not ; n9565
g9310 and b[30]_not n9565_not ; n9566
g9311 and n9077_not n9454 ; n9567
g9312 and n9450_not n9567 ; n9568
g9313 and n9451_not n9454_not ; n9569
g9314 and n9568_not n9569_not ; n9570
g9315 and quotient[28] n9570_not ; n9571
g9316 and n9067_not n9500_not ; n9572
g9317 and n9499_not n9572 ; n9573
g9318 and n9571_not n9573_not ; n9574
g9319 and b[29]_not n9574_not ; n9575
g9320 and n9086_not n9449 ; n9576
g9321 and n9445_not n9576 ; n9577
g9322 and n9446_not n9449_not ; n9578
g9323 and n9577_not n9578_not ; n9579
g9324 and quotient[28] n9579_not ; n9580
g9325 and n9076_not n9500_not ; n9581
g9326 and n9499_not n9581 ; n9582
g9327 and n9580_not n9582_not ; n9583
g9328 and b[28]_not n9583_not ; n9584
g9329 and n9095_not n9444 ; n9585
g9330 and n9440_not n9585 ; n9586
g9331 and n9441_not n9444_not ; n9587
g9332 and n9586_not n9587_not ; n9588
g9333 and quotient[28] n9588_not ; n9589
g9334 and n9085_not n9500_not ; n9590
g9335 and n9499_not n9590 ; n9591
g9336 and n9589_not n9591_not ; n9592
g9337 and b[27]_not n9592_not ; n9593
g9338 and n9104_not n9439 ; n9594
g9339 and n9435_not n9594 ; n9595
g9340 and n9436_not n9439_not ; n9596
g9341 and n9595_not n9596_not ; n9597
g9342 and quotient[28] n9597_not ; n9598
g9343 and n9094_not n9500_not ; n9599
g9344 and n9499_not n9599 ; n9600
g9345 and n9598_not n9600_not ; n9601
g9346 and b[26]_not n9601_not ; n9602
g9347 and n9113_not n9434 ; n9603
g9348 and n9430_not n9603 ; n9604
g9349 and n9431_not n9434_not ; n9605
g9350 and n9604_not n9605_not ; n9606
g9351 and quotient[28] n9606_not ; n9607
g9352 and n9103_not n9500_not ; n9608
g9353 and n9499_not n9608 ; n9609
g9354 and n9607_not n9609_not ; n9610
g9355 and b[25]_not n9610_not ; n9611
g9356 and n9122_not n9429 ; n9612
g9357 and n9425_not n9612 ; n9613
g9358 and n9426_not n9429_not ; n9614
g9359 and n9613_not n9614_not ; n9615
g9360 and quotient[28] n9615_not ; n9616
g9361 and n9112_not n9500_not ; n9617
g9362 and n9499_not n9617 ; n9618
g9363 and n9616_not n9618_not ; n9619
g9364 and b[24]_not n9619_not ; n9620
g9365 and n9131_not n9424 ; n9621
g9366 and n9420_not n9621 ; n9622
g9367 and n9421_not n9424_not ; n9623
g9368 and n9622_not n9623_not ; n9624
g9369 and quotient[28] n9624_not ; n9625
g9370 and n9121_not n9500_not ; n9626
g9371 and n9499_not n9626 ; n9627
g9372 and n9625_not n9627_not ; n9628
g9373 and b[23]_not n9628_not ; n9629
g9374 and n9140_not n9419 ; n9630
g9375 and n9415_not n9630 ; n9631
g9376 and n9416_not n9419_not ; n9632
g9377 and n9631_not n9632_not ; n9633
g9378 and quotient[28] n9633_not ; n9634
g9379 and n9130_not n9500_not ; n9635
g9380 and n9499_not n9635 ; n9636
g9381 and n9634_not n9636_not ; n9637
g9382 and b[22]_not n9637_not ; n9638
g9383 and n9149_not n9414 ; n9639
g9384 and n9410_not n9639 ; n9640
g9385 and n9411_not n9414_not ; n9641
g9386 and n9640_not n9641_not ; n9642
g9387 and quotient[28] n9642_not ; n9643
g9388 and n9139_not n9500_not ; n9644
g9389 and n9499_not n9644 ; n9645
g9390 and n9643_not n9645_not ; n9646
g9391 and b[21]_not n9646_not ; n9647
g9392 and n9158_not n9409 ; n9648
g9393 and n9405_not n9648 ; n9649
g9394 and n9406_not n9409_not ; n9650
g9395 and n9649_not n9650_not ; n9651
g9396 and quotient[28] n9651_not ; n9652
g9397 and n9148_not n9500_not ; n9653
g9398 and n9499_not n9653 ; n9654
g9399 and n9652_not n9654_not ; n9655
g9400 and b[20]_not n9655_not ; n9656
g9401 and n9167_not n9404 ; n9657
g9402 and n9400_not n9657 ; n9658
g9403 and n9401_not n9404_not ; n9659
g9404 and n9658_not n9659_not ; n9660
g9405 and quotient[28] n9660_not ; n9661
g9406 and n9157_not n9500_not ; n9662
g9407 and n9499_not n9662 ; n9663
g9408 and n9661_not n9663_not ; n9664
g9409 and b[19]_not n9664_not ; n9665
g9410 and n9176_not n9399 ; n9666
g9411 and n9395_not n9666 ; n9667
g9412 and n9396_not n9399_not ; n9668
g9413 and n9667_not n9668_not ; n9669
g9414 and quotient[28] n9669_not ; n9670
g9415 and n9166_not n9500_not ; n9671
g9416 and n9499_not n9671 ; n9672
g9417 and n9670_not n9672_not ; n9673
g9418 and b[18]_not n9673_not ; n9674
g9419 and n9185_not n9394 ; n9675
g9420 and n9390_not n9675 ; n9676
g9421 and n9391_not n9394_not ; n9677
g9422 and n9676_not n9677_not ; n9678
g9423 and quotient[28] n9678_not ; n9679
g9424 and n9175_not n9500_not ; n9680
g9425 and n9499_not n9680 ; n9681
g9426 and n9679_not n9681_not ; n9682
g9427 and b[17]_not n9682_not ; n9683
g9428 and n9194_not n9389 ; n9684
g9429 and n9385_not n9684 ; n9685
g9430 and n9386_not n9389_not ; n9686
g9431 and n9685_not n9686_not ; n9687
g9432 and quotient[28] n9687_not ; n9688
g9433 and n9184_not n9500_not ; n9689
g9434 and n9499_not n9689 ; n9690
g9435 and n9688_not n9690_not ; n9691
g9436 and b[16]_not n9691_not ; n9692
g9437 and n9203_not n9384 ; n9693
g9438 and n9380_not n9693 ; n9694
g9439 and n9381_not n9384_not ; n9695
g9440 and n9694_not n9695_not ; n9696
g9441 and quotient[28] n9696_not ; n9697
g9442 and n9193_not n9500_not ; n9698
g9443 and n9499_not n9698 ; n9699
g9444 and n9697_not n9699_not ; n9700
g9445 and b[15]_not n9700_not ; n9701
g9446 and n9212_not n9379 ; n9702
g9447 and n9375_not n9702 ; n9703
g9448 and n9376_not n9379_not ; n9704
g9449 and n9703_not n9704_not ; n9705
g9450 and quotient[28] n9705_not ; n9706
g9451 and n9202_not n9500_not ; n9707
g9452 and n9499_not n9707 ; n9708
g9453 and n9706_not n9708_not ; n9709
g9454 and b[14]_not n9709_not ; n9710
g9455 and n9221_not n9374 ; n9711
g9456 and n9370_not n9711 ; n9712
g9457 and n9371_not n9374_not ; n9713
g9458 and n9712_not n9713_not ; n9714
g9459 and quotient[28] n9714_not ; n9715
g9460 and n9211_not n9500_not ; n9716
g9461 and n9499_not n9716 ; n9717
g9462 and n9715_not n9717_not ; n9718
g9463 and b[13]_not n9718_not ; n9719
g9464 and n9230_not n9369 ; n9720
g9465 and n9365_not n9720 ; n9721
g9466 and n9366_not n9369_not ; n9722
g9467 and n9721_not n9722_not ; n9723
g9468 and quotient[28] n9723_not ; n9724
g9469 and n9220_not n9500_not ; n9725
g9470 and n9499_not n9725 ; n9726
g9471 and n9724_not n9726_not ; n9727
g9472 and b[12]_not n9727_not ; n9728
g9473 and n9239_not n9364 ; n9729
g9474 and n9360_not n9729 ; n9730
g9475 and n9361_not n9364_not ; n9731
g9476 and n9730_not n9731_not ; n9732
g9477 and quotient[28] n9732_not ; n9733
g9478 and n9229_not n9500_not ; n9734
g9479 and n9499_not n9734 ; n9735
g9480 and n9733_not n9735_not ; n9736
g9481 and b[11]_not n9736_not ; n9737
g9482 and n9248_not n9359 ; n9738
g9483 and n9355_not n9738 ; n9739
g9484 and n9356_not n9359_not ; n9740
g9485 and n9739_not n9740_not ; n9741
g9486 and quotient[28] n9741_not ; n9742
g9487 and n9238_not n9500_not ; n9743
g9488 and n9499_not n9743 ; n9744
g9489 and n9742_not n9744_not ; n9745
g9490 and b[10]_not n9745_not ; n9746
g9491 and n9257_not n9354 ; n9747
g9492 and n9350_not n9747 ; n9748
g9493 and n9351_not n9354_not ; n9749
g9494 and n9748_not n9749_not ; n9750
g9495 and quotient[28] n9750_not ; n9751
g9496 and n9247_not n9500_not ; n9752
g9497 and n9499_not n9752 ; n9753
g9498 and n9751_not n9753_not ; n9754
g9499 and b[9]_not n9754_not ; n9755
g9500 and n9266_not n9349 ; n9756
g9501 and n9345_not n9756 ; n9757
g9502 and n9346_not n9349_not ; n9758
g9503 and n9757_not n9758_not ; n9759
g9504 and quotient[28] n9759_not ; n9760
g9505 and n9256_not n9500_not ; n9761
g9506 and n9499_not n9761 ; n9762
g9507 and n9760_not n9762_not ; n9763
g9508 and b[8]_not n9763_not ; n9764
g9509 and n9275_not n9344 ; n9765
g9510 and n9340_not n9765 ; n9766
g9511 and n9341_not n9344_not ; n9767
g9512 and n9766_not n9767_not ; n9768
g9513 and quotient[28] n9768_not ; n9769
g9514 and n9265_not n9500_not ; n9770
g9515 and n9499_not n9770 ; n9771
g9516 and n9769_not n9771_not ; n9772
g9517 and b[7]_not n9772_not ; n9773
g9518 and n9284_not n9339 ; n9774
g9519 and n9335_not n9774 ; n9775
g9520 and n9336_not n9339_not ; n9776
g9521 and n9775_not n9776_not ; n9777
g9522 and quotient[28] n9777_not ; n9778
g9523 and n9274_not n9500_not ; n9779
g9524 and n9499_not n9779 ; n9780
g9525 and n9778_not n9780_not ; n9781
g9526 and b[6]_not n9781_not ; n9782
g9527 and n9293_not n9334 ; n9783
g9528 and n9330_not n9783 ; n9784
g9529 and n9331_not n9334_not ; n9785
g9530 and n9784_not n9785_not ; n9786
g9531 and quotient[28] n9786_not ; n9787
g9532 and n9283_not n9500_not ; n9788
g9533 and n9499_not n9788 ; n9789
g9534 and n9787_not n9789_not ; n9790
g9535 and b[5]_not n9790_not ; n9791
g9536 and n9301_not n9329 ; n9792
g9537 and n9325_not n9792 ; n9793
g9538 and n9326_not n9329_not ; n9794
g9539 and n9793_not n9794_not ; n9795
g9540 and quotient[28] n9795_not ; n9796
g9541 and n9292_not n9500_not ; n9797
g9542 and n9499_not n9797 ; n9798
g9543 and n9796_not n9798_not ; n9799
g9544 and b[4]_not n9799_not ; n9800
g9545 and n9320_not n9324 ; n9801
g9546 and n9319_not n9801 ; n9802
g9547 and n9321_not n9324_not ; n9803
g9548 and n9802_not n9803_not ; n9804
g9549 and quotient[28] n9804_not ; n9805
g9550 and n9300_not n9500_not ; n9806
g9551 and n9499_not n9806 ; n9807
g9552 and n9805_not n9807_not ; n9808
g9553 and b[3]_not n9808_not ; n9809
g9554 and n9316_not n9318 ; n9810
g9555 and n9314_not n9810 ; n9811
g9556 and n9319_not n9811_not ; n9812
g9557 and quotient[28] n9812 ; n9813
g9558 and n9313_not n9500_not ; n9814
g9559 and n9499_not n9814 ; n9815
g9560 and n9813_not n9815_not ; n9816
g9561 and b[2]_not n9816_not ; n9817
g9562 and b[0] quotient[28] ; n9818
g9563 and a[28] n9818_not ; n9819
g9564 and n9318 quotient[28] ; n9820
g9565 and n9819_not n9820_not ; n9821
g9566 and b[1] n9821_not ; n9822
g9567 and b[1]_not n9820_not ; n9823
g9568 and n9819_not n9823 ; n9824
g9569 and n9822_not n9824_not ; n9825
g9570 and a[27]_not b[0] ; n9826
g9571 and n9825_not n9826_not ; n9827
g9572 and b[1]_not n9821_not ; n9828
g9573 and n9827_not n9828_not ; n9829
g9574 and b[2] n9815_not ; n9830
g9575 and n9813_not n9830 ; n9831
g9576 and n9817_not n9831_not ; n9832
g9577 and n9829_not n9832 ; n9833
g9578 and n9817_not n9833_not ; n9834
g9579 and b[3] n9807_not ; n9835
g9580 and n9805_not n9835 ; n9836
g9581 and n9809_not n9836_not ; n9837
g9582 and n9834_not n9837 ; n9838
g9583 and n9809_not n9838_not ; n9839
g9584 and b[4] n9798_not ; n9840
g9585 and n9796_not n9840 ; n9841
g9586 and n9800_not n9841_not ; n9842
g9587 and n9839_not n9842 ; n9843
g9588 and n9800_not n9843_not ; n9844
g9589 and b[5] n9789_not ; n9845
g9590 and n9787_not n9845 ; n9846
g9591 and n9791_not n9846_not ; n9847
g9592 and n9844_not n9847 ; n9848
g9593 and n9791_not n9848_not ; n9849
g9594 and b[6] n9780_not ; n9850
g9595 and n9778_not n9850 ; n9851
g9596 and n9782_not n9851_not ; n9852
g9597 and n9849_not n9852 ; n9853
g9598 and n9782_not n9853_not ; n9854
g9599 and b[7] n9771_not ; n9855
g9600 and n9769_not n9855 ; n9856
g9601 and n9773_not n9856_not ; n9857
g9602 and n9854_not n9857 ; n9858
g9603 and n9773_not n9858_not ; n9859
g9604 and b[8] n9762_not ; n9860
g9605 and n9760_not n9860 ; n9861
g9606 and n9764_not n9861_not ; n9862
g9607 and n9859_not n9862 ; n9863
g9608 and n9764_not n9863_not ; n9864
g9609 and b[9] n9753_not ; n9865
g9610 and n9751_not n9865 ; n9866
g9611 and n9755_not n9866_not ; n9867
g9612 and n9864_not n9867 ; n9868
g9613 and n9755_not n9868_not ; n9869
g9614 and b[10] n9744_not ; n9870
g9615 and n9742_not n9870 ; n9871
g9616 and n9746_not n9871_not ; n9872
g9617 and n9869_not n9872 ; n9873
g9618 and n9746_not n9873_not ; n9874
g9619 and b[11] n9735_not ; n9875
g9620 and n9733_not n9875 ; n9876
g9621 and n9737_not n9876_not ; n9877
g9622 and n9874_not n9877 ; n9878
g9623 and n9737_not n9878_not ; n9879
g9624 and b[12] n9726_not ; n9880
g9625 and n9724_not n9880 ; n9881
g9626 and n9728_not n9881_not ; n9882
g9627 and n9879_not n9882 ; n9883
g9628 and n9728_not n9883_not ; n9884
g9629 and b[13] n9717_not ; n9885
g9630 and n9715_not n9885 ; n9886
g9631 and n9719_not n9886_not ; n9887
g9632 and n9884_not n9887 ; n9888
g9633 and n9719_not n9888_not ; n9889
g9634 and b[14] n9708_not ; n9890
g9635 and n9706_not n9890 ; n9891
g9636 and n9710_not n9891_not ; n9892
g9637 and n9889_not n9892 ; n9893
g9638 and n9710_not n9893_not ; n9894
g9639 and b[15] n9699_not ; n9895
g9640 and n9697_not n9895 ; n9896
g9641 and n9701_not n9896_not ; n9897
g9642 and n9894_not n9897 ; n9898
g9643 and n9701_not n9898_not ; n9899
g9644 and b[16] n9690_not ; n9900
g9645 and n9688_not n9900 ; n9901
g9646 and n9692_not n9901_not ; n9902
g9647 and n9899_not n9902 ; n9903
g9648 and n9692_not n9903_not ; n9904
g9649 and b[17] n9681_not ; n9905
g9650 and n9679_not n9905 ; n9906
g9651 and n9683_not n9906_not ; n9907
g9652 and n9904_not n9907 ; n9908
g9653 and n9683_not n9908_not ; n9909
g9654 and b[18] n9672_not ; n9910
g9655 and n9670_not n9910 ; n9911
g9656 and n9674_not n9911_not ; n9912
g9657 and n9909_not n9912 ; n9913
g9658 and n9674_not n9913_not ; n9914
g9659 and b[19] n9663_not ; n9915
g9660 and n9661_not n9915 ; n9916
g9661 and n9665_not n9916_not ; n9917
g9662 and n9914_not n9917 ; n9918
g9663 and n9665_not n9918_not ; n9919
g9664 and b[20] n9654_not ; n9920
g9665 and n9652_not n9920 ; n9921
g9666 and n9656_not n9921_not ; n9922
g9667 and n9919_not n9922 ; n9923
g9668 and n9656_not n9923_not ; n9924
g9669 and b[21] n9645_not ; n9925
g9670 and n9643_not n9925 ; n9926
g9671 and n9647_not n9926_not ; n9927
g9672 and n9924_not n9927 ; n9928
g9673 and n9647_not n9928_not ; n9929
g9674 and b[22] n9636_not ; n9930
g9675 and n9634_not n9930 ; n9931
g9676 and n9638_not n9931_not ; n9932
g9677 and n9929_not n9932 ; n9933
g9678 and n9638_not n9933_not ; n9934
g9679 and b[23] n9627_not ; n9935
g9680 and n9625_not n9935 ; n9936
g9681 and n9629_not n9936_not ; n9937
g9682 and n9934_not n9937 ; n9938
g9683 and n9629_not n9938_not ; n9939
g9684 and b[24] n9618_not ; n9940
g9685 and n9616_not n9940 ; n9941
g9686 and n9620_not n9941_not ; n9942
g9687 and n9939_not n9942 ; n9943
g9688 and n9620_not n9943_not ; n9944
g9689 and b[25] n9609_not ; n9945
g9690 and n9607_not n9945 ; n9946
g9691 and n9611_not n9946_not ; n9947
g9692 and n9944_not n9947 ; n9948
g9693 and n9611_not n9948_not ; n9949
g9694 and b[26] n9600_not ; n9950
g9695 and n9598_not n9950 ; n9951
g9696 and n9602_not n9951_not ; n9952
g9697 and n9949_not n9952 ; n9953
g9698 and n9602_not n9953_not ; n9954
g9699 and b[27] n9591_not ; n9955
g9700 and n9589_not n9955 ; n9956
g9701 and n9593_not n9956_not ; n9957
g9702 and n9954_not n9957 ; n9958
g9703 and n9593_not n9958_not ; n9959
g9704 and b[28] n9582_not ; n9960
g9705 and n9580_not n9960 ; n9961
g9706 and n9584_not n9961_not ; n9962
g9707 and n9959_not n9962 ; n9963
g9708 and n9584_not n9963_not ; n9964
g9709 and b[29] n9573_not ; n9965
g9710 and n9571_not n9965 ; n9966
g9711 and n9575_not n9966_not ; n9967
g9712 and n9964_not n9967 ; n9968
g9713 and n9575_not n9968_not ; n9969
g9714 and b[30] n9564_not ; n9970
g9715 and n9562_not n9970 ; n9971
g9716 and n9566_not n9971_not ; n9972
g9717 and n9969_not n9972 ; n9973
g9718 and n9566_not n9973_not ; n9974
g9719 and b[31] n9555_not ; n9975
g9720 and n9553_not n9975 ; n9976
g9721 and n9557_not n9976_not ; n9977
g9722 and n9974_not n9977 ; n9978
g9723 and n9557_not n9978_not ; n9979
g9724 and b[32] n9546_not ; n9980
g9725 and n9544_not n9980 ; n9981
g9726 and n9548_not n9981_not ; n9982
g9727 and n9979_not n9982 ; n9983
g9728 and n9548_not n9983_not ; n9984
g9729 and b[33] n9537_not ; n9985
g9730 and n9535_not n9985 ; n9986
g9731 and n9539_not n9986_not ; n9987
g9732 and n9984_not n9987 ; n9988
g9733 and n9539_not n9988_not ; n9989
g9734 and b[34] n9528_not ; n9990
g9735 and n9526_not n9990 ; n9991
g9736 and n9530_not n9991_not ; n9992
g9737 and n9989_not n9992 ; n9993
g9738 and n9530_not n9993_not ; n9994
g9739 and b[35] n9508_not ; n9995
g9740 and n9506_not n9995 ; n9996
g9741 and n9521_not n9996_not ; n9997
g9742 and n9994_not n9997 ; n9998
g9743 and n9521_not n9998_not ; n9999
g9744 and b[36] n9518_not ; n10000
g9745 and n9516_not n10000 ; n10001
g9746 and n9520_not n10001_not ; n10002
g9747 and n9999_not n10002 ; n10003
g9748 and n9520_not n10003_not ; n10004
g9749 and n599 n10004_not ; quotient[27]
g9750 and n9509_not quotient[27]_not ; n10006
g9751 and n9530_not n9997 ; n10007
g9752 and n9993_not n10007 ; n10008
g9753 and n9994_not n9997_not ; n10009
g9754 and n10008_not n10009_not ; n10010
g9755 and n599 n10010_not ; n10011
g9756 and n10004_not n10011 ; n10012
g9757 and n10006_not n10012_not ; n10013
g9758 and n9519_not quotient[27]_not ; n10014
g9759 and n9521_not n10002 ; n10015
g9760 and n9998_not n10015 ; n10016
g9761 and n9999_not n10002_not ; n10017
g9762 and n10016_not n10017_not ; n10018
g9763 and quotient[27] n10018_not ; n10019
g9764 and n10014_not n10019_not ; n10020
g9765 and b[37]_not n10020_not ; n10021
g9766 and b[36]_not n10013_not ; n10022
g9767 and n9529_not quotient[27]_not ; n10023
g9768 and n9539_not n9992 ; n10024
g9769 and n9988_not n10024 ; n10025
g9770 and n9989_not n9992_not ; n10026
g9771 and n10025_not n10026_not ; n10027
g9772 and n599 n10027_not ; n10028
g9773 and n10004_not n10028 ; n10029
g9774 and n10023_not n10029_not ; n10030
g9775 and b[35]_not n10030_not ; n10031
g9776 and n9538_not quotient[27]_not ; n10032
g9777 and n9548_not n9987 ; n10033
g9778 and n9983_not n10033 ; n10034
g9779 and n9984_not n9987_not ; n10035
g9780 and n10034_not n10035_not ; n10036
g9781 and n599 n10036_not ; n10037
g9782 and n10004_not n10037 ; n10038
g9783 and n10032_not n10038_not ; n10039
g9784 and b[34]_not n10039_not ; n10040
g9785 and n9547_not quotient[27]_not ; n10041
g9786 and n9557_not n9982 ; n10042
g9787 and n9978_not n10042 ; n10043
g9788 and n9979_not n9982_not ; n10044
g9789 and n10043_not n10044_not ; n10045
g9790 and n599 n10045_not ; n10046
g9791 and n10004_not n10046 ; n10047
g9792 and n10041_not n10047_not ; n10048
g9793 and b[33]_not n10048_not ; n10049
g9794 and n9556_not quotient[27]_not ; n10050
g9795 and n9566_not n9977 ; n10051
g9796 and n9973_not n10051 ; n10052
g9797 and n9974_not n9977_not ; n10053
g9798 and n10052_not n10053_not ; n10054
g9799 and n599 n10054_not ; n10055
g9800 and n10004_not n10055 ; n10056
g9801 and n10050_not n10056_not ; n10057
g9802 and b[32]_not n10057_not ; n10058
g9803 and n9565_not quotient[27]_not ; n10059
g9804 and n9575_not n9972 ; n10060
g9805 and n9968_not n10060 ; n10061
g9806 and n9969_not n9972_not ; n10062
g9807 and n10061_not n10062_not ; n10063
g9808 and n599 n10063_not ; n10064
g9809 and n10004_not n10064 ; n10065
g9810 and n10059_not n10065_not ; n10066
g9811 and b[31]_not n10066_not ; n10067
g9812 and n9574_not quotient[27]_not ; n10068
g9813 and n9584_not n9967 ; n10069
g9814 and n9963_not n10069 ; n10070
g9815 and n9964_not n9967_not ; n10071
g9816 and n10070_not n10071_not ; n10072
g9817 and n599 n10072_not ; n10073
g9818 and n10004_not n10073 ; n10074
g9819 and n10068_not n10074_not ; n10075
g9820 and b[30]_not n10075_not ; n10076
g9821 and n9583_not quotient[27]_not ; n10077
g9822 and n9593_not n9962 ; n10078
g9823 and n9958_not n10078 ; n10079
g9824 and n9959_not n9962_not ; n10080
g9825 and n10079_not n10080_not ; n10081
g9826 and n599 n10081_not ; n10082
g9827 and n10004_not n10082 ; n10083
g9828 and n10077_not n10083_not ; n10084
g9829 and b[29]_not n10084_not ; n10085
g9830 and n9592_not quotient[27]_not ; n10086
g9831 and n9602_not n9957 ; n10087
g9832 and n9953_not n10087 ; n10088
g9833 and n9954_not n9957_not ; n10089
g9834 and n10088_not n10089_not ; n10090
g9835 and n599 n10090_not ; n10091
g9836 and n10004_not n10091 ; n10092
g9837 and n10086_not n10092_not ; n10093
g9838 and b[28]_not n10093_not ; n10094
g9839 and n9601_not quotient[27]_not ; n10095
g9840 and n9611_not n9952 ; n10096
g9841 and n9948_not n10096 ; n10097
g9842 and n9949_not n9952_not ; n10098
g9843 and n10097_not n10098_not ; n10099
g9844 and n599 n10099_not ; n10100
g9845 and n10004_not n10100 ; n10101
g9846 and n10095_not n10101_not ; n10102
g9847 and b[27]_not n10102_not ; n10103
g9848 and n9610_not quotient[27]_not ; n10104
g9849 and n9620_not n9947 ; n10105
g9850 and n9943_not n10105 ; n10106
g9851 and n9944_not n9947_not ; n10107
g9852 and n10106_not n10107_not ; n10108
g9853 and n599 n10108_not ; n10109
g9854 and n10004_not n10109 ; n10110
g9855 and n10104_not n10110_not ; n10111
g9856 and b[26]_not n10111_not ; n10112
g9857 and n9619_not quotient[27]_not ; n10113
g9858 and n9629_not n9942 ; n10114
g9859 and n9938_not n10114 ; n10115
g9860 and n9939_not n9942_not ; n10116
g9861 and n10115_not n10116_not ; n10117
g9862 and n599 n10117_not ; n10118
g9863 and n10004_not n10118 ; n10119
g9864 and n10113_not n10119_not ; n10120
g9865 and b[25]_not n10120_not ; n10121
g9866 and n9628_not quotient[27]_not ; n10122
g9867 and n9638_not n9937 ; n10123
g9868 and n9933_not n10123 ; n10124
g9869 and n9934_not n9937_not ; n10125
g9870 and n10124_not n10125_not ; n10126
g9871 and n599 n10126_not ; n10127
g9872 and n10004_not n10127 ; n10128
g9873 and n10122_not n10128_not ; n10129
g9874 and b[24]_not n10129_not ; n10130
g9875 and n9637_not quotient[27]_not ; n10131
g9876 and n9647_not n9932 ; n10132
g9877 and n9928_not n10132 ; n10133
g9878 and n9929_not n9932_not ; n10134
g9879 and n10133_not n10134_not ; n10135
g9880 and n599 n10135_not ; n10136
g9881 and n10004_not n10136 ; n10137
g9882 and n10131_not n10137_not ; n10138
g9883 and b[23]_not n10138_not ; n10139
g9884 and n9646_not quotient[27]_not ; n10140
g9885 and n9656_not n9927 ; n10141
g9886 and n9923_not n10141 ; n10142
g9887 and n9924_not n9927_not ; n10143
g9888 and n10142_not n10143_not ; n10144
g9889 and n599 n10144_not ; n10145
g9890 and n10004_not n10145 ; n10146
g9891 and n10140_not n10146_not ; n10147
g9892 and b[22]_not n10147_not ; n10148
g9893 and n9655_not quotient[27]_not ; n10149
g9894 and n9665_not n9922 ; n10150
g9895 and n9918_not n10150 ; n10151
g9896 and n9919_not n9922_not ; n10152
g9897 and n10151_not n10152_not ; n10153
g9898 and n599 n10153_not ; n10154
g9899 and n10004_not n10154 ; n10155
g9900 and n10149_not n10155_not ; n10156
g9901 and b[21]_not n10156_not ; n10157
g9902 and n9664_not quotient[27]_not ; n10158
g9903 and n9674_not n9917 ; n10159
g9904 and n9913_not n10159 ; n10160
g9905 and n9914_not n9917_not ; n10161
g9906 and n10160_not n10161_not ; n10162
g9907 and n599 n10162_not ; n10163
g9908 and n10004_not n10163 ; n10164
g9909 and n10158_not n10164_not ; n10165
g9910 and b[20]_not n10165_not ; n10166
g9911 and n9673_not quotient[27]_not ; n10167
g9912 and n9683_not n9912 ; n10168
g9913 and n9908_not n10168 ; n10169
g9914 and n9909_not n9912_not ; n10170
g9915 and n10169_not n10170_not ; n10171
g9916 and n599 n10171_not ; n10172
g9917 and n10004_not n10172 ; n10173
g9918 and n10167_not n10173_not ; n10174
g9919 and b[19]_not n10174_not ; n10175
g9920 and n9682_not quotient[27]_not ; n10176
g9921 and n9692_not n9907 ; n10177
g9922 and n9903_not n10177 ; n10178
g9923 and n9904_not n9907_not ; n10179
g9924 and n10178_not n10179_not ; n10180
g9925 and n599 n10180_not ; n10181
g9926 and n10004_not n10181 ; n10182
g9927 and n10176_not n10182_not ; n10183
g9928 and b[18]_not n10183_not ; n10184
g9929 and n9691_not quotient[27]_not ; n10185
g9930 and n9701_not n9902 ; n10186
g9931 and n9898_not n10186 ; n10187
g9932 and n9899_not n9902_not ; n10188
g9933 and n10187_not n10188_not ; n10189
g9934 and n599 n10189_not ; n10190
g9935 and n10004_not n10190 ; n10191
g9936 and n10185_not n10191_not ; n10192
g9937 and b[17]_not n10192_not ; n10193
g9938 and n9700_not quotient[27]_not ; n10194
g9939 and n9710_not n9897 ; n10195
g9940 and n9893_not n10195 ; n10196
g9941 and n9894_not n9897_not ; n10197
g9942 and n10196_not n10197_not ; n10198
g9943 and n599 n10198_not ; n10199
g9944 and n10004_not n10199 ; n10200
g9945 and n10194_not n10200_not ; n10201
g9946 and b[16]_not n10201_not ; n10202
g9947 and n9709_not quotient[27]_not ; n10203
g9948 and n9719_not n9892 ; n10204
g9949 and n9888_not n10204 ; n10205
g9950 and n9889_not n9892_not ; n10206
g9951 and n10205_not n10206_not ; n10207
g9952 and n599 n10207_not ; n10208
g9953 and n10004_not n10208 ; n10209
g9954 and n10203_not n10209_not ; n10210
g9955 and b[15]_not n10210_not ; n10211
g9956 and n9718_not quotient[27]_not ; n10212
g9957 and n9728_not n9887 ; n10213
g9958 and n9883_not n10213 ; n10214
g9959 and n9884_not n9887_not ; n10215
g9960 and n10214_not n10215_not ; n10216
g9961 and n599 n10216_not ; n10217
g9962 and n10004_not n10217 ; n10218
g9963 and n10212_not n10218_not ; n10219
g9964 and b[14]_not n10219_not ; n10220
g9965 and n9727_not quotient[27]_not ; n10221
g9966 and n9737_not n9882 ; n10222
g9967 and n9878_not n10222 ; n10223
g9968 and n9879_not n9882_not ; n10224
g9969 and n10223_not n10224_not ; n10225
g9970 and n599 n10225_not ; n10226
g9971 and n10004_not n10226 ; n10227
g9972 and n10221_not n10227_not ; n10228
g9973 and b[13]_not n10228_not ; n10229
g9974 and n9736_not quotient[27]_not ; n10230
g9975 and n9746_not n9877 ; n10231
g9976 and n9873_not n10231 ; n10232
g9977 and n9874_not n9877_not ; n10233
g9978 and n10232_not n10233_not ; n10234
g9979 and n599 n10234_not ; n10235
g9980 and n10004_not n10235 ; n10236
g9981 and n10230_not n10236_not ; n10237
g9982 and b[12]_not n10237_not ; n10238
g9983 and n9745_not quotient[27]_not ; n10239
g9984 and n9755_not n9872 ; n10240
g9985 and n9868_not n10240 ; n10241
g9986 and n9869_not n9872_not ; n10242
g9987 and n10241_not n10242_not ; n10243
g9988 and n599 n10243_not ; n10244
g9989 and n10004_not n10244 ; n10245
g9990 and n10239_not n10245_not ; n10246
g9991 and b[11]_not n10246_not ; n10247
g9992 and n9754_not quotient[27]_not ; n10248
g9993 and n9764_not n9867 ; n10249
g9994 and n9863_not n10249 ; n10250
g9995 and n9864_not n9867_not ; n10251
g9996 and n10250_not n10251_not ; n10252
g9997 and n599 n10252_not ; n10253
g9998 and n10004_not n10253 ; n10254
g9999 and n10248_not n10254_not ; n10255
g10000 and b[10]_not n10255_not ; n10256
g10001 and n9763_not quotient[27]_not ; n10257
g10002 and n9773_not n9862 ; n10258
g10003 and n9858_not n10258 ; n10259
g10004 and n9859_not n9862_not ; n10260
g10005 and n10259_not n10260_not ; n10261
g10006 and n599 n10261_not ; n10262
g10007 and n10004_not n10262 ; n10263
g10008 and n10257_not n10263_not ; n10264
g10009 and b[9]_not n10264_not ; n10265
g10010 and n9772_not quotient[27]_not ; n10266
g10011 and n9782_not n9857 ; n10267
g10012 and n9853_not n10267 ; n10268
g10013 and n9854_not n9857_not ; n10269
g10014 and n10268_not n10269_not ; n10270
g10015 and n599 n10270_not ; n10271
g10016 and n10004_not n10271 ; n10272
g10017 and n10266_not n10272_not ; n10273
g10018 and b[8]_not n10273_not ; n10274
g10019 and n9781_not quotient[27]_not ; n10275
g10020 and n9791_not n9852 ; n10276
g10021 and n9848_not n10276 ; n10277
g10022 and n9849_not n9852_not ; n10278
g10023 and n10277_not n10278_not ; n10279
g10024 and n599 n10279_not ; n10280
g10025 and n10004_not n10280 ; n10281
g10026 and n10275_not n10281_not ; n10282
g10027 and b[7]_not n10282_not ; n10283
g10028 and n9790_not quotient[27]_not ; n10284
g10029 and n9800_not n9847 ; n10285
g10030 and n9843_not n10285 ; n10286
g10031 and n9844_not n9847_not ; n10287
g10032 and n10286_not n10287_not ; n10288
g10033 and n599 n10288_not ; n10289
g10034 and n10004_not n10289 ; n10290
g10035 and n10284_not n10290_not ; n10291
g10036 and b[6]_not n10291_not ; n10292
g10037 and n9799_not quotient[27]_not ; n10293
g10038 and n9809_not n9842 ; n10294
g10039 and n9838_not n10294 ; n10295
g10040 and n9839_not n9842_not ; n10296
g10041 and n10295_not n10296_not ; n10297
g10042 and n599 n10297_not ; n10298
g10043 and n10004_not n10298 ; n10299
g10044 and n10293_not n10299_not ; n10300
g10045 and b[5]_not n10300_not ; n10301
g10046 and n9808_not quotient[27]_not ; n10302
g10047 and n9817_not n9837 ; n10303
g10048 and n9833_not n10303 ; n10304
g10049 and n9834_not n9837_not ; n10305
g10050 and n10304_not n10305_not ; n10306
g10051 and n599 n10306_not ; n10307
g10052 and n10004_not n10307 ; n10308
g10053 and n10302_not n10308_not ; n10309
g10054 and b[4]_not n10309_not ; n10310
g10055 and n9816_not quotient[27]_not ; n10311
g10056 and n9828_not n9832 ; n10312
g10057 and n9827_not n10312 ; n10313
g10058 and n9829_not n9832_not ; n10314
g10059 and n10313_not n10314_not ; n10315
g10060 and n599 n10315_not ; n10316
g10061 and n10004_not n10316 ; n10317
g10062 and n10311_not n10317_not ; n10318
g10063 and b[3]_not n10318_not ; n10319
g10064 and n9821_not quotient[27]_not ; n10320
g10065 and n9824_not n9826 ; n10321
g10066 and n9822_not n10321 ; n10322
g10067 and n599 n10322_not ; n10323
g10068 and n9827_not n10323 ; n10324
g10069 and n10004_not n10324 ; n10325
g10070 and n10320_not n10325_not ; n10326
g10071 and b[2]_not n10326_not ; n10327
g10072 and b[0] b[37]_not ; n10328
g10073 and n293 n10328 ; n10329
g10074 and n291 n10329 ; n10330
g10075 and n302 n10330 ; n10331
g10076 and n288 n10331 ; n10332
g10077 and n10004_not n10332 ; n10333
g10078 and a[27] n10333_not ; n10334
g10079 and n411 n9826 ; n10335
g10080 and n422 n10335 ; n10336
g10081 and n408 n10336 ; n10337
g10082 and n10004_not n10337 ; n10338
g10083 and n10334_not n10338_not ; n10339
g10084 and b[1] n10339_not ; n10340
g10085 and b[1]_not n10338_not ; n10341
g10086 and n10334_not n10341 ; n10342
g10087 and n10340_not n10342_not ; n10343
g10088 and a[26]_not b[0] ; n10344
g10089 and n10343_not n10344_not ; n10345
g10090 and b[1]_not n10339_not ; n10346
g10091 and n10345_not n10346_not ; n10347
g10092 and b[2] n10325_not ; n10348
g10093 and n10320_not n10348 ; n10349
g10094 and n10327_not n10349_not ; n10350
g10095 and n10347_not n10350 ; n10351
g10096 and n10327_not n10351_not ; n10352
g10097 and b[3] n10317_not ; n10353
g10098 and n10311_not n10353 ; n10354
g10099 and n10319_not n10354_not ; n10355
g10100 and n10352_not n10355 ; n10356
g10101 and n10319_not n10356_not ; n10357
g10102 and b[4] n10308_not ; n10358
g10103 and n10302_not n10358 ; n10359
g10104 and n10310_not n10359_not ; n10360
g10105 and n10357_not n10360 ; n10361
g10106 and n10310_not n10361_not ; n10362
g10107 and b[5] n10299_not ; n10363
g10108 and n10293_not n10363 ; n10364
g10109 and n10301_not n10364_not ; n10365
g10110 and n10362_not n10365 ; n10366
g10111 and n10301_not n10366_not ; n10367
g10112 and b[6] n10290_not ; n10368
g10113 and n10284_not n10368 ; n10369
g10114 and n10292_not n10369_not ; n10370
g10115 and n10367_not n10370 ; n10371
g10116 and n10292_not n10371_not ; n10372
g10117 and b[7] n10281_not ; n10373
g10118 and n10275_not n10373 ; n10374
g10119 and n10283_not n10374_not ; n10375
g10120 and n10372_not n10375 ; n10376
g10121 and n10283_not n10376_not ; n10377
g10122 and b[8] n10272_not ; n10378
g10123 and n10266_not n10378 ; n10379
g10124 and n10274_not n10379_not ; n10380
g10125 and n10377_not n10380 ; n10381
g10126 and n10274_not n10381_not ; n10382
g10127 and b[9] n10263_not ; n10383
g10128 and n10257_not n10383 ; n10384
g10129 and n10265_not n10384_not ; n10385
g10130 and n10382_not n10385 ; n10386
g10131 and n10265_not n10386_not ; n10387
g10132 and b[10] n10254_not ; n10388
g10133 and n10248_not n10388 ; n10389
g10134 and n10256_not n10389_not ; n10390
g10135 and n10387_not n10390 ; n10391
g10136 and n10256_not n10391_not ; n10392
g10137 and b[11] n10245_not ; n10393
g10138 and n10239_not n10393 ; n10394
g10139 and n10247_not n10394_not ; n10395
g10140 and n10392_not n10395 ; n10396
g10141 and n10247_not n10396_not ; n10397
g10142 and b[12] n10236_not ; n10398
g10143 and n10230_not n10398 ; n10399
g10144 and n10238_not n10399_not ; n10400
g10145 and n10397_not n10400 ; n10401
g10146 and n10238_not n10401_not ; n10402
g10147 and b[13] n10227_not ; n10403
g10148 and n10221_not n10403 ; n10404
g10149 and n10229_not n10404_not ; n10405
g10150 and n10402_not n10405 ; n10406
g10151 and n10229_not n10406_not ; n10407
g10152 and b[14] n10218_not ; n10408
g10153 and n10212_not n10408 ; n10409
g10154 and n10220_not n10409_not ; n10410
g10155 and n10407_not n10410 ; n10411
g10156 and n10220_not n10411_not ; n10412
g10157 and b[15] n10209_not ; n10413
g10158 and n10203_not n10413 ; n10414
g10159 and n10211_not n10414_not ; n10415
g10160 and n10412_not n10415 ; n10416
g10161 and n10211_not n10416_not ; n10417
g10162 and b[16] n10200_not ; n10418
g10163 and n10194_not n10418 ; n10419
g10164 and n10202_not n10419_not ; n10420
g10165 and n10417_not n10420 ; n10421
g10166 and n10202_not n10421_not ; n10422
g10167 and b[17] n10191_not ; n10423
g10168 and n10185_not n10423 ; n10424
g10169 and n10193_not n10424_not ; n10425
g10170 and n10422_not n10425 ; n10426
g10171 and n10193_not n10426_not ; n10427
g10172 and b[18] n10182_not ; n10428
g10173 and n10176_not n10428 ; n10429
g10174 and n10184_not n10429_not ; n10430
g10175 and n10427_not n10430 ; n10431
g10176 and n10184_not n10431_not ; n10432
g10177 and b[19] n10173_not ; n10433
g10178 and n10167_not n10433 ; n10434
g10179 and n10175_not n10434_not ; n10435
g10180 and n10432_not n10435 ; n10436
g10181 and n10175_not n10436_not ; n10437
g10182 and b[20] n10164_not ; n10438
g10183 and n10158_not n10438 ; n10439
g10184 and n10166_not n10439_not ; n10440
g10185 and n10437_not n10440 ; n10441
g10186 and n10166_not n10441_not ; n10442
g10187 and b[21] n10155_not ; n10443
g10188 and n10149_not n10443 ; n10444
g10189 and n10157_not n10444_not ; n10445
g10190 and n10442_not n10445 ; n10446
g10191 and n10157_not n10446_not ; n10447
g10192 and b[22] n10146_not ; n10448
g10193 and n10140_not n10448 ; n10449
g10194 and n10148_not n10449_not ; n10450
g10195 and n10447_not n10450 ; n10451
g10196 and n10148_not n10451_not ; n10452
g10197 and b[23] n10137_not ; n10453
g10198 and n10131_not n10453 ; n10454
g10199 and n10139_not n10454_not ; n10455
g10200 and n10452_not n10455 ; n10456
g10201 and n10139_not n10456_not ; n10457
g10202 and b[24] n10128_not ; n10458
g10203 and n10122_not n10458 ; n10459
g10204 and n10130_not n10459_not ; n10460
g10205 and n10457_not n10460 ; n10461
g10206 and n10130_not n10461_not ; n10462
g10207 and b[25] n10119_not ; n10463
g10208 and n10113_not n10463 ; n10464
g10209 and n10121_not n10464_not ; n10465
g10210 and n10462_not n10465 ; n10466
g10211 and n10121_not n10466_not ; n10467
g10212 and b[26] n10110_not ; n10468
g10213 and n10104_not n10468 ; n10469
g10214 and n10112_not n10469_not ; n10470
g10215 and n10467_not n10470 ; n10471
g10216 and n10112_not n10471_not ; n10472
g10217 and b[27] n10101_not ; n10473
g10218 and n10095_not n10473 ; n10474
g10219 and n10103_not n10474_not ; n10475
g10220 and n10472_not n10475 ; n10476
g10221 and n10103_not n10476_not ; n10477
g10222 and b[28] n10092_not ; n10478
g10223 and n10086_not n10478 ; n10479
g10224 and n10094_not n10479_not ; n10480
g10225 and n10477_not n10480 ; n10481
g10226 and n10094_not n10481_not ; n10482
g10227 and b[29] n10083_not ; n10483
g10228 and n10077_not n10483 ; n10484
g10229 and n10085_not n10484_not ; n10485
g10230 and n10482_not n10485 ; n10486
g10231 and n10085_not n10486_not ; n10487
g10232 and b[30] n10074_not ; n10488
g10233 and n10068_not n10488 ; n10489
g10234 and n10076_not n10489_not ; n10490
g10235 and n10487_not n10490 ; n10491
g10236 and n10076_not n10491_not ; n10492
g10237 and b[31] n10065_not ; n10493
g10238 and n10059_not n10493 ; n10494
g10239 and n10067_not n10494_not ; n10495
g10240 and n10492_not n10495 ; n10496
g10241 and n10067_not n10496_not ; n10497
g10242 and b[32] n10056_not ; n10498
g10243 and n10050_not n10498 ; n10499
g10244 and n10058_not n10499_not ; n10500
g10245 and n10497_not n10500 ; n10501
g10246 and n10058_not n10501_not ; n10502
g10247 and b[33] n10047_not ; n10503
g10248 and n10041_not n10503 ; n10504
g10249 and n10049_not n10504_not ; n10505
g10250 and n10502_not n10505 ; n10506
g10251 and n10049_not n10506_not ; n10507
g10252 and b[34] n10038_not ; n10508
g10253 and n10032_not n10508 ; n10509
g10254 and n10040_not n10509_not ; n10510
g10255 and n10507_not n10510 ; n10511
g10256 and n10040_not n10511_not ; n10512
g10257 and b[35] n10029_not ; n10513
g10258 and n10023_not n10513 ; n10514
g10259 and n10031_not n10514_not ; n10515
g10260 and n10512_not n10515 ; n10516
g10261 and n10031_not n10516_not ; n10517
g10262 and b[36] n10012_not ; n10518
g10263 and n10006_not n10518 ; n10519
g10264 and n10022_not n10519_not ; n10520
g10265 and n10517_not n10520 ; n10521
g10266 and n10022_not n10521_not ; n10522
g10267 and b[37] n10014_not ; n10523
g10268 and n10019_not n10523 ; n10524
g10269 and n10021_not n10524_not ; n10525
g10270 and n10522_not n10525 ; n10526
g10271 and n10021_not n10526_not ; n10527
g10272 and n291 n293 ; n10528
g10273 and n302 n10528 ; n10529
g10274 and n288 n10529 ; n10530
g10275 and n10527_not n10530 ; quotient[26]
g10276 and n10013_not quotient[26]_not ; n10532
g10277 and n10031_not n10520 ; n10533
g10278 and n10516_not n10533 ; n10534
g10279 and n10517_not n10520_not ; n10535
g10280 and n10534_not n10535_not ; n10536
g10281 and n10530 n10536_not ; n10537
g10282 and n10527_not n10537 ; n10538
g10283 and n10532_not n10538_not ; n10539
g10284 and b[37]_not n10539_not ; n10540
g10285 and n10030_not quotient[26]_not ; n10541
g10286 and n10040_not n10515 ; n10542
g10287 and n10511_not n10542 ; n10543
g10288 and n10512_not n10515_not ; n10544
g10289 and n10543_not n10544_not ; n10545
g10290 and n10530 n10545_not ; n10546
g10291 and n10527_not n10546 ; n10547
g10292 and n10541_not n10547_not ; n10548
g10293 and b[36]_not n10548_not ; n10549
g10294 and n10039_not quotient[26]_not ; n10550
g10295 and n10049_not n10510 ; n10551
g10296 and n10506_not n10551 ; n10552
g10297 and n10507_not n10510_not ; n10553
g10298 and n10552_not n10553_not ; n10554
g10299 and n10530 n10554_not ; n10555
g10300 and n10527_not n10555 ; n10556
g10301 and n10550_not n10556_not ; n10557
g10302 and b[35]_not n10557_not ; n10558
g10303 and n10048_not quotient[26]_not ; n10559
g10304 and n10058_not n10505 ; n10560
g10305 and n10501_not n10560 ; n10561
g10306 and n10502_not n10505_not ; n10562
g10307 and n10561_not n10562_not ; n10563
g10308 and n10530 n10563_not ; n10564
g10309 and n10527_not n10564 ; n10565
g10310 and n10559_not n10565_not ; n10566
g10311 and b[34]_not n10566_not ; n10567
g10312 and n10057_not quotient[26]_not ; n10568
g10313 and n10067_not n10500 ; n10569
g10314 and n10496_not n10569 ; n10570
g10315 and n10497_not n10500_not ; n10571
g10316 and n10570_not n10571_not ; n10572
g10317 and n10530 n10572_not ; n10573
g10318 and n10527_not n10573 ; n10574
g10319 and n10568_not n10574_not ; n10575
g10320 and b[33]_not n10575_not ; n10576
g10321 and n10066_not quotient[26]_not ; n10577
g10322 and n10076_not n10495 ; n10578
g10323 and n10491_not n10578 ; n10579
g10324 and n10492_not n10495_not ; n10580
g10325 and n10579_not n10580_not ; n10581
g10326 and n10530 n10581_not ; n10582
g10327 and n10527_not n10582 ; n10583
g10328 and n10577_not n10583_not ; n10584
g10329 and b[32]_not n10584_not ; n10585
g10330 and n10075_not quotient[26]_not ; n10586
g10331 and n10085_not n10490 ; n10587
g10332 and n10486_not n10587 ; n10588
g10333 and n10487_not n10490_not ; n10589
g10334 and n10588_not n10589_not ; n10590
g10335 and n10530 n10590_not ; n10591
g10336 and n10527_not n10591 ; n10592
g10337 and n10586_not n10592_not ; n10593
g10338 and b[31]_not n10593_not ; n10594
g10339 and n10084_not quotient[26]_not ; n10595
g10340 and n10094_not n10485 ; n10596
g10341 and n10481_not n10596 ; n10597
g10342 and n10482_not n10485_not ; n10598
g10343 and n10597_not n10598_not ; n10599
g10344 and n10530 n10599_not ; n10600
g10345 and n10527_not n10600 ; n10601
g10346 and n10595_not n10601_not ; n10602
g10347 and b[30]_not n10602_not ; n10603
g10348 and n10093_not quotient[26]_not ; n10604
g10349 and n10103_not n10480 ; n10605
g10350 and n10476_not n10605 ; n10606
g10351 and n10477_not n10480_not ; n10607
g10352 and n10606_not n10607_not ; n10608
g10353 and n10530 n10608_not ; n10609
g10354 and n10527_not n10609 ; n10610
g10355 and n10604_not n10610_not ; n10611
g10356 and b[29]_not n10611_not ; n10612
g10357 and n10102_not quotient[26]_not ; n10613
g10358 and n10112_not n10475 ; n10614
g10359 and n10471_not n10614 ; n10615
g10360 and n10472_not n10475_not ; n10616
g10361 and n10615_not n10616_not ; n10617
g10362 and n10530 n10617_not ; n10618
g10363 and n10527_not n10618 ; n10619
g10364 and n10613_not n10619_not ; n10620
g10365 and b[28]_not n10620_not ; n10621
g10366 and n10111_not quotient[26]_not ; n10622
g10367 and n10121_not n10470 ; n10623
g10368 and n10466_not n10623 ; n10624
g10369 and n10467_not n10470_not ; n10625
g10370 and n10624_not n10625_not ; n10626
g10371 and n10530 n10626_not ; n10627
g10372 and n10527_not n10627 ; n10628
g10373 and n10622_not n10628_not ; n10629
g10374 and b[27]_not n10629_not ; n10630
g10375 and n10120_not quotient[26]_not ; n10631
g10376 and n10130_not n10465 ; n10632
g10377 and n10461_not n10632 ; n10633
g10378 and n10462_not n10465_not ; n10634
g10379 and n10633_not n10634_not ; n10635
g10380 and n10530 n10635_not ; n10636
g10381 and n10527_not n10636 ; n10637
g10382 and n10631_not n10637_not ; n10638
g10383 and b[26]_not n10638_not ; n10639
g10384 and n10129_not quotient[26]_not ; n10640
g10385 and n10139_not n10460 ; n10641
g10386 and n10456_not n10641 ; n10642
g10387 and n10457_not n10460_not ; n10643
g10388 and n10642_not n10643_not ; n10644
g10389 and n10530 n10644_not ; n10645
g10390 and n10527_not n10645 ; n10646
g10391 and n10640_not n10646_not ; n10647
g10392 and b[25]_not n10647_not ; n10648
g10393 and n10138_not quotient[26]_not ; n10649
g10394 and n10148_not n10455 ; n10650
g10395 and n10451_not n10650 ; n10651
g10396 and n10452_not n10455_not ; n10652
g10397 and n10651_not n10652_not ; n10653
g10398 and n10530 n10653_not ; n10654
g10399 and n10527_not n10654 ; n10655
g10400 and n10649_not n10655_not ; n10656
g10401 and b[24]_not n10656_not ; n10657
g10402 and n10147_not quotient[26]_not ; n10658
g10403 and n10157_not n10450 ; n10659
g10404 and n10446_not n10659 ; n10660
g10405 and n10447_not n10450_not ; n10661
g10406 and n10660_not n10661_not ; n10662
g10407 and n10530 n10662_not ; n10663
g10408 and n10527_not n10663 ; n10664
g10409 and n10658_not n10664_not ; n10665
g10410 and b[23]_not n10665_not ; n10666
g10411 and n10156_not quotient[26]_not ; n10667
g10412 and n10166_not n10445 ; n10668
g10413 and n10441_not n10668 ; n10669
g10414 and n10442_not n10445_not ; n10670
g10415 and n10669_not n10670_not ; n10671
g10416 and n10530 n10671_not ; n10672
g10417 and n10527_not n10672 ; n10673
g10418 and n10667_not n10673_not ; n10674
g10419 and b[22]_not n10674_not ; n10675
g10420 and n10165_not quotient[26]_not ; n10676
g10421 and n10175_not n10440 ; n10677
g10422 and n10436_not n10677 ; n10678
g10423 and n10437_not n10440_not ; n10679
g10424 and n10678_not n10679_not ; n10680
g10425 and n10530 n10680_not ; n10681
g10426 and n10527_not n10681 ; n10682
g10427 and n10676_not n10682_not ; n10683
g10428 and b[21]_not n10683_not ; n10684
g10429 and n10174_not quotient[26]_not ; n10685
g10430 and n10184_not n10435 ; n10686
g10431 and n10431_not n10686 ; n10687
g10432 and n10432_not n10435_not ; n10688
g10433 and n10687_not n10688_not ; n10689
g10434 and n10530 n10689_not ; n10690
g10435 and n10527_not n10690 ; n10691
g10436 and n10685_not n10691_not ; n10692
g10437 and b[20]_not n10692_not ; n10693
g10438 and n10183_not quotient[26]_not ; n10694
g10439 and n10193_not n10430 ; n10695
g10440 and n10426_not n10695 ; n10696
g10441 and n10427_not n10430_not ; n10697
g10442 and n10696_not n10697_not ; n10698
g10443 and n10530 n10698_not ; n10699
g10444 and n10527_not n10699 ; n10700
g10445 and n10694_not n10700_not ; n10701
g10446 and b[19]_not n10701_not ; n10702
g10447 and n10192_not quotient[26]_not ; n10703
g10448 and n10202_not n10425 ; n10704
g10449 and n10421_not n10704 ; n10705
g10450 and n10422_not n10425_not ; n10706
g10451 and n10705_not n10706_not ; n10707
g10452 and n10530 n10707_not ; n10708
g10453 and n10527_not n10708 ; n10709
g10454 and n10703_not n10709_not ; n10710
g10455 and b[18]_not n10710_not ; n10711
g10456 and n10201_not quotient[26]_not ; n10712
g10457 and n10211_not n10420 ; n10713
g10458 and n10416_not n10713 ; n10714
g10459 and n10417_not n10420_not ; n10715
g10460 and n10714_not n10715_not ; n10716
g10461 and n10530 n10716_not ; n10717
g10462 and n10527_not n10717 ; n10718
g10463 and n10712_not n10718_not ; n10719
g10464 and b[17]_not n10719_not ; n10720
g10465 and n10210_not quotient[26]_not ; n10721
g10466 and n10220_not n10415 ; n10722
g10467 and n10411_not n10722 ; n10723
g10468 and n10412_not n10415_not ; n10724
g10469 and n10723_not n10724_not ; n10725
g10470 and n10530 n10725_not ; n10726
g10471 and n10527_not n10726 ; n10727
g10472 and n10721_not n10727_not ; n10728
g10473 and b[16]_not n10728_not ; n10729
g10474 and n10219_not quotient[26]_not ; n10730
g10475 and n10229_not n10410 ; n10731
g10476 and n10406_not n10731 ; n10732
g10477 and n10407_not n10410_not ; n10733
g10478 and n10732_not n10733_not ; n10734
g10479 and n10530 n10734_not ; n10735
g10480 and n10527_not n10735 ; n10736
g10481 and n10730_not n10736_not ; n10737
g10482 and b[15]_not n10737_not ; n10738
g10483 and n10228_not quotient[26]_not ; n10739
g10484 and n10238_not n10405 ; n10740
g10485 and n10401_not n10740 ; n10741
g10486 and n10402_not n10405_not ; n10742
g10487 and n10741_not n10742_not ; n10743
g10488 and n10530 n10743_not ; n10744
g10489 and n10527_not n10744 ; n10745
g10490 and n10739_not n10745_not ; n10746
g10491 and b[14]_not n10746_not ; n10747
g10492 and n10237_not quotient[26]_not ; n10748
g10493 and n10247_not n10400 ; n10749
g10494 and n10396_not n10749 ; n10750
g10495 and n10397_not n10400_not ; n10751
g10496 and n10750_not n10751_not ; n10752
g10497 and n10530 n10752_not ; n10753
g10498 and n10527_not n10753 ; n10754
g10499 and n10748_not n10754_not ; n10755
g10500 and b[13]_not n10755_not ; n10756
g10501 and n10246_not quotient[26]_not ; n10757
g10502 and n10256_not n10395 ; n10758
g10503 and n10391_not n10758 ; n10759
g10504 and n10392_not n10395_not ; n10760
g10505 and n10759_not n10760_not ; n10761
g10506 and n10530 n10761_not ; n10762
g10507 and n10527_not n10762 ; n10763
g10508 and n10757_not n10763_not ; n10764
g10509 and b[12]_not n10764_not ; n10765
g10510 and n10255_not quotient[26]_not ; n10766
g10511 and n10265_not n10390 ; n10767
g10512 and n10386_not n10767 ; n10768
g10513 and n10387_not n10390_not ; n10769
g10514 and n10768_not n10769_not ; n10770
g10515 and n10530 n10770_not ; n10771
g10516 and n10527_not n10771 ; n10772
g10517 and n10766_not n10772_not ; n10773
g10518 and b[11]_not n10773_not ; n10774
g10519 and n10264_not quotient[26]_not ; n10775
g10520 and n10274_not n10385 ; n10776
g10521 and n10381_not n10776 ; n10777
g10522 and n10382_not n10385_not ; n10778
g10523 and n10777_not n10778_not ; n10779
g10524 and n10530 n10779_not ; n10780
g10525 and n10527_not n10780 ; n10781
g10526 and n10775_not n10781_not ; n10782
g10527 and b[10]_not n10782_not ; n10783
g10528 and n10273_not quotient[26]_not ; n10784
g10529 and n10283_not n10380 ; n10785
g10530 and n10376_not n10785 ; n10786
g10531 and n10377_not n10380_not ; n10787
g10532 and n10786_not n10787_not ; n10788
g10533 and n10530 n10788_not ; n10789
g10534 and n10527_not n10789 ; n10790
g10535 and n10784_not n10790_not ; n10791
g10536 and b[9]_not n10791_not ; n10792
g10537 and n10282_not quotient[26]_not ; n10793
g10538 and n10292_not n10375 ; n10794
g10539 and n10371_not n10794 ; n10795
g10540 and n10372_not n10375_not ; n10796
g10541 and n10795_not n10796_not ; n10797
g10542 and n10530 n10797_not ; n10798
g10543 and n10527_not n10798 ; n10799
g10544 and n10793_not n10799_not ; n10800
g10545 and b[8]_not n10800_not ; n10801
g10546 and n10291_not quotient[26]_not ; n10802
g10547 and n10301_not n10370 ; n10803
g10548 and n10366_not n10803 ; n10804
g10549 and n10367_not n10370_not ; n10805
g10550 and n10804_not n10805_not ; n10806
g10551 and n10530 n10806_not ; n10807
g10552 and n10527_not n10807 ; n10808
g10553 and n10802_not n10808_not ; n10809
g10554 and b[7]_not n10809_not ; n10810
g10555 and n10300_not quotient[26]_not ; n10811
g10556 and n10310_not n10365 ; n10812
g10557 and n10361_not n10812 ; n10813
g10558 and n10362_not n10365_not ; n10814
g10559 and n10813_not n10814_not ; n10815
g10560 and n10530 n10815_not ; n10816
g10561 and n10527_not n10816 ; n10817
g10562 and n10811_not n10817_not ; n10818
g10563 and b[6]_not n10818_not ; n10819
g10564 and n10309_not quotient[26]_not ; n10820
g10565 and n10319_not n10360 ; n10821
g10566 and n10356_not n10821 ; n10822
g10567 and n10357_not n10360_not ; n10823
g10568 and n10822_not n10823_not ; n10824
g10569 and n10530 n10824_not ; n10825
g10570 and n10527_not n10825 ; n10826
g10571 and n10820_not n10826_not ; n10827
g10572 and b[5]_not n10827_not ; n10828
g10573 and n10318_not quotient[26]_not ; n10829
g10574 and n10327_not n10355 ; n10830
g10575 and n10351_not n10830 ; n10831
g10576 and n10352_not n10355_not ; n10832
g10577 and n10831_not n10832_not ; n10833
g10578 and n10530 n10833_not ; n10834
g10579 and n10527_not n10834 ; n10835
g10580 and n10829_not n10835_not ; n10836
g10581 and b[4]_not n10836_not ; n10837
g10582 and n10326_not quotient[26]_not ; n10838
g10583 and n10346_not n10350 ; n10839
g10584 and n10345_not n10839 ; n10840
g10585 and n10347_not n10350_not ; n10841
g10586 and n10840_not n10841_not ; n10842
g10587 and n10530 n10842_not ; n10843
g10588 and n10527_not n10843 ; n10844
g10589 and n10838_not n10844_not ; n10845
g10590 and b[3]_not n10845_not ; n10846
g10591 and n10339_not quotient[26]_not ; n10847
g10592 and n10342_not n10344 ; n10848
g10593 and n10340_not n10848 ; n10849
g10594 and n10530 n10849_not ; n10850
g10595 and n10345_not n10850 ; n10851
g10596 and n10527_not n10851 ; n10852
g10597 and n10847_not n10852_not ; n10853
g10598 and b[2]_not n10853_not ; n10854
g10599 and b[0] b[38]_not ; n10855
g10600 and n410 n10855 ; n10856
g10601 and n421 n10856 ; n10857
g10602 and n597 n10857 ; n10858
g10603 and n595 n10858 ; n10859
g10604 and n10527_not n10859 ; n10860
g10605 and a[26] n10860_not ; n10861
g10606 and n293 n10344 ; n10862
g10607 and n291 n10862 ; n10863
g10608 and n302 n10863 ; n10864
g10609 and n288 n10864 ; n10865
g10610 and n10527_not n10865 ; n10866
g10611 and n10861_not n10866_not ; n10867
g10612 and b[1] n10867_not ; n10868
g10613 and b[1]_not n10866_not ; n10869
g10614 and n10861_not n10869 ; n10870
g10615 and n10868_not n10870_not ; n10871
g10616 and a[25]_not b[0] ; n10872
g10617 and n10871_not n10872_not ; n10873
g10618 and b[1]_not n10867_not ; n10874
g10619 and n10873_not n10874_not ; n10875
g10620 and b[2] n10852_not ; n10876
g10621 and n10847_not n10876 ; n10877
g10622 and n10854_not n10877_not ; n10878
g10623 and n10875_not n10878 ; n10879
g10624 and n10854_not n10879_not ; n10880
g10625 and b[3] n10844_not ; n10881
g10626 and n10838_not n10881 ; n10882
g10627 and n10846_not n10882_not ; n10883
g10628 and n10880_not n10883 ; n10884
g10629 and n10846_not n10884_not ; n10885
g10630 and b[4] n10835_not ; n10886
g10631 and n10829_not n10886 ; n10887
g10632 and n10837_not n10887_not ; n10888
g10633 and n10885_not n10888 ; n10889
g10634 and n10837_not n10889_not ; n10890
g10635 and b[5] n10826_not ; n10891
g10636 and n10820_not n10891 ; n10892
g10637 and n10828_not n10892_not ; n10893
g10638 and n10890_not n10893 ; n10894
g10639 and n10828_not n10894_not ; n10895
g10640 and b[6] n10817_not ; n10896
g10641 and n10811_not n10896 ; n10897
g10642 and n10819_not n10897_not ; n10898
g10643 and n10895_not n10898 ; n10899
g10644 and n10819_not n10899_not ; n10900
g10645 and b[7] n10808_not ; n10901
g10646 and n10802_not n10901 ; n10902
g10647 and n10810_not n10902_not ; n10903
g10648 and n10900_not n10903 ; n10904
g10649 and n10810_not n10904_not ; n10905
g10650 and b[8] n10799_not ; n10906
g10651 and n10793_not n10906 ; n10907
g10652 and n10801_not n10907_not ; n10908
g10653 and n10905_not n10908 ; n10909
g10654 and n10801_not n10909_not ; n10910
g10655 and b[9] n10790_not ; n10911
g10656 and n10784_not n10911 ; n10912
g10657 and n10792_not n10912_not ; n10913
g10658 and n10910_not n10913 ; n10914
g10659 and n10792_not n10914_not ; n10915
g10660 and b[10] n10781_not ; n10916
g10661 and n10775_not n10916 ; n10917
g10662 and n10783_not n10917_not ; n10918
g10663 and n10915_not n10918 ; n10919
g10664 and n10783_not n10919_not ; n10920
g10665 and b[11] n10772_not ; n10921
g10666 and n10766_not n10921 ; n10922
g10667 and n10774_not n10922_not ; n10923
g10668 and n10920_not n10923 ; n10924
g10669 and n10774_not n10924_not ; n10925
g10670 and b[12] n10763_not ; n10926
g10671 and n10757_not n10926 ; n10927
g10672 and n10765_not n10927_not ; n10928
g10673 and n10925_not n10928 ; n10929
g10674 and n10765_not n10929_not ; n10930
g10675 and b[13] n10754_not ; n10931
g10676 and n10748_not n10931 ; n10932
g10677 and n10756_not n10932_not ; n10933
g10678 and n10930_not n10933 ; n10934
g10679 and n10756_not n10934_not ; n10935
g10680 and b[14] n10745_not ; n10936
g10681 and n10739_not n10936 ; n10937
g10682 and n10747_not n10937_not ; n10938
g10683 and n10935_not n10938 ; n10939
g10684 and n10747_not n10939_not ; n10940
g10685 and b[15] n10736_not ; n10941
g10686 and n10730_not n10941 ; n10942
g10687 and n10738_not n10942_not ; n10943
g10688 and n10940_not n10943 ; n10944
g10689 and n10738_not n10944_not ; n10945
g10690 and b[16] n10727_not ; n10946
g10691 and n10721_not n10946 ; n10947
g10692 and n10729_not n10947_not ; n10948
g10693 and n10945_not n10948 ; n10949
g10694 and n10729_not n10949_not ; n10950
g10695 and b[17] n10718_not ; n10951
g10696 and n10712_not n10951 ; n10952
g10697 and n10720_not n10952_not ; n10953
g10698 and n10950_not n10953 ; n10954
g10699 and n10720_not n10954_not ; n10955
g10700 and b[18] n10709_not ; n10956
g10701 and n10703_not n10956 ; n10957
g10702 and n10711_not n10957_not ; n10958
g10703 and n10955_not n10958 ; n10959
g10704 and n10711_not n10959_not ; n10960
g10705 and b[19] n10700_not ; n10961
g10706 and n10694_not n10961 ; n10962
g10707 and n10702_not n10962_not ; n10963
g10708 and n10960_not n10963 ; n10964
g10709 and n10702_not n10964_not ; n10965
g10710 and b[20] n10691_not ; n10966
g10711 and n10685_not n10966 ; n10967
g10712 and n10693_not n10967_not ; n10968
g10713 and n10965_not n10968 ; n10969
g10714 and n10693_not n10969_not ; n10970
g10715 and b[21] n10682_not ; n10971
g10716 and n10676_not n10971 ; n10972
g10717 and n10684_not n10972_not ; n10973
g10718 and n10970_not n10973 ; n10974
g10719 and n10684_not n10974_not ; n10975
g10720 and b[22] n10673_not ; n10976
g10721 and n10667_not n10976 ; n10977
g10722 and n10675_not n10977_not ; n10978
g10723 and n10975_not n10978 ; n10979
g10724 and n10675_not n10979_not ; n10980
g10725 and b[23] n10664_not ; n10981
g10726 and n10658_not n10981 ; n10982
g10727 and n10666_not n10982_not ; n10983
g10728 and n10980_not n10983 ; n10984
g10729 and n10666_not n10984_not ; n10985
g10730 and b[24] n10655_not ; n10986
g10731 and n10649_not n10986 ; n10987
g10732 and n10657_not n10987_not ; n10988
g10733 and n10985_not n10988 ; n10989
g10734 and n10657_not n10989_not ; n10990
g10735 and b[25] n10646_not ; n10991
g10736 and n10640_not n10991 ; n10992
g10737 and n10648_not n10992_not ; n10993
g10738 and n10990_not n10993 ; n10994
g10739 and n10648_not n10994_not ; n10995
g10740 and b[26] n10637_not ; n10996
g10741 and n10631_not n10996 ; n10997
g10742 and n10639_not n10997_not ; n10998
g10743 and n10995_not n10998 ; n10999
g10744 and n10639_not n10999_not ; n11000
g10745 and b[27] n10628_not ; n11001
g10746 and n10622_not n11001 ; n11002
g10747 and n10630_not n11002_not ; n11003
g10748 and n11000_not n11003 ; n11004
g10749 and n10630_not n11004_not ; n11005
g10750 and b[28] n10619_not ; n11006
g10751 and n10613_not n11006 ; n11007
g10752 and n10621_not n11007_not ; n11008
g10753 and n11005_not n11008 ; n11009
g10754 and n10621_not n11009_not ; n11010
g10755 and b[29] n10610_not ; n11011
g10756 and n10604_not n11011 ; n11012
g10757 and n10612_not n11012_not ; n11013
g10758 and n11010_not n11013 ; n11014
g10759 and n10612_not n11014_not ; n11015
g10760 and b[30] n10601_not ; n11016
g10761 and n10595_not n11016 ; n11017
g10762 and n10603_not n11017_not ; n11018
g10763 and n11015_not n11018 ; n11019
g10764 and n10603_not n11019_not ; n11020
g10765 and b[31] n10592_not ; n11021
g10766 and n10586_not n11021 ; n11022
g10767 and n10594_not n11022_not ; n11023
g10768 and n11020_not n11023 ; n11024
g10769 and n10594_not n11024_not ; n11025
g10770 and b[32] n10583_not ; n11026
g10771 and n10577_not n11026 ; n11027
g10772 and n10585_not n11027_not ; n11028
g10773 and n11025_not n11028 ; n11029
g10774 and n10585_not n11029_not ; n11030
g10775 and b[33] n10574_not ; n11031
g10776 and n10568_not n11031 ; n11032
g10777 and n10576_not n11032_not ; n11033
g10778 and n11030_not n11033 ; n11034
g10779 and n10576_not n11034_not ; n11035
g10780 and b[34] n10565_not ; n11036
g10781 and n10559_not n11036 ; n11037
g10782 and n10567_not n11037_not ; n11038
g10783 and n11035_not n11038 ; n11039
g10784 and n10567_not n11039_not ; n11040
g10785 and b[35] n10556_not ; n11041
g10786 and n10550_not n11041 ; n11042
g10787 and n10558_not n11042_not ; n11043
g10788 and n11040_not n11043 ; n11044
g10789 and n10558_not n11044_not ; n11045
g10790 and b[36] n10547_not ; n11046
g10791 and n10541_not n11046 ; n11047
g10792 and n10549_not n11047_not ; n11048
g10793 and n11045_not n11048 ; n11049
g10794 and n10549_not n11049_not ; n11050
g10795 and b[37] n10538_not ; n11051
g10796 and n10532_not n11051 ; n11052
g10797 and n10540_not n11052_not ; n11053
g10798 and n11050_not n11053 ; n11054
g10799 and n10540_not n11054_not ; n11055
g10800 and n10020_not quotient[26]_not ; n11056
g10801 and n10022_not n10525 ; n11057
g10802 and n10521_not n11057 ; n11058
g10803 and n10522_not n10525_not ; n11059
g10804 and n11058_not n11059_not ; n11060
g10805 and quotient[26] n11060_not ; n11061
g10806 and n11056_not n11061_not ; n11062
g10807 and b[38]_not n11062_not ; n11063
g10808 and b[38] n11056_not ; n11064
g10809 and n11061_not n11064 ; n11065
g10810 and n410 n421 ; n11066
g10811 and n597 n11066 ; n11067
g10812 and n595 n11067 ; n11068
g10813 and n11065_not n11068 ; n11069
g10814 and n11063_not n11069 ; n11070
g10815 and n11055_not n11070 ; n11071
g10816 and n10530 n11062_not ; n11072
g10817 and n11071_not n11072_not ; quotient[25]
g10818 and n10549_not n11053 ; n11074
g10819 and n11049_not n11074 ; n11075
g10820 and n11050_not n11053_not ; n11076
g10821 and n11075_not n11076_not ; n11077
g10822 and quotient[25] n11077_not ; n11078
g10823 and n10539_not n11072_not ; n11079
g10824 and n11071_not n11079 ; n11080
g10825 and n11078_not n11080_not ; n11081
g10826 and n10540_not n11065_not ; n11082
g10827 and n11063_not n11082 ; n11083
g10828 and n11054_not n11083 ; n11084
g10829 and n11063_not n11065_not ; n11085
g10830 and n11055_not n11085_not ; n11086
g10831 and n11084_not n11086_not ; n11087
g10832 and quotient[25] n11087_not ; n11088
g10833 and n11062_not n11072_not ; n11089
g10834 and n11071_not n11089 ; n11090
g10835 and n11088_not n11090_not ; n11091
g10836 and b[39]_not n11091_not ; n11092
g10837 and b[38]_not n11081_not ; n11093
g10838 and n10558_not n11048 ; n11094
g10839 and n11044_not n11094 ; n11095
g10840 and n11045_not n11048_not ; n11096
g10841 and n11095_not n11096_not ; n11097
g10842 and quotient[25] n11097_not ; n11098
g10843 and n10548_not n11072_not ; n11099
g10844 and n11071_not n11099 ; n11100
g10845 and n11098_not n11100_not ; n11101
g10846 and b[37]_not n11101_not ; n11102
g10847 and n10567_not n11043 ; n11103
g10848 and n11039_not n11103 ; n11104
g10849 and n11040_not n11043_not ; n11105
g10850 and n11104_not n11105_not ; n11106
g10851 and quotient[25] n11106_not ; n11107
g10852 and n10557_not n11072_not ; n11108
g10853 and n11071_not n11108 ; n11109
g10854 and n11107_not n11109_not ; n11110
g10855 and b[36]_not n11110_not ; n11111
g10856 and n10576_not n11038 ; n11112
g10857 and n11034_not n11112 ; n11113
g10858 and n11035_not n11038_not ; n11114
g10859 and n11113_not n11114_not ; n11115
g10860 and quotient[25] n11115_not ; n11116
g10861 and n10566_not n11072_not ; n11117
g10862 and n11071_not n11117 ; n11118
g10863 and n11116_not n11118_not ; n11119
g10864 and b[35]_not n11119_not ; n11120
g10865 and n10585_not n11033 ; n11121
g10866 and n11029_not n11121 ; n11122
g10867 and n11030_not n11033_not ; n11123
g10868 and n11122_not n11123_not ; n11124
g10869 and quotient[25] n11124_not ; n11125
g10870 and n10575_not n11072_not ; n11126
g10871 and n11071_not n11126 ; n11127
g10872 and n11125_not n11127_not ; n11128
g10873 and b[34]_not n11128_not ; n11129
g10874 and n10594_not n11028 ; n11130
g10875 and n11024_not n11130 ; n11131
g10876 and n11025_not n11028_not ; n11132
g10877 and n11131_not n11132_not ; n11133
g10878 and quotient[25] n11133_not ; n11134
g10879 and n10584_not n11072_not ; n11135
g10880 and n11071_not n11135 ; n11136
g10881 and n11134_not n11136_not ; n11137
g10882 and b[33]_not n11137_not ; n11138
g10883 and n10603_not n11023 ; n11139
g10884 and n11019_not n11139 ; n11140
g10885 and n11020_not n11023_not ; n11141
g10886 and n11140_not n11141_not ; n11142
g10887 and quotient[25] n11142_not ; n11143
g10888 and n10593_not n11072_not ; n11144
g10889 and n11071_not n11144 ; n11145
g10890 and n11143_not n11145_not ; n11146
g10891 and b[32]_not n11146_not ; n11147
g10892 and n10612_not n11018 ; n11148
g10893 and n11014_not n11148 ; n11149
g10894 and n11015_not n11018_not ; n11150
g10895 and n11149_not n11150_not ; n11151
g10896 and quotient[25] n11151_not ; n11152
g10897 and n10602_not n11072_not ; n11153
g10898 and n11071_not n11153 ; n11154
g10899 and n11152_not n11154_not ; n11155
g10900 and b[31]_not n11155_not ; n11156
g10901 and n10621_not n11013 ; n11157
g10902 and n11009_not n11157 ; n11158
g10903 and n11010_not n11013_not ; n11159
g10904 and n11158_not n11159_not ; n11160
g10905 and quotient[25] n11160_not ; n11161
g10906 and n10611_not n11072_not ; n11162
g10907 and n11071_not n11162 ; n11163
g10908 and n11161_not n11163_not ; n11164
g10909 and b[30]_not n11164_not ; n11165
g10910 and n10630_not n11008 ; n11166
g10911 and n11004_not n11166 ; n11167
g10912 and n11005_not n11008_not ; n11168
g10913 and n11167_not n11168_not ; n11169
g10914 and quotient[25] n11169_not ; n11170
g10915 and n10620_not n11072_not ; n11171
g10916 and n11071_not n11171 ; n11172
g10917 and n11170_not n11172_not ; n11173
g10918 and b[29]_not n11173_not ; n11174
g10919 and n10639_not n11003 ; n11175
g10920 and n10999_not n11175 ; n11176
g10921 and n11000_not n11003_not ; n11177
g10922 and n11176_not n11177_not ; n11178
g10923 and quotient[25] n11178_not ; n11179
g10924 and n10629_not n11072_not ; n11180
g10925 and n11071_not n11180 ; n11181
g10926 and n11179_not n11181_not ; n11182
g10927 and b[28]_not n11182_not ; n11183
g10928 and n10648_not n10998 ; n11184
g10929 and n10994_not n11184 ; n11185
g10930 and n10995_not n10998_not ; n11186
g10931 and n11185_not n11186_not ; n11187
g10932 and quotient[25] n11187_not ; n11188
g10933 and n10638_not n11072_not ; n11189
g10934 and n11071_not n11189 ; n11190
g10935 and n11188_not n11190_not ; n11191
g10936 and b[27]_not n11191_not ; n11192
g10937 and n10657_not n10993 ; n11193
g10938 and n10989_not n11193 ; n11194
g10939 and n10990_not n10993_not ; n11195
g10940 and n11194_not n11195_not ; n11196
g10941 and quotient[25] n11196_not ; n11197
g10942 and n10647_not n11072_not ; n11198
g10943 and n11071_not n11198 ; n11199
g10944 and n11197_not n11199_not ; n11200
g10945 and b[26]_not n11200_not ; n11201
g10946 and n10666_not n10988 ; n11202
g10947 and n10984_not n11202 ; n11203
g10948 and n10985_not n10988_not ; n11204
g10949 and n11203_not n11204_not ; n11205
g10950 and quotient[25] n11205_not ; n11206
g10951 and n10656_not n11072_not ; n11207
g10952 and n11071_not n11207 ; n11208
g10953 and n11206_not n11208_not ; n11209
g10954 and b[25]_not n11209_not ; n11210
g10955 and n10675_not n10983 ; n11211
g10956 and n10979_not n11211 ; n11212
g10957 and n10980_not n10983_not ; n11213
g10958 and n11212_not n11213_not ; n11214
g10959 and quotient[25] n11214_not ; n11215
g10960 and n10665_not n11072_not ; n11216
g10961 and n11071_not n11216 ; n11217
g10962 and n11215_not n11217_not ; n11218
g10963 and b[24]_not n11218_not ; n11219
g10964 and n10684_not n10978 ; n11220
g10965 and n10974_not n11220 ; n11221
g10966 and n10975_not n10978_not ; n11222
g10967 and n11221_not n11222_not ; n11223
g10968 and quotient[25] n11223_not ; n11224
g10969 and n10674_not n11072_not ; n11225
g10970 and n11071_not n11225 ; n11226
g10971 and n11224_not n11226_not ; n11227
g10972 and b[23]_not n11227_not ; n11228
g10973 and n10693_not n10973 ; n11229
g10974 and n10969_not n11229 ; n11230
g10975 and n10970_not n10973_not ; n11231
g10976 and n11230_not n11231_not ; n11232
g10977 and quotient[25] n11232_not ; n11233
g10978 and n10683_not n11072_not ; n11234
g10979 and n11071_not n11234 ; n11235
g10980 and n11233_not n11235_not ; n11236
g10981 and b[22]_not n11236_not ; n11237
g10982 and n10702_not n10968 ; n11238
g10983 and n10964_not n11238 ; n11239
g10984 and n10965_not n10968_not ; n11240
g10985 and n11239_not n11240_not ; n11241
g10986 and quotient[25] n11241_not ; n11242
g10987 and n10692_not n11072_not ; n11243
g10988 and n11071_not n11243 ; n11244
g10989 and n11242_not n11244_not ; n11245
g10990 and b[21]_not n11245_not ; n11246
g10991 and n10711_not n10963 ; n11247
g10992 and n10959_not n11247 ; n11248
g10993 and n10960_not n10963_not ; n11249
g10994 and n11248_not n11249_not ; n11250
g10995 and quotient[25] n11250_not ; n11251
g10996 and n10701_not n11072_not ; n11252
g10997 and n11071_not n11252 ; n11253
g10998 and n11251_not n11253_not ; n11254
g10999 and b[20]_not n11254_not ; n11255
g11000 and n10720_not n10958 ; n11256
g11001 and n10954_not n11256 ; n11257
g11002 and n10955_not n10958_not ; n11258
g11003 and n11257_not n11258_not ; n11259
g11004 and quotient[25] n11259_not ; n11260
g11005 and n10710_not n11072_not ; n11261
g11006 and n11071_not n11261 ; n11262
g11007 and n11260_not n11262_not ; n11263
g11008 and b[19]_not n11263_not ; n11264
g11009 and n10729_not n10953 ; n11265
g11010 and n10949_not n11265 ; n11266
g11011 and n10950_not n10953_not ; n11267
g11012 and n11266_not n11267_not ; n11268
g11013 and quotient[25] n11268_not ; n11269
g11014 and n10719_not n11072_not ; n11270
g11015 and n11071_not n11270 ; n11271
g11016 and n11269_not n11271_not ; n11272
g11017 and b[18]_not n11272_not ; n11273
g11018 and n10738_not n10948 ; n11274
g11019 and n10944_not n11274 ; n11275
g11020 and n10945_not n10948_not ; n11276
g11021 and n11275_not n11276_not ; n11277
g11022 and quotient[25] n11277_not ; n11278
g11023 and n10728_not n11072_not ; n11279
g11024 and n11071_not n11279 ; n11280
g11025 and n11278_not n11280_not ; n11281
g11026 and b[17]_not n11281_not ; n11282
g11027 and n10747_not n10943 ; n11283
g11028 and n10939_not n11283 ; n11284
g11029 and n10940_not n10943_not ; n11285
g11030 and n11284_not n11285_not ; n11286
g11031 and quotient[25] n11286_not ; n11287
g11032 and n10737_not n11072_not ; n11288
g11033 and n11071_not n11288 ; n11289
g11034 and n11287_not n11289_not ; n11290
g11035 and b[16]_not n11290_not ; n11291
g11036 and n10756_not n10938 ; n11292
g11037 and n10934_not n11292 ; n11293
g11038 and n10935_not n10938_not ; n11294
g11039 and n11293_not n11294_not ; n11295
g11040 and quotient[25] n11295_not ; n11296
g11041 and n10746_not n11072_not ; n11297
g11042 and n11071_not n11297 ; n11298
g11043 and n11296_not n11298_not ; n11299
g11044 and b[15]_not n11299_not ; n11300
g11045 and n10765_not n10933 ; n11301
g11046 and n10929_not n11301 ; n11302
g11047 and n10930_not n10933_not ; n11303
g11048 and n11302_not n11303_not ; n11304
g11049 and quotient[25] n11304_not ; n11305
g11050 and n10755_not n11072_not ; n11306
g11051 and n11071_not n11306 ; n11307
g11052 and n11305_not n11307_not ; n11308
g11053 and b[14]_not n11308_not ; n11309
g11054 and n10774_not n10928 ; n11310
g11055 and n10924_not n11310 ; n11311
g11056 and n10925_not n10928_not ; n11312
g11057 and n11311_not n11312_not ; n11313
g11058 and quotient[25] n11313_not ; n11314
g11059 and n10764_not n11072_not ; n11315
g11060 and n11071_not n11315 ; n11316
g11061 and n11314_not n11316_not ; n11317
g11062 and b[13]_not n11317_not ; n11318
g11063 and n10783_not n10923 ; n11319
g11064 and n10919_not n11319 ; n11320
g11065 and n10920_not n10923_not ; n11321
g11066 and n11320_not n11321_not ; n11322
g11067 and quotient[25] n11322_not ; n11323
g11068 and n10773_not n11072_not ; n11324
g11069 and n11071_not n11324 ; n11325
g11070 and n11323_not n11325_not ; n11326
g11071 and b[12]_not n11326_not ; n11327
g11072 and n10792_not n10918 ; n11328
g11073 and n10914_not n11328 ; n11329
g11074 and n10915_not n10918_not ; n11330
g11075 and n11329_not n11330_not ; n11331
g11076 and quotient[25] n11331_not ; n11332
g11077 and n10782_not n11072_not ; n11333
g11078 and n11071_not n11333 ; n11334
g11079 and n11332_not n11334_not ; n11335
g11080 and b[11]_not n11335_not ; n11336
g11081 and n10801_not n10913 ; n11337
g11082 and n10909_not n11337 ; n11338
g11083 and n10910_not n10913_not ; n11339
g11084 and n11338_not n11339_not ; n11340
g11085 and quotient[25] n11340_not ; n11341
g11086 and n10791_not n11072_not ; n11342
g11087 and n11071_not n11342 ; n11343
g11088 and n11341_not n11343_not ; n11344
g11089 and b[10]_not n11344_not ; n11345
g11090 and n10810_not n10908 ; n11346
g11091 and n10904_not n11346 ; n11347
g11092 and n10905_not n10908_not ; n11348
g11093 and n11347_not n11348_not ; n11349
g11094 and quotient[25] n11349_not ; n11350
g11095 and n10800_not n11072_not ; n11351
g11096 and n11071_not n11351 ; n11352
g11097 and n11350_not n11352_not ; n11353
g11098 and b[9]_not n11353_not ; n11354
g11099 and n10819_not n10903 ; n11355
g11100 and n10899_not n11355 ; n11356
g11101 and n10900_not n10903_not ; n11357
g11102 and n11356_not n11357_not ; n11358
g11103 and quotient[25] n11358_not ; n11359
g11104 and n10809_not n11072_not ; n11360
g11105 and n11071_not n11360 ; n11361
g11106 and n11359_not n11361_not ; n11362
g11107 and b[8]_not n11362_not ; n11363
g11108 and n10828_not n10898 ; n11364
g11109 and n10894_not n11364 ; n11365
g11110 and n10895_not n10898_not ; n11366
g11111 and n11365_not n11366_not ; n11367
g11112 and quotient[25] n11367_not ; n11368
g11113 and n10818_not n11072_not ; n11369
g11114 and n11071_not n11369 ; n11370
g11115 and n11368_not n11370_not ; n11371
g11116 and b[7]_not n11371_not ; n11372
g11117 and n10837_not n10893 ; n11373
g11118 and n10889_not n11373 ; n11374
g11119 and n10890_not n10893_not ; n11375
g11120 and n11374_not n11375_not ; n11376
g11121 and quotient[25] n11376_not ; n11377
g11122 and n10827_not n11072_not ; n11378
g11123 and n11071_not n11378 ; n11379
g11124 and n11377_not n11379_not ; n11380
g11125 and b[6]_not n11380_not ; n11381
g11126 and n10846_not n10888 ; n11382
g11127 and n10884_not n11382 ; n11383
g11128 and n10885_not n10888_not ; n11384
g11129 and n11383_not n11384_not ; n11385
g11130 and quotient[25] n11385_not ; n11386
g11131 and n10836_not n11072_not ; n11387
g11132 and n11071_not n11387 ; n11388
g11133 and n11386_not n11388_not ; n11389
g11134 and b[5]_not n11389_not ; n11390
g11135 and n10854_not n10883 ; n11391
g11136 and n10879_not n11391 ; n11392
g11137 and n10880_not n10883_not ; n11393
g11138 and n11392_not n11393_not ; n11394
g11139 and quotient[25] n11394_not ; n11395
g11140 and n10845_not n11072_not ; n11396
g11141 and n11071_not n11396 ; n11397
g11142 and n11395_not n11397_not ; n11398
g11143 and b[4]_not n11398_not ; n11399
g11144 and n10874_not n10878 ; n11400
g11145 and n10873_not n11400 ; n11401
g11146 and n10875_not n10878_not ; n11402
g11147 and n11401_not n11402_not ; n11403
g11148 and quotient[25] n11403_not ; n11404
g11149 and n10853_not n11072_not ; n11405
g11150 and n11071_not n11405 ; n11406
g11151 and n11404_not n11406_not ; n11407
g11152 and b[3]_not n11407_not ; n11408
g11153 and n10870_not n10872 ; n11409
g11154 and n10868_not n11409 ; n11410
g11155 and n10873_not n11410_not ; n11411
g11156 and quotient[25] n11411 ; n11412
g11157 and n10867_not n11072_not ; n11413
g11158 and n11071_not n11413 ; n11414
g11159 and n11412_not n11414_not ; n11415
g11160 and b[2]_not n11415_not ; n11416
g11161 and b[0] quotient[25] ; n11417
g11162 and a[25] n11417_not ; n11418
g11163 and n10872 quotient[25] ; n11419
g11164 and n11418_not n11419_not ; n11420
g11165 and b[1] n11420_not ; n11421
g11166 and b[1]_not n11419_not ; n11422
g11167 and n11418_not n11422 ; n11423
g11168 and n11421_not n11423_not ; n11424
g11169 and a[24]_not b[0] ; n11425
g11170 and n11424_not n11425_not ; n11426
g11171 and b[1]_not n11420_not ; n11427
g11172 and n11426_not n11427_not ; n11428
g11173 and b[2] n11414_not ; n11429
g11174 and n11412_not n11429 ; n11430
g11175 and n11416_not n11430_not ; n11431
g11176 and n11428_not n11431 ; n11432
g11177 and n11416_not n11432_not ; n11433
g11178 and b[3] n11406_not ; n11434
g11179 and n11404_not n11434 ; n11435
g11180 and n11408_not n11435_not ; n11436
g11181 and n11433_not n11436 ; n11437
g11182 and n11408_not n11437_not ; n11438
g11183 and b[4] n11397_not ; n11439
g11184 and n11395_not n11439 ; n11440
g11185 and n11399_not n11440_not ; n11441
g11186 and n11438_not n11441 ; n11442
g11187 and n11399_not n11442_not ; n11443
g11188 and b[5] n11388_not ; n11444
g11189 and n11386_not n11444 ; n11445
g11190 and n11390_not n11445_not ; n11446
g11191 and n11443_not n11446 ; n11447
g11192 and n11390_not n11447_not ; n11448
g11193 and b[6] n11379_not ; n11449
g11194 and n11377_not n11449 ; n11450
g11195 and n11381_not n11450_not ; n11451
g11196 and n11448_not n11451 ; n11452
g11197 and n11381_not n11452_not ; n11453
g11198 and b[7] n11370_not ; n11454
g11199 and n11368_not n11454 ; n11455
g11200 and n11372_not n11455_not ; n11456
g11201 and n11453_not n11456 ; n11457
g11202 and n11372_not n11457_not ; n11458
g11203 and b[8] n11361_not ; n11459
g11204 and n11359_not n11459 ; n11460
g11205 and n11363_not n11460_not ; n11461
g11206 and n11458_not n11461 ; n11462
g11207 and n11363_not n11462_not ; n11463
g11208 and b[9] n11352_not ; n11464
g11209 and n11350_not n11464 ; n11465
g11210 and n11354_not n11465_not ; n11466
g11211 and n11463_not n11466 ; n11467
g11212 and n11354_not n11467_not ; n11468
g11213 and b[10] n11343_not ; n11469
g11214 and n11341_not n11469 ; n11470
g11215 and n11345_not n11470_not ; n11471
g11216 and n11468_not n11471 ; n11472
g11217 and n11345_not n11472_not ; n11473
g11218 and b[11] n11334_not ; n11474
g11219 and n11332_not n11474 ; n11475
g11220 and n11336_not n11475_not ; n11476
g11221 and n11473_not n11476 ; n11477
g11222 and n11336_not n11477_not ; n11478
g11223 and b[12] n11325_not ; n11479
g11224 and n11323_not n11479 ; n11480
g11225 and n11327_not n11480_not ; n11481
g11226 and n11478_not n11481 ; n11482
g11227 and n11327_not n11482_not ; n11483
g11228 and b[13] n11316_not ; n11484
g11229 and n11314_not n11484 ; n11485
g11230 and n11318_not n11485_not ; n11486
g11231 and n11483_not n11486 ; n11487
g11232 and n11318_not n11487_not ; n11488
g11233 and b[14] n11307_not ; n11489
g11234 and n11305_not n11489 ; n11490
g11235 and n11309_not n11490_not ; n11491
g11236 and n11488_not n11491 ; n11492
g11237 and n11309_not n11492_not ; n11493
g11238 and b[15] n11298_not ; n11494
g11239 and n11296_not n11494 ; n11495
g11240 and n11300_not n11495_not ; n11496
g11241 and n11493_not n11496 ; n11497
g11242 and n11300_not n11497_not ; n11498
g11243 and b[16] n11289_not ; n11499
g11244 and n11287_not n11499 ; n11500
g11245 and n11291_not n11500_not ; n11501
g11246 and n11498_not n11501 ; n11502
g11247 and n11291_not n11502_not ; n11503
g11248 and b[17] n11280_not ; n11504
g11249 and n11278_not n11504 ; n11505
g11250 and n11282_not n11505_not ; n11506
g11251 and n11503_not n11506 ; n11507
g11252 and n11282_not n11507_not ; n11508
g11253 and b[18] n11271_not ; n11509
g11254 and n11269_not n11509 ; n11510
g11255 and n11273_not n11510_not ; n11511
g11256 and n11508_not n11511 ; n11512
g11257 and n11273_not n11512_not ; n11513
g11258 and b[19] n11262_not ; n11514
g11259 and n11260_not n11514 ; n11515
g11260 and n11264_not n11515_not ; n11516
g11261 and n11513_not n11516 ; n11517
g11262 and n11264_not n11517_not ; n11518
g11263 and b[20] n11253_not ; n11519
g11264 and n11251_not n11519 ; n11520
g11265 and n11255_not n11520_not ; n11521
g11266 and n11518_not n11521 ; n11522
g11267 and n11255_not n11522_not ; n11523
g11268 and b[21] n11244_not ; n11524
g11269 and n11242_not n11524 ; n11525
g11270 and n11246_not n11525_not ; n11526
g11271 and n11523_not n11526 ; n11527
g11272 and n11246_not n11527_not ; n11528
g11273 and b[22] n11235_not ; n11529
g11274 and n11233_not n11529 ; n11530
g11275 and n11237_not n11530_not ; n11531
g11276 and n11528_not n11531 ; n11532
g11277 and n11237_not n11532_not ; n11533
g11278 and b[23] n11226_not ; n11534
g11279 and n11224_not n11534 ; n11535
g11280 and n11228_not n11535_not ; n11536
g11281 and n11533_not n11536 ; n11537
g11282 and n11228_not n11537_not ; n11538
g11283 and b[24] n11217_not ; n11539
g11284 and n11215_not n11539 ; n11540
g11285 and n11219_not n11540_not ; n11541
g11286 and n11538_not n11541 ; n11542
g11287 and n11219_not n11542_not ; n11543
g11288 and b[25] n11208_not ; n11544
g11289 and n11206_not n11544 ; n11545
g11290 and n11210_not n11545_not ; n11546
g11291 and n11543_not n11546 ; n11547
g11292 and n11210_not n11547_not ; n11548
g11293 and b[26] n11199_not ; n11549
g11294 and n11197_not n11549 ; n11550
g11295 and n11201_not n11550_not ; n11551
g11296 and n11548_not n11551 ; n11552
g11297 and n11201_not n11552_not ; n11553
g11298 and b[27] n11190_not ; n11554
g11299 and n11188_not n11554 ; n11555
g11300 and n11192_not n11555_not ; n11556
g11301 and n11553_not n11556 ; n11557
g11302 and n11192_not n11557_not ; n11558
g11303 and b[28] n11181_not ; n11559
g11304 and n11179_not n11559 ; n11560
g11305 and n11183_not n11560_not ; n11561
g11306 and n11558_not n11561 ; n11562
g11307 and n11183_not n11562_not ; n11563
g11308 and b[29] n11172_not ; n11564
g11309 and n11170_not n11564 ; n11565
g11310 and n11174_not n11565_not ; n11566
g11311 and n11563_not n11566 ; n11567
g11312 and n11174_not n11567_not ; n11568
g11313 and b[30] n11163_not ; n11569
g11314 and n11161_not n11569 ; n11570
g11315 and n11165_not n11570_not ; n11571
g11316 and n11568_not n11571 ; n11572
g11317 and n11165_not n11572_not ; n11573
g11318 and b[31] n11154_not ; n11574
g11319 and n11152_not n11574 ; n11575
g11320 and n11156_not n11575_not ; n11576
g11321 and n11573_not n11576 ; n11577
g11322 and n11156_not n11577_not ; n11578
g11323 and b[32] n11145_not ; n11579
g11324 and n11143_not n11579 ; n11580
g11325 and n11147_not n11580_not ; n11581
g11326 and n11578_not n11581 ; n11582
g11327 and n11147_not n11582_not ; n11583
g11328 and b[33] n11136_not ; n11584
g11329 and n11134_not n11584 ; n11585
g11330 and n11138_not n11585_not ; n11586
g11331 and n11583_not n11586 ; n11587
g11332 and n11138_not n11587_not ; n11588
g11333 and b[34] n11127_not ; n11589
g11334 and n11125_not n11589 ; n11590
g11335 and n11129_not n11590_not ; n11591
g11336 and n11588_not n11591 ; n11592
g11337 and n11129_not n11592_not ; n11593
g11338 and b[35] n11118_not ; n11594
g11339 and n11116_not n11594 ; n11595
g11340 and n11120_not n11595_not ; n11596
g11341 and n11593_not n11596 ; n11597
g11342 and n11120_not n11597_not ; n11598
g11343 and b[36] n11109_not ; n11599
g11344 and n11107_not n11599 ; n11600
g11345 and n11111_not n11600_not ; n11601
g11346 and n11598_not n11601 ; n11602
g11347 and n11111_not n11602_not ; n11603
g11348 and b[37] n11100_not ; n11604
g11349 and n11098_not n11604 ; n11605
g11350 and n11102_not n11605_not ; n11606
g11351 and n11603_not n11606 ; n11607
g11352 and n11102_not n11607_not ; n11608
g11353 and b[38] n11080_not ; n11609
g11354 and n11078_not n11609 ; n11610
g11355 and n11093_not n11610_not ; n11611
g11356 and n11608_not n11611 ; n11612
g11357 and n11093_not n11612_not ; n11613
g11358 and b[39] n11090_not ; n11614
g11359 and n11088_not n11614 ; n11615
g11360 and n11092_not n11615_not ; n11616
g11361 and n11613_not n11616 ; n11617
g11362 and n11092_not n11617_not ; n11618
g11363 and n338 n340 ; n11619
g11364 and n11618_not n11619 ; quotient[24]
g11365 and n11081_not quotient[24]_not ; n11621
g11366 and n11102_not n11611 ; n11622
g11367 and n11607_not n11622 ; n11623
g11368 and n11608_not n11611_not ; n11624
g11369 and n11623_not n11624_not ; n11625
g11370 and n11619 n11625_not ; n11626
g11371 and n11618_not n11626 ; n11627
g11372 and n11621_not n11627_not ; n11628
g11373 and n11091_not quotient[24]_not ; n11629
g11374 and n11093_not n11616 ; n11630
g11375 and n11612_not n11630 ; n11631
g11376 and n11613_not n11616_not ; n11632
g11377 and n11631_not n11632_not ; n11633
g11378 and quotient[24] n11633_not ; n11634
g11379 and n11629_not n11634_not ; n11635
g11380 and b[40]_not n11635_not ; n11636
g11381 and b[39]_not n11628_not ; n11637
g11382 and n11101_not quotient[24]_not ; n11638
g11383 and n11111_not n11606 ; n11639
g11384 and n11602_not n11639 ; n11640
g11385 and n11603_not n11606_not ; n11641
g11386 and n11640_not n11641_not ; n11642
g11387 and n11619 n11642_not ; n11643
g11388 and n11618_not n11643 ; n11644
g11389 and n11638_not n11644_not ; n11645
g11390 and b[38]_not n11645_not ; n11646
g11391 and n11110_not quotient[24]_not ; n11647
g11392 and n11120_not n11601 ; n11648
g11393 and n11597_not n11648 ; n11649
g11394 and n11598_not n11601_not ; n11650
g11395 and n11649_not n11650_not ; n11651
g11396 and n11619 n11651_not ; n11652
g11397 and n11618_not n11652 ; n11653
g11398 and n11647_not n11653_not ; n11654
g11399 and b[37]_not n11654_not ; n11655
g11400 and n11119_not quotient[24]_not ; n11656
g11401 and n11129_not n11596 ; n11657
g11402 and n11592_not n11657 ; n11658
g11403 and n11593_not n11596_not ; n11659
g11404 and n11658_not n11659_not ; n11660
g11405 and n11619 n11660_not ; n11661
g11406 and n11618_not n11661 ; n11662
g11407 and n11656_not n11662_not ; n11663
g11408 and b[36]_not n11663_not ; n11664
g11409 and n11128_not quotient[24]_not ; n11665
g11410 and n11138_not n11591 ; n11666
g11411 and n11587_not n11666 ; n11667
g11412 and n11588_not n11591_not ; n11668
g11413 and n11667_not n11668_not ; n11669
g11414 and n11619 n11669_not ; n11670
g11415 and n11618_not n11670 ; n11671
g11416 and n11665_not n11671_not ; n11672
g11417 and b[35]_not n11672_not ; n11673
g11418 and n11137_not quotient[24]_not ; n11674
g11419 and n11147_not n11586 ; n11675
g11420 and n11582_not n11675 ; n11676
g11421 and n11583_not n11586_not ; n11677
g11422 and n11676_not n11677_not ; n11678
g11423 and n11619 n11678_not ; n11679
g11424 and n11618_not n11679 ; n11680
g11425 and n11674_not n11680_not ; n11681
g11426 and b[34]_not n11681_not ; n11682
g11427 and n11146_not quotient[24]_not ; n11683
g11428 and n11156_not n11581 ; n11684
g11429 and n11577_not n11684 ; n11685
g11430 and n11578_not n11581_not ; n11686
g11431 and n11685_not n11686_not ; n11687
g11432 and n11619 n11687_not ; n11688
g11433 and n11618_not n11688 ; n11689
g11434 and n11683_not n11689_not ; n11690
g11435 and b[33]_not n11690_not ; n11691
g11436 and n11155_not quotient[24]_not ; n11692
g11437 and n11165_not n11576 ; n11693
g11438 and n11572_not n11693 ; n11694
g11439 and n11573_not n11576_not ; n11695
g11440 and n11694_not n11695_not ; n11696
g11441 and n11619 n11696_not ; n11697
g11442 and n11618_not n11697 ; n11698
g11443 and n11692_not n11698_not ; n11699
g11444 and b[32]_not n11699_not ; n11700
g11445 and n11164_not quotient[24]_not ; n11701
g11446 and n11174_not n11571 ; n11702
g11447 and n11567_not n11702 ; n11703
g11448 and n11568_not n11571_not ; n11704
g11449 and n11703_not n11704_not ; n11705
g11450 and n11619 n11705_not ; n11706
g11451 and n11618_not n11706 ; n11707
g11452 and n11701_not n11707_not ; n11708
g11453 and b[31]_not n11708_not ; n11709
g11454 and n11173_not quotient[24]_not ; n11710
g11455 and n11183_not n11566 ; n11711
g11456 and n11562_not n11711 ; n11712
g11457 and n11563_not n11566_not ; n11713
g11458 and n11712_not n11713_not ; n11714
g11459 and n11619 n11714_not ; n11715
g11460 and n11618_not n11715 ; n11716
g11461 and n11710_not n11716_not ; n11717
g11462 and b[30]_not n11717_not ; n11718
g11463 and n11182_not quotient[24]_not ; n11719
g11464 and n11192_not n11561 ; n11720
g11465 and n11557_not n11720 ; n11721
g11466 and n11558_not n11561_not ; n11722
g11467 and n11721_not n11722_not ; n11723
g11468 and n11619 n11723_not ; n11724
g11469 and n11618_not n11724 ; n11725
g11470 and n11719_not n11725_not ; n11726
g11471 and b[29]_not n11726_not ; n11727
g11472 and n11191_not quotient[24]_not ; n11728
g11473 and n11201_not n11556 ; n11729
g11474 and n11552_not n11729 ; n11730
g11475 and n11553_not n11556_not ; n11731
g11476 and n11730_not n11731_not ; n11732
g11477 and n11619 n11732_not ; n11733
g11478 and n11618_not n11733 ; n11734
g11479 and n11728_not n11734_not ; n11735
g11480 and b[28]_not n11735_not ; n11736
g11481 and n11200_not quotient[24]_not ; n11737
g11482 and n11210_not n11551 ; n11738
g11483 and n11547_not n11738 ; n11739
g11484 and n11548_not n11551_not ; n11740
g11485 and n11739_not n11740_not ; n11741
g11486 and n11619 n11741_not ; n11742
g11487 and n11618_not n11742 ; n11743
g11488 and n11737_not n11743_not ; n11744
g11489 and b[27]_not n11744_not ; n11745
g11490 and n11209_not quotient[24]_not ; n11746
g11491 and n11219_not n11546 ; n11747
g11492 and n11542_not n11747 ; n11748
g11493 and n11543_not n11546_not ; n11749
g11494 and n11748_not n11749_not ; n11750
g11495 and n11619 n11750_not ; n11751
g11496 and n11618_not n11751 ; n11752
g11497 and n11746_not n11752_not ; n11753
g11498 and b[26]_not n11753_not ; n11754
g11499 and n11218_not quotient[24]_not ; n11755
g11500 and n11228_not n11541 ; n11756
g11501 and n11537_not n11756 ; n11757
g11502 and n11538_not n11541_not ; n11758
g11503 and n11757_not n11758_not ; n11759
g11504 and n11619 n11759_not ; n11760
g11505 and n11618_not n11760 ; n11761
g11506 and n11755_not n11761_not ; n11762
g11507 and b[25]_not n11762_not ; n11763
g11508 and n11227_not quotient[24]_not ; n11764
g11509 and n11237_not n11536 ; n11765
g11510 and n11532_not n11765 ; n11766
g11511 and n11533_not n11536_not ; n11767
g11512 and n11766_not n11767_not ; n11768
g11513 and n11619 n11768_not ; n11769
g11514 and n11618_not n11769 ; n11770
g11515 and n11764_not n11770_not ; n11771
g11516 and b[24]_not n11771_not ; n11772
g11517 and n11236_not quotient[24]_not ; n11773
g11518 and n11246_not n11531 ; n11774
g11519 and n11527_not n11774 ; n11775
g11520 and n11528_not n11531_not ; n11776
g11521 and n11775_not n11776_not ; n11777
g11522 and n11619 n11777_not ; n11778
g11523 and n11618_not n11778 ; n11779
g11524 and n11773_not n11779_not ; n11780
g11525 and b[23]_not n11780_not ; n11781
g11526 and n11245_not quotient[24]_not ; n11782
g11527 and n11255_not n11526 ; n11783
g11528 and n11522_not n11783 ; n11784
g11529 and n11523_not n11526_not ; n11785
g11530 and n11784_not n11785_not ; n11786
g11531 and n11619 n11786_not ; n11787
g11532 and n11618_not n11787 ; n11788
g11533 and n11782_not n11788_not ; n11789
g11534 and b[22]_not n11789_not ; n11790
g11535 and n11254_not quotient[24]_not ; n11791
g11536 and n11264_not n11521 ; n11792
g11537 and n11517_not n11792 ; n11793
g11538 and n11518_not n11521_not ; n11794
g11539 and n11793_not n11794_not ; n11795
g11540 and n11619 n11795_not ; n11796
g11541 and n11618_not n11796 ; n11797
g11542 and n11791_not n11797_not ; n11798
g11543 and b[21]_not n11798_not ; n11799
g11544 and n11263_not quotient[24]_not ; n11800
g11545 and n11273_not n11516 ; n11801
g11546 and n11512_not n11801 ; n11802
g11547 and n11513_not n11516_not ; n11803
g11548 and n11802_not n11803_not ; n11804
g11549 and n11619 n11804_not ; n11805
g11550 and n11618_not n11805 ; n11806
g11551 and n11800_not n11806_not ; n11807
g11552 and b[20]_not n11807_not ; n11808
g11553 and n11272_not quotient[24]_not ; n11809
g11554 and n11282_not n11511 ; n11810
g11555 and n11507_not n11810 ; n11811
g11556 and n11508_not n11511_not ; n11812
g11557 and n11811_not n11812_not ; n11813
g11558 and n11619 n11813_not ; n11814
g11559 and n11618_not n11814 ; n11815
g11560 and n11809_not n11815_not ; n11816
g11561 and b[19]_not n11816_not ; n11817
g11562 and n11281_not quotient[24]_not ; n11818
g11563 and n11291_not n11506 ; n11819
g11564 and n11502_not n11819 ; n11820
g11565 and n11503_not n11506_not ; n11821
g11566 and n11820_not n11821_not ; n11822
g11567 and n11619 n11822_not ; n11823
g11568 and n11618_not n11823 ; n11824
g11569 and n11818_not n11824_not ; n11825
g11570 and b[18]_not n11825_not ; n11826
g11571 and n11290_not quotient[24]_not ; n11827
g11572 and n11300_not n11501 ; n11828
g11573 and n11497_not n11828 ; n11829
g11574 and n11498_not n11501_not ; n11830
g11575 and n11829_not n11830_not ; n11831
g11576 and n11619 n11831_not ; n11832
g11577 and n11618_not n11832 ; n11833
g11578 and n11827_not n11833_not ; n11834
g11579 and b[17]_not n11834_not ; n11835
g11580 and n11299_not quotient[24]_not ; n11836
g11581 and n11309_not n11496 ; n11837
g11582 and n11492_not n11837 ; n11838
g11583 and n11493_not n11496_not ; n11839
g11584 and n11838_not n11839_not ; n11840
g11585 and n11619 n11840_not ; n11841
g11586 and n11618_not n11841 ; n11842
g11587 and n11836_not n11842_not ; n11843
g11588 and b[16]_not n11843_not ; n11844
g11589 and n11308_not quotient[24]_not ; n11845
g11590 and n11318_not n11491 ; n11846
g11591 and n11487_not n11846 ; n11847
g11592 and n11488_not n11491_not ; n11848
g11593 and n11847_not n11848_not ; n11849
g11594 and n11619 n11849_not ; n11850
g11595 and n11618_not n11850 ; n11851
g11596 and n11845_not n11851_not ; n11852
g11597 and b[15]_not n11852_not ; n11853
g11598 and n11317_not quotient[24]_not ; n11854
g11599 and n11327_not n11486 ; n11855
g11600 and n11482_not n11855 ; n11856
g11601 and n11483_not n11486_not ; n11857
g11602 and n11856_not n11857_not ; n11858
g11603 and n11619 n11858_not ; n11859
g11604 and n11618_not n11859 ; n11860
g11605 and n11854_not n11860_not ; n11861
g11606 and b[14]_not n11861_not ; n11862
g11607 and n11326_not quotient[24]_not ; n11863
g11608 and n11336_not n11481 ; n11864
g11609 and n11477_not n11864 ; n11865
g11610 and n11478_not n11481_not ; n11866
g11611 and n11865_not n11866_not ; n11867
g11612 and n11619 n11867_not ; n11868
g11613 and n11618_not n11868 ; n11869
g11614 and n11863_not n11869_not ; n11870
g11615 and b[13]_not n11870_not ; n11871
g11616 and n11335_not quotient[24]_not ; n11872
g11617 and n11345_not n11476 ; n11873
g11618 and n11472_not n11873 ; n11874
g11619 and n11473_not n11476_not ; n11875
g11620 and n11874_not n11875_not ; n11876
g11621 and n11619 n11876_not ; n11877
g11622 and n11618_not n11877 ; n11878
g11623 and n11872_not n11878_not ; n11879
g11624 and b[12]_not n11879_not ; n11880
g11625 and n11344_not quotient[24]_not ; n11881
g11626 and n11354_not n11471 ; n11882
g11627 and n11467_not n11882 ; n11883
g11628 and n11468_not n11471_not ; n11884
g11629 and n11883_not n11884_not ; n11885
g11630 and n11619 n11885_not ; n11886
g11631 and n11618_not n11886 ; n11887
g11632 and n11881_not n11887_not ; n11888
g11633 and b[11]_not n11888_not ; n11889
g11634 and n11353_not quotient[24]_not ; n11890
g11635 and n11363_not n11466 ; n11891
g11636 and n11462_not n11891 ; n11892
g11637 and n11463_not n11466_not ; n11893
g11638 and n11892_not n11893_not ; n11894
g11639 and n11619 n11894_not ; n11895
g11640 and n11618_not n11895 ; n11896
g11641 and n11890_not n11896_not ; n11897
g11642 and b[10]_not n11897_not ; n11898
g11643 and n11362_not quotient[24]_not ; n11899
g11644 and n11372_not n11461 ; n11900
g11645 and n11457_not n11900 ; n11901
g11646 and n11458_not n11461_not ; n11902
g11647 and n11901_not n11902_not ; n11903
g11648 and n11619 n11903_not ; n11904
g11649 and n11618_not n11904 ; n11905
g11650 and n11899_not n11905_not ; n11906
g11651 and b[9]_not n11906_not ; n11907
g11652 and n11371_not quotient[24]_not ; n11908
g11653 and n11381_not n11456 ; n11909
g11654 and n11452_not n11909 ; n11910
g11655 and n11453_not n11456_not ; n11911
g11656 and n11910_not n11911_not ; n11912
g11657 and n11619 n11912_not ; n11913
g11658 and n11618_not n11913 ; n11914
g11659 and n11908_not n11914_not ; n11915
g11660 and b[8]_not n11915_not ; n11916
g11661 and n11380_not quotient[24]_not ; n11917
g11662 and n11390_not n11451 ; n11918
g11663 and n11447_not n11918 ; n11919
g11664 and n11448_not n11451_not ; n11920
g11665 and n11919_not n11920_not ; n11921
g11666 and n11619 n11921_not ; n11922
g11667 and n11618_not n11922 ; n11923
g11668 and n11917_not n11923_not ; n11924
g11669 and b[7]_not n11924_not ; n11925
g11670 and n11389_not quotient[24]_not ; n11926
g11671 and n11399_not n11446 ; n11927
g11672 and n11442_not n11927 ; n11928
g11673 and n11443_not n11446_not ; n11929
g11674 and n11928_not n11929_not ; n11930
g11675 and n11619 n11930_not ; n11931
g11676 and n11618_not n11931 ; n11932
g11677 and n11926_not n11932_not ; n11933
g11678 and b[6]_not n11933_not ; n11934
g11679 and n11398_not quotient[24]_not ; n11935
g11680 and n11408_not n11441 ; n11936
g11681 and n11437_not n11936 ; n11937
g11682 and n11438_not n11441_not ; n11938
g11683 and n11937_not n11938_not ; n11939
g11684 and n11619 n11939_not ; n11940
g11685 and n11618_not n11940 ; n11941
g11686 and n11935_not n11941_not ; n11942
g11687 and b[5]_not n11942_not ; n11943
g11688 and n11407_not quotient[24]_not ; n11944
g11689 and n11416_not n11436 ; n11945
g11690 and n11432_not n11945 ; n11946
g11691 and n11433_not n11436_not ; n11947
g11692 and n11946_not n11947_not ; n11948
g11693 and n11619 n11948_not ; n11949
g11694 and n11618_not n11949 ; n11950
g11695 and n11944_not n11950_not ; n11951
g11696 and b[4]_not n11951_not ; n11952
g11697 and n11415_not quotient[24]_not ; n11953
g11698 and n11427_not n11431 ; n11954
g11699 and n11426_not n11954 ; n11955
g11700 and n11428_not n11431_not ; n11956
g11701 and n11955_not n11956_not ; n11957
g11702 and n11619 n11957_not ; n11958
g11703 and n11618_not n11958 ; n11959
g11704 and n11953_not n11959_not ; n11960
g11705 and b[3]_not n11960_not ; n11961
g11706 and n11420_not quotient[24]_not ; n11962
g11707 and n11423_not n11425 ; n11963
g11708 and n11421_not n11963 ; n11964
g11709 and n11619 n11964_not ; n11965
g11710 and n11426_not n11965 ; n11966
g11711 and n11618_not n11966 ; n11967
g11712 and n11962_not n11967_not ; n11968
g11713 and b[2]_not n11968_not ; n11969
g11714 and b[0] b[40]_not ; n11970
g11715 and n421 n11970 ; n11971
g11716 and n597 n11971 ; n11972
g11717 and n595 n11972 ; n11973
g11718 and n11618_not n11973 ; n11974
g11719 and a[24] n11974_not ; n11975
g11720 and n291 n11425 ; n11976
g11721 and n302 n11976 ; n11977
g11722 and n288 n11977 ; n11978
g11723 and n11618_not n11978 ; n11979
g11724 and n11975_not n11979_not ; n11980
g11725 and b[1] n11980_not ; n11981
g11726 and b[1]_not n11979_not ; n11982
g11727 and n11975_not n11982 ; n11983
g11728 and n11981_not n11983_not ; n11984
g11729 and a[23]_not b[0] ; n11985
g11730 and n11984_not n11985_not ; n11986
g11731 and b[1]_not n11980_not ; n11987
g11732 and n11986_not n11987_not ; n11988
g11733 and b[2] n11967_not ; n11989
g11734 and n11962_not n11989 ; n11990
g11735 and n11969_not n11990_not ; n11991
g11736 and n11988_not n11991 ; n11992
g11737 and n11969_not n11992_not ; n11993
g11738 and b[3] n11959_not ; n11994
g11739 and n11953_not n11994 ; n11995
g11740 and n11961_not n11995_not ; n11996
g11741 and n11993_not n11996 ; n11997
g11742 and n11961_not n11997_not ; n11998
g11743 and b[4] n11950_not ; n11999
g11744 and n11944_not n11999 ; n12000
g11745 and n11952_not n12000_not ; n12001
g11746 and n11998_not n12001 ; n12002
g11747 and n11952_not n12002_not ; n12003
g11748 and b[5] n11941_not ; n12004
g11749 and n11935_not n12004 ; n12005
g11750 and n11943_not n12005_not ; n12006
g11751 and n12003_not n12006 ; n12007
g11752 and n11943_not n12007_not ; n12008
g11753 and b[6] n11932_not ; n12009
g11754 and n11926_not n12009 ; n12010
g11755 and n11934_not n12010_not ; n12011
g11756 and n12008_not n12011 ; n12012
g11757 and n11934_not n12012_not ; n12013
g11758 and b[7] n11923_not ; n12014
g11759 and n11917_not n12014 ; n12015
g11760 and n11925_not n12015_not ; n12016
g11761 and n12013_not n12016 ; n12017
g11762 and n11925_not n12017_not ; n12018
g11763 and b[8] n11914_not ; n12019
g11764 and n11908_not n12019 ; n12020
g11765 and n11916_not n12020_not ; n12021
g11766 and n12018_not n12021 ; n12022
g11767 and n11916_not n12022_not ; n12023
g11768 and b[9] n11905_not ; n12024
g11769 and n11899_not n12024 ; n12025
g11770 and n11907_not n12025_not ; n12026
g11771 and n12023_not n12026 ; n12027
g11772 and n11907_not n12027_not ; n12028
g11773 and b[10] n11896_not ; n12029
g11774 and n11890_not n12029 ; n12030
g11775 and n11898_not n12030_not ; n12031
g11776 and n12028_not n12031 ; n12032
g11777 and n11898_not n12032_not ; n12033
g11778 and b[11] n11887_not ; n12034
g11779 and n11881_not n12034 ; n12035
g11780 and n11889_not n12035_not ; n12036
g11781 and n12033_not n12036 ; n12037
g11782 and n11889_not n12037_not ; n12038
g11783 and b[12] n11878_not ; n12039
g11784 and n11872_not n12039 ; n12040
g11785 and n11880_not n12040_not ; n12041
g11786 and n12038_not n12041 ; n12042
g11787 and n11880_not n12042_not ; n12043
g11788 and b[13] n11869_not ; n12044
g11789 and n11863_not n12044 ; n12045
g11790 and n11871_not n12045_not ; n12046
g11791 and n12043_not n12046 ; n12047
g11792 and n11871_not n12047_not ; n12048
g11793 and b[14] n11860_not ; n12049
g11794 and n11854_not n12049 ; n12050
g11795 and n11862_not n12050_not ; n12051
g11796 and n12048_not n12051 ; n12052
g11797 and n11862_not n12052_not ; n12053
g11798 and b[15] n11851_not ; n12054
g11799 and n11845_not n12054 ; n12055
g11800 and n11853_not n12055_not ; n12056
g11801 and n12053_not n12056 ; n12057
g11802 and n11853_not n12057_not ; n12058
g11803 and b[16] n11842_not ; n12059
g11804 and n11836_not n12059 ; n12060
g11805 and n11844_not n12060_not ; n12061
g11806 and n12058_not n12061 ; n12062
g11807 and n11844_not n12062_not ; n12063
g11808 and b[17] n11833_not ; n12064
g11809 and n11827_not n12064 ; n12065
g11810 and n11835_not n12065_not ; n12066
g11811 and n12063_not n12066 ; n12067
g11812 and n11835_not n12067_not ; n12068
g11813 and b[18] n11824_not ; n12069
g11814 and n11818_not n12069 ; n12070
g11815 and n11826_not n12070_not ; n12071
g11816 and n12068_not n12071 ; n12072
g11817 and n11826_not n12072_not ; n12073
g11818 and b[19] n11815_not ; n12074
g11819 and n11809_not n12074 ; n12075
g11820 and n11817_not n12075_not ; n12076
g11821 and n12073_not n12076 ; n12077
g11822 and n11817_not n12077_not ; n12078
g11823 and b[20] n11806_not ; n12079
g11824 and n11800_not n12079 ; n12080
g11825 and n11808_not n12080_not ; n12081
g11826 and n12078_not n12081 ; n12082
g11827 and n11808_not n12082_not ; n12083
g11828 and b[21] n11797_not ; n12084
g11829 and n11791_not n12084 ; n12085
g11830 and n11799_not n12085_not ; n12086
g11831 and n12083_not n12086 ; n12087
g11832 and n11799_not n12087_not ; n12088
g11833 and b[22] n11788_not ; n12089
g11834 and n11782_not n12089 ; n12090
g11835 and n11790_not n12090_not ; n12091
g11836 and n12088_not n12091 ; n12092
g11837 and n11790_not n12092_not ; n12093
g11838 and b[23] n11779_not ; n12094
g11839 and n11773_not n12094 ; n12095
g11840 and n11781_not n12095_not ; n12096
g11841 and n12093_not n12096 ; n12097
g11842 and n11781_not n12097_not ; n12098
g11843 and b[24] n11770_not ; n12099
g11844 and n11764_not n12099 ; n12100
g11845 and n11772_not n12100_not ; n12101
g11846 and n12098_not n12101 ; n12102
g11847 and n11772_not n12102_not ; n12103
g11848 and b[25] n11761_not ; n12104
g11849 and n11755_not n12104 ; n12105
g11850 and n11763_not n12105_not ; n12106
g11851 and n12103_not n12106 ; n12107
g11852 and n11763_not n12107_not ; n12108
g11853 and b[26] n11752_not ; n12109
g11854 and n11746_not n12109 ; n12110
g11855 and n11754_not n12110_not ; n12111
g11856 and n12108_not n12111 ; n12112
g11857 and n11754_not n12112_not ; n12113
g11858 and b[27] n11743_not ; n12114
g11859 and n11737_not n12114 ; n12115
g11860 and n11745_not n12115_not ; n12116
g11861 and n12113_not n12116 ; n12117
g11862 and n11745_not n12117_not ; n12118
g11863 and b[28] n11734_not ; n12119
g11864 and n11728_not n12119 ; n12120
g11865 and n11736_not n12120_not ; n12121
g11866 and n12118_not n12121 ; n12122
g11867 and n11736_not n12122_not ; n12123
g11868 and b[29] n11725_not ; n12124
g11869 and n11719_not n12124 ; n12125
g11870 and n11727_not n12125_not ; n12126
g11871 and n12123_not n12126 ; n12127
g11872 and n11727_not n12127_not ; n12128
g11873 and b[30] n11716_not ; n12129
g11874 and n11710_not n12129 ; n12130
g11875 and n11718_not n12130_not ; n12131
g11876 and n12128_not n12131 ; n12132
g11877 and n11718_not n12132_not ; n12133
g11878 and b[31] n11707_not ; n12134
g11879 and n11701_not n12134 ; n12135
g11880 and n11709_not n12135_not ; n12136
g11881 and n12133_not n12136 ; n12137
g11882 and n11709_not n12137_not ; n12138
g11883 and b[32] n11698_not ; n12139
g11884 and n11692_not n12139 ; n12140
g11885 and n11700_not n12140_not ; n12141
g11886 and n12138_not n12141 ; n12142
g11887 and n11700_not n12142_not ; n12143
g11888 and b[33] n11689_not ; n12144
g11889 and n11683_not n12144 ; n12145
g11890 and n11691_not n12145_not ; n12146
g11891 and n12143_not n12146 ; n12147
g11892 and n11691_not n12147_not ; n12148
g11893 and b[34] n11680_not ; n12149
g11894 and n11674_not n12149 ; n12150
g11895 and n11682_not n12150_not ; n12151
g11896 and n12148_not n12151 ; n12152
g11897 and n11682_not n12152_not ; n12153
g11898 and b[35] n11671_not ; n12154
g11899 and n11665_not n12154 ; n12155
g11900 and n11673_not n12155_not ; n12156
g11901 and n12153_not n12156 ; n12157
g11902 and n11673_not n12157_not ; n12158
g11903 and b[36] n11662_not ; n12159
g11904 and n11656_not n12159 ; n12160
g11905 and n11664_not n12160_not ; n12161
g11906 and n12158_not n12161 ; n12162
g11907 and n11664_not n12162_not ; n12163
g11908 and b[37] n11653_not ; n12164
g11909 and n11647_not n12164 ; n12165
g11910 and n11655_not n12165_not ; n12166
g11911 and n12163_not n12166 ; n12167
g11912 and n11655_not n12167_not ; n12168
g11913 and b[38] n11644_not ; n12169
g11914 and n11638_not n12169 ; n12170
g11915 and n11646_not n12170_not ; n12171
g11916 and n12168_not n12171 ; n12172
g11917 and n11646_not n12172_not ; n12173
g11918 and b[39] n11627_not ; n12174
g11919 and n11621_not n12174 ; n12175
g11920 and n11637_not n12175_not ; n12176
g11921 and n12173_not n12176 ; n12177
g11922 and n11637_not n12177_not ; n12178
g11923 and b[40] n11629_not ; n12179
g11924 and n11634_not n12179 ; n12180
g11925 and n11636_not n12180_not ; n12181
g11926 and n12178_not n12181 ; n12182
g11927 and n11636_not n12182_not ; n12183
g11928 and n408 n422 ; n12184
g11929 and n12183_not n12184 ; quotient[23]
g11930 and n11628_not quotient[23]_not ; n12186
g11931 and n11646_not n12176 ; n12187
g11932 and n12172_not n12187 ; n12188
g11933 and n12173_not n12176_not ; n12189
g11934 and n12188_not n12189_not ; n12190
g11935 and n12184 n12190_not ; n12191
g11936 and n12183_not n12191 ; n12192
g11937 and n12186_not n12192_not ; n12193
g11938 and b[40]_not n12193_not ; n12194
g11939 and n11645_not quotient[23]_not ; n12195
g11940 and n11655_not n12171 ; n12196
g11941 and n12167_not n12196 ; n12197
g11942 and n12168_not n12171_not ; n12198
g11943 and n12197_not n12198_not ; n12199
g11944 and n12184 n12199_not ; n12200
g11945 and n12183_not n12200 ; n12201
g11946 and n12195_not n12201_not ; n12202
g11947 and b[39]_not n12202_not ; n12203
g11948 and n11654_not quotient[23]_not ; n12204
g11949 and n11664_not n12166 ; n12205
g11950 and n12162_not n12205 ; n12206
g11951 and n12163_not n12166_not ; n12207
g11952 and n12206_not n12207_not ; n12208
g11953 and n12184 n12208_not ; n12209
g11954 and n12183_not n12209 ; n12210
g11955 and n12204_not n12210_not ; n12211
g11956 and b[38]_not n12211_not ; n12212
g11957 and n11663_not quotient[23]_not ; n12213
g11958 and n11673_not n12161 ; n12214
g11959 and n12157_not n12214 ; n12215
g11960 and n12158_not n12161_not ; n12216
g11961 and n12215_not n12216_not ; n12217
g11962 and n12184 n12217_not ; n12218
g11963 and n12183_not n12218 ; n12219
g11964 and n12213_not n12219_not ; n12220
g11965 and b[37]_not n12220_not ; n12221
g11966 and n11672_not quotient[23]_not ; n12222
g11967 and n11682_not n12156 ; n12223
g11968 and n12152_not n12223 ; n12224
g11969 and n12153_not n12156_not ; n12225
g11970 and n12224_not n12225_not ; n12226
g11971 and n12184 n12226_not ; n12227
g11972 and n12183_not n12227 ; n12228
g11973 and n12222_not n12228_not ; n12229
g11974 and b[36]_not n12229_not ; n12230
g11975 and n11681_not quotient[23]_not ; n12231
g11976 and n11691_not n12151 ; n12232
g11977 and n12147_not n12232 ; n12233
g11978 and n12148_not n12151_not ; n12234
g11979 and n12233_not n12234_not ; n12235
g11980 and n12184 n12235_not ; n12236
g11981 and n12183_not n12236 ; n12237
g11982 and n12231_not n12237_not ; n12238
g11983 and b[35]_not n12238_not ; n12239
g11984 and n11690_not quotient[23]_not ; n12240
g11985 and n11700_not n12146 ; n12241
g11986 and n12142_not n12241 ; n12242
g11987 and n12143_not n12146_not ; n12243
g11988 and n12242_not n12243_not ; n12244
g11989 and n12184 n12244_not ; n12245
g11990 and n12183_not n12245 ; n12246
g11991 and n12240_not n12246_not ; n12247
g11992 and b[34]_not n12247_not ; n12248
g11993 and n11699_not quotient[23]_not ; n12249
g11994 and n11709_not n12141 ; n12250
g11995 and n12137_not n12250 ; n12251
g11996 and n12138_not n12141_not ; n12252
g11997 and n12251_not n12252_not ; n12253
g11998 and n12184 n12253_not ; n12254
g11999 and n12183_not n12254 ; n12255
g12000 and n12249_not n12255_not ; n12256
g12001 and b[33]_not n12256_not ; n12257
g12002 and n11708_not quotient[23]_not ; n12258
g12003 and n11718_not n12136 ; n12259
g12004 and n12132_not n12259 ; n12260
g12005 and n12133_not n12136_not ; n12261
g12006 and n12260_not n12261_not ; n12262
g12007 and n12184 n12262_not ; n12263
g12008 and n12183_not n12263 ; n12264
g12009 and n12258_not n12264_not ; n12265
g12010 and b[32]_not n12265_not ; n12266
g12011 and n11717_not quotient[23]_not ; n12267
g12012 and n11727_not n12131 ; n12268
g12013 and n12127_not n12268 ; n12269
g12014 and n12128_not n12131_not ; n12270
g12015 and n12269_not n12270_not ; n12271
g12016 and n12184 n12271_not ; n12272
g12017 and n12183_not n12272 ; n12273
g12018 and n12267_not n12273_not ; n12274
g12019 and b[31]_not n12274_not ; n12275
g12020 and n11726_not quotient[23]_not ; n12276
g12021 and n11736_not n12126 ; n12277
g12022 and n12122_not n12277 ; n12278
g12023 and n12123_not n12126_not ; n12279
g12024 and n12278_not n12279_not ; n12280
g12025 and n12184 n12280_not ; n12281
g12026 and n12183_not n12281 ; n12282
g12027 and n12276_not n12282_not ; n12283
g12028 and b[30]_not n12283_not ; n12284
g12029 and n11735_not quotient[23]_not ; n12285
g12030 and n11745_not n12121 ; n12286
g12031 and n12117_not n12286 ; n12287
g12032 and n12118_not n12121_not ; n12288
g12033 and n12287_not n12288_not ; n12289
g12034 and n12184 n12289_not ; n12290
g12035 and n12183_not n12290 ; n12291
g12036 and n12285_not n12291_not ; n12292
g12037 and b[29]_not n12292_not ; n12293
g12038 and n11744_not quotient[23]_not ; n12294
g12039 and n11754_not n12116 ; n12295
g12040 and n12112_not n12295 ; n12296
g12041 and n12113_not n12116_not ; n12297
g12042 and n12296_not n12297_not ; n12298
g12043 and n12184 n12298_not ; n12299
g12044 and n12183_not n12299 ; n12300
g12045 and n12294_not n12300_not ; n12301
g12046 and b[28]_not n12301_not ; n12302
g12047 and n11753_not quotient[23]_not ; n12303
g12048 and n11763_not n12111 ; n12304
g12049 and n12107_not n12304 ; n12305
g12050 and n12108_not n12111_not ; n12306
g12051 and n12305_not n12306_not ; n12307
g12052 and n12184 n12307_not ; n12308
g12053 and n12183_not n12308 ; n12309
g12054 and n12303_not n12309_not ; n12310
g12055 and b[27]_not n12310_not ; n12311
g12056 and n11762_not quotient[23]_not ; n12312
g12057 and n11772_not n12106 ; n12313
g12058 and n12102_not n12313 ; n12314
g12059 and n12103_not n12106_not ; n12315
g12060 and n12314_not n12315_not ; n12316
g12061 and n12184 n12316_not ; n12317
g12062 and n12183_not n12317 ; n12318
g12063 and n12312_not n12318_not ; n12319
g12064 and b[26]_not n12319_not ; n12320
g12065 and n11771_not quotient[23]_not ; n12321
g12066 and n11781_not n12101 ; n12322
g12067 and n12097_not n12322 ; n12323
g12068 and n12098_not n12101_not ; n12324
g12069 and n12323_not n12324_not ; n12325
g12070 and n12184 n12325_not ; n12326
g12071 and n12183_not n12326 ; n12327
g12072 and n12321_not n12327_not ; n12328
g12073 and b[25]_not n12328_not ; n12329
g12074 and n11780_not quotient[23]_not ; n12330
g12075 and n11790_not n12096 ; n12331
g12076 and n12092_not n12331 ; n12332
g12077 and n12093_not n12096_not ; n12333
g12078 and n12332_not n12333_not ; n12334
g12079 and n12184 n12334_not ; n12335
g12080 and n12183_not n12335 ; n12336
g12081 and n12330_not n12336_not ; n12337
g12082 and b[24]_not n12337_not ; n12338
g12083 and n11789_not quotient[23]_not ; n12339
g12084 and n11799_not n12091 ; n12340
g12085 and n12087_not n12340 ; n12341
g12086 and n12088_not n12091_not ; n12342
g12087 and n12341_not n12342_not ; n12343
g12088 and n12184 n12343_not ; n12344
g12089 and n12183_not n12344 ; n12345
g12090 and n12339_not n12345_not ; n12346
g12091 and b[23]_not n12346_not ; n12347
g12092 and n11798_not quotient[23]_not ; n12348
g12093 and n11808_not n12086 ; n12349
g12094 and n12082_not n12349 ; n12350
g12095 and n12083_not n12086_not ; n12351
g12096 and n12350_not n12351_not ; n12352
g12097 and n12184 n12352_not ; n12353
g12098 and n12183_not n12353 ; n12354
g12099 and n12348_not n12354_not ; n12355
g12100 and b[22]_not n12355_not ; n12356
g12101 and n11807_not quotient[23]_not ; n12357
g12102 and n11817_not n12081 ; n12358
g12103 and n12077_not n12358 ; n12359
g12104 and n12078_not n12081_not ; n12360
g12105 and n12359_not n12360_not ; n12361
g12106 and n12184 n12361_not ; n12362
g12107 and n12183_not n12362 ; n12363
g12108 and n12357_not n12363_not ; n12364
g12109 and b[21]_not n12364_not ; n12365
g12110 and n11816_not quotient[23]_not ; n12366
g12111 and n11826_not n12076 ; n12367
g12112 and n12072_not n12367 ; n12368
g12113 and n12073_not n12076_not ; n12369
g12114 and n12368_not n12369_not ; n12370
g12115 and n12184 n12370_not ; n12371
g12116 and n12183_not n12371 ; n12372
g12117 and n12366_not n12372_not ; n12373
g12118 and b[20]_not n12373_not ; n12374
g12119 and n11825_not quotient[23]_not ; n12375
g12120 and n11835_not n12071 ; n12376
g12121 and n12067_not n12376 ; n12377
g12122 and n12068_not n12071_not ; n12378
g12123 and n12377_not n12378_not ; n12379
g12124 and n12184 n12379_not ; n12380
g12125 and n12183_not n12380 ; n12381
g12126 and n12375_not n12381_not ; n12382
g12127 and b[19]_not n12382_not ; n12383
g12128 and n11834_not quotient[23]_not ; n12384
g12129 and n11844_not n12066 ; n12385
g12130 and n12062_not n12385 ; n12386
g12131 and n12063_not n12066_not ; n12387
g12132 and n12386_not n12387_not ; n12388
g12133 and n12184 n12388_not ; n12389
g12134 and n12183_not n12389 ; n12390
g12135 and n12384_not n12390_not ; n12391
g12136 and b[18]_not n12391_not ; n12392
g12137 and n11843_not quotient[23]_not ; n12393
g12138 and n11853_not n12061 ; n12394
g12139 and n12057_not n12394 ; n12395
g12140 and n12058_not n12061_not ; n12396
g12141 and n12395_not n12396_not ; n12397
g12142 and n12184 n12397_not ; n12398
g12143 and n12183_not n12398 ; n12399
g12144 and n12393_not n12399_not ; n12400
g12145 and b[17]_not n12400_not ; n12401
g12146 and n11852_not quotient[23]_not ; n12402
g12147 and n11862_not n12056 ; n12403
g12148 and n12052_not n12403 ; n12404
g12149 and n12053_not n12056_not ; n12405
g12150 and n12404_not n12405_not ; n12406
g12151 and n12184 n12406_not ; n12407
g12152 and n12183_not n12407 ; n12408
g12153 and n12402_not n12408_not ; n12409
g12154 and b[16]_not n12409_not ; n12410
g12155 and n11861_not quotient[23]_not ; n12411
g12156 and n11871_not n12051 ; n12412
g12157 and n12047_not n12412 ; n12413
g12158 and n12048_not n12051_not ; n12414
g12159 and n12413_not n12414_not ; n12415
g12160 and n12184 n12415_not ; n12416
g12161 and n12183_not n12416 ; n12417
g12162 and n12411_not n12417_not ; n12418
g12163 and b[15]_not n12418_not ; n12419
g12164 and n11870_not quotient[23]_not ; n12420
g12165 and n11880_not n12046 ; n12421
g12166 and n12042_not n12421 ; n12422
g12167 and n12043_not n12046_not ; n12423
g12168 and n12422_not n12423_not ; n12424
g12169 and n12184 n12424_not ; n12425
g12170 and n12183_not n12425 ; n12426
g12171 and n12420_not n12426_not ; n12427
g12172 and b[14]_not n12427_not ; n12428
g12173 and n11879_not quotient[23]_not ; n12429
g12174 and n11889_not n12041 ; n12430
g12175 and n12037_not n12430 ; n12431
g12176 and n12038_not n12041_not ; n12432
g12177 and n12431_not n12432_not ; n12433
g12178 and n12184 n12433_not ; n12434
g12179 and n12183_not n12434 ; n12435
g12180 and n12429_not n12435_not ; n12436
g12181 and b[13]_not n12436_not ; n12437
g12182 and n11888_not quotient[23]_not ; n12438
g12183 and n11898_not n12036 ; n12439
g12184 and n12032_not n12439 ; n12440
g12185 and n12033_not n12036_not ; n12441
g12186 and n12440_not n12441_not ; n12442
g12187 and n12184 n12442_not ; n12443
g12188 and n12183_not n12443 ; n12444
g12189 and n12438_not n12444_not ; n12445
g12190 and b[12]_not n12445_not ; n12446
g12191 and n11897_not quotient[23]_not ; n12447
g12192 and n11907_not n12031 ; n12448
g12193 and n12027_not n12448 ; n12449
g12194 and n12028_not n12031_not ; n12450
g12195 and n12449_not n12450_not ; n12451
g12196 and n12184 n12451_not ; n12452
g12197 and n12183_not n12452 ; n12453
g12198 and n12447_not n12453_not ; n12454
g12199 and b[11]_not n12454_not ; n12455
g12200 and n11906_not quotient[23]_not ; n12456
g12201 and n11916_not n12026 ; n12457
g12202 and n12022_not n12457 ; n12458
g12203 and n12023_not n12026_not ; n12459
g12204 and n12458_not n12459_not ; n12460
g12205 and n12184 n12460_not ; n12461
g12206 and n12183_not n12461 ; n12462
g12207 and n12456_not n12462_not ; n12463
g12208 and b[10]_not n12463_not ; n12464
g12209 and n11915_not quotient[23]_not ; n12465
g12210 and n11925_not n12021 ; n12466
g12211 and n12017_not n12466 ; n12467
g12212 and n12018_not n12021_not ; n12468
g12213 and n12467_not n12468_not ; n12469
g12214 and n12184 n12469_not ; n12470
g12215 and n12183_not n12470 ; n12471
g12216 and n12465_not n12471_not ; n12472
g12217 and b[9]_not n12472_not ; n12473
g12218 and n11924_not quotient[23]_not ; n12474
g12219 and n11934_not n12016 ; n12475
g12220 and n12012_not n12475 ; n12476
g12221 and n12013_not n12016_not ; n12477
g12222 and n12476_not n12477_not ; n12478
g12223 and n12184 n12478_not ; n12479
g12224 and n12183_not n12479 ; n12480
g12225 and n12474_not n12480_not ; n12481
g12226 and b[8]_not n12481_not ; n12482
g12227 and n11933_not quotient[23]_not ; n12483
g12228 and n11943_not n12011 ; n12484
g12229 and n12007_not n12484 ; n12485
g12230 and n12008_not n12011_not ; n12486
g12231 and n12485_not n12486_not ; n12487
g12232 and n12184 n12487_not ; n12488
g12233 and n12183_not n12488 ; n12489
g12234 and n12483_not n12489_not ; n12490
g12235 and b[7]_not n12490_not ; n12491
g12236 and n11942_not quotient[23]_not ; n12492
g12237 and n11952_not n12006 ; n12493
g12238 and n12002_not n12493 ; n12494
g12239 and n12003_not n12006_not ; n12495
g12240 and n12494_not n12495_not ; n12496
g12241 and n12184 n12496_not ; n12497
g12242 and n12183_not n12497 ; n12498
g12243 and n12492_not n12498_not ; n12499
g12244 and b[6]_not n12499_not ; n12500
g12245 and n11951_not quotient[23]_not ; n12501
g12246 and n11961_not n12001 ; n12502
g12247 and n11997_not n12502 ; n12503
g12248 and n11998_not n12001_not ; n12504
g12249 and n12503_not n12504_not ; n12505
g12250 and n12184 n12505_not ; n12506
g12251 and n12183_not n12506 ; n12507
g12252 and n12501_not n12507_not ; n12508
g12253 and b[5]_not n12508_not ; n12509
g12254 and n11960_not quotient[23]_not ; n12510
g12255 and n11969_not n11996 ; n12511
g12256 and n11992_not n12511 ; n12512
g12257 and n11993_not n11996_not ; n12513
g12258 and n12512_not n12513_not ; n12514
g12259 and n12184 n12514_not ; n12515
g12260 and n12183_not n12515 ; n12516
g12261 and n12510_not n12516_not ; n12517
g12262 and b[4]_not n12517_not ; n12518
g12263 and n11968_not quotient[23]_not ; n12519
g12264 and n11987_not n11991 ; n12520
g12265 and n11986_not n12520 ; n12521
g12266 and n11988_not n11991_not ; n12522
g12267 and n12521_not n12522_not ; n12523
g12268 and n12184 n12523_not ; n12524
g12269 and n12183_not n12524 ; n12525
g12270 and n12519_not n12525_not ; n12526
g12271 and b[3]_not n12526_not ; n12527
g12272 and n11980_not quotient[23]_not ; n12528
g12273 and n11983_not n11985 ; n12529
g12274 and n11981_not n12529 ; n12530
g12275 and n12184 n12530_not ; n12531
g12276 and n11986_not n12531 ; n12532
g12277 and n12183_not n12532 ; n12533
g12278 and n12528_not n12533_not ; n12534
g12279 and b[2]_not n12534_not ; n12535
g12280 and b[0] b[41]_not ; n12536
g12281 and n290 n12536 ; n12537
g12282 and n301 n12537 ; n12538
g12283 and n338 n12538 ; n12539
g12284 and n12183_not n12539 ; n12540
g12285 and a[23] n12540_not ; n12541
g12286 and n421 n11985 ; n12542
g12287 and n597 n12542 ; n12543
g12288 and n595 n12543 ; n12544
g12289 and n12183_not n12544 ; n12545
g12290 and n12541_not n12545_not ; n12546
g12291 and b[1] n12546_not ; n12547
g12292 and b[1]_not n12545_not ; n12548
g12293 and n12541_not n12548 ; n12549
g12294 and n12547_not n12549_not ; n12550
g12295 and a[22]_not b[0] ; n12551
g12296 and n12550_not n12551_not ; n12552
g12297 and b[1]_not n12546_not ; n12553
g12298 and n12552_not n12553_not ; n12554
g12299 and b[2] n12533_not ; n12555
g12300 and n12528_not n12555 ; n12556
g12301 and n12535_not n12556_not ; n12557
g12302 and n12554_not n12557 ; n12558
g12303 and n12535_not n12558_not ; n12559
g12304 and b[3] n12525_not ; n12560
g12305 and n12519_not n12560 ; n12561
g12306 and n12527_not n12561_not ; n12562
g12307 and n12559_not n12562 ; n12563
g12308 and n12527_not n12563_not ; n12564
g12309 and b[4] n12516_not ; n12565
g12310 and n12510_not n12565 ; n12566
g12311 and n12518_not n12566_not ; n12567
g12312 and n12564_not n12567 ; n12568
g12313 and n12518_not n12568_not ; n12569
g12314 and b[5] n12507_not ; n12570
g12315 and n12501_not n12570 ; n12571
g12316 and n12509_not n12571_not ; n12572
g12317 and n12569_not n12572 ; n12573
g12318 and n12509_not n12573_not ; n12574
g12319 and b[6] n12498_not ; n12575
g12320 and n12492_not n12575 ; n12576
g12321 and n12500_not n12576_not ; n12577
g12322 and n12574_not n12577 ; n12578
g12323 and n12500_not n12578_not ; n12579
g12324 and b[7] n12489_not ; n12580
g12325 and n12483_not n12580 ; n12581
g12326 and n12491_not n12581_not ; n12582
g12327 and n12579_not n12582 ; n12583
g12328 and n12491_not n12583_not ; n12584
g12329 and b[8] n12480_not ; n12585
g12330 and n12474_not n12585 ; n12586
g12331 and n12482_not n12586_not ; n12587
g12332 and n12584_not n12587 ; n12588
g12333 and n12482_not n12588_not ; n12589
g12334 and b[9] n12471_not ; n12590
g12335 and n12465_not n12590 ; n12591
g12336 and n12473_not n12591_not ; n12592
g12337 and n12589_not n12592 ; n12593
g12338 and n12473_not n12593_not ; n12594
g12339 and b[10] n12462_not ; n12595
g12340 and n12456_not n12595 ; n12596
g12341 and n12464_not n12596_not ; n12597
g12342 and n12594_not n12597 ; n12598
g12343 and n12464_not n12598_not ; n12599
g12344 and b[11] n12453_not ; n12600
g12345 and n12447_not n12600 ; n12601
g12346 and n12455_not n12601_not ; n12602
g12347 and n12599_not n12602 ; n12603
g12348 and n12455_not n12603_not ; n12604
g12349 and b[12] n12444_not ; n12605
g12350 and n12438_not n12605 ; n12606
g12351 and n12446_not n12606_not ; n12607
g12352 and n12604_not n12607 ; n12608
g12353 and n12446_not n12608_not ; n12609
g12354 and b[13] n12435_not ; n12610
g12355 and n12429_not n12610 ; n12611
g12356 and n12437_not n12611_not ; n12612
g12357 and n12609_not n12612 ; n12613
g12358 and n12437_not n12613_not ; n12614
g12359 and b[14] n12426_not ; n12615
g12360 and n12420_not n12615 ; n12616
g12361 and n12428_not n12616_not ; n12617
g12362 and n12614_not n12617 ; n12618
g12363 and n12428_not n12618_not ; n12619
g12364 and b[15] n12417_not ; n12620
g12365 and n12411_not n12620 ; n12621
g12366 and n12419_not n12621_not ; n12622
g12367 and n12619_not n12622 ; n12623
g12368 and n12419_not n12623_not ; n12624
g12369 and b[16] n12408_not ; n12625
g12370 and n12402_not n12625 ; n12626
g12371 and n12410_not n12626_not ; n12627
g12372 and n12624_not n12627 ; n12628
g12373 and n12410_not n12628_not ; n12629
g12374 and b[17] n12399_not ; n12630
g12375 and n12393_not n12630 ; n12631
g12376 and n12401_not n12631_not ; n12632
g12377 and n12629_not n12632 ; n12633
g12378 and n12401_not n12633_not ; n12634
g12379 and b[18] n12390_not ; n12635
g12380 and n12384_not n12635 ; n12636
g12381 and n12392_not n12636_not ; n12637
g12382 and n12634_not n12637 ; n12638
g12383 and n12392_not n12638_not ; n12639
g12384 and b[19] n12381_not ; n12640
g12385 and n12375_not n12640 ; n12641
g12386 and n12383_not n12641_not ; n12642
g12387 and n12639_not n12642 ; n12643
g12388 and n12383_not n12643_not ; n12644
g12389 and b[20] n12372_not ; n12645
g12390 and n12366_not n12645 ; n12646
g12391 and n12374_not n12646_not ; n12647
g12392 and n12644_not n12647 ; n12648
g12393 and n12374_not n12648_not ; n12649
g12394 and b[21] n12363_not ; n12650
g12395 and n12357_not n12650 ; n12651
g12396 and n12365_not n12651_not ; n12652
g12397 and n12649_not n12652 ; n12653
g12398 and n12365_not n12653_not ; n12654
g12399 and b[22] n12354_not ; n12655
g12400 and n12348_not n12655 ; n12656
g12401 and n12356_not n12656_not ; n12657
g12402 and n12654_not n12657 ; n12658
g12403 and n12356_not n12658_not ; n12659
g12404 and b[23] n12345_not ; n12660
g12405 and n12339_not n12660 ; n12661
g12406 and n12347_not n12661_not ; n12662
g12407 and n12659_not n12662 ; n12663
g12408 and n12347_not n12663_not ; n12664
g12409 and b[24] n12336_not ; n12665
g12410 and n12330_not n12665 ; n12666
g12411 and n12338_not n12666_not ; n12667
g12412 and n12664_not n12667 ; n12668
g12413 and n12338_not n12668_not ; n12669
g12414 and b[25] n12327_not ; n12670
g12415 and n12321_not n12670 ; n12671
g12416 and n12329_not n12671_not ; n12672
g12417 and n12669_not n12672 ; n12673
g12418 and n12329_not n12673_not ; n12674
g12419 and b[26] n12318_not ; n12675
g12420 and n12312_not n12675 ; n12676
g12421 and n12320_not n12676_not ; n12677
g12422 and n12674_not n12677 ; n12678
g12423 and n12320_not n12678_not ; n12679
g12424 and b[27] n12309_not ; n12680
g12425 and n12303_not n12680 ; n12681
g12426 and n12311_not n12681_not ; n12682
g12427 and n12679_not n12682 ; n12683
g12428 and n12311_not n12683_not ; n12684
g12429 and b[28] n12300_not ; n12685
g12430 and n12294_not n12685 ; n12686
g12431 and n12302_not n12686_not ; n12687
g12432 and n12684_not n12687 ; n12688
g12433 and n12302_not n12688_not ; n12689
g12434 and b[29] n12291_not ; n12690
g12435 and n12285_not n12690 ; n12691
g12436 and n12293_not n12691_not ; n12692
g12437 and n12689_not n12692 ; n12693
g12438 and n12293_not n12693_not ; n12694
g12439 and b[30] n12282_not ; n12695
g12440 and n12276_not n12695 ; n12696
g12441 and n12284_not n12696_not ; n12697
g12442 and n12694_not n12697 ; n12698
g12443 and n12284_not n12698_not ; n12699
g12444 and b[31] n12273_not ; n12700
g12445 and n12267_not n12700 ; n12701
g12446 and n12275_not n12701_not ; n12702
g12447 and n12699_not n12702 ; n12703
g12448 and n12275_not n12703_not ; n12704
g12449 and b[32] n12264_not ; n12705
g12450 and n12258_not n12705 ; n12706
g12451 and n12266_not n12706_not ; n12707
g12452 and n12704_not n12707 ; n12708
g12453 and n12266_not n12708_not ; n12709
g12454 and b[33] n12255_not ; n12710
g12455 and n12249_not n12710 ; n12711
g12456 and n12257_not n12711_not ; n12712
g12457 and n12709_not n12712 ; n12713
g12458 and n12257_not n12713_not ; n12714
g12459 and b[34] n12246_not ; n12715
g12460 and n12240_not n12715 ; n12716
g12461 and n12248_not n12716_not ; n12717
g12462 and n12714_not n12717 ; n12718
g12463 and n12248_not n12718_not ; n12719
g12464 and b[35] n12237_not ; n12720
g12465 and n12231_not n12720 ; n12721
g12466 and n12239_not n12721_not ; n12722
g12467 and n12719_not n12722 ; n12723
g12468 and n12239_not n12723_not ; n12724
g12469 and b[36] n12228_not ; n12725
g12470 and n12222_not n12725 ; n12726
g12471 and n12230_not n12726_not ; n12727
g12472 and n12724_not n12727 ; n12728
g12473 and n12230_not n12728_not ; n12729
g12474 and b[37] n12219_not ; n12730
g12475 and n12213_not n12730 ; n12731
g12476 and n12221_not n12731_not ; n12732
g12477 and n12729_not n12732 ; n12733
g12478 and n12221_not n12733_not ; n12734
g12479 and b[38] n12210_not ; n12735
g12480 and n12204_not n12735 ; n12736
g12481 and n12212_not n12736_not ; n12737
g12482 and n12734_not n12737 ; n12738
g12483 and n12212_not n12738_not ; n12739
g12484 and b[39] n12201_not ; n12740
g12485 and n12195_not n12740 ; n12741
g12486 and n12203_not n12741_not ; n12742
g12487 and n12739_not n12742 ; n12743
g12488 and n12203_not n12743_not ; n12744
g12489 and b[40] n12192_not ; n12745
g12490 and n12186_not n12745 ; n12746
g12491 and n12194_not n12746_not ; n12747
g12492 and n12744_not n12747 ; n12748
g12493 and n12194_not n12748_not ; n12749
g12494 and n11635_not quotient[23]_not ; n12750
g12495 and n11637_not n12181 ; n12751
g12496 and n12177_not n12751 ; n12752
g12497 and n12178_not n12181_not ; n12753
g12498 and n12752_not n12753_not ; n12754
g12499 and quotient[23] n12754_not ; n12755
g12500 and n12750_not n12755_not ; n12756
g12501 and b[41]_not n12756_not ; n12757
g12502 and b[41] n12750_not ; n12758
g12503 and n12755_not n12758 ; n12759
g12504 and n290 n301 ; n12760
g12505 and n338 n12760 ; n12761
g12506 and n12759_not n12761 ; n12762
g12507 and n12757_not n12762 ; n12763
g12508 and n12749_not n12763 ; n12764
g12509 and n12184 n12756_not ; n12765
g12510 and n12764_not n12765_not ; quotient[22]
g12511 and n12203_not n12747 ; n12767
g12512 and n12743_not n12767 ; n12768
g12513 and n12744_not n12747_not ; n12769
g12514 and n12768_not n12769_not ; n12770
g12515 and quotient[22] n12770_not ; n12771
g12516 and n12193_not n12765_not ; n12772
g12517 and n12764_not n12772 ; n12773
g12518 and n12771_not n12773_not ; n12774
g12519 and n12194_not n12759_not ; n12775
g12520 and n12757_not n12775 ; n12776
g12521 and n12748_not n12776 ; n12777
g12522 and n12757_not n12759_not ; n12778
g12523 and n12749_not n12778_not ; n12779
g12524 and n12777_not n12779_not ; n12780
g12525 and quotient[22] n12780_not ; n12781
g12526 and n12756_not n12765_not ; n12782
g12527 and n12764_not n12782 ; n12783
g12528 and n12781_not n12783_not ; n12784
g12529 and b[42]_not n12784_not ; n12785
g12530 and b[41]_not n12774_not ; n12786
g12531 and n12212_not n12742 ; n12787
g12532 and n12738_not n12787 ; n12788
g12533 and n12739_not n12742_not ; n12789
g12534 and n12788_not n12789_not ; n12790
g12535 and quotient[22] n12790_not ; n12791
g12536 and n12202_not n12765_not ; n12792
g12537 and n12764_not n12792 ; n12793
g12538 and n12791_not n12793_not ; n12794
g12539 and b[40]_not n12794_not ; n12795
g12540 and n12221_not n12737 ; n12796
g12541 and n12733_not n12796 ; n12797
g12542 and n12734_not n12737_not ; n12798
g12543 and n12797_not n12798_not ; n12799
g12544 and quotient[22] n12799_not ; n12800
g12545 and n12211_not n12765_not ; n12801
g12546 and n12764_not n12801 ; n12802
g12547 and n12800_not n12802_not ; n12803
g12548 and b[39]_not n12803_not ; n12804
g12549 and n12230_not n12732 ; n12805
g12550 and n12728_not n12805 ; n12806
g12551 and n12729_not n12732_not ; n12807
g12552 and n12806_not n12807_not ; n12808
g12553 and quotient[22] n12808_not ; n12809
g12554 and n12220_not n12765_not ; n12810
g12555 and n12764_not n12810 ; n12811
g12556 and n12809_not n12811_not ; n12812
g12557 and b[38]_not n12812_not ; n12813
g12558 and n12239_not n12727 ; n12814
g12559 and n12723_not n12814 ; n12815
g12560 and n12724_not n12727_not ; n12816
g12561 and n12815_not n12816_not ; n12817
g12562 and quotient[22] n12817_not ; n12818
g12563 and n12229_not n12765_not ; n12819
g12564 and n12764_not n12819 ; n12820
g12565 and n12818_not n12820_not ; n12821
g12566 and b[37]_not n12821_not ; n12822
g12567 and n12248_not n12722 ; n12823
g12568 and n12718_not n12823 ; n12824
g12569 and n12719_not n12722_not ; n12825
g12570 and n12824_not n12825_not ; n12826
g12571 and quotient[22] n12826_not ; n12827
g12572 and n12238_not n12765_not ; n12828
g12573 and n12764_not n12828 ; n12829
g12574 and n12827_not n12829_not ; n12830
g12575 and b[36]_not n12830_not ; n12831
g12576 and n12257_not n12717 ; n12832
g12577 and n12713_not n12832 ; n12833
g12578 and n12714_not n12717_not ; n12834
g12579 and n12833_not n12834_not ; n12835
g12580 and quotient[22] n12835_not ; n12836
g12581 and n12247_not n12765_not ; n12837
g12582 and n12764_not n12837 ; n12838
g12583 and n12836_not n12838_not ; n12839
g12584 and b[35]_not n12839_not ; n12840
g12585 and n12266_not n12712 ; n12841
g12586 and n12708_not n12841 ; n12842
g12587 and n12709_not n12712_not ; n12843
g12588 and n12842_not n12843_not ; n12844
g12589 and quotient[22] n12844_not ; n12845
g12590 and n12256_not n12765_not ; n12846
g12591 and n12764_not n12846 ; n12847
g12592 and n12845_not n12847_not ; n12848
g12593 and b[34]_not n12848_not ; n12849
g12594 and n12275_not n12707 ; n12850
g12595 and n12703_not n12850 ; n12851
g12596 and n12704_not n12707_not ; n12852
g12597 and n12851_not n12852_not ; n12853
g12598 and quotient[22] n12853_not ; n12854
g12599 and n12265_not n12765_not ; n12855
g12600 and n12764_not n12855 ; n12856
g12601 and n12854_not n12856_not ; n12857
g12602 and b[33]_not n12857_not ; n12858
g12603 and n12284_not n12702 ; n12859
g12604 and n12698_not n12859 ; n12860
g12605 and n12699_not n12702_not ; n12861
g12606 and n12860_not n12861_not ; n12862
g12607 and quotient[22] n12862_not ; n12863
g12608 and n12274_not n12765_not ; n12864
g12609 and n12764_not n12864 ; n12865
g12610 and n12863_not n12865_not ; n12866
g12611 and b[32]_not n12866_not ; n12867
g12612 and n12293_not n12697 ; n12868
g12613 and n12693_not n12868 ; n12869
g12614 and n12694_not n12697_not ; n12870
g12615 and n12869_not n12870_not ; n12871
g12616 and quotient[22] n12871_not ; n12872
g12617 and n12283_not n12765_not ; n12873
g12618 and n12764_not n12873 ; n12874
g12619 and n12872_not n12874_not ; n12875
g12620 and b[31]_not n12875_not ; n12876
g12621 and n12302_not n12692 ; n12877
g12622 and n12688_not n12877 ; n12878
g12623 and n12689_not n12692_not ; n12879
g12624 and n12878_not n12879_not ; n12880
g12625 and quotient[22] n12880_not ; n12881
g12626 and n12292_not n12765_not ; n12882
g12627 and n12764_not n12882 ; n12883
g12628 and n12881_not n12883_not ; n12884
g12629 and b[30]_not n12884_not ; n12885
g12630 and n12311_not n12687 ; n12886
g12631 and n12683_not n12886 ; n12887
g12632 and n12684_not n12687_not ; n12888
g12633 and n12887_not n12888_not ; n12889
g12634 and quotient[22] n12889_not ; n12890
g12635 and n12301_not n12765_not ; n12891
g12636 and n12764_not n12891 ; n12892
g12637 and n12890_not n12892_not ; n12893
g12638 and b[29]_not n12893_not ; n12894
g12639 and n12320_not n12682 ; n12895
g12640 and n12678_not n12895 ; n12896
g12641 and n12679_not n12682_not ; n12897
g12642 and n12896_not n12897_not ; n12898
g12643 and quotient[22] n12898_not ; n12899
g12644 and n12310_not n12765_not ; n12900
g12645 and n12764_not n12900 ; n12901
g12646 and n12899_not n12901_not ; n12902
g12647 and b[28]_not n12902_not ; n12903
g12648 and n12329_not n12677 ; n12904
g12649 and n12673_not n12904 ; n12905
g12650 and n12674_not n12677_not ; n12906
g12651 and n12905_not n12906_not ; n12907
g12652 and quotient[22] n12907_not ; n12908
g12653 and n12319_not n12765_not ; n12909
g12654 and n12764_not n12909 ; n12910
g12655 and n12908_not n12910_not ; n12911
g12656 and b[27]_not n12911_not ; n12912
g12657 and n12338_not n12672 ; n12913
g12658 and n12668_not n12913 ; n12914
g12659 and n12669_not n12672_not ; n12915
g12660 and n12914_not n12915_not ; n12916
g12661 and quotient[22] n12916_not ; n12917
g12662 and n12328_not n12765_not ; n12918
g12663 and n12764_not n12918 ; n12919
g12664 and n12917_not n12919_not ; n12920
g12665 and b[26]_not n12920_not ; n12921
g12666 and n12347_not n12667 ; n12922
g12667 and n12663_not n12922 ; n12923
g12668 and n12664_not n12667_not ; n12924
g12669 and n12923_not n12924_not ; n12925
g12670 and quotient[22] n12925_not ; n12926
g12671 and n12337_not n12765_not ; n12927
g12672 and n12764_not n12927 ; n12928
g12673 and n12926_not n12928_not ; n12929
g12674 and b[25]_not n12929_not ; n12930
g12675 and n12356_not n12662 ; n12931
g12676 and n12658_not n12931 ; n12932
g12677 and n12659_not n12662_not ; n12933
g12678 and n12932_not n12933_not ; n12934
g12679 and quotient[22] n12934_not ; n12935
g12680 and n12346_not n12765_not ; n12936
g12681 and n12764_not n12936 ; n12937
g12682 and n12935_not n12937_not ; n12938
g12683 and b[24]_not n12938_not ; n12939
g12684 and n12365_not n12657 ; n12940
g12685 and n12653_not n12940 ; n12941
g12686 and n12654_not n12657_not ; n12942
g12687 and n12941_not n12942_not ; n12943
g12688 and quotient[22] n12943_not ; n12944
g12689 and n12355_not n12765_not ; n12945
g12690 and n12764_not n12945 ; n12946
g12691 and n12944_not n12946_not ; n12947
g12692 and b[23]_not n12947_not ; n12948
g12693 and n12374_not n12652 ; n12949
g12694 and n12648_not n12949 ; n12950
g12695 and n12649_not n12652_not ; n12951
g12696 and n12950_not n12951_not ; n12952
g12697 and quotient[22] n12952_not ; n12953
g12698 and n12364_not n12765_not ; n12954
g12699 and n12764_not n12954 ; n12955
g12700 and n12953_not n12955_not ; n12956
g12701 and b[22]_not n12956_not ; n12957
g12702 and n12383_not n12647 ; n12958
g12703 and n12643_not n12958 ; n12959
g12704 and n12644_not n12647_not ; n12960
g12705 and n12959_not n12960_not ; n12961
g12706 and quotient[22] n12961_not ; n12962
g12707 and n12373_not n12765_not ; n12963
g12708 and n12764_not n12963 ; n12964
g12709 and n12962_not n12964_not ; n12965
g12710 and b[21]_not n12965_not ; n12966
g12711 and n12392_not n12642 ; n12967
g12712 and n12638_not n12967 ; n12968
g12713 and n12639_not n12642_not ; n12969
g12714 and n12968_not n12969_not ; n12970
g12715 and quotient[22] n12970_not ; n12971
g12716 and n12382_not n12765_not ; n12972
g12717 and n12764_not n12972 ; n12973
g12718 and n12971_not n12973_not ; n12974
g12719 and b[20]_not n12974_not ; n12975
g12720 and n12401_not n12637 ; n12976
g12721 and n12633_not n12976 ; n12977
g12722 and n12634_not n12637_not ; n12978
g12723 and n12977_not n12978_not ; n12979
g12724 and quotient[22] n12979_not ; n12980
g12725 and n12391_not n12765_not ; n12981
g12726 and n12764_not n12981 ; n12982
g12727 and n12980_not n12982_not ; n12983
g12728 and b[19]_not n12983_not ; n12984
g12729 and n12410_not n12632 ; n12985
g12730 and n12628_not n12985 ; n12986
g12731 and n12629_not n12632_not ; n12987
g12732 and n12986_not n12987_not ; n12988
g12733 and quotient[22] n12988_not ; n12989
g12734 and n12400_not n12765_not ; n12990
g12735 and n12764_not n12990 ; n12991
g12736 and n12989_not n12991_not ; n12992
g12737 and b[18]_not n12992_not ; n12993
g12738 and n12419_not n12627 ; n12994
g12739 and n12623_not n12994 ; n12995
g12740 and n12624_not n12627_not ; n12996
g12741 and n12995_not n12996_not ; n12997
g12742 and quotient[22] n12997_not ; n12998
g12743 and n12409_not n12765_not ; n12999
g12744 and n12764_not n12999 ; n13000
g12745 and n12998_not n13000_not ; n13001
g12746 and b[17]_not n13001_not ; n13002
g12747 and n12428_not n12622 ; n13003
g12748 and n12618_not n13003 ; n13004
g12749 and n12619_not n12622_not ; n13005
g12750 and n13004_not n13005_not ; n13006
g12751 and quotient[22] n13006_not ; n13007
g12752 and n12418_not n12765_not ; n13008
g12753 and n12764_not n13008 ; n13009
g12754 and n13007_not n13009_not ; n13010
g12755 and b[16]_not n13010_not ; n13011
g12756 and n12437_not n12617 ; n13012
g12757 and n12613_not n13012 ; n13013
g12758 and n12614_not n12617_not ; n13014
g12759 and n13013_not n13014_not ; n13015
g12760 and quotient[22] n13015_not ; n13016
g12761 and n12427_not n12765_not ; n13017
g12762 and n12764_not n13017 ; n13018
g12763 and n13016_not n13018_not ; n13019
g12764 and b[15]_not n13019_not ; n13020
g12765 and n12446_not n12612 ; n13021
g12766 and n12608_not n13021 ; n13022
g12767 and n12609_not n12612_not ; n13023
g12768 and n13022_not n13023_not ; n13024
g12769 and quotient[22] n13024_not ; n13025
g12770 and n12436_not n12765_not ; n13026
g12771 and n12764_not n13026 ; n13027
g12772 and n13025_not n13027_not ; n13028
g12773 and b[14]_not n13028_not ; n13029
g12774 and n12455_not n12607 ; n13030
g12775 and n12603_not n13030 ; n13031
g12776 and n12604_not n12607_not ; n13032
g12777 and n13031_not n13032_not ; n13033
g12778 and quotient[22] n13033_not ; n13034
g12779 and n12445_not n12765_not ; n13035
g12780 and n12764_not n13035 ; n13036
g12781 and n13034_not n13036_not ; n13037
g12782 and b[13]_not n13037_not ; n13038
g12783 and n12464_not n12602 ; n13039
g12784 and n12598_not n13039 ; n13040
g12785 and n12599_not n12602_not ; n13041
g12786 and n13040_not n13041_not ; n13042
g12787 and quotient[22] n13042_not ; n13043
g12788 and n12454_not n12765_not ; n13044
g12789 and n12764_not n13044 ; n13045
g12790 and n13043_not n13045_not ; n13046
g12791 and b[12]_not n13046_not ; n13047
g12792 and n12473_not n12597 ; n13048
g12793 and n12593_not n13048 ; n13049
g12794 and n12594_not n12597_not ; n13050
g12795 and n13049_not n13050_not ; n13051
g12796 and quotient[22] n13051_not ; n13052
g12797 and n12463_not n12765_not ; n13053
g12798 and n12764_not n13053 ; n13054
g12799 and n13052_not n13054_not ; n13055
g12800 and b[11]_not n13055_not ; n13056
g12801 and n12482_not n12592 ; n13057
g12802 and n12588_not n13057 ; n13058
g12803 and n12589_not n12592_not ; n13059
g12804 and n13058_not n13059_not ; n13060
g12805 and quotient[22] n13060_not ; n13061
g12806 and n12472_not n12765_not ; n13062
g12807 and n12764_not n13062 ; n13063
g12808 and n13061_not n13063_not ; n13064
g12809 and b[10]_not n13064_not ; n13065
g12810 and n12491_not n12587 ; n13066
g12811 and n12583_not n13066 ; n13067
g12812 and n12584_not n12587_not ; n13068
g12813 and n13067_not n13068_not ; n13069
g12814 and quotient[22] n13069_not ; n13070
g12815 and n12481_not n12765_not ; n13071
g12816 and n12764_not n13071 ; n13072
g12817 and n13070_not n13072_not ; n13073
g12818 and b[9]_not n13073_not ; n13074
g12819 and n12500_not n12582 ; n13075
g12820 and n12578_not n13075 ; n13076
g12821 and n12579_not n12582_not ; n13077
g12822 and n13076_not n13077_not ; n13078
g12823 and quotient[22] n13078_not ; n13079
g12824 and n12490_not n12765_not ; n13080
g12825 and n12764_not n13080 ; n13081
g12826 and n13079_not n13081_not ; n13082
g12827 and b[8]_not n13082_not ; n13083
g12828 and n12509_not n12577 ; n13084
g12829 and n12573_not n13084 ; n13085
g12830 and n12574_not n12577_not ; n13086
g12831 and n13085_not n13086_not ; n13087
g12832 and quotient[22] n13087_not ; n13088
g12833 and n12499_not n12765_not ; n13089
g12834 and n12764_not n13089 ; n13090
g12835 and n13088_not n13090_not ; n13091
g12836 and b[7]_not n13091_not ; n13092
g12837 and n12518_not n12572 ; n13093
g12838 and n12568_not n13093 ; n13094
g12839 and n12569_not n12572_not ; n13095
g12840 and n13094_not n13095_not ; n13096
g12841 and quotient[22] n13096_not ; n13097
g12842 and n12508_not n12765_not ; n13098
g12843 and n12764_not n13098 ; n13099
g12844 and n13097_not n13099_not ; n13100
g12845 and b[6]_not n13100_not ; n13101
g12846 and n12527_not n12567 ; n13102
g12847 and n12563_not n13102 ; n13103
g12848 and n12564_not n12567_not ; n13104
g12849 and n13103_not n13104_not ; n13105
g12850 and quotient[22] n13105_not ; n13106
g12851 and n12517_not n12765_not ; n13107
g12852 and n12764_not n13107 ; n13108
g12853 and n13106_not n13108_not ; n13109
g12854 and b[5]_not n13109_not ; n13110
g12855 and n12535_not n12562 ; n13111
g12856 and n12558_not n13111 ; n13112
g12857 and n12559_not n12562_not ; n13113
g12858 and n13112_not n13113_not ; n13114
g12859 and quotient[22] n13114_not ; n13115
g12860 and n12526_not n12765_not ; n13116
g12861 and n12764_not n13116 ; n13117
g12862 and n13115_not n13117_not ; n13118
g12863 and b[4]_not n13118_not ; n13119
g12864 and n12553_not n12557 ; n13120
g12865 and n12552_not n13120 ; n13121
g12866 and n12554_not n12557_not ; n13122
g12867 and n13121_not n13122_not ; n13123
g12868 and quotient[22] n13123_not ; n13124
g12869 and n12534_not n12765_not ; n13125
g12870 and n12764_not n13125 ; n13126
g12871 and n13124_not n13126_not ; n13127
g12872 and b[3]_not n13127_not ; n13128
g12873 and n12549_not n12551 ; n13129
g12874 and n12547_not n13129 ; n13130
g12875 and n12552_not n13130_not ; n13131
g12876 and quotient[22] n13131 ; n13132
g12877 and n12546_not n12765_not ; n13133
g12878 and n12764_not n13133 ; n13134
g12879 and n13132_not n13134_not ; n13135
g12880 and b[2]_not n13135_not ; n13136
g12881 and b[0] quotient[22] ; n13137
g12882 and a[22] n13137_not ; n13138
g12883 and n12551 quotient[22] ; n13139
g12884 and n13138_not n13139_not ; n13140
g12885 and b[1] n13140_not ; n13141
g12886 and b[1]_not n13139_not ; n13142
g12887 and n13138_not n13142 ; n13143
g12888 and n13141_not n13143_not ; n13144
g12889 and a[21]_not b[0] ; n13145
g12890 and n13144_not n13145_not ; n13146
g12891 and b[1]_not n13140_not ; n13147
g12892 and n13146_not n13147_not ; n13148
g12893 and b[2] n13134_not ; n13149
g12894 and n13132_not n13149 ; n13150
g12895 and n13136_not n13150_not ; n13151
g12896 and n13148_not n13151 ; n13152
g12897 and n13136_not n13152_not ; n13153
g12898 and b[3] n13126_not ; n13154
g12899 and n13124_not n13154 ; n13155
g12900 and n13128_not n13155_not ; n13156
g12901 and n13153_not n13156 ; n13157
g12902 and n13128_not n13157_not ; n13158
g12903 and b[4] n13117_not ; n13159
g12904 and n13115_not n13159 ; n13160
g12905 and n13119_not n13160_not ; n13161
g12906 and n13158_not n13161 ; n13162
g12907 and n13119_not n13162_not ; n13163
g12908 and b[5] n13108_not ; n13164
g12909 and n13106_not n13164 ; n13165
g12910 and n13110_not n13165_not ; n13166
g12911 and n13163_not n13166 ; n13167
g12912 and n13110_not n13167_not ; n13168
g12913 and b[6] n13099_not ; n13169
g12914 and n13097_not n13169 ; n13170
g12915 and n13101_not n13170_not ; n13171
g12916 and n13168_not n13171 ; n13172
g12917 and n13101_not n13172_not ; n13173
g12918 and b[7] n13090_not ; n13174
g12919 and n13088_not n13174 ; n13175
g12920 and n13092_not n13175_not ; n13176
g12921 and n13173_not n13176 ; n13177
g12922 and n13092_not n13177_not ; n13178
g12923 and b[8] n13081_not ; n13179
g12924 and n13079_not n13179 ; n13180
g12925 and n13083_not n13180_not ; n13181
g12926 and n13178_not n13181 ; n13182
g12927 and n13083_not n13182_not ; n13183
g12928 and b[9] n13072_not ; n13184
g12929 and n13070_not n13184 ; n13185
g12930 and n13074_not n13185_not ; n13186
g12931 and n13183_not n13186 ; n13187
g12932 and n13074_not n13187_not ; n13188
g12933 and b[10] n13063_not ; n13189
g12934 and n13061_not n13189 ; n13190
g12935 and n13065_not n13190_not ; n13191
g12936 and n13188_not n13191 ; n13192
g12937 and n13065_not n13192_not ; n13193
g12938 and b[11] n13054_not ; n13194
g12939 and n13052_not n13194 ; n13195
g12940 and n13056_not n13195_not ; n13196
g12941 and n13193_not n13196 ; n13197
g12942 and n13056_not n13197_not ; n13198
g12943 and b[12] n13045_not ; n13199
g12944 and n13043_not n13199 ; n13200
g12945 and n13047_not n13200_not ; n13201
g12946 and n13198_not n13201 ; n13202
g12947 and n13047_not n13202_not ; n13203
g12948 and b[13] n13036_not ; n13204
g12949 and n13034_not n13204 ; n13205
g12950 and n13038_not n13205_not ; n13206
g12951 and n13203_not n13206 ; n13207
g12952 and n13038_not n13207_not ; n13208
g12953 and b[14] n13027_not ; n13209
g12954 and n13025_not n13209 ; n13210
g12955 and n13029_not n13210_not ; n13211
g12956 and n13208_not n13211 ; n13212
g12957 and n13029_not n13212_not ; n13213
g12958 and b[15] n13018_not ; n13214
g12959 and n13016_not n13214 ; n13215
g12960 and n13020_not n13215_not ; n13216
g12961 and n13213_not n13216 ; n13217
g12962 and n13020_not n13217_not ; n13218
g12963 and b[16] n13009_not ; n13219
g12964 and n13007_not n13219 ; n13220
g12965 and n13011_not n13220_not ; n13221
g12966 and n13218_not n13221 ; n13222
g12967 and n13011_not n13222_not ; n13223
g12968 and b[17] n13000_not ; n13224
g12969 and n12998_not n13224 ; n13225
g12970 and n13002_not n13225_not ; n13226
g12971 and n13223_not n13226 ; n13227
g12972 and n13002_not n13227_not ; n13228
g12973 and b[18] n12991_not ; n13229
g12974 and n12989_not n13229 ; n13230
g12975 and n12993_not n13230_not ; n13231
g12976 and n13228_not n13231 ; n13232
g12977 and n12993_not n13232_not ; n13233
g12978 and b[19] n12982_not ; n13234
g12979 and n12980_not n13234 ; n13235
g12980 and n12984_not n13235_not ; n13236
g12981 and n13233_not n13236 ; n13237
g12982 and n12984_not n13237_not ; n13238
g12983 and b[20] n12973_not ; n13239
g12984 and n12971_not n13239 ; n13240
g12985 and n12975_not n13240_not ; n13241
g12986 and n13238_not n13241 ; n13242
g12987 and n12975_not n13242_not ; n13243
g12988 and b[21] n12964_not ; n13244
g12989 and n12962_not n13244 ; n13245
g12990 and n12966_not n13245_not ; n13246
g12991 and n13243_not n13246 ; n13247
g12992 and n12966_not n13247_not ; n13248
g12993 and b[22] n12955_not ; n13249
g12994 and n12953_not n13249 ; n13250
g12995 and n12957_not n13250_not ; n13251
g12996 and n13248_not n13251 ; n13252
g12997 and n12957_not n13252_not ; n13253
g12998 and b[23] n12946_not ; n13254
g12999 and n12944_not n13254 ; n13255
g13000 and n12948_not n13255_not ; n13256
g13001 and n13253_not n13256 ; n13257
g13002 and n12948_not n13257_not ; n13258
g13003 and b[24] n12937_not ; n13259
g13004 and n12935_not n13259 ; n13260
g13005 and n12939_not n13260_not ; n13261
g13006 and n13258_not n13261 ; n13262
g13007 and n12939_not n13262_not ; n13263
g13008 and b[25] n12928_not ; n13264
g13009 and n12926_not n13264 ; n13265
g13010 and n12930_not n13265_not ; n13266
g13011 and n13263_not n13266 ; n13267
g13012 and n12930_not n13267_not ; n13268
g13013 and b[26] n12919_not ; n13269
g13014 and n12917_not n13269 ; n13270
g13015 and n12921_not n13270_not ; n13271
g13016 and n13268_not n13271 ; n13272
g13017 and n12921_not n13272_not ; n13273
g13018 and b[27] n12910_not ; n13274
g13019 and n12908_not n13274 ; n13275
g13020 and n12912_not n13275_not ; n13276
g13021 and n13273_not n13276 ; n13277
g13022 and n12912_not n13277_not ; n13278
g13023 and b[28] n12901_not ; n13279
g13024 and n12899_not n13279 ; n13280
g13025 and n12903_not n13280_not ; n13281
g13026 and n13278_not n13281 ; n13282
g13027 and n12903_not n13282_not ; n13283
g13028 and b[29] n12892_not ; n13284
g13029 and n12890_not n13284 ; n13285
g13030 and n12894_not n13285_not ; n13286
g13031 and n13283_not n13286 ; n13287
g13032 and n12894_not n13287_not ; n13288
g13033 and b[30] n12883_not ; n13289
g13034 and n12881_not n13289 ; n13290
g13035 and n12885_not n13290_not ; n13291
g13036 and n13288_not n13291 ; n13292
g13037 and n12885_not n13292_not ; n13293
g13038 and b[31] n12874_not ; n13294
g13039 and n12872_not n13294 ; n13295
g13040 and n12876_not n13295_not ; n13296
g13041 and n13293_not n13296 ; n13297
g13042 and n12876_not n13297_not ; n13298
g13043 and b[32] n12865_not ; n13299
g13044 and n12863_not n13299 ; n13300
g13045 and n12867_not n13300_not ; n13301
g13046 and n13298_not n13301 ; n13302
g13047 and n12867_not n13302_not ; n13303
g13048 and b[33] n12856_not ; n13304
g13049 and n12854_not n13304 ; n13305
g13050 and n12858_not n13305_not ; n13306
g13051 and n13303_not n13306 ; n13307
g13052 and n12858_not n13307_not ; n13308
g13053 and b[34] n12847_not ; n13309
g13054 and n12845_not n13309 ; n13310
g13055 and n12849_not n13310_not ; n13311
g13056 and n13308_not n13311 ; n13312
g13057 and n12849_not n13312_not ; n13313
g13058 and b[35] n12838_not ; n13314
g13059 and n12836_not n13314 ; n13315
g13060 and n12840_not n13315_not ; n13316
g13061 and n13313_not n13316 ; n13317
g13062 and n12840_not n13317_not ; n13318
g13063 and b[36] n12829_not ; n13319
g13064 and n12827_not n13319 ; n13320
g13065 and n12831_not n13320_not ; n13321
g13066 and n13318_not n13321 ; n13322
g13067 and n12831_not n13322_not ; n13323
g13068 and b[37] n12820_not ; n13324
g13069 and n12818_not n13324 ; n13325
g13070 and n12822_not n13325_not ; n13326
g13071 and n13323_not n13326 ; n13327
g13072 and n12822_not n13327_not ; n13328
g13073 and b[38] n12811_not ; n13329
g13074 and n12809_not n13329 ; n13330
g13075 and n12813_not n13330_not ; n13331
g13076 and n13328_not n13331 ; n13332
g13077 and n12813_not n13332_not ; n13333
g13078 and b[39] n12802_not ; n13334
g13079 and n12800_not n13334 ; n13335
g13080 and n12804_not n13335_not ; n13336
g13081 and n13333_not n13336 ; n13337
g13082 and n12804_not n13337_not ; n13338
g13083 and b[40] n12793_not ; n13339
g13084 and n12791_not n13339 ; n13340
g13085 and n12795_not n13340_not ; n13341
g13086 and n13338_not n13341 ; n13342
g13087 and n12795_not n13342_not ; n13343
g13088 and b[41] n12773_not ; n13344
g13089 and n12771_not n13344 ; n13345
g13090 and n12786_not n13345_not ; n13346
g13091 and n13343_not n13346 ; n13347
g13092 and n12786_not n13347_not ; n13348
g13093 and b[42] n12783_not ; n13349
g13094 and n12781_not n13349 ; n13350
g13095 and n12785_not n13350_not ; n13351
g13096 and n13348_not n13351 ; n13352
g13097 and n12785_not n13352_not ; n13353
g13098 and n418 n420 ; n13354
g13099 and n408 n13354 ; n13355
g13100 and n13353_not n13355 ; quotient[21]
g13101 and n12774_not quotient[21]_not ; n13357
g13102 and n12795_not n13346 ; n13358
g13103 and n13342_not n13358 ; n13359
g13104 and n13343_not n13346_not ; n13360
g13105 and n13359_not n13360_not ; n13361
g13106 and n13355 n13361_not ; n13362
g13107 and n13353_not n13362 ; n13363
g13108 and n13357_not n13363_not ; n13364
g13109 and b[42]_not n13364_not ; n13365
g13110 and n12794_not quotient[21]_not ; n13366
g13111 and n12804_not n13341 ; n13367
g13112 and n13337_not n13367 ; n13368
g13113 and n13338_not n13341_not ; n13369
g13114 and n13368_not n13369_not ; n13370
g13115 and n13355 n13370_not ; n13371
g13116 and n13353_not n13371 ; n13372
g13117 and n13366_not n13372_not ; n13373
g13118 and b[41]_not n13373_not ; n13374
g13119 and n12803_not quotient[21]_not ; n13375
g13120 and n12813_not n13336 ; n13376
g13121 and n13332_not n13376 ; n13377
g13122 and n13333_not n13336_not ; n13378
g13123 and n13377_not n13378_not ; n13379
g13124 and n13355 n13379_not ; n13380
g13125 and n13353_not n13380 ; n13381
g13126 and n13375_not n13381_not ; n13382
g13127 and b[40]_not n13382_not ; n13383
g13128 and n12812_not quotient[21]_not ; n13384
g13129 and n12822_not n13331 ; n13385
g13130 and n13327_not n13385 ; n13386
g13131 and n13328_not n13331_not ; n13387
g13132 and n13386_not n13387_not ; n13388
g13133 and n13355 n13388_not ; n13389
g13134 and n13353_not n13389 ; n13390
g13135 and n13384_not n13390_not ; n13391
g13136 and b[39]_not n13391_not ; n13392
g13137 and n12821_not quotient[21]_not ; n13393
g13138 and n12831_not n13326 ; n13394
g13139 and n13322_not n13394 ; n13395
g13140 and n13323_not n13326_not ; n13396
g13141 and n13395_not n13396_not ; n13397
g13142 and n13355 n13397_not ; n13398
g13143 and n13353_not n13398 ; n13399
g13144 and n13393_not n13399_not ; n13400
g13145 and b[38]_not n13400_not ; n13401
g13146 and n12830_not quotient[21]_not ; n13402
g13147 and n12840_not n13321 ; n13403
g13148 and n13317_not n13403 ; n13404
g13149 and n13318_not n13321_not ; n13405
g13150 and n13404_not n13405_not ; n13406
g13151 and n13355 n13406_not ; n13407
g13152 and n13353_not n13407 ; n13408
g13153 and n13402_not n13408_not ; n13409
g13154 and b[37]_not n13409_not ; n13410
g13155 and n12839_not quotient[21]_not ; n13411
g13156 and n12849_not n13316 ; n13412
g13157 and n13312_not n13412 ; n13413
g13158 and n13313_not n13316_not ; n13414
g13159 and n13413_not n13414_not ; n13415
g13160 and n13355 n13415_not ; n13416
g13161 and n13353_not n13416 ; n13417
g13162 and n13411_not n13417_not ; n13418
g13163 and b[36]_not n13418_not ; n13419
g13164 and n12848_not quotient[21]_not ; n13420
g13165 and n12858_not n13311 ; n13421
g13166 and n13307_not n13421 ; n13422
g13167 and n13308_not n13311_not ; n13423
g13168 and n13422_not n13423_not ; n13424
g13169 and n13355 n13424_not ; n13425
g13170 and n13353_not n13425 ; n13426
g13171 and n13420_not n13426_not ; n13427
g13172 and b[35]_not n13427_not ; n13428
g13173 and n12857_not quotient[21]_not ; n13429
g13174 and n12867_not n13306 ; n13430
g13175 and n13302_not n13430 ; n13431
g13176 and n13303_not n13306_not ; n13432
g13177 and n13431_not n13432_not ; n13433
g13178 and n13355 n13433_not ; n13434
g13179 and n13353_not n13434 ; n13435
g13180 and n13429_not n13435_not ; n13436
g13181 and b[34]_not n13436_not ; n13437
g13182 and n12866_not quotient[21]_not ; n13438
g13183 and n12876_not n13301 ; n13439
g13184 and n13297_not n13439 ; n13440
g13185 and n13298_not n13301_not ; n13441
g13186 and n13440_not n13441_not ; n13442
g13187 and n13355 n13442_not ; n13443
g13188 and n13353_not n13443 ; n13444
g13189 and n13438_not n13444_not ; n13445
g13190 and b[33]_not n13445_not ; n13446
g13191 and n12875_not quotient[21]_not ; n13447
g13192 and n12885_not n13296 ; n13448
g13193 and n13292_not n13448 ; n13449
g13194 and n13293_not n13296_not ; n13450
g13195 and n13449_not n13450_not ; n13451
g13196 and n13355 n13451_not ; n13452
g13197 and n13353_not n13452 ; n13453
g13198 and n13447_not n13453_not ; n13454
g13199 and b[32]_not n13454_not ; n13455
g13200 and n12884_not quotient[21]_not ; n13456
g13201 and n12894_not n13291 ; n13457
g13202 and n13287_not n13457 ; n13458
g13203 and n13288_not n13291_not ; n13459
g13204 and n13458_not n13459_not ; n13460
g13205 and n13355 n13460_not ; n13461
g13206 and n13353_not n13461 ; n13462
g13207 and n13456_not n13462_not ; n13463
g13208 and b[31]_not n13463_not ; n13464
g13209 and n12893_not quotient[21]_not ; n13465
g13210 and n12903_not n13286 ; n13466
g13211 and n13282_not n13466 ; n13467
g13212 and n13283_not n13286_not ; n13468
g13213 and n13467_not n13468_not ; n13469
g13214 and n13355 n13469_not ; n13470
g13215 and n13353_not n13470 ; n13471
g13216 and n13465_not n13471_not ; n13472
g13217 and b[30]_not n13472_not ; n13473
g13218 and n12902_not quotient[21]_not ; n13474
g13219 and n12912_not n13281 ; n13475
g13220 and n13277_not n13475 ; n13476
g13221 and n13278_not n13281_not ; n13477
g13222 and n13476_not n13477_not ; n13478
g13223 and n13355 n13478_not ; n13479
g13224 and n13353_not n13479 ; n13480
g13225 and n13474_not n13480_not ; n13481
g13226 and b[29]_not n13481_not ; n13482
g13227 and n12911_not quotient[21]_not ; n13483
g13228 and n12921_not n13276 ; n13484
g13229 and n13272_not n13484 ; n13485
g13230 and n13273_not n13276_not ; n13486
g13231 and n13485_not n13486_not ; n13487
g13232 and n13355 n13487_not ; n13488
g13233 and n13353_not n13488 ; n13489
g13234 and n13483_not n13489_not ; n13490
g13235 and b[28]_not n13490_not ; n13491
g13236 and n12920_not quotient[21]_not ; n13492
g13237 and n12930_not n13271 ; n13493
g13238 and n13267_not n13493 ; n13494
g13239 and n13268_not n13271_not ; n13495
g13240 and n13494_not n13495_not ; n13496
g13241 and n13355 n13496_not ; n13497
g13242 and n13353_not n13497 ; n13498
g13243 and n13492_not n13498_not ; n13499
g13244 and b[27]_not n13499_not ; n13500
g13245 and n12929_not quotient[21]_not ; n13501
g13246 and n12939_not n13266 ; n13502
g13247 and n13262_not n13502 ; n13503
g13248 and n13263_not n13266_not ; n13504
g13249 and n13503_not n13504_not ; n13505
g13250 and n13355 n13505_not ; n13506
g13251 and n13353_not n13506 ; n13507
g13252 and n13501_not n13507_not ; n13508
g13253 and b[26]_not n13508_not ; n13509
g13254 and n12938_not quotient[21]_not ; n13510
g13255 and n12948_not n13261 ; n13511
g13256 and n13257_not n13511 ; n13512
g13257 and n13258_not n13261_not ; n13513
g13258 and n13512_not n13513_not ; n13514
g13259 and n13355 n13514_not ; n13515
g13260 and n13353_not n13515 ; n13516
g13261 and n13510_not n13516_not ; n13517
g13262 and b[25]_not n13517_not ; n13518
g13263 and n12947_not quotient[21]_not ; n13519
g13264 and n12957_not n13256 ; n13520
g13265 and n13252_not n13520 ; n13521
g13266 and n13253_not n13256_not ; n13522
g13267 and n13521_not n13522_not ; n13523
g13268 and n13355 n13523_not ; n13524
g13269 and n13353_not n13524 ; n13525
g13270 and n13519_not n13525_not ; n13526
g13271 and b[24]_not n13526_not ; n13527
g13272 and n12956_not quotient[21]_not ; n13528
g13273 and n12966_not n13251 ; n13529
g13274 and n13247_not n13529 ; n13530
g13275 and n13248_not n13251_not ; n13531
g13276 and n13530_not n13531_not ; n13532
g13277 and n13355 n13532_not ; n13533
g13278 and n13353_not n13533 ; n13534
g13279 and n13528_not n13534_not ; n13535
g13280 and b[23]_not n13535_not ; n13536
g13281 and n12965_not quotient[21]_not ; n13537
g13282 and n12975_not n13246 ; n13538
g13283 and n13242_not n13538 ; n13539
g13284 and n13243_not n13246_not ; n13540
g13285 and n13539_not n13540_not ; n13541
g13286 and n13355 n13541_not ; n13542
g13287 and n13353_not n13542 ; n13543
g13288 and n13537_not n13543_not ; n13544
g13289 and b[22]_not n13544_not ; n13545
g13290 and n12974_not quotient[21]_not ; n13546
g13291 and n12984_not n13241 ; n13547
g13292 and n13237_not n13547 ; n13548
g13293 and n13238_not n13241_not ; n13549
g13294 and n13548_not n13549_not ; n13550
g13295 and n13355 n13550_not ; n13551
g13296 and n13353_not n13551 ; n13552
g13297 and n13546_not n13552_not ; n13553
g13298 and b[21]_not n13553_not ; n13554
g13299 and n12983_not quotient[21]_not ; n13555
g13300 and n12993_not n13236 ; n13556
g13301 and n13232_not n13556 ; n13557
g13302 and n13233_not n13236_not ; n13558
g13303 and n13557_not n13558_not ; n13559
g13304 and n13355 n13559_not ; n13560
g13305 and n13353_not n13560 ; n13561
g13306 and n13555_not n13561_not ; n13562
g13307 and b[20]_not n13562_not ; n13563
g13308 and n12992_not quotient[21]_not ; n13564
g13309 and n13002_not n13231 ; n13565
g13310 and n13227_not n13565 ; n13566
g13311 and n13228_not n13231_not ; n13567
g13312 and n13566_not n13567_not ; n13568
g13313 and n13355 n13568_not ; n13569
g13314 and n13353_not n13569 ; n13570
g13315 and n13564_not n13570_not ; n13571
g13316 and b[19]_not n13571_not ; n13572
g13317 and n13001_not quotient[21]_not ; n13573
g13318 and n13011_not n13226 ; n13574
g13319 and n13222_not n13574 ; n13575
g13320 and n13223_not n13226_not ; n13576
g13321 and n13575_not n13576_not ; n13577
g13322 and n13355 n13577_not ; n13578
g13323 and n13353_not n13578 ; n13579
g13324 and n13573_not n13579_not ; n13580
g13325 and b[18]_not n13580_not ; n13581
g13326 and n13010_not quotient[21]_not ; n13582
g13327 and n13020_not n13221 ; n13583
g13328 and n13217_not n13583 ; n13584
g13329 and n13218_not n13221_not ; n13585
g13330 and n13584_not n13585_not ; n13586
g13331 and n13355 n13586_not ; n13587
g13332 and n13353_not n13587 ; n13588
g13333 and n13582_not n13588_not ; n13589
g13334 and b[17]_not n13589_not ; n13590
g13335 and n13019_not quotient[21]_not ; n13591
g13336 and n13029_not n13216 ; n13592
g13337 and n13212_not n13592 ; n13593
g13338 and n13213_not n13216_not ; n13594
g13339 and n13593_not n13594_not ; n13595
g13340 and n13355 n13595_not ; n13596
g13341 and n13353_not n13596 ; n13597
g13342 and n13591_not n13597_not ; n13598
g13343 and b[16]_not n13598_not ; n13599
g13344 and n13028_not quotient[21]_not ; n13600
g13345 and n13038_not n13211 ; n13601
g13346 and n13207_not n13601 ; n13602
g13347 and n13208_not n13211_not ; n13603
g13348 and n13602_not n13603_not ; n13604
g13349 and n13355 n13604_not ; n13605
g13350 and n13353_not n13605 ; n13606
g13351 and n13600_not n13606_not ; n13607
g13352 and b[15]_not n13607_not ; n13608
g13353 and n13037_not quotient[21]_not ; n13609
g13354 and n13047_not n13206 ; n13610
g13355 and n13202_not n13610 ; n13611
g13356 and n13203_not n13206_not ; n13612
g13357 and n13611_not n13612_not ; n13613
g13358 and n13355 n13613_not ; n13614
g13359 and n13353_not n13614 ; n13615
g13360 and n13609_not n13615_not ; n13616
g13361 and b[14]_not n13616_not ; n13617
g13362 and n13046_not quotient[21]_not ; n13618
g13363 and n13056_not n13201 ; n13619
g13364 and n13197_not n13619 ; n13620
g13365 and n13198_not n13201_not ; n13621
g13366 and n13620_not n13621_not ; n13622
g13367 and n13355 n13622_not ; n13623
g13368 and n13353_not n13623 ; n13624
g13369 and n13618_not n13624_not ; n13625
g13370 and b[13]_not n13625_not ; n13626
g13371 and n13055_not quotient[21]_not ; n13627
g13372 and n13065_not n13196 ; n13628
g13373 and n13192_not n13628 ; n13629
g13374 and n13193_not n13196_not ; n13630
g13375 and n13629_not n13630_not ; n13631
g13376 and n13355 n13631_not ; n13632
g13377 and n13353_not n13632 ; n13633
g13378 and n13627_not n13633_not ; n13634
g13379 and b[12]_not n13634_not ; n13635
g13380 and n13064_not quotient[21]_not ; n13636
g13381 and n13074_not n13191 ; n13637
g13382 and n13187_not n13637 ; n13638
g13383 and n13188_not n13191_not ; n13639
g13384 and n13638_not n13639_not ; n13640
g13385 and n13355 n13640_not ; n13641
g13386 and n13353_not n13641 ; n13642
g13387 and n13636_not n13642_not ; n13643
g13388 and b[11]_not n13643_not ; n13644
g13389 and n13073_not quotient[21]_not ; n13645
g13390 and n13083_not n13186 ; n13646
g13391 and n13182_not n13646 ; n13647
g13392 and n13183_not n13186_not ; n13648
g13393 and n13647_not n13648_not ; n13649
g13394 and n13355 n13649_not ; n13650
g13395 and n13353_not n13650 ; n13651
g13396 and n13645_not n13651_not ; n13652
g13397 and b[10]_not n13652_not ; n13653
g13398 and n13082_not quotient[21]_not ; n13654
g13399 and n13092_not n13181 ; n13655
g13400 and n13177_not n13655 ; n13656
g13401 and n13178_not n13181_not ; n13657
g13402 and n13656_not n13657_not ; n13658
g13403 and n13355 n13658_not ; n13659
g13404 and n13353_not n13659 ; n13660
g13405 and n13654_not n13660_not ; n13661
g13406 and b[9]_not n13661_not ; n13662
g13407 and n13091_not quotient[21]_not ; n13663
g13408 and n13101_not n13176 ; n13664
g13409 and n13172_not n13664 ; n13665
g13410 and n13173_not n13176_not ; n13666
g13411 and n13665_not n13666_not ; n13667
g13412 and n13355 n13667_not ; n13668
g13413 and n13353_not n13668 ; n13669
g13414 and n13663_not n13669_not ; n13670
g13415 and b[8]_not n13670_not ; n13671
g13416 and n13100_not quotient[21]_not ; n13672
g13417 and n13110_not n13171 ; n13673
g13418 and n13167_not n13673 ; n13674
g13419 and n13168_not n13171_not ; n13675
g13420 and n13674_not n13675_not ; n13676
g13421 and n13355 n13676_not ; n13677
g13422 and n13353_not n13677 ; n13678
g13423 and n13672_not n13678_not ; n13679
g13424 and b[7]_not n13679_not ; n13680
g13425 and n13109_not quotient[21]_not ; n13681
g13426 and n13119_not n13166 ; n13682
g13427 and n13162_not n13682 ; n13683
g13428 and n13163_not n13166_not ; n13684
g13429 and n13683_not n13684_not ; n13685
g13430 and n13355 n13685_not ; n13686
g13431 and n13353_not n13686 ; n13687
g13432 and n13681_not n13687_not ; n13688
g13433 and b[6]_not n13688_not ; n13689
g13434 and n13118_not quotient[21]_not ; n13690
g13435 and n13128_not n13161 ; n13691
g13436 and n13157_not n13691 ; n13692
g13437 and n13158_not n13161_not ; n13693
g13438 and n13692_not n13693_not ; n13694
g13439 and n13355 n13694_not ; n13695
g13440 and n13353_not n13695 ; n13696
g13441 and n13690_not n13696_not ; n13697
g13442 and b[5]_not n13697_not ; n13698
g13443 and n13127_not quotient[21]_not ; n13699
g13444 and n13136_not n13156 ; n13700
g13445 and n13152_not n13700 ; n13701
g13446 and n13153_not n13156_not ; n13702
g13447 and n13701_not n13702_not ; n13703
g13448 and n13355 n13703_not ; n13704
g13449 and n13353_not n13704 ; n13705
g13450 and n13699_not n13705_not ; n13706
g13451 and b[4]_not n13706_not ; n13707
g13452 and n13135_not quotient[21]_not ; n13708
g13453 and n13147_not n13151 ; n13709
g13454 and n13146_not n13709 ; n13710
g13455 and n13148_not n13151_not ; n13711
g13456 and n13710_not n13711_not ; n13712
g13457 and n13355 n13712_not ; n13713
g13458 and n13353_not n13713 ; n13714
g13459 and n13708_not n13714_not ; n13715
g13460 and b[3]_not n13715_not ; n13716
g13461 and n13140_not quotient[21]_not ; n13717
g13462 and n13143_not n13145 ; n13718
g13463 and n13141_not n13718 ; n13719
g13464 and n13355 n13719_not ; n13720
g13465 and n13146_not n13720 ; n13721
g13466 and n13353_not n13721 ; n13722
g13467 and n13717_not n13722_not ; n13723
g13468 and b[2]_not n13723_not ; n13724
g13469 and b[0] b[43]_not ; n13725
g13470 and n301 n13725 ; n13726
g13471 and n338 n13726 ; n13727
g13472 and n13353_not n13727 ; n13728
g13473 and a[21] n13728_not ; n13729
g13474 and n420 n13145 ; n13730
g13475 and n418 n13730 ; n13731
g13476 and n408 n13731 ; n13732
g13477 and n13353_not n13732 ; n13733
g13478 and n13729_not n13733_not ; n13734
g13479 and b[1] n13734_not ; n13735
g13480 and b[1]_not n13733_not ; n13736
g13481 and n13729_not n13736 ; n13737
g13482 and n13735_not n13737_not ; n13738
g13483 and a[20]_not b[0] ; n13739
g13484 and n13738_not n13739_not ; n13740
g13485 and b[1]_not n13734_not ; n13741
g13486 and n13740_not n13741_not ; n13742
g13487 and b[2] n13722_not ; n13743
g13488 and n13717_not n13743 ; n13744
g13489 and n13724_not n13744_not ; n13745
g13490 and n13742_not n13745 ; n13746
g13491 and n13724_not n13746_not ; n13747
g13492 and b[3] n13714_not ; n13748
g13493 and n13708_not n13748 ; n13749
g13494 and n13716_not n13749_not ; n13750
g13495 and n13747_not n13750 ; n13751
g13496 and n13716_not n13751_not ; n13752
g13497 and b[4] n13705_not ; n13753
g13498 and n13699_not n13753 ; n13754
g13499 and n13707_not n13754_not ; n13755
g13500 and n13752_not n13755 ; n13756
g13501 and n13707_not n13756_not ; n13757
g13502 and b[5] n13696_not ; n13758
g13503 and n13690_not n13758 ; n13759
g13504 and n13698_not n13759_not ; n13760
g13505 and n13757_not n13760 ; n13761
g13506 and n13698_not n13761_not ; n13762
g13507 and b[6] n13687_not ; n13763
g13508 and n13681_not n13763 ; n13764
g13509 and n13689_not n13764_not ; n13765
g13510 and n13762_not n13765 ; n13766
g13511 and n13689_not n13766_not ; n13767
g13512 and b[7] n13678_not ; n13768
g13513 and n13672_not n13768 ; n13769
g13514 and n13680_not n13769_not ; n13770
g13515 and n13767_not n13770 ; n13771
g13516 and n13680_not n13771_not ; n13772
g13517 and b[8] n13669_not ; n13773
g13518 and n13663_not n13773 ; n13774
g13519 and n13671_not n13774_not ; n13775
g13520 and n13772_not n13775 ; n13776
g13521 and n13671_not n13776_not ; n13777
g13522 and b[9] n13660_not ; n13778
g13523 and n13654_not n13778 ; n13779
g13524 and n13662_not n13779_not ; n13780
g13525 and n13777_not n13780 ; n13781
g13526 and n13662_not n13781_not ; n13782
g13527 and b[10] n13651_not ; n13783
g13528 and n13645_not n13783 ; n13784
g13529 and n13653_not n13784_not ; n13785
g13530 and n13782_not n13785 ; n13786
g13531 and n13653_not n13786_not ; n13787
g13532 and b[11] n13642_not ; n13788
g13533 and n13636_not n13788 ; n13789
g13534 and n13644_not n13789_not ; n13790
g13535 and n13787_not n13790 ; n13791
g13536 and n13644_not n13791_not ; n13792
g13537 and b[12] n13633_not ; n13793
g13538 and n13627_not n13793 ; n13794
g13539 and n13635_not n13794_not ; n13795
g13540 and n13792_not n13795 ; n13796
g13541 and n13635_not n13796_not ; n13797
g13542 and b[13] n13624_not ; n13798
g13543 and n13618_not n13798 ; n13799
g13544 and n13626_not n13799_not ; n13800
g13545 and n13797_not n13800 ; n13801
g13546 and n13626_not n13801_not ; n13802
g13547 and b[14] n13615_not ; n13803
g13548 and n13609_not n13803 ; n13804
g13549 and n13617_not n13804_not ; n13805
g13550 and n13802_not n13805 ; n13806
g13551 and n13617_not n13806_not ; n13807
g13552 and b[15] n13606_not ; n13808
g13553 and n13600_not n13808 ; n13809
g13554 and n13608_not n13809_not ; n13810
g13555 and n13807_not n13810 ; n13811
g13556 and n13608_not n13811_not ; n13812
g13557 and b[16] n13597_not ; n13813
g13558 and n13591_not n13813 ; n13814
g13559 and n13599_not n13814_not ; n13815
g13560 and n13812_not n13815 ; n13816
g13561 and n13599_not n13816_not ; n13817
g13562 and b[17] n13588_not ; n13818
g13563 and n13582_not n13818 ; n13819
g13564 and n13590_not n13819_not ; n13820
g13565 and n13817_not n13820 ; n13821
g13566 and n13590_not n13821_not ; n13822
g13567 and b[18] n13579_not ; n13823
g13568 and n13573_not n13823 ; n13824
g13569 and n13581_not n13824_not ; n13825
g13570 and n13822_not n13825 ; n13826
g13571 and n13581_not n13826_not ; n13827
g13572 and b[19] n13570_not ; n13828
g13573 and n13564_not n13828 ; n13829
g13574 and n13572_not n13829_not ; n13830
g13575 and n13827_not n13830 ; n13831
g13576 and n13572_not n13831_not ; n13832
g13577 and b[20] n13561_not ; n13833
g13578 and n13555_not n13833 ; n13834
g13579 and n13563_not n13834_not ; n13835
g13580 and n13832_not n13835 ; n13836
g13581 and n13563_not n13836_not ; n13837
g13582 and b[21] n13552_not ; n13838
g13583 and n13546_not n13838 ; n13839
g13584 and n13554_not n13839_not ; n13840
g13585 and n13837_not n13840 ; n13841
g13586 and n13554_not n13841_not ; n13842
g13587 and b[22] n13543_not ; n13843
g13588 and n13537_not n13843 ; n13844
g13589 and n13545_not n13844_not ; n13845
g13590 and n13842_not n13845 ; n13846
g13591 and n13545_not n13846_not ; n13847
g13592 and b[23] n13534_not ; n13848
g13593 and n13528_not n13848 ; n13849
g13594 and n13536_not n13849_not ; n13850
g13595 and n13847_not n13850 ; n13851
g13596 and n13536_not n13851_not ; n13852
g13597 and b[24] n13525_not ; n13853
g13598 and n13519_not n13853 ; n13854
g13599 and n13527_not n13854_not ; n13855
g13600 and n13852_not n13855 ; n13856
g13601 and n13527_not n13856_not ; n13857
g13602 and b[25] n13516_not ; n13858
g13603 and n13510_not n13858 ; n13859
g13604 and n13518_not n13859_not ; n13860
g13605 and n13857_not n13860 ; n13861
g13606 and n13518_not n13861_not ; n13862
g13607 and b[26] n13507_not ; n13863
g13608 and n13501_not n13863 ; n13864
g13609 and n13509_not n13864_not ; n13865
g13610 and n13862_not n13865 ; n13866
g13611 and n13509_not n13866_not ; n13867
g13612 and b[27] n13498_not ; n13868
g13613 and n13492_not n13868 ; n13869
g13614 and n13500_not n13869_not ; n13870
g13615 and n13867_not n13870 ; n13871
g13616 and n13500_not n13871_not ; n13872
g13617 and b[28] n13489_not ; n13873
g13618 and n13483_not n13873 ; n13874
g13619 and n13491_not n13874_not ; n13875
g13620 and n13872_not n13875 ; n13876
g13621 and n13491_not n13876_not ; n13877
g13622 and b[29] n13480_not ; n13878
g13623 and n13474_not n13878 ; n13879
g13624 and n13482_not n13879_not ; n13880
g13625 and n13877_not n13880 ; n13881
g13626 and n13482_not n13881_not ; n13882
g13627 and b[30] n13471_not ; n13883
g13628 and n13465_not n13883 ; n13884
g13629 and n13473_not n13884_not ; n13885
g13630 and n13882_not n13885 ; n13886
g13631 and n13473_not n13886_not ; n13887
g13632 and b[31] n13462_not ; n13888
g13633 and n13456_not n13888 ; n13889
g13634 and n13464_not n13889_not ; n13890
g13635 and n13887_not n13890 ; n13891
g13636 and n13464_not n13891_not ; n13892
g13637 and b[32] n13453_not ; n13893
g13638 and n13447_not n13893 ; n13894
g13639 and n13455_not n13894_not ; n13895
g13640 and n13892_not n13895 ; n13896
g13641 and n13455_not n13896_not ; n13897
g13642 and b[33] n13444_not ; n13898
g13643 and n13438_not n13898 ; n13899
g13644 and n13446_not n13899_not ; n13900
g13645 and n13897_not n13900 ; n13901
g13646 and n13446_not n13901_not ; n13902
g13647 and b[34] n13435_not ; n13903
g13648 and n13429_not n13903 ; n13904
g13649 and n13437_not n13904_not ; n13905
g13650 and n13902_not n13905 ; n13906
g13651 and n13437_not n13906_not ; n13907
g13652 and b[35] n13426_not ; n13908
g13653 and n13420_not n13908 ; n13909
g13654 and n13428_not n13909_not ; n13910
g13655 and n13907_not n13910 ; n13911
g13656 and n13428_not n13911_not ; n13912
g13657 and b[36] n13417_not ; n13913
g13658 and n13411_not n13913 ; n13914
g13659 and n13419_not n13914_not ; n13915
g13660 and n13912_not n13915 ; n13916
g13661 and n13419_not n13916_not ; n13917
g13662 and b[37] n13408_not ; n13918
g13663 and n13402_not n13918 ; n13919
g13664 and n13410_not n13919_not ; n13920
g13665 and n13917_not n13920 ; n13921
g13666 and n13410_not n13921_not ; n13922
g13667 and b[38] n13399_not ; n13923
g13668 and n13393_not n13923 ; n13924
g13669 and n13401_not n13924_not ; n13925
g13670 and n13922_not n13925 ; n13926
g13671 and n13401_not n13926_not ; n13927
g13672 and b[39] n13390_not ; n13928
g13673 and n13384_not n13928 ; n13929
g13674 and n13392_not n13929_not ; n13930
g13675 and n13927_not n13930 ; n13931
g13676 and n13392_not n13931_not ; n13932
g13677 and b[40] n13381_not ; n13933
g13678 and n13375_not n13933 ; n13934
g13679 and n13383_not n13934_not ; n13935
g13680 and n13932_not n13935 ; n13936
g13681 and n13383_not n13936_not ; n13937
g13682 and b[41] n13372_not ; n13938
g13683 and n13366_not n13938 ; n13939
g13684 and n13374_not n13939_not ; n13940
g13685 and n13937_not n13940 ; n13941
g13686 and n13374_not n13941_not ; n13942
g13687 and b[42] n13363_not ; n13943
g13688 and n13357_not n13943 ; n13944
g13689 and n13365_not n13944_not ; n13945
g13690 and n13942_not n13945 ; n13946
g13691 and n13365_not n13946_not ; n13947
g13692 and n12784_not quotient[21]_not ; n13948
g13693 and n12786_not n13351 ; n13949
g13694 and n13347_not n13949 ; n13950
g13695 and n13348_not n13351_not ; n13951
g13696 and n13950_not n13951_not ; n13952
g13697 and quotient[21] n13952_not ; n13953
g13698 and n13948_not n13953_not ; n13954
g13699 and b[43]_not n13954_not ; n13955
g13700 and b[43] n13948_not ; n13956
g13701 and n13953_not n13956 ; n13957
g13702 and n288 n302 ; n13958
g13703 and n13957_not n13958 ; n13959
g13704 and n13955_not n13959 ; n13960
g13705 and n13947_not n13960 ; n13961
g13706 and n13355 n13954_not ; n13962
g13707 and n13961_not n13962_not ; quotient[20]
g13708 and n13374_not n13945 ; n13964
g13709 and n13941_not n13964 ; n13965
g13710 and n13942_not n13945_not ; n13966
g13711 and n13965_not n13966_not ; n13967
g13712 and quotient[20] n13967_not ; n13968
g13713 and n13364_not n13962_not ; n13969
g13714 and n13961_not n13969 ; n13970
g13715 and n13968_not n13970_not ; n13971
g13716 and b[43]_not n13971_not ; n13972
g13717 and n13383_not n13940 ; n13973
g13718 and n13936_not n13973 ; n13974
g13719 and n13937_not n13940_not ; n13975
g13720 and n13974_not n13975_not ; n13976
g13721 and quotient[20] n13976_not ; n13977
g13722 and n13373_not n13962_not ; n13978
g13723 and n13961_not n13978 ; n13979
g13724 and n13977_not n13979_not ; n13980
g13725 and b[42]_not n13980_not ; n13981
g13726 and n13392_not n13935 ; n13982
g13727 and n13931_not n13982 ; n13983
g13728 and n13932_not n13935_not ; n13984
g13729 and n13983_not n13984_not ; n13985
g13730 and quotient[20] n13985_not ; n13986
g13731 and n13382_not n13962_not ; n13987
g13732 and n13961_not n13987 ; n13988
g13733 and n13986_not n13988_not ; n13989
g13734 and b[41]_not n13989_not ; n13990
g13735 and n13401_not n13930 ; n13991
g13736 and n13926_not n13991 ; n13992
g13737 and n13927_not n13930_not ; n13993
g13738 and n13992_not n13993_not ; n13994
g13739 and quotient[20] n13994_not ; n13995
g13740 and n13391_not n13962_not ; n13996
g13741 and n13961_not n13996 ; n13997
g13742 and n13995_not n13997_not ; n13998
g13743 and b[40]_not n13998_not ; n13999
g13744 and n13410_not n13925 ; n14000
g13745 and n13921_not n14000 ; n14001
g13746 and n13922_not n13925_not ; n14002
g13747 and n14001_not n14002_not ; n14003
g13748 and quotient[20] n14003_not ; n14004
g13749 and n13400_not n13962_not ; n14005
g13750 and n13961_not n14005 ; n14006
g13751 and n14004_not n14006_not ; n14007
g13752 and b[39]_not n14007_not ; n14008
g13753 and n13419_not n13920 ; n14009
g13754 and n13916_not n14009 ; n14010
g13755 and n13917_not n13920_not ; n14011
g13756 and n14010_not n14011_not ; n14012
g13757 and quotient[20] n14012_not ; n14013
g13758 and n13409_not n13962_not ; n14014
g13759 and n13961_not n14014 ; n14015
g13760 and n14013_not n14015_not ; n14016
g13761 and b[38]_not n14016_not ; n14017
g13762 and n13428_not n13915 ; n14018
g13763 and n13911_not n14018 ; n14019
g13764 and n13912_not n13915_not ; n14020
g13765 and n14019_not n14020_not ; n14021
g13766 and quotient[20] n14021_not ; n14022
g13767 and n13418_not n13962_not ; n14023
g13768 and n13961_not n14023 ; n14024
g13769 and n14022_not n14024_not ; n14025
g13770 and b[37]_not n14025_not ; n14026
g13771 and n13437_not n13910 ; n14027
g13772 and n13906_not n14027 ; n14028
g13773 and n13907_not n13910_not ; n14029
g13774 and n14028_not n14029_not ; n14030
g13775 and quotient[20] n14030_not ; n14031
g13776 and n13427_not n13962_not ; n14032
g13777 and n13961_not n14032 ; n14033
g13778 and n14031_not n14033_not ; n14034
g13779 and b[36]_not n14034_not ; n14035
g13780 and n13446_not n13905 ; n14036
g13781 and n13901_not n14036 ; n14037
g13782 and n13902_not n13905_not ; n14038
g13783 and n14037_not n14038_not ; n14039
g13784 and quotient[20] n14039_not ; n14040
g13785 and n13436_not n13962_not ; n14041
g13786 and n13961_not n14041 ; n14042
g13787 and n14040_not n14042_not ; n14043
g13788 and b[35]_not n14043_not ; n14044
g13789 and n13455_not n13900 ; n14045
g13790 and n13896_not n14045 ; n14046
g13791 and n13897_not n13900_not ; n14047
g13792 and n14046_not n14047_not ; n14048
g13793 and quotient[20] n14048_not ; n14049
g13794 and n13445_not n13962_not ; n14050
g13795 and n13961_not n14050 ; n14051
g13796 and n14049_not n14051_not ; n14052
g13797 and b[34]_not n14052_not ; n14053
g13798 and n13464_not n13895 ; n14054
g13799 and n13891_not n14054 ; n14055
g13800 and n13892_not n13895_not ; n14056
g13801 and n14055_not n14056_not ; n14057
g13802 and quotient[20] n14057_not ; n14058
g13803 and n13454_not n13962_not ; n14059
g13804 and n13961_not n14059 ; n14060
g13805 and n14058_not n14060_not ; n14061
g13806 and b[33]_not n14061_not ; n14062
g13807 and n13473_not n13890 ; n14063
g13808 and n13886_not n14063 ; n14064
g13809 and n13887_not n13890_not ; n14065
g13810 and n14064_not n14065_not ; n14066
g13811 and quotient[20] n14066_not ; n14067
g13812 and n13463_not n13962_not ; n14068
g13813 and n13961_not n14068 ; n14069
g13814 and n14067_not n14069_not ; n14070
g13815 and b[32]_not n14070_not ; n14071
g13816 and n13482_not n13885 ; n14072
g13817 and n13881_not n14072 ; n14073
g13818 and n13882_not n13885_not ; n14074
g13819 and n14073_not n14074_not ; n14075
g13820 and quotient[20] n14075_not ; n14076
g13821 and n13472_not n13962_not ; n14077
g13822 and n13961_not n14077 ; n14078
g13823 and n14076_not n14078_not ; n14079
g13824 and b[31]_not n14079_not ; n14080
g13825 and n13491_not n13880 ; n14081
g13826 and n13876_not n14081 ; n14082
g13827 and n13877_not n13880_not ; n14083
g13828 and n14082_not n14083_not ; n14084
g13829 and quotient[20] n14084_not ; n14085
g13830 and n13481_not n13962_not ; n14086
g13831 and n13961_not n14086 ; n14087
g13832 and n14085_not n14087_not ; n14088
g13833 and b[30]_not n14088_not ; n14089
g13834 and n13500_not n13875 ; n14090
g13835 and n13871_not n14090 ; n14091
g13836 and n13872_not n13875_not ; n14092
g13837 and n14091_not n14092_not ; n14093
g13838 and quotient[20] n14093_not ; n14094
g13839 and n13490_not n13962_not ; n14095
g13840 and n13961_not n14095 ; n14096
g13841 and n14094_not n14096_not ; n14097
g13842 and b[29]_not n14097_not ; n14098
g13843 and n13509_not n13870 ; n14099
g13844 and n13866_not n14099 ; n14100
g13845 and n13867_not n13870_not ; n14101
g13846 and n14100_not n14101_not ; n14102
g13847 and quotient[20] n14102_not ; n14103
g13848 and n13499_not n13962_not ; n14104
g13849 and n13961_not n14104 ; n14105
g13850 and n14103_not n14105_not ; n14106
g13851 and b[28]_not n14106_not ; n14107
g13852 and n13518_not n13865 ; n14108
g13853 and n13861_not n14108 ; n14109
g13854 and n13862_not n13865_not ; n14110
g13855 and n14109_not n14110_not ; n14111
g13856 and quotient[20] n14111_not ; n14112
g13857 and n13508_not n13962_not ; n14113
g13858 and n13961_not n14113 ; n14114
g13859 and n14112_not n14114_not ; n14115
g13860 and b[27]_not n14115_not ; n14116
g13861 and n13527_not n13860 ; n14117
g13862 and n13856_not n14117 ; n14118
g13863 and n13857_not n13860_not ; n14119
g13864 and n14118_not n14119_not ; n14120
g13865 and quotient[20] n14120_not ; n14121
g13866 and n13517_not n13962_not ; n14122
g13867 and n13961_not n14122 ; n14123
g13868 and n14121_not n14123_not ; n14124
g13869 and b[26]_not n14124_not ; n14125
g13870 and n13536_not n13855 ; n14126
g13871 and n13851_not n14126 ; n14127
g13872 and n13852_not n13855_not ; n14128
g13873 and n14127_not n14128_not ; n14129
g13874 and quotient[20] n14129_not ; n14130
g13875 and n13526_not n13962_not ; n14131
g13876 and n13961_not n14131 ; n14132
g13877 and n14130_not n14132_not ; n14133
g13878 and b[25]_not n14133_not ; n14134
g13879 and n13545_not n13850 ; n14135
g13880 and n13846_not n14135 ; n14136
g13881 and n13847_not n13850_not ; n14137
g13882 and n14136_not n14137_not ; n14138
g13883 and quotient[20] n14138_not ; n14139
g13884 and n13535_not n13962_not ; n14140
g13885 and n13961_not n14140 ; n14141
g13886 and n14139_not n14141_not ; n14142
g13887 and b[24]_not n14142_not ; n14143
g13888 and n13554_not n13845 ; n14144
g13889 and n13841_not n14144 ; n14145
g13890 and n13842_not n13845_not ; n14146
g13891 and n14145_not n14146_not ; n14147
g13892 and quotient[20] n14147_not ; n14148
g13893 and n13544_not n13962_not ; n14149
g13894 and n13961_not n14149 ; n14150
g13895 and n14148_not n14150_not ; n14151
g13896 and b[23]_not n14151_not ; n14152
g13897 and n13563_not n13840 ; n14153
g13898 and n13836_not n14153 ; n14154
g13899 and n13837_not n13840_not ; n14155
g13900 and n14154_not n14155_not ; n14156
g13901 and quotient[20] n14156_not ; n14157
g13902 and n13553_not n13962_not ; n14158
g13903 and n13961_not n14158 ; n14159
g13904 and n14157_not n14159_not ; n14160
g13905 and b[22]_not n14160_not ; n14161
g13906 and n13572_not n13835 ; n14162
g13907 and n13831_not n14162 ; n14163
g13908 and n13832_not n13835_not ; n14164
g13909 and n14163_not n14164_not ; n14165
g13910 and quotient[20] n14165_not ; n14166
g13911 and n13562_not n13962_not ; n14167
g13912 and n13961_not n14167 ; n14168
g13913 and n14166_not n14168_not ; n14169
g13914 and b[21]_not n14169_not ; n14170
g13915 and n13581_not n13830 ; n14171
g13916 and n13826_not n14171 ; n14172
g13917 and n13827_not n13830_not ; n14173
g13918 and n14172_not n14173_not ; n14174
g13919 and quotient[20] n14174_not ; n14175
g13920 and n13571_not n13962_not ; n14176
g13921 and n13961_not n14176 ; n14177
g13922 and n14175_not n14177_not ; n14178
g13923 and b[20]_not n14178_not ; n14179
g13924 and n13590_not n13825 ; n14180
g13925 and n13821_not n14180 ; n14181
g13926 and n13822_not n13825_not ; n14182
g13927 and n14181_not n14182_not ; n14183
g13928 and quotient[20] n14183_not ; n14184
g13929 and n13580_not n13962_not ; n14185
g13930 and n13961_not n14185 ; n14186
g13931 and n14184_not n14186_not ; n14187
g13932 and b[19]_not n14187_not ; n14188
g13933 and n13599_not n13820 ; n14189
g13934 and n13816_not n14189 ; n14190
g13935 and n13817_not n13820_not ; n14191
g13936 and n14190_not n14191_not ; n14192
g13937 and quotient[20] n14192_not ; n14193
g13938 and n13589_not n13962_not ; n14194
g13939 and n13961_not n14194 ; n14195
g13940 and n14193_not n14195_not ; n14196
g13941 and b[18]_not n14196_not ; n14197
g13942 and n13608_not n13815 ; n14198
g13943 and n13811_not n14198 ; n14199
g13944 and n13812_not n13815_not ; n14200
g13945 and n14199_not n14200_not ; n14201
g13946 and quotient[20] n14201_not ; n14202
g13947 and n13598_not n13962_not ; n14203
g13948 and n13961_not n14203 ; n14204
g13949 and n14202_not n14204_not ; n14205
g13950 and b[17]_not n14205_not ; n14206
g13951 and n13617_not n13810 ; n14207
g13952 and n13806_not n14207 ; n14208
g13953 and n13807_not n13810_not ; n14209
g13954 and n14208_not n14209_not ; n14210
g13955 and quotient[20] n14210_not ; n14211
g13956 and n13607_not n13962_not ; n14212
g13957 and n13961_not n14212 ; n14213
g13958 and n14211_not n14213_not ; n14214
g13959 and b[16]_not n14214_not ; n14215
g13960 and n13626_not n13805 ; n14216
g13961 and n13801_not n14216 ; n14217
g13962 and n13802_not n13805_not ; n14218
g13963 and n14217_not n14218_not ; n14219
g13964 and quotient[20] n14219_not ; n14220
g13965 and n13616_not n13962_not ; n14221
g13966 and n13961_not n14221 ; n14222
g13967 and n14220_not n14222_not ; n14223
g13968 and b[15]_not n14223_not ; n14224
g13969 and n13635_not n13800 ; n14225
g13970 and n13796_not n14225 ; n14226
g13971 and n13797_not n13800_not ; n14227
g13972 and n14226_not n14227_not ; n14228
g13973 and quotient[20] n14228_not ; n14229
g13974 and n13625_not n13962_not ; n14230
g13975 and n13961_not n14230 ; n14231
g13976 and n14229_not n14231_not ; n14232
g13977 and b[14]_not n14232_not ; n14233
g13978 and n13644_not n13795 ; n14234
g13979 and n13791_not n14234 ; n14235
g13980 and n13792_not n13795_not ; n14236
g13981 and n14235_not n14236_not ; n14237
g13982 and quotient[20] n14237_not ; n14238
g13983 and n13634_not n13962_not ; n14239
g13984 and n13961_not n14239 ; n14240
g13985 and n14238_not n14240_not ; n14241
g13986 and b[13]_not n14241_not ; n14242
g13987 and n13653_not n13790 ; n14243
g13988 and n13786_not n14243 ; n14244
g13989 and n13787_not n13790_not ; n14245
g13990 and n14244_not n14245_not ; n14246
g13991 and quotient[20] n14246_not ; n14247
g13992 and n13643_not n13962_not ; n14248
g13993 and n13961_not n14248 ; n14249
g13994 and n14247_not n14249_not ; n14250
g13995 and b[12]_not n14250_not ; n14251
g13996 and n13662_not n13785 ; n14252
g13997 and n13781_not n14252 ; n14253
g13998 and n13782_not n13785_not ; n14254
g13999 and n14253_not n14254_not ; n14255
g14000 and quotient[20] n14255_not ; n14256
g14001 and n13652_not n13962_not ; n14257
g14002 and n13961_not n14257 ; n14258
g14003 and n14256_not n14258_not ; n14259
g14004 and b[11]_not n14259_not ; n14260
g14005 and n13671_not n13780 ; n14261
g14006 and n13776_not n14261 ; n14262
g14007 and n13777_not n13780_not ; n14263
g14008 and n14262_not n14263_not ; n14264
g14009 and quotient[20] n14264_not ; n14265
g14010 and n13661_not n13962_not ; n14266
g14011 and n13961_not n14266 ; n14267
g14012 and n14265_not n14267_not ; n14268
g14013 and b[10]_not n14268_not ; n14269
g14014 and n13680_not n13775 ; n14270
g14015 and n13771_not n14270 ; n14271
g14016 and n13772_not n13775_not ; n14272
g14017 and n14271_not n14272_not ; n14273
g14018 and quotient[20] n14273_not ; n14274
g14019 and n13670_not n13962_not ; n14275
g14020 and n13961_not n14275 ; n14276
g14021 and n14274_not n14276_not ; n14277
g14022 and b[9]_not n14277_not ; n14278
g14023 and n13689_not n13770 ; n14279
g14024 and n13766_not n14279 ; n14280
g14025 and n13767_not n13770_not ; n14281
g14026 and n14280_not n14281_not ; n14282
g14027 and quotient[20] n14282_not ; n14283
g14028 and n13679_not n13962_not ; n14284
g14029 and n13961_not n14284 ; n14285
g14030 and n14283_not n14285_not ; n14286
g14031 and b[8]_not n14286_not ; n14287
g14032 and n13698_not n13765 ; n14288
g14033 and n13761_not n14288 ; n14289
g14034 and n13762_not n13765_not ; n14290
g14035 and n14289_not n14290_not ; n14291
g14036 and quotient[20] n14291_not ; n14292
g14037 and n13688_not n13962_not ; n14293
g14038 and n13961_not n14293 ; n14294
g14039 and n14292_not n14294_not ; n14295
g14040 and b[7]_not n14295_not ; n14296
g14041 and n13707_not n13760 ; n14297
g14042 and n13756_not n14297 ; n14298
g14043 and n13757_not n13760_not ; n14299
g14044 and n14298_not n14299_not ; n14300
g14045 and quotient[20] n14300_not ; n14301
g14046 and n13697_not n13962_not ; n14302
g14047 and n13961_not n14302 ; n14303
g14048 and n14301_not n14303_not ; n14304
g14049 and b[6]_not n14304_not ; n14305
g14050 and n13716_not n13755 ; n14306
g14051 and n13751_not n14306 ; n14307
g14052 and n13752_not n13755_not ; n14308
g14053 and n14307_not n14308_not ; n14309
g14054 and quotient[20] n14309_not ; n14310
g14055 and n13706_not n13962_not ; n14311
g14056 and n13961_not n14311 ; n14312
g14057 and n14310_not n14312_not ; n14313
g14058 and b[5]_not n14313_not ; n14314
g14059 and n13724_not n13750 ; n14315
g14060 and n13746_not n14315 ; n14316
g14061 and n13747_not n13750_not ; n14317
g14062 and n14316_not n14317_not ; n14318
g14063 and quotient[20] n14318_not ; n14319
g14064 and n13715_not n13962_not ; n14320
g14065 and n13961_not n14320 ; n14321
g14066 and n14319_not n14321_not ; n14322
g14067 and b[4]_not n14322_not ; n14323
g14068 and n13741_not n13745 ; n14324
g14069 and n13740_not n14324 ; n14325
g14070 and n13742_not n13745_not ; n14326
g14071 and n14325_not n14326_not ; n14327
g14072 and quotient[20] n14327_not ; n14328
g14073 and n13723_not n13962_not ; n14329
g14074 and n13961_not n14329 ; n14330
g14075 and n14328_not n14330_not ; n14331
g14076 and b[3]_not n14331_not ; n14332
g14077 and n13737_not n13739 ; n14333
g14078 and n13735_not n14333 ; n14334
g14079 and n13740_not n14334_not ; n14335
g14080 and quotient[20] n14335 ; n14336
g14081 and n13734_not n13962_not ; n14337
g14082 and n13961_not n14337 ; n14338
g14083 and n14336_not n14338_not ; n14339
g14084 and b[2]_not n14339_not ; n14340
g14085 and b[0] quotient[20] ; n14341
g14086 and a[20] n14341_not ; n14342
g14087 and n13739 quotient[20] ; n14343
g14088 and n14342_not n14343_not ; n14344
g14089 and b[1] n14344_not ; n14345
g14090 and b[1]_not n14343_not ; n14346
g14091 and n14342_not n14346 ; n14347
g14092 and n14345_not n14347_not ; n14348
g14093 and a[19]_not b[0] ; n14349
g14094 and n14348_not n14349_not ; n14350
g14095 and b[1]_not n14344_not ; n14351
g14096 and n14350_not n14351_not ; n14352
g14097 and b[2] n14338_not ; n14353
g14098 and n14336_not n14353 ; n14354
g14099 and n14340_not n14354_not ; n14355
g14100 and n14352_not n14355 ; n14356
g14101 and n14340_not n14356_not ; n14357
g14102 and b[3] n14330_not ; n14358
g14103 and n14328_not n14358 ; n14359
g14104 and n14332_not n14359_not ; n14360
g14105 and n14357_not n14360 ; n14361
g14106 and n14332_not n14361_not ; n14362
g14107 and b[4] n14321_not ; n14363
g14108 and n14319_not n14363 ; n14364
g14109 and n14323_not n14364_not ; n14365
g14110 and n14362_not n14365 ; n14366
g14111 and n14323_not n14366_not ; n14367
g14112 and b[5] n14312_not ; n14368
g14113 and n14310_not n14368 ; n14369
g14114 and n14314_not n14369_not ; n14370
g14115 and n14367_not n14370 ; n14371
g14116 and n14314_not n14371_not ; n14372
g14117 and b[6] n14303_not ; n14373
g14118 and n14301_not n14373 ; n14374
g14119 and n14305_not n14374_not ; n14375
g14120 and n14372_not n14375 ; n14376
g14121 and n14305_not n14376_not ; n14377
g14122 and b[7] n14294_not ; n14378
g14123 and n14292_not n14378 ; n14379
g14124 and n14296_not n14379_not ; n14380
g14125 and n14377_not n14380 ; n14381
g14126 and n14296_not n14381_not ; n14382
g14127 and b[8] n14285_not ; n14383
g14128 and n14283_not n14383 ; n14384
g14129 and n14287_not n14384_not ; n14385
g14130 and n14382_not n14385 ; n14386
g14131 and n14287_not n14386_not ; n14387
g14132 and b[9] n14276_not ; n14388
g14133 and n14274_not n14388 ; n14389
g14134 and n14278_not n14389_not ; n14390
g14135 and n14387_not n14390 ; n14391
g14136 and n14278_not n14391_not ; n14392
g14137 and b[10] n14267_not ; n14393
g14138 and n14265_not n14393 ; n14394
g14139 and n14269_not n14394_not ; n14395
g14140 and n14392_not n14395 ; n14396
g14141 and n14269_not n14396_not ; n14397
g14142 and b[11] n14258_not ; n14398
g14143 and n14256_not n14398 ; n14399
g14144 and n14260_not n14399_not ; n14400
g14145 and n14397_not n14400 ; n14401
g14146 and n14260_not n14401_not ; n14402
g14147 and b[12] n14249_not ; n14403
g14148 and n14247_not n14403 ; n14404
g14149 and n14251_not n14404_not ; n14405
g14150 and n14402_not n14405 ; n14406
g14151 and n14251_not n14406_not ; n14407
g14152 and b[13] n14240_not ; n14408
g14153 and n14238_not n14408 ; n14409
g14154 and n14242_not n14409_not ; n14410
g14155 and n14407_not n14410 ; n14411
g14156 and n14242_not n14411_not ; n14412
g14157 and b[14] n14231_not ; n14413
g14158 and n14229_not n14413 ; n14414
g14159 and n14233_not n14414_not ; n14415
g14160 and n14412_not n14415 ; n14416
g14161 and n14233_not n14416_not ; n14417
g14162 and b[15] n14222_not ; n14418
g14163 and n14220_not n14418 ; n14419
g14164 and n14224_not n14419_not ; n14420
g14165 and n14417_not n14420 ; n14421
g14166 and n14224_not n14421_not ; n14422
g14167 and b[16] n14213_not ; n14423
g14168 and n14211_not n14423 ; n14424
g14169 and n14215_not n14424_not ; n14425
g14170 and n14422_not n14425 ; n14426
g14171 and n14215_not n14426_not ; n14427
g14172 and b[17] n14204_not ; n14428
g14173 and n14202_not n14428 ; n14429
g14174 and n14206_not n14429_not ; n14430
g14175 and n14427_not n14430 ; n14431
g14176 and n14206_not n14431_not ; n14432
g14177 and b[18] n14195_not ; n14433
g14178 and n14193_not n14433 ; n14434
g14179 and n14197_not n14434_not ; n14435
g14180 and n14432_not n14435 ; n14436
g14181 and n14197_not n14436_not ; n14437
g14182 and b[19] n14186_not ; n14438
g14183 and n14184_not n14438 ; n14439
g14184 and n14188_not n14439_not ; n14440
g14185 and n14437_not n14440 ; n14441
g14186 and n14188_not n14441_not ; n14442
g14187 and b[20] n14177_not ; n14443
g14188 and n14175_not n14443 ; n14444
g14189 and n14179_not n14444_not ; n14445
g14190 and n14442_not n14445 ; n14446
g14191 and n14179_not n14446_not ; n14447
g14192 and b[21] n14168_not ; n14448
g14193 and n14166_not n14448 ; n14449
g14194 and n14170_not n14449_not ; n14450
g14195 and n14447_not n14450 ; n14451
g14196 and n14170_not n14451_not ; n14452
g14197 and b[22] n14159_not ; n14453
g14198 and n14157_not n14453 ; n14454
g14199 and n14161_not n14454_not ; n14455
g14200 and n14452_not n14455 ; n14456
g14201 and n14161_not n14456_not ; n14457
g14202 and b[23] n14150_not ; n14458
g14203 and n14148_not n14458 ; n14459
g14204 and n14152_not n14459_not ; n14460
g14205 and n14457_not n14460 ; n14461
g14206 and n14152_not n14461_not ; n14462
g14207 and b[24] n14141_not ; n14463
g14208 and n14139_not n14463 ; n14464
g14209 and n14143_not n14464_not ; n14465
g14210 and n14462_not n14465 ; n14466
g14211 and n14143_not n14466_not ; n14467
g14212 and b[25] n14132_not ; n14468
g14213 and n14130_not n14468 ; n14469
g14214 and n14134_not n14469_not ; n14470
g14215 and n14467_not n14470 ; n14471
g14216 and n14134_not n14471_not ; n14472
g14217 and b[26] n14123_not ; n14473
g14218 and n14121_not n14473 ; n14474
g14219 and n14125_not n14474_not ; n14475
g14220 and n14472_not n14475 ; n14476
g14221 and n14125_not n14476_not ; n14477
g14222 and b[27] n14114_not ; n14478
g14223 and n14112_not n14478 ; n14479
g14224 and n14116_not n14479_not ; n14480
g14225 and n14477_not n14480 ; n14481
g14226 and n14116_not n14481_not ; n14482
g14227 and b[28] n14105_not ; n14483
g14228 and n14103_not n14483 ; n14484
g14229 and n14107_not n14484_not ; n14485
g14230 and n14482_not n14485 ; n14486
g14231 and n14107_not n14486_not ; n14487
g14232 and b[29] n14096_not ; n14488
g14233 and n14094_not n14488 ; n14489
g14234 and n14098_not n14489_not ; n14490
g14235 and n14487_not n14490 ; n14491
g14236 and n14098_not n14491_not ; n14492
g14237 and b[30] n14087_not ; n14493
g14238 and n14085_not n14493 ; n14494
g14239 and n14089_not n14494_not ; n14495
g14240 and n14492_not n14495 ; n14496
g14241 and n14089_not n14496_not ; n14497
g14242 and b[31] n14078_not ; n14498
g14243 and n14076_not n14498 ; n14499
g14244 and n14080_not n14499_not ; n14500
g14245 and n14497_not n14500 ; n14501
g14246 and n14080_not n14501_not ; n14502
g14247 and b[32] n14069_not ; n14503
g14248 and n14067_not n14503 ; n14504
g14249 and n14071_not n14504_not ; n14505
g14250 and n14502_not n14505 ; n14506
g14251 and n14071_not n14506_not ; n14507
g14252 and b[33] n14060_not ; n14508
g14253 and n14058_not n14508 ; n14509
g14254 and n14062_not n14509_not ; n14510
g14255 and n14507_not n14510 ; n14511
g14256 and n14062_not n14511_not ; n14512
g14257 and b[34] n14051_not ; n14513
g14258 and n14049_not n14513 ; n14514
g14259 and n14053_not n14514_not ; n14515
g14260 and n14512_not n14515 ; n14516
g14261 and n14053_not n14516_not ; n14517
g14262 and b[35] n14042_not ; n14518
g14263 and n14040_not n14518 ; n14519
g14264 and n14044_not n14519_not ; n14520
g14265 and n14517_not n14520 ; n14521
g14266 and n14044_not n14521_not ; n14522
g14267 and b[36] n14033_not ; n14523
g14268 and n14031_not n14523 ; n14524
g14269 and n14035_not n14524_not ; n14525
g14270 and n14522_not n14525 ; n14526
g14271 and n14035_not n14526_not ; n14527
g14272 and b[37] n14024_not ; n14528
g14273 and n14022_not n14528 ; n14529
g14274 and n14026_not n14529_not ; n14530
g14275 and n14527_not n14530 ; n14531
g14276 and n14026_not n14531_not ; n14532
g14277 and b[38] n14015_not ; n14533
g14278 and n14013_not n14533 ; n14534
g14279 and n14017_not n14534_not ; n14535
g14280 and n14532_not n14535 ; n14536
g14281 and n14017_not n14536_not ; n14537
g14282 and b[39] n14006_not ; n14538
g14283 and n14004_not n14538 ; n14539
g14284 and n14008_not n14539_not ; n14540
g14285 and n14537_not n14540 ; n14541
g14286 and n14008_not n14541_not ; n14542
g14287 and b[40] n13997_not ; n14543
g14288 and n13995_not n14543 ; n14544
g14289 and n13999_not n14544_not ; n14545
g14290 and n14542_not n14545 ; n14546
g14291 and n13999_not n14546_not ; n14547
g14292 and b[41] n13988_not ; n14548
g14293 and n13986_not n14548 ; n14549
g14294 and n13990_not n14549_not ; n14550
g14295 and n14547_not n14550 ; n14551
g14296 and n13990_not n14551_not ; n14552
g14297 and b[42] n13979_not ; n14553
g14298 and n13977_not n14553 ; n14554
g14299 and n13981_not n14554_not ; n14555
g14300 and n14552_not n14555 ; n14556
g14301 and n13981_not n14556_not ; n14557
g14302 and b[43] n13970_not ; n14558
g14303 and n13968_not n14558 ; n14559
g14304 and n13972_not n14559_not ; n14560
g14305 and n14557_not n14560 ; n14561
g14306 and n13972_not n14561_not ; n14562
g14307 and n13365_not n13957_not ; n14563
g14308 and n13955_not n14563 ; n14564
g14309 and n13946_not n14564 ; n14565
g14310 and n13955_not n13957_not ; n14566
g14311 and n13947_not n14566_not ; n14567
g14312 and n14565_not n14567_not ; n14568
g14313 and quotient[20] n14568_not ; n14569
g14314 and n13954_not n13962_not ; n14570
g14315 and n13961_not n14570 ; n14571
g14316 and n14569_not n14571_not ; n14572
g14317 and b[44]_not n14572_not ; n14573
g14318 and b[44] n14571_not ; n14574
g14319 and n14569_not n14574 ; n14575
g14320 and n595 n597 ; n14576
g14321 and n14575_not n14576 ; n14577
g14322 and n14573_not n14577 ; n14578
g14323 and n14562_not n14578 ; n14579
g14324 and n13958 n14572_not ; n14580
g14325 and n14579_not n14580_not ; quotient[19]
g14326 and n13981_not n14560 ; n14582
g14327 and n14556_not n14582 ; n14583
g14328 and n14557_not n14560_not ; n14584
g14329 and n14583_not n14584_not ; n14585
g14330 and quotient[19] n14585_not ; n14586
g14331 and n13971_not n14580_not ; n14587
g14332 and n14579_not n14587 ; n14588
g14333 and n14586_not n14588_not ; n14589
g14334 and n13972_not n14575_not ; n14590
g14335 and n14573_not n14590 ; n14591
g14336 and n14561_not n14591 ; n14592
g14337 and n14573_not n14575_not ; n14593
g14338 and n14562_not n14593_not ; n14594
g14339 and n14592_not n14594_not ; n14595
g14340 and quotient[19] n14595_not ; n14596
g14341 and n14572_not n14580_not ; n14597
g14342 and n14579_not n14597 ; n14598
g14343 and n14596_not n14598_not ; n14599
g14344 and b[45]_not n14599_not ; n14600
g14345 and b[44]_not n14589_not ; n14601
g14346 and n13990_not n14555 ; n14602
g14347 and n14551_not n14602 ; n14603
g14348 and n14552_not n14555_not ; n14604
g14349 and n14603_not n14604_not ; n14605
g14350 and quotient[19] n14605_not ; n14606
g14351 and n13980_not n14580_not ; n14607
g14352 and n14579_not n14607 ; n14608
g14353 and n14606_not n14608_not ; n14609
g14354 and b[43]_not n14609_not ; n14610
g14355 and n13999_not n14550 ; n14611
g14356 and n14546_not n14611 ; n14612
g14357 and n14547_not n14550_not ; n14613
g14358 and n14612_not n14613_not ; n14614
g14359 and quotient[19] n14614_not ; n14615
g14360 and n13989_not n14580_not ; n14616
g14361 and n14579_not n14616 ; n14617
g14362 and n14615_not n14617_not ; n14618
g14363 and b[42]_not n14618_not ; n14619
g14364 and n14008_not n14545 ; n14620
g14365 and n14541_not n14620 ; n14621
g14366 and n14542_not n14545_not ; n14622
g14367 and n14621_not n14622_not ; n14623
g14368 and quotient[19] n14623_not ; n14624
g14369 and n13998_not n14580_not ; n14625
g14370 and n14579_not n14625 ; n14626
g14371 and n14624_not n14626_not ; n14627
g14372 and b[41]_not n14627_not ; n14628
g14373 and n14017_not n14540 ; n14629
g14374 and n14536_not n14629 ; n14630
g14375 and n14537_not n14540_not ; n14631
g14376 and n14630_not n14631_not ; n14632
g14377 and quotient[19] n14632_not ; n14633
g14378 and n14007_not n14580_not ; n14634
g14379 and n14579_not n14634 ; n14635
g14380 and n14633_not n14635_not ; n14636
g14381 and b[40]_not n14636_not ; n14637
g14382 and n14026_not n14535 ; n14638
g14383 and n14531_not n14638 ; n14639
g14384 and n14532_not n14535_not ; n14640
g14385 and n14639_not n14640_not ; n14641
g14386 and quotient[19] n14641_not ; n14642
g14387 and n14016_not n14580_not ; n14643
g14388 and n14579_not n14643 ; n14644
g14389 and n14642_not n14644_not ; n14645
g14390 and b[39]_not n14645_not ; n14646
g14391 and n14035_not n14530 ; n14647
g14392 and n14526_not n14647 ; n14648
g14393 and n14527_not n14530_not ; n14649
g14394 and n14648_not n14649_not ; n14650
g14395 and quotient[19] n14650_not ; n14651
g14396 and n14025_not n14580_not ; n14652
g14397 and n14579_not n14652 ; n14653
g14398 and n14651_not n14653_not ; n14654
g14399 and b[38]_not n14654_not ; n14655
g14400 and n14044_not n14525 ; n14656
g14401 and n14521_not n14656 ; n14657
g14402 and n14522_not n14525_not ; n14658
g14403 and n14657_not n14658_not ; n14659
g14404 and quotient[19] n14659_not ; n14660
g14405 and n14034_not n14580_not ; n14661
g14406 and n14579_not n14661 ; n14662
g14407 and n14660_not n14662_not ; n14663
g14408 and b[37]_not n14663_not ; n14664
g14409 and n14053_not n14520 ; n14665
g14410 and n14516_not n14665 ; n14666
g14411 and n14517_not n14520_not ; n14667
g14412 and n14666_not n14667_not ; n14668
g14413 and quotient[19] n14668_not ; n14669
g14414 and n14043_not n14580_not ; n14670
g14415 and n14579_not n14670 ; n14671
g14416 and n14669_not n14671_not ; n14672
g14417 and b[36]_not n14672_not ; n14673
g14418 and n14062_not n14515 ; n14674
g14419 and n14511_not n14674 ; n14675
g14420 and n14512_not n14515_not ; n14676
g14421 and n14675_not n14676_not ; n14677
g14422 and quotient[19] n14677_not ; n14678
g14423 and n14052_not n14580_not ; n14679
g14424 and n14579_not n14679 ; n14680
g14425 and n14678_not n14680_not ; n14681
g14426 and b[35]_not n14681_not ; n14682
g14427 and n14071_not n14510 ; n14683
g14428 and n14506_not n14683 ; n14684
g14429 and n14507_not n14510_not ; n14685
g14430 and n14684_not n14685_not ; n14686
g14431 and quotient[19] n14686_not ; n14687
g14432 and n14061_not n14580_not ; n14688
g14433 and n14579_not n14688 ; n14689
g14434 and n14687_not n14689_not ; n14690
g14435 and b[34]_not n14690_not ; n14691
g14436 and n14080_not n14505 ; n14692
g14437 and n14501_not n14692 ; n14693
g14438 and n14502_not n14505_not ; n14694
g14439 and n14693_not n14694_not ; n14695
g14440 and quotient[19] n14695_not ; n14696
g14441 and n14070_not n14580_not ; n14697
g14442 and n14579_not n14697 ; n14698
g14443 and n14696_not n14698_not ; n14699
g14444 and b[33]_not n14699_not ; n14700
g14445 and n14089_not n14500 ; n14701
g14446 and n14496_not n14701 ; n14702
g14447 and n14497_not n14500_not ; n14703
g14448 and n14702_not n14703_not ; n14704
g14449 and quotient[19] n14704_not ; n14705
g14450 and n14079_not n14580_not ; n14706
g14451 and n14579_not n14706 ; n14707
g14452 and n14705_not n14707_not ; n14708
g14453 and b[32]_not n14708_not ; n14709
g14454 and n14098_not n14495 ; n14710
g14455 and n14491_not n14710 ; n14711
g14456 and n14492_not n14495_not ; n14712
g14457 and n14711_not n14712_not ; n14713
g14458 and quotient[19] n14713_not ; n14714
g14459 and n14088_not n14580_not ; n14715
g14460 and n14579_not n14715 ; n14716
g14461 and n14714_not n14716_not ; n14717
g14462 and b[31]_not n14717_not ; n14718
g14463 and n14107_not n14490 ; n14719
g14464 and n14486_not n14719 ; n14720
g14465 and n14487_not n14490_not ; n14721
g14466 and n14720_not n14721_not ; n14722
g14467 and quotient[19] n14722_not ; n14723
g14468 and n14097_not n14580_not ; n14724
g14469 and n14579_not n14724 ; n14725
g14470 and n14723_not n14725_not ; n14726
g14471 and b[30]_not n14726_not ; n14727
g14472 and n14116_not n14485 ; n14728
g14473 and n14481_not n14728 ; n14729
g14474 and n14482_not n14485_not ; n14730
g14475 and n14729_not n14730_not ; n14731
g14476 and quotient[19] n14731_not ; n14732
g14477 and n14106_not n14580_not ; n14733
g14478 and n14579_not n14733 ; n14734
g14479 and n14732_not n14734_not ; n14735
g14480 and b[29]_not n14735_not ; n14736
g14481 and n14125_not n14480 ; n14737
g14482 and n14476_not n14737 ; n14738
g14483 and n14477_not n14480_not ; n14739
g14484 and n14738_not n14739_not ; n14740
g14485 and quotient[19] n14740_not ; n14741
g14486 and n14115_not n14580_not ; n14742
g14487 and n14579_not n14742 ; n14743
g14488 and n14741_not n14743_not ; n14744
g14489 and b[28]_not n14744_not ; n14745
g14490 and n14134_not n14475 ; n14746
g14491 and n14471_not n14746 ; n14747
g14492 and n14472_not n14475_not ; n14748
g14493 and n14747_not n14748_not ; n14749
g14494 and quotient[19] n14749_not ; n14750
g14495 and n14124_not n14580_not ; n14751
g14496 and n14579_not n14751 ; n14752
g14497 and n14750_not n14752_not ; n14753
g14498 and b[27]_not n14753_not ; n14754
g14499 and n14143_not n14470 ; n14755
g14500 and n14466_not n14755 ; n14756
g14501 and n14467_not n14470_not ; n14757
g14502 and n14756_not n14757_not ; n14758
g14503 and quotient[19] n14758_not ; n14759
g14504 and n14133_not n14580_not ; n14760
g14505 and n14579_not n14760 ; n14761
g14506 and n14759_not n14761_not ; n14762
g14507 and b[26]_not n14762_not ; n14763
g14508 and n14152_not n14465 ; n14764
g14509 and n14461_not n14764 ; n14765
g14510 and n14462_not n14465_not ; n14766
g14511 and n14765_not n14766_not ; n14767
g14512 and quotient[19] n14767_not ; n14768
g14513 and n14142_not n14580_not ; n14769
g14514 and n14579_not n14769 ; n14770
g14515 and n14768_not n14770_not ; n14771
g14516 and b[25]_not n14771_not ; n14772
g14517 and n14161_not n14460 ; n14773
g14518 and n14456_not n14773 ; n14774
g14519 and n14457_not n14460_not ; n14775
g14520 and n14774_not n14775_not ; n14776
g14521 and quotient[19] n14776_not ; n14777
g14522 and n14151_not n14580_not ; n14778
g14523 and n14579_not n14778 ; n14779
g14524 and n14777_not n14779_not ; n14780
g14525 and b[24]_not n14780_not ; n14781
g14526 and n14170_not n14455 ; n14782
g14527 and n14451_not n14782 ; n14783
g14528 and n14452_not n14455_not ; n14784
g14529 and n14783_not n14784_not ; n14785
g14530 and quotient[19] n14785_not ; n14786
g14531 and n14160_not n14580_not ; n14787
g14532 and n14579_not n14787 ; n14788
g14533 and n14786_not n14788_not ; n14789
g14534 and b[23]_not n14789_not ; n14790
g14535 and n14179_not n14450 ; n14791
g14536 and n14446_not n14791 ; n14792
g14537 and n14447_not n14450_not ; n14793
g14538 and n14792_not n14793_not ; n14794
g14539 and quotient[19] n14794_not ; n14795
g14540 and n14169_not n14580_not ; n14796
g14541 and n14579_not n14796 ; n14797
g14542 and n14795_not n14797_not ; n14798
g14543 and b[22]_not n14798_not ; n14799
g14544 and n14188_not n14445 ; n14800
g14545 and n14441_not n14800 ; n14801
g14546 and n14442_not n14445_not ; n14802
g14547 and n14801_not n14802_not ; n14803
g14548 and quotient[19] n14803_not ; n14804
g14549 and n14178_not n14580_not ; n14805
g14550 and n14579_not n14805 ; n14806
g14551 and n14804_not n14806_not ; n14807
g14552 and b[21]_not n14807_not ; n14808
g14553 and n14197_not n14440 ; n14809
g14554 and n14436_not n14809 ; n14810
g14555 and n14437_not n14440_not ; n14811
g14556 and n14810_not n14811_not ; n14812
g14557 and quotient[19] n14812_not ; n14813
g14558 and n14187_not n14580_not ; n14814
g14559 and n14579_not n14814 ; n14815
g14560 and n14813_not n14815_not ; n14816
g14561 and b[20]_not n14816_not ; n14817
g14562 and n14206_not n14435 ; n14818
g14563 and n14431_not n14818 ; n14819
g14564 and n14432_not n14435_not ; n14820
g14565 and n14819_not n14820_not ; n14821
g14566 and quotient[19] n14821_not ; n14822
g14567 and n14196_not n14580_not ; n14823
g14568 and n14579_not n14823 ; n14824
g14569 and n14822_not n14824_not ; n14825
g14570 and b[19]_not n14825_not ; n14826
g14571 and n14215_not n14430 ; n14827
g14572 and n14426_not n14827 ; n14828
g14573 and n14427_not n14430_not ; n14829
g14574 and n14828_not n14829_not ; n14830
g14575 and quotient[19] n14830_not ; n14831
g14576 and n14205_not n14580_not ; n14832
g14577 and n14579_not n14832 ; n14833
g14578 and n14831_not n14833_not ; n14834
g14579 and b[18]_not n14834_not ; n14835
g14580 and n14224_not n14425 ; n14836
g14581 and n14421_not n14836 ; n14837
g14582 and n14422_not n14425_not ; n14838
g14583 and n14837_not n14838_not ; n14839
g14584 and quotient[19] n14839_not ; n14840
g14585 and n14214_not n14580_not ; n14841
g14586 and n14579_not n14841 ; n14842
g14587 and n14840_not n14842_not ; n14843
g14588 and b[17]_not n14843_not ; n14844
g14589 and n14233_not n14420 ; n14845
g14590 and n14416_not n14845 ; n14846
g14591 and n14417_not n14420_not ; n14847
g14592 and n14846_not n14847_not ; n14848
g14593 and quotient[19] n14848_not ; n14849
g14594 and n14223_not n14580_not ; n14850
g14595 and n14579_not n14850 ; n14851
g14596 and n14849_not n14851_not ; n14852
g14597 and b[16]_not n14852_not ; n14853
g14598 and n14242_not n14415 ; n14854
g14599 and n14411_not n14854 ; n14855
g14600 and n14412_not n14415_not ; n14856
g14601 and n14855_not n14856_not ; n14857
g14602 and quotient[19] n14857_not ; n14858
g14603 and n14232_not n14580_not ; n14859
g14604 and n14579_not n14859 ; n14860
g14605 and n14858_not n14860_not ; n14861
g14606 and b[15]_not n14861_not ; n14862
g14607 and n14251_not n14410 ; n14863
g14608 and n14406_not n14863 ; n14864
g14609 and n14407_not n14410_not ; n14865
g14610 and n14864_not n14865_not ; n14866
g14611 and quotient[19] n14866_not ; n14867
g14612 and n14241_not n14580_not ; n14868
g14613 and n14579_not n14868 ; n14869
g14614 and n14867_not n14869_not ; n14870
g14615 and b[14]_not n14870_not ; n14871
g14616 and n14260_not n14405 ; n14872
g14617 and n14401_not n14872 ; n14873
g14618 and n14402_not n14405_not ; n14874
g14619 and n14873_not n14874_not ; n14875
g14620 and quotient[19] n14875_not ; n14876
g14621 and n14250_not n14580_not ; n14877
g14622 and n14579_not n14877 ; n14878
g14623 and n14876_not n14878_not ; n14879
g14624 and b[13]_not n14879_not ; n14880
g14625 and n14269_not n14400 ; n14881
g14626 and n14396_not n14881 ; n14882
g14627 and n14397_not n14400_not ; n14883
g14628 and n14882_not n14883_not ; n14884
g14629 and quotient[19] n14884_not ; n14885
g14630 and n14259_not n14580_not ; n14886
g14631 and n14579_not n14886 ; n14887
g14632 and n14885_not n14887_not ; n14888
g14633 and b[12]_not n14888_not ; n14889
g14634 and n14278_not n14395 ; n14890
g14635 and n14391_not n14890 ; n14891
g14636 and n14392_not n14395_not ; n14892
g14637 and n14891_not n14892_not ; n14893
g14638 and quotient[19] n14893_not ; n14894
g14639 and n14268_not n14580_not ; n14895
g14640 and n14579_not n14895 ; n14896
g14641 and n14894_not n14896_not ; n14897
g14642 and b[11]_not n14897_not ; n14898
g14643 and n14287_not n14390 ; n14899
g14644 and n14386_not n14899 ; n14900
g14645 and n14387_not n14390_not ; n14901
g14646 and n14900_not n14901_not ; n14902
g14647 and quotient[19] n14902_not ; n14903
g14648 and n14277_not n14580_not ; n14904
g14649 and n14579_not n14904 ; n14905
g14650 and n14903_not n14905_not ; n14906
g14651 and b[10]_not n14906_not ; n14907
g14652 and n14296_not n14385 ; n14908
g14653 and n14381_not n14908 ; n14909
g14654 and n14382_not n14385_not ; n14910
g14655 and n14909_not n14910_not ; n14911
g14656 and quotient[19] n14911_not ; n14912
g14657 and n14286_not n14580_not ; n14913
g14658 and n14579_not n14913 ; n14914
g14659 and n14912_not n14914_not ; n14915
g14660 and b[9]_not n14915_not ; n14916
g14661 and n14305_not n14380 ; n14917
g14662 and n14376_not n14917 ; n14918
g14663 and n14377_not n14380_not ; n14919
g14664 and n14918_not n14919_not ; n14920
g14665 and quotient[19] n14920_not ; n14921
g14666 and n14295_not n14580_not ; n14922
g14667 and n14579_not n14922 ; n14923
g14668 and n14921_not n14923_not ; n14924
g14669 and b[8]_not n14924_not ; n14925
g14670 and n14314_not n14375 ; n14926
g14671 and n14371_not n14926 ; n14927
g14672 and n14372_not n14375_not ; n14928
g14673 and n14927_not n14928_not ; n14929
g14674 and quotient[19] n14929_not ; n14930
g14675 and n14304_not n14580_not ; n14931
g14676 and n14579_not n14931 ; n14932
g14677 and n14930_not n14932_not ; n14933
g14678 and b[7]_not n14933_not ; n14934
g14679 and n14323_not n14370 ; n14935
g14680 and n14366_not n14935 ; n14936
g14681 and n14367_not n14370_not ; n14937
g14682 and n14936_not n14937_not ; n14938
g14683 and quotient[19] n14938_not ; n14939
g14684 and n14313_not n14580_not ; n14940
g14685 and n14579_not n14940 ; n14941
g14686 and n14939_not n14941_not ; n14942
g14687 and b[6]_not n14942_not ; n14943
g14688 and n14332_not n14365 ; n14944
g14689 and n14361_not n14944 ; n14945
g14690 and n14362_not n14365_not ; n14946
g14691 and n14945_not n14946_not ; n14947
g14692 and quotient[19] n14947_not ; n14948
g14693 and n14322_not n14580_not ; n14949
g14694 and n14579_not n14949 ; n14950
g14695 and n14948_not n14950_not ; n14951
g14696 and b[5]_not n14951_not ; n14952
g14697 and n14340_not n14360 ; n14953
g14698 and n14356_not n14953 ; n14954
g14699 and n14357_not n14360_not ; n14955
g14700 and n14954_not n14955_not ; n14956
g14701 and quotient[19] n14956_not ; n14957
g14702 and n14331_not n14580_not ; n14958
g14703 and n14579_not n14958 ; n14959
g14704 and n14957_not n14959_not ; n14960
g14705 and b[4]_not n14960_not ; n14961
g14706 and n14351_not n14355 ; n14962
g14707 and n14350_not n14962 ; n14963
g14708 and n14352_not n14355_not ; n14964
g14709 and n14963_not n14964_not ; n14965
g14710 and quotient[19] n14965_not ; n14966
g14711 and n14339_not n14580_not ; n14967
g14712 and n14579_not n14967 ; n14968
g14713 and n14966_not n14968_not ; n14969
g14714 and b[3]_not n14969_not ; n14970
g14715 and n14347_not n14349 ; n14971
g14716 and n14345_not n14971 ; n14972
g14717 and n14350_not n14972_not ; n14973
g14718 and quotient[19] n14973 ; n14974
g14719 and n14344_not n14580_not ; n14975
g14720 and n14579_not n14975 ; n14976
g14721 and n14974_not n14976_not ; n14977
g14722 and b[2]_not n14977_not ; n14978
g14723 and b[0] quotient[19] ; n14979
g14724 and a[19] n14979_not ; n14980
g14725 and n14349 quotient[19] ; n14981
g14726 and n14980_not n14981_not ; n14982
g14727 and b[1] n14982_not ; n14983
g14728 and b[1]_not n14981_not ; n14984
g14729 and n14980_not n14984 ; n14985
g14730 and n14983_not n14985_not ; n14986
g14731 and a[18]_not b[0] ; n14987
g14732 and n14986_not n14987_not ; n14988
g14733 and b[1]_not n14982_not ; n14989
g14734 and n14988_not n14989_not ; n14990
g14735 and b[2] n14976_not ; n14991
g14736 and n14974_not n14991 ; n14992
g14737 and n14978_not n14992_not ; n14993
g14738 and n14990_not n14993 ; n14994
g14739 and n14978_not n14994_not ; n14995
g14740 and b[3] n14968_not ; n14996
g14741 and n14966_not n14996 ; n14997
g14742 and n14970_not n14997_not ; n14998
g14743 and n14995_not n14998 ; n14999
g14744 and n14970_not n14999_not ; n15000
g14745 and b[4] n14959_not ; n15001
g14746 and n14957_not n15001 ; n15002
g14747 and n14961_not n15002_not ; n15003
g14748 and n15000_not n15003 ; n15004
g14749 and n14961_not n15004_not ; n15005
g14750 and b[5] n14950_not ; n15006
g14751 and n14948_not n15006 ; n15007
g14752 and n14952_not n15007_not ; n15008
g14753 and n15005_not n15008 ; n15009
g14754 and n14952_not n15009_not ; n15010
g14755 and b[6] n14941_not ; n15011
g14756 and n14939_not n15011 ; n15012
g14757 and n14943_not n15012_not ; n15013
g14758 and n15010_not n15013 ; n15014
g14759 and n14943_not n15014_not ; n15015
g14760 and b[7] n14932_not ; n15016
g14761 and n14930_not n15016 ; n15017
g14762 and n14934_not n15017_not ; n15018
g14763 and n15015_not n15018 ; n15019
g14764 and n14934_not n15019_not ; n15020
g14765 and b[8] n14923_not ; n15021
g14766 and n14921_not n15021 ; n15022
g14767 and n14925_not n15022_not ; n15023
g14768 and n15020_not n15023 ; n15024
g14769 and n14925_not n15024_not ; n15025
g14770 and b[9] n14914_not ; n15026
g14771 and n14912_not n15026 ; n15027
g14772 and n14916_not n15027_not ; n15028
g14773 and n15025_not n15028 ; n15029
g14774 and n14916_not n15029_not ; n15030
g14775 and b[10] n14905_not ; n15031
g14776 and n14903_not n15031 ; n15032
g14777 and n14907_not n15032_not ; n15033
g14778 and n15030_not n15033 ; n15034
g14779 and n14907_not n15034_not ; n15035
g14780 and b[11] n14896_not ; n15036
g14781 and n14894_not n15036 ; n15037
g14782 and n14898_not n15037_not ; n15038
g14783 and n15035_not n15038 ; n15039
g14784 and n14898_not n15039_not ; n15040
g14785 and b[12] n14887_not ; n15041
g14786 and n14885_not n15041 ; n15042
g14787 and n14889_not n15042_not ; n15043
g14788 and n15040_not n15043 ; n15044
g14789 and n14889_not n15044_not ; n15045
g14790 and b[13] n14878_not ; n15046
g14791 and n14876_not n15046 ; n15047
g14792 and n14880_not n15047_not ; n15048
g14793 and n15045_not n15048 ; n15049
g14794 and n14880_not n15049_not ; n15050
g14795 and b[14] n14869_not ; n15051
g14796 and n14867_not n15051 ; n15052
g14797 and n14871_not n15052_not ; n15053
g14798 and n15050_not n15053 ; n15054
g14799 and n14871_not n15054_not ; n15055
g14800 and b[15] n14860_not ; n15056
g14801 and n14858_not n15056 ; n15057
g14802 and n14862_not n15057_not ; n15058
g14803 and n15055_not n15058 ; n15059
g14804 and n14862_not n15059_not ; n15060
g14805 and b[16] n14851_not ; n15061
g14806 and n14849_not n15061 ; n15062
g14807 and n14853_not n15062_not ; n15063
g14808 and n15060_not n15063 ; n15064
g14809 and n14853_not n15064_not ; n15065
g14810 and b[17] n14842_not ; n15066
g14811 and n14840_not n15066 ; n15067
g14812 and n14844_not n15067_not ; n15068
g14813 and n15065_not n15068 ; n15069
g14814 and n14844_not n15069_not ; n15070
g14815 and b[18] n14833_not ; n15071
g14816 and n14831_not n15071 ; n15072
g14817 and n14835_not n15072_not ; n15073
g14818 and n15070_not n15073 ; n15074
g14819 and n14835_not n15074_not ; n15075
g14820 and b[19] n14824_not ; n15076
g14821 and n14822_not n15076 ; n15077
g14822 and n14826_not n15077_not ; n15078
g14823 and n15075_not n15078 ; n15079
g14824 and n14826_not n15079_not ; n15080
g14825 and b[20] n14815_not ; n15081
g14826 and n14813_not n15081 ; n15082
g14827 and n14817_not n15082_not ; n15083
g14828 and n15080_not n15083 ; n15084
g14829 and n14817_not n15084_not ; n15085
g14830 and b[21] n14806_not ; n15086
g14831 and n14804_not n15086 ; n15087
g14832 and n14808_not n15087_not ; n15088
g14833 and n15085_not n15088 ; n15089
g14834 and n14808_not n15089_not ; n15090
g14835 and b[22] n14797_not ; n15091
g14836 and n14795_not n15091 ; n15092
g14837 and n14799_not n15092_not ; n15093
g14838 and n15090_not n15093 ; n15094
g14839 and n14799_not n15094_not ; n15095
g14840 and b[23] n14788_not ; n15096
g14841 and n14786_not n15096 ; n15097
g14842 and n14790_not n15097_not ; n15098
g14843 and n15095_not n15098 ; n15099
g14844 and n14790_not n15099_not ; n15100
g14845 and b[24] n14779_not ; n15101
g14846 and n14777_not n15101 ; n15102
g14847 and n14781_not n15102_not ; n15103
g14848 and n15100_not n15103 ; n15104
g14849 and n14781_not n15104_not ; n15105
g14850 and b[25] n14770_not ; n15106
g14851 and n14768_not n15106 ; n15107
g14852 and n14772_not n15107_not ; n15108
g14853 and n15105_not n15108 ; n15109
g14854 and n14772_not n15109_not ; n15110
g14855 and b[26] n14761_not ; n15111
g14856 and n14759_not n15111 ; n15112
g14857 and n14763_not n15112_not ; n15113
g14858 and n15110_not n15113 ; n15114
g14859 and n14763_not n15114_not ; n15115
g14860 and b[27] n14752_not ; n15116
g14861 and n14750_not n15116 ; n15117
g14862 and n14754_not n15117_not ; n15118
g14863 and n15115_not n15118 ; n15119
g14864 and n14754_not n15119_not ; n15120
g14865 and b[28] n14743_not ; n15121
g14866 and n14741_not n15121 ; n15122
g14867 and n14745_not n15122_not ; n15123
g14868 and n15120_not n15123 ; n15124
g14869 and n14745_not n15124_not ; n15125
g14870 and b[29] n14734_not ; n15126
g14871 and n14732_not n15126 ; n15127
g14872 and n14736_not n15127_not ; n15128
g14873 and n15125_not n15128 ; n15129
g14874 and n14736_not n15129_not ; n15130
g14875 and b[30] n14725_not ; n15131
g14876 and n14723_not n15131 ; n15132
g14877 and n14727_not n15132_not ; n15133
g14878 and n15130_not n15133 ; n15134
g14879 and n14727_not n15134_not ; n15135
g14880 and b[31] n14716_not ; n15136
g14881 and n14714_not n15136 ; n15137
g14882 and n14718_not n15137_not ; n15138
g14883 and n15135_not n15138 ; n15139
g14884 and n14718_not n15139_not ; n15140
g14885 and b[32] n14707_not ; n15141
g14886 and n14705_not n15141 ; n15142
g14887 and n14709_not n15142_not ; n15143
g14888 and n15140_not n15143 ; n15144
g14889 and n14709_not n15144_not ; n15145
g14890 and b[33] n14698_not ; n15146
g14891 and n14696_not n15146 ; n15147
g14892 and n14700_not n15147_not ; n15148
g14893 and n15145_not n15148 ; n15149
g14894 and n14700_not n15149_not ; n15150
g14895 and b[34] n14689_not ; n15151
g14896 and n14687_not n15151 ; n15152
g14897 and n14691_not n15152_not ; n15153
g14898 and n15150_not n15153 ; n15154
g14899 and n14691_not n15154_not ; n15155
g14900 and b[35] n14680_not ; n15156
g14901 and n14678_not n15156 ; n15157
g14902 and n14682_not n15157_not ; n15158
g14903 and n15155_not n15158 ; n15159
g14904 and n14682_not n15159_not ; n15160
g14905 and b[36] n14671_not ; n15161
g14906 and n14669_not n15161 ; n15162
g14907 and n14673_not n15162_not ; n15163
g14908 and n15160_not n15163 ; n15164
g14909 and n14673_not n15164_not ; n15165
g14910 and b[37] n14662_not ; n15166
g14911 and n14660_not n15166 ; n15167
g14912 and n14664_not n15167_not ; n15168
g14913 and n15165_not n15168 ; n15169
g14914 and n14664_not n15169_not ; n15170
g14915 and b[38] n14653_not ; n15171
g14916 and n14651_not n15171 ; n15172
g14917 and n14655_not n15172_not ; n15173
g14918 and n15170_not n15173 ; n15174
g14919 and n14655_not n15174_not ; n15175
g14920 and b[39] n14644_not ; n15176
g14921 and n14642_not n15176 ; n15177
g14922 and n14646_not n15177_not ; n15178
g14923 and n15175_not n15178 ; n15179
g14924 and n14646_not n15179_not ; n15180
g14925 and b[40] n14635_not ; n15181
g14926 and n14633_not n15181 ; n15182
g14927 and n14637_not n15182_not ; n15183
g14928 and n15180_not n15183 ; n15184
g14929 and n14637_not n15184_not ; n15185
g14930 and b[41] n14626_not ; n15186
g14931 and n14624_not n15186 ; n15187
g14932 and n14628_not n15187_not ; n15188
g14933 and n15185_not n15188 ; n15189
g14934 and n14628_not n15189_not ; n15190
g14935 and b[42] n14617_not ; n15191
g14936 and n14615_not n15191 ; n15192
g14937 and n14619_not n15192_not ; n15193
g14938 and n15190_not n15193 ; n15194
g14939 and n14619_not n15194_not ; n15195
g14940 and b[43] n14608_not ; n15196
g14941 and n14606_not n15196 ; n15197
g14942 and n14610_not n15197_not ; n15198
g14943 and n15195_not n15198 ; n15199
g14944 and n14610_not n15199_not ; n15200
g14945 and b[44] n14588_not ; n15201
g14946 and n14586_not n15201 ; n15202
g14947 and n14601_not n15202_not ; n15203
g14948 and n15200_not n15203 ; n15204
g14949 and n14601_not n15204_not ; n15205
g14950 and b[45] n14598_not ; n15206
g14951 and n14596_not n15206 ; n15207
g14952 and n14600_not n15207_not ; n15208
g14953 and n15205_not n15208 ; n15209
g14954 and n14600_not n15209_not ; n15210
g14955 and n298 n300 ; n15211
g14956 and n288 n15211 ; n15212
g14957 and n15210_not n15212 ; quotient[18]
g14958 and n14589_not quotient[18]_not ; n15214
g14959 and n14610_not n15203 ; n15215
g14960 and n15199_not n15215 ; n15216
g14961 and n15200_not n15203_not ; n15217
g14962 and n15216_not n15217_not ; n15218
g14963 and n15212 n15218_not ; n15219
g14964 and n15210_not n15219 ; n15220
g14965 and n15214_not n15220_not ; n15221
g14966 and b[45]_not n15221_not ; n15222
g14967 and n14609_not quotient[18]_not ; n15223
g14968 and n14619_not n15198 ; n15224
g14969 and n15194_not n15224 ; n15225
g14970 and n15195_not n15198_not ; n15226
g14971 and n15225_not n15226_not ; n15227
g14972 and n15212 n15227_not ; n15228
g14973 and n15210_not n15228 ; n15229
g14974 and n15223_not n15229_not ; n15230
g14975 and b[44]_not n15230_not ; n15231
g14976 and n14618_not quotient[18]_not ; n15232
g14977 and n14628_not n15193 ; n15233
g14978 and n15189_not n15233 ; n15234
g14979 and n15190_not n15193_not ; n15235
g14980 and n15234_not n15235_not ; n15236
g14981 and n15212 n15236_not ; n15237
g14982 and n15210_not n15237 ; n15238
g14983 and n15232_not n15238_not ; n15239
g14984 and b[43]_not n15239_not ; n15240
g14985 and n14627_not quotient[18]_not ; n15241
g14986 and n14637_not n15188 ; n15242
g14987 and n15184_not n15242 ; n15243
g14988 and n15185_not n15188_not ; n15244
g14989 and n15243_not n15244_not ; n15245
g14990 and n15212 n15245_not ; n15246
g14991 and n15210_not n15246 ; n15247
g14992 and n15241_not n15247_not ; n15248
g14993 and b[42]_not n15248_not ; n15249
g14994 and n14636_not quotient[18]_not ; n15250
g14995 and n14646_not n15183 ; n15251
g14996 and n15179_not n15251 ; n15252
g14997 and n15180_not n15183_not ; n15253
g14998 and n15252_not n15253_not ; n15254
g14999 and n15212 n15254_not ; n15255
g15000 and n15210_not n15255 ; n15256
g15001 and n15250_not n15256_not ; n15257
g15002 and b[41]_not n15257_not ; n15258
g15003 and n14645_not quotient[18]_not ; n15259
g15004 and n14655_not n15178 ; n15260
g15005 and n15174_not n15260 ; n15261
g15006 and n15175_not n15178_not ; n15262
g15007 and n15261_not n15262_not ; n15263
g15008 and n15212 n15263_not ; n15264
g15009 and n15210_not n15264 ; n15265
g15010 and n15259_not n15265_not ; n15266
g15011 and b[40]_not n15266_not ; n15267
g15012 and n14654_not quotient[18]_not ; n15268
g15013 and n14664_not n15173 ; n15269
g15014 and n15169_not n15269 ; n15270
g15015 and n15170_not n15173_not ; n15271
g15016 and n15270_not n15271_not ; n15272
g15017 and n15212 n15272_not ; n15273
g15018 and n15210_not n15273 ; n15274
g15019 and n15268_not n15274_not ; n15275
g15020 and b[39]_not n15275_not ; n15276
g15021 and n14663_not quotient[18]_not ; n15277
g15022 and n14673_not n15168 ; n15278
g15023 and n15164_not n15278 ; n15279
g15024 and n15165_not n15168_not ; n15280
g15025 and n15279_not n15280_not ; n15281
g15026 and n15212 n15281_not ; n15282
g15027 and n15210_not n15282 ; n15283
g15028 and n15277_not n15283_not ; n15284
g15029 and b[38]_not n15284_not ; n15285
g15030 and n14672_not quotient[18]_not ; n15286
g15031 and n14682_not n15163 ; n15287
g15032 and n15159_not n15287 ; n15288
g15033 and n15160_not n15163_not ; n15289
g15034 and n15288_not n15289_not ; n15290
g15035 and n15212 n15290_not ; n15291
g15036 and n15210_not n15291 ; n15292
g15037 and n15286_not n15292_not ; n15293
g15038 and b[37]_not n15293_not ; n15294
g15039 and n14681_not quotient[18]_not ; n15295
g15040 and n14691_not n15158 ; n15296
g15041 and n15154_not n15296 ; n15297
g15042 and n15155_not n15158_not ; n15298
g15043 and n15297_not n15298_not ; n15299
g15044 and n15212 n15299_not ; n15300
g15045 and n15210_not n15300 ; n15301
g15046 and n15295_not n15301_not ; n15302
g15047 and b[36]_not n15302_not ; n15303
g15048 and n14690_not quotient[18]_not ; n15304
g15049 and n14700_not n15153 ; n15305
g15050 and n15149_not n15305 ; n15306
g15051 and n15150_not n15153_not ; n15307
g15052 and n15306_not n15307_not ; n15308
g15053 and n15212 n15308_not ; n15309
g15054 and n15210_not n15309 ; n15310
g15055 and n15304_not n15310_not ; n15311
g15056 and b[35]_not n15311_not ; n15312
g15057 and n14699_not quotient[18]_not ; n15313
g15058 and n14709_not n15148 ; n15314
g15059 and n15144_not n15314 ; n15315
g15060 and n15145_not n15148_not ; n15316
g15061 and n15315_not n15316_not ; n15317
g15062 and n15212 n15317_not ; n15318
g15063 and n15210_not n15318 ; n15319
g15064 and n15313_not n15319_not ; n15320
g15065 and b[34]_not n15320_not ; n15321
g15066 and n14708_not quotient[18]_not ; n15322
g15067 and n14718_not n15143 ; n15323
g15068 and n15139_not n15323 ; n15324
g15069 and n15140_not n15143_not ; n15325
g15070 and n15324_not n15325_not ; n15326
g15071 and n15212 n15326_not ; n15327
g15072 and n15210_not n15327 ; n15328
g15073 and n15322_not n15328_not ; n15329
g15074 and b[33]_not n15329_not ; n15330
g15075 and n14717_not quotient[18]_not ; n15331
g15076 and n14727_not n15138 ; n15332
g15077 and n15134_not n15332 ; n15333
g15078 and n15135_not n15138_not ; n15334
g15079 and n15333_not n15334_not ; n15335
g15080 and n15212 n15335_not ; n15336
g15081 and n15210_not n15336 ; n15337
g15082 and n15331_not n15337_not ; n15338
g15083 and b[32]_not n15338_not ; n15339
g15084 and n14726_not quotient[18]_not ; n15340
g15085 and n14736_not n15133 ; n15341
g15086 and n15129_not n15341 ; n15342
g15087 and n15130_not n15133_not ; n15343
g15088 and n15342_not n15343_not ; n15344
g15089 and n15212 n15344_not ; n15345
g15090 and n15210_not n15345 ; n15346
g15091 and n15340_not n15346_not ; n15347
g15092 and b[31]_not n15347_not ; n15348
g15093 and n14735_not quotient[18]_not ; n15349
g15094 and n14745_not n15128 ; n15350
g15095 and n15124_not n15350 ; n15351
g15096 and n15125_not n15128_not ; n15352
g15097 and n15351_not n15352_not ; n15353
g15098 and n15212 n15353_not ; n15354
g15099 and n15210_not n15354 ; n15355
g15100 and n15349_not n15355_not ; n15356
g15101 and b[30]_not n15356_not ; n15357
g15102 and n14744_not quotient[18]_not ; n15358
g15103 and n14754_not n15123 ; n15359
g15104 and n15119_not n15359 ; n15360
g15105 and n15120_not n15123_not ; n15361
g15106 and n15360_not n15361_not ; n15362
g15107 and n15212 n15362_not ; n15363
g15108 and n15210_not n15363 ; n15364
g15109 and n15358_not n15364_not ; n15365
g15110 and b[29]_not n15365_not ; n15366
g15111 and n14753_not quotient[18]_not ; n15367
g15112 and n14763_not n15118 ; n15368
g15113 and n15114_not n15368 ; n15369
g15114 and n15115_not n15118_not ; n15370
g15115 and n15369_not n15370_not ; n15371
g15116 and n15212 n15371_not ; n15372
g15117 and n15210_not n15372 ; n15373
g15118 and n15367_not n15373_not ; n15374
g15119 and b[28]_not n15374_not ; n15375
g15120 and n14762_not quotient[18]_not ; n15376
g15121 and n14772_not n15113 ; n15377
g15122 and n15109_not n15377 ; n15378
g15123 and n15110_not n15113_not ; n15379
g15124 and n15378_not n15379_not ; n15380
g15125 and n15212 n15380_not ; n15381
g15126 and n15210_not n15381 ; n15382
g15127 and n15376_not n15382_not ; n15383
g15128 and b[27]_not n15383_not ; n15384
g15129 and n14771_not quotient[18]_not ; n15385
g15130 and n14781_not n15108 ; n15386
g15131 and n15104_not n15386 ; n15387
g15132 and n15105_not n15108_not ; n15388
g15133 and n15387_not n15388_not ; n15389
g15134 and n15212 n15389_not ; n15390
g15135 and n15210_not n15390 ; n15391
g15136 and n15385_not n15391_not ; n15392
g15137 and b[26]_not n15392_not ; n15393
g15138 and n14780_not quotient[18]_not ; n15394
g15139 and n14790_not n15103 ; n15395
g15140 and n15099_not n15395 ; n15396
g15141 and n15100_not n15103_not ; n15397
g15142 and n15396_not n15397_not ; n15398
g15143 and n15212 n15398_not ; n15399
g15144 and n15210_not n15399 ; n15400
g15145 and n15394_not n15400_not ; n15401
g15146 and b[25]_not n15401_not ; n15402
g15147 and n14789_not quotient[18]_not ; n15403
g15148 and n14799_not n15098 ; n15404
g15149 and n15094_not n15404 ; n15405
g15150 and n15095_not n15098_not ; n15406
g15151 and n15405_not n15406_not ; n15407
g15152 and n15212 n15407_not ; n15408
g15153 and n15210_not n15408 ; n15409
g15154 and n15403_not n15409_not ; n15410
g15155 and b[24]_not n15410_not ; n15411
g15156 and n14798_not quotient[18]_not ; n15412
g15157 and n14808_not n15093 ; n15413
g15158 and n15089_not n15413 ; n15414
g15159 and n15090_not n15093_not ; n15415
g15160 and n15414_not n15415_not ; n15416
g15161 and n15212 n15416_not ; n15417
g15162 and n15210_not n15417 ; n15418
g15163 and n15412_not n15418_not ; n15419
g15164 and b[23]_not n15419_not ; n15420
g15165 and n14807_not quotient[18]_not ; n15421
g15166 and n14817_not n15088 ; n15422
g15167 and n15084_not n15422 ; n15423
g15168 and n15085_not n15088_not ; n15424
g15169 and n15423_not n15424_not ; n15425
g15170 and n15212 n15425_not ; n15426
g15171 and n15210_not n15426 ; n15427
g15172 and n15421_not n15427_not ; n15428
g15173 and b[22]_not n15428_not ; n15429
g15174 and n14816_not quotient[18]_not ; n15430
g15175 and n14826_not n15083 ; n15431
g15176 and n15079_not n15431 ; n15432
g15177 and n15080_not n15083_not ; n15433
g15178 and n15432_not n15433_not ; n15434
g15179 and n15212 n15434_not ; n15435
g15180 and n15210_not n15435 ; n15436
g15181 and n15430_not n15436_not ; n15437
g15182 and b[21]_not n15437_not ; n15438
g15183 and n14825_not quotient[18]_not ; n15439
g15184 and n14835_not n15078 ; n15440
g15185 and n15074_not n15440 ; n15441
g15186 and n15075_not n15078_not ; n15442
g15187 and n15441_not n15442_not ; n15443
g15188 and n15212 n15443_not ; n15444
g15189 and n15210_not n15444 ; n15445
g15190 and n15439_not n15445_not ; n15446
g15191 and b[20]_not n15446_not ; n15447
g15192 and n14834_not quotient[18]_not ; n15448
g15193 and n14844_not n15073 ; n15449
g15194 and n15069_not n15449 ; n15450
g15195 and n15070_not n15073_not ; n15451
g15196 and n15450_not n15451_not ; n15452
g15197 and n15212 n15452_not ; n15453
g15198 and n15210_not n15453 ; n15454
g15199 and n15448_not n15454_not ; n15455
g15200 and b[19]_not n15455_not ; n15456
g15201 and n14843_not quotient[18]_not ; n15457
g15202 and n14853_not n15068 ; n15458
g15203 and n15064_not n15458 ; n15459
g15204 and n15065_not n15068_not ; n15460
g15205 and n15459_not n15460_not ; n15461
g15206 and n15212 n15461_not ; n15462
g15207 and n15210_not n15462 ; n15463
g15208 and n15457_not n15463_not ; n15464
g15209 and b[18]_not n15464_not ; n15465
g15210 and n14852_not quotient[18]_not ; n15466
g15211 and n14862_not n15063 ; n15467
g15212 and n15059_not n15467 ; n15468
g15213 and n15060_not n15063_not ; n15469
g15214 and n15468_not n15469_not ; n15470
g15215 and n15212 n15470_not ; n15471
g15216 and n15210_not n15471 ; n15472
g15217 and n15466_not n15472_not ; n15473
g15218 and b[17]_not n15473_not ; n15474
g15219 and n14861_not quotient[18]_not ; n15475
g15220 and n14871_not n15058 ; n15476
g15221 and n15054_not n15476 ; n15477
g15222 and n15055_not n15058_not ; n15478
g15223 and n15477_not n15478_not ; n15479
g15224 and n15212 n15479_not ; n15480
g15225 and n15210_not n15480 ; n15481
g15226 and n15475_not n15481_not ; n15482
g15227 and b[16]_not n15482_not ; n15483
g15228 and n14870_not quotient[18]_not ; n15484
g15229 and n14880_not n15053 ; n15485
g15230 and n15049_not n15485 ; n15486
g15231 and n15050_not n15053_not ; n15487
g15232 and n15486_not n15487_not ; n15488
g15233 and n15212 n15488_not ; n15489
g15234 and n15210_not n15489 ; n15490
g15235 and n15484_not n15490_not ; n15491
g15236 and b[15]_not n15491_not ; n15492
g15237 and n14879_not quotient[18]_not ; n15493
g15238 and n14889_not n15048 ; n15494
g15239 and n15044_not n15494 ; n15495
g15240 and n15045_not n15048_not ; n15496
g15241 and n15495_not n15496_not ; n15497
g15242 and n15212 n15497_not ; n15498
g15243 and n15210_not n15498 ; n15499
g15244 and n15493_not n15499_not ; n15500
g15245 and b[14]_not n15500_not ; n15501
g15246 and n14888_not quotient[18]_not ; n15502
g15247 and n14898_not n15043 ; n15503
g15248 and n15039_not n15503 ; n15504
g15249 and n15040_not n15043_not ; n15505
g15250 and n15504_not n15505_not ; n15506
g15251 and n15212 n15506_not ; n15507
g15252 and n15210_not n15507 ; n15508
g15253 and n15502_not n15508_not ; n15509
g15254 and b[13]_not n15509_not ; n15510
g15255 and n14897_not quotient[18]_not ; n15511
g15256 and n14907_not n15038 ; n15512
g15257 and n15034_not n15512 ; n15513
g15258 and n15035_not n15038_not ; n15514
g15259 and n15513_not n15514_not ; n15515
g15260 and n15212 n15515_not ; n15516
g15261 and n15210_not n15516 ; n15517
g15262 and n15511_not n15517_not ; n15518
g15263 and b[12]_not n15518_not ; n15519
g15264 and n14906_not quotient[18]_not ; n15520
g15265 and n14916_not n15033 ; n15521
g15266 and n15029_not n15521 ; n15522
g15267 and n15030_not n15033_not ; n15523
g15268 and n15522_not n15523_not ; n15524
g15269 and n15212 n15524_not ; n15525
g15270 and n15210_not n15525 ; n15526
g15271 and n15520_not n15526_not ; n15527
g15272 and b[11]_not n15527_not ; n15528
g15273 and n14915_not quotient[18]_not ; n15529
g15274 and n14925_not n15028 ; n15530
g15275 and n15024_not n15530 ; n15531
g15276 and n15025_not n15028_not ; n15532
g15277 and n15531_not n15532_not ; n15533
g15278 and n15212 n15533_not ; n15534
g15279 and n15210_not n15534 ; n15535
g15280 and n15529_not n15535_not ; n15536
g15281 and b[10]_not n15536_not ; n15537
g15282 and n14924_not quotient[18]_not ; n15538
g15283 and n14934_not n15023 ; n15539
g15284 and n15019_not n15539 ; n15540
g15285 and n15020_not n15023_not ; n15541
g15286 and n15540_not n15541_not ; n15542
g15287 and n15212 n15542_not ; n15543
g15288 and n15210_not n15543 ; n15544
g15289 and n15538_not n15544_not ; n15545
g15290 and b[9]_not n15545_not ; n15546
g15291 and n14933_not quotient[18]_not ; n15547
g15292 and n14943_not n15018 ; n15548
g15293 and n15014_not n15548 ; n15549
g15294 and n15015_not n15018_not ; n15550
g15295 and n15549_not n15550_not ; n15551
g15296 and n15212 n15551_not ; n15552
g15297 and n15210_not n15552 ; n15553
g15298 and n15547_not n15553_not ; n15554
g15299 and b[8]_not n15554_not ; n15555
g15300 and n14942_not quotient[18]_not ; n15556
g15301 and n14952_not n15013 ; n15557
g15302 and n15009_not n15557 ; n15558
g15303 and n15010_not n15013_not ; n15559
g15304 and n15558_not n15559_not ; n15560
g15305 and n15212 n15560_not ; n15561
g15306 and n15210_not n15561 ; n15562
g15307 and n15556_not n15562_not ; n15563
g15308 and b[7]_not n15563_not ; n15564
g15309 and n14951_not quotient[18]_not ; n15565
g15310 and n14961_not n15008 ; n15566
g15311 and n15004_not n15566 ; n15567
g15312 and n15005_not n15008_not ; n15568
g15313 and n15567_not n15568_not ; n15569
g15314 and n15212 n15569_not ; n15570
g15315 and n15210_not n15570 ; n15571
g15316 and n15565_not n15571_not ; n15572
g15317 and b[6]_not n15572_not ; n15573
g15318 and n14960_not quotient[18]_not ; n15574
g15319 and n14970_not n15003 ; n15575
g15320 and n14999_not n15575 ; n15576
g15321 and n15000_not n15003_not ; n15577
g15322 and n15576_not n15577_not ; n15578
g15323 and n15212 n15578_not ; n15579
g15324 and n15210_not n15579 ; n15580
g15325 and n15574_not n15580_not ; n15581
g15326 and b[5]_not n15581_not ; n15582
g15327 and n14969_not quotient[18]_not ; n15583
g15328 and n14978_not n14998 ; n15584
g15329 and n14994_not n15584 ; n15585
g15330 and n14995_not n14998_not ; n15586
g15331 and n15585_not n15586_not ; n15587
g15332 and n15212 n15587_not ; n15588
g15333 and n15210_not n15588 ; n15589
g15334 and n15583_not n15589_not ; n15590
g15335 and b[4]_not n15590_not ; n15591
g15336 and n14977_not quotient[18]_not ; n15592
g15337 and n14989_not n14993 ; n15593
g15338 and n14988_not n15593 ; n15594
g15339 and n14990_not n14993_not ; n15595
g15340 and n15594_not n15595_not ; n15596
g15341 and n15212 n15596_not ; n15597
g15342 and n15210_not n15597 ; n15598
g15343 and n15592_not n15598_not ; n15599
g15344 and b[3]_not n15599_not ; n15600
g15345 and n14982_not quotient[18]_not ; n15601
g15346 and n14985_not n14987 ; n15602
g15347 and n14983_not n15602 ; n15603
g15348 and n15212 n15603_not ; n15604
g15349 and n14988_not n15604 ; n15605
g15350 and n15210_not n15605 ; n15606
g15351 and n15601_not n15606_not ; n15607
g15352 and b[2]_not n15607_not ; n15608
g15353 and b[0] b[46]_not ; n15609
g15354 and n417 n15609 ; n15610
g15355 and n400 n15610 ; n15611
g15356 and n595 n15611 ; n15612
g15357 and n15210_not n15612 ; n15613
g15358 and a[18] n15613_not ; n15614
g15359 and n300 n14987 ; n15615
g15360 and n298 n15615 ; n15616
g15361 and n288 n15616 ; n15617
g15362 and n15210_not n15617 ; n15618
g15363 and n15614_not n15618_not ; n15619
g15364 and b[1] n15619_not ; n15620
g15365 and b[1]_not n15618_not ; n15621
g15366 and n15614_not n15621 ; n15622
g15367 and n15620_not n15622_not ; n15623
g15368 and a[17]_not b[0] ; n15624
g15369 and n15623_not n15624_not ; n15625
g15370 and b[1]_not n15619_not ; n15626
g15371 and n15625_not n15626_not ; n15627
g15372 and b[2] n15606_not ; n15628
g15373 and n15601_not n15628 ; n15629
g15374 and n15608_not n15629_not ; n15630
g15375 and n15627_not n15630 ; n15631
g15376 and n15608_not n15631_not ; n15632
g15377 and b[3] n15598_not ; n15633
g15378 and n15592_not n15633 ; n15634
g15379 and n15600_not n15634_not ; n15635
g15380 and n15632_not n15635 ; n15636
g15381 and n15600_not n15636_not ; n15637
g15382 and b[4] n15589_not ; n15638
g15383 and n15583_not n15638 ; n15639
g15384 and n15591_not n15639_not ; n15640
g15385 and n15637_not n15640 ; n15641
g15386 and n15591_not n15641_not ; n15642
g15387 and b[5] n15580_not ; n15643
g15388 and n15574_not n15643 ; n15644
g15389 and n15582_not n15644_not ; n15645
g15390 and n15642_not n15645 ; n15646
g15391 and n15582_not n15646_not ; n15647
g15392 and b[6] n15571_not ; n15648
g15393 and n15565_not n15648 ; n15649
g15394 and n15573_not n15649_not ; n15650
g15395 and n15647_not n15650 ; n15651
g15396 and n15573_not n15651_not ; n15652
g15397 and b[7] n15562_not ; n15653
g15398 and n15556_not n15653 ; n15654
g15399 and n15564_not n15654_not ; n15655
g15400 and n15652_not n15655 ; n15656
g15401 and n15564_not n15656_not ; n15657
g15402 and b[8] n15553_not ; n15658
g15403 and n15547_not n15658 ; n15659
g15404 and n15555_not n15659_not ; n15660
g15405 and n15657_not n15660 ; n15661
g15406 and n15555_not n15661_not ; n15662
g15407 and b[9] n15544_not ; n15663
g15408 and n15538_not n15663 ; n15664
g15409 and n15546_not n15664_not ; n15665
g15410 and n15662_not n15665 ; n15666
g15411 and n15546_not n15666_not ; n15667
g15412 and b[10] n15535_not ; n15668
g15413 and n15529_not n15668 ; n15669
g15414 and n15537_not n15669_not ; n15670
g15415 and n15667_not n15670 ; n15671
g15416 and n15537_not n15671_not ; n15672
g15417 and b[11] n15526_not ; n15673
g15418 and n15520_not n15673 ; n15674
g15419 and n15528_not n15674_not ; n15675
g15420 and n15672_not n15675 ; n15676
g15421 and n15528_not n15676_not ; n15677
g15422 and b[12] n15517_not ; n15678
g15423 and n15511_not n15678 ; n15679
g15424 and n15519_not n15679_not ; n15680
g15425 and n15677_not n15680 ; n15681
g15426 and n15519_not n15681_not ; n15682
g15427 and b[13] n15508_not ; n15683
g15428 and n15502_not n15683 ; n15684
g15429 and n15510_not n15684_not ; n15685
g15430 and n15682_not n15685 ; n15686
g15431 and n15510_not n15686_not ; n15687
g15432 and b[14] n15499_not ; n15688
g15433 and n15493_not n15688 ; n15689
g15434 and n15501_not n15689_not ; n15690
g15435 and n15687_not n15690 ; n15691
g15436 and n15501_not n15691_not ; n15692
g15437 and b[15] n15490_not ; n15693
g15438 and n15484_not n15693 ; n15694
g15439 and n15492_not n15694_not ; n15695
g15440 and n15692_not n15695 ; n15696
g15441 and n15492_not n15696_not ; n15697
g15442 and b[16] n15481_not ; n15698
g15443 and n15475_not n15698 ; n15699
g15444 and n15483_not n15699_not ; n15700
g15445 and n15697_not n15700 ; n15701
g15446 and n15483_not n15701_not ; n15702
g15447 and b[17] n15472_not ; n15703
g15448 and n15466_not n15703 ; n15704
g15449 and n15474_not n15704_not ; n15705
g15450 and n15702_not n15705 ; n15706
g15451 and n15474_not n15706_not ; n15707
g15452 and b[18] n15463_not ; n15708
g15453 and n15457_not n15708 ; n15709
g15454 and n15465_not n15709_not ; n15710
g15455 and n15707_not n15710 ; n15711
g15456 and n15465_not n15711_not ; n15712
g15457 and b[19] n15454_not ; n15713
g15458 and n15448_not n15713 ; n15714
g15459 and n15456_not n15714_not ; n15715
g15460 and n15712_not n15715 ; n15716
g15461 and n15456_not n15716_not ; n15717
g15462 and b[20] n15445_not ; n15718
g15463 and n15439_not n15718 ; n15719
g15464 and n15447_not n15719_not ; n15720
g15465 and n15717_not n15720 ; n15721
g15466 and n15447_not n15721_not ; n15722
g15467 and b[21] n15436_not ; n15723
g15468 and n15430_not n15723 ; n15724
g15469 and n15438_not n15724_not ; n15725
g15470 and n15722_not n15725 ; n15726
g15471 and n15438_not n15726_not ; n15727
g15472 and b[22] n15427_not ; n15728
g15473 and n15421_not n15728 ; n15729
g15474 and n15429_not n15729_not ; n15730
g15475 and n15727_not n15730 ; n15731
g15476 and n15429_not n15731_not ; n15732
g15477 and b[23] n15418_not ; n15733
g15478 and n15412_not n15733 ; n15734
g15479 and n15420_not n15734_not ; n15735
g15480 and n15732_not n15735 ; n15736
g15481 and n15420_not n15736_not ; n15737
g15482 and b[24] n15409_not ; n15738
g15483 and n15403_not n15738 ; n15739
g15484 and n15411_not n15739_not ; n15740
g15485 and n15737_not n15740 ; n15741
g15486 and n15411_not n15741_not ; n15742
g15487 and b[25] n15400_not ; n15743
g15488 and n15394_not n15743 ; n15744
g15489 and n15402_not n15744_not ; n15745
g15490 and n15742_not n15745 ; n15746
g15491 and n15402_not n15746_not ; n15747
g15492 and b[26] n15391_not ; n15748
g15493 and n15385_not n15748 ; n15749
g15494 and n15393_not n15749_not ; n15750
g15495 and n15747_not n15750 ; n15751
g15496 and n15393_not n15751_not ; n15752
g15497 and b[27] n15382_not ; n15753
g15498 and n15376_not n15753 ; n15754
g15499 and n15384_not n15754_not ; n15755
g15500 and n15752_not n15755 ; n15756
g15501 and n15384_not n15756_not ; n15757
g15502 and b[28] n15373_not ; n15758
g15503 and n15367_not n15758 ; n15759
g15504 and n15375_not n15759_not ; n15760
g15505 and n15757_not n15760 ; n15761
g15506 and n15375_not n15761_not ; n15762
g15507 and b[29] n15364_not ; n15763
g15508 and n15358_not n15763 ; n15764
g15509 and n15366_not n15764_not ; n15765
g15510 and n15762_not n15765 ; n15766
g15511 and n15366_not n15766_not ; n15767
g15512 and b[30] n15355_not ; n15768
g15513 and n15349_not n15768 ; n15769
g15514 and n15357_not n15769_not ; n15770
g15515 and n15767_not n15770 ; n15771
g15516 and n15357_not n15771_not ; n15772
g15517 and b[31] n15346_not ; n15773
g15518 and n15340_not n15773 ; n15774
g15519 and n15348_not n15774_not ; n15775
g15520 and n15772_not n15775 ; n15776
g15521 and n15348_not n15776_not ; n15777
g15522 and b[32] n15337_not ; n15778
g15523 and n15331_not n15778 ; n15779
g15524 and n15339_not n15779_not ; n15780
g15525 and n15777_not n15780 ; n15781
g15526 and n15339_not n15781_not ; n15782
g15527 and b[33] n15328_not ; n15783
g15528 and n15322_not n15783 ; n15784
g15529 and n15330_not n15784_not ; n15785
g15530 and n15782_not n15785 ; n15786
g15531 and n15330_not n15786_not ; n15787
g15532 and b[34] n15319_not ; n15788
g15533 and n15313_not n15788 ; n15789
g15534 and n15321_not n15789_not ; n15790
g15535 and n15787_not n15790 ; n15791
g15536 and n15321_not n15791_not ; n15792
g15537 and b[35] n15310_not ; n15793
g15538 and n15304_not n15793 ; n15794
g15539 and n15312_not n15794_not ; n15795
g15540 and n15792_not n15795 ; n15796
g15541 and n15312_not n15796_not ; n15797
g15542 and b[36] n15301_not ; n15798
g15543 and n15295_not n15798 ; n15799
g15544 and n15303_not n15799_not ; n15800
g15545 and n15797_not n15800 ; n15801
g15546 and n15303_not n15801_not ; n15802
g15547 and b[37] n15292_not ; n15803
g15548 and n15286_not n15803 ; n15804
g15549 and n15294_not n15804_not ; n15805
g15550 and n15802_not n15805 ; n15806
g15551 and n15294_not n15806_not ; n15807
g15552 and b[38] n15283_not ; n15808
g15553 and n15277_not n15808 ; n15809
g15554 and n15285_not n15809_not ; n15810
g15555 and n15807_not n15810 ; n15811
g15556 and n15285_not n15811_not ; n15812
g15557 and b[39] n15274_not ; n15813
g15558 and n15268_not n15813 ; n15814
g15559 and n15276_not n15814_not ; n15815
g15560 and n15812_not n15815 ; n15816
g15561 and n15276_not n15816_not ; n15817
g15562 and b[40] n15265_not ; n15818
g15563 and n15259_not n15818 ; n15819
g15564 and n15267_not n15819_not ; n15820
g15565 and n15817_not n15820 ; n15821
g15566 and n15267_not n15821_not ; n15822
g15567 and b[41] n15256_not ; n15823
g15568 and n15250_not n15823 ; n15824
g15569 and n15258_not n15824_not ; n15825
g15570 and n15822_not n15825 ; n15826
g15571 and n15258_not n15826_not ; n15827
g15572 and b[42] n15247_not ; n15828
g15573 and n15241_not n15828 ; n15829
g15574 and n15249_not n15829_not ; n15830
g15575 and n15827_not n15830 ; n15831
g15576 and n15249_not n15831_not ; n15832
g15577 and b[43] n15238_not ; n15833
g15578 and n15232_not n15833 ; n15834
g15579 and n15240_not n15834_not ; n15835
g15580 and n15832_not n15835 ; n15836
g15581 and n15240_not n15836_not ; n15837
g15582 and b[44] n15229_not ; n15838
g15583 and n15223_not n15838 ; n15839
g15584 and n15231_not n15839_not ; n15840
g15585 and n15837_not n15840 ; n15841
g15586 and n15231_not n15841_not ; n15842
g15587 and b[45] n15220_not ; n15843
g15588 and n15214_not n15843 ; n15844
g15589 and n15222_not n15844_not ; n15845
g15590 and n15842_not n15845 ; n15846
g15591 and n15222_not n15846_not ; n15847
g15592 and n14599_not quotient[18]_not ; n15848
g15593 and n14601_not n15208 ; n15849
g15594 and n15204_not n15849 ; n15850
g15595 and n15205_not n15208_not ; n15851
g15596 and n15850_not n15851_not ; n15852
g15597 and quotient[18] n15852_not ; n15853
g15598 and n15848_not n15853_not ; n15854
g15599 and b[46]_not n15854_not ; n15855
g15600 and b[46] n15848_not ; n15856
g15601 and n15853_not n15856 ; n15857
g15602 and n400 n417 ; n15858
g15603 and n595 n15858 ; n15859
g15604 and n15857_not n15859 ; n15860
g15605 and n15855_not n15860 ; n15861
g15606 and n15847_not n15861 ; n15862
g15607 and n15212 n15854_not ; n15863
g15608 and n15862_not n15863_not ; quotient[17]
g15609 and n15231_not n15845 ; n15865
g15610 and n15841_not n15865 ; n15866
g15611 and n15842_not n15845_not ; n15867
g15612 and n15866_not n15867_not ; n15868
g15613 and quotient[17] n15868_not ; n15869
g15614 and n15221_not n15863_not ; n15870
g15615 and n15862_not n15870 ; n15871
g15616 and n15869_not n15871_not ; n15872
g15617 and b[46]_not n15872_not ; n15873
g15618 and n15240_not n15840 ; n15874
g15619 and n15836_not n15874 ; n15875
g15620 and n15837_not n15840_not ; n15876
g15621 and n15875_not n15876_not ; n15877
g15622 and quotient[17] n15877_not ; n15878
g15623 and n15230_not n15863_not ; n15879
g15624 and n15862_not n15879 ; n15880
g15625 and n15878_not n15880_not ; n15881
g15626 and b[45]_not n15881_not ; n15882
g15627 and n15249_not n15835 ; n15883
g15628 and n15831_not n15883 ; n15884
g15629 and n15832_not n15835_not ; n15885
g15630 and n15884_not n15885_not ; n15886
g15631 and quotient[17] n15886_not ; n15887
g15632 and n15239_not n15863_not ; n15888
g15633 and n15862_not n15888 ; n15889
g15634 and n15887_not n15889_not ; n15890
g15635 and b[44]_not n15890_not ; n15891
g15636 and n15258_not n15830 ; n15892
g15637 and n15826_not n15892 ; n15893
g15638 and n15827_not n15830_not ; n15894
g15639 and n15893_not n15894_not ; n15895
g15640 and quotient[17] n15895_not ; n15896
g15641 and n15248_not n15863_not ; n15897
g15642 and n15862_not n15897 ; n15898
g15643 and n15896_not n15898_not ; n15899
g15644 and b[43]_not n15899_not ; n15900
g15645 and n15267_not n15825 ; n15901
g15646 and n15821_not n15901 ; n15902
g15647 and n15822_not n15825_not ; n15903
g15648 and n15902_not n15903_not ; n15904
g15649 and quotient[17] n15904_not ; n15905
g15650 and n15257_not n15863_not ; n15906
g15651 and n15862_not n15906 ; n15907
g15652 and n15905_not n15907_not ; n15908
g15653 and b[42]_not n15908_not ; n15909
g15654 and n15276_not n15820 ; n15910
g15655 and n15816_not n15910 ; n15911
g15656 and n15817_not n15820_not ; n15912
g15657 and n15911_not n15912_not ; n15913
g15658 and quotient[17] n15913_not ; n15914
g15659 and n15266_not n15863_not ; n15915
g15660 and n15862_not n15915 ; n15916
g15661 and n15914_not n15916_not ; n15917
g15662 and b[41]_not n15917_not ; n15918
g15663 and n15285_not n15815 ; n15919
g15664 and n15811_not n15919 ; n15920
g15665 and n15812_not n15815_not ; n15921
g15666 and n15920_not n15921_not ; n15922
g15667 and quotient[17] n15922_not ; n15923
g15668 and n15275_not n15863_not ; n15924
g15669 and n15862_not n15924 ; n15925
g15670 and n15923_not n15925_not ; n15926
g15671 and b[40]_not n15926_not ; n15927
g15672 and n15294_not n15810 ; n15928
g15673 and n15806_not n15928 ; n15929
g15674 and n15807_not n15810_not ; n15930
g15675 and n15929_not n15930_not ; n15931
g15676 and quotient[17] n15931_not ; n15932
g15677 and n15284_not n15863_not ; n15933
g15678 and n15862_not n15933 ; n15934
g15679 and n15932_not n15934_not ; n15935
g15680 and b[39]_not n15935_not ; n15936
g15681 and n15303_not n15805 ; n15937
g15682 and n15801_not n15937 ; n15938
g15683 and n15802_not n15805_not ; n15939
g15684 and n15938_not n15939_not ; n15940
g15685 and quotient[17] n15940_not ; n15941
g15686 and n15293_not n15863_not ; n15942
g15687 and n15862_not n15942 ; n15943
g15688 and n15941_not n15943_not ; n15944
g15689 and b[38]_not n15944_not ; n15945
g15690 and n15312_not n15800 ; n15946
g15691 and n15796_not n15946 ; n15947
g15692 and n15797_not n15800_not ; n15948
g15693 and n15947_not n15948_not ; n15949
g15694 and quotient[17] n15949_not ; n15950
g15695 and n15302_not n15863_not ; n15951
g15696 and n15862_not n15951 ; n15952
g15697 and n15950_not n15952_not ; n15953
g15698 and b[37]_not n15953_not ; n15954
g15699 and n15321_not n15795 ; n15955
g15700 and n15791_not n15955 ; n15956
g15701 and n15792_not n15795_not ; n15957
g15702 and n15956_not n15957_not ; n15958
g15703 and quotient[17] n15958_not ; n15959
g15704 and n15311_not n15863_not ; n15960
g15705 and n15862_not n15960 ; n15961
g15706 and n15959_not n15961_not ; n15962
g15707 and b[36]_not n15962_not ; n15963
g15708 and n15330_not n15790 ; n15964
g15709 and n15786_not n15964 ; n15965
g15710 and n15787_not n15790_not ; n15966
g15711 and n15965_not n15966_not ; n15967
g15712 and quotient[17] n15967_not ; n15968
g15713 and n15320_not n15863_not ; n15969
g15714 and n15862_not n15969 ; n15970
g15715 and n15968_not n15970_not ; n15971
g15716 and b[35]_not n15971_not ; n15972
g15717 and n15339_not n15785 ; n15973
g15718 and n15781_not n15973 ; n15974
g15719 and n15782_not n15785_not ; n15975
g15720 and n15974_not n15975_not ; n15976
g15721 and quotient[17] n15976_not ; n15977
g15722 and n15329_not n15863_not ; n15978
g15723 and n15862_not n15978 ; n15979
g15724 and n15977_not n15979_not ; n15980
g15725 and b[34]_not n15980_not ; n15981
g15726 and n15348_not n15780 ; n15982
g15727 and n15776_not n15982 ; n15983
g15728 and n15777_not n15780_not ; n15984
g15729 and n15983_not n15984_not ; n15985
g15730 and quotient[17] n15985_not ; n15986
g15731 and n15338_not n15863_not ; n15987
g15732 and n15862_not n15987 ; n15988
g15733 and n15986_not n15988_not ; n15989
g15734 and b[33]_not n15989_not ; n15990
g15735 and n15357_not n15775 ; n15991
g15736 and n15771_not n15991 ; n15992
g15737 and n15772_not n15775_not ; n15993
g15738 and n15992_not n15993_not ; n15994
g15739 and quotient[17] n15994_not ; n15995
g15740 and n15347_not n15863_not ; n15996
g15741 and n15862_not n15996 ; n15997
g15742 and n15995_not n15997_not ; n15998
g15743 and b[32]_not n15998_not ; n15999
g15744 and n15366_not n15770 ; n16000
g15745 and n15766_not n16000 ; n16001
g15746 and n15767_not n15770_not ; n16002
g15747 and n16001_not n16002_not ; n16003
g15748 and quotient[17] n16003_not ; n16004
g15749 and n15356_not n15863_not ; n16005
g15750 and n15862_not n16005 ; n16006
g15751 and n16004_not n16006_not ; n16007
g15752 and b[31]_not n16007_not ; n16008
g15753 and n15375_not n15765 ; n16009
g15754 and n15761_not n16009 ; n16010
g15755 and n15762_not n15765_not ; n16011
g15756 and n16010_not n16011_not ; n16012
g15757 and quotient[17] n16012_not ; n16013
g15758 and n15365_not n15863_not ; n16014
g15759 and n15862_not n16014 ; n16015
g15760 and n16013_not n16015_not ; n16016
g15761 and b[30]_not n16016_not ; n16017
g15762 and n15384_not n15760 ; n16018
g15763 and n15756_not n16018 ; n16019
g15764 and n15757_not n15760_not ; n16020
g15765 and n16019_not n16020_not ; n16021
g15766 and quotient[17] n16021_not ; n16022
g15767 and n15374_not n15863_not ; n16023
g15768 and n15862_not n16023 ; n16024
g15769 and n16022_not n16024_not ; n16025
g15770 and b[29]_not n16025_not ; n16026
g15771 and n15393_not n15755 ; n16027
g15772 and n15751_not n16027 ; n16028
g15773 and n15752_not n15755_not ; n16029
g15774 and n16028_not n16029_not ; n16030
g15775 and quotient[17] n16030_not ; n16031
g15776 and n15383_not n15863_not ; n16032
g15777 and n15862_not n16032 ; n16033
g15778 and n16031_not n16033_not ; n16034
g15779 and b[28]_not n16034_not ; n16035
g15780 and n15402_not n15750 ; n16036
g15781 and n15746_not n16036 ; n16037
g15782 and n15747_not n15750_not ; n16038
g15783 and n16037_not n16038_not ; n16039
g15784 and quotient[17] n16039_not ; n16040
g15785 and n15392_not n15863_not ; n16041
g15786 and n15862_not n16041 ; n16042
g15787 and n16040_not n16042_not ; n16043
g15788 and b[27]_not n16043_not ; n16044
g15789 and n15411_not n15745 ; n16045
g15790 and n15741_not n16045 ; n16046
g15791 and n15742_not n15745_not ; n16047
g15792 and n16046_not n16047_not ; n16048
g15793 and quotient[17] n16048_not ; n16049
g15794 and n15401_not n15863_not ; n16050
g15795 and n15862_not n16050 ; n16051
g15796 and n16049_not n16051_not ; n16052
g15797 and b[26]_not n16052_not ; n16053
g15798 and n15420_not n15740 ; n16054
g15799 and n15736_not n16054 ; n16055
g15800 and n15737_not n15740_not ; n16056
g15801 and n16055_not n16056_not ; n16057
g15802 and quotient[17] n16057_not ; n16058
g15803 and n15410_not n15863_not ; n16059
g15804 and n15862_not n16059 ; n16060
g15805 and n16058_not n16060_not ; n16061
g15806 and b[25]_not n16061_not ; n16062
g15807 and n15429_not n15735 ; n16063
g15808 and n15731_not n16063 ; n16064
g15809 and n15732_not n15735_not ; n16065
g15810 and n16064_not n16065_not ; n16066
g15811 and quotient[17] n16066_not ; n16067
g15812 and n15419_not n15863_not ; n16068
g15813 and n15862_not n16068 ; n16069
g15814 and n16067_not n16069_not ; n16070
g15815 and b[24]_not n16070_not ; n16071
g15816 and n15438_not n15730 ; n16072
g15817 and n15726_not n16072 ; n16073
g15818 and n15727_not n15730_not ; n16074
g15819 and n16073_not n16074_not ; n16075
g15820 and quotient[17] n16075_not ; n16076
g15821 and n15428_not n15863_not ; n16077
g15822 and n15862_not n16077 ; n16078
g15823 and n16076_not n16078_not ; n16079
g15824 and b[23]_not n16079_not ; n16080
g15825 and n15447_not n15725 ; n16081
g15826 and n15721_not n16081 ; n16082
g15827 and n15722_not n15725_not ; n16083
g15828 and n16082_not n16083_not ; n16084
g15829 and quotient[17] n16084_not ; n16085
g15830 and n15437_not n15863_not ; n16086
g15831 and n15862_not n16086 ; n16087
g15832 and n16085_not n16087_not ; n16088
g15833 and b[22]_not n16088_not ; n16089
g15834 and n15456_not n15720 ; n16090
g15835 and n15716_not n16090 ; n16091
g15836 and n15717_not n15720_not ; n16092
g15837 and n16091_not n16092_not ; n16093
g15838 and quotient[17] n16093_not ; n16094
g15839 and n15446_not n15863_not ; n16095
g15840 and n15862_not n16095 ; n16096
g15841 and n16094_not n16096_not ; n16097
g15842 and b[21]_not n16097_not ; n16098
g15843 and n15465_not n15715 ; n16099
g15844 and n15711_not n16099 ; n16100
g15845 and n15712_not n15715_not ; n16101
g15846 and n16100_not n16101_not ; n16102
g15847 and quotient[17] n16102_not ; n16103
g15848 and n15455_not n15863_not ; n16104
g15849 and n15862_not n16104 ; n16105
g15850 and n16103_not n16105_not ; n16106
g15851 and b[20]_not n16106_not ; n16107
g15852 and n15474_not n15710 ; n16108
g15853 and n15706_not n16108 ; n16109
g15854 and n15707_not n15710_not ; n16110
g15855 and n16109_not n16110_not ; n16111
g15856 and quotient[17] n16111_not ; n16112
g15857 and n15464_not n15863_not ; n16113
g15858 and n15862_not n16113 ; n16114
g15859 and n16112_not n16114_not ; n16115
g15860 and b[19]_not n16115_not ; n16116
g15861 and n15483_not n15705 ; n16117
g15862 and n15701_not n16117 ; n16118
g15863 and n15702_not n15705_not ; n16119
g15864 and n16118_not n16119_not ; n16120
g15865 and quotient[17] n16120_not ; n16121
g15866 and n15473_not n15863_not ; n16122
g15867 and n15862_not n16122 ; n16123
g15868 and n16121_not n16123_not ; n16124
g15869 and b[18]_not n16124_not ; n16125
g15870 and n15492_not n15700 ; n16126
g15871 and n15696_not n16126 ; n16127
g15872 and n15697_not n15700_not ; n16128
g15873 and n16127_not n16128_not ; n16129
g15874 and quotient[17] n16129_not ; n16130
g15875 and n15482_not n15863_not ; n16131
g15876 and n15862_not n16131 ; n16132
g15877 and n16130_not n16132_not ; n16133
g15878 and b[17]_not n16133_not ; n16134
g15879 and n15501_not n15695 ; n16135
g15880 and n15691_not n16135 ; n16136
g15881 and n15692_not n15695_not ; n16137
g15882 and n16136_not n16137_not ; n16138
g15883 and quotient[17] n16138_not ; n16139
g15884 and n15491_not n15863_not ; n16140
g15885 and n15862_not n16140 ; n16141
g15886 and n16139_not n16141_not ; n16142
g15887 and b[16]_not n16142_not ; n16143
g15888 and n15510_not n15690 ; n16144
g15889 and n15686_not n16144 ; n16145
g15890 and n15687_not n15690_not ; n16146
g15891 and n16145_not n16146_not ; n16147
g15892 and quotient[17] n16147_not ; n16148
g15893 and n15500_not n15863_not ; n16149
g15894 and n15862_not n16149 ; n16150
g15895 and n16148_not n16150_not ; n16151
g15896 and b[15]_not n16151_not ; n16152
g15897 and n15519_not n15685 ; n16153
g15898 and n15681_not n16153 ; n16154
g15899 and n15682_not n15685_not ; n16155
g15900 and n16154_not n16155_not ; n16156
g15901 and quotient[17] n16156_not ; n16157
g15902 and n15509_not n15863_not ; n16158
g15903 and n15862_not n16158 ; n16159
g15904 and n16157_not n16159_not ; n16160
g15905 and b[14]_not n16160_not ; n16161
g15906 and n15528_not n15680 ; n16162
g15907 and n15676_not n16162 ; n16163
g15908 and n15677_not n15680_not ; n16164
g15909 and n16163_not n16164_not ; n16165
g15910 and quotient[17] n16165_not ; n16166
g15911 and n15518_not n15863_not ; n16167
g15912 and n15862_not n16167 ; n16168
g15913 and n16166_not n16168_not ; n16169
g15914 and b[13]_not n16169_not ; n16170
g15915 and n15537_not n15675 ; n16171
g15916 and n15671_not n16171 ; n16172
g15917 and n15672_not n15675_not ; n16173
g15918 and n16172_not n16173_not ; n16174
g15919 and quotient[17] n16174_not ; n16175
g15920 and n15527_not n15863_not ; n16176
g15921 and n15862_not n16176 ; n16177
g15922 and n16175_not n16177_not ; n16178
g15923 and b[12]_not n16178_not ; n16179
g15924 and n15546_not n15670 ; n16180
g15925 and n15666_not n16180 ; n16181
g15926 and n15667_not n15670_not ; n16182
g15927 and n16181_not n16182_not ; n16183
g15928 and quotient[17] n16183_not ; n16184
g15929 and n15536_not n15863_not ; n16185
g15930 and n15862_not n16185 ; n16186
g15931 and n16184_not n16186_not ; n16187
g15932 and b[11]_not n16187_not ; n16188
g15933 and n15555_not n15665 ; n16189
g15934 and n15661_not n16189 ; n16190
g15935 and n15662_not n15665_not ; n16191
g15936 and n16190_not n16191_not ; n16192
g15937 and quotient[17] n16192_not ; n16193
g15938 and n15545_not n15863_not ; n16194
g15939 and n15862_not n16194 ; n16195
g15940 and n16193_not n16195_not ; n16196
g15941 and b[10]_not n16196_not ; n16197
g15942 and n15564_not n15660 ; n16198
g15943 and n15656_not n16198 ; n16199
g15944 and n15657_not n15660_not ; n16200
g15945 and n16199_not n16200_not ; n16201
g15946 and quotient[17] n16201_not ; n16202
g15947 and n15554_not n15863_not ; n16203
g15948 and n15862_not n16203 ; n16204
g15949 and n16202_not n16204_not ; n16205
g15950 and b[9]_not n16205_not ; n16206
g15951 and n15573_not n15655 ; n16207
g15952 and n15651_not n16207 ; n16208
g15953 and n15652_not n15655_not ; n16209
g15954 and n16208_not n16209_not ; n16210
g15955 and quotient[17] n16210_not ; n16211
g15956 and n15563_not n15863_not ; n16212
g15957 and n15862_not n16212 ; n16213
g15958 and n16211_not n16213_not ; n16214
g15959 and b[8]_not n16214_not ; n16215
g15960 and n15582_not n15650 ; n16216
g15961 and n15646_not n16216 ; n16217
g15962 and n15647_not n15650_not ; n16218
g15963 and n16217_not n16218_not ; n16219
g15964 and quotient[17] n16219_not ; n16220
g15965 and n15572_not n15863_not ; n16221
g15966 and n15862_not n16221 ; n16222
g15967 and n16220_not n16222_not ; n16223
g15968 and b[7]_not n16223_not ; n16224
g15969 and n15591_not n15645 ; n16225
g15970 and n15641_not n16225 ; n16226
g15971 and n15642_not n15645_not ; n16227
g15972 and n16226_not n16227_not ; n16228
g15973 and quotient[17] n16228_not ; n16229
g15974 and n15581_not n15863_not ; n16230
g15975 and n15862_not n16230 ; n16231
g15976 and n16229_not n16231_not ; n16232
g15977 and b[6]_not n16232_not ; n16233
g15978 and n15600_not n15640 ; n16234
g15979 and n15636_not n16234 ; n16235
g15980 and n15637_not n15640_not ; n16236
g15981 and n16235_not n16236_not ; n16237
g15982 and quotient[17] n16237_not ; n16238
g15983 and n15590_not n15863_not ; n16239
g15984 and n15862_not n16239 ; n16240
g15985 and n16238_not n16240_not ; n16241
g15986 and b[5]_not n16241_not ; n16242
g15987 and n15608_not n15635 ; n16243
g15988 and n15631_not n16243 ; n16244
g15989 and n15632_not n15635_not ; n16245
g15990 and n16244_not n16245_not ; n16246
g15991 and quotient[17] n16246_not ; n16247
g15992 and n15599_not n15863_not ; n16248
g15993 and n15862_not n16248 ; n16249
g15994 and n16247_not n16249_not ; n16250
g15995 and b[4]_not n16250_not ; n16251
g15996 and n15626_not n15630 ; n16252
g15997 and n15625_not n16252 ; n16253
g15998 and n15627_not n15630_not ; n16254
g15999 and n16253_not n16254_not ; n16255
g16000 and quotient[17] n16255_not ; n16256
g16001 and n15607_not n15863_not ; n16257
g16002 and n15862_not n16257 ; n16258
g16003 and n16256_not n16258_not ; n16259
g16004 and b[3]_not n16259_not ; n16260
g16005 and n15622_not n15624 ; n16261
g16006 and n15620_not n16261 ; n16262
g16007 and n15625_not n16262_not ; n16263
g16008 and quotient[17] n16263 ; n16264
g16009 and n15619_not n15863_not ; n16265
g16010 and n15862_not n16265 ; n16266
g16011 and n16264_not n16266_not ; n16267
g16012 and b[2]_not n16267_not ; n16268
g16013 and b[0] quotient[17] ; n16269
g16014 and a[17] n16269_not ; n16270
g16015 and n15624 quotient[17] ; n16271
g16016 and n16270_not n16271_not ; n16272
g16017 and b[1] n16272_not ; n16273
g16018 and b[1]_not n16271_not ; n16274
g16019 and n16270_not n16274 ; n16275
g16020 and n16273_not n16275_not ; n16276
g16021 and a[16]_not b[0] ; n16277
g16022 and n16276_not n16277_not ; n16278
g16023 and b[1]_not n16272_not ; n16279
g16024 and n16278_not n16279_not ; n16280
g16025 and b[2] n16266_not ; n16281
g16026 and n16264_not n16281 ; n16282
g16027 and n16268_not n16282_not ; n16283
g16028 and n16280_not n16283 ; n16284
g16029 and n16268_not n16284_not ; n16285
g16030 and b[3] n16258_not ; n16286
g16031 and n16256_not n16286 ; n16287
g16032 and n16260_not n16287_not ; n16288
g16033 and n16285_not n16288 ; n16289
g16034 and n16260_not n16289_not ; n16290
g16035 and b[4] n16249_not ; n16291
g16036 and n16247_not n16291 ; n16292
g16037 and n16251_not n16292_not ; n16293
g16038 and n16290_not n16293 ; n16294
g16039 and n16251_not n16294_not ; n16295
g16040 and b[5] n16240_not ; n16296
g16041 and n16238_not n16296 ; n16297
g16042 and n16242_not n16297_not ; n16298
g16043 and n16295_not n16298 ; n16299
g16044 and n16242_not n16299_not ; n16300
g16045 and b[6] n16231_not ; n16301
g16046 and n16229_not n16301 ; n16302
g16047 and n16233_not n16302_not ; n16303
g16048 and n16300_not n16303 ; n16304
g16049 and n16233_not n16304_not ; n16305
g16050 and b[7] n16222_not ; n16306
g16051 and n16220_not n16306 ; n16307
g16052 and n16224_not n16307_not ; n16308
g16053 and n16305_not n16308 ; n16309
g16054 and n16224_not n16309_not ; n16310
g16055 and b[8] n16213_not ; n16311
g16056 and n16211_not n16311 ; n16312
g16057 and n16215_not n16312_not ; n16313
g16058 and n16310_not n16313 ; n16314
g16059 and n16215_not n16314_not ; n16315
g16060 and b[9] n16204_not ; n16316
g16061 and n16202_not n16316 ; n16317
g16062 and n16206_not n16317_not ; n16318
g16063 and n16315_not n16318 ; n16319
g16064 and n16206_not n16319_not ; n16320
g16065 and b[10] n16195_not ; n16321
g16066 and n16193_not n16321 ; n16322
g16067 and n16197_not n16322_not ; n16323
g16068 and n16320_not n16323 ; n16324
g16069 and n16197_not n16324_not ; n16325
g16070 and b[11] n16186_not ; n16326
g16071 and n16184_not n16326 ; n16327
g16072 and n16188_not n16327_not ; n16328
g16073 and n16325_not n16328 ; n16329
g16074 and n16188_not n16329_not ; n16330
g16075 and b[12] n16177_not ; n16331
g16076 and n16175_not n16331 ; n16332
g16077 and n16179_not n16332_not ; n16333
g16078 and n16330_not n16333 ; n16334
g16079 and n16179_not n16334_not ; n16335
g16080 and b[13] n16168_not ; n16336
g16081 and n16166_not n16336 ; n16337
g16082 and n16170_not n16337_not ; n16338
g16083 and n16335_not n16338 ; n16339
g16084 and n16170_not n16339_not ; n16340
g16085 and b[14] n16159_not ; n16341
g16086 and n16157_not n16341 ; n16342
g16087 and n16161_not n16342_not ; n16343
g16088 and n16340_not n16343 ; n16344
g16089 and n16161_not n16344_not ; n16345
g16090 and b[15] n16150_not ; n16346
g16091 and n16148_not n16346 ; n16347
g16092 and n16152_not n16347_not ; n16348
g16093 and n16345_not n16348 ; n16349
g16094 and n16152_not n16349_not ; n16350
g16095 and b[16] n16141_not ; n16351
g16096 and n16139_not n16351 ; n16352
g16097 and n16143_not n16352_not ; n16353
g16098 and n16350_not n16353 ; n16354
g16099 and n16143_not n16354_not ; n16355
g16100 and b[17] n16132_not ; n16356
g16101 and n16130_not n16356 ; n16357
g16102 and n16134_not n16357_not ; n16358
g16103 and n16355_not n16358 ; n16359
g16104 and n16134_not n16359_not ; n16360
g16105 and b[18] n16123_not ; n16361
g16106 and n16121_not n16361 ; n16362
g16107 and n16125_not n16362_not ; n16363
g16108 and n16360_not n16363 ; n16364
g16109 and n16125_not n16364_not ; n16365
g16110 and b[19] n16114_not ; n16366
g16111 and n16112_not n16366 ; n16367
g16112 and n16116_not n16367_not ; n16368
g16113 and n16365_not n16368 ; n16369
g16114 and n16116_not n16369_not ; n16370
g16115 and b[20] n16105_not ; n16371
g16116 and n16103_not n16371 ; n16372
g16117 and n16107_not n16372_not ; n16373
g16118 and n16370_not n16373 ; n16374
g16119 and n16107_not n16374_not ; n16375
g16120 and b[21] n16096_not ; n16376
g16121 and n16094_not n16376 ; n16377
g16122 and n16098_not n16377_not ; n16378
g16123 and n16375_not n16378 ; n16379
g16124 and n16098_not n16379_not ; n16380
g16125 and b[22] n16087_not ; n16381
g16126 and n16085_not n16381 ; n16382
g16127 and n16089_not n16382_not ; n16383
g16128 and n16380_not n16383 ; n16384
g16129 and n16089_not n16384_not ; n16385
g16130 and b[23] n16078_not ; n16386
g16131 and n16076_not n16386 ; n16387
g16132 and n16080_not n16387_not ; n16388
g16133 and n16385_not n16388 ; n16389
g16134 and n16080_not n16389_not ; n16390
g16135 and b[24] n16069_not ; n16391
g16136 and n16067_not n16391 ; n16392
g16137 and n16071_not n16392_not ; n16393
g16138 and n16390_not n16393 ; n16394
g16139 and n16071_not n16394_not ; n16395
g16140 and b[25] n16060_not ; n16396
g16141 and n16058_not n16396 ; n16397
g16142 and n16062_not n16397_not ; n16398
g16143 and n16395_not n16398 ; n16399
g16144 and n16062_not n16399_not ; n16400
g16145 and b[26] n16051_not ; n16401
g16146 and n16049_not n16401 ; n16402
g16147 and n16053_not n16402_not ; n16403
g16148 and n16400_not n16403 ; n16404
g16149 and n16053_not n16404_not ; n16405
g16150 and b[27] n16042_not ; n16406
g16151 and n16040_not n16406 ; n16407
g16152 and n16044_not n16407_not ; n16408
g16153 and n16405_not n16408 ; n16409
g16154 and n16044_not n16409_not ; n16410
g16155 and b[28] n16033_not ; n16411
g16156 and n16031_not n16411 ; n16412
g16157 and n16035_not n16412_not ; n16413
g16158 and n16410_not n16413 ; n16414
g16159 and n16035_not n16414_not ; n16415
g16160 and b[29] n16024_not ; n16416
g16161 and n16022_not n16416 ; n16417
g16162 and n16026_not n16417_not ; n16418
g16163 and n16415_not n16418 ; n16419
g16164 and n16026_not n16419_not ; n16420
g16165 and b[30] n16015_not ; n16421
g16166 and n16013_not n16421 ; n16422
g16167 and n16017_not n16422_not ; n16423
g16168 and n16420_not n16423 ; n16424
g16169 and n16017_not n16424_not ; n16425
g16170 and b[31] n16006_not ; n16426
g16171 and n16004_not n16426 ; n16427
g16172 and n16008_not n16427_not ; n16428
g16173 and n16425_not n16428 ; n16429
g16174 and n16008_not n16429_not ; n16430
g16175 and b[32] n15997_not ; n16431
g16176 and n15995_not n16431 ; n16432
g16177 and n15999_not n16432_not ; n16433
g16178 and n16430_not n16433 ; n16434
g16179 and n15999_not n16434_not ; n16435
g16180 and b[33] n15988_not ; n16436
g16181 and n15986_not n16436 ; n16437
g16182 and n15990_not n16437_not ; n16438
g16183 and n16435_not n16438 ; n16439
g16184 and n15990_not n16439_not ; n16440
g16185 and b[34] n15979_not ; n16441
g16186 and n15977_not n16441 ; n16442
g16187 and n15981_not n16442_not ; n16443
g16188 and n16440_not n16443 ; n16444
g16189 and n15981_not n16444_not ; n16445
g16190 and b[35] n15970_not ; n16446
g16191 and n15968_not n16446 ; n16447
g16192 and n15972_not n16447_not ; n16448
g16193 and n16445_not n16448 ; n16449
g16194 and n15972_not n16449_not ; n16450
g16195 and b[36] n15961_not ; n16451
g16196 and n15959_not n16451 ; n16452
g16197 and n15963_not n16452_not ; n16453
g16198 and n16450_not n16453 ; n16454
g16199 and n15963_not n16454_not ; n16455
g16200 and b[37] n15952_not ; n16456
g16201 and n15950_not n16456 ; n16457
g16202 and n15954_not n16457_not ; n16458
g16203 and n16455_not n16458 ; n16459
g16204 and n15954_not n16459_not ; n16460
g16205 and b[38] n15943_not ; n16461
g16206 and n15941_not n16461 ; n16462
g16207 and n15945_not n16462_not ; n16463
g16208 and n16460_not n16463 ; n16464
g16209 and n15945_not n16464_not ; n16465
g16210 and b[39] n15934_not ; n16466
g16211 and n15932_not n16466 ; n16467
g16212 and n15936_not n16467_not ; n16468
g16213 and n16465_not n16468 ; n16469
g16214 and n15936_not n16469_not ; n16470
g16215 and b[40] n15925_not ; n16471
g16216 and n15923_not n16471 ; n16472
g16217 and n15927_not n16472_not ; n16473
g16218 and n16470_not n16473 ; n16474
g16219 and n15927_not n16474_not ; n16475
g16220 and b[41] n15916_not ; n16476
g16221 and n15914_not n16476 ; n16477
g16222 and n15918_not n16477_not ; n16478
g16223 and n16475_not n16478 ; n16479
g16224 and n15918_not n16479_not ; n16480
g16225 and b[42] n15907_not ; n16481
g16226 and n15905_not n16481 ; n16482
g16227 and n15909_not n16482_not ; n16483
g16228 and n16480_not n16483 ; n16484
g16229 and n15909_not n16484_not ; n16485
g16230 and b[43] n15898_not ; n16486
g16231 and n15896_not n16486 ; n16487
g16232 and n15900_not n16487_not ; n16488
g16233 and n16485_not n16488 ; n16489
g16234 and n15900_not n16489_not ; n16490
g16235 and b[44] n15889_not ; n16491
g16236 and n15887_not n16491 ; n16492
g16237 and n15891_not n16492_not ; n16493
g16238 and n16490_not n16493 ; n16494
g16239 and n15891_not n16494_not ; n16495
g16240 and b[45] n15880_not ; n16496
g16241 and n15878_not n16496 ; n16497
g16242 and n15882_not n16497_not ; n16498
g16243 and n16495_not n16498 ; n16499
g16244 and n15882_not n16499_not ; n16500
g16245 and b[46] n15871_not ; n16501
g16246 and n15869_not n16501 ; n16502
g16247 and n15873_not n16502_not ; n16503
g16248 and n16500_not n16503 ; n16504
g16249 and n15873_not n16504_not ; n16505
g16250 and n15222_not n15857_not ; n16506
g16251 and n15855_not n16506 ; n16507
g16252 and n15846_not n16507 ; n16508
g16253 and n15855_not n15857_not ; n16509
g16254 and n15847_not n16509_not ; n16510
g16255 and n16508_not n16510_not ; n16511
g16256 and quotient[17] n16511_not ; n16512
g16257 and n15854_not n15863_not ; n16513
g16258 and n15862_not n16513 ; n16514
g16259 and n16512_not n16514_not ; n16515
g16260 and b[47]_not n16515_not ; n16516
g16261 and b[47] n16514_not ; n16517
g16262 and n16512_not n16517 ; n16518
g16263 and n338 n16518_not ; n16519
g16264 and n16516_not n16519 ; n16520
g16265 and n16505_not n16520 ; n16521
g16266 and n15859 n16515_not ; n16522
g16267 and n16521_not n16522_not ; quotient[16]
g16268 and n15882_not n16503 ; n16524
g16269 and n16499_not n16524 ; n16525
g16270 and n16500_not n16503_not ; n16526
g16271 and n16525_not n16526_not ; n16527
g16272 and quotient[16] n16527_not ; n16528
g16273 and n15872_not n16522_not ; n16529
g16274 and n16521_not n16529 ; n16530
g16275 and n16528_not n16530_not ; n16531
g16276 and n15873_not n16518_not ; n16532
g16277 and n16516_not n16532 ; n16533
g16278 and n16504_not n16533 ; n16534
g16279 and n16516_not n16518_not ; n16535
g16280 and n16505_not n16535_not ; n16536
g16281 and n16534_not n16536_not ; n16537
g16282 and quotient[16] n16537_not ; n16538
g16283 and n16515_not n16522_not ; n16539
g16284 and n16521_not n16539 ; n16540
g16285 and n16538_not n16540_not ; n16541
g16286 and b[48]_not n16541_not ; n16542
g16287 and b[47]_not n16531_not ; n16543
g16288 and n15891_not n16498 ; n16544
g16289 and n16494_not n16544 ; n16545
g16290 and n16495_not n16498_not ; n16546
g16291 and n16545_not n16546_not ; n16547
g16292 and quotient[16] n16547_not ; n16548
g16293 and n15881_not n16522_not ; n16549
g16294 and n16521_not n16549 ; n16550
g16295 and n16548_not n16550_not ; n16551
g16296 and b[46]_not n16551_not ; n16552
g16297 and n15900_not n16493 ; n16553
g16298 and n16489_not n16553 ; n16554
g16299 and n16490_not n16493_not ; n16555
g16300 and n16554_not n16555_not ; n16556
g16301 and quotient[16] n16556_not ; n16557
g16302 and n15890_not n16522_not ; n16558
g16303 and n16521_not n16558 ; n16559
g16304 and n16557_not n16559_not ; n16560
g16305 and b[45]_not n16560_not ; n16561
g16306 and n15909_not n16488 ; n16562
g16307 and n16484_not n16562 ; n16563
g16308 and n16485_not n16488_not ; n16564
g16309 and n16563_not n16564_not ; n16565
g16310 and quotient[16] n16565_not ; n16566
g16311 and n15899_not n16522_not ; n16567
g16312 and n16521_not n16567 ; n16568
g16313 and n16566_not n16568_not ; n16569
g16314 and b[44]_not n16569_not ; n16570
g16315 and n15918_not n16483 ; n16571
g16316 and n16479_not n16571 ; n16572
g16317 and n16480_not n16483_not ; n16573
g16318 and n16572_not n16573_not ; n16574
g16319 and quotient[16] n16574_not ; n16575
g16320 and n15908_not n16522_not ; n16576
g16321 and n16521_not n16576 ; n16577
g16322 and n16575_not n16577_not ; n16578
g16323 and b[43]_not n16578_not ; n16579
g16324 and n15927_not n16478 ; n16580
g16325 and n16474_not n16580 ; n16581
g16326 and n16475_not n16478_not ; n16582
g16327 and n16581_not n16582_not ; n16583
g16328 and quotient[16] n16583_not ; n16584
g16329 and n15917_not n16522_not ; n16585
g16330 and n16521_not n16585 ; n16586
g16331 and n16584_not n16586_not ; n16587
g16332 and b[42]_not n16587_not ; n16588
g16333 and n15936_not n16473 ; n16589
g16334 and n16469_not n16589 ; n16590
g16335 and n16470_not n16473_not ; n16591
g16336 and n16590_not n16591_not ; n16592
g16337 and quotient[16] n16592_not ; n16593
g16338 and n15926_not n16522_not ; n16594
g16339 and n16521_not n16594 ; n16595
g16340 and n16593_not n16595_not ; n16596
g16341 and b[41]_not n16596_not ; n16597
g16342 and n15945_not n16468 ; n16598
g16343 and n16464_not n16598 ; n16599
g16344 and n16465_not n16468_not ; n16600
g16345 and n16599_not n16600_not ; n16601
g16346 and quotient[16] n16601_not ; n16602
g16347 and n15935_not n16522_not ; n16603
g16348 and n16521_not n16603 ; n16604
g16349 and n16602_not n16604_not ; n16605
g16350 and b[40]_not n16605_not ; n16606
g16351 and n15954_not n16463 ; n16607
g16352 and n16459_not n16607 ; n16608
g16353 and n16460_not n16463_not ; n16609
g16354 and n16608_not n16609_not ; n16610
g16355 and quotient[16] n16610_not ; n16611
g16356 and n15944_not n16522_not ; n16612
g16357 and n16521_not n16612 ; n16613
g16358 and n16611_not n16613_not ; n16614
g16359 and b[39]_not n16614_not ; n16615
g16360 and n15963_not n16458 ; n16616
g16361 and n16454_not n16616 ; n16617
g16362 and n16455_not n16458_not ; n16618
g16363 and n16617_not n16618_not ; n16619
g16364 and quotient[16] n16619_not ; n16620
g16365 and n15953_not n16522_not ; n16621
g16366 and n16521_not n16621 ; n16622
g16367 and n16620_not n16622_not ; n16623
g16368 and b[38]_not n16623_not ; n16624
g16369 and n15972_not n16453 ; n16625
g16370 and n16449_not n16625 ; n16626
g16371 and n16450_not n16453_not ; n16627
g16372 and n16626_not n16627_not ; n16628
g16373 and quotient[16] n16628_not ; n16629
g16374 and n15962_not n16522_not ; n16630
g16375 and n16521_not n16630 ; n16631
g16376 and n16629_not n16631_not ; n16632
g16377 and b[37]_not n16632_not ; n16633
g16378 and n15981_not n16448 ; n16634
g16379 and n16444_not n16634 ; n16635
g16380 and n16445_not n16448_not ; n16636
g16381 and n16635_not n16636_not ; n16637
g16382 and quotient[16] n16637_not ; n16638
g16383 and n15971_not n16522_not ; n16639
g16384 and n16521_not n16639 ; n16640
g16385 and n16638_not n16640_not ; n16641
g16386 and b[36]_not n16641_not ; n16642
g16387 and n15990_not n16443 ; n16643
g16388 and n16439_not n16643 ; n16644
g16389 and n16440_not n16443_not ; n16645
g16390 and n16644_not n16645_not ; n16646
g16391 and quotient[16] n16646_not ; n16647
g16392 and n15980_not n16522_not ; n16648
g16393 and n16521_not n16648 ; n16649
g16394 and n16647_not n16649_not ; n16650
g16395 and b[35]_not n16650_not ; n16651
g16396 and n15999_not n16438 ; n16652
g16397 and n16434_not n16652 ; n16653
g16398 and n16435_not n16438_not ; n16654
g16399 and n16653_not n16654_not ; n16655
g16400 and quotient[16] n16655_not ; n16656
g16401 and n15989_not n16522_not ; n16657
g16402 and n16521_not n16657 ; n16658
g16403 and n16656_not n16658_not ; n16659
g16404 and b[34]_not n16659_not ; n16660
g16405 and n16008_not n16433 ; n16661
g16406 and n16429_not n16661 ; n16662
g16407 and n16430_not n16433_not ; n16663
g16408 and n16662_not n16663_not ; n16664
g16409 and quotient[16] n16664_not ; n16665
g16410 and n15998_not n16522_not ; n16666
g16411 and n16521_not n16666 ; n16667
g16412 and n16665_not n16667_not ; n16668
g16413 and b[33]_not n16668_not ; n16669
g16414 and n16017_not n16428 ; n16670
g16415 and n16424_not n16670 ; n16671
g16416 and n16425_not n16428_not ; n16672
g16417 and n16671_not n16672_not ; n16673
g16418 and quotient[16] n16673_not ; n16674
g16419 and n16007_not n16522_not ; n16675
g16420 and n16521_not n16675 ; n16676
g16421 and n16674_not n16676_not ; n16677
g16422 and b[32]_not n16677_not ; n16678
g16423 and n16026_not n16423 ; n16679
g16424 and n16419_not n16679 ; n16680
g16425 and n16420_not n16423_not ; n16681
g16426 and n16680_not n16681_not ; n16682
g16427 and quotient[16] n16682_not ; n16683
g16428 and n16016_not n16522_not ; n16684
g16429 and n16521_not n16684 ; n16685
g16430 and n16683_not n16685_not ; n16686
g16431 and b[31]_not n16686_not ; n16687
g16432 and n16035_not n16418 ; n16688
g16433 and n16414_not n16688 ; n16689
g16434 and n16415_not n16418_not ; n16690
g16435 and n16689_not n16690_not ; n16691
g16436 and quotient[16] n16691_not ; n16692
g16437 and n16025_not n16522_not ; n16693
g16438 and n16521_not n16693 ; n16694
g16439 and n16692_not n16694_not ; n16695
g16440 and b[30]_not n16695_not ; n16696
g16441 and n16044_not n16413 ; n16697
g16442 and n16409_not n16697 ; n16698
g16443 and n16410_not n16413_not ; n16699
g16444 and n16698_not n16699_not ; n16700
g16445 and quotient[16] n16700_not ; n16701
g16446 and n16034_not n16522_not ; n16702
g16447 and n16521_not n16702 ; n16703
g16448 and n16701_not n16703_not ; n16704
g16449 and b[29]_not n16704_not ; n16705
g16450 and n16053_not n16408 ; n16706
g16451 and n16404_not n16706 ; n16707
g16452 and n16405_not n16408_not ; n16708
g16453 and n16707_not n16708_not ; n16709
g16454 and quotient[16] n16709_not ; n16710
g16455 and n16043_not n16522_not ; n16711
g16456 and n16521_not n16711 ; n16712
g16457 and n16710_not n16712_not ; n16713
g16458 and b[28]_not n16713_not ; n16714
g16459 and n16062_not n16403 ; n16715
g16460 and n16399_not n16715 ; n16716
g16461 and n16400_not n16403_not ; n16717
g16462 and n16716_not n16717_not ; n16718
g16463 and quotient[16] n16718_not ; n16719
g16464 and n16052_not n16522_not ; n16720
g16465 and n16521_not n16720 ; n16721
g16466 and n16719_not n16721_not ; n16722
g16467 and b[27]_not n16722_not ; n16723
g16468 and n16071_not n16398 ; n16724
g16469 and n16394_not n16724 ; n16725
g16470 and n16395_not n16398_not ; n16726
g16471 and n16725_not n16726_not ; n16727
g16472 and quotient[16] n16727_not ; n16728
g16473 and n16061_not n16522_not ; n16729
g16474 and n16521_not n16729 ; n16730
g16475 and n16728_not n16730_not ; n16731
g16476 and b[26]_not n16731_not ; n16732
g16477 and n16080_not n16393 ; n16733
g16478 and n16389_not n16733 ; n16734
g16479 and n16390_not n16393_not ; n16735
g16480 and n16734_not n16735_not ; n16736
g16481 and quotient[16] n16736_not ; n16737
g16482 and n16070_not n16522_not ; n16738
g16483 and n16521_not n16738 ; n16739
g16484 and n16737_not n16739_not ; n16740
g16485 and b[25]_not n16740_not ; n16741
g16486 and n16089_not n16388 ; n16742
g16487 and n16384_not n16742 ; n16743
g16488 and n16385_not n16388_not ; n16744
g16489 and n16743_not n16744_not ; n16745
g16490 and quotient[16] n16745_not ; n16746
g16491 and n16079_not n16522_not ; n16747
g16492 and n16521_not n16747 ; n16748
g16493 and n16746_not n16748_not ; n16749
g16494 and b[24]_not n16749_not ; n16750
g16495 and n16098_not n16383 ; n16751
g16496 and n16379_not n16751 ; n16752
g16497 and n16380_not n16383_not ; n16753
g16498 and n16752_not n16753_not ; n16754
g16499 and quotient[16] n16754_not ; n16755
g16500 and n16088_not n16522_not ; n16756
g16501 and n16521_not n16756 ; n16757
g16502 and n16755_not n16757_not ; n16758
g16503 and b[23]_not n16758_not ; n16759
g16504 and n16107_not n16378 ; n16760
g16505 and n16374_not n16760 ; n16761
g16506 and n16375_not n16378_not ; n16762
g16507 and n16761_not n16762_not ; n16763
g16508 and quotient[16] n16763_not ; n16764
g16509 and n16097_not n16522_not ; n16765
g16510 and n16521_not n16765 ; n16766
g16511 and n16764_not n16766_not ; n16767
g16512 and b[22]_not n16767_not ; n16768
g16513 and n16116_not n16373 ; n16769
g16514 and n16369_not n16769 ; n16770
g16515 and n16370_not n16373_not ; n16771
g16516 and n16770_not n16771_not ; n16772
g16517 and quotient[16] n16772_not ; n16773
g16518 and n16106_not n16522_not ; n16774
g16519 and n16521_not n16774 ; n16775
g16520 and n16773_not n16775_not ; n16776
g16521 and b[21]_not n16776_not ; n16777
g16522 and n16125_not n16368 ; n16778
g16523 and n16364_not n16778 ; n16779
g16524 and n16365_not n16368_not ; n16780
g16525 and n16779_not n16780_not ; n16781
g16526 and quotient[16] n16781_not ; n16782
g16527 and n16115_not n16522_not ; n16783
g16528 and n16521_not n16783 ; n16784
g16529 and n16782_not n16784_not ; n16785
g16530 and b[20]_not n16785_not ; n16786
g16531 and n16134_not n16363 ; n16787
g16532 and n16359_not n16787 ; n16788
g16533 and n16360_not n16363_not ; n16789
g16534 and n16788_not n16789_not ; n16790
g16535 and quotient[16] n16790_not ; n16791
g16536 and n16124_not n16522_not ; n16792
g16537 and n16521_not n16792 ; n16793
g16538 and n16791_not n16793_not ; n16794
g16539 and b[19]_not n16794_not ; n16795
g16540 and n16143_not n16358 ; n16796
g16541 and n16354_not n16796 ; n16797
g16542 and n16355_not n16358_not ; n16798
g16543 and n16797_not n16798_not ; n16799
g16544 and quotient[16] n16799_not ; n16800
g16545 and n16133_not n16522_not ; n16801
g16546 and n16521_not n16801 ; n16802
g16547 and n16800_not n16802_not ; n16803
g16548 and b[18]_not n16803_not ; n16804
g16549 and n16152_not n16353 ; n16805
g16550 and n16349_not n16805 ; n16806
g16551 and n16350_not n16353_not ; n16807
g16552 and n16806_not n16807_not ; n16808
g16553 and quotient[16] n16808_not ; n16809
g16554 and n16142_not n16522_not ; n16810
g16555 and n16521_not n16810 ; n16811
g16556 and n16809_not n16811_not ; n16812
g16557 and b[17]_not n16812_not ; n16813
g16558 and n16161_not n16348 ; n16814
g16559 and n16344_not n16814 ; n16815
g16560 and n16345_not n16348_not ; n16816
g16561 and n16815_not n16816_not ; n16817
g16562 and quotient[16] n16817_not ; n16818
g16563 and n16151_not n16522_not ; n16819
g16564 and n16521_not n16819 ; n16820
g16565 and n16818_not n16820_not ; n16821
g16566 and b[16]_not n16821_not ; n16822
g16567 and n16170_not n16343 ; n16823
g16568 and n16339_not n16823 ; n16824
g16569 and n16340_not n16343_not ; n16825
g16570 and n16824_not n16825_not ; n16826
g16571 and quotient[16] n16826_not ; n16827
g16572 and n16160_not n16522_not ; n16828
g16573 and n16521_not n16828 ; n16829
g16574 and n16827_not n16829_not ; n16830
g16575 and b[15]_not n16830_not ; n16831
g16576 and n16179_not n16338 ; n16832
g16577 and n16334_not n16832 ; n16833
g16578 and n16335_not n16338_not ; n16834
g16579 and n16833_not n16834_not ; n16835
g16580 and quotient[16] n16835_not ; n16836
g16581 and n16169_not n16522_not ; n16837
g16582 and n16521_not n16837 ; n16838
g16583 and n16836_not n16838_not ; n16839
g16584 and b[14]_not n16839_not ; n16840
g16585 and n16188_not n16333 ; n16841
g16586 and n16329_not n16841 ; n16842
g16587 and n16330_not n16333_not ; n16843
g16588 and n16842_not n16843_not ; n16844
g16589 and quotient[16] n16844_not ; n16845
g16590 and n16178_not n16522_not ; n16846
g16591 and n16521_not n16846 ; n16847
g16592 and n16845_not n16847_not ; n16848
g16593 and b[13]_not n16848_not ; n16849
g16594 and n16197_not n16328 ; n16850
g16595 and n16324_not n16850 ; n16851
g16596 and n16325_not n16328_not ; n16852
g16597 and n16851_not n16852_not ; n16853
g16598 and quotient[16] n16853_not ; n16854
g16599 and n16187_not n16522_not ; n16855
g16600 and n16521_not n16855 ; n16856
g16601 and n16854_not n16856_not ; n16857
g16602 and b[12]_not n16857_not ; n16858
g16603 and n16206_not n16323 ; n16859
g16604 and n16319_not n16859 ; n16860
g16605 and n16320_not n16323_not ; n16861
g16606 and n16860_not n16861_not ; n16862
g16607 and quotient[16] n16862_not ; n16863
g16608 and n16196_not n16522_not ; n16864
g16609 and n16521_not n16864 ; n16865
g16610 and n16863_not n16865_not ; n16866
g16611 and b[11]_not n16866_not ; n16867
g16612 and n16215_not n16318 ; n16868
g16613 and n16314_not n16868 ; n16869
g16614 and n16315_not n16318_not ; n16870
g16615 and n16869_not n16870_not ; n16871
g16616 and quotient[16] n16871_not ; n16872
g16617 and n16205_not n16522_not ; n16873
g16618 and n16521_not n16873 ; n16874
g16619 and n16872_not n16874_not ; n16875
g16620 and b[10]_not n16875_not ; n16876
g16621 and n16224_not n16313 ; n16877
g16622 and n16309_not n16877 ; n16878
g16623 and n16310_not n16313_not ; n16879
g16624 and n16878_not n16879_not ; n16880
g16625 and quotient[16] n16880_not ; n16881
g16626 and n16214_not n16522_not ; n16882
g16627 and n16521_not n16882 ; n16883
g16628 and n16881_not n16883_not ; n16884
g16629 and b[9]_not n16884_not ; n16885
g16630 and n16233_not n16308 ; n16886
g16631 and n16304_not n16886 ; n16887
g16632 and n16305_not n16308_not ; n16888
g16633 and n16887_not n16888_not ; n16889
g16634 and quotient[16] n16889_not ; n16890
g16635 and n16223_not n16522_not ; n16891
g16636 and n16521_not n16891 ; n16892
g16637 and n16890_not n16892_not ; n16893
g16638 and b[8]_not n16893_not ; n16894
g16639 and n16242_not n16303 ; n16895
g16640 and n16299_not n16895 ; n16896
g16641 and n16300_not n16303_not ; n16897
g16642 and n16896_not n16897_not ; n16898
g16643 and quotient[16] n16898_not ; n16899
g16644 and n16232_not n16522_not ; n16900
g16645 and n16521_not n16900 ; n16901
g16646 and n16899_not n16901_not ; n16902
g16647 and b[7]_not n16902_not ; n16903
g16648 and n16251_not n16298 ; n16904
g16649 and n16294_not n16904 ; n16905
g16650 and n16295_not n16298_not ; n16906
g16651 and n16905_not n16906_not ; n16907
g16652 and quotient[16] n16907_not ; n16908
g16653 and n16241_not n16522_not ; n16909
g16654 and n16521_not n16909 ; n16910
g16655 and n16908_not n16910_not ; n16911
g16656 and b[6]_not n16911_not ; n16912
g16657 and n16260_not n16293 ; n16913
g16658 and n16289_not n16913 ; n16914
g16659 and n16290_not n16293_not ; n16915
g16660 and n16914_not n16915_not ; n16916
g16661 and quotient[16] n16916_not ; n16917
g16662 and n16250_not n16522_not ; n16918
g16663 and n16521_not n16918 ; n16919
g16664 and n16917_not n16919_not ; n16920
g16665 and b[5]_not n16920_not ; n16921
g16666 and n16268_not n16288 ; n16922
g16667 and n16284_not n16922 ; n16923
g16668 and n16285_not n16288_not ; n16924
g16669 and n16923_not n16924_not ; n16925
g16670 and quotient[16] n16925_not ; n16926
g16671 and n16259_not n16522_not ; n16927
g16672 and n16521_not n16927 ; n16928
g16673 and n16926_not n16928_not ; n16929
g16674 and b[4]_not n16929_not ; n16930
g16675 and n16279_not n16283 ; n16931
g16676 and n16278_not n16931 ; n16932
g16677 and n16280_not n16283_not ; n16933
g16678 and n16932_not n16933_not ; n16934
g16679 and quotient[16] n16934_not ; n16935
g16680 and n16267_not n16522_not ; n16936
g16681 and n16521_not n16936 ; n16937
g16682 and n16935_not n16937_not ; n16938
g16683 and b[3]_not n16938_not ; n16939
g16684 and n16275_not n16277 ; n16940
g16685 and n16273_not n16940 ; n16941
g16686 and n16278_not n16941_not ; n16942
g16687 and quotient[16] n16942 ; n16943
g16688 and n16272_not n16522_not ; n16944
g16689 and n16521_not n16944 ; n16945
g16690 and n16943_not n16945_not ; n16946
g16691 and b[2]_not n16946_not ; n16947
g16692 and b[0] quotient[16] ; n16948
g16693 and a[16] n16948_not ; n16949
g16694 and n16277 quotient[16] ; n16950
g16695 and n16949_not n16950_not ; n16951
g16696 and b[1] n16951_not ; n16952
g16697 and b[1]_not n16950_not ; n16953
g16698 and n16949_not n16953 ; n16954
g16699 and n16952_not n16954_not ; n16955
g16700 and a[15]_not b[0] ; n16956
g16701 and n16955_not n16956_not ; n16957
g16702 and b[1]_not n16951_not ; n16958
g16703 and n16957_not n16958_not ; n16959
g16704 and b[2] n16945_not ; n16960
g16705 and n16943_not n16960 ; n16961
g16706 and n16947_not n16961_not ; n16962
g16707 and n16959_not n16962 ; n16963
g16708 and n16947_not n16963_not ; n16964
g16709 and b[3] n16937_not ; n16965
g16710 and n16935_not n16965 ; n16966
g16711 and n16939_not n16966_not ; n16967
g16712 and n16964_not n16967 ; n16968
g16713 and n16939_not n16968_not ; n16969
g16714 and b[4] n16928_not ; n16970
g16715 and n16926_not n16970 ; n16971
g16716 and n16930_not n16971_not ; n16972
g16717 and n16969_not n16972 ; n16973
g16718 and n16930_not n16973_not ; n16974
g16719 and b[5] n16919_not ; n16975
g16720 and n16917_not n16975 ; n16976
g16721 and n16921_not n16976_not ; n16977
g16722 and n16974_not n16977 ; n16978
g16723 and n16921_not n16978_not ; n16979
g16724 and b[6] n16910_not ; n16980
g16725 and n16908_not n16980 ; n16981
g16726 and n16912_not n16981_not ; n16982
g16727 and n16979_not n16982 ; n16983
g16728 and n16912_not n16983_not ; n16984
g16729 and b[7] n16901_not ; n16985
g16730 and n16899_not n16985 ; n16986
g16731 and n16903_not n16986_not ; n16987
g16732 and n16984_not n16987 ; n16988
g16733 and n16903_not n16988_not ; n16989
g16734 and b[8] n16892_not ; n16990
g16735 and n16890_not n16990 ; n16991
g16736 and n16894_not n16991_not ; n16992
g16737 and n16989_not n16992 ; n16993
g16738 and n16894_not n16993_not ; n16994
g16739 and b[9] n16883_not ; n16995
g16740 and n16881_not n16995 ; n16996
g16741 and n16885_not n16996_not ; n16997
g16742 and n16994_not n16997 ; n16998
g16743 and n16885_not n16998_not ; n16999
g16744 and b[10] n16874_not ; n17000
g16745 and n16872_not n17000 ; n17001
g16746 and n16876_not n17001_not ; n17002
g16747 and n16999_not n17002 ; n17003
g16748 and n16876_not n17003_not ; n17004
g16749 and b[11] n16865_not ; n17005
g16750 and n16863_not n17005 ; n17006
g16751 and n16867_not n17006_not ; n17007
g16752 and n17004_not n17007 ; n17008
g16753 and n16867_not n17008_not ; n17009
g16754 and b[12] n16856_not ; n17010
g16755 and n16854_not n17010 ; n17011
g16756 and n16858_not n17011_not ; n17012
g16757 and n17009_not n17012 ; n17013
g16758 and n16858_not n17013_not ; n17014
g16759 and b[13] n16847_not ; n17015
g16760 and n16845_not n17015 ; n17016
g16761 and n16849_not n17016_not ; n17017
g16762 and n17014_not n17017 ; n17018
g16763 and n16849_not n17018_not ; n17019
g16764 and b[14] n16838_not ; n17020
g16765 and n16836_not n17020 ; n17021
g16766 and n16840_not n17021_not ; n17022
g16767 and n17019_not n17022 ; n17023
g16768 and n16840_not n17023_not ; n17024
g16769 and b[15] n16829_not ; n17025
g16770 and n16827_not n17025 ; n17026
g16771 and n16831_not n17026_not ; n17027
g16772 and n17024_not n17027 ; n17028
g16773 and n16831_not n17028_not ; n17029
g16774 and b[16] n16820_not ; n17030
g16775 and n16818_not n17030 ; n17031
g16776 and n16822_not n17031_not ; n17032
g16777 and n17029_not n17032 ; n17033
g16778 and n16822_not n17033_not ; n17034
g16779 and b[17] n16811_not ; n17035
g16780 and n16809_not n17035 ; n17036
g16781 and n16813_not n17036_not ; n17037
g16782 and n17034_not n17037 ; n17038
g16783 and n16813_not n17038_not ; n17039
g16784 and b[18] n16802_not ; n17040
g16785 and n16800_not n17040 ; n17041
g16786 and n16804_not n17041_not ; n17042
g16787 and n17039_not n17042 ; n17043
g16788 and n16804_not n17043_not ; n17044
g16789 and b[19] n16793_not ; n17045
g16790 and n16791_not n17045 ; n17046
g16791 and n16795_not n17046_not ; n17047
g16792 and n17044_not n17047 ; n17048
g16793 and n16795_not n17048_not ; n17049
g16794 and b[20] n16784_not ; n17050
g16795 and n16782_not n17050 ; n17051
g16796 and n16786_not n17051_not ; n17052
g16797 and n17049_not n17052 ; n17053
g16798 and n16786_not n17053_not ; n17054
g16799 and b[21] n16775_not ; n17055
g16800 and n16773_not n17055 ; n17056
g16801 and n16777_not n17056_not ; n17057
g16802 and n17054_not n17057 ; n17058
g16803 and n16777_not n17058_not ; n17059
g16804 and b[22] n16766_not ; n17060
g16805 and n16764_not n17060 ; n17061
g16806 and n16768_not n17061_not ; n17062
g16807 and n17059_not n17062 ; n17063
g16808 and n16768_not n17063_not ; n17064
g16809 and b[23] n16757_not ; n17065
g16810 and n16755_not n17065 ; n17066
g16811 and n16759_not n17066_not ; n17067
g16812 and n17064_not n17067 ; n17068
g16813 and n16759_not n17068_not ; n17069
g16814 and b[24] n16748_not ; n17070
g16815 and n16746_not n17070 ; n17071
g16816 and n16750_not n17071_not ; n17072
g16817 and n17069_not n17072 ; n17073
g16818 and n16750_not n17073_not ; n17074
g16819 and b[25] n16739_not ; n17075
g16820 and n16737_not n17075 ; n17076
g16821 and n16741_not n17076_not ; n17077
g16822 and n17074_not n17077 ; n17078
g16823 and n16741_not n17078_not ; n17079
g16824 and b[26] n16730_not ; n17080
g16825 and n16728_not n17080 ; n17081
g16826 and n16732_not n17081_not ; n17082
g16827 and n17079_not n17082 ; n17083
g16828 and n16732_not n17083_not ; n17084
g16829 and b[27] n16721_not ; n17085
g16830 and n16719_not n17085 ; n17086
g16831 and n16723_not n17086_not ; n17087
g16832 and n17084_not n17087 ; n17088
g16833 and n16723_not n17088_not ; n17089
g16834 and b[28] n16712_not ; n17090
g16835 and n16710_not n17090 ; n17091
g16836 and n16714_not n17091_not ; n17092
g16837 and n17089_not n17092 ; n17093
g16838 and n16714_not n17093_not ; n17094
g16839 and b[29] n16703_not ; n17095
g16840 and n16701_not n17095 ; n17096
g16841 and n16705_not n17096_not ; n17097
g16842 and n17094_not n17097 ; n17098
g16843 and n16705_not n17098_not ; n17099
g16844 and b[30] n16694_not ; n17100
g16845 and n16692_not n17100 ; n17101
g16846 and n16696_not n17101_not ; n17102
g16847 and n17099_not n17102 ; n17103
g16848 and n16696_not n17103_not ; n17104
g16849 and b[31] n16685_not ; n17105
g16850 and n16683_not n17105 ; n17106
g16851 and n16687_not n17106_not ; n17107
g16852 and n17104_not n17107 ; n17108
g16853 and n16687_not n17108_not ; n17109
g16854 and b[32] n16676_not ; n17110
g16855 and n16674_not n17110 ; n17111
g16856 and n16678_not n17111_not ; n17112
g16857 and n17109_not n17112 ; n17113
g16858 and n16678_not n17113_not ; n17114
g16859 and b[33] n16667_not ; n17115
g16860 and n16665_not n17115 ; n17116
g16861 and n16669_not n17116_not ; n17117
g16862 and n17114_not n17117 ; n17118
g16863 and n16669_not n17118_not ; n17119
g16864 and b[34] n16658_not ; n17120
g16865 and n16656_not n17120 ; n17121
g16866 and n16660_not n17121_not ; n17122
g16867 and n17119_not n17122 ; n17123
g16868 and n16660_not n17123_not ; n17124
g16869 and b[35] n16649_not ; n17125
g16870 and n16647_not n17125 ; n17126
g16871 and n16651_not n17126_not ; n17127
g16872 and n17124_not n17127 ; n17128
g16873 and n16651_not n17128_not ; n17129
g16874 and b[36] n16640_not ; n17130
g16875 and n16638_not n17130 ; n17131
g16876 and n16642_not n17131_not ; n17132
g16877 and n17129_not n17132 ; n17133
g16878 and n16642_not n17133_not ; n17134
g16879 and b[37] n16631_not ; n17135
g16880 and n16629_not n17135 ; n17136
g16881 and n16633_not n17136_not ; n17137
g16882 and n17134_not n17137 ; n17138
g16883 and n16633_not n17138_not ; n17139
g16884 and b[38] n16622_not ; n17140
g16885 and n16620_not n17140 ; n17141
g16886 and n16624_not n17141_not ; n17142
g16887 and n17139_not n17142 ; n17143
g16888 and n16624_not n17143_not ; n17144
g16889 and b[39] n16613_not ; n17145
g16890 and n16611_not n17145 ; n17146
g16891 and n16615_not n17146_not ; n17147
g16892 and n17144_not n17147 ; n17148
g16893 and n16615_not n17148_not ; n17149
g16894 and b[40] n16604_not ; n17150
g16895 and n16602_not n17150 ; n17151
g16896 and n16606_not n17151_not ; n17152
g16897 and n17149_not n17152 ; n17153
g16898 and n16606_not n17153_not ; n17154
g16899 and b[41] n16595_not ; n17155
g16900 and n16593_not n17155 ; n17156
g16901 and n16597_not n17156_not ; n17157
g16902 and n17154_not n17157 ; n17158
g16903 and n16597_not n17158_not ; n17159
g16904 and b[42] n16586_not ; n17160
g16905 and n16584_not n17160 ; n17161
g16906 and n16588_not n17161_not ; n17162
g16907 and n17159_not n17162 ; n17163
g16908 and n16588_not n17163_not ; n17164
g16909 and b[43] n16577_not ; n17165
g16910 and n16575_not n17165 ; n17166
g16911 and n16579_not n17166_not ; n17167
g16912 and n17164_not n17167 ; n17168
g16913 and n16579_not n17168_not ; n17169
g16914 and b[44] n16568_not ; n17170
g16915 and n16566_not n17170 ; n17171
g16916 and n16570_not n17171_not ; n17172
g16917 and n17169_not n17172 ; n17173
g16918 and n16570_not n17173_not ; n17174
g16919 and b[45] n16559_not ; n17175
g16920 and n16557_not n17175 ; n17176
g16921 and n16561_not n17176_not ; n17177
g16922 and n17174_not n17177 ; n17178
g16923 and n16561_not n17178_not ; n17179
g16924 and b[46] n16550_not ; n17180
g16925 and n16548_not n17180 ; n17181
g16926 and n16552_not n17181_not ; n17182
g16927 and n17179_not n17182 ; n17183
g16928 and n16552_not n17183_not ; n17184
g16929 and b[47] n16530_not ; n17185
g16930 and n16528_not n17185 ; n17186
g16931 and n16543_not n17186_not ; n17187
g16932 and n17184_not n17187 ; n17188
g16933 and n16543_not n17188_not ; n17189
g16934 and b[48] n16540_not ; n17190
g16935 and n16538_not n17190 ; n17191
g16936 and n16542_not n17191_not ; n17192
g16937 and n17189_not n17192 ; n17193
g16938 and n16542_not n17193_not ; n17194
g16939 and n408 n17194_not ; quotient[15]
g16940 and n16531_not quotient[15]_not ; n17196
g16941 and n16552_not n17187 ; n17197
g16942 and n17183_not n17197 ; n17198
g16943 and n17184_not n17187_not ; n17199
g16944 and n17198_not n17199_not ; n17200
g16945 and n408 n17200_not ; n17201
g16946 and n17194_not n17201 ; n17202
g16947 and n17196_not n17202_not ; n17203
g16948 and b[48]_not n17203_not ; n17204
g16949 and n16551_not quotient[15]_not ; n17205
g16950 and n16561_not n17182 ; n17206
g16951 and n17178_not n17206 ; n17207
g16952 and n17179_not n17182_not ; n17208
g16953 and n17207_not n17208_not ; n17209
g16954 and n408 n17209_not ; n17210
g16955 and n17194_not n17210 ; n17211
g16956 and n17205_not n17211_not ; n17212
g16957 and b[47]_not n17212_not ; n17213
g16958 and n16560_not quotient[15]_not ; n17214
g16959 and n16570_not n17177 ; n17215
g16960 and n17173_not n17215 ; n17216
g16961 and n17174_not n17177_not ; n17217
g16962 and n17216_not n17217_not ; n17218
g16963 and n408 n17218_not ; n17219
g16964 and n17194_not n17219 ; n17220
g16965 and n17214_not n17220_not ; n17221
g16966 and b[46]_not n17221_not ; n17222
g16967 and n16569_not quotient[15]_not ; n17223
g16968 and n16579_not n17172 ; n17224
g16969 and n17168_not n17224 ; n17225
g16970 and n17169_not n17172_not ; n17226
g16971 and n17225_not n17226_not ; n17227
g16972 and n408 n17227_not ; n17228
g16973 and n17194_not n17228 ; n17229
g16974 and n17223_not n17229_not ; n17230
g16975 and b[45]_not n17230_not ; n17231
g16976 and n16578_not quotient[15]_not ; n17232
g16977 and n16588_not n17167 ; n17233
g16978 and n17163_not n17233 ; n17234
g16979 and n17164_not n17167_not ; n17235
g16980 and n17234_not n17235_not ; n17236
g16981 and n408 n17236_not ; n17237
g16982 and n17194_not n17237 ; n17238
g16983 and n17232_not n17238_not ; n17239
g16984 and b[44]_not n17239_not ; n17240
g16985 and n16587_not quotient[15]_not ; n17241
g16986 and n16597_not n17162 ; n17242
g16987 and n17158_not n17242 ; n17243
g16988 and n17159_not n17162_not ; n17244
g16989 and n17243_not n17244_not ; n17245
g16990 and n408 n17245_not ; n17246
g16991 and n17194_not n17246 ; n17247
g16992 and n17241_not n17247_not ; n17248
g16993 and b[43]_not n17248_not ; n17249
g16994 and n16596_not quotient[15]_not ; n17250
g16995 and n16606_not n17157 ; n17251
g16996 and n17153_not n17251 ; n17252
g16997 and n17154_not n17157_not ; n17253
g16998 and n17252_not n17253_not ; n17254
g16999 and n408 n17254_not ; n17255
g17000 and n17194_not n17255 ; n17256
g17001 and n17250_not n17256_not ; n17257
g17002 and b[42]_not n17257_not ; n17258
g17003 and n16605_not quotient[15]_not ; n17259
g17004 and n16615_not n17152 ; n17260
g17005 and n17148_not n17260 ; n17261
g17006 and n17149_not n17152_not ; n17262
g17007 and n17261_not n17262_not ; n17263
g17008 and n408 n17263_not ; n17264
g17009 and n17194_not n17264 ; n17265
g17010 and n17259_not n17265_not ; n17266
g17011 and b[41]_not n17266_not ; n17267
g17012 and n16614_not quotient[15]_not ; n17268
g17013 and n16624_not n17147 ; n17269
g17014 and n17143_not n17269 ; n17270
g17015 and n17144_not n17147_not ; n17271
g17016 and n17270_not n17271_not ; n17272
g17017 and n408 n17272_not ; n17273
g17018 and n17194_not n17273 ; n17274
g17019 and n17268_not n17274_not ; n17275
g17020 and b[40]_not n17275_not ; n17276
g17021 and n16623_not quotient[15]_not ; n17277
g17022 and n16633_not n17142 ; n17278
g17023 and n17138_not n17278 ; n17279
g17024 and n17139_not n17142_not ; n17280
g17025 and n17279_not n17280_not ; n17281
g17026 and n408 n17281_not ; n17282
g17027 and n17194_not n17282 ; n17283
g17028 and n17277_not n17283_not ; n17284
g17029 and b[39]_not n17284_not ; n17285
g17030 and n16632_not quotient[15]_not ; n17286
g17031 and n16642_not n17137 ; n17287
g17032 and n17133_not n17287 ; n17288
g17033 and n17134_not n17137_not ; n17289
g17034 and n17288_not n17289_not ; n17290
g17035 and n408 n17290_not ; n17291
g17036 and n17194_not n17291 ; n17292
g17037 and n17286_not n17292_not ; n17293
g17038 and b[38]_not n17293_not ; n17294
g17039 and n16641_not quotient[15]_not ; n17295
g17040 and n16651_not n17132 ; n17296
g17041 and n17128_not n17296 ; n17297
g17042 and n17129_not n17132_not ; n17298
g17043 and n17297_not n17298_not ; n17299
g17044 and n408 n17299_not ; n17300
g17045 and n17194_not n17300 ; n17301
g17046 and n17295_not n17301_not ; n17302
g17047 and b[37]_not n17302_not ; n17303
g17048 and n16650_not quotient[15]_not ; n17304
g17049 and n16660_not n17127 ; n17305
g17050 and n17123_not n17305 ; n17306
g17051 and n17124_not n17127_not ; n17307
g17052 and n17306_not n17307_not ; n17308
g17053 and n408 n17308_not ; n17309
g17054 and n17194_not n17309 ; n17310
g17055 and n17304_not n17310_not ; n17311
g17056 and b[36]_not n17311_not ; n17312
g17057 and n16659_not quotient[15]_not ; n17313
g17058 and n16669_not n17122 ; n17314
g17059 and n17118_not n17314 ; n17315
g17060 and n17119_not n17122_not ; n17316
g17061 and n17315_not n17316_not ; n17317
g17062 and n408 n17317_not ; n17318
g17063 and n17194_not n17318 ; n17319
g17064 and n17313_not n17319_not ; n17320
g17065 and b[35]_not n17320_not ; n17321
g17066 and n16668_not quotient[15]_not ; n17322
g17067 and n16678_not n17117 ; n17323
g17068 and n17113_not n17323 ; n17324
g17069 and n17114_not n17117_not ; n17325
g17070 and n17324_not n17325_not ; n17326
g17071 and n408 n17326_not ; n17327
g17072 and n17194_not n17327 ; n17328
g17073 and n17322_not n17328_not ; n17329
g17074 and b[34]_not n17329_not ; n17330
g17075 and n16677_not quotient[15]_not ; n17331
g17076 and n16687_not n17112 ; n17332
g17077 and n17108_not n17332 ; n17333
g17078 and n17109_not n17112_not ; n17334
g17079 and n17333_not n17334_not ; n17335
g17080 and n408 n17335_not ; n17336
g17081 and n17194_not n17336 ; n17337
g17082 and n17331_not n17337_not ; n17338
g17083 and b[33]_not n17338_not ; n17339
g17084 and n16686_not quotient[15]_not ; n17340
g17085 and n16696_not n17107 ; n17341
g17086 and n17103_not n17341 ; n17342
g17087 and n17104_not n17107_not ; n17343
g17088 and n17342_not n17343_not ; n17344
g17089 and n408 n17344_not ; n17345
g17090 and n17194_not n17345 ; n17346
g17091 and n17340_not n17346_not ; n17347
g17092 and b[32]_not n17347_not ; n17348
g17093 and n16695_not quotient[15]_not ; n17349
g17094 and n16705_not n17102 ; n17350
g17095 and n17098_not n17350 ; n17351
g17096 and n17099_not n17102_not ; n17352
g17097 and n17351_not n17352_not ; n17353
g17098 and n408 n17353_not ; n17354
g17099 and n17194_not n17354 ; n17355
g17100 and n17349_not n17355_not ; n17356
g17101 and b[31]_not n17356_not ; n17357
g17102 and n16704_not quotient[15]_not ; n17358
g17103 and n16714_not n17097 ; n17359
g17104 and n17093_not n17359 ; n17360
g17105 and n17094_not n17097_not ; n17361
g17106 and n17360_not n17361_not ; n17362
g17107 and n408 n17362_not ; n17363
g17108 and n17194_not n17363 ; n17364
g17109 and n17358_not n17364_not ; n17365
g17110 and b[30]_not n17365_not ; n17366
g17111 and n16713_not quotient[15]_not ; n17367
g17112 and n16723_not n17092 ; n17368
g17113 and n17088_not n17368 ; n17369
g17114 and n17089_not n17092_not ; n17370
g17115 and n17369_not n17370_not ; n17371
g17116 and n408 n17371_not ; n17372
g17117 and n17194_not n17372 ; n17373
g17118 and n17367_not n17373_not ; n17374
g17119 and b[29]_not n17374_not ; n17375
g17120 and n16722_not quotient[15]_not ; n17376
g17121 and n16732_not n17087 ; n17377
g17122 and n17083_not n17377 ; n17378
g17123 and n17084_not n17087_not ; n17379
g17124 and n17378_not n17379_not ; n17380
g17125 and n408 n17380_not ; n17381
g17126 and n17194_not n17381 ; n17382
g17127 and n17376_not n17382_not ; n17383
g17128 and b[28]_not n17383_not ; n17384
g17129 and n16731_not quotient[15]_not ; n17385
g17130 and n16741_not n17082 ; n17386
g17131 and n17078_not n17386 ; n17387
g17132 and n17079_not n17082_not ; n17388
g17133 and n17387_not n17388_not ; n17389
g17134 and n408 n17389_not ; n17390
g17135 and n17194_not n17390 ; n17391
g17136 and n17385_not n17391_not ; n17392
g17137 and b[27]_not n17392_not ; n17393
g17138 and n16740_not quotient[15]_not ; n17394
g17139 and n16750_not n17077 ; n17395
g17140 and n17073_not n17395 ; n17396
g17141 and n17074_not n17077_not ; n17397
g17142 and n17396_not n17397_not ; n17398
g17143 and n408 n17398_not ; n17399
g17144 and n17194_not n17399 ; n17400
g17145 and n17394_not n17400_not ; n17401
g17146 and b[26]_not n17401_not ; n17402
g17147 and n16749_not quotient[15]_not ; n17403
g17148 and n16759_not n17072 ; n17404
g17149 and n17068_not n17404 ; n17405
g17150 and n17069_not n17072_not ; n17406
g17151 and n17405_not n17406_not ; n17407
g17152 and n408 n17407_not ; n17408
g17153 and n17194_not n17408 ; n17409
g17154 and n17403_not n17409_not ; n17410
g17155 and b[25]_not n17410_not ; n17411
g17156 and n16758_not quotient[15]_not ; n17412
g17157 and n16768_not n17067 ; n17413
g17158 and n17063_not n17413 ; n17414
g17159 and n17064_not n17067_not ; n17415
g17160 and n17414_not n17415_not ; n17416
g17161 and n408 n17416_not ; n17417
g17162 and n17194_not n17417 ; n17418
g17163 and n17412_not n17418_not ; n17419
g17164 and b[24]_not n17419_not ; n17420
g17165 and n16767_not quotient[15]_not ; n17421
g17166 and n16777_not n17062 ; n17422
g17167 and n17058_not n17422 ; n17423
g17168 and n17059_not n17062_not ; n17424
g17169 and n17423_not n17424_not ; n17425
g17170 and n408 n17425_not ; n17426
g17171 and n17194_not n17426 ; n17427
g17172 and n17421_not n17427_not ; n17428
g17173 and b[23]_not n17428_not ; n17429
g17174 and n16776_not quotient[15]_not ; n17430
g17175 and n16786_not n17057 ; n17431
g17176 and n17053_not n17431 ; n17432
g17177 and n17054_not n17057_not ; n17433
g17178 and n17432_not n17433_not ; n17434
g17179 and n408 n17434_not ; n17435
g17180 and n17194_not n17435 ; n17436
g17181 and n17430_not n17436_not ; n17437
g17182 and b[22]_not n17437_not ; n17438
g17183 and n16785_not quotient[15]_not ; n17439
g17184 and n16795_not n17052 ; n17440
g17185 and n17048_not n17440 ; n17441
g17186 and n17049_not n17052_not ; n17442
g17187 and n17441_not n17442_not ; n17443
g17188 and n408 n17443_not ; n17444
g17189 and n17194_not n17444 ; n17445
g17190 and n17439_not n17445_not ; n17446
g17191 and b[21]_not n17446_not ; n17447
g17192 and n16794_not quotient[15]_not ; n17448
g17193 and n16804_not n17047 ; n17449
g17194 and n17043_not n17449 ; n17450
g17195 and n17044_not n17047_not ; n17451
g17196 and n17450_not n17451_not ; n17452
g17197 and n408 n17452_not ; n17453
g17198 and n17194_not n17453 ; n17454
g17199 and n17448_not n17454_not ; n17455
g17200 and b[20]_not n17455_not ; n17456
g17201 and n16803_not quotient[15]_not ; n17457
g17202 and n16813_not n17042 ; n17458
g17203 and n17038_not n17458 ; n17459
g17204 and n17039_not n17042_not ; n17460
g17205 and n17459_not n17460_not ; n17461
g17206 and n408 n17461_not ; n17462
g17207 and n17194_not n17462 ; n17463
g17208 and n17457_not n17463_not ; n17464
g17209 and b[19]_not n17464_not ; n17465
g17210 and n16812_not quotient[15]_not ; n17466
g17211 and n16822_not n17037 ; n17467
g17212 and n17033_not n17467 ; n17468
g17213 and n17034_not n17037_not ; n17469
g17214 and n17468_not n17469_not ; n17470
g17215 and n408 n17470_not ; n17471
g17216 and n17194_not n17471 ; n17472
g17217 and n17466_not n17472_not ; n17473
g17218 and b[18]_not n17473_not ; n17474
g17219 and n16821_not quotient[15]_not ; n17475
g17220 and n16831_not n17032 ; n17476
g17221 and n17028_not n17476 ; n17477
g17222 and n17029_not n17032_not ; n17478
g17223 and n17477_not n17478_not ; n17479
g17224 and n408 n17479_not ; n17480
g17225 and n17194_not n17480 ; n17481
g17226 and n17475_not n17481_not ; n17482
g17227 and b[17]_not n17482_not ; n17483
g17228 and n16830_not quotient[15]_not ; n17484
g17229 and n16840_not n17027 ; n17485
g17230 and n17023_not n17485 ; n17486
g17231 and n17024_not n17027_not ; n17487
g17232 and n17486_not n17487_not ; n17488
g17233 and n408 n17488_not ; n17489
g17234 and n17194_not n17489 ; n17490
g17235 and n17484_not n17490_not ; n17491
g17236 and b[16]_not n17491_not ; n17492
g17237 and n16839_not quotient[15]_not ; n17493
g17238 and n16849_not n17022 ; n17494
g17239 and n17018_not n17494 ; n17495
g17240 and n17019_not n17022_not ; n17496
g17241 and n17495_not n17496_not ; n17497
g17242 and n408 n17497_not ; n17498
g17243 and n17194_not n17498 ; n17499
g17244 and n17493_not n17499_not ; n17500
g17245 and b[15]_not n17500_not ; n17501
g17246 and n16848_not quotient[15]_not ; n17502
g17247 and n16858_not n17017 ; n17503
g17248 and n17013_not n17503 ; n17504
g17249 and n17014_not n17017_not ; n17505
g17250 and n17504_not n17505_not ; n17506
g17251 and n408 n17506_not ; n17507
g17252 and n17194_not n17507 ; n17508
g17253 and n17502_not n17508_not ; n17509
g17254 and b[14]_not n17509_not ; n17510
g17255 and n16857_not quotient[15]_not ; n17511
g17256 and n16867_not n17012 ; n17512
g17257 and n17008_not n17512 ; n17513
g17258 and n17009_not n17012_not ; n17514
g17259 and n17513_not n17514_not ; n17515
g17260 and n408 n17515_not ; n17516
g17261 and n17194_not n17516 ; n17517
g17262 and n17511_not n17517_not ; n17518
g17263 and b[13]_not n17518_not ; n17519
g17264 and n16866_not quotient[15]_not ; n17520
g17265 and n16876_not n17007 ; n17521
g17266 and n17003_not n17521 ; n17522
g17267 and n17004_not n17007_not ; n17523
g17268 and n17522_not n17523_not ; n17524
g17269 and n408 n17524_not ; n17525
g17270 and n17194_not n17525 ; n17526
g17271 and n17520_not n17526_not ; n17527
g17272 and b[12]_not n17527_not ; n17528
g17273 and n16875_not quotient[15]_not ; n17529
g17274 and n16885_not n17002 ; n17530
g17275 and n16998_not n17530 ; n17531
g17276 and n16999_not n17002_not ; n17532
g17277 and n17531_not n17532_not ; n17533
g17278 and n408 n17533_not ; n17534
g17279 and n17194_not n17534 ; n17535
g17280 and n17529_not n17535_not ; n17536
g17281 and b[11]_not n17536_not ; n17537
g17282 and n16884_not quotient[15]_not ; n17538
g17283 and n16894_not n16997 ; n17539
g17284 and n16993_not n17539 ; n17540
g17285 and n16994_not n16997_not ; n17541
g17286 and n17540_not n17541_not ; n17542
g17287 and n408 n17542_not ; n17543
g17288 and n17194_not n17543 ; n17544
g17289 and n17538_not n17544_not ; n17545
g17290 and b[10]_not n17545_not ; n17546
g17291 and n16893_not quotient[15]_not ; n17547
g17292 and n16903_not n16992 ; n17548
g17293 and n16988_not n17548 ; n17549
g17294 and n16989_not n16992_not ; n17550
g17295 and n17549_not n17550_not ; n17551
g17296 and n408 n17551_not ; n17552
g17297 and n17194_not n17552 ; n17553
g17298 and n17547_not n17553_not ; n17554
g17299 and b[9]_not n17554_not ; n17555
g17300 and n16902_not quotient[15]_not ; n17556
g17301 and n16912_not n16987 ; n17557
g17302 and n16983_not n17557 ; n17558
g17303 and n16984_not n16987_not ; n17559
g17304 and n17558_not n17559_not ; n17560
g17305 and n408 n17560_not ; n17561
g17306 and n17194_not n17561 ; n17562
g17307 and n17556_not n17562_not ; n17563
g17308 and b[8]_not n17563_not ; n17564
g17309 and n16911_not quotient[15]_not ; n17565
g17310 and n16921_not n16982 ; n17566
g17311 and n16978_not n17566 ; n17567
g17312 and n16979_not n16982_not ; n17568
g17313 and n17567_not n17568_not ; n17569
g17314 and n408 n17569_not ; n17570
g17315 and n17194_not n17570 ; n17571
g17316 and n17565_not n17571_not ; n17572
g17317 and b[7]_not n17572_not ; n17573
g17318 and n16920_not quotient[15]_not ; n17574
g17319 and n16930_not n16977 ; n17575
g17320 and n16973_not n17575 ; n17576
g17321 and n16974_not n16977_not ; n17577
g17322 and n17576_not n17577_not ; n17578
g17323 and n408 n17578_not ; n17579
g17324 and n17194_not n17579 ; n17580
g17325 and n17574_not n17580_not ; n17581
g17326 and b[6]_not n17581_not ; n17582
g17327 and n16929_not quotient[15]_not ; n17583
g17328 and n16939_not n16972 ; n17584
g17329 and n16968_not n17584 ; n17585
g17330 and n16969_not n16972_not ; n17586
g17331 and n17585_not n17586_not ; n17587
g17332 and n408 n17587_not ; n17588
g17333 and n17194_not n17588 ; n17589
g17334 and n17583_not n17589_not ; n17590
g17335 and b[5]_not n17590_not ; n17591
g17336 and n16938_not quotient[15]_not ; n17592
g17337 and n16947_not n16967 ; n17593
g17338 and n16963_not n17593 ; n17594
g17339 and n16964_not n16967_not ; n17595
g17340 and n17594_not n17595_not ; n17596
g17341 and n408 n17596_not ; n17597
g17342 and n17194_not n17597 ; n17598
g17343 and n17592_not n17598_not ; n17599
g17344 and b[4]_not n17599_not ; n17600
g17345 and n16946_not quotient[15]_not ; n17601
g17346 and n16958_not n16962 ; n17602
g17347 and n16957_not n17602 ; n17603
g17348 and n16959_not n16962_not ; n17604
g17349 and n17603_not n17604_not ; n17605
g17350 and n408 n17605_not ; n17606
g17351 and n17194_not n17606 ; n17607
g17352 and n17601_not n17607_not ; n17608
g17353 and b[3]_not n17608_not ; n17609
g17354 and n16951_not quotient[15]_not ; n17610
g17355 and n16954_not n16956 ; n17611
g17356 and n16952_not n17611 ; n17612
g17357 and n408 n17612_not ; n17613
g17358 and n16957_not n17613 ; n17614
g17359 and n17194_not n17614 ; n17615
g17360 and n17610_not n17615_not ; n17616
g17361 and b[2]_not n17616_not ; n17617
g17362 and b[0] b[49]_not ; n17618
g17363 and n297 n17618 ; n17619
g17364 and n286 n17619 ; n17620
g17365 and n337 n17620 ; n17621
g17366 and n17194_not n17621 ; n17622
g17367 and a[15] n17622_not ; n17623
g17368 and n400 n16956 ; n17624
g17369 and n595 n17624 ; n17625
g17370 and n17194_not n17625 ; n17626
g17371 and n17623_not n17626_not ; n17627
g17372 and b[1] n17627_not ; n17628
g17373 and b[1]_not n17626_not ; n17629
g17374 and n17623_not n17629 ; n17630
g17375 and n17628_not n17630_not ; n17631
g17376 and a[14]_not b[0] ; n17632
g17377 and n17631_not n17632_not ; n17633
g17378 and b[1]_not n17627_not ; n17634
g17379 and n17633_not n17634_not ; n17635
g17380 and b[2] n17615_not ; n17636
g17381 and n17610_not n17636 ; n17637
g17382 and n17617_not n17637_not ; n17638
g17383 and n17635_not n17638 ; n17639
g17384 and n17617_not n17639_not ; n17640
g17385 and b[3] n17607_not ; n17641
g17386 and n17601_not n17641 ; n17642
g17387 and n17609_not n17642_not ; n17643
g17388 and n17640_not n17643 ; n17644
g17389 and n17609_not n17644_not ; n17645
g17390 and b[4] n17598_not ; n17646
g17391 and n17592_not n17646 ; n17647
g17392 and n17600_not n17647_not ; n17648
g17393 and n17645_not n17648 ; n17649
g17394 and n17600_not n17649_not ; n17650
g17395 and b[5] n17589_not ; n17651
g17396 and n17583_not n17651 ; n17652
g17397 and n17591_not n17652_not ; n17653
g17398 and n17650_not n17653 ; n17654
g17399 and n17591_not n17654_not ; n17655
g17400 and b[6] n17580_not ; n17656
g17401 and n17574_not n17656 ; n17657
g17402 and n17582_not n17657_not ; n17658
g17403 and n17655_not n17658 ; n17659
g17404 and n17582_not n17659_not ; n17660
g17405 and b[7] n17571_not ; n17661
g17406 and n17565_not n17661 ; n17662
g17407 and n17573_not n17662_not ; n17663
g17408 and n17660_not n17663 ; n17664
g17409 and n17573_not n17664_not ; n17665
g17410 and b[8] n17562_not ; n17666
g17411 and n17556_not n17666 ; n17667
g17412 and n17564_not n17667_not ; n17668
g17413 and n17665_not n17668 ; n17669
g17414 and n17564_not n17669_not ; n17670
g17415 and b[9] n17553_not ; n17671
g17416 and n17547_not n17671 ; n17672
g17417 and n17555_not n17672_not ; n17673
g17418 and n17670_not n17673 ; n17674
g17419 and n17555_not n17674_not ; n17675
g17420 and b[10] n17544_not ; n17676
g17421 and n17538_not n17676 ; n17677
g17422 and n17546_not n17677_not ; n17678
g17423 and n17675_not n17678 ; n17679
g17424 and n17546_not n17679_not ; n17680
g17425 and b[11] n17535_not ; n17681
g17426 and n17529_not n17681 ; n17682
g17427 and n17537_not n17682_not ; n17683
g17428 and n17680_not n17683 ; n17684
g17429 and n17537_not n17684_not ; n17685
g17430 and b[12] n17526_not ; n17686
g17431 and n17520_not n17686 ; n17687
g17432 and n17528_not n17687_not ; n17688
g17433 and n17685_not n17688 ; n17689
g17434 and n17528_not n17689_not ; n17690
g17435 and b[13] n17517_not ; n17691
g17436 and n17511_not n17691 ; n17692
g17437 and n17519_not n17692_not ; n17693
g17438 and n17690_not n17693 ; n17694
g17439 and n17519_not n17694_not ; n17695
g17440 and b[14] n17508_not ; n17696
g17441 and n17502_not n17696 ; n17697
g17442 and n17510_not n17697_not ; n17698
g17443 and n17695_not n17698 ; n17699
g17444 and n17510_not n17699_not ; n17700
g17445 and b[15] n17499_not ; n17701
g17446 and n17493_not n17701 ; n17702
g17447 and n17501_not n17702_not ; n17703
g17448 and n17700_not n17703 ; n17704
g17449 and n17501_not n17704_not ; n17705
g17450 and b[16] n17490_not ; n17706
g17451 and n17484_not n17706 ; n17707
g17452 and n17492_not n17707_not ; n17708
g17453 and n17705_not n17708 ; n17709
g17454 and n17492_not n17709_not ; n17710
g17455 and b[17] n17481_not ; n17711
g17456 and n17475_not n17711 ; n17712
g17457 and n17483_not n17712_not ; n17713
g17458 and n17710_not n17713 ; n17714
g17459 and n17483_not n17714_not ; n17715
g17460 and b[18] n17472_not ; n17716
g17461 and n17466_not n17716 ; n17717
g17462 and n17474_not n17717_not ; n17718
g17463 and n17715_not n17718 ; n17719
g17464 and n17474_not n17719_not ; n17720
g17465 and b[19] n17463_not ; n17721
g17466 and n17457_not n17721 ; n17722
g17467 and n17465_not n17722_not ; n17723
g17468 and n17720_not n17723 ; n17724
g17469 and n17465_not n17724_not ; n17725
g17470 and b[20] n17454_not ; n17726
g17471 and n17448_not n17726 ; n17727
g17472 and n17456_not n17727_not ; n17728
g17473 and n17725_not n17728 ; n17729
g17474 and n17456_not n17729_not ; n17730
g17475 and b[21] n17445_not ; n17731
g17476 and n17439_not n17731 ; n17732
g17477 and n17447_not n17732_not ; n17733
g17478 and n17730_not n17733 ; n17734
g17479 and n17447_not n17734_not ; n17735
g17480 and b[22] n17436_not ; n17736
g17481 and n17430_not n17736 ; n17737
g17482 and n17438_not n17737_not ; n17738
g17483 and n17735_not n17738 ; n17739
g17484 and n17438_not n17739_not ; n17740
g17485 and b[23] n17427_not ; n17741
g17486 and n17421_not n17741 ; n17742
g17487 and n17429_not n17742_not ; n17743
g17488 and n17740_not n17743 ; n17744
g17489 and n17429_not n17744_not ; n17745
g17490 and b[24] n17418_not ; n17746
g17491 and n17412_not n17746 ; n17747
g17492 and n17420_not n17747_not ; n17748
g17493 and n17745_not n17748 ; n17749
g17494 and n17420_not n17749_not ; n17750
g17495 and b[25] n17409_not ; n17751
g17496 and n17403_not n17751 ; n17752
g17497 and n17411_not n17752_not ; n17753
g17498 and n17750_not n17753 ; n17754
g17499 and n17411_not n17754_not ; n17755
g17500 and b[26] n17400_not ; n17756
g17501 and n17394_not n17756 ; n17757
g17502 and n17402_not n17757_not ; n17758
g17503 and n17755_not n17758 ; n17759
g17504 and n17402_not n17759_not ; n17760
g17505 and b[27] n17391_not ; n17761
g17506 and n17385_not n17761 ; n17762
g17507 and n17393_not n17762_not ; n17763
g17508 and n17760_not n17763 ; n17764
g17509 and n17393_not n17764_not ; n17765
g17510 and b[28] n17382_not ; n17766
g17511 and n17376_not n17766 ; n17767
g17512 and n17384_not n17767_not ; n17768
g17513 and n17765_not n17768 ; n17769
g17514 and n17384_not n17769_not ; n17770
g17515 and b[29] n17373_not ; n17771
g17516 and n17367_not n17771 ; n17772
g17517 and n17375_not n17772_not ; n17773
g17518 and n17770_not n17773 ; n17774
g17519 and n17375_not n17774_not ; n17775
g17520 and b[30] n17364_not ; n17776
g17521 and n17358_not n17776 ; n17777
g17522 and n17366_not n17777_not ; n17778
g17523 and n17775_not n17778 ; n17779
g17524 and n17366_not n17779_not ; n17780
g17525 and b[31] n17355_not ; n17781
g17526 and n17349_not n17781 ; n17782
g17527 and n17357_not n17782_not ; n17783
g17528 and n17780_not n17783 ; n17784
g17529 and n17357_not n17784_not ; n17785
g17530 and b[32] n17346_not ; n17786
g17531 and n17340_not n17786 ; n17787
g17532 and n17348_not n17787_not ; n17788
g17533 and n17785_not n17788 ; n17789
g17534 and n17348_not n17789_not ; n17790
g17535 and b[33] n17337_not ; n17791
g17536 and n17331_not n17791 ; n17792
g17537 and n17339_not n17792_not ; n17793
g17538 and n17790_not n17793 ; n17794
g17539 and n17339_not n17794_not ; n17795
g17540 and b[34] n17328_not ; n17796
g17541 and n17322_not n17796 ; n17797
g17542 and n17330_not n17797_not ; n17798
g17543 and n17795_not n17798 ; n17799
g17544 and n17330_not n17799_not ; n17800
g17545 and b[35] n17319_not ; n17801
g17546 and n17313_not n17801 ; n17802
g17547 and n17321_not n17802_not ; n17803
g17548 and n17800_not n17803 ; n17804
g17549 and n17321_not n17804_not ; n17805
g17550 and b[36] n17310_not ; n17806
g17551 and n17304_not n17806 ; n17807
g17552 and n17312_not n17807_not ; n17808
g17553 and n17805_not n17808 ; n17809
g17554 and n17312_not n17809_not ; n17810
g17555 and b[37] n17301_not ; n17811
g17556 and n17295_not n17811 ; n17812
g17557 and n17303_not n17812_not ; n17813
g17558 and n17810_not n17813 ; n17814
g17559 and n17303_not n17814_not ; n17815
g17560 and b[38] n17292_not ; n17816
g17561 and n17286_not n17816 ; n17817
g17562 and n17294_not n17817_not ; n17818
g17563 and n17815_not n17818 ; n17819
g17564 and n17294_not n17819_not ; n17820
g17565 and b[39] n17283_not ; n17821
g17566 and n17277_not n17821 ; n17822
g17567 and n17285_not n17822_not ; n17823
g17568 and n17820_not n17823 ; n17824
g17569 and n17285_not n17824_not ; n17825
g17570 and b[40] n17274_not ; n17826
g17571 and n17268_not n17826 ; n17827
g17572 and n17276_not n17827_not ; n17828
g17573 and n17825_not n17828 ; n17829
g17574 and n17276_not n17829_not ; n17830
g17575 and b[41] n17265_not ; n17831
g17576 and n17259_not n17831 ; n17832
g17577 and n17267_not n17832_not ; n17833
g17578 and n17830_not n17833 ; n17834
g17579 and n17267_not n17834_not ; n17835
g17580 and b[42] n17256_not ; n17836
g17581 and n17250_not n17836 ; n17837
g17582 and n17258_not n17837_not ; n17838
g17583 and n17835_not n17838 ; n17839
g17584 and n17258_not n17839_not ; n17840
g17585 and b[43] n17247_not ; n17841
g17586 and n17241_not n17841 ; n17842
g17587 and n17249_not n17842_not ; n17843
g17588 and n17840_not n17843 ; n17844
g17589 and n17249_not n17844_not ; n17845
g17590 and b[44] n17238_not ; n17846
g17591 and n17232_not n17846 ; n17847
g17592 and n17240_not n17847_not ; n17848
g17593 and n17845_not n17848 ; n17849
g17594 and n17240_not n17849_not ; n17850
g17595 and b[45] n17229_not ; n17851
g17596 and n17223_not n17851 ; n17852
g17597 and n17231_not n17852_not ; n17853
g17598 and n17850_not n17853 ; n17854
g17599 and n17231_not n17854_not ; n17855
g17600 and b[46] n17220_not ; n17856
g17601 and n17214_not n17856 ; n17857
g17602 and n17222_not n17857_not ; n17858
g17603 and n17855_not n17858 ; n17859
g17604 and n17222_not n17859_not ; n17860
g17605 and b[47] n17211_not ; n17861
g17606 and n17205_not n17861 ; n17862
g17607 and n17213_not n17862_not ; n17863
g17608 and n17860_not n17863 ; n17864
g17609 and n17213_not n17864_not ; n17865
g17610 and b[48] n17202_not ; n17866
g17611 and n17196_not n17866 ; n17867
g17612 and n17204_not n17867_not ; n17868
g17613 and n17865_not n17868 ; n17869
g17614 and n17204_not n17869_not ; n17870
g17615 and n16541_not quotient[15]_not ; n17871
g17616 and n16543_not n17192 ; n17872
g17617 and n17188_not n17872 ; n17873
g17618 and n17189_not n17192_not ; n17874
g17619 and n17873_not n17874_not ; n17875
g17620 and quotient[15] n17875_not ; n17876
g17621 and n17871_not n17876_not ; n17877
g17622 and b[49]_not n17877_not ; n17878
g17623 and b[49] n17871_not ; n17879
g17624 and n17876_not n17879 ; n17880
g17625 and n286 n297 ; n17881
g17626 and n337 n17881 ; n17882
g17627 and n17880_not n17882 ; n17883
g17628 and n17878_not n17883 ; n17884
g17629 and n17870_not n17884 ; n17885
g17630 and n408 n17877_not ; n17886
g17631 and n17885_not n17886_not ; quotient[14]
g17632 and n17213_not n17868 ; n17888
g17633 and n17864_not n17888 ; n17889
g17634 and n17865_not n17868_not ; n17890
g17635 and n17889_not n17890_not ; n17891
g17636 and quotient[14] n17891_not ; n17892
g17637 and n17203_not n17886_not ; n17893
g17638 and n17885_not n17893 ; n17894
g17639 and n17892_not n17894_not ; n17895
g17640 and b[49]_not n17895_not ; n17896
g17641 and n17222_not n17863 ; n17897
g17642 and n17859_not n17897 ; n17898
g17643 and n17860_not n17863_not ; n17899
g17644 and n17898_not n17899_not ; n17900
g17645 and quotient[14] n17900_not ; n17901
g17646 and n17212_not n17886_not ; n17902
g17647 and n17885_not n17902 ; n17903
g17648 and n17901_not n17903_not ; n17904
g17649 and b[48]_not n17904_not ; n17905
g17650 and n17231_not n17858 ; n17906
g17651 and n17854_not n17906 ; n17907
g17652 and n17855_not n17858_not ; n17908
g17653 and n17907_not n17908_not ; n17909
g17654 and quotient[14] n17909_not ; n17910
g17655 and n17221_not n17886_not ; n17911
g17656 and n17885_not n17911 ; n17912
g17657 and n17910_not n17912_not ; n17913
g17658 and b[47]_not n17913_not ; n17914
g17659 and n17240_not n17853 ; n17915
g17660 and n17849_not n17915 ; n17916
g17661 and n17850_not n17853_not ; n17917
g17662 and n17916_not n17917_not ; n17918
g17663 and quotient[14] n17918_not ; n17919
g17664 and n17230_not n17886_not ; n17920
g17665 and n17885_not n17920 ; n17921
g17666 and n17919_not n17921_not ; n17922
g17667 and b[46]_not n17922_not ; n17923
g17668 and n17249_not n17848 ; n17924
g17669 and n17844_not n17924 ; n17925
g17670 and n17845_not n17848_not ; n17926
g17671 and n17925_not n17926_not ; n17927
g17672 and quotient[14] n17927_not ; n17928
g17673 and n17239_not n17886_not ; n17929
g17674 and n17885_not n17929 ; n17930
g17675 and n17928_not n17930_not ; n17931
g17676 and b[45]_not n17931_not ; n17932
g17677 and n17258_not n17843 ; n17933
g17678 and n17839_not n17933 ; n17934
g17679 and n17840_not n17843_not ; n17935
g17680 and n17934_not n17935_not ; n17936
g17681 and quotient[14] n17936_not ; n17937
g17682 and n17248_not n17886_not ; n17938
g17683 and n17885_not n17938 ; n17939
g17684 and n17937_not n17939_not ; n17940
g17685 and b[44]_not n17940_not ; n17941
g17686 and n17267_not n17838 ; n17942
g17687 and n17834_not n17942 ; n17943
g17688 and n17835_not n17838_not ; n17944
g17689 and n17943_not n17944_not ; n17945
g17690 and quotient[14] n17945_not ; n17946
g17691 and n17257_not n17886_not ; n17947
g17692 and n17885_not n17947 ; n17948
g17693 and n17946_not n17948_not ; n17949
g17694 and b[43]_not n17949_not ; n17950
g17695 and n17276_not n17833 ; n17951
g17696 and n17829_not n17951 ; n17952
g17697 and n17830_not n17833_not ; n17953
g17698 and n17952_not n17953_not ; n17954
g17699 and quotient[14] n17954_not ; n17955
g17700 and n17266_not n17886_not ; n17956
g17701 and n17885_not n17956 ; n17957
g17702 and n17955_not n17957_not ; n17958
g17703 and b[42]_not n17958_not ; n17959
g17704 and n17285_not n17828 ; n17960
g17705 and n17824_not n17960 ; n17961
g17706 and n17825_not n17828_not ; n17962
g17707 and n17961_not n17962_not ; n17963
g17708 and quotient[14] n17963_not ; n17964
g17709 and n17275_not n17886_not ; n17965
g17710 and n17885_not n17965 ; n17966
g17711 and n17964_not n17966_not ; n17967
g17712 and b[41]_not n17967_not ; n17968
g17713 and n17294_not n17823 ; n17969
g17714 and n17819_not n17969 ; n17970
g17715 and n17820_not n17823_not ; n17971
g17716 and n17970_not n17971_not ; n17972
g17717 and quotient[14] n17972_not ; n17973
g17718 and n17284_not n17886_not ; n17974
g17719 and n17885_not n17974 ; n17975
g17720 and n17973_not n17975_not ; n17976
g17721 and b[40]_not n17976_not ; n17977
g17722 and n17303_not n17818 ; n17978
g17723 and n17814_not n17978 ; n17979
g17724 and n17815_not n17818_not ; n17980
g17725 and n17979_not n17980_not ; n17981
g17726 and quotient[14] n17981_not ; n17982
g17727 and n17293_not n17886_not ; n17983
g17728 and n17885_not n17983 ; n17984
g17729 and n17982_not n17984_not ; n17985
g17730 and b[39]_not n17985_not ; n17986
g17731 and n17312_not n17813 ; n17987
g17732 and n17809_not n17987 ; n17988
g17733 and n17810_not n17813_not ; n17989
g17734 and n17988_not n17989_not ; n17990
g17735 and quotient[14] n17990_not ; n17991
g17736 and n17302_not n17886_not ; n17992
g17737 and n17885_not n17992 ; n17993
g17738 and n17991_not n17993_not ; n17994
g17739 and b[38]_not n17994_not ; n17995
g17740 and n17321_not n17808 ; n17996
g17741 and n17804_not n17996 ; n17997
g17742 and n17805_not n17808_not ; n17998
g17743 and n17997_not n17998_not ; n17999
g17744 and quotient[14] n17999_not ; n18000
g17745 and n17311_not n17886_not ; n18001
g17746 and n17885_not n18001 ; n18002
g17747 and n18000_not n18002_not ; n18003
g17748 and b[37]_not n18003_not ; n18004
g17749 and n17330_not n17803 ; n18005
g17750 and n17799_not n18005 ; n18006
g17751 and n17800_not n17803_not ; n18007
g17752 and n18006_not n18007_not ; n18008
g17753 and quotient[14] n18008_not ; n18009
g17754 and n17320_not n17886_not ; n18010
g17755 and n17885_not n18010 ; n18011
g17756 and n18009_not n18011_not ; n18012
g17757 and b[36]_not n18012_not ; n18013
g17758 and n17339_not n17798 ; n18014
g17759 and n17794_not n18014 ; n18015
g17760 and n17795_not n17798_not ; n18016
g17761 and n18015_not n18016_not ; n18017
g17762 and quotient[14] n18017_not ; n18018
g17763 and n17329_not n17886_not ; n18019
g17764 and n17885_not n18019 ; n18020
g17765 and n18018_not n18020_not ; n18021
g17766 and b[35]_not n18021_not ; n18022
g17767 and n17348_not n17793 ; n18023
g17768 and n17789_not n18023 ; n18024
g17769 and n17790_not n17793_not ; n18025
g17770 and n18024_not n18025_not ; n18026
g17771 and quotient[14] n18026_not ; n18027
g17772 and n17338_not n17886_not ; n18028
g17773 and n17885_not n18028 ; n18029
g17774 and n18027_not n18029_not ; n18030
g17775 and b[34]_not n18030_not ; n18031
g17776 and n17357_not n17788 ; n18032
g17777 and n17784_not n18032 ; n18033
g17778 and n17785_not n17788_not ; n18034
g17779 and n18033_not n18034_not ; n18035
g17780 and quotient[14] n18035_not ; n18036
g17781 and n17347_not n17886_not ; n18037
g17782 and n17885_not n18037 ; n18038
g17783 and n18036_not n18038_not ; n18039
g17784 and b[33]_not n18039_not ; n18040
g17785 and n17366_not n17783 ; n18041
g17786 and n17779_not n18041 ; n18042
g17787 and n17780_not n17783_not ; n18043
g17788 and n18042_not n18043_not ; n18044
g17789 and quotient[14] n18044_not ; n18045
g17790 and n17356_not n17886_not ; n18046
g17791 and n17885_not n18046 ; n18047
g17792 and n18045_not n18047_not ; n18048
g17793 and b[32]_not n18048_not ; n18049
g17794 and n17375_not n17778 ; n18050
g17795 and n17774_not n18050 ; n18051
g17796 and n17775_not n17778_not ; n18052
g17797 and n18051_not n18052_not ; n18053
g17798 and quotient[14] n18053_not ; n18054
g17799 and n17365_not n17886_not ; n18055
g17800 and n17885_not n18055 ; n18056
g17801 and n18054_not n18056_not ; n18057
g17802 and b[31]_not n18057_not ; n18058
g17803 and n17384_not n17773 ; n18059
g17804 and n17769_not n18059 ; n18060
g17805 and n17770_not n17773_not ; n18061
g17806 and n18060_not n18061_not ; n18062
g17807 and quotient[14] n18062_not ; n18063
g17808 and n17374_not n17886_not ; n18064
g17809 and n17885_not n18064 ; n18065
g17810 and n18063_not n18065_not ; n18066
g17811 and b[30]_not n18066_not ; n18067
g17812 and n17393_not n17768 ; n18068
g17813 and n17764_not n18068 ; n18069
g17814 and n17765_not n17768_not ; n18070
g17815 and n18069_not n18070_not ; n18071
g17816 and quotient[14] n18071_not ; n18072
g17817 and n17383_not n17886_not ; n18073
g17818 and n17885_not n18073 ; n18074
g17819 and n18072_not n18074_not ; n18075
g17820 and b[29]_not n18075_not ; n18076
g17821 and n17402_not n17763 ; n18077
g17822 and n17759_not n18077 ; n18078
g17823 and n17760_not n17763_not ; n18079
g17824 and n18078_not n18079_not ; n18080
g17825 and quotient[14] n18080_not ; n18081
g17826 and n17392_not n17886_not ; n18082
g17827 and n17885_not n18082 ; n18083
g17828 and n18081_not n18083_not ; n18084
g17829 and b[28]_not n18084_not ; n18085
g17830 and n17411_not n17758 ; n18086
g17831 and n17754_not n18086 ; n18087
g17832 and n17755_not n17758_not ; n18088
g17833 and n18087_not n18088_not ; n18089
g17834 and quotient[14] n18089_not ; n18090
g17835 and n17401_not n17886_not ; n18091
g17836 and n17885_not n18091 ; n18092
g17837 and n18090_not n18092_not ; n18093
g17838 and b[27]_not n18093_not ; n18094
g17839 and n17420_not n17753 ; n18095
g17840 and n17749_not n18095 ; n18096
g17841 and n17750_not n17753_not ; n18097
g17842 and n18096_not n18097_not ; n18098
g17843 and quotient[14] n18098_not ; n18099
g17844 and n17410_not n17886_not ; n18100
g17845 and n17885_not n18100 ; n18101
g17846 and n18099_not n18101_not ; n18102
g17847 and b[26]_not n18102_not ; n18103
g17848 and n17429_not n17748 ; n18104
g17849 and n17744_not n18104 ; n18105
g17850 and n17745_not n17748_not ; n18106
g17851 and n18105_not n18106_not ; n18107
g17852 and quotient[14] n18107_not ; n18108
g17853 and n17419_not n17886_not ; n18109
g17854 and n17885_not n18109 ; n18110
g17855 and n18108_not n18110_not ; n18111
g17856 and b[25]_not n18111_not ; n18112
g17857 and n17438_not n17743 ; n18113
g17858 and n17739_not n18113 ; n18114
g17859 and n17740_not n17743_not ; n18115
g17860 and n18114_not n18115_not ; n18116
g17861 and quotient[14] n18116_not ; n18117
g17862 and n17428_not n17886_not ; n18118
g17863 and n17885_not n18118 ; n18119
g17864 and n18117_not n18119_not ; n18120
g17865 and b[24]_not n18120_not ; n18121
g17866 and n17447_not n17738 ; n18122
g17867 and n17734_not n18122 ; n18123
g17868 and n17735_not n17738_not ; n18124
g17869 and n18123_not n18124_not ; n18125
g17870 and quotient[14] n18125_not ; n18126
g17871 and n17437_not n17886_not ; n18127
g17872 and n17885_not n18127 ; n18128
g17873 and n18126_not n18128_not ; n18129
g17874 and b[23]_not n18129_not ; n18130
g17875 and n17456_not n17733 ; n18131
g17876 and n17729_not n18131 ; n18132
g17877 and n17730_not n17733_not ; n18133
g17878 and n18132_not n18133_not ; n18134
g17879 and quotient[14] n18134_not ; n18135
g17880 and n17446_not n17886_not ; n18136
g17881 and n17885_not n18136 ; n18137
g17882 and n18135_not n18137_not ; n18138
g17883 and b[22]_not n18138_not ; n18139
g17884 and n17465_not n17728 ; n18140
g17885 and n17724_not n18140 ; n18141
g17886 and n17725_not n17728_not ; n18142
g17887 and n18141_not n18142_not ; n18143
g17888 and quotient[14] n18143_not ; n18144
g17889 and n17455_not n17886_not ; n18145
g17890 and n17885_not n18145 ; n18146
g17891 and n18144_not n18146_not ; n18147
g17892 and b[21]_not n18147_not ; n18148
g17893 and n17474_not n17723 ; n18149
g17894 and n17719_not n18149 ; n18150
g17895 and n17720_not n17723_not ; n18151
g17896 and n18150_not n18151_not ; n18152
g17897 and quotient[14] n18152_not ; n18153
g17898 and n17464_not n17886_not ; n18154
g17899 and n17885_not n18154 ; n18155
g17900 and n18153_not n18155_not ; n18156
g17901 and b[20]_not n18156_not ; n18157
g17902 and n17483_not n17718 ; n18158
g17903 and n17714_not n18158 ; n18159
g17904 and n17715_not n17718_not ; n18160
g17905 and n18159_not n18160_not ; n18161
g17906 and quotient[14] n18161_not ; n18162
g17907 and n17473_not n17886_not ; n18163
g17908 and n17885_not n18163 ; n18164
g17909 and n18162_not n18164_not ; n18165
g17910 and b[19]_not n18165_not ; n18166
g17911 and n17492_not n17713 ; n18167
g17912 and n17709_not n18167 ; n18168
g17913 and n17710_not n17713_not ; n18169
g17914 and n18168_not n18169_not ; n18170
g17915 and quotient[14] n18170_not ; n18171
g17916 and n17482_not n17886_not ; n18172
g17917 and n17885_not n18172 ; n18173
g17918 and n18171_not n18173_not ; n18174
g17919 and b[18]_not n18174_not ; n18175
g17920 and n17501_not n17708 ; n18176
g17921 and n17704_not n18176 ; n18177
g17922 and n17705_not n17708_not ; n18178
g17923 and n18177_not n18178_not ; n18179
g17924 and quotient[14] n18179_not ; n18180
g17925 and n17491_not n17886_not ; n18181
g17926 and n17885_not n18181 ; n18182
g17927 and n18180_not n18182_not ; n18183
g17928 and b[17]_not n18183_not ; n18184
g17929 and n17510_not n17703 ; n18185
g17930 and n17699_not n18185 ; n18186
g17931 and n17700_not n17703_not ; n18187
g17932 and n18186_not n18187_not ; n18188
g17933 and quotient[14] n18188_not ; n18189
g17934 and n17500_not n17886_not ; n18190
g17935 and n17885_not n18190 ; n18191
g17936 and n18189_not n18191_not ; n18192
g17937 and b[16]_not n18192_not ; n18193
g17938 and n17519_not n17698 ; n18194
g17939 and n17694_not n18194 ; n18195
g17940 and n17695_not n17698_not ; n18196
g17941 and n18195_not n18196_not ; n18197
g17942 and quotient[14] n18197_not ; n18198
g17943 and n17509_not n17886_not ; n18199
g17944 and n17885_not n18199 ; n18200
g17945 and n18198_not n18200_not ; n18201
g17946 and b[15]_not n18201_not ; n18202
g17947 and n17528_not n17693 ; n18203
g17948 and n17689_not n18203 ; n18204
g17949 and n17690_not n17693_not ; n18205
g17950 and n18204_not n18205_not ; n18206
g17951 and quotient[14] n18206_not ; n18207
g17952 and n17518_not n17886_not ; n18208
g17953 and n17885_not n18208 ; n18209
g17954 and n18207_not n18209_not ; n18210
g17955 and b[14]_not n18210_not ; n18211
g17956 and n17537_not n17688 ; n18212
g17957 and n17684_not n18212 ; n18213
g17958 and n17685_not n17688_not ; n18214
g17959 and n18213_not n18214_not ; n18215
g17960 and quotient[14] n18215_not ; n18216
g17961 and n17527_not n17886_not ; n18217
g17962 and n17885_not n18217 ; n18218
g17963 and n18216_not n18218_not ; n18219
g17964 and b[13]_not n18219_not ; n18220
g17965 and n17546_not n17683 ; n18221
g17966 and n17679_not n18221 ; n18222
g17967 and n17680_not n17683_not ; n18223
g17968 and n18222_not n18223_not ; n18224
g17969 and quotient[14] n18224_not ; n18225
g17970 and n17536_not n17886_not ; n18226
g17971 and n17885_not n18226 ; n18227
g17972 and n18225_not n18227_not ; n18228
g17973 and b[12]_not n18228_not ; n18229
g17974 and n17555_not n17678 ; n18230
g17975 and n17674_not n18230 ; n18231
g17976 and n17675_not n17678_not ; n18232
g17977 and n18231_not n18232_not ; n18233
g17978 and quotient[14] n18233_not ; n18234
g17979 and n17545_not n17886_not ; n18235
g17980 and n17885_not n18235 ; n18236
g17981 and n18234_not n18236_not ; n18237
g17982 and b[11]_not n18237_not ; n18238
g17983 and n17564_not n17673 ; n18239
g17984 and n17669_not n18239 ; n18240
g17985 and n17670_not n17673_not ; n18241
g17986 and n18240_not n18241_not ; n18242
g17987 and quotient[14] n18242_not ; n18243
g17988 and n17554_not n17886_not ; n18244
g17989 and n17885_not n18244 ; n18245
g17990 and n18243_not n18245_not ; n18246
g17991 and b[10]_not n18246_not ; n18247
g17992 and n17573_not n17668 ; n18248
g17993 and n17664_not n18248 ; n18249
g17994 and n17665_not n17668_not ; n18250
g17995 and n18249_not n18250_not ; n18251
g17996 and quotient[14] n18251_not ; n18252
g17997 and n17563_not n17886_not ; n18253
g17998 and n17885_not n18253 ; n18254
g17999 and n18252_not n18254_not ; n18255
g18000 and b[9]_not n18255_not ; n18256
g18001 and n17582_not n17663 ; n18257
g18002 and n17659_not n18257 ; n18258
g18003 and n17660_not n17663_not ; n18259
g18004 and n18258_not n18259_not ; n18260
g18005 and quotient[14] n18260_not ; n18261
g18006 and n17572_not n17886_not ; n18262
g18007 and n17885_not n18262 ; n18263
g18008 and n18261_not n18263_not ; n18264
g18009 and b[8]_not n18264_not ; n18265
g18010 and n17591_not n17658 ; n18266
g18011 and n17654_not n18266 ; n18267
g18012 and n17655_not n17658_not ; n18268
g18013 and n18267_not n18268_not ; n18269
g18014 and quotient[14] n18269_not ; n18270
g18015 and n17581_not n17886_not ; n18271
g18016 and n17885_not n18271 ; n18272
g18017 and n18270_not n18272_not ; n18273
g18018 and b[7]_not n18273_not ; n18274
g18019 and n17600_not n17653 ; n18275
g18020 and n17649_not n18275 ; n18276
g18021 and n17650_not n17653_not ; n18277
g18022 and n18276_not n18277_not ; n18278
g18023 and quotient[14] n18278_not ; n18279
g18024 and n17590_not n17886_not ; n18280
g18025 and n17885_not n18280 ; n18281
g18026 and n18279_not n18281_not ; n18282
g18027 and b[6]_not n18282_not ; n18283
g18028 and n17609_not n17648 ; n18284
g18029 and n17644_not n18284 ; n18285
g18030 and n17645_not n17648_not ; n18286
g18031 and n18285_not n18286_not ; n18287
g18032 and quotient[14] n18287_not ; n18288
g18033 and n17599_not n17886_not ; n18289
g18034 and n17885_not n18289 ; n18290
g18035 and n18288_not n18290_not ; n18291
g18036 and b[5]_not n18291_not ; n18292
g18037 and n17617_not n17643 ; n18293
g18038 and n17639_not n18293 ; n18294
g18039 and n17640_not n17643_not ; n18295
g18040 and n18294_not n18295_not ; n18296
g18041 and quotient[14] n18296_not ; n18297
g18042 and n17608_not n17886_not ; n18298
g18043 and n17885_not n18298 ; n18299
g18044 and n18297_not n18299_not ; n18300
g18045 and b[4]_not n18300_not ; n18301
g18046 and n17634_not n17638 ; n18302
g18047 and n17633_not n18302 ; n18303
g18048 and n17635_not n17638_not ; n18304
g18049 and n18303_not n18304_not ; n18305
g18050 and quotient[14] n18305_not ; n18306
g18051 and n17616_not n17886_not ; n18307
g18052 and n17885_not n18307 ; n18308
g18053 and n18306_not n18308_not ; n18309
g18054 and b[3]_not n18309_not ; n18310
g18055 and n17630_not n17632 ; n18311
g18056 and n17628_not n18311 ; n18312
g18057 and n17633_not n18312_not ; n18313
g18058 and quotient[14] n18313 ; n18314
g18059 and n17627_not n17886_not ; n18315
g18060 and n17885_not n18315 ; n18316
g18061 and n18314_not n18316_not ; n18317
g18062 and b[2]_not n18317_not ; n18318
g18063 and b[0] quotient[14] ; n18319
g18064 and a[14] n18319_not ; n18320
g18065 and n17632 quotient[14] ; n18321
g18066 and n18320_not n18321_not ; n18322
g18067 and b[1] n18322_not ; n18323
g18068 and b[1]_not n18321_not ; n18324
g18069 and n18320_not n18324 ; n18325
g18070 and n18323_not n18325_not ; n18326
g18071 and a[13]_not b[0] ; n18327
g18072 and n18326_not n18327_not ; n18328
g18073 and b[1]_not n18322_not ; n18329
g18074 and n18328_not n18329_not ; n18330
g18075 and b[2] n18316_not ; n18331
g18076 and n18314_not n18331 ; n18332
g18077 and n18318_not n18332_not ; n18333
g18078 and n18330_not n18333 ; n18334
g18079 and n18318_not n18334_not ; n18335
g18080 and b[3] n18308_not ; n18336
g18081 and n18306_not n18336 ; n18337
g18082 and n18310_not n18337_not ; n18338
g18083 and n18335_not n18338 ; n18339
g18084 and n18310_not n18339_not ; n18340
g18085 and b[4] n18299_not ; n18341
g18086 and n18297_not n18341 ; n18342
g18087 and n18301_not n18342_not ; n18343
g18088 and n18340_not n18343 ; n18344
g18089 and n18301_not n18344_not ; n18345
g18090 and b[5] n18290_not ; n18346
g18091 and n18288_not n18346 ; n18347
g18092 and n18292_not n18347_not ; n18348
g18093 and n18345_not n18348 ; n18349
g18094 and n18292_not n18349_not ; n18350
g18095 and b[6] n18281_not ; n18351
g18096 and n18279_not n18351 ; n18352
g18097 and n18283_not n18352_not ; n18353
g18098 and n18350_not n18353 ; n18354
g18099 and n18283_not n18354_not ; n18355
g18100 and b[7] n18272_not ; n18356
g18101 and n18270_not n18356 ; n18357
g18102 and n18274_not n18357_not ; n18358
g18103 and n18355_not n18358 ; n18359
g18104 and n18274_not n18359_not ; n18360
g18105 and b[8] n18263_not ; n18361
g18106 and n18261_not n18361 ; n18362
g18107 and n18265_not n18362_not ; n18363
g18108 and n18360_not n18363 ; n18364
g18109 and n18265_not n18364_not ; n18365
g18110 and b[9] n18254_not ; n18366
g18111 and n18252_not n18366 ; n18367
g18112 and n18256_not n18367_not ; n18368
g18113 and n18365_not n18368 ; n18369
g18114 and n18256_not n18369_not ; n18370
g18115 and b[10] n18245_not ; n18371
g18116 and n18243_not n18371 ; n18372
g18117 and n18247_not n18372_not ; n18373
g18118 and n18370_not n18373 ; n18374
g18119 and n18247_not n18374_not ; n18375
g18120 and b[11] n18236_not ; n18376
g18121 and n18234_not n18376 ; n18377
g18122 and n18238_not n18377_not ; n18378
g18123 and n18375_not n18378 ; n18379
g18124 and n18238_not n18379_not ; n18380
g18125 and b[12] n18227_not ; n18381
g18126 and n18225_not n18381 ; n18382
g18127 and n18229_not n18382_not ; n18383
g18128 and n18380_not n18383 ; n18384
g18129 and n18229_not n18384_not ; n18385
g18130 and b[13] n18218_not ; n18386
g18131 and n18216_not n18386 ; n18387
g18132 and n18220_not n18387_not ; n18388
g18133 and n18385_not n18388 ; n18389
g18134 and n18220_not n18389_not ; n18390
g18135 and b[14] n18209_not ; n18391
g18136 and n18207_not n18391 ; n18392
g18137 and n18211_not n18392_not ; n18393
g18138 and n18390_not n18393 ; n18394
g18139 and n18211_not n18394_not ; n18395
g18140 and b[15] n18200_not ; n18396
g18141 and n18198_not n18396 ; n18397
g18142 and n18202_not n18397_not ; n18398
g18143 and n18395_not n18398 ; n18399
g18144 and n18202_not n18399_not ; n18400
g18145 and b[16] n18191_not ; n18401
g18146 and n18189_not n18401 ; n18402
g18147 and n18193_not n18402_not ; n18403
g18148 and n18400_not n18403 ; n18404
g18149 and n18193_not n18404_not ; n18405
g18150 and b[17] n18182_not ; n18406
g18151 and n18180_not n18406 ; n18407
g18152 and n18184_not n18407_not ; n18408
g18153 and n18405_not n18408 ; n18409
g18154 and n18184_not n18409_not ; n18410
g18155 and b[18] n18173_not ; n18411
g18156 and n18171_not n18411 ; n18412
g18157 and n18175_not n18412_not ; n18413
g18158 and n18410_not n18413 ; n18414
g18159 and n18175_not n18414_not ; n18415
g18160 and b[19] n18164_not ; n18416
g18161 and n18162_not n18416 ; n18417
g18162 and n18166_not n18417_not ; n18418
g18163 and n18415_not n18418 ; n18419
g18164 and n18166_not n18419_not ; n18420
g18165 and b[20] n18155_not ; n18421
g18166 and n18153_not n18421 ; n18422
g18167 and n18157_not n18422_not ; n18423
g18168 and n18420_not n18423 ; n18424
g18169 and n18157_not n18424_not ; n18425
g18170 and b[21] n18146_not ; n18426
g18171 and n18144_not n18426 ; n18427
g18172 and n18148_not n18427_not ; n18428
g18173 and n18425_not n18428 ; n18429
g18174 and n18148_not n18429_not ; n18430
g18175 and b[22] n18137_not ; n18431
g18176 and n18135_not n18431 ; n18432
g18177 and n18139_not n18432_not ; n18433
g18178 and n18430_not n18433 ; n18434
g18179 and n18139_not n18434_not ; n18435
g18180 and b[23] n18128_not ; n18436
g18181 and n18126_not n18436 ; n18437
g18182 and n18130_not n18437_not ; n18438
g18183 and n18435_not n18438 ; n18439
g18184 and n18130_not n18439_not ; n18440
g18185 and b[24] n18119_not ; n18441
g18186 and n18117_not n18441 ; n18442
g18187 and n18121_not n18442_not ; n18443
g18188 and n18440_not n18443 ; n18444
g18189 and n18121_not n18444_not ; n18445
g18190 and b[25] n18110_not ; n18446
g18191 and n18108_not n18446 ; n18447
g18192 and n18112_not n18447_not ; n18448
g18193 and n18445_not n18448 ; n18449
g18194 and n18112_not n18449_not ; n18450
g18195 and b[26] n18101_not ; n18451
g18196 and n18099_not n18451 ; n18452
g18197 and n18103_not n18452_not ; n18453
g18198 and n18450_not n18453 ; n18454
g18199 and n18103_not n18454_not ; n18455
g18200 and b[27] n18092_not ; n18456
g18201 and n18090_not n18456 ; n18457
g18202 and n18094_not n18457_not ; n18458
g18203 and n18455_not n18458 ; n18459
g18204 and n18094_not n18459_not ; n18460
g18205 and b[28] n18083_not ; n18461
g18206 and n18081_not n18461 ; n18462
g18207 and n18085_not n18462_not ; n18463
g18208 and n18460_not n18463 ; n18464
g18209 and n18085_not n18464_not ; n18465
g18210 and b[29] n18074_not ; n18466
g18211 and n18072_not n18466 ; n18467
g18212 and n18076_not n18467_not ; n18468
g18213 and n18465_not n18468 ; n18469
g18214 and n18076_not n18469_not ; n18470
g18215 and b[30] n18065_not ; n18471
g18216 and n18063_not n18471 ; n18472
g18217 and n18067_not n18472_not ; n18473
g18218 and n18470_not n18473 ; n18474
g18219 and n18067_not n18474_not ; n18475
g18220 and b[31] n18056_not ; n18476
g18221 and n18054_not n18476 ; n18477
g18222 and n18058_not n18477_not ; n18478
g18223 and n18475_not n18478 ; n18479
g18224 and n18058_not n18479_not ; n18480
g18225 and b[32] n18047_not ; n18481
g18226 and n18045_not n18481 ; n18482
g18227 and n18049_not n18482_not ; n18483
g18228 and n18480_not n18483 ; n18484
g18229 and n18049_not n18484_not ; n18485
g18230 and b[33] n18038_not ; n18486
g18231 and n18036_not n18486 ; n18487
g18232 and n18040_not n18487_not ; n18488
g18233 and n18485_not n18488 ; n18489
g18234 and n18040_not n18489_not ; n18490
g18235 and b[34] n18029_not ; n18491
g18236 and n18027_not n18491 ; n18492
g18237 and n18031_not n18492_not ; n18493
g18238 and n18490_not n18493 ; n18494
g18239 and n18031_not n18494_not ; n18495
g18240 and b[35] n18020_not ; n18496
g18241 and n18018_not n18496 ; n18497
g18242 and n18022_not n18497_not ; n18498
g18243 and n18495_not n18498 ; n18499
g18244 and n18022_not n18499_not ; n18500
g18245 and b[36] n18011_not ; n18501
g18246 and n18009_not n18501 ; n18502
g18247 and n18013_not n18502_not ; n18503
g18248 and n18500_not n18503 ; n18504
g18249 and n18013_not n18504_not ; n18505
g18250 and b[37] n18002_not ; n18506
g18251 and n18000_not n18506 ; n18507
g18252 and n18004_not n18507_not ; n18508
g18253 and n18505_not n18508 ; n18509
g18254 and n18004_not n18509_not ; n18510
g18255 and b[38] n17993_not ; n18511
g18256 and n17991_not n18511 ; n18512
g18257 and n17995_not n18512_not ; n18513
g18258 and n18510_not n18513 ; n18514
g18259 and n17995_not n18514_not ; n18515
g18260 and b[39] n17984_not ; n18516
g18261 and n17982_not n18516 ; n18517
g18262 and n17986_not n18517_not ; n18518
g18263 and n18515_not n18518 ; n18519
g18264 and n17986_not n18519_not ; n18520
g18265 and b[40] n17975_not ; n18521
g18266 and n17973_not n18521 ; n18522
g18267 and n17977_not n18522_not ; n18523
g18268 and n18520_not n18523 ; n18524
g18269 and n17977_not n18524_not ; n18525
g18270 and b[41] n17966_not ; n18526
g18271 and n17964_not n18526 ; n18527
g18272 and n17968_not n18527_not ; n18528
g18273 and n18525_not n18528 ; n18529
g18274 and n17968_not n18529_not ; n18530
g18275 and b[42] n17957_not ; n18531
g18276 and n17955_not n18531 ; n18532
g18277 and n17959_not n18532_not ; n18533
g18278 and n18530_not n18533 ; n18534
g18279 and n17959_not n18534_not ; n18535
g18280 and b[43] n17948_not ; n18536
g18281 and n17946_not n18536 ; n18537
g18282 and n17950_not n18537_not ; n18538
g18283 and n18535_not n18538 ; n18539
g18284 and n17950_not n18539_not ; n18540
g18285 and b[44] n17939_not ; n18541
g18286 and n17937_not n18541 ; n18542
g18287 and n17941_not n18542_not ; n18543
g18288 and n18540_not n18543 ; n18544
g18289 and n17941_not n18544_not ; n18545
g18290 and b[45] n17930_not ; n18546
g18291 and n17928_not n18546 ; n18547
g18292 and n17932_not n18547_not ; n18548
g18293 and n18545_not n18548 ; n18549
g18294 and n17932_not n18549_not ; n18550
g18295 and b[46] n17921_not ; n18551
g18296 and n17919_not n18551 ; n18552
g18297 and n17923_not n18552_not ; n18553
g18298 and n18550_not n18553 ; n18554
g18299 and n17923_not n18554_not ; n18555
g18300 and b[47] n17912_not ; n18556
g18301 and n17910_not n18556 ; n18557
g18302 and n17914_not n18557_not ; n18558
g18303 and n18555_not n18558 ; n18559
g18304 and n17914_not n18559_not ; n18560
g18305 and b[48] n17903_not ; n18561
g18306 and n17901_not n18561 ; n18562
g18307 and n17905_not n18562_not ; n18563
g18308 and n18560_not n18563 ; n18564
g18309 and n17905_not n18564_not ; n18565
g18310 and b[49] n17894_not ; n18566
g18311 and n17892_not n18566 ; n18567
g18312 and n17896_not n18567_not ; n18568
g18313 and n18565_not n18568 ; n18569
g18314 and n17896_not n18569_not ; n18570
g18315 and n17204_not n17880_not ; n18571
g18316 and n17878_not n18571 ; n18572
g18317 and n17869_not n18572 ; n18573
g18318 and n17878_not n17880_not ; n18574
g18319 and n17870_not n18574_not ; n18575
g18320 and n18573_not n18575_not ; n18576
g18321 and quotient[14] n18576_not ; n18577
g18322 and n17877_not n17886_not ; n18578
g18323 and n17885_not n18578 ; n18579
g18324 and n18577_not n18579_not ; n18580
g18325 and b[50]_not n18580_not ; n18581
g18326 and b[50] n18579_not ; n18582
g18327 and n18577_not n18582 ; n18583
g18328 and n397 n399 ; n18584
g18329 and n407 n18584 ; n18585
g18330 and n18583_not n18585 ; n18586
g18331 and n18581_not n18586 ; n18587
g18332 and n18570_not n18587 ; n18588
g18333 and n17882 n18580_not ; n18589
g18334 and n18588_not n18589_not ; quotient[13]
g18335 and n17905_not n18568 ; n18591
g18336 and n18564_not n18591 ; n18592
g18337 and n18565_not n18568_not ; n18593
g18338 and n18592_not n18593_not ; n18594
g18339 and quotient[13] n18594_not ; n18595
g18340 and n17895_not n18589_not ; n18596
g18341 and n18588_not n18596 ; n18597
g18342 and n18595_not n18597_not ; n18598
g18343 and n17896_not n18583_not ; n18599
g18344 and n18581_not n18599 ; n18600
g18345 and n18569_not n18600 ; n18601
g18346 and n18581_not n18583_not ; n18602
g18347 and n18570_not n18602_not ; n18603
g18348 and n18601_not n18603_not ; n18604
g18349 and quotient[13] n18604_not ; n18605
g18350 and n18580_not n18589_not ; n18606
g18351 and n18588_not n18606 ; n18607
g18352 and n18605_not n18607_not ; n18608
g18353 and b[51]_not n18608_not ; n18609
g18354 and b[50]_not n18598_not ; n18610
g18355 and n17914_not n18563 ; n18611
g18356 and n18559_not n18611 ; n18612
g18357 and n18560_not n18563_not ; n18613
g18358 and n18612_not n18613_not ; n18614
g18359 and quotient[13] n18614_not ; n18615
g18360 and n17904_not n18589_not ; n18616
g18361 and n18588_not n18616 ; n18617
g18362 and n18615_not n18617_not ; n18618
g18363 and b[49]_not n18618_not ; n18619
g18364 and n17923_not n18558 ; n18620
g18365 and n18554_not n18620 ; n18621
g18366 and n18555_not n18558_not ; n18622
g18367 and n18621_not n18622_not ; n18623
g18368 and quotient[13] n18623_not ; n18624
g18369 and n17913_not n18589_not ; n18625
g18370 and n18588_not n18625 ; n18626
g18371 and n18624_not n18626_not ; n18627
g18372 and b[48]_not n18627_not ; n18628
g18373 and n17932_not n18553 ; n18629
g18374 and n18549_not n18629 ; n18630
g18375 and n18550_not n18553_not ; n18631
g18376 and n18630_not n18631_not ; n18632
g18377 and quotient[13] n18632_not ; n18633
g18378 and n17922_not n18589_not ; n18634
g18379 and n18588_not n18634 ; n18635
g18380 and n18633_not n18635_not ; n18636
g18381 and b[47]_not n18636_not ; n18637
g18382 and n17941_not n18548 ; n18638
g18383 and n18544_not n18638 ; n18639
g18384 and n18545_not n18548_not ; n18640
g18385 and n18639_not n18640_not ; n18641
g18386 and quotient[13] n18641_not ; n18642
g18387 and n17931_not n18589_not ; n18643
g18388 and n18588_not n18643 ; n18644
g18389 and n18642_not n18644_not ; n18645
g18390 and b[46]_not n18645_not ; n18646
g18391 and n17950_not n18543 ; n18647
g18392 and n18539_not n18647 ; n18648
g18393 and n18540_not n18543_not ; n18649
g18394 and n18648_not n18649_not ; n18650
g18395 and quotient[13] n18650_not ; n18651
g18396 and n17940_not n18589_not ; n18652
g18397 and n18588_not n18652 ; n18653
g18398 and n18651_not n18653_not ; n18654
g18399 and b[45]_not n18654_not ; n18655
g18400 and n17959_not n18538 ; n18656
g18401 and n18534_not n18656 ; n18657
g18402 and n18535_not n18538_not ; n18658
g18403 and n18657_not n18658_not ; n18659
g18404 and quotient[13] n18659_not ; n18660
g18405 and n17949_not n18589_not ; n18661
g18406 and n18588_not n18661 ; n18662
g18407 and n18660_not n18662_not ; n18663
g18408 and b[44]_not n18663_not ; n18664
g18409 and n17968_not n18533 ; n18665
g18410 and n18529_not n18665 ; n18666
g18411 and n18530_not n18533_not ; n18667
g18412 and n18666_not n18667_not ; n18668
g18413 and quotient[13] n18668_not ; n18669
g18414 and n17958_not n18589_not ; n18670
g18415 and n18588_not n18670 ; n18671
g18416 and n18669_not n18671_not ; n18672
g18417 and b[43]_not n18672_not ; n18673
g18418 and n17977_not n18528 ; n18674
g18419 and n18524_not n18674 ; n18675
g18420 and n18525_not n18528_not ; n18676
g18421 and n18675_not n18676_not ; n18677
g18422 and quotient[13] n18677_not ; n18678
g18423 and n17967_not n18589_not ; n18679
g18424 and n18588_not n18679 ; n18680
g18425 and n18678_not n18680_not ; n18681
g18426 and b[42]_not n18681_not ; n18682
g18427 and n17986_not n18523 ; n18683
g18428 and n18519_not n18683 ; n18684
g18429 and n18520_not n18523_not ; n18685
g18430 and n18684_not n18685_not ; n18686
g18431 and quotient[13] n18686_not ; n18687
g18432 and n17976_not n18589_not ; n18688
g18433 and n18588_not n18688 ; n18689
g18434 and n18687_not n18689_not ; n18690
g18435 and b[41]_not n18690_not ; n18691
g18436 and n17995_not n18518 ; n18692
g18437 and n18514_not n18692 ; n18693
g18438 and n18515_not n18518_not ; n18694
g18439 and n18693_not n18694_not ; n18695
g18440 and quotient[13] n18695_not ; n18696
g18441 and n17985_not n18589_not ; n18697
g18442 and n18588_not n18697 ; n18698
g18443 and n18696_not n18698_not ; n18699
g18444 and b[40]_not n18699_not ; n18700
g18445 and n18004_not n18513 ; n18701
g18446 and n18509_not n18701 ; n18702
g18447 and n18510_not n18513_not ; n18703
g18448 and n18702_not n18703_not ; n18704
g18449 and quotient[13] n18704_not ; n18705
g18450 and n17994_not n18589_not ; n18706
g18451 and n18588_not n18706 ; n18707
g18452 and n18705_not n18707_not ; n18708
g18453 and b[39]_not n18708_not ; n18709
g18454 and n18013_not n18508 ; n18710
g18455 and n18504_not n18710 ; n18711
g18456 and n18505_not n18508_not ; n18712
g18457 and n18711_not n18712_not ; n18713
g18458 and quotient[13] n18713_not ; n18714
g18459 and n18003_not n18589_not ; n18715
g18460 and n18588_not n18715 ; n18716
g18461 and n18714_not n18716_not ; n18717
g18462 and b[38]_not n18717_not ; n18718
g18463 and n18022_not n18503 ; n18719
g18464 and n18499_not n18719 ; n18720
g18465 and n18500_not n18503_not ; n18721
g18466 and n18720_not n18721_not ; n18722
g18467 and quotient[13] n18722_not ; n18723
g18468 and n18012_not n18589_not ; n18724
g18469 and n18588_not n18724 ; n18725
g18470 and n18723_not n18725_not ; n18726
g18471 and b[37]_not n18726_not ; n18727
g18472 and n18031_not n18498 ; n18728
g18473 and n18494_not n18728 ; n18729
g18474 and n18495_not n18498_not ; n18730
g18475 and n18729_not n18730_not ; n18731
g18476 and quotient[13] n18731_not ; n18732
g18477 and n18021_not n18589_not ; n18733
g18478 and n18588_not n18733 ; n18734
g18479 and n18732_not n18734_not ; n18735
g18480 and b[36]_not n18735_not ; n18736
g18481 and n18040_not n18493 ; n18737
g18482 and n18489_not n18737 ; n18738
g18483 and n18490_not n18493_not ; n18739
g18484 and n18738_not n18739_not ; n18740
g18485 and quotient[13] n18740_not ; n18741
g18486 and n18030_not n18589_not ; n18742
g18487 and n18588_not n18742 ; n18743
g18488 and n18741_not n18743_not ; n18744
g18489 and b[35]_not n18744_not ; n18745
g18490 and n18049_not n18488 ; n18746
g18491 and n18484_not n18746 ; n18747
g18492 and n18485_not n18488_not ; n18748
g18493 and n18747_not n18748_not ; n18749
g18494 and quotient[13] n18749_not ; n18750
g18495 and n18039_not n18589_not ; n18751
g18496 and n18588_not n18751 ; n18752
g18497 and n18750_not n18752_not ; n18753
g18498 and b[34]_not n18753_not ; n18754
g18499 and n18058_not n18483 ; n18755
g18500 and n18479_not n18755 ; n18756
g18501 and n18480_not n18483_not ; n18757
g18502 and n18756_not n18757_not ; n18758
g18503 and quotient[13] n18758_not ; n18759
g18504 and n18048_not n18589_not ; n18760
g18505 and n18588_not n18760 ; n18761
g18506 and n18759_not n18761_not ; n18762
g18507 and b[33]_not n18762_not ; n18763
g18508 and n18067_not n18478 ; n18764
g18509 and n18474_not n18764 ; n18765
g18510 and n18475_not n18478_not ; n18766
g18511 and n18765_not n18766_not ; n18767
g18512 and quotient[13] n18767_not ; n18768
g18513 and n18057_not n18589_not ; n18769
g18514 and n18588_not n18769 ; n18770
g18515 and n18768_not n18770_not ; n18771
g18516 and b[32]_not n18771_not ; n18772
g18517 and n18076_not n18473 ; n18773
g18518 and n18469_not n18773 ; n18774
g18519 and n18470_not n18473_not ; n18775
g18520 and n18774_not n18775_not ; n18776
g18521 and quotient[13] n18776_not ; n18777
g18522 and n18066_not n18589_not ; n18778
g18523 and n18588_not n18778 ; n18779
g18524 and n18777_not n18779_not ; n18780
g18525 and b[31]_not n18780_not ; n18781
g18526 and n18085_not n18468 ; n18782
g18527 and n18464_not n18782 ; n18783
g18528 and n18465_not n18468_not ; n18784
g18529 and n18783_not n18784_not ; n18785
g18530 and quotient[13] n18785_not ; n18786
g18531 and n18075_not n18589_not ; n18787
g18532 and n18588_not n18787 ; n18788
g18533 and n18786_not n18788_not ; n18789
g18534 and b[30]_not n18789_not ; n18790
g18535 and n18094_not n18463 ; n18791
g18536 and n18459_not n18791 ; n18792
g18537 and n18460_not n18463_not ; n18793
g18538 and n18792_not n18793_not ; n18794
g18539 and quotient[13] n18794_not ; n18795
g18540 and n18084_not n18589_not ; n18796
g18541 and n18588_not n18796 ; n18797
g18542 and n18795_not n18797_not ; n18798
g18543 and b[29]_not n18798_not ; n18799
g18544 and n18103_not n18458 ; n18800
g18545 and n18454_not n18800 ; n18801
g18546 and n18455_not n18458_not ; n18802
g18547 and n18801_not n18802_not ; n18803
g18548 and quotient[13] n18803_not ; n18804
g18549 and n18093_not n18589_not ; n18805
g18550 and n18588_not n18805 ; n18806
g18551 and n18804_not n18806_not ; n18807
g18552 and b[28]_not n18807_not ; n18808
g18553 and n18112_not n18453 ; n18809
g18554 and n18449_not n18809 ; n18810
g18555 and n18450_not n18453_not ; n18811
g18556 and n18810_not n18811_not ; n18812
g18557 and quotient[13] n18812_not ; n18813
g18558 and n18102_not n18589_not ; n18814
g18559 and n18588_not n18814 ; n18815
g18560 and n18813_not n18815_not ; n18816
g18561 and b[27]_not n18816_not ; n18817
g18562 and n18121_not n18448 ; n18818
g18563 and n18444_not n18818 ; n18819
g18564 and n18445_not n18448_not ; n18820
g18565 and n18819_not n18820_not ; n18821
g18566 and quotient[13] n18821_not ; n18822
g18567 and n18111_not n18589_not ; n18823
g18568 and n18588_not n18823 ; n18824
g18569 and n18822_not n18824_not ; n18825
g18570 and b[26]_not n18825_not ; n18826
g18571 and n18130_not n18443 ; n18827
g18572 and n18439_not n18827 ; n18828
g18573 and n18440_not n18443_not ; n18829
g18574 and n18828_not n18829_not ; n18830
g18575 and quotient[13] n18830_not ; n18831
g18576 and n18120_not n18589_not ; n18832
g18577 and n18588_not n18832 ; n18833
g18578 and n18831_not n18833_not ; n18834
g18579 and b[25]_not n18834_not ; n18835
g18580 and n18139_not n18438 ; n18836
g18581 and n18434_not n18836 ; n18837
g18582 and n18435_not n18438_not ; n18838
g18583 and n18837_not n18838_not ; n18839
g18584 and quotient[13] n18839_not ; n18840
g18585 and n18129_not n18589_not ; n18841
g18586 and n18588_not n18841 ; n18842
g18587 and n18840_not n18842_not ; n18843
g18588 and b[24]_not n18843_not ; n18844
g18589 and n18148_not n18433 ; n18845
g18590 and n18429_not n18845 ; n18846
g18591 and n18430_not n18433_not ; n18847
g18592 and n18846_not n18847_not ; n18848
g18593 and quotient[13] n18848_not ; n18849
g18594 and n18138_not n18589_not ; n18850
g18595 and n18588_not n18850 ; n18851
g18596 and n18849_not n18851_not ; n18852
g18597 and b[23]_not n18852_not ; n18853
g18598 and n18157_not n18428 ; n18854
g18599 and n18424_not n18854 ; n18855
g18600 and n18425_not n18428_not ; n18856
g18601 and n18855_not n18856_not ; n18857
g18602 and quotient[13] n18857_not ; n18858
g18603 and n18147_not n18589_not ; n18859
g18604 and n18588_not n18859 ; n18860
g18605 and n18858_not n18860_not ; n18861
g18606 and b[22]_not n18861_not ; n18862
g18607 and n18166_not n18423 ; n18863
g18608 and n18419_not n18863 ; n18864
g18609 and n18420_not n18423_not ; n18865
g18610 and n18864_not n18865_not ; n18866
g18611 and quotient[13] n18866_not ; n18867
g18612 and n18156_not n18589_not ; n18868
g18613 and n18588_not n18868 ; n18869
g18614 and n18867_not n18869_not ; n18870
g18615 and b[21]_not n18870_not ; n18871
g18616 and n18175_not n18418 ; n18872
g18617 and n18414_not n18872 ; n18873
g18618 and n18415_not n18418_not ; n18874
g18619 and n18873_not n18874_not ; n18875
g18620 and quotient[13] n18875_not ; n18876
g18621 and n18165_not n18589_not ; n18877
g18622 and n18588_not n18877 ; n18878
g18623 and n18876_not n18878_not ; n18879
g18624 and b[20]_not n18879_not ; n18880
g18625 and n18184_not n18413 ; n18881
g18626 and n18409_not n18881 ; n18882
g18627 and n18410_not n18413_not ; n18883
g18628 and n18882_not n18883_not ; n18884
g18629 and quotient[13] n18884_not ; n18885
g18630 and n18174_not n18589_not ; n18886
g18631 and n18588_not n18886 ; n18887
g18632 and n18885_not n18887_not ; n18888
g18633 and b[19]_not n18888_not ; n18889
g18634 and n18193_not n18408 ; n18890
g18635 and n18404_not n18890 ; n18891
g18636 and n18405_not n18408_not ; n18892
g18637 and n18891_not n18892_not ; n18893
g18638 and quotient[13] n18893_not ; n18894
g18639 and n18183_not n18589_not ; n18895
g18640 and n18588_not n18895 ; n18896
g18641 and n18894_not n18896_not ; n18897
g18642 and b[18]_not n18897_not ; n18898
g18643 and n18202_not n18403 ; n18899
g18644 and n18399_not n18899 ; n18900
g18645 and n18400_not n18403_not ; n18901
g18646 and n18900_not n18901_not ; n18902
g18647 and quotient[13] n18902_not ; n18903
g18648 and n18192_not n18589_not ; n18904
g18649 and n18588_not n18904 ; n18905
g18650 and n18903_not n18905_not ; n18906
g18651 and b[17]_not n18906_not ; n18907
g18652 and n18211_not n18398 ; n18908
g18653 and n18394_not n18908 ; n18909
g18654 and n18395_not n18398_not ; n18910
g18655 and n18909_not n18910_not ; n18911
g18656 and quotient[13] n18911_not ; n18912
g18657 and n18201_not n18589_not ; n18913
g18658 and n18588_not n18913 ; n18914
g18659 and n18912_not n18914_not ; n18915
g18660 and b[16]_not n18915_not ; n18916
g18661 and n18220_not n18393 ; n18917
g18662 and n18389_not n18917 ; n18918
g18663 and n18390_not n18393_not ; n18919
g18664 and n18918_not n18919_not ; n18920
g18665 and quotient[13] n18920_not ; n18921
g18666 and n18210_not n18589_not ; n18922
g18667 and n18588_not n18922 ; n18923
g18668 and n18921_not n18923_not ; n18924
g18669 and b[15]_not n18924_not ; n18925
g18670 and n18229_not n18388 ; n18926
g18671 and n18384_not n18926 ; n18927
g18672 and n18385_not n18388_not ; n18928
g18673 and n18927_not n18928_not ; n18929
g18674 and quotient[13] n18929_not ; n18930
g18675 and n18219_not n18589_not ; n18931
g18676 and n18588_not n18931 ; n18932
g18677 and n18930_not n18932_not ; n18933
g18678 and b[14]_not n18933_not ; n18934
g18679 and n18238_not n18383 ; n18935
g18680 and n18379_not n18935 ; n18936
g18681 and n18380_not n18383_not ; n18937
g18682 and n18936_not n18937_not ; n18938
g18683 and quotient[13] n18938_not ; n18939
g18684 and n18228_not n18589_not ; n18940
g18685 and n18588_not n18940 ; n18941
g18686 and n18939_not n18941_not ; n18942
g18687 and b[13]_not n18942_not ; n18943
g18688 and n18247_not n18378 ; n18944
g18689 and n18374_not n18944 ; n18945
g18690 and n18375_not n18378_not ; n18946
g18691 and n18945_not n18946_not ; n18947
g18692 and quotient[13] n18947_not ; n18948
g18693 and n18237_not n18589_not ; n18949
g18694 and n18588_not n18949 ; n18950
g18695 and n18948_not n18950_not ; n18951
g18696 and b[12]_not n18951_not ; n18952
g18697 and n18256_not n18373 ; n18953
g18698 and n18369_not n18953 ; n18954
g18699 and n18370_not n18373_not ; n18955
g18700 and n18954_not n18955_not ; n18956
g18701 and quotient[13] n18956_not ; n18957
g18702 and n18246_not n18589_not ; n18958
g18703 and n18588_not n18958 ; n18959
g18704 and n18957_not n18959_not ; n18960
g18705 and b[11]_not n18960_not ; n18961
g18706 and n18265_not n18368 ; n18962
g18707 and n18364_not n18962 ; n18963
g18708 and n18365_not n18368_not ; n18964
g18709 and n18963_not n18964_not ; n18965
g18710 and quotient[13] n18965_not ; n18966
g18711 and n18255_not n18589_not ; n18967
g18712 and n18588_not n18967 ; n18968
g18713 and n18966_not n18968_not ; n18969
g18714 and b[10]_not n18969_not ; n18970
g18715 and n18274_not n18363 ; n18971
g18716 and n18359_not n18971 ; n18972
g18717 and n18360_not n18363_not ; n18973
g18718 and n18972_not n18973_not ; n18974
g18719 and quotient[13] n18974_not ; n18975
g18720 and n18264_not n18589_not ; n18976
g18721 and n18588_not n18976 ; n18977
g18722 and n18975_not n18977_not ; n18978
g18723 and b[9]_not n18978_not ; n18979
g18724 and n18283_not n18358 ; n18980
g18725 and n18354_not n18980 ; n18981
g18726 and n18355_not n18358_not ; n18982
g18727 and n18981_not n18982_not ; n18983
g18728 and quotient[13] n18983_not ; n18984
g18729 and n18273_not n18589_not ; n18985
g18730 and n18588_not n18985 ; n18986
g18731 and n18984_not n18986_not ; n18987
g18732 and b[8]_not n18987_not ; n18988
g18733 and n18292_not n18353 ; n18989
g18734 and n18349_not n18989 ; n18990
g18735 and n18350_not n18353_not ; n18991
g18736 and n18990_not n18991_not ; n18992
g18737 and quotient[13] n18992_not ; n18993
g18738 and n18282_not n18589_not ; n18994
g18739 and n18588_not n18994 ; n18995
g18740 and n18993_not n18995_not ; n18996
g18741 and b[7]_not n18996_not ; n18997
g18742 and n18301_not n18348 ; n18998
g18743 and n18344_not n18998 ; n18999
g18744 and n18345_not n18348_not ; n19000
g18745 and n18999_not n19000_not ; n19001
g18746 and quotient[13] n19001_not ; n19002
g18747 and n18291_not n18589_not ; n19003
g18748 and n18588_not n19003 ; n19004
g18749 and n19002_not n19004_not ; n19005
g18750 and b[6]_not n19005_not ; n19006
g18751 and n18310_not n18343 ; n19007
g18752 and n18339_not n19007 ; n19008
g18753 and n18340_not n18343_not ; n19009
g18754 and n19008_not n19009_not ; n19010
g18755 and quotient[13] n19010_not ; n19011
g18756 and n18300_not n18589_not ; n19012
g18757 and n18588_not n19012 ; n19013
g18758 and n19011_not n19013_not ; n19014
g18759 and b[5]_not n19014_not ; n19015
g18760 and n18318_not n18338 ; n19016
g18761 and n18334_not n19016 ; n19017
g18762 and n18335_not n18338_not ; n19018
g18763 and n19017_not n19018_not ; n19019
g18764 and quotient[13] n19019_not ; n19020
g18765 and n18309_not n18589_not ; n19021
g18766 and n18588_not n19021 ; n19022
g18767 and n19020_not n19022_not ; n19023
g18768 and b[4]_not n19023_not ; n19024
g18769 and n18329_not n18333 ; n19025
g18770 and n18328_not n19025 ; n19026
g18771 and n18330_not n18333_not ; n19027
g18772 and n19026_not n19027_not ; n19028
g18773 and quotient[13] n19028_not ; n19029
g18774 and n18317_not n18589_not ; n19030
g18775 and n18588_not n19030 ; n19031
g18776 and n19029_not n19031_not ; n19032
g18777 and b[3]_not n19032_not ; n19033
g18778 and n18325_not n18327 ; n19034
g18779 and n18323_not n19034 ; n19035
g18780 and n18328_not n19035_not ; n19036
g18781 and quotient[13] n19036 ; n19037
g18782 and n18322_not n18589_not ; n19038
g18783 and n18588_not n19038 ; n19039
g18784 and n19037_not n19039_not ; n19040
g18785 and b[2]_not n19040_not ; n19041
g18786 and b[0] quotient[13] ; n19042
g18787 and a[13] n19042_not ; n19043
g18788 and n18327 quotient[13] ; n19044
g18789 and n19043_not n19044_not ; n19045
g18790 and b[1] n19045_not ; n19046
g18791 and b[1]_not n19044_not ; n19047
g18792 and n19043_not n19047 ; n19048
g18793 and n19046_not n19048_not ; n19049
g18794 and a[12]_not b[0] ; n19050
g18795 and n19049_not n19050_not ; n19051
g18796 and b[1]_not n19045_not ; n19052
g18797 and n19051_not n19052_not ; n19053
g18798 and b[2] n19039_not ; n19054
g18799 and n19037_not n19054 ; n19055
g18800 and n19041_not n19055_not ; n19056
g18801 and n19053_not n19056 ; n19057
g18802 and n19041_not n19057_not ; n19058
g18803 and b[3] n19031_not ; n19059
g18804 and n19029_not n19059 ; n19060
g18805 and n19033_not n19060_not ; n19061
g18806 and n19058_not n19061 ; n19062
g18807 and n19033_not n19062_not ; n19063
g18808 and b[4] n19022_not ; n19064
g18809 and n19020_not n19064 ; n19065
g18810 and n19024_not n19065_not ; n19066
g18811 and n19063_not n19066 ; n19067
g18812 and n19024_not n19067_not ; n19068
g18813 and b[5] n19013_not ; n19069
g18814 and n19011_not n19069 ; n19070
g18815 and n19015_not n19070_not ; n19071
g18816 and n19068_not n19071 ; n19072
g18817 and n19015_not n19072_not ; n19073
g18818 and b[6] n19004_not ; n19074
g18819 and n19002_not n19074 ; n19075
g18820 and n19006_not n19075_not ; n19076
g18821 and n19073_not n19076 ; n19077
g18822 and n19006_not n19077_not ; n19078
g18823 and b[7] n18995_not ; n19079
g18824 and n18993_not n19079 ; n19080
g18825 and n18997_not n19080_not ; n19081
g18826 and n19078_not n19081 ; n19082
g18827 and n18997_not n19082_not ; n19083
g18828 and b[8] n18986_not ; n19084
g18829 and n18984_not n19084 ; n19085
g18830 and n18988_not n19085_not ; n19086
g18831 and n19083_not n19086 ; n19087
g18832 and n18988_not n19087_not ; n19088
g18833 and b[9] n18977_not ; n19089
g18834 and n18975_not n19089 ; n19090
g18835 and n18979_not n19090_not ; n19091
g18836 and n19088_not n19091 ; n19092
g18837 and n18979_not n19092_not ; n19093
g18838 and b[10] n18968_not ; n19094
g18839 and n18966_not n19094 ; n19095
g18840 and n18970_not n19095_not ; n19096
g18841 and n19093_not n19096 ; n19097
g18842 and n18970_not n19097_not ; n19098
g18843 and b[11] n18959_not ; n19099
g18844 and n18957_not n19099 ; n19100
g18845 and n18961_not n19100_not ; n19101
g18846 and n19098_not n19101 ; n19102
g18847 and n18961_not n19102_not ; n19103
g18848 and b[12] n18950_not ; n19104
g18849 and n18948_not n19104 ; n19105
g18850 and n18952_not n19105_not ; n19106
g18851 and n19103_not n19106 ; n19107
g18852 and n18952_not n19107_not ; n19108
g18853 and b[13] n18941_not ; n19109
g18854 and n18939_not n19109 ; n19110
g18855 and n18943_not n19110_not ; n19111
g18856 and n19108_not n19111 ; n19112
g18857 and n18943_not n19112_not ; n19113
g18858 and b[14] n18932_not ; n19114
g18859 and n18930_not n19114 ; n19115
g18860 and n18934_not n19115_not ; n19116
g18861 and n19113_not n19116 ; n19117
g18862 and n18934_not n19117_not ; n19118
g18863 and b[15] n18923_not ; n19119
g18864 and n18921_not n19119 ; n19120
g18865 and n18925_not n19120_not ; n19121
g18866 and n19118_not n19121 ; n19122
g18867 and n18925_not n19122_not ; n19123
g18868 and b[16] n18914_not ; n19124
g18869 and n18912_not n19124 ; n19125
g18870 and n18916_not n19125_not ; n19126
g18871 and n19123_not n19126 ; n19127
g18872 and n18916_not n19127_not ; n19128
g18873 and b[17] n18905_not ; n19129
g18874 and n18903_not n19129 ; n19130
g18875 and n18907_not n19130_not ; n19131
g18876 and n19128_not n19131 ; n19132
g18877 and n18907_not n19132_not ; n19133
g18878 and b[18] n18896_not ; n19134
g18879 and n18894_not n19134 ; n19135
g18880 and n18898_not n19135_not ; n19136
g18881 and n19133_not n19136 ; n19137
g18882 and n18898_not n19137_not ; n19138
g18883 and b[19] n18887_not ; n19139
g18884 and n18885_not n19139 ; n19140
g18885 and n18889_not n19140_not ; n19141
g18886 and n19138_not n19141 ; n19142
g18887 and n18889_not n19142_not ; n19143
g18888 and b[20] n18878_not ; n19144
g18889 and n18876_not n19144 ; n19145
g18890 and n18880_not n19145_not ; n19146
g18891 and n19143_not n19146 ; n19147
g18892 and n18880_not n19147_not ; n19148
g18893 and b[21] n18869_not ; n19149
g18894 and n18867_not n19149 ; n19150
g18895 and n18871_not n19150_not ; n19151
g18896 and n19148_not n19151 ; n19152
g18897 and n18871_not n19152_not ; n19153
g18898 and b[22] n18860_not ; n19154
g18899 and n18858_not n19154 ; n19155
g18900 and n18862_not n19155_not ; n19156
g18901 and n19153_not n19156 ; n19157
g18902 and n18862_not n19157_not ; n19158
g18903 and b[23] n18851_not ; n19159
g18904 and n18849_not n19159 ; n19160
g18905 and n18853_not n19160_not ; n19161
g18906 and n19158_not n19161 ; n19162
g18907 and n18853_not n19162_not ; n19163
g18908 and b[24] n18842_not ; n19164
g18909 and n18840_not n19164 ; n19165
g18910 and n18844_not n19165_not ; n19166
g18911 and n19163_not n19166 ; n19167
g18912 and n18844_not n19167_not ; n19168
g18913 and b[25] n18833_not ; n19169
g18914 and n18831_not n19169 ; n19170
g18915 and n18835_not n19170_not ; n19171
g18916 and n19168_not n19171 ; n19172
g18917 and n18835_not n19172_not ; n19173
g18918 and b[26] n18824_not ; n19174
g18919 and n18822_not n19174 ; n19175
g18920 and n18826_not n19175_not ; n19176
g18921 and n19173_not n19176 ; n19177
g18922 and n18826_not n19177_not ; n19178
g18923 and b[27] n18815_not ; n19179
g18924 and n18813_not n19179 ; n19180
g18925 and n18817_not n19180_not ; n19181
g18926 and n19178_not n19181 ; n19182
g18927 and n18817_not n19182_not ; n19183
g18928 and b[28] n18806_not ; n19184
g18929 and n18804_not n19184 ; n19185
g18930 and n18808_not n19185_not ; n19186
g18931 and n19183_not n19186 ; n19187
g18932 and n18808_not n19187_not ; n19188
g18933 and b[29] n18797_not ; n19189
g18934 and n18795_not n19189 ; n19190
g18935 and n18799_not n19190_not ; n19191
g18936 and n19188_not n19191 ; n19192
g18937 and n18799_not n19192_not ; n19193
g18938 and b[30] n18788_not ; n19194
g18939 and n18786_not n19194 ; n19195
g18940 and n18790_not n19195_not ; n19196
g18941 and n19193_not n19196 ; n19197
g18942 and n18790_not n19197_not ; n19198
g18943 and b[31] n18779_not ; n19199
g18944 and n18777_not n19199 ; n19200
g18945 and n18781_not n19200_not ; n19201
g18946 and n19198_not n19201 ; n19202
g18947 and n18781_not n19202_not ; n19203
g18948 and b[32] n18770_not ; n19204
g18949 and n18768_not n19204 ; n19205
g18950 and n18772_not n19205_not ; n19206
g18951 and n19203_not n19206 ; n19207
g18952 and n18772_not n19207_not ; n19208
g18953 and b[33] n18761_not ; n19209
g18954 and n18759_not n19209 ; n19210
g18955 and n18763_not n19210_not ; n19211
g18956 and n19208_not n19211 ; n19212
g18957 and n18763_not n19212_not ; n19213
g18958 and b[34] n18752_not ; n19214
g18959 and n18750_not n19214 ; n19215
g18960 and n18754_not n19215_not ; n19216
g18961 and n19213_not n19216 ; n19217
g18962 and n18754_not n19217_not ; n19218
g18963 and b[35] n18743_not ; n19219
g18964 and n18741_not n19219 ; n19220
g18965 and n18745_not n19220_not ; n19221
g18966 and n19218_not n19221 ; n19222
g18967 and n18745_not n19222_not ; n19223
g18968 and b[36] n18734_not ; n19224
g18969 and n18732_not n19224 ; n19225
g18970 and n18736_not n19225_not ; n19226
g18971 and n19223_not n19226 ; n19227
g18972 and n18736_not n19227_not ; n19228
g18973 and b[37] n18725_not ; n19229
g18974 and n18723_not n19229 ; n19230
g18975 and n18727_not n19230_not ; n19231
g18976 and n19228_not n19231 ; n19232
g18977 and n18727_not n19232_not ; n19233
g18978 and b[38] n18716_not ; n19234
g18979 and n18714_not n19234 ; n19235
g18980 and n18718_not n19235_not ; n19236
g18981 and n19233_not n19236 ; n19237
g18982 and n18718_not n19237_not ; n19238
g18983 and b[39] n18707_not ; n19239
g18984 and n18705_not n19239 ; n19240
g18985 and n18709_not n19240_not ; n19241
g18986 and n19238_not n19241 ; n19242
g18987 and n18709_not n19242_not ; n19243
g18988 and b[40] n18698_not ; n19244
g18989 and n18696_not n19244 ; n19245
g18990 and n18700_not n19245_not ; n19246
g18991 and n19243_not n19246 ; n19247
g18992 and n18700_not n19247_not ; n19248
g18993 and b[41] n18689_not ; n19249
g18994 and n18687_not n19249 ; n19250
g18995 and n18691_not n19250_not ; n19251
g18996 and n19248_not n19251 ; n19252
g18997 and n18691_not n19252_not ; n19253
g18998 and b[42] n18680_not ; n19254
g18999 and n18678_not n19254 ; n19255
g19000 and n18682_not n19255_not ; n19256
g19001 and n19253_not n19256 ; n19257
g19002 and n18682_not n19257_not ; n19258
g19003 and b[43] n18671_not ; n19259
g19004 and n18669_not n19259 ; n19260
g19005 and n18673_not n19260_not ; n19261
g19006 and n19258_not n19261 ; n19262
g19007 and n18673_not n19262_not ; n19263
g19008 and b[44] n18662_not ; n19264
g19009 and n18660_not n19264 ; n19265
g19010 and n18664_not n19265_not ; n19266
g19011 and n19263_not n19266 ; n19267
g19012 and n18664_not n19267_not ; n19268
g19013 and b[45] n18653_not ; n19269
g19014 and n18651_not n19269 ; n19270
g19015 and n18655_not n19270_not ; n19271
g19016 and n19268_not n19271 ; n19272
g19017 and n18655_not n19272_not ; n19273
g19018 and b[46] n18644_not ; n19274
g19019 and n18642_not n19274 ; n19275
g19020 and n18646_not n19275_not ; n19276
g19021 and n19273_not n19276 ; n19277
g19022 and n18646_not n19277_not ; n19278
g19023 and b[47] n18635_not ; n19279
g19024 and n18633_not n19279 ; n19280
g19025 and n18637_not n19280_not ; n19281
g19026 and n19278_not n19281 ; n19282
g19027 and n18637_not n19282_not ; n19283
g19028 and b[48] n18626_not ; n19284
g19029 and n18624_not n19284 ; n19285
g19030 and n18628_not n19285_not ; n19286
g19031 and n19283_not n19286 ; n19287
g19032 and n18628_not n19287_not ; n19288
g19033 and b[49] n18617_not ; n19289
g19034 and n18615_not n19289 ; n19290
g19035 and n18619_not n19290_not ; n19291
g19036 and n19288_not n19291 ; n19292
g19037 and n18619_not n19292_not ; n19293
g19038 and b[50] n18597_not ; n19294
g19039 and n18595_not n19294 ; n19295
g19040 and n18610_not n19295_not ; n19296
g19041 and n19293_not n19296 ; n19297
g19042 and n18610_not n19297_not ; n19298
g19043 and b[51] n18607_not ; n19299
g19044 and n18605_not n19299 ; n19300
g19045 and n18609_not n19300_not ; n19301
g19046 and n19298_not n19301 ; n19302
g19047 and n18609_not n19302_not ; n19303
g19048 and n288 n19303_not ; quotient[12]
g19049 and n18598_not quotient[12]_not ; n19305
g19050 and n18619_not n19296 ; n19306
g19051 and n19292_not n19306 ; n19307
g19052 and n19293_not n19296_not ; n19308
g19053 and n19307_not n19308_not ; n19309
g19054 and n288 n19309_not ; n19310
g19055 and n19303_not n19310 ; n19311
g19056 and n19305_not n19311_not ; n19312
g19057 and b[51]_not n19312_not ; n19313
g19058 and n18618_not quotient[12]_not ; n19314
g19059 and n18628_not n19291 ; n19315
g19060 and n19287_not n19315 ; n19316
g19061 and n19288_not n19291_not ; n19317
g19062 and n19316_not n19317_not ; n19318
g19063 and n288 n19318_not ; n19319
g19064 and n19303_not n19319 ; n19320
g19065 and n19314_not n19320_not ; n19321
g19066 and b[50]_not n19321_not ; n19322
g19067 and n18627_not quotient[12]_not ; n19323
g19068 and n18637_not n19286 ; n19324
g19069 and n19282_not n19324 ; n19325
g19070 and n19283_not n19286_not ; n19326
g19071 and n19325_not n19326_not ; n19327
g19072 and n288 n19327_not ; n19328
g19073 and n19303_not n19328 ; n19329
g19074 and n19323_not n19329_not ; n19330
g19075 and b[49]_not n19330_not ; n19331
g19076 and n18636_not quotient[12]_not ; n19332
g19077 and n18646_not n19281 ; n19333
g19078 and n19277_not n19333 ; n19334
g19079 and n19278_not n19281_not ; n19335
g19080 and n19334_not n19335_not ; n19336
g19081 and n288 n19336_not ; n19337
g19082 and n19303_not n19337 ; n19338
g19083 and n19332_not n19338_not ; n19339
g19084 and b[48]_not n19339_not ; n19340
g19085 and n18645_not quotient[12]_not ; n19341
g19086 and n18655_not n19276 ; n19342
g19087 and n19272_not n19342 ; n19343
g19088 and n19273_not n19276_not ; n19344
g19089 and n19343_not n19344_not ; n19345
g19090 and n288 n19345_not ; n19346
g19091 and n19303_not n19346 ; n19347
g19092 and n19341_not n19347_not ; n19348
g19093 and b[47]_not n19348_not ; n19349
g19094 and n18654_not quotient[12]_not ; n19350
g19095 and n18664_not n19271 ; n19351
g19096 and n19267_not n19351 ; n19352
g19097 and n19268_not n19271_not ; n19353
g19098 and n19352_not n19353_not ; n19354
g19099 and n288 n19354_not ; n19355
g19100 and n19303_not n19355 ; n19356
g19101 and n19350_not n19356_not ; n19357
g19102 and b[46]_not n19357_not ; n19358
g19103 and n18663_not quotient[12]_not ; n19359
g19104 and n18673_not n19266 ; n19360
g19105 and n19262_not n19360 ; n19361
g19106 and n19263_not n19266_not ; n19362
g19107 and n19361_not n19362_not ; n19363
g19108 and n288 n19363_not ; n19364
g19109 and n19303_not n19364 ; n19365
g19110 and n19359_not n19365_not ; n19366
g19111 and b[45]_not n19366_not ; n19367
g19112 and n18672_not quotient[12]_not ; n19368
g19113 and n18682_not n19261 ; n19369
g19114 and n19257_not n19369 ; n19370
g19115 and n19258_not n19261_not ; n19371
g19116 and n19370_not n19371_not ; n19372
g19117 and n288 n19372_not ; n19373
g19118 and n19303_not n19373 ; n19374
g19119 and n19368_not n19374_not ; n19375
g19120 and b[44]_not n19375_not ; n19376
g19121 and n18681_not quotient[12]_not ; n19377
g19122 and n18691_not n19256 ; n19378
g19123 and n19252_not n19378 ; n19379
g19124 and n19253_not n19256_not ; n19380
g19125 and n19379_not n19380_not ; n19381
g19126 and n288 n19381_not ; n19382
g19127 and n19303_not n19382 ; n19383
g19128 and n19377_not n19383_not ; n19384
g19129 and b[43]_not n19384_not ; n19385
g19130 and n18690_not quotient[12]_not ; n19386
g19131 and n18700_not n19251 ; n19387
g19132 and n19247_not n19387 ; n19388
g19133 and n19248_not n19251_not ; n19389
g19134 and n19388_not n19389_not ; n19390
g19135 and n288 n19390_not ; n19391
g19136 and n19303_not n19391 ; n19392
g19137 and n19386_not n19392_not ; n19393
g19138 and b[42]_not n19393_not ; n19394
g19139 and n18699_not quotient[12]_not ; n19395
g19140 and n18709_not n19246 ; n19396
g19141 and n19242_not n19396 ; n19397
g19142 and n19243_not n19246_not ; n19398
g19143 and n19397_not n19398_not ; n19399
g19144 and n288 n19399_not ; n19400
g19145 and n19303_not n19400 ; n19401
g19146 and n19395_not n19401_not ; n19402
g19147 and b[41]_not n19402_not ; n19403
g19148 and n18708_not quotient[12]_not ; n19404
g19149 and n18718_not n19241 ; n19405
g19150 and n19237_not n19405 ; n19406
g19151 and n19238_not n19241_not ; n19407
g19152 and n19406_not n19407_not ; n19408
g19153 and n288 n19408_not ; n19409
g19154 and n19303_not n19409 ; n19410
g19155 and n19404_not n19410_not ; n19411
g19156 and b[40]_not n19411_not ; n19412
g19157 and n18717_not quotient[12]_not ; n19413
g19158 and n18727_not n19236 ; n19414
g19159 and n19232_not n19414 ; n19415
g19160 and n19233_not n19236_not ; n19416
g19161 and n19415_not n19416_not ; n19417
g19162 and n288 n19417_not ; n19418
g19163 and n19303_not n19418 ; n19419
g19164 and n19413_not n19419_not ; n19420
g19165 and b[39]_not n19420_not ; n19421
g19166 and n18726_not quotient[12]_not ; n19422
g19167 and n18736_not n19231 ; n19423
g19168 and n19227_not n19423 ; n19424
g19169 and n19228_not n19231_not ; n19425
g19170 and n19424_not n19425_not ; n19426
g19171 and n288 n19426_not ; n19427
g19172 and n19303_not n19427 ; n19428
g19173 and n19422_not n19428_not ; n19429
g19174 and b[38]_not n19429_not ; n19430
g19175 and n18735_not quotient[12]_not ; n19431
g19176 and n18745_not n19226 ; n19432
g19177 and n19222_not n19432 ; n19433
g19178 and n19223_not n19226_not ; n19434
g19179 and n19433_not n19434_not ; n19435
g19180 and n288 n19435_not ; n19436
g19181 and n19303_not n19436 ; n19437
g19182 and n19431_not n19437_not ; n19438
g19183 and b[37]_not n19438_not ; n19439
g19184 and n18744_not quotient[12]_not ; n19440
g19185 and n18754_not n19221 ; n19441
g19186 and n19217_not n19441 ; n19442
g19187 and n19218_not n19221_not ; n19443
g19188 and n19442_not n19443_not ; n19444
g19189 and n288 n19444_not ; n19445
g19190 and n19303_not n19445 ; n19446
g19191 and n19440_not n19446_not ; n19447
g19192 and b[36]_not n19447_not ; n19448
g19193 and n18753_not quotient[12]_not ; n19449
g19194 and n18763_not n19216 ; n19450
g19195 and n19212_not n19450 ; n19451
g19196 and n19213_not n19216_not ; n19452
g19197 and n19451_not n19452_not ; n19453
g19198 and n288 n19453_not ; n19454
g19199 and n19303_not n19454 ; n19455
g19200 and n19449_not n19455_not ; n19456
g19201 and b[35]_not n19456_not ; n19457
g19202 and n18762_not quotient[12]_not ; n19458
g19203 and n18772_not n19211 ; n19459
g19204 and n19207_not n19459 ; n19460
g19205 and n19208_not n19211_not ; n19461
g19206 and n19460_not n19461_not ; n19462
g19207 and n288 n19462_not ; n19463
g19208 and n19303_not n19463 ; n19464
g19209 and n19458_not n19464_not ; n19465
g19210 and b[34]_not n19465_not ; n19466
g19211 and n18771_not quotient[12]_not ; n19467
g19212 and n18781_not n19206 ; n19468
g19213 and n19202_not n19468 ; n19469
g19214 and n19203_not n19206_not ; n19470
g19215 and n19469_not n19470_not ; n19471
g19216 and n288 n19471_not ; n19472
g19217 and n19303_not n19472 ; n19473
g19218 and n19467_not n19473_not ; n19474
g19219 and b[33]_not n19474_not ; n19475
g19220 and n18780_not quotient[12]_not ; n19476
g19221 and n18790_not n19201 ; n19477
g19222 and n19197_not n19477 ; n19478
g19223 and n19198_not n19201_not ; n19479
g19224 and n19478_not n19479_not ; n19480
g19225 and n288 n19480_not ; n19481
g19226 and n19303_not n19481 ; n19482
g19227 and n19476_not n19482_not ; n19483
g19228 and b[32]_not n19483_not ; n19484
g19229 and n18789_not quotient[12]_not ; n19485
g19230 and n18799_not n19196 ; n19486
g19231 and n19192_not n19486 ; n19487
g19232 and n19193_not n19196_not ; n19488
g19233 and n19487_not n19488_not ; n19489
g19234 and n288 n19489_not ; n19490
g19235 and n19303_not n19490 ; n19491
g19236 and n19485_not n19491_not ; n19492
g19237 and b[31]_not n19492_not ; n19493
g19238 and n18798_not quotient[12]_not ; n19494
g19239 and n18808_not n19191 ; n19495
g19240 and n19187_not n19495 ; n19496
g19241 and n19188_not n19191_not ; n19497
g19242 and n19496_not n19497_not ; n19498
g19243 and n288 n19498_not ; n19499
g19244 and n19303_not n19499 ; n19500
g19245 and n19494_not n19500_not ; n19501
g19246 and b[30]_not n19501_not ; n19502
g19247 and n18807_not quotient[12]_not ; n19503
g19248 and n18817_not n19186 ; n19504
g19249 and n19182_not n19504 ; n19505
g19250 and n19183_not n19186_not ; n19506
g19251 and n19505_not n19506_not ; n19507
g19252 and n288 n19507_not ; n19508
g19253 and n19303_not n19508 ; n19509
g19254 and n19503_not n19509_not ; n19510
g19255 and b[29]_not n19510_not ; n19511
g19256 and n18816_not quotient[12]_not ; n19512
g19257 and n18826_not n19181 ; n19513
g19258 and n19177_not n19513 ; n19514
g19259 and n19178_not n19181_not ; n19515
g19260 and n19514_not n19515_not ; n19516
g19261 and n288 n19516_not ; n19517
g19262 and n19303_not n19517 ; n19518
g19263 and n19512_not n19518_not ; n19519
g19264 and b[28]_not n19519_not ; n19520
g19265 and n18825_not quotient[12]_not ; n19521
g19266 and n18835_not n19176 ; n19522
g19267 and n19172_not n19522 ; n19523
g19268 and n19173_not n19176_not ; n19524
g19269 and n19523_not n19524_not ; n19525
g19270 and n288 n19525_not ; n19526
g19271 and n19303_not n19526 ; n19527
g19272 and n19521_not n19527_not ; n19528
g19273 and b[27]_not n19528_not ; n19529
g19274 and n18834_not quotient[12]_not ; n19530
g19275 and n18844_not n19171 ; n19531
g19276 and n19167_not n19531 ; n19532
g19277 and n19168_not n19171_not ; n19533
g19278 and n19532_not n19533_not ; n19534
g19279 and n288 n19534_not ; n19535
g19280 and n19303_not n19535 ; n19536
g19281 and n19530_not n19536_not ; n19537
g19282 and b[26]_not n19537_not ; n19538
g19283 and n18843_not quotient[12]_not ; n19539
g19284 and n18853_not n19166 ; n19540
g19285 and n19162_not n19540 ; n19541
g19286 and n19163_not n19166_not ; n19542
g19287 and n19541_not n19542_not ; n19543
g19288 and n288 n19543_not ; n19544
g19289 and n19303_not n19544 ; n19545
g19290 and n19539_not n19545_not ; n19546
g19291 and b[25]_not n19546_not ; n19547
g19292 and n18852_not quotient[12]_not ; n19548
g19293 and n18862_not n19161 ; n19549
g19294 and n19157_not n19549 ; n19550
g19295 and n19158_not n19161_not ; n19551
g19296 and n19550_not n19551_not ; n19552
g19297 and n288 n19552_not ; n19553
g19298 and n19303_not n19553 ; n19554
g19299 and n19548_not n19554_not ; n19555
g19300 and b[24]_not n19555_not ; n19556
g19301 and n18861_not quotient[12]_not ; n19557
g19302 and n18871_not n19156 ; n19558
g19303 and n19152_not n19558 ; n19559
g19304 and n19153_not n19156_not ; n19560
g19305 and n19559_not n19560_not ; n19561
g19306 and n288 n19561_not ; n19562
g19307 and n19303_not n19562 ; n19563
g19308 and n19557_not n19563_not ; n19564
g19309 and b[23]_not n19564_not ; n19565
g19310 and n18870_not quotient[12]_not ; n19566
g19311 and n18880_not n19151 ; n19567
g19312 and n19147_not n19567 ; n19568
g19313 and n19148_not n19151_not ; n19569
g19314 and n19568_not n19569_not ; n19570
g19315 and n288 n19570_not ; n19571
g19316 and n19303_not n19571 ; n19572
g19317 and n19566_not n19572_not ; n19573
g19318 and b[22]_not n19573_not ; n19574
g19319 and n18879_not quotient[12]_not ; n19575
g19320 and n18889_not n19146 ; n19576
g19321 and n19142_not n19576 ; n19577
g19322 and n19143_not n19146_not ; n19578
g19323 and n19577_not n19578_not ; n19579
g19324 and n288 n19579_not ; n19580
g19325 and n19303_not n19580 ; n19581
g19326 and n19575_not n19581_not ; n19582
g19327 and b[21]_not n19582_not ; n19583
g19328 and n18888_not quotient[12]_not ; n19584
g19329 and n18898_not n19141 ; n19585
g19330 and n19137_not n19585 ; n19586
g19331 and n19138_not n19141_not ; n19587
g19332 and n19586_not n19587_not ; n19588
g19333 and n288 n19588_not ; n19589
g19334 and n19303_not n19589 ; n19590
g19335 and n19584_not n19590_not ; n19591
g19336 and b[20]_not n19591_not ; n19592
g19337 and n18897_not quotient[12]_not ; n19593
g19338 and n18907_not n19136 ; n19594
g19339 and n19132_not n19594 ; n19595
g19340 and n19133_not n19136_not ; n19596
g19341 and n19595_not n19596_not ; n19597
g19342 and n288 n19597_not ; n19598
g19343 and n19303_not n19598 ; n19599
g19344 and n19593_not n19599_not ; n19600
g19345 and b[19]_not n19600_not ; n19601
g19346 and n18906_not quotient[12]_not ; n19602
g19347 and n18916_not n19131 ; n19603
g19348 and n19127_not n19603 ; n19604
g19349 and n19128_not n19131_not ; n19605
g19350 and n19604_not n19605_not ; n19606
g19351 and n288 n19606_not ; n19607
g19352 and n19303_not n19607 ; n19608
g19353 and n19602_not n19608_not ; n19609
g19354 and b[18]_not n19609_not ; n19610
g19355 and n18915_not quotient[12]_not ; n19611
g19356 and n18925_not n19126 ; n19612
g19357 and n19122_not n19612 ; n19613
g19358 and n19123_not n19126_not ; n19614
g19359 and n19613_not n19614_not ; n19615
g19360 and n288 n19615_not ; n19616
g19361 and n19303_not n19616 ; n19617
g19362 and n19611_not n19617_not ; n19618
g19363 and b[17]_not n19618_not ; n19619
g19364 and n18924_not quotient[12]_not ; n19620
g19365 and n18934_not n19121 ; n19621
g19366 and n19117_not n19621 ; n19622
g19367 and n19118_not n19121_not ; n19623
g19368 and n19622_not n19623_not ; n19624
g19369 and n288 n19624_not ; n19625
g19370 and n19303_not n19625 ; n19626
g19371 and n19620_not n19626_not ; n19627
g19372 and b[16]_not n19627_not ; n19628
g19373 and n18933_not quotient[12]_not ; n19629
g19374 and n18943_not n19116 ; n19630
g19375 and n19112_not n19630 ; n19631
g19376 and n19113_not n19116_not ; n19632
g19377 and n19631_not n19632_not ; n19633
g19378 and n288 n19633_not ; n19634
g19379 and n19303_not n19634 ; n19635
g19380 and n19629_not n19635_not ; n19636
g19381 and b[15]_not n19636_not ; n19637
g19382 and n18942_not quotient[12]_not ; n19638
g19383 and n18952_not n19111 ; n19639
g19384 and n19107_not n19639 ; n19640
g19385 and n19108_not n19111_not ; n19641
g19386 and n19640_not n19641_not ; n19642
g19387 and n288 n19642_not ; n19643
g19388 and n19303_not n19643 ; n19644
g19389 and n19638_not n19644_not ; n19645
g19390 and b[14]_not n19645_not ; n19646
g19391 and n18951_not quotient[12]_not ; n19647
g19392 and n18961_not n19106 ; n19648
g19393 and n19102_not n19648 ; n19649
g19394 and n19103_not n19106_not ; n19650
g19395 and n19649_not n19650_not ; n19651
g19396 and n288 n19651_not ; n19652
g19397 and n19303_not n19652 ; n19653
g19398 and n19647_not n19653_not ; n19654
g19399 and b[13]_not n19654_not ; n19655
g19400 and n18960_not quotient[12]_not ; n19656
g19401 and n18970_not n19101 ; n19657
g19402 and n19097_not n19657 ; n19658
g19403 and n19098_not n19101_not ; n19659
g19404 and n19658_not n19659_not ; n19660
g19405 and n288 n19660_not ; n19661
g19406 and n19303_not n19661 ; n19662
g19407 and n19656_not n19662_not ; n19663
g19408 and b[12]_not n19663_not ; n19664
g19409 and n18969_not quotient[12]_not ; n19665
g19410 and n18979_not n19096 ; n19666
g19411 and n19092_not n19666 ; n19667
g19412 and n19093_not n19096_not ; n19668
g19413 and n19667_not n19668_not ; n19669
g19414 and n288 n19669_not ; n19670
g19415 and n19303_not n19670 ; n19671
g19416 and n19665_not n19671_not ; n19672
g19417 and b[11]_not n19672_not ; n19673
g19418 and n18978_not quotient[12]_not ; n19674
g19419 and n18988_not n19091 ; n19675
g19420 and n19087_not n19675 ; n19676
g19421 and n19088_not n19091_not ; n19677
g19422 and n19676_not n19677_not ; n19678
g19423 and n288 n19678_not ; n19679
g19424 and n19303_not n19679 ; n19680
g19425 and n19674_not n19680_not ; n19681
g19426 and b[10]_not n19681_not ; n19682
g19427 and n18987_not quotient[12]_not ; n19683
g19428 and n18997_not n19086 ; n19684
g19429 and n19082_not n19684 ; n19685
g19430 and n19083_not n19086_not ; n19686
g19431 and n19685_not n19686_not ; n19687
g19432 and n288 n19687_not ; n19688
g19433 and n19303_not n19688 ; n19689
g19434 and n19683_not n19689_not ; n19690
g19435 and b[9]_not n19690_not ; n19691
g19436 and n18996_not quotient[12]_not ; n19692
g19437 and n19006_not n19081 ; n19693
g19438 and n19077_not n19693 ; n19694
g19439 and n19078_not n19081_not ; n19695
g19440 and n19694_not n19695_not ; n19696
g19441 and n288 n19696_not ; n19697
g19442 and n19303_not n19697 ; n19698
g19443 and n19692_not n19698_not ; n19699
g19444 and b[8]_not n19699_not ; n19700
g19445 and n19005_not quotient[12]_not ; n19701
g19446 and n19015_not n19076 ; n19702
g19447 and n19072_not n19702 ; n19703
g19448 and n19073_not n19076_not ; n19704
g19449 and n19703_not n19704_not ; n19705
g19450 and n288 n19705_not ; n19706
g19451 and n19303_not n19706 ; n19707
g19452 and n19701_not n19707_not ; n19708
g19453 and b[7]_not n19708_not ; n19709
g19454 and n19014_not quotient[12]_not ; n19710
g19455 and n19024_not n19071 ; n19711
g19456 and n19067_not n19711 ; n19712
g19457 and n19068_not n19071_not ; n19713
g19458 and n19712_not n19713_not ; n19714
g19459 and n288 n19714_not ; n19715
g19460 and n19303_not n19715 ; n19716
g19461 and n19710_not n19716_not ; n19717
g19462 and b[6]_not n19717_not ; n19718
g19463 and n19023_not quotient[12]_not ; n19719
g19464 and n19033_not n19066 ; n19720
g19465 and n19062_not n19720 ; n19721
g19466 and n19063_not n19066_not ; n19722
g19467 and n19721_not n19722_not ; n19723
g19468 and n288 n19723_not ; n19724
g19469 and n19303_not n19724 ; n19725
g19470 and n19719_not n19725_not ; n19726
g19471 and b[5]_not n19726_not ; n19727
g19472 and n19032_not quotient[12]_not ; n19728
g19473 and n19041_not n19061 ; n19729
g19474 and n19057_not n19729 ; n19730
g19475 and n19058_not n19061_not ; n19731
g19476 and n19730_not n19731_not ; n19732
g19477 and n288 n19732_not ; n19733
g19478 and n19303_not n19733 ; n19734
g19479 and n19728_not n19734_not ; n19735
g19480 and b[4]_not n19735_not ; n19736
g19481 and n19040_not quotient[12]_not ; n19737
g19482 and n19052_not n19056 ; n19738
g19483 and n19051_not n19738 ; n19739
g19484 and n19053_not n19056_not ; n19740
g19485 and n19739_not n19740_not ; n19741
g19486 and n288 n19741_not ; n19742
g19487 and n19303_not n19742 ; n19743
g19488 and n19737_not n19743_not ; n19744
g19489 and b[3]_not n19744_not ; n19745
g19490 and n19045_not quotient[12]_not ; n19746
g19491 and n19048_not n19050 ; n19747
g19492 and n19046_not n19747 ; n19748
g19493 and n288 n19748_not ; n19749
g19494 and n19051_not n19749 ; n19750
g19495 and n19303_not n19750 ; n19751
g19496 and n19746_not n19751_not ; n19752
g19497 and b[2]_not n19752_not ; n19753
g19498 and b[0] b[52]_not ; n19754
g19499 and n397 n19754 ; n19755
g19500 and n407 n19755 ; n19756
g19501 and n19303_not n19756 ; n19757
g19502 and a[12] n19757_not ; n19758
g19503 and n286 n19050 ; n19759
g19504 and n337 n19759 ; n19760
g19505 and n19303_not n19760 ; n19761
g19506 and n19758_not n19761_not ; n19762
g19507 and b[1] n19762_not ; n19763
g19508 and b[1]_not n19761_not ; n19764
g19509 and n19758_not n19764 ; n19765
g19510 and n19763_not n19765_not ; n19766
g19511 and a[11]_not b[0] ; n19767
g19512 and n19766_not n19767_not ; n19768
g19513 and b[1]_not n19762_not ; n19769
g19514 and n19768_not n19769_not ; n19770
g19515 and b[2] n19751_not ; n19771
g19516 and n19746_not n19771 ; n19772
g19517 and n19753_not n19772_not ; n19773
g19518 and n19770_not n19773 ; n19774
g19519 and n19753_not n19774_not ; n19775
g19520 and b[3] n19743_not ; n19776
g19521 and n19737_not n19776 ; n19777
g19522 and n19745_not n19777_not ; n19778
g19523 and n19775_not n19778 ; n19779
g19524 and n19745_not n19779_not ; n19780
g19525 and b[4] n19734_not ; n19781
g19526 and n19728_not n19781 ; n19782
g19527 and n19736_not n19782_not ; n19783
g19528 and n19780_not n19783 ; n19784
g19529 and n19736_not n19784_not ; n19785
g19530 and b[5] n19725_not ; n19786
g19531 and n19719_not n19786 ; n19787
g19532 and n19727_not n19787_not ; n19788
g19533 and n19785_not n19788 ; n19789
g19534 and n19727_not n19789_not ; n19790
g19535 and b[6] n19716_not ; n19791
g19536 and n19710_not n19791 ; n19792
g19537 and n19718_not n19792_not ; n19793
g19538 and n19790_not n19793 ; n19794
g19539 and n19718_not n19794_not ; n19795
g19540 and b[7] n19707_not ; n19796
g19541 and n19701_not n19796 ; n19797
g19542 and n19709_not n19797_not ; n19798
g19543 and n19795_not n19798 ; n19799
g19544 and n19709_not n19799_not ; n19800
g19545 and b[8] n19698_not ; n19801
g19546 and n19692_not n19801 ; n19802
g19547 and n19700_not n19802_not ; n19803
g19548 and n19800_not n19803 ; n19804
g19549 and n19700_not n19804_not ; n19805
g19550 and b[9] n19689_not ; n19806
g19551 and n19683_not n19806 ; n19807
g19552 and n19691_not n19807_not ; n19808
g19553 and n19805_not n19808 ; n19809
g19554 and n19691_not n19809_not ; n19810
g19555 and b[10] n19680_not ; n19811
g19556 and n19674_not n19811 ; n19812
g19557 and n19682_not n19812_not ; n19813
g19558 and n19810_not n19813 ; n19814
g19559 and n19682_not n19814_not ; n19815
g19560 and b[11] n19671_not ; n19816
g19561 and n19665_not n19816 ; n19817
g19562 and n19673_not n19817_not ; n19818
g19563 and n19815_not n19818 ; n19819
g19564 and n19673_not n19819_not ; n19820
g19565 and b[12] n19662_not ; n19821
g19566 and n19656_not n19821 ; n19822
g19567 and n19664_not n19822_not ; n19823
g19568 and n19820_not n19823 ; n19824
g19569 and n19664_not n19824_not ; n19825
g19570 and b[13] n19653_not ; n19826
g19571 and n19647_not n19826 ; n19827
g19572 and n19655_not n19827_not ; n19828
g19573 and n19825_not n19828 ; n19829
g19574 and n19655_not n19829_not ; n19830
g19575 and b[14] n19644_not ; n19831
g19576 and n19638_not n19831 ; n19832
g19577 and n19646_not n19832_not ; n19833
g19578 and n19830_not n19833 ; n19834
g19579 and n19646_not n19834_not ; n19835
g19580 and b[15] n19635_not ; n19836
g19581 and n19629_not n19836 ; n19837
g19582 and n19637_not n19837_not ; n19838
g19583 and n19835_not n19838 ; n19839
g19584 and n19637_not n19839_not ; n19840
g19585 and b[16] n19626_not ; n19841
g19586 and n19620_not n19841 ; n19842
g19587 and n19628_not n19842_not ; n19843
g19588 and n19840_not n19843 ; n19844
g19589 and n19628_not n19844_not ; n19845
g19590 and b[17] n19617_not ; n19846
g19591 and n19611_not n19846 ; n19847
g19592 and n19619_not n19847_not ; n19848
g19593 and n19845_not n19848 ; n19849
g19594 and n19619_not n19849_not ; n19850
g19595 and b[18] n19608_not ; n19851
g19596 and n19602_not n19851 ; n19852
g19597 and n19610_not n19852_not ; n19853
g19598 and n19850_not n19853 ; n19854
g19599 and n19610_not n19854_not ; n19855
g19600 and b[19] n19599_not ; n19856
g19601 and n19593_not n19856 ; n19857
g19602 and n19601_not n19857_not ; n19858
g19603 and n19855_not n19858 ; n19859
g19604 and n19601_not n19859_not ; n19860
g19605 and b[20] n19590_not ; n19861
g19606 and n19584_not n19861 ; n19862
g19607 and n19592_not n19862_not ; n19863
g19608 and n19860_not n19863 ; n19864
g19609 and n19592_not n19864_not ; n19865
g19610 and b[21] n19581_not ; n19866
g19611 and n19575_not n19866 ; n19867
g19612 and n19583_not n19867_not ; n19868
g19613 and n19865_not n19868 ; n19869
g19614 and n19583_not n19869_not ; n19870
g19615 and b[22] n19572_not ; n19871
g19616 and n19566_not n19871 ; n19872
g19617 and n19574_not n19872_not ; n19873
g19618 and n19870_not n19873 ; n19874
g19619 and n19574_not n19874_not ; n19875
g19620 and b[23] n19563_not ; n19876
g19621 and n19557_not n19876 ; n19877
g19622 and n19565_not n19877_not ; n19878
g19623 and n19875_not n19878 ; n19879
g19624 and n19565_not n19879_not ; n19880
g19625 and b[24] n19554_not ; n19881
g19626 and n19548_not n19881 ; n19882
g19627 and n19556_not n19882_not ; n19883
g19628 and n19880_not n19883 ; n19884
g19629 and n19556_not n19884_not ; n19885
g19630 and b[25] n19545_not ; n19886
g19631 and n19539_not n19886 ; n19887
g19632 and n19547_not n19887_not ; n19888
g19633 and n19885_not n19888 ; n19889
g19634 and n19547_not n19889_not ; n19890
g19635 and b[26] n19536_not ; n19891
g19636 and n19530_not n19891 ; n19892
g19637 and n19538_not n19892_not ; n19893
g19638 and n19890_not n19893 ; n19894
g19639 and n19538_not n19894_not ; n19895
g19640 and b[27] n19527_not ; n19896
g19641 and n19521_not n19896 ; n19897
g19642 and n19529_not n19897_not ; n19898
g19643 and n19895_not n19898 ; n19899
g19644 and n19529_not n19899_not ; n19900
g19645 and b[28] n19518_not ; n19901
g19646 and n19512_not n19901 ; n19902
g19647 and n19520_not n19902_not ; n19903
g19648 and n19900_not n19903 ; n19904
g19649 and n19520_not n19904_not ; n19905
g19650 and b[29] n19509_not ; n19906
g19651 and n19503_not n19906 ; n19907
g19652 and n19511_not n19907_not ; n19908
g19653 and n19905_not n19908 ; n19909
g19654 and n19511_not n19909_not ; n19910
g19655 and b[30] n19500_not ; n19911
g19656 and n19494_not n19911 ; n19912
g19657 and n19502_not n19912_not ; n19913
g19658 and n19910_not n19913 ; n19914
g19659 and n19502_not n19914_not ; n19915
g19660 and b[31] n19491_not ; n19916
g19661 and n19485_not n19916 ; n19917
g19662 and n19493_not n19917_not ; n19918
g19663 and n19915_not n19918 ; n19919
g19664 and n19493_not n19919_not ; n19920
g19665 and b[32] n19482_not ; n19921
g19666 and n19476_not n19921 ; n19922
g19667 and n19484_not n19922_not ; n19923
g19668 and n19920_not n19923 ; n19924
g19669 and n19484_not n19924_not ; n19925
g19670 and b[33] n19473_not ; n19926
g19671 and n19467_not n19926 ; n19927
g19672 and n19475_not n19927_not ; n19928
g19673 and n19925_not n19928 ; n19929
g19674 and n19475_not n19929_not ; n19930
g19675 and b[34] n19464_not ; n19931
g19676 and n19458_not n19931 ; n19932
g19677 and n19466_not n19932_not ; n19933
g19678 and n19930_not n19933 ; n19934
g19679 and n19466_not n19934_not ; n19935
g19680 and b[35] n19455_not ; n19936
g19681 and n19449_not n19936 ; n19937
g19682 and n19457_not n19937_not ; n19938
g19683 and n19935_not n19938 ; n19939
g19684 and n19457_not n19939_not ; n19940
g19685 and b[36] n19446_not ; n19941
g19686 and n19440_not n19941 ; n19942
g19687 and n19448_not n19942_not ; n19943
g19688 and n19940_not n19943 ; n19944
g19689 and n19448_not n19944_not ; n19945
g19690 and b[37] n19437_not ; n19946
g19691 and n19431_not n19946 ; n19947
g19692 and n19439_not n19947_not ; n19948
g19693 and n19945_not n19948 ; n19949
g19694 and n19439_not n19949_not ; n19950
g19695 and b[38] n19428_not ; n19951
g19696 and n19422_not n19951 ; n19952
g19697 and n19430_not n19952_not ; n19953
g19698 and n19950_not n19953 ; n19954
g19699 and n19430_not n19954_not ; n19955
g19700 and b[39] n19419_not ; n19956
g19701 and n19413_not n19956 ; n19957
g19702 and n19421_not n19957_not ; n19958
g19703 and n19955_not n19958 ; n19959
g19704 and n19421_not n19959_not ; n19960
g19705 and b[40] n19410_not ; n19961
g19706 and n19404_not n19961 ; n19962
g19707 and n19412_not n19962_not ; n19963
g19708 and n19960_not n19963 ; n19964
g19709 and n19412_not n19964_not ; n19965
g19710 and b[41] n19401_not ; n19966
g19711 and n19395_not n19966 ; n19967
g19712 and n19403_not n19967_not ; n19968
g19713 and n19965_not n19968 ; n19969
g19714 and n19403_not n19969_not ; n19970
g19715 and b[42] n19392_not ; n19971
g19716 and n19386_not n19971 ; n19972
g19717 and n19394_not n19972_not ; n19973
g19718 and n19970_not n19973 ; n19974
g19719 and n19394_not n19974_not ; n19975
g19720 and b[43] n19383_not ; n19976
g19721 and n19377_not n19976 ; n19977
g19722 and n19385_not n19977_not ; n19978
g19723 and n19975_not n19978 ; n19979
g19724 and n19385_not n19979_not ; n19980
g19725 and b[44] n19374_not ; n19981
g19726 and n19368_not n19981 ; n19982
g19727 and n19376_not n19982_not ; n19983
g19728 and n19980_not n19983 ; n19984
g19729 and n19376_not n19984_not ; n19985
g19730 and b[45] n19365_not ; n19986
g19731 and n19359_not n19986 ; n19987
g19732 and n19367_not n19987_not ; n19988
g19733 and n19985_not n19988 ; n19989
g19734 and n19367_not n19989_not ; n19990
g19735 and b[46] n19356_not ; n19991
g19736 and n19350_not n19991 ; n19992
g19737 and n19358_not n19992_not ; n19993
g19738 and n19990_not n19993 ; n19994
g19739 and n19358_not n19994_not ; n19995
g19740 and b[47] n19347_not ; n19996
g19741 and n19341_not n19996 ; n19997
g19742 and n19349_not n19997_not ; n19998
g19743 and n19995_not n19998 ; n19999
g19744 and n19349_not n19999_not ; n20000
g19745 and b[48] n19338_not ; n20001
g19746 and n19332_not n20001 ; n20002
g19747 and n19340_not n20002_not ; n20003
g19748 and n20000_not n20003 ; n20004
g19749 and n19340_not n20004_not ; n20005
g19750 and b[49] n19329_not ; n20006
g19751 and n19323_not n20006 ; n20007
g19752 and n19331_not n20007_not ; n20008
g19753 and n20005_not n20008 ; n20009
g19754 and n19331_not n20009_not ; n20010
g19755 and b[50] n19320_not ; n20011
g19756 and n19314_not n20011 ; n20012
g19757 and n19322_not n20012_not ; n20013
g19758 and n20010_not n20013 ; n20014
g19759 and n19322_not n20014_not ; n20015
g19760 and b[51] n19311_not ; n20016
g19761 and n19305_not n20016 ; n20017
g19762 and n19313_not n20017_not ; n20018
g19763 and n20015_not n20018 ; n20019
g19764 and n19313_not n20019_not ; n20020
g19765 and n18608_not quotient[12]_not ; n20021
g19766 and n18610_not n19301 ; n20022
g19767 and n19297_not n20022 ; n20023
g19768 and n19298_not n19301_not ; n20024
g19769 and n20023_not n20024_not ; n20025
g19770 and quotient[12] n20025_not ; n20026
g19771 and n20021_not n20026_not ; n20027
g19772 and b[52]_not n20027_not ; n20028
g19773 and b[52] n20021_not ; n20029
g19774 and n20026_not n20029 ; n20030
g19775 and n595 n20030_not ; n20031
g19776 and n20028_not n20031 ; n20032
g19777 and n20020_not n20032 ; n20033
g19778 and n288 n20027_not ; n20034
g19779 and n20033_not n20034_not ; quotient[11]
g19780 and n19322_not n20018 ; n20036
g19781 and n20014_not n20036 ; n20037
g19782 and n20015_not n20018_not ; n20038
g19783 and n20037_not n20038_not ; n20039
g19784 and quotient[11] n20039_not ; n20040
g19785 and n19312_not n20034_not ; n20041
g19786 and n20033_not n20041 ; n20042
g19787 and n20040_not n20042_not ; n20043
g19788 and b[52]_not n20043_not ; n20044
g19789 and n19331_not n20013 ; n20045
g19790 and n20009_not n20045 ; n20046
g19791 and n20010_not n20013_not ; n20047
g19792 and n20046_not n20047_not ; n20048
g19793 and quotient[11] n20048_not ; n20049
g19794 and n19321_not n20034_not ; n20050
g19795 and n20033_not n20050 ; n20051
g19796 and n20049_not n20051_not ; n20052
g19797 and b[51]_not n20052_not ; n20053
g19798 and n19340_not n20008 ; n20054
g19799 and n20004_not n20054 ; n20055
g19800 and n20005_not n20008_not ; n20056
g19801 and n20055_not n20056_not ; n20057
g19802 and quotient[11] n20057_not ; n20058
g19803 and n19330_not n20034_not ; n20059
g19804 and n20033_not n20059 ; n20060
g19805 and n20058_not n20060_not ; n20061
g19806 and b[50]_not n20061_not ; n20062
g19807 and n19349_not n20003 ; n20063
g19808 and n19999_not n20063 ; n20064
g19809 and n20000_not n20003_not ; n20065
g19810 and n20064_not n20065_not ; n20066
g19811 and quotient[11] n20066_not ; n20067
g19812 and n19339_not n20034_not ; n20068
g19813 and n20033_not n20068 ; n20069
g19814 and n20067_not n20069_not ; n20070
g19815 and b[49]_not n20070_not ; n20071
g19816 and n19358_not n19998 ; n20072
g19817 and n19994_not n20072 ; n20073
g19818 and n19995_not n19998_not ; n20074
g19819 and n20073_not n20074_not ; n20075
g19820 and quotient[11] n20075_not ; n20076
g19821 and n19348_not n20034_not ; n20077
g19822 and n20033_not n20077 ; n20078
g19823 and n20076_not n20078_not ; n20079
g19824 and b[48]_not n20079_not ; n20080
g19825 and n19367_not n19993 ; n20081
g19826 and n19989_not n20081 ; n20082
g19827 and n19990_not n19993_not ; n20083
g19828 and n20082_not n20083_not ; n20084
g19829 and quotient[11] n20084_not ; n20085
g19830 and n19357_not n20034_not ; n20086
g19831 and n20033_not n20086 ; n20087
g19832 and n20085_not n20087_not ; n20088
g19833 and b[47]_not n20088_not ; n20089
g19834 and n19376_not n19988 ; n20090
g19835 and n19984_not n20090 ; n20091
g19836 and n19985_not n19988_not ; n20092
g19837 and n20091_not n20092_not ; n20093
g19838 and quotient[11] n20093_not ; n20094
g19839 and n19366_not n20034_not ; n20095
g19840 and n20033_not n20095 ; n20096
g19841 and n20094_not n20096_not ; n20097
g19842 and b[46]_not n20097_not ; n20098
g19843 and n19385_not n19983 ; n20099
g19844 and n19979_not n20099 ; n20100
g19845 and n19980_not n19983_not ; n20101
g19846 and n20100_not n20101_not ; n20102
g19847 and quotient[11] n20102_not ; n20103
g19848 and n19375_not n20034_not ; n20104
g19849 and n20033_not n20104 ; n20105
g19850 and n20103_not n20105_not ; n20106
g19851 and b[45]_not n20106_not ; n20107
g19852 and n19394_not n19978 ; n20108
g19853 and n19974_not n20108 ; n20109
g19854 and n19975_not n19978_not ; n20110
g19855 and n20109_not n20110_not ; n20111
g19856 and quotient[11] n20111_not ; n20112
g19857 and n19384_not n20034_not ; n20113
g19858 and n20033_not n20113 ; n20114
g19859 and n20112_not n20114_not ; n20115
g19860 and b[44]_not n20115_not ; n20116
g19861 and n19403_not n19973 ; n20117
g19862 and n19969_not n20117 ; n20118
g19863 and n19970_not n19973_not ; n20119
g19864 and n20118_not n20119_not ; n20120
g19865 and quotient[11] n20120_not ; n20121
g19866 and n19393_not n20034_not ; n20122
g19867 and n20033_not n20122 ; n20123
g19868 and n20121_not n20123_not ; n20124
g19869 and b[43]_not n20124_not ; n20125
g19870 and n19412_not n19968 ; n20126
g19871 and n19964_not n20126 ; n20127
g19872 and n19965_not n19968_not ; n20128
g19873 and n20127_not n20128_not ; n20129
g19874 and quotient[11] n20129_not ; n20130
g19875 and n19402_not n20034_not ; n20131
g19876 and n20033_not n20131 ; n20132
g19877 and n20130_not n20132_not ; n20133
g19878 and b[42]_not n20133_not ; n20134
g19879 and n19421_not n19963 ; n20135
g19880 and n19959_not n20135 ; n20136
g19881 and n19960_not n19963_not ; n20137
g19882 and n20136_not n20137_not ; n20138
g19883 and quotient[11] n20138_not ; n20139
g19884 and n19411_not n20034_not ; n20140
g19885 and n20033_not n20140 ; n20141
g19886 and n20139_not n20141_not ; n20142
g19887 and b[41]_not n20142_not ; n20143
g19888 and n19430_not n19958 ; n20144
g19889 and n19954_not n20144 ; n20145
g19890 and n19955_not n19958_not ; n20146
g19891 and n20145_not n20146_not ; n20147
g19892 and quotient[11] n20147_not ; n20148
g19893 and n19420_not n20034_not ; n20149
g19894 and n20033_not n20149 ; n20150
g19895 and n20148_not n20150_not ; n20151
g19896 and b[40]_not n20151_not ; n20152
g19897 and n19439_not n19953 ; n20153
g19898 and n19949_not n20153 ; n20154
g19899 and n19950_not n19953_not ; n20155
g19900 and n20154_not n20155_not ; n20156
g19901 and quotient[11] n20156_not ; n20157
g19902 and n19429_not n20034_not ; n20158
g19903 and n20033_not n20158 ; n20159
g19904 and n20157_not n20159_not ; n20160
g19905 and b[39]_not n20160_not ; n20161
g19906 and n19448_not n19948 ; n20162
g19907 and n19944_not n20162 ; n20163
g19908 and n19945_not n19948_not ; n20164
g19909 and n20163_not n20164_not ; n20165
g19910 and quotient[11] n20165_not ; n20166
g19911 and n19438_not n20034_not ; n20167
g19912 and n20033_not n20167 ; n20168
g19913 and n20166_not n20168_not ; n20169
g19914 and b[38]_not n20169_not ; n20170
g19915 and n19457_not n19943 ; n20171
g19916 and n19939_not n20171 ; n20172
g19917 and n19940_not n19943_not ; n20173
g19918 and n20172_not n20173_not ; n20174
g19919 and quotient[11] n20174_not ; n20175
g19920 and n19447_not n20034_not ; n20176
g19921 and n20033_not n20176 ; n20177
g19922 and n20175_not n20177_not ; n20178
g19923 and b[37]_not n20178_not ; n20179
g19924 and n19466_not n19938 ; n20180
g19925 and n19934_not n20180 ; n20181
g19926 and n19935_not n19938_not ; n20182
g19927 and n20181_not n20182_not ; n20183
g19928 and quotient[11] n20183_not ; n20184
g19929 and n19456_not n20034_not ; n20185
g19930 and n20033_not n20185 ; n20186
g19931 and n20184_not n20186_not ; n20187
g19932 and b[36]_not n20187_not ; n20188
g19933 and n19475_not n19933 ; n20189
g19934 and n19929_not n20189 ; n20190
g19935 and n19930_not n19933_not ; n20191
g19936 and n20190_not n20191_not ; n20192
g19937 and quotient[11] n20192_not ; n20193
g19938 and n19465_not n20034_not ; n20194
g19939 and n20033_not n20194 ; n20195
g19940 and n20193_not n20195_not ; n20196
g19941 and b[35]_not n20196_not ; n20197
g19942 and n19484_not n19928 ; n20198
g19943 and n19924_not n20198 ; n20199
g19944 and n19925_not n19928_not ; n20200
g19945 and n20199_not n20200_not ; n20201
g19946 and quotient[11] n20201_not ; n20202
g19947 and n19474_not n20034_not ; n20203
g19948 and n20033_not n20203 ; n20204
g19949 and n20202_not n20204_not ; n20205
g19950 and b[34]_not n20205_not ; n20206
g19951 and n19493_not n19923 ; n20207
g19952 and n19919_not n20207 ; n20208
g19953 and n19920_not n19923_not ; n20209
g19954 and n20208_not n20209_not ; n20210
g19955 and quotient[11] n20210_not ; n20211
g19956 and n19483_not n20034_not ; n20212
g19957 and n20033_not n20212 ; n20213
g19958 and n20211_not n20213_not ; n20214
g19959 and b[33]_not n20214_not ; n20215
g19960 and n19502_not n19918 ; n20216
g19961 and n19914_not n20216 ; n20217
g19962 and n19915_not n19918_not ; n20218
g19963 and n20217_not n20218_not ; n20219
g19964 and quotient[11] n20219_not ; n20220
g19965 and n19492_not n20034_not ; n20221
g19966 and n20033_not n20221 ; n20222
g19967 and n20220_not n20222_not ; n20223
g19968 and b[32]_not n20223_not ; n20224
g19969 and n19511_not n19913 ; n20225
g19970 and n19909_not n20225 ; n20226
g19971 and n19910_not n19913_not ; n20227
g19972 and n20226_not n20227_not ; n20228
g19973 and quotient[11] n20228_not ; n20229
g19974 and n19501_not n20034_not ; n20230
g19975 and n20033_not n20230 ; n20231
g19976 and n20229_not n20231_not ; n20232
g19977 and b[31]_not n20232_not ; n20233
g19978 and n19520_not n19908 ; n20234
g19979 and n19904_not n20234 ; n20235
g19980 and n19905_not n19908_not ; n20236
g19981 and n20235_not n20236_not ; n20237
g19982 and quotient[11] n20237_not ; n20238
g19983 and n19510_not n20034_not ; n20239
g19984 and n20033_not n20239 ; n20240
g19985 and n20238_not n20240_not ; n20241
g19986 and b[30]_not n20241_not ; n20242
g19987 and n19529_not n19903 ; n20243
g19988 and n19899_not n20243 ; n20244
g19989 and n19900_not n19903_not ; n20245
g19990 and n20244_not n20245_not ; n20246
g19991 and quotient[11] n20246_not ; n20247
g19992 and n19519_not n20034_not ; n20248
g19993 and n20033_not n20248 ; n20249
g19994 and n20247_not n20249_not ; n20250
g19995 and b[29]_not n20250_not ; n20251
g19996 and n19538_not n19898 ; n20252
g19997 and n19894_not n20252 ; n20253
g19998 and n19895_not n19898_not ; n20254
g19999 and n20253_not n20254_not ; n20255
g20000 and quotient[11] n20255_not ; n20256
g20001 and n19528_not n20034_not ; n20257
g20002 and n20033_not n20257 ; n20258
g20003 and n20256_not n20258_not ; n20259
g20004 and b[28]_not n20259_not ; n20260
g20005 and n19547_not n19893 ; n20261
g20006 and n19889_not n20261 ; n20262
g20007 and n19890_not n19893_not ; n20263
g20008 and n20262_not n20263_not ; n20264
g20009 and quotient[11] n20264_not ; n20265
g20010 and n19537_not n20034_not ; n20266
g20011 and n20033_not n20266 ; n20267
g20012 and n20265_not n20267_not ; n20268
g20013 and b[27]_not n20268_not ; n20269
g20014 and n19556_not n19888 ; n20270
g20015 and n19884_not n20270 ; n20271
g20016 and n19885_not n19888_not ; n20272
g20017 and n20271_not n20272_not ; n20273
g20018 and quotient[11] n20273_not ; n20274
g20019 and n19546_not n20034_not ; n20275
g20020 and n20033_not n20275 ; n20276
g20021 and n20274_not n20276_not ; n20277
g20022 and b[26]_not n20277_not ; n20278
g20023 and n19565_not n19883 ; n20279
g20024 and n19879_not n20279 ; n20280
g20025 and n19880_not n19883_not ; n20281
g20026 and n20280_not n20281_not ; n20282
g20027 and quotient[11] n20282_not ; n20283
g20028 and n19555_not n20034_not ; n20284
g20029 and n20033_not n20284 ; n20285
g20030 and n20283_not n20285_not ; n20286
g20031 and b[25]_not n20286_not ; n20287
g20032 and n19574_not n19878 ; n20288
g20033 and n19874_not n20288 ; n20289
g20034 and n19875_not n19878_not ; n20290
g20035 and n20289_not n20290_not ; n20291
g20036 and quotient[11] n20291_not ; n20292
g20037 and n19564_not n20034_not ; n20293
g20038 and n20033_not n20293 ; n20294
g20039 and n20292_not n20294_not ; n20295
g20040 and b[24]_not n20295_not ; n20296
g20041 and n19583_not n19873 ; n20297
g20042 and n19869_not n20297 ; n20298
g20043 and n19870_not n19873_not ; n20299
g20044 and n20298_not n20299_not ; n20300
g20045 and quotient[11] n20300_not ; n20301
g20046 and n19573_not n20034_not ; n20302
g20047 and n20033_not n20302 ; n20303
g20048 and n20301_not n20303_not ; n20304
g20049 and b[23]_not n20304_not ; n20305
g20050 and n19592_not n19868 ; n20306
g20051 and n19864_not n20306 ; n20307
g20052 and n19865_not n19868_not ; n20308
g20053 and n20307_not n20308_not ; n20309
g20054 and quotient[11] n20309_not ; n20310
g20055 and n19582_not n20034_not ; n20311
g20056 and n20033_not n20311 ; n20312
g20057 and n20310_not n20312_not ; n20313
g20058 and b[22]_not n20313_not ; n20314
g20059 and n19601_not n19863 ; n20315
g20060 and n19859_not n20315 ; n20316
g20061 and n19860_not n19863_not ; n20317
g20062 and n20316_not n20317_not ; n20318
g20063 and quotient[11] n20318_not ; n20319
g20064 and n19591_not n20034_not ; n20320
g20065 and n20033_not n20320 ; n20321
g20066 and n20319_not n20321_not ; n20322
g20067 and b[21]_not n20322_not ; n20323
g20068 and n19610_not n19858 ; n20324
g20069 and n19854_not n20324 ; n20325
g20070 and n19855_not n19858_not ; n20326
g20071 and n20325_not n20326_not ; n20327
g20072 and quotient[11] n20327_not ; n20328
g20073 and n19600_not n20034_not ; n20329
g20074 and n20033_not n20329 ; n20330
g20075 and n20328_not n20330_not ; n20331
g20076 and b[20]_not n20331_not ; n20332
g20077 and n19619_not n19853 ; n20333
g20078 and n19849_not n20333 ; n20334
g20079 and n19850_not n19853_not ; n20335
g20080 and n20334_not n20335_not ; n20336
g20081 and quotient[11] n20336_not ; n20337
g20082 and n19609_not n20034_not ; n20338
g20083 and n20033_not n20338 ; n20339
g20084 and n20337_not n20339_not ; n20340
g20085 and b[19]_not n20340_not ; n20341
g20086 and n19628_not n19848 ; n20342
g20087 and n19844_not n20342 ; n20343
g20088 and n19845_not n19848_not ; n20344
g20089 and n20343_not n20344_not ; n20345
g20090 and quotient[11] n20345_not ; n20346
g20091 and n19618_not n20034_not ; n20347
g20092 and n20033_not n20347 ; n20348
g20093 and n20346_not n20348_not ; n20349
g20094 and b[18]_not n20349_not ; n20350
g20095 and n19637_not n19843 ; n20351
g20096 and n19839_not n20351 ; n20352
g20097 and n19840_not n19843_not ; n20353
g20098 and n20352_not n20353_not ; n20354
g20099 and quotient[11] n20354_not ; n20355
g20100 and n19627_not n20034_not ; n20356
g20101 and n20033_not n20356 ; n20357
g20102 and n20355_not n20357_not ; n20358
g20103 and b[17]_not n20358_not ; n20359
g20104 and n19646_not n19838 ; n20360
g20105 and n19834_not n20360 ; n20361
g20106 and n19835_not n19838_not ; n20362
g20107 and n20361_not n20362_not ; n20363
g20108 and quotient[11] n20363_not ; n20364
g20109 and n19636_not n20034_not ; n20365
g20110 and n20033_not n20365 ; n20366
g20111 and n20364_not n20366_not ; n20367
g20112 and b[16]_not n20367_not ; n20368
g20113 and n19655_not n19833 ; n20369
g20114 and n19829_not n20369 ; n20370
g20115 and n19830_not n19833_not ; n20371
g20116 and n20370_not n20371_not ; n20372
g20117 and quotient[11] n20372_not ; n20373
g20118 and n19645_not n20034_not ; n20374
g20119 and n20033_not n20374 ; n20375
g20120 and n20373_not n20375_not ; n20376
g20121 and b[15]_not n20376_not ; n20377
g20122 and n19664_not n19828 ; n20378
g20123 and n19824_not n20378 ; n20379
g20124 and n19825_not n19828_not ; n20380
g20125 and n20379_not n20380_not ; n20381
g20126 and quotient[11] n20381_not ; n20382
g20127 and n19654_not n20034_not ; n20383
g20128 and n20033_not n20383 ; n20384
g20129 and n20382_not n20384_not ; n20385
g20130 and b[14]_not n20385_not ; n20386
g20131 and n19673_not n19823 ; n20387
g20132 and n19819_not n20387 ; n20388
g20133 and n19820_not n19823_not ; n20389
g20134 and n20388_not n20389_not ; n20390
g20135 and quotient[11] n20390_not ; n20391
g20136 and n19663_not n20034_not ; n20392
g20137 and n20033_not n20392 ; n20393
g20138 and n20391_not n20393_not ; n20394
g20139 and b[13]_not n20394_not ; n20395
g20140 and n19682_not n19818 ; n20396
g20141 and n19814_not n20396 ; n20397
g20142 and n19815_not n19818_not ; n20398
g20143 and n20397_not n20398_not ; n20399
g20144 and quotient[11] n20399_not ; n20400
g20145 and n19672_not n20034_not ; n20401
g20146 and n20033_not n20401 ; n20402
g20147 and n20400_not n20402_not ; n20403
g20148 and b[12]_not n20403_not ; n20404
g20149 and n19691_not n19813 ; n20405
g20150 and n19809_not n20405 ; n20406
g20151 and n19810_not n19813_not ; n20407
g20152 and n20406_not n20407_not ; n20408
g20153 and quotient[11] n20408_not ; n20409
g20154 and n19681_not n20034_not ; n20410
g20155 and n20033_not n20410 ; n20411
g20156 and n20409_not n20411_not ; n20412
g20157 and b[11]_not n20412_not ; n20413
g20158 and n19700_not n19808 ; n20414
g20159 and n19804_not n20414 ; n20415
g20160 and n19805_not n19808_not ; n20416
g20161 and n20415_not n20416_not ; n20417
g20162 and quotient[11] n20417_not ; n20418
g20163 and n19690_not n20034_not ; n20419
g20164 and n20033_not n20419 ; n20420
g20165 and n20418_not n20420_not ; n20421
g20166 and b[10]_not n20421_not ; n20422
g20167 and n19709_not n19803 ; n20423
g20168 and n19799_not n20423 ; n20424
g20169 and n19800_not n19803_not ; n20425
g20170 and n20424_not n20425_not ; n20426
g20171 and quotient[11] n20426_not ; n20427
g20172 and n19699_not n20034_not ; n20428
g20173 and n20033_not n20428 ; n20429
g20174 and n20427_not n20429_not ; n20430
g20175 and b[9]_not n20430_not ; n20431
g20176 and n19718_not n19798 ; n20432
g20177 and n19794_not n20432 ; n20433
g20178 and n19795_not n19798_not ; n20434
g20179 and n20433_not n20434_not ; n20435
g20180 and quotient[11] n20435_not ; n20436
g20181 and n19708_not n20034_not ; n20437
g20182 and n20033_not n20437 ; n20438
g20183 and n20436_not n20438_not ; n20439
g20184 and b[8]_not n20439_not ; n20440
g20185 and n19727_not n19793 ; n20441
g20186 and n19789_not n20441 ; n20442
g20187 and n19790_not n19793_not ; n20443
g20188 and n20442_not n20443_not ; n20444
g20189 and quotient[11] n20444_not ; n20445
g20190 and n19717_not n20034_not ; n20446
g20191 and n20033_not n20446 ; n20447
g20192 and n20445_not n20447_not ; n20448
g20193 and b[7]_not n20448_not ; n20449
g20194 and n19736_not n19788 ; n20450
g20195 and n19784_not n20450 ; n20451
g20196 and n19785_not n19788_not ; n20452
g20197 and n20451_not n20452_not ; n20453
g20198 and quotient[11] n20453_not ; n20454
g20199 and n19726_not n20034_not ; n20455
g20200 and n20033_not n20455 ; n20456
g20201 and n20454_not n20456_not ; n20457
g20202 and b[6]_not n20457_not ; n20458
g20203 and n19745_not n19783 ; n20459
g20204 and n19779_not n20459 ; n20460
g20205 and n19780_not n19783_not ; n20461
g20206 and n20460_not n20461_not ; n20462
g20207 and quotient[11] n20462_not ; n20463
g20208 and n19735_not n20034_not ; n20464
g20209 and n20033_not n20464 ; n20465
g20210 and n20463_not n20465_not ; n20466
g20211 and b[5]_not n20466_not ; n20467
g20212 and n19753_not n19778 ; n20468
g20213 and n19774_not n20468 ; n20469
g20214 and n19775_not n19778_not ; n20470
g20215 and n20469_not n20470_not ; n20471
g20216 and quotient[11] n20471_not ; n20472
g20217 and n19744_not n20034_not ; n20473
g20218 and n20033_not n20473 ; n20474
g20219 and n20472_not n20474_not ; n20475
g20220 and b[4]_not n20475_not ; n20476
g20221 and n19769_not n19773 ; n20477
g20222 and n19768_not n20477 ; n20478
g20223 and n19770_not n19773_not ; n20479
g20224 and n20478_not n20479_not ; n20480
g20225 and quotient[11] n20480_not ; n20481
g20226 and n19752_not n20034_not ; n20482
g20227 and n20033_not n20482 ; n20483
g20228 and n20481_not n20483_not ; n20484
g20229 and b[3]_not n20484_not ; n20485
g20230 and n19765_not n19767 ; n20486
g20231 and n19763_not n20486 ; n20487
g20232 and n19768_not n20487_not ; n20488
g20233 and quotient[11] n20488 ; n20489
g20234 and n19762_not n20034_not ; n20490
g20235 and n20033_not n20490 ; n20491
g20236 and n20489_not n20491_not ; n20492
g20237 and b[2]_not n20492_not ; n20493
g20238 and b[0] quotient[11] ; n20494
g20239 and a[11] n20494_not ; n20495
g20240 and n19767 quotient[11] ; n20496
g20241 and n20495_not n20496_not ; n20497
g20242 and b[1] n20497_not ; n20498
g20243 and b[1]_not n20496_not ; n20499
g20244 and n20495_not n20499 ; n20500
g20245 and n20498_not n20500_not ; n20501
g20246 and a[10]_not b[0] ; n20502
g20247 and n20501_not n20502_not ; n20503
g20248 and b[1]_not n20497_not ; n20504
g20249 and n20503_not n20504_not ; n20505
g20250 and b[2] n20491_not ; n20506
g20251 and n20489_not n20506 ; n20507
g20252 and n20493_not n20507_not ; n20508
g20253 and n20505_not n20508 ; n20509
g20254 and n20493_not n20509_not ; n20510
g20255 and b[3] n20483_not ; n20511
g20256 and n20481_not n20511 ; n20512
g20257 and n20485_not n20512_not ; n20513
g20258 and n20510_not n20513 ; n20514
g20259 and n20485_not n20514_not ; n20515
g20260 and b[4] n20474_not ; n20516
g20261 and n20472_not n20516 ; n20517
g20262 and n20476_not n20517_not ; n20518
g20263 and n20515_not n20518 ; n20519
g20264 and n20476_not n20519_not ; n20520
g20265 and b[5] n20465_not ; n20521
g20266 and n20463_not n20521 ; n20522
g20267 and n20467_not n20522_not ; n20523
g20268 and n20520_not n20523 ; n20524
g20269 and n20467_not n20524_not ; n20525
g20270 and b[6] n20456_not ; n20526
g20271 and n20454_not n20526 ; n20527
g20272 and n20458_not n20527_not ; n20528
g20273 and n20525_not n20528 ; n20529
g20274 and n20458_not n20529_not ; n20530
g20275 and b[7] n20447_not ; n20531
g20276 and n20445_not n20531 ; n20532
g20277 and n20449_not n20532_not ; n20533
g20278 and n20530_not n20533 ; n20534
g20279 and n20449_not n20534_not ; n20535
g20280 and b[8] n20438_not ; n20536
g20281 and n20436_not n20536 ; n20537
g20282 and n20440_not n20537_not ; n20538
g20283 and n20535_not n20538 ; n20539
g20284 and n20440_not n20539_not ; n20540
g20285 and b[9] n20429_not ; n20541
g20286 and n20427_not n20541 ; n20542
g20287 and n20431_not n20542_not ; n20543
g20288 and n20540_not n20543 ; n20544
g20289 and n20431_not n20544_not ; n20545
g20290 and b[10] n20420_not ; n20546
g20291 and n20418_not n20546 ; n20547
g20292 and n20422_not n20547_not ; n20548
g20293 and n20545_not n20548 ; n20549
g20294 and n20422_not n20549_not ; n20550
g20295 and b[11] n20411_not ; n20551
g20296 and n20409_not n20551 ; n20552
g20297 and n20413_not n20552_not ; n20553
g20298 and n20550_not n20553 ; n20554
g20299 and n20413_not n20554_not ; n20555
g20300 and b[12] n20402_not ; n20556
g20301 and n20400_not n20556 ; n20557
g20302 and n20404_not n20557_not ; n20558
g20303 and n20555_not n20558 ; n20559
g20304 and n20404_not n20559_not ; n20560
g20305 and b[13] n20393_not ; n20561
g20306 and n20391_not n20561 ; n20562
g20307 and n20395_not n20562_not ; n20563
g20308 and n20560_not n20563 ; n20564
g20309 and n20395_not n20564_not ; n20565
g20310 and b[14] n20384_not ; n20566
g20311 and n20382_not n20566 ; n20567
g20312 and n20386_not n20567_not ; n20568
g20313 and n20565_not n20568 ; n20569
g20314 and n20386_not n20569_not ; n20570
g20315 and b[15] n20375_not ; n20571
g20316 and n20373_not n20571 ; n20572
g20317 and n20377_not n20572_not ; n20573
g20318 and n20570_not n20573 ; n20574
g20319 and n20377_not n20574_not ; n20575
g20320 and b[16] n20366_not ; n20576
g20321 and n20364_not n20576 ; n20577
g20322 and n20368_not n20577_not ; n20578
g20323 and n20575_not n20578 ; n20579
g20324 and n20368_not n20579_not ; n20580
g20325 and b[17] n20357_not ; n20581
g20326 and n20355_not n20581 ; n20582
g20327 and n20359_not n20582_not ; n20583
g20328 and n20580_not n20583 ; n20584
g20329 and n20359_not n20584_not ; n20585
g20330 and b[18] n20348_not ; n20586
g20331 and n20346_not n20586 ; n20587
g20332 and n20350_not n20587_not ; n20588
g20333 and n20585_not n20588 ; n20589
g20334 and n20350_not n20589_not ; n20590
g20335 and b[19] n20339_not ; n20591
g20336 and n20337_not n20591 ; n20592
g20337 and n20341_not n20592_not ; n20593
g20338 and n20590_not n20593 ; n20594
g20339 and n20341_not n20594_not ; n20595
g20340 and b[20] n20330_not ; n20596
g20341 and n20328_not n20596 ; n20597
g20342 and n20332_not n20597_not ; n20598
g20343 and n20595_not n20598 ; n20599
g20344 and n20332_not n20599_not ; n20600
g20345 and b[21] n20321_not ; n20601
g20346 and n20319_not n20601 ; n20602
g20347 and n20323_not n20602_not ; n20603
g20348 and n20600_not n20603 ; n20604
g20349 and n20323_not n20604_not ; n20605
g20350 and b[22] n20312_not ; n20606
g20351 and n20310_not n20606 ; n20607
g20352 and n20314_not n20607_not ; n20608
g20353 and n20605_not n20608 ; n20609
g20354 and n20314_not n20609_not ; n20610
g20355 and b[23] n20303_not ; n20611
g20356 and n20301_not n20611 ; n20612
g20357 and n20305_not n20612_not ; n20613
g20358 and n20610_not n20613 ; n20614
g20359 and n20305_not n20614_not ; n20615
g20360 and b[24] n20294_not ; n20616
g20361 and n20292_not n20616 ; n20617
g20362 and n20296_not n20617_not ; n20618
g20363 and n20615_not n20618 ; n20619
g20364 and n20296_not n20619_not ; n20620
g20365 and b[25] n20285_not ; n20621
g20366 and n20283_not n20621 ; n20622
g20367 and n20287_not n20622_not ; n20623
g20368 and n20620_not n20623 ; n20624
g20369 and n20287_not n20624_not ; n20625
g20370 and b[26] n20276_not ; n20626
g20371 and n20274_not n20626 ; n20627
g20372 and n20278_not n20627_not ; n20628
g20373 and n20625_not n20628 ; n20629
g20374 and n20278_not n20629_not ; n20630
g20375 and b[27] n20267_not ; n20631
g20376 and n20265_not n20631 ; n20632
g20377 and n20269_not n20632_not ; n20633
g20378 and n20630_not n20633 ; n20634
g20379 and n20269_not n20634_not ; n20635
g20380 and b[28] n20258_not ; n20636
g20381 and n20256_not n20636 ; n20637
g20382 and n20260_not n20637_not ; n20638
g20383 and n20635_not n20638 ; n20639
g20384 and n20260_not n20639_not ; n20640
g20385 and b[29] n20249_not ; n20641
g20386 and n20247_not n20641 ; n20642
g20387 and n20251_not n20642_not ; n20643
g20388 and n20640_not n20643 ; n20644
g20389 and n20251_not n20644_not ; n20645
g20390 and b[30] n20240_not ; n20646
g20391 and n20238_not n20646 ; n20647
g20392 and n20242_not n20647_not ; n20648
g20393 and n20645_not n20648 ; n20649
g20394 and n20242_not n20649_not ; n20650
g20395 and b[31] n20231_not ; n20651
g20396 and n20229_not n20651 ; n20652
g20397 and n20233_not n20652_not ; n20653
g20398 and n20650_not n20653 ; n20654
g20399 and n20233_not n20654_not ; n20655
g20400 and b[32] n20222_not ; n20656
g20401 and n20220_not n20656 ; n20657
g20402 and n20224_not n20657_not ; n20658
g20403 and n20655_not n20658 ; n20659
g20404 and n20224_not n20659_not ; n20660
g20405 and b[33] n20213_not ; n20661
g20406 and n20211_not n20661 ; n20662
g20407 and n20215_not n20662_not ; n20663
g20408 and n20660_not n20663 ; n20664
g20409 and n20215_not n20664_not ; n20665
g20410 and b[34] n20204_not ; n20666
g20411 and n20202_not n20666 ; n20667
g20412 and n20206_not n20667_not ; n20668
g20413 and n20665_not n20668 ; n20669
g20414 and n20206_not n20669_not ; n20670
g20415 and b[35] n20195_not ; n20671
g20416 and n20193_not n20671 ; n20672
g20417 and n20197_not n20672_not ; n20673
g20418 and n20670_not n20673 ; n20674
g20419 and n20197_not n20674_not ; n20675
g20420 and b[36] n20186_not ; n20676
g20421 and n20184_not n20676 ; n20677
g20422 and n20188_not n20677_not ; n20678
g20423 and n20675_not n20678 ; n20679
g20424 and n20188_not n20679_not ; n20680
g20425 and b[37] n20177_not ; n20681
g20426 and n20175_not n20681 ; n20682
g20427 and n20179_not n20682_not ; n20683
g20428 and n20680_not n20683 ; n20684
g20429 and n20179_not n20684_not ; n20685
g20430 and b[38] n20168_not ; n20686
g20431 and n20166_not n20686 ; n20687
g20432 and n20170_not n20687_not ; n20688
g20433 and n20685_not n20688 ; n20689
g20434 and n20170_not n20689_not ; n20690
g20435 and b[39] n20159_not ; n20691
g20436 and n20157_not n20691 ; n20692
g20437 and n20161_not n20692_not ; n20693
g20438 and n20690_not n20693 ; n20694
g20439 and n20161_not n20694_not ; n20695
g20440 and b[40] n20150_not ; n20696
g20441 and n20148_not n20696 ; n20697
g20442 and n20152_not n20697_not ; n20698
g20443 and n20695_not n20698 ; n20699
g20444 and n20152_not n20699_not ; n20700
g20445 and b[41] n20141_not ; n20701
g20446 and n20139_not n20701 ; n20702
g20447 and n20143_not n20702_not ; n20703
g20448 and n20700_not n20703 ; n20704
g20449 and n20143_not n20704_not ; n20705
g20450 and b[42] n20132_not ; n20706
g20451 and n20130_not n20706 ; n20707
g20452 and n20134_not n20707_not ; n20708
g20453 and n20705_not n20708 ; n20709
g20454 and n20134_not n20709_not ; n20710
g20455 and b[43] n20123_not ; n20711
g20456 and n20121_not n20711 ; n20712
g20457 and n20125_not n20712_not ; n20713
g20458 and n20710_not n20713 ; n20714
g20459 and n20125_not n20714_not ; n20715
g20460 and b[44] n20114_not ; n20716
g20461 and n20112_not n20716 ; n20717
g20462 and n20116_not n20717_not ; n20718
g20463 and n20715_not n20718 ; n20719
g20464 and n20116_not n20719_not ; n20720
g20465 and b[45] n20105_not ; n20721
g20466 and n20103_not n20721 ; n20722
g20467 and n20107_not n20722_not ; n20723
g20468 and n20720_not n20723 ; n20724
g20469 and n20107_not n20724_not ; n20725
g20470 and b[46] n20096_not ; n20726
g20471 and n20094_not n20726 ; n20727
g20472 and n20098_not n20727_not ; n20728
g20473 and n20725_not n20728 ; n20729
g20474 and n20098_not n20729_not ; n20730
g20475 and b[47] n20087_not ; n20731
g20476 and n20085_not n20731 ; n20732
g20477 and n20089_not n20732_not ; n20733
g20478 and n20730_not n20733 ; n20734
g20479 and n20089_not n20734_not ; n20735
g20480 and b[48] n20078_not ; n20736
g20481 and n20076_not n20736 ; n20737
g20482 and n20080_not n20737_not ; n20738
g20483 and n20735_not n20738 ; n20739
g20484 and n20080_not n20739_not ; n20740
g20485 and b[49] n20069_not ; n20741
g20486 and n20067_not n20741 ; n20742
g20487 and n20071_not n20742_not ; n20743
g20488 and n20740_not n20743 ; n20744
g20489 and n20071_not n20744_not ; n20745
g20490 and b[50] n20060_not ; n20746
g20491 and n20058_not n20746 ; n20747
g20492 and n20062_not n20747_not ; n20748
g20493 and n20745_not n20748 ; n20749
g20494 and n20062_not n20749_not ; n20750
g20495 and b[51] n20051_not ; n20751
g20496 and n20049_not n20751 ; n20752
g20497 and n20053_not n20752_not ; n20753
g20498 and n20750_not n20753 ; n20754
g20499 and n20053_not n20754_not ; n20755
g20500 and b[52] n20042_not ; n20756
g20501 and n20040_not n20756 ; n20757
g20502 and n20044_not n20757_not ; n20758
g20503 and n20755_not n20758 ; n20759
g20504 and n20044_not n20759_not ; n20760
g20505 and n19313_not n20030_not ; n20761
g20506 and n20028_not n20761 ; n20762
g20507 and n20019_not n20762 ; n20763
g20508 and n20028_not n20030_not ; n20764
g20509 and n20020_not n20764_not ; n20765
g20510 and n20763_not n20765_not ; n20766
g20511 and quotient[11] n20766_not ; n20767
g20512 and n20027_not n20034_not ; n20768
g20513 and n20033_not n20768 ; n20769
g20514 and n20767_not n20769_not ; n20770
g20515 and b[53]_not n20770_not ; n20771
g20516 and b[53] n20769_not ; n20772
g20517 and n20767_not n20772 ; n20773
g20518 and n283 n285 ; n20774
g20519 and n280 n20774 ; n20775
g20520 and n20773_not n20775 ; n20776
g20521 and n20771_not n20776 ; n20777
g20522 and n20760_not n20777 ; n20778
g20523 and n595 n20770_not ; n20779
g20524 and n20778_not n20779_not ; quotient[10]
g20525 and n20053_not n20758 ; n20781
g20526 and n20754_not n20781 ; n20782
g20527 and n20755_not n20758_not ; n20783
g20528 and n20782_not n20783_not ; n20784
g20529 and quotient[10] n20784_not ; n20785
g20530 and n20043_not n20779_not ; n20786
g20531 and n20778_not n20786 ; n20787
g20532 and n20785_not n20787_not ; n20788
g20533 and n20044_not n20773_not ; n20789
g20534 and n20771_not n20789 ; n20790
g20535 and n20759_not n20790 ; n20791
g20536 and n20771_not n20773_not ; n20792
g20537 and n20760_not n20792_not ; n20793
g20538 and n20791_not n20793_not ; n20794
g20539 and quotient[10] n20794_not ; n20795
g20540 and n20770_not n20779_not ; n20796
g20541 and n20778_not n20796 ; n20797
g20542 and n20795_not n20797_not ; n20798
g20543 and b[54]_not n20798_not ; n20799
g20544 and b[53]_not n20788_not ; n20800
g20545 and n20062_not n20753 ; n20801
g20546 and n20749_not n20801 ; n20802
g20547 and n20750_not n20753_not ; n20803
g20548 and n20802_not n20803_not ; n20804
g20549 and quotient[10] n20804_not ; n20805
g20550 and n20052_not n20779_not ; n20806
g20551 and n20778_not n20806 ; n20807
g20552 and n20805_not n20807_not ; n20808
g20553 and b[52]_not n20808_not ; n20809
g20554 and n20071_not n20748 ; n20810
g20555 and n20744_not n20810 ; n20811
g20556 and n20745_not n20748_not ; n20812
g20557 and n20811_not n20812_not ; n20813
g20558 and quotient[10] n20813_not ; n20814
g20559 and n20061_not n20779_not ; n20815
g20560 and n20778_not n20815 ; n20816
g20561 and n20814_not n20816_not ; n20817
g20562 and b[51]_not n20817_not ; n20818
g20563 and n20080_not n20743 ; n20819
g20564 and n20739_not n20819 ; n20820
g20565 and n20740_not n20743_not ; n20821
g20566 and n20820_not n20821_not ; n20822
g20567 and quotient[10] n20822_not ; n20823
g20568 and n20070_not n20779_not ; n20824
g20569 and n20778_not n20824 ; n20825
g20570 and n20823_not n20825_not ; n20826
g20571 and b[50]_not n20826_not ; n20827
g20572 and n20089_not n20738 ; n20828
g20573 and n20734_not n20828 ; n20829
g20574 and n20735_not n20738_not ; n20830
g20575 and n20829_not n20830_not ; n20831
g20576 and quotient[10] n20831_not ; n20832
g20577 and n20079_not n20779_not ; n20833
g20578 and n20778_not n20833 ; n20834
g20579 and n20832_not n20834_not ; n20835
g20580 and b[49]_not n20835_not ; n20836
g20581 and n20098_not n20733 ; n20837
g20582 and n20729_not n20837 ; n20838
g20583 and n20730_not n20733_not ; n20839
g20584 and n20838_not n20839_not ; n20840
g20585 and quotient[10] n20840_not ; n20841
g20586 and n20088_not n20779_not ; n20842
g20587 and n20778_not n20842 ; n20843
g20588 and n20841_not n20843_not ; n20844
g20589 and b[48]_not n20844_not ; n20845
g20590 and n20107_not n20728 ; n20846
g20591 and n20724_not n20846 ; n20847
g20592 and n20725_not n20728_not ; n20848
g20593 and n20847_not n20848_not ; n20849
g20594 and quotient[10] n20849_not ; n20850
g20595 and n20097_not n20779_not ; n20851
g20596 and n20778_not n20851 ; n20852
g20597 and n20850_not n20852_not ; n20853
g20598 and b[47]_not n20853_not ; n20854
g20599 and n20116_not n20723 ; n20855
g20600 and n20719_not n20855 ; n20856
g20601 and n20720_not n20723_not ; n20857
g20602 and n20856_not n20857_not ; n20858
g20603 and quotient[10] n20858_not ; n20859
g20604 and n20106_not n20779_not ; n20860
g20605 and n20778_not n20860 ; n20861
g20606 and n20859_not n20861_not ; n20862
g20607 and b[46]_not n20862_not ; n20863
g20608 and n20125_not n20718 ; n20864
g20609 and n20714_not n20864 ; n20865
g20610 and n20715_not n20718_not ; n20866
g20611 and n20865_not n20866_not ; n20867
g20612 and quotient[10] n20867_not ; n20868
g20613 and n20115_not n20779_not ; n20869
g20614 and n20778_not n20869 ; n20870
g20615 and n20868_not n20870_not ; n20871
g20616 and b[45]_not n20871_not ; n20872
g20617 and n20134_not n20713 ; n20873
g20618 and n20709_not n20873 ; n20874
g20619 and n20710_not n20713_not ; n20875
g20620 and n20874_not n20875_not ; n20876
g20621 and quotient[10] n20876_not ; n20877
g20622 and n20124_not n20779_not ; n20878
g20623 and n20778_not n20878 ; n20879
g20624 and n20877_not n20879_not ; n20880
g20625 and b[44]_not n20880_not ; n20881
g20626 and n20143_not n20708 ; n20882
g20627 and n20704_not n20882 ; n20883
g20628 and n20705_not n20708_not ; n20884
g20629 and n20883_not n20884_not ; n20885
g20630 and quotient[10] n20885_not ; n20886
g20631 and n20133_not n20779_not ; n20887
g20632 and n20778_not n20887 ; n20888
g20633 and n20886_not n20888_not ; n20889
g20634 and b[43]_not n20889_not ; n20890
g20635 and n20152_not n20703 ; n20891
g20636 and n20699_not n20891 ; n20892
g20637 and n20700_not n20703_not ; n20893
g20638 and n20892_not n20893_not ; n20894
g20639 and quotient[10] n20894_not ; n20895
g20640 and n20142_not n20779_not ; n20896
g20641 and n20778_not n20896 ; n20897
g20642 and n20895_not n20897_not ; n20898
g20643 and b[42]_not n20898_not ; n20899
g20644 and n20161_not n20698 ; n20900
g20645 and n20694_not n20900 ; n20901
g20646 and n20695_not n20698_not ; n20902
g20647 and n20901_not n20902_not ; n20903
g20648 and quotient[10] n20903_not ; n20904
g20649 and n20151_not n20779_not ; n20905
g20650 and n20778_not n20905 ; n20906
g20651 and n20904_not n20906_not ; n20907
g20652 and b[41]_not n20907_not ; n20908
g20653 and n20170_not n20693 ; n20909
g20654 and n20689_not n20909 ; n20910
g20655 and n20690_not n20693_not ; n20911
g20656 and n20910_not n20911_not ; n20912
g20657 and quotient[10] n20912_not ; n20913
g20658 and n20160_not n20779_not ; n20914
g20659 and n20778_not n20914 ; n20915
g20660 and n20913_not n20915_not ; n20916
g20661 and b[40]_not n20916_not ; n20917
g20662 and n20179_not n20688 ; n20918
g20663 and n20684_not n20918 ; n20919
g20664 and n20685_not n20688_not ; n20920
g20665 and n20919_not n20920_not ; n20921
g20666 and quotient[10] n20921_not ; n20922
g20667 and n20169_not n20779_not ; n20923
g20668 and n20778_not n20923 ; n20924
g20669 and n20922_not n20924_not ; n20925
g20670 and b[39]_not n20925_not ; n20926
g20671 and n20188_not n20683 ; n20927
g20672 and n20679_not n20927 ; n20928
g20673 and n20680_not n20683_not ; n20929
g20674 and n20928_not n20929_not ; n20930
g20675 and quotient[10] n20930_not ; n20931
g20676 and n20178_not n20779_not ; n20932
g20677 and n20778_not n20932 ; n20933
g20678 and n20931_not n20933_not ; n20934
g20679 and b[38]_not n20934_not ; n20935
g20680 and n20197_not n20678 ; n20936
g20681 and n20674_not n20936 ; n20937
g20682 and n20675_not n20678_not ; n20938
g20683 and n20937_not n20938_not ; n20939
g20684 and quotient[10] n20939_not ; n20940
g20685 and n20187_not n20779_not ; n20941
g20686 and n20778_not n20941 ; n20942
g20687 and n20940_not n20942_not ; n20943
g20688 and b[37]_not n20943_not ; n20944
g20689 and n20206_not n20673 ; n20945
g20690 and n20669_not n20945 ; n20946
g20691 and n20670_not n20673_not ; n20947
g20692 and n20946_not n20947_not ; n20948
g20693 and quotient[10] n20948_not ; n20949
g20694 and n20196_not n20779_not ; n20950
g20695 and n20778_not n20950 ; n20951
g20696 and n20949_not n20951_not ; n20952
g20697 and b[36]_not n20952_not ; n20953
g20698 and n20215_not n20668 ; n20954
g20699 and n20664_not n20954 ; n20955
g20700 and n20665_not n20668_not ; n20956
g20701 and n20955_not n20956_not ; n20957
g20702 and quotient[10] n20957_not ; n20958
g20703 and n20205_not n20779_not ; n20959
g20704 and n20778_not n20959 ; n20960
g20705 and n20958_not n20960_not ; n20961
g20706 and b[35]_not n20961_not ; n20962
g20707 and n20224_not n20663 ; n20963
g20708 and n20659_not n20963 ; n20964
g20709 and n20660_not n20663_not ; n20965
g20710 and n20964_not n20965_not ; n20966
g20711 and quotient[10] n20966_not ; n20967
g20712 and n20214_not n20779_not ; n20968
g20713 and n20778_not n20968 ; n20969
g20714 and n20967_not n20969_not ; n20970
g20715 and b[34]_not n20970_not ; n20971
g20716 and n20233_not n20658 ; n20972
g20717 and n20654_not n20972 ; n20973
g20718 and n20655_not n20658_not ; n20974
g20719 and n20973_not n20974_not ; n20975
g20720 and quotient[10] n20975_not ; n20976
g20721 and n20223_not n20779_not ; n20977
g20722 and n20778_not n20977 ; n20978
g20723 and n20976_not n20978_not ; n20979
g20724 and b[33]_not n20979_not ; n20980
g20725 and n20242_not n20653 ; n20981
g20726 and n20649_not n20981 ; n20982
g20727 and n20650_not n20653_not ; n20983
g20728 and n20982_not n20983_not ; n20984
g20729 and quotient[10] n20984_not ; n20985
g20730 and n20232_not n20779_not ; n20986
g20731 and n20778_not n20986 ; n20987
g20732 and n20985_not n20987_not ; n20988
g20733 and b[32]_not n20988_not ; n20989
g20734 and n20251_not n20648 ; n20990
g20735 and n20644_not n20990 ; n20991
g20736 and n20645_not n20648_not ; n20992
g20737 and n20991_not n20992_not ; n20993
g20738 and quotient[10] n20993_not ; n20994
g20739 and n20241_not n20779_not ; n20995
g20740 and n20778_not n20995 ; n20996
g20741 and n20994_not n20996_not ; n20997
g20742 and b[31]_not n20997_not ; n20998
g20743 and n20260_not n20643 ; n20999
g20744 and n20639_not n20999 ; n21000
g20745 and n20640_not n20643_not ; n21001
g20746 and n21000_not n21001_not ; n21002
g20747 and quotient[10] n21002_not ; n21003
g20748 and n20250_not n20779_not ; n21004
g20749 and n20778_not n21004 ; n21005
g20750 and n21003_not n21005_not ; n21006
g20751 and b[30]_not n21006_not ; n21007
g20752 and n20269_not n20638 ; n21008
g20753 and n20634_not n21008 ; n21009
g20754 and n20635_not n20638_not ; n21010
g20755 and n21009_not n21010_not ; n21011
g20756 and quotient[10] n21011_not ; n21012
g20757 and n20259_not n20779_not ; n21013
g20758 and n20778_not n21013 ; n21014
g20759 and n21012_not n21014_not ; n21015
g20760 and b[29]_not n21015_not ; n21016
g20761 and n20278_not n20633 ; n21017
g20762 and n20629_not n21017 ; n21018
g20763 and n20630_not n20633_not ; n21019
g20764 and n21018_not n21019_not ; n21020
g20765 and quotient[10] n21020_not ; n21021
g20766 and n20268_not n20779_not ; n21022
g20767 and n20778_not n21022 ; n21023
g20768 and n21021_not n21023_not ; n21024
g20769 and b[28]_not n21024_not ; n21025
g20770 and n20287_not n20628 ; n21026
g20771 and n20624_not n21026 ; n21027
g20772 and n20625_not n20628_not ; n21028
g20773 and n21027_not n21028_not ; n21029
g20774 and quotient[10] n21029_not ; n21030
g20775 and n20277_not n20779_not ; n21031
g20776 and n20778_not n21031 ; n21032
g20777 and n21030_not n21032_not ; n21033
g20778 and b[27]_not n21033_not ; n21034
g20779 and n20296_not n20623 ; n21035
g20780 and n20619_not n21035 ; n21036
g20781 and n20620_not n20623_not ; n21037
g20782 and n21036_not n21037_not ; n21038
g20783 and quotient[10] n21038_not ; n21039
g20784 and n20286_not n20779_not ; n21040
g20785 and n20778_not n21040 ; n21041
g20786 and n21039_not n21041_not ; n21042
g20787 and b[26]_not n21042_not ; n21043
g20788 and n20305_not n20618 ; n21044
g20789 and n20614_not n21044 ; n21045
g20790 and n20615_not n20618_not ; n21046
g20791 and n21045_not n21046_not ; n21047
g20792 and quotient[10] n21047_not ; n21048
g20793 and n20295_not n20779_not ; n21049
g20794 and n20778_not n21049 ; n21050
g20795 and n21048_not n21050_not ; n21051
g20796 and b[25]_not n21051_not ; n21052
g20797 and n20314_not n20613 ; n21053
g20798 and n20609_not n21053 ; n21054
g20799 and n20610_not n20613_not ; n21055
g20800 and n21054_not n21055_not ; n21056
g20801 and quotient[10] n21056_not ; n21057
g20802 and n20304_not n20779_not ; n21058
g20803 and n20778_not n21058 ; n21059
g20804 and n21057_not n21059_not ; n21060
g20805 and b[24]_not n21060_not ; n21061
g20806 and n20323_not n20608 ; n21062
g20807 and n20604_not n21062 ; n21063
g20808 and n20605_not n20608_not ; n21064
g20809 and n21063_not n21064_not ; n21065
g20810 and quotient[10] n21065_not ; n21066
g20811 and n20313_not n20779_not ; n21067
g20812 and n20778_not n21067 ; n21068
g20813 and n21066_not n21068_not ; n21069
g20814 and b[23]_not n21069_not ; n21070
g20815 and n20332_not n20603 ; n21071
g20816 and n20599_not n21071 ; n21072
g20817 and n20600_not n20603_not ; n21073
g20818 and n21072_not n21073_not ; n21074
g20819 and quotient[10] n21074_not ; n21075
g20820 and n20322_not n20779_not ; n21076
g20821 and n20778_not n21076 ; n21077
g20822 and n21075_not n21077_not ; n21078
g20823 and b[22]_not n21078_not ; n21079
g20824 and n20341_not n20598 ; n21080
g20825 and n20594_not n21080 ; n21081
g20826 and n20595_not n20598_not ; n21082
g20827 and n21081_not n21082_not ; n21083
g20828 and quotient[10] n21083_not ; n21084
g20829 and n20331_not n20779_not ; n21085
g20830 and n20778_not n21085 ; n21086
g20831 and n21084_not n21086_not ; n21087
g20832 and b[21]_not n21087_not ; n21088
g20833 and n20350_not n20593 ; n21089
g20834 and n20589_not n21089 ; n21090
g20835 and n20590_not n20593_not ; n21091
g20836 and n21090_not n21091_not ; n21092
g20837 and quotient[10] n21092_not ; n21093
g20838 and n20340_not n20779_not ; n21094
g20839 and n20778_not n21094 ; n21095
g20840 and n21093_not n21095_not ; n21096
g20841 and b[20]_not n21096_not ; n21097
g20842 and n20359_not n20588 ; n21098
g20843 and n20584_not n21098 ; n21099
g20844 and n20585_not n20588_not ; n21100
g20845 and n21099_not n21100_not ; n21101
g20846 and quotient[10] n21101_not ; n21102
g20847 and n20349_not n20779_not ; n21103
g20848 and n20778_not n21103 ; n21104
g20849 and n21102_not n21104_not ; n21105
g20850 and b[19]_not n21105_not ; n21106
g20851 and n20368_not n20583 ; n21107
g20852 and n20579_not n21107 ; n21108
g20853 and n20580_not n20583_not ; n21109
g20854 and n21108_not n21109_not ; n21110
g20855 and quotient[10] n21110_not ; n21111
g20856 and n20358_not n20779_not ; n21112
g20857 and n20778_not n21112 ; n21113
g20858 and n21111_not n21113_not ; n21114
g20859 and b[18]_not n21114_not ; n21115
g20860 and n20377_not n20578 ; n21116
g20861 and n20574_not n21116 ; n21117
g20862 and n20575_not n20578_not ; n21118
g20863 and n21117_not n21118_not ; n21119
g20864 and quotient[10] n21119_not ; n21120
g20865 and n20367_not n20779_not ; n21121
g20866 and n20778_not n21121 ; n21122
g20867 and n21120_not n21122_not ; n21123
g20868 and b[17]_not n21123_not ; n21124
g20869 and n20386_not n20573 ; n21125
g20870 and n20569_not n21125 ; n21126
g20871 and n20570_not n20573_not ; n21127
g20872 and n21126_not n21127_not ; n21128
g20873 and quotient[10] n21128_not ; n21129
g20874 and n20376_not n20779_not ; n21130
g20875 and n20778_not n21130 ; n21131
g20876 and n21129_not n21131_not ; n21132
g20877 and b[16]_not n21132_not ; n21133
g20878 and n20395_not n20568 ; n21134
g20879 and n20564_not n21134 ; n21135
g20880 and n20565_not n20568_not ; n21136
g20881 and n21135_not n21136_not ; n21137
g20882 and quotient[10] n21137_not ; n21138
g20883 and n20385_not n20779_not ; n21139
g20884 and n20778_not n21139 ; n21140
g20885 and n21138_not n21140_not ; n21141
g20886 and b[15]_not n21141_not ; n21142
g20887 and n20404_not n20563 ; n21143
g20888 and n20559_not n21143 ; n21144
g20889 and n20560_not n20563_not ; n21145
g20890 and n21144_not n21145_not ; n21146
g20891 and quotient[10] n21146_not ; n21147
g20892 and n20394_not n20779_not ; n21148
g20893 and n20778_not n21148 ; n21149
g20894 and n21147_not n21149_not ; n21150
g20895 and b[14]_not n21150_not ; n21151
g20896 and n20413_not n20558 ; n21152
g20897 and n20554_not n21152 ; n21153
g20898 and n20555_not n20558_not ; n21154
g20899 and n21153_not n21154_not ; n21155
g20900 and quotient[10] n21155_not ; n21156
g20901 and n20403_not n20779_not ; n21157
g20902 and n20778_not n21157 ; n21158
g20903 and n21156_not n21158_not ; n21159
g20904 and b[13]_not n21159_not ; n21160
g20905 and n20422_not n20553 ; n21161
g20906 and n20549_not n21161 ; n21162
g20907 and n20550_not n20553_not ; n21163
g20908 and n21162_not n21163_not ; n21164
g20909 and quotient[10] n21164_not ; n21165
g20910 and n20412_not n20779_not ; n21166
g20911 and n20778_not n21166 ; n21167
g20912 and n21165_not n21167_not ; n21168
g20913 and b[12]_not n21168_not ; n21169
g20914 and n20431_not n20548 ; n21170
g20915 and n20544_not n21170 ; n21171
g20916 and n20545_not n20548_not ; n21172
g20917 and n21171_not n21172_not ; n21173
g20918 and quotient[10] n21173_not ; n21174
g20919 and n20421_not n20779_not ; n21175
g20920 and n20778_not n21175 ; n21176
g20921 and n21174_not n21176_not ; n21177
g20922 and b[11]_not n21177_not ; n21178
g20923 and n20440_not n20543 ; n21179
g20924 and n20539_not n21179 ; n21180
g20925 and n20540_not n20543_not ; n21181
g20926 and n21180_not n21181_not ; n21182
g20927 and quotient[10] n21182_not ; n21183
g20928 and n20430_not n20779_not ; n21184
g20929 and n20778_not n21184 ; n21185
g20930 and n21183_not n21185_not ; n21186
g20931 and b[10]_not n21186_not ; n21187
g20932 and n20449_not n20538 ; n21188
g20933 and n20534_not n21188 ; n21189
g20934 and n20535_not n20538_not ; n21190
g20935 and n21189_not n21190_not ; n21191
g20936 and quotient[10] n21191_not ; n21192
g20937 and n20439_not n20779_not ; n21193
g20938 and n20778_not n21193 ; n21194
g20939 and n21192_not n21194_not ; n21195
g20940 and b[9]_not n21195_not ; n21196
g20941 and n20458_not n20533 ; n21197
g20942 and n20529_not n21197 ; n21198
g20943 and n20530_not n20533_not ; n21199
g20944 and n21198_not n21199_not ; n21200
g20945 and quotient[10] n21200_not ; n21201
g20946 and n20448_not n20779_not ; n21202
g20947 and n20778_not n21202 ; n21203
g20948 and n21201_not n21203_not ; n21204
g20949 and b[8]_not n21204_not ; n21205
g20950 and n20467_not n20528 ; n21206
g20951 and n20524_not n21206 ; n21207
g20952 and n20525_not n20528_not ; n21208
g20953 and n21207_not n21208_not ; n21209
g20954 and quotient[10] n21209_not ; n21210
g20955 and n20457_not n20779_not ; n21211
g20956 and n20778_not n21211 ; n21212
g20957 and n21210_not n21212_not ; n21213
g20958 and b[7]_not n21213_not ; n21214
g20959 and n20476_not n20523 ; n21215
g20960 and n20519_not n21215 ; n21216
g20961 and n20520_not n20523_not ; n21217
g20962 and n21216_not n21217_not ; n21218
g20963 and quotient[10] n21218_not ; n21219
g20964 and n20466_not n20779_not ; n21220
g20965 and n20778_not n21220 ; n21221
g20966 and n21219_not n21221_not ; n21222
g20967 and b[6]_not n21222_not ; n21223
g20968 and n20485_not n20518 ; n21224
g20969 and n20514_not n21224 ; n21225
g20970 and n20515_not n20518_not ; n21226
g20971 and n21225_not n21226_not ; n21227
g20972 and quotient[10] n21227_not ; n21228
g20973 and n20475_not n20779_not ; n21229
g20974 and n20778_not n21229 ; n21230
g20975 and n21228_not n21230_not ; n21231
g20976 and b[5]_not n21231_not ; n21232
g20977 and n20493_not n20513 ; n21233
g20978 and n20509_not n21233 ; n21234
g20979 and n20510_not n20513_not ; n21235
g20980 and n21234_not n21235_not ; n21236
g20981 and quotient[10] n21236_not ; n21237
g20982 and n20484_not n20779_not ; n21238
g20983 and n20778_not n21238 ; n21239
g20984 and n21237_not n21239_not ; n21240
g20985 and b[4]_not n21240_not ; n21241
g20986 and n20504_not n20508 ; n21242
g20987 and n20503_not n21242 ; n21243
g20988 and n20505_not n20508_not ; n21244
g20989 and n21243_not n21244_not ; n21245
g20990 and quotient[10] n21245_not ; n21246
g20991 and n20492_not n20779_not ; n21247
g20992 and n20778_not n21247 ; n21248
g20993 and n21246_not n21248_not ; n21249
g20994 and b[3]_not n21249_not ; n21250
g20995 and n20500_not n20502 ; n21251
g20996 and n20498_not n21251 ; n21252
g20997 and n20503_not n21252_not ; n21253
g20998 and quotient[10] n21253 ; n21254
g20999 and n20497_not n20779_not ; n21255
g21000 and n20778_not n21255 ; n21256
g21001 and n21254_not n21256_not ; n21257
g21002 and b[2]_not n21257_not ; n21258
g21003 and b[0] quotient[10] ; n21259
g21004 and a[10] n21259_not ; n21260
g21005 and n20502 quotient[10] ; n21261
g21006 and n21260_not n21261_not ; n21262
g21007 and b[1] n21262_not ; n21263
g21008 and b[1]_not n21261_not ; n21264
g21009 and n21260_not n21264 ; n21265
g21010 and n21263_not n21265_not ; n21266
g21011 and a[9]_not b[0] ; n21267
g21012 and n21266_not n21267_not ; n21268
g21013 and b[1]_not n21262_not ; n21269
g21014 and n21268_not n21269_not ; n21270
g21015 and b[2] n21256_not ; n21271
g21016 and n21254_not n21271 ; n21272
g21017 and n21258_not n21272_not ; n21273
g21018 and n21270_not n21273 ; n21274
g21019 and n21258_not n21274_not ; n21275
g21020 and b[3] n21248_not ; n21276
g21021 and n21246_not n21276 ; n21277
g21022 and n21250_not n21277_not ; n21278
g21023 and n21275_not n21278 ; n21279
g21024 and n21250_not n21279_not ; n21280
g21025 and b[4] n21239_not ; n21281
g21026 and n21237_not n21281 ; n21282
g21027 and n21241_not n21282_not ; n21283
g21028 and n21280_not n21283 ; n21284
g21029 and n21241_not n21284_not ; n21285
g21030 and b[5] n21230_not ; n21286
g21031 and n21228_not n21286 ; n21287
g21032 and n21232_not n21287_not ; n21288
g21033 and n21285_not n21288 ; n21289
g21034 and n21232_not n21289_not ; n21290
g21035 and b[6] n21221_not ; n21291
g21036 and n21219_not n21291 ; n21292
g21037 and n21223_not n21292_not ; n21293
g21038 and n21290_not n21293 ; n21294
g21039 and n21223_not n21294_not ; n21295
g21040 and b[7] n21212_not ; n21296
g21041 and n21210_not n21296 ; n21297
g21042 and n21214_not n21297_not ; n21298
g21043 and n21295_not n21298 ; n21299
g21044 and n21214_not n21299_not ; n21300
g21045 and b[8] n21203_not ; n21301
g21046 and n21201_not n21301 ; n21302
g21047 and n21205_not n21302_not ; n21303
g21048 and n21300_not n21303 ; n21304
g21049 and n21205_not n21304_not ; n21305
g21050 and b[9] n21194_not ; n21306
g21051 and n21192_not n21306 ; n21307
g21052 and n21196_not n21307_not ; n21308
g21053 and n21305_not n21308 ; n21309
g21054 and n21196_not n21309_not ; n21310
g21055 and b[10] n21185_not ; n21311
g21056 and n21183_not n21311 ; n21312
g21057 and n21187_not n21312_not ; n21313
g21058 and n21310_not n21313 ; n21314
g21059 and n21187_not n21314_not ; n21315
g21060 and b[11] n21176_not ; n21316
g21061 and n21174_not n21316 ; n21317
g21062 and n21178_not n21317_not ; n21318
g21063 and n21315_not n21318 ; n21319
g21064 and n21178_not n21319_not ; n21320
g21065 and b[12] n21167_not ; n21321
g21066 and n21165_not n21321 ; n21322
g21067 and n21169_not n21322_not ; n21323
g21068 and n21320_not n21323 ; n21324
g21069 and n21169_not n21324_not ; n21325
g21070 and b[13] n21158_not ; n21326
g21071 and n21156_not n21326 ; n21327
g21072 and n21160_not n21327_not ; n21328
g21073 and n21325_not n21328 ; n21329
g21074 and n21160_not n21329_not ; n21330
g21075 and b[14] n21149_not ; n21331
g21076 and n21147_not n21331 ; n21332
g21077 and n21151_not n21332_not ; n21333
g21078 and n21330_not n21333 ; n21334
g21079 and n21151_not n21334_not ; n21335
g21080 and b[15] n21140_not ; n21336
g21081 and n21138_not n21336 ; n21337
g21082 and n21142_not n21337_not ; n21338
g21083 and n21335_not n21338 ; n21339
g21084 and n21142_not n21339_not ; n21340
g21085 and b[16] n21131_not ; n21341
g21086 and n21129_not n21341 ; n21342
g21087 and n21133_not n21342_not ; n21343
g21088 and n21340_not n21343 ; n21344
g21089 and n21133_not n21344_not ; n21345
g21090 and b[17] n21122_not ; n21346
g21091 and n21120_not n21346 ; n21347
g21092 and n21124_not n21347_not ; n21348
g21093 and n21345_not n21348 ; n21349
g21094 and n21124_not n21349_not ; n21350
g21095 and b[18] n21113_not ; n21351
g21096 and n21111_not n21351 ; n21352
g21097 and n21115_not n21352_not ; n21353
g21098 and n21350_not n21353 ; n21354
g21099 and n21115_not n21354_not ; n21355
g21100 and b[19] n21104_not ; n21356
g21101 and n21102_not n21356 ; n21357
g21102 and n21106_not n21357_not ; n21358
g21103 and n21355_not n21358 ; n21359
g21104 and n21106_not n21359_not ; n21360
g21105 and b[20] n21095_not ; n21361
g21106 and n21093_not n21361 ; n21362
g21107 and n21097_not n21362_not ; n21363
g21108 and n21360_not n21363 ; n21364
g21109 and n21097_not n21364_not ; n21365
g21110 and b[21] n21086_not ; n21366
g21111 and n21084_not n21366 ; n21367
g21112 and n21088_not n21367_not ; n21368
g21113 and n21365_not n21368 ; n21369
g21114 and n21088_not n21369_not ; n21370
g21115 and b[22] n21077_not ; n21371
g21116 and n21075_not n21371 ; n21372
g21117 and n21079_not n21372_not ; n21373
g21118 and n21370_not n21373 ; n21374
g21119 and n21079_not n21374_not ; n21375
g21120 and b[23] n21068_not ; n21376
g21121 and n21066_not n21376 ; n21377
g21122 and n21070_not n21377_not ; n21378
g21123 and n21375_not n21378 ; n21379
g21124 and n21070_not n21379_not ; n21380
g21125 and b[24] n21059_not ; n21381
g21126 and n21057_not n21381 ; n21382
g21127 and n21061_not n21382_not ; n21383
g21128 and n21380_not n21383 ; n21384
g21129 and n21061_not n21384_not ; n21385
g21130 and b[25] n21050_not ; n21386
g21131 and n21048_not n21386 ; n21387
g21132 and n21052_not n21387_not ; n21388
g21133 and n21385_not n21388 ; n21389
g21134 and n21052_not n21389_not ; n21390
g21135 and b[26] n21041_not ; n21391
g21136 and n21039_not n21391 ; n21392
g21137 and n21043_not n21392_not ; n21393
g21138 and n21390_not n21393 ; n21394
g21139 and n21043_not n21394_not ; n21395
g21140 and b[27] n21032_not ; n21396
g21141 and n21030_not n21396 ; n21397
g21142 and n21034_not n21397_not ; n21398
g21143 and n21395_not n21398 ; n21399
g21144 and n21034_not n21399_not ; n21400
g21145 and b[28] n21023_not ; n21401
g21146 and n21021_not n21401 ; n21402
g21147 and n21025_not n21402_not ; n21403
g21148 and n21400_not n21403 ; n21404
g21149 and n21025_not n21404_not ; n21405
g21150 and b[29] n21014_not ; n21406
g21151 and n21012_not n21406 ; n21407
g21152 and n21016_not n21407_not ; n21408
g21153 and n21405_not n21408 ; n21409
g21154 and n21016_not n21409_not ; n21410
g21155 and b[30] n21005_not ; n21411
g21156 and n21003_not n21411 ; n21412
g21157 and n21007_not n21412_not ; n21413
g21158 and n21410_not n21413 ; n21414
g21159 and n21007_not n21414_not ; n21415
g21160 and b[31] n20996_not ; n21416
g21161 and n20994_not n21416 ; n21417
g21162 and n20998_not n21417_not ; n21418
g21163 and n21415_not n21418 ; n21419
g21164 and n20998_not n21419_not ; n21420
g21165 and b[32] n20987_not ; n21421
g21166 and n20985_not n21421 ; n21422
g21167 and n20989_not n21422_not ; n21423
g21168 and n21420_not n21423 ; n21424
g21169 and n20989_not n21424_not ; n21425
g21170 and b[33] n20978_not ; n21426
g21171 and n20976_not n21426 ; n21427
g21172 and n20980_not n21427_not ; n21428
g21173 and n21425_not n21428 ; n21429
g21174 and n20980_not n21429_not ; n21430
g21175 and b[34] n20969_not ; n21431
g21176 and n20967_not n21431 ; n21432
g21177 and n20971_not n21432_not ; n21433
g21178 and n21430_not n21433 ; n21434
g21179 and n20971_not n21434_not ; n21435
g21180 and b[35] n20960_not ; n21436
g21181 and n20958_not n21436 ; n21437
g21182 and n20962_not n21437_not ; n21438
g21183 and n21435_not n21438 ; n21439
g21184 and n20962_not n21439_not ; n21440
g21185 and b[36] n20951_not ; n21441
g21186 and n20949_not n21441 ; n21442
g21187 and n20953_not n21442_not ; n21443
g21188 and n21440_not n21443 ; n21444
g21189 and n20953_not n21444_not ; n21445
g21190 and b[37] n20942_not ; n21446
g21191 and n20940_not n21446 ; n21447
g21192 and n20944_not n21447_not ; n21448
g21193 and n21445_not n21448 ; n21449
g21194 and n20944_not n21449_not ; n21450
g21195 and b[38] n20933_not ; n21451
g21196 and n20931_not n21451 ; n21452
g21197 and n20935_not n21452_not ; n21453
g21198 and n21450_not n21453 ; n21454
g21199 and n20935_not n21454_not ; n21455
g21200 and b[39] n20924_not ; n21456
g21201 and n20922_not n21456 ; n21457
g21202 and n20926_not n21457_not ; n21458
g21203 and n21455_not n21458 ; n21459
g21204 and n20926_not n21459_not ; n21460
g21205 and b[40] n20915_not ; n21461
g21206 and n20913_not n21461 ; n21462
g21207 and n20917_not n21462_not ; n21463
g21208 and n21460_not n21463 ; n21464
g21209 and n20917_not n21464_not ; n21465
g21210 and b[41] n20906_not ; n21466
g21211 and n20904_not n21466 ; n21467
g21212 and n20908_not n21467_not ; n21468
g21213 and n21465_not n21468 ; n21469
g21214 and n20908_not n21469_not ; n21470
g21215 and b[42] n20897_not ; n21471
g21216 and n20895_not n21471 ; n21472
g21217 and n20899_not n21472_not ; n21473
g21218 and n21470_not n21473 ; n21474
g21219 and n20899_not n21474_not ; n21475
g21220 and b[43] n20888_not ; n21476
g21221 and n20886_not n21476 ; n21477
g21222 and n20890_not n21477_not ; n21478
g21223 and n21475_not n21478 ; n21479
g21224 and n20890_not n21479_not ; n21480
g21225 and b[44] n20879_not ; n21481
g21226 and n20877_not n21481 ; n21482
g21227 and n20881_not n21482_not ; n21483
g21228 and n21480_not n21483 ; n21484
g21229 and n20881_not n21484_not ; n21485
g21230 and b[45] n20870_not ; n21486
g21231 and n20868_not n21486 ; n21487
g21232 and n20872_not n21487_not ; n21488
g21233 and n21485_not n21488 ; n21489
g21234 and n20872_not n21489_not ; n21490
g21235 and b[46] n20861_not ; n21491
g21236 and n20859_not n21491 ; n21492
g21237 and n20863_not n21492_not ; n21493
g21238 and n21490_not n21493 ; n21494
g21239 and n20863_not n21494_not ; n21495
g21240 and b[47] n20852_not ; n21496
g21241 and n20850_not n21496 ; n21497
g21242 and n20854_not n21497_not ; n21498
g21243 and n21495_not n21498 ; n21499
g21244 and n20854_not n21499_not ; n21500
g21245 and b[48] n20843_not ; n21501
g21246 and n20841_not n21501 ; n21502
g21247 and n20845_not n21502_not ; n21503
g21248 and n21500_not n21503 ; n21504
g21249 and n20845_not n21504_not ; n21505
g21250 and b[49] n20834_not ; n21506
g21251 and n20832_not n21506 ; n21507
g21252 and n20836_not n21507_not ; n21508
g21253 and n21505_not n21508 ; n21509
g21254 and n20836_not n21509_not ; n21510
g21255 and b[50] n20825_not ; n21511
g21256 and n20823_not n21511 ; n21512
g21257 and n20827_not n21512_not ; n21513
g21258 and n21510_not n21513 ; n21514
g21259 and n20827_not n21514_not ; n21515
g21260 and b[51] n20816_not ; n21516
g21261 and n20814_not n21516 ; n21517
g21262 and n20818_not n21517_not ; n21518
g21263 and n21515_not n21518 ; n21519
g21264 and n20818_not n21519_not ; n21520
g21265 and b[52] n20807_not ; n21521
g21266 and n20805_not n21521 ; n21522
g21267 and n20809_not n21522_not ; n21523
g21268 and n21520_not n21523 ; n21524
g21269 and n20809_not n21524_not ; n21525
g21270 and b[53] n20787_not ; n21526
g21271 and n20785_not n21526 ; n21527
g21272 and n20800_not n21527_not ; n21528
g21273 and n21525_not n21528 ; n21529
g21274 and n20800_not n21529_not ; n21530
g21275 and b[54] n20797_not ; n21531
g21276 and n20795_not n21531 ; n21532
g21277 and n20799_not n21532_not ; n21533
g21278 and n21530_not n21533 ; n21534
g21279 and n20799_not n21534_not ; n21535
g21280 and n396 n406 ; n21536
g21281 and n403 n21536 ; n21537
g21282 and n21535_not n21537 ; quotient[9]
g21283 and n20788_not quotient[9]_not ; n21539
g21284 and n20809_not n21528 ; n21540
g21285 and n21524_not n21540 ; n21541
g21286 and n21525_not n21528_not ; n21542
g21287 and n21541_not n21542_not ; n21543
g21288 and n21537 n21543_not ; n21544
g21289 and n21535_not n21544 ; n21545
g21290 and n21539_not n21545_not ; n21546
g21291 and b[54]_not n21546_not ; n21547
g21292 and n20808_not quotient[9]_not ; n21548
g21293 and n20818_not n21523 ; n21549
g21294 and n21519_not n21549 ; n21550
g21295 and n21520_not n21523_not ; n21551
g21296 and n21550_not n21551_not ; n21552
g21297 and n21537 n21552_not ; n21553
g21298 and n21535_not n21553 ; n21554
g21299 and n21548_not n21554_not ; n21555
g21300 and b[53]_not n21555_not ; n21556
g21301 and n20817_not quotient[9]_not ; n21557
g21302 and n20827_not n21518 ; n21558
g21303 and n21514_not n21558 ; n21559
g21304 and n21515_not n21518_not ; n21560
g21305 and n21559_not n21560_not ; n21561
g21306 and n21537 n21561_not ; n21562
g21307 and n21535_not n21562 ; n21563
g21308 and n21557_not n21563_not ; n21564
g21309 and b[52]_not n21564_not ; n21565
g21310 and n20826_not quotient[9]_not ; n21566
g21311 and n20836_not n21513 ; n21567
g21312 and n21509_not n21567 ; n21568
g21313 and n21510_not n21513_not ; n21569
g21314 and n21568_not n21569_not ; n21570
g21315 and n21537 n21570_not ; n21571
g21316 and n21535_not n21571 ; n21572
g21317 and n21566_not n21572_not ; n21573
g21318 and b[51]_not n21573_not ; n21574
g21319 and n20835_not quotient[9]_not ; n21575
g21320 and n20845_not n21508 ; n21576
g21321 and n21504_not n21576 ; n21577
g21322 and n21505_not n21508_not ; n21578
g21323 and n21577_not n21578_not ; n21579
g21324 and n21537 n21579_not ; n21580
g21325 and n21535_not n21580 ; n21581
g21326 and n21575_not n21581_not ; n21582
g21327 and b[50]_not n21582_not ; n21583
g21328 and n20844_not quotient[9]_not ; n21584
g21329 and n20854_not n21503 ; n21585
g21330 and n21499_not n21585 ; n21586
g21331 and n21500_not n21503_not ; n21587
g21332 and n21586_not n21587_not ; n21588
g21333 and n21537 n21588_not ; n21589
g21334 and n21535_not n21589 ; n21590
g21335 and n21584_not n21590_not ; n21591
g21336 and b[49]_not n21591_not ; n21592
g21337 and n20853_not quotient[9]_not ; n21593
g21338 and n20863_not n21498 ; n21594
g21339 and n21494_not n21594 ; n21595
g21340 and n21495_not n21498_not ; n21596
g21341 and n21595_not n21596_not ; n21597
g21342 and n21537 n21597_not ; n21598
g21343 and n21535_not n21598 ; n21599
g21344 and n21593_not n21599_not ; n21600
g21345 and b[48]_not n21600_not ; n21601
g21346 and n20862_not quotient[9]_not ; n21602
g21347 and n20872_not n21493 ; n21603
g21348 and n21489_not n21603 ; n21604
g21349 and n21490_not n21493_not ; n21605
g21350 and n21604_not n21605_not ; n21606
g21351 and n21537 n21606_not ; n21607
g21352 and n21535_not n21607 ; n21608
g21353 and n21602_not n21608_not ; n21609
g21354 and b[47]_not n21609_not ; n21610
g21355 and n20871_not quotient[9]_not ; n21611
g21356 and n20881_not n21488 ; n21612
g21357 and n21484_not n21612 ; n21613
g21358 and n21485_not n21488_not ; n21614
g21359 and n21613_not n21614_not ; n21615
g21360 and n21537 n21615_not ; n21616
g21361 and n21535_not n21616 ; n21617
g21362 and n21611_not n21617_not ; n21618
g21363 and b[46]_not n21618_not ; n21619
g21364 and n20880_not quotient[9]_not ; n21620
g21365 and n20890_not n21483 ; n21621
g21366 and n21479_not n21621 ; n21622
g21367 and n21480_not n21483_not ; n21623
g21368 and n21622_not n21623_not ; n21624
g21369 and n21537 n21624_not ; n21625
g21370 and n21535_not n21625 ; n21626
g21371 and n21620_not n21626_not ; n21627
g21372 and b[45]_not n21627_not ; n21628
g21373 and n20889_not quotient[9]_not ; n21629
g21374 and n20899_not n21478 ; n21630
g21375 and n21474_not n21630 ; n21631
g21376 and n21475_not n21478_not ; n21632
g21377 and n21631_not n21632_not ; n21633
g21378 and n21537 n21633_not ; n21634
g21379 and n21535_not n21634 ; n21635
g21380 and n21629_not n21635_not ; n21636
g21381 and b[44]_not n21636_not ; n21637
g21382 and n20898_not quotient[9]_not ; n21638
g21383 and n20908_not n21473 ; n21639
g21384 and n21469_not n21639 ; n21640
g21385 and n21470_not n21473_not ; n21641
g21386 and n21640_not n21641_not ; n21642
g21387 and n21537 n21642_not ; n21643
g21388 and n21535_not n21643 ; n21644
g21389 and n21638_not n21644_not ; n21645
g21390 and b[43]_not n21645_not ; n21646
g21391 and n20907_not quotient[9]_not ; n21647
g21392 and n20917_not n21468 ; n21648
g21393 and n21464_not n21648 ; n21649
g21394 and n21465_not n21468_not ; n21650
g21395 and n21649_not n21650_not ; n21651
g21396 and n21537 n21651_not ; n21652
g21397 and n21535_not n21652 ; n21653
g21398 and n21647_not n21653_not ; n21654
g21399 and b[42]_not n21654_not ; n21655
g21400 and n20916_not quotient[9]_not ; n21656
g21401 and n20926_not n21463 ; n21657
g21402 and n21459_not n21657 ; n21658
g21403 and n21460_not n21463_not ; n21659
g21404 and n21658_not n21659_not ; n21660
g21405 and n21537 n21660_not ; n21661
g21406 and n21535_not n21661 ; n21662
g21407 and n21656_not n21662_not ; n21663
g21408 and b[41]_not n21663_not ; n21664
g21409 and n20925_not quotient[9]_not ; n21665
g21410 and n20935_not n21458 ; n21666
g21411 and n21454_not n21666 ; n21667
g21412 and n21455_not n21458_not ; n21668
g21413 and n21667_not n21668_not ; n21669
g21414 and n21537 n21669_not ; n21670
g21415 and n21535_not n21670 ; n21671
g21416 and n21665_not n21671_not ; n21672
g21417 and b[40]_not n21672_not ; n21673
g21418 and n20934_not quotient[9]_not ; n21674
g21419 and n20944_not n21453 ; n21675
g21420 and n21449_not n21675 ; n21676
g21421 and n21450_not n21453_not ; n21677
g21422 and n21676_not n21677_not ; n21678
g21423 and n21537 n21678_not ; n21679
g21424 and n21535_not n21679 ; n21680
g21425 and n21674_not n21680_not ; n21681
g21426 and b[39]_not n21681_not ; n21682
g21427 and n20943_not quotient[9]_not ; n21683
g21428 and n20953_not n21448 ; n21684
g21429 and n21444_not n21684 ; n21685
g21430 and n21445_not n21448_not ; n21686
g21431 and n21685_not n21686_not ; n21687
g21432 and n21537 n21687_not ; n21688
g21433 and n21535_not n21688 ; n21689
g21434 and n21683_not n21689_not ; n21690
g21435 and b[38]_not n21690_not ; n21691
g21436 and n20952_not quotient[9]_not ; n21692
g21437 and n20962_not n21443 ; n21693
g21438 and n21439_not n21693 ; n21694
g21439 and n21440_not n21443_not ; n21695
g21440 and n21694_not n21695_not ; n21696
g21441 and n21537 n21696_not ; n21697
g21442 and n21535_not n21697 ; n21698
g21443 and n21692_not n21698_not ; n21699
g21444 and b[37]_not n21699_not ; n21700
g21445 and n20961_not quotient[9]_not ; n21701
g21446 and n20971_not n21438 ; n21702
g21447 and n21434_not n21702 ; n21703
g21448 and n21435_not n21438_not ; n21704
g21449 and n21703_not n21704_not ; n21705
g21450 and n21537 n21705_not ; n21706
g21451 and n21535_not n21706 ; n21707
g21452 and n21701_not n21707_not ; n21708
g21453 and b[36]_not n21708_not ; n21709
g21454 and n20970_not quotient[9]_not ; n21710
g21455 and n20980_not n21433 ; n21711
g21456 and n21429_not n21711 ; n21712
g21457 and n21430_not n21433_not ; n21713
g21458 and n21712_not n21713_not ; n21714
g21459 and n21537 n21714_not ; n21715
g21460 and n21535_not n21715 ; n21716
g21461 and n21710_not n21716_not ; n21717
g21462 and b[35]_not n21717_not ; n21718
g21463 and n20979_not quotient[9]_not ; n21719
g21464 and n20989_not n21428 ; n21720
g21465 and n21424_not n21720 ; n21721
g21466 and n21425_not n21428_not ; n21722
g21467 and n21721_not n21722_not ; n21723
g21468 and n21537 n21723_not ; n21724
g21469 and n21535_not n21724 ; n21725
g21470 and n21719_not n21725_not ; n21726
g21471 and b[34]_not n21726_not ; n21727
g21472 and n20988_not quotient[9]_not ; n21728
g21473 and n20998_not n21423 ; n21729
g21474 and n21419_not n21729 ; n21730
g21475 and n21420_not n21423_not ; n21731
g21476 and n21730_not n21731_not ; n21732
g21477 and n21537 n21732_not ; n21733
g21478 and n21535_not n21733 ; n21734
g21479 and n21728_not n21734_not ; n21735
g21480 and b[33]_not n21735_not ; n21736
g21481 and n20997_not quotient[9]_not ; n21737
g21482 and n21007_not n21418 ; n21738
g21483 and n21414_not n21738 ; n21739
g21484 and n21415_not n21418_not ; n21740
g21485 and n21739_not n21740_not ; n21741
g21486 and n21537 n21741_not ; n21742
g21487 and n21535_not n21742 ; n21743
g21488 and n21737_not n21743_not ; n21744
g21489 and b[32]_not n21744_not ; n21745
g21490 and n21006_not quotient[9]_not ; n21746
g21491 and n21016_not n21413 ; n21747
g21492 and n21409_not n21747 ; n21748
g21493 and n21410_not n21413_not ; n21749
g21494 and n21748_not n21749_not ; n21750
g21495 and n21537 n21750_not ; n21751
g21496 and n21535_not n21751 ; n21752
g21497 and n21746_not n21752_not ; n21753
g21498 and b[31]_not n21753_not ; n21754
g21499 and n21015_not quotient[9]_not ; n21755
g21500 and n21025_not n21408 ; n21756
g21501 and n21404_not n21756 ; n21757
g21502 and n21405_not n21408_not ; n21758
g21503 and n21757_not n21758_not ; n21759
g21504 and n21537 n21759_not ; n21760
g21505 and n21535_not n21760 ; n21761
g21506 and n21755_not n21761_not ; n21762
g21507 and b[30]_not n21762_not ; n21763
g21508 and n21024_not quotient[9]_not ; n21764
g21509 and n21034_not n21403 ; n21765
g21510 and n21399_not n21765 ; n21766
g21511 and n21400_not n21403_not ; n21767
g21512 and n21766_not n21767_not ; n21768
g21513 and n21537 n21768_not ; n21769
g21514 and n21535_not n21769 ; n21770
g21515 and n21764_not n21770_not ; n21771
g21516 and b[29]_not n21771_not ; n21772
g21517 and n21033_not quotient[9]_not ; n21773
g21518 and n21043_not n21398 ; n21774
g21519 and n21394_not n21774 ; n21775
g21520 and n21395_not n21398_not ; n21776
g21521 and n21775_not n21776_not ; n21777
g21522 and n21537 n21777_not ; n21778
g21523 and n21535_not n21778 ; n21779
g21524 and n21773_not n21779_not ; n21780
g21525 and b[28]_not n21780_not ; n21781
g21526 and n21042_not quotient[9]_not ; n21782
g21527 and n21052_not n21393 ; n21783
g21528 and n21389_not n21783 ; n21784
g21529 and n21390_not n21393_not ; n21785
g21530 and n21784_not n21785_not ; n21786
g21531 and n21537 n21786_not ; n21787
g21532 and n21535_not n21787 ; n21788
g21533 and n21782_not n21788_not ; n21789
g21534 and b[27]_not n21789_not ; n21790
g21535 and n21051_not quotient[9]_not ; n21791
g21536 and n21061_not n21388 ; n21792
g21537 and n21384_not n21792 ; n21793
g21538 and n21385_not n21388_not ; n21794
g21539 and n21793_not n21794_not ; n21795
g21540 and n21537 n21795_not ; n21796
g21541 and n21535_not n21796 ; n21797
g21542 and n21791_not n21797_not ; n21798
g21543 and b[26]_not n21798_not ; n21799
g21544 and n21060_not quotient[9]_not ; n21800
g21545 and n21070_not n21383 ; n21801
g21546 and n21379_not n21801 ; n21802
g21547 and n21380_not n21383_not ; n21803
g21548 and n21802_not n21803_not ; n21804
g21549 and n21537 n21804_not ; n21805
g21550 and n21535_not n21805 ; n21806
g21551 and n21800_not n21806_not ; n21807
g21552 and b[25]_not n21807_not ; n21808
g21553 and n21069_not quotient[9]_not ; n21809
g21554 and n21079_not n21378 ; n21810
g21555 and n21374_not n21810 ; n21811
g21556 and n21375_not n21378_not ; n21812
g21557 and n21811_not n21812_not ; n21813
g21558 and n21537 n21813_not ; n21814
g21559 and n21535_not n21814 ; n21815
g21560 and n21809_not n21815_not ; n21816
g21561 and b[24]_not n21816_not ; n21817
g21562 and n21078_not quotient[9]_not ; n21818
g21563 and n21088_not n21373 ; n21819
g21564 and n21369_not n21819 ; n21820
g21565 and n21370_not n21373_not ; n21821
g21566 and n21820_not n21821_not ; n21822
g21567 and n21537 n21822_not ; n21823
g21568 and n21535_not n21823 ; n21824
g21569 and n21818_not n21824_not ; n21825
g21570 and b[23]_not n21825_not ; n21826
g21571 and n21087_not quotient[9]_not ; n21827
g21572 and n21097_not n21368 ; n21828
g21573 and n21364_not n21828 ; n21829
g21574 and n21365_not n21368_not ; n21830
g21575 and n21829_not n21830_not ; n21831
g21576 and n21537 n21831_not ; n21832
g21577 and n21535_not n21832 ; n21833
g21578 and n21827_not n21833_not ; n21834
g21579 and b[22]_not n21834_not ; n21835
g21580 and n21096_not quotient[9]_not ; n21836
g21581 and n21106_not n21363 ; n21837
g21582 and n21359_not n21837 ; n21838
g21583 and n21360_not n21363_not ; n21839
g21584 and n21838_not n21839_not ; n21840
g21585 and n21537 n21840_not ; n21841
g21586 and n21535_not n21841 ; n21842
g21587 and n21836_not n21842_not ; n21843
g21588 and b[21]_not n21843_not ; n21844
g21589 and n21105_not quotient[9]_not ; n21845
g21590 and n21115_not n21358 ; n21846
g21591 and n21354_not n21846 ; n21847
g21592 and n21355_not n21358_not ; n21848
g21593 and n21847_not n21848_not ; n21849
g21594 and n21537 n21849_not ; n21850
g21595 and n21535_not n21850 ; n21851
g21596 and n21845_not n21851_not ; n21852
g21597 and b[20]_not n21852_not ; n21853
g21598 and n21114_not quotient[9]_not ; n21854
g21599 and n21124_not n21353 ; n21855
g21600 and n21349_not n21855 ; n21856
g21601 and n21350_not n21353_not ; n21857
g21602 and n21856_not n21857_not ; n21858
g21603 and n21537 n21858_not ; n21859
g21604 and n21535_not n21859 ; n21860
g21605 and n21854_not n21860_not ; n21861
g21606 and b[19]_not n21861_not ; n21862
g21607 and n21123_not quotient[9]_not ; n21863
g21608 and n21133_not n21348 ; n21864
g21609 and n21344_not n21864 ; n21865
g21610 and n21345_not n21348_not ; n21866
g21611 and n21865_not n21866_not ; n21867
g21612 and n21537 n21867_not ; n21868
g21613 and n21535_not n21868 ; n21869
g21614 and n21863_not n21869_not ; n21870
g21615 and b[18]_not n21870_not ; n21871
g21616 and n21132_not quotient[9]_not ; n21872
g21617 and n21142_not n21343 ; n21873
g21618 and n21339_not n21873 ; n21874
g21619 and n21340_not n21343_not ; n21875
g21620 and n21874_not n21875_not ; n21876
g21621 and n21537 n21876_not ; n21877
g21622 and n21535_not n21877 ; n21878
g21623 and n21872_not n21878_not ; n21879
g21624 and b[17]_not n21879_not ; n21880
g21625 and n21141_not quotient[9]_not ; n21881
g21626 and n21151_not n21338 ; n21882
g21627 and n21334_not n21882 ; n21883
g21628 and n21335_not n21338_not ; n21884
g21629 and n21883_not n21884_not ; n21885
g21630 and n21537 n21885_not ; n21886
g21631 and n21535_not n21886 ; n21887
g21632 and n21881_not n21887_not ; n21888
g21633 and b[16]_not n21888_not ; n21889
g21634 and n21150_not quotient[9]_not ; n21890
g21635 and n21160_not n21333 ; n21891
g21636 and n21329_not n21891 ; n21892
g21637 and n21330_not n21333_not ; n21893
g21638 and n21892_not n21893_not ; n21894
g21639 and n21537 n21894_not ; n21895
g21640 and n21535_not n21895 ; n21896
g21641 and n21890_not n21896_not ; n21897
g21642 and b[15]_not n21897_not ; n21898
g21643 and n21159_not quotient[9]_not ; n21899
g21644 and n21169_not n21328 ; n21900
g21645 and n21324_not n21900 ; n21901
g21646 and n21325_not n21328_not ; n21902
g21647 and n21901_not n21902_not ; n21903
g21648 and n21537 n21903_not ; n21904
g21649 and n21535_not n21904 ; n21905
g21650 and n21899_not n21905_not ; n21906
g21651 and b[14]_not n21906_not ; n21907
g21652 and n21168_not quotient[9]_not ; n21908
g21653 and n21178_not n21323 ; n21909
g21654 and n21319_not n21909 ; n21910
g21655 and n21320_not n21323_not ; n21911
g21656 and n21910_not n21911_not ; n21912
g21657 and n21537 n21912_not ; n21913
g21658 and n21535_not n21913 ; n21914
g21659 and n21908_not n21914_not ; n21915
g21660 and b[13]_not n21915_not ; n21916
g21661 and n21177_not quotient[9]_not ; n21917
g21662 and n21187_not n21318 ; n21918
g21663 and n21314_not n21918 ; n21919
g21664 and n21315_not n21318_not ; n21920
g21665 and n21919_not n21920_not ; n21921
g21666 and n21537 n21921_not ; n21922
g21667 and n21535_not n21922 ; n21923
g21668 and n21917_not n21923_not ; n21924
g21669 and b[12]_not n21924_not ; n21925
g21670 and n21186_not quotient[9]_not ; n21926
g21671 and n21196_not n21313 ; n21927
g21672 and n21309_not n21927 ; n21928
g21673 and n21310_not n21313_not ; n21929
g21674 and n21928_not n21929_not ; n21930
g21675 and n21537 n21930_not ; n21931
g21676 and n21535_not n21931 ; n21932
g21677 and n21926_not n21932_not ; n21933
g21678 and b[11]_not n21933_not ; n21934
g21679 and n21195_not quotient[9]_not ; n21935
g21680 and n21205_not n21308 ; n21936
g21681 and n21304_not n21936 ; n21937
g21682 and n21305_not n21308_not ; n21938
g21683 and n21937_not n21938_not ; n21939
g21684 and n21537 n21939_not ; n21940
g21685 and n21535_not n21940 ; n21941
g21686 and n21935_not n21941_not ; n21942
g21687 and b[10]_not n21942_not ; n21943
g21688 and n21204_not quotient[9]_not ; n21944
g21689 and n21214_not n21303 ; n21945
g21690 and n21299_not n21945 ; n21946
g21691 and n21300_not n21303_not ; n21947
g21692 and n21946_not n21947_not ; n21948
g21693 and n21537 n21948_not ; n21949
g21694 and n21535_not n21949 ; n21950
g21695 and n21944_not n21950_not ; n21951
g21696 and b[9]_not n21951_not ; n21952
g21697 and n21213_not quotient[9]_not ; n21953
g21698 and n21223_not n21298 ; n21954
g21699 and n21294_not n21954 ; n21955
g21700 and n21295_not n21298_not ; n21956
g21701 and n21955_not n21956_not ; n21957
g21702 and n21537 n21957_not ; n21958
g21703 and n21535_not n21958 ; n21959
g21704 and n21953_not n21959_not ; n21960
g21705 and b[8]_not n21960_not ; n21961
g21706 and n21222_not quotient[9]_not ; n21962
g21707 and n21232_not n21293 ; n21963
g21708 and n21289_not n21963 ; n21964
g21709 and n21290_not n21293_not ; n21965
g21710 and n21964_not n21965_not ; n21966
g21711 and n21537 n21966_not ; n21967
g21712 and n21535_not n21967 ; n21968
g21713 and n21962_not n21968_not ; n21969
g21714 and b[7]_not n21969_not ; n21970
g21715 and n21231_not quotient[9]_not ; n21971
g21716 and n21241_not n21288 ; n21972
g21717 and n21284_not n21972 ; n21973
g21718 and n21285_not n21288_not ; n21974
g21719 and n21973_not n21974_not ; n21975
g21720 and n21537 n21975_not ; n21976
g21721 and n21535_not n21976 ; n21977
g21722 and n21971_not n21977_not ; n21978
g21723 and b[6]_not n21978_not ; n21979
g21724 and n21240_not quotient[9]_not ; n21980
g21725 and n21250_not n21283 ; n21981
g21726 and n21279_not n21981 ; n21982
g21727 and n21280_not n21283_not ; n21983
g21728 and n21982_not n21983_not ; n21984
g21729 and n21537 n21984_not ; n21985
g21730 and n21535_not n21985 ; n21986
g21731 and n21980_not n21986_not ; n21987
g21732 and b[5]_not n21987_not ; n21988
g21733 and n21249_not quotient[9]_not ; n21989
g21734 and n21258_not n21278 ; n21990
g21735 and n21274_not n21990 ; n21991
g21736 and n21275_not n21278_not ; n21992
g21737 and n21991_not n21992_not ; n21993
g21738 and n21537 n21993_not ; n21994
g21739 and n21535_not n21994 ; n21995
g21740 and n21989_not n21995_not ; n21996
g21741 and b[4]_not n21996_not ; n21997
g21742 and n21257_not quotient[9]_not ; n21998
g21743 and n21269_not n21273 ; n21999
g21744 and n21268_not n21999 ; n22000
g21745 and n21270_not n21273_not ; n22001
g21746 and n22000_not n22001_not ; n22002
g21747 and n21537 n22002_not ; n22003
g21748 and n21535_not n22003 ; n22004
g21749 and n21998_not n22004_not ; n22005
g21750 and b[3]_not n22005_not ; n22006
g21751 and n21262_not quotient[9]_not ; n22007
g21752 and n21265_not n21267 ; n22008
g21753 and n21263_not n22008 ; n22009
g21754 and n21537 n22009_not ; n22010
g21755 and n21268_not n22010 ; n22011
g21756 and n21535_not n22011 ; n22012
g21757 and n22007_not n22012_not ; n22013
g21758 and b[2]_not n22013_not ; n22014
g21759 and b[0] b[55]_not ; n22015
g21760 and n283 n22015 ; n22016
g21761 and n280 n22016 ; n22017
g21762 and n21535_not n22017 ; n22018
g21763 and a[9] n22018_not ; n22019
g21764 and n396 n21267 ; n22020
g21765 and n406 n22020 ; n22021
g21766 and n403 n22021 ; n22022
g21767 and n21535_not n22022 ; n22023
g21768 and n22019_not n22023_not ; n22024
g21769 and b[1] n22024_not ; n22025
g21770 and b[1]_not n22023_not ; n22026
g21771 and n22019_not n22026 ; n22027
g21772 and n22025_not n22027_not ; n22028
g21773 and a[8]_not b[0] ; n22029
g21774 and n22028_not n22029_not ; n22030
g21775 and b[1]_not n22024_not ; n22031
g21776 and n22030_not n22031_not ; n22032
g21777 and b[2] n22012_not ; n22033
g21778 and n22007_not n22033 ; n22034
g21779 and n22014_not n22034_not ; n22035
g21780 and n22032_not n22035 ; n22036
g21781 and n22014_not n22036_not ; n22037
g21782 and b[3] n22004_not ; n22038
g21783 and n21998_not n22038 ; n22039
g21784 and n22006_not n22039_not ; n22040
g21785 and n22037_not n22040 ; n22041
g21786 and n22006_not n22041_not ; n22042
g21787 and b[4] n21995_not ; n22043
g21788 and n21989_not n22043 ; n22044
g21789 and n21997_not n22044_not ; n22045
g21790 and n22042_not n22045 ; n22046
g21791 and n21997_not n22046_not ; n22047
g21792 and b[5] n21986_not ; n22048
g21793 and n21980_not n22048 ; n22049
g21794 and n21988_not n22049_not ; n22050
g21795 and n22047_not n22050 ; n22051
g21796 and n21988_not n22051_not ; n22052
g21797 and b[6] n21977_not ; n22053
g21798 and n21971_not n22053 ; n22054
g21799 and n21979_not n22054_not ; n22055
g21800 and n22052_not n22055 ; n22056
g21801 and n21979_not n22056_not ; n22057
g21802 and b[7] n21968_not ; n22058
g21803 and n21962_not n22058 ; n22059
g21804 and n21970_not n22059_not ; n22060
g21805 and n22057_not n22060 ; n22061
g21806 and n21970_not n22061_not ; n22062
g21807 and b[8] n21959_not ; n22063
g21808 and n21953_not n22063 ; n22064
g21809 and n21961_not n22064_not ; n22065
g21810 and n22062_not n22065 ; n22066
g21811 and n21961_not n22066_not ; n22067
g21812 and b[9] n21950_not ; n22068
g21813 and n21944_not n22068 ; n22069
g21814 and n21952_not n22069_not ; n22070
g21815 and n22067_not n22070 ; n22071
g21816 and n21952_not n22071_not ; n22072
g21817 and b[10] n21941_not ; n22073
g21818 and n21935_not n22073 ; n22074
g21819 and n21943_not n22074_not ; n22075
g21820 and n22072_not n22075 ; n22076
g21821 and n21943_not n22076_not ; n22077
g21822 and b[11] n21932_not ; n22078
g21823 and n21926_not n22078 ; n22079
g21824 and n21934_not n22079_not ; n22080
g21825 and n22077_not n22080 ; n22081
g21826 and n21934_not n22081_not ; n22082
g21827 and b[12] n21923_not ; n22083
g21828 and n21917_not n22083 ; n22084
g21829 and n21925_not n22084_not ; n22085
g21830 and n22082_not n22085 ; n22086
g21831 and n21925_not n22086_not ; n22087
g21832 and b[13] n21914_not ; n22088
g21833 and n21908_not n22088 ; n22089
g21834 and n21916_not n22089_not ; n22090
g21835 and n22087_not n22090 ; n22091
g21836 and n21916_not n22091_not ; n22092
g21837 and b[14] n21905_not ; n22093
g21838 and n21899_not n22093 ; n22094
g21839 and n21907_not n22094_not ; n22095
g21840 and n22092_not n22095 ; n22096
g21841 and n21907_not n22096_not ; n22097
g21842 and b[15] n21896_not ; n22098
g21843 and n21890_not n22098 ; n22099
g21844 and n21898_not n22099_not ; n22100
g21845 and n22097_not n22100 ; n22101
g21846 and n21898_not n22101_not ; n22102
g21847 and b[16] n21887_not ; n22103
g21848 and n21881_not n22103 ; n22104
g21849 and n21889_not n22104_not ; n22105
g21850 and n22102_not n22105 ; n22106
g21851 and n21889_not n22106_not ; n22107
g21852 and b[17] n21878_not ; n22108
g21853 and n21872_not n22108 ; n22109
g21854 and n21880_not n22109_not ; n22110
g21855 and n22107_not n22110 ; n22111
g21856 and n21880_not n22111_not ; n22112
g21857 and b[18] n21869_not ; n22113
g21858 and n21863_not n22113 ; n22114
g21859 and n21871_not n22114_not ; n22115
g21860 and n22112_not n22115 ; n22116
g21861 and n21871_not n22116_not ; n22117
g21862 and b[19] n21860_not ; n22118
g21863 and n21854_not n22118 ; n22119
g21864 and n21862_not n22119_not ; n22120
g21865 and n22117_not n22120 ; n22121
g21866 and n21862_not n22121_not ; n22122
g21867 and b[20] n21851_not ; n22123
g21868 and n21845_not n22123 ; n22124
g21869 and n21853_not n22124_not ; n22125
g21870 and n22122_not n22125 ; n22126
g21871 and n21853_not n22126_not ; n22127
g21872 and b[21] n21842_not ; n22128
g21873 and n21836_not n22128 ; n22129
g21874 and n21844_not n22129_not ; n22130
g21875 and n22127_not n22130 ; n22131
g21876 and n21844_not n22131_not ; n22132
g21877 and b[22] n21833_not ; n22133
g21878 and n21827_not n22133 ; n22134
g21879 and n21835_not n22134_not ; n22135
g21880 and n22132_not n22135 ; n22136
g21881 and n21835_not n22136_not ; n22137
g21882 and b[23] n21824_not ; n22138
g21883 and n21818_not n22138 ; n22139
g21884 and n21826_not n22139_not ; n22140
g21885 and n22137_not n22140 ; n22141
g21886 and n21826_not n22141_not ; n22142
g21887 and b[24] n21815_not ; n22143
g21888 and n21809_not n22143 ; n22144
g21889 and n21817_not n22144_not ; n22145
g21890 and n22142_not n22145 ; n22146
g21891 and n21817_not n22146_not ; n22147
g21892 and b[25] n21806_not ; n22148
g21893 and n21800_not n22148 ; n22149
g21894 and n21808_not n22149_not ; n22150
g21895 and n22147_not n22150 ; n22151
g21896 and n21808_not n22151_not ; n22152
g21897 and b[26] n21797_not ; n22153
g21898 and n21791_not n22153 ; n22154
g21899 and n21799_not n22154_not ; n22155
g21900 and n22152_not n22155 ; n22156
g21901 and n21799_not n22156_not ; n22157
g21902 and b[27] n21788_not ; n22158
g21903 and n21782_not n22158 ; n22159
g21904 and n21790_not n22159_not ; n22160
g21905 and n22157_not n22160 ; n22161
g21906 and n21790_not n22161_not ; n22162
g21907 and b[28] n21779_not ; n22163
g21908 and n21773_not n22163 ; n22164
g21909 and n21781_not n22164_not ; n22165
g21910 and n22162_not n22165 ; n22166
g21911 and n21781_not n22166_not ; n22167
g21912 and b[29] n21770_not ; n22168
g21913 and n21764_not n22168 ; n22169
g21914 and n21772_not n22169_not ; n22170
g21915 and n22167_not n22170 ; n22171
g21916 and n21772_not n22171_not ; n22172
g21917 and b[30] n21761_not ; n22173
g21918 and n21755_not n22173 ; n22174
g21919 and n21763_not n22174_not ; n22175
g21920 and n22172_not n22175 ; n22176
g21921 and n21763_not n22176_not ; n22177
g21922 and b[31] n21752_not ; n22178
g21923 and n21746_not n22178 ; n22179
g21924 and n21754_not n22179_not ; n22180
g21925 and n22177_not n22180 ; n22181
g21926 and n21754_not n22181_not ; n22182
g21927 and b[32] n21743_not ; n22183
g21928 and n21737_not n22183 ; n22184
g21929 and n21745_not n22184_not ; n22185
g21930 and n22182_not n22185 ; n22186
g21931 and n21745_not n22186_not ; n22187
g21932 and b[33] n21734_not ; n22188
g21933 and n21728_not n22188 ; n22189
g21934 and n21736_not n22189_not ; n22190
g21935 and n22187_not n22190 ; n22191
g21936 and n21736_not n22191_not ; n22192
g21937 and b[34] n21725_not ; n22193
g21938 and n21719_not n22193 ; n22194
g21939 and n21727_not n22194_not ; n22195
g21940 and n22192_not n22195 ; n22196
g21941 and n21727_not n22196_not ; n22197
g21942 and b[35] n21716_not ; n22198
g21943 and n21710_not n22198 ; n22199
g21944 and n21718_not n22199_not ; n22200
g21945 and n22197_not n22200 ; n22201
g21946 and n21718_not n22201_not ; n22202
g21947 and b[36] n21707_not ; n22203
g21948 and n21701_not n22203 ; n22204
g21949 and n21709_not n22204_not ; n22205
g21950 and n22202_not n22205 ; n22206
g21951 and n21709_not n22206_not ; n22207
g21952 and b[37] n21698_not ; n22208
g21953 and n21692_not n22208 ; n22209
g21954 and n21700_not n22209_not ; n22210
g21955 and n22207_not n22210 ; n22211
g21956 and n21700_not n22211_not ; n22212
g21957 and b[38] n21689_not ; n22213
g21958 and n21683_not n22213 ; n22214
g21959 and n21691_not n22214_not ; n22215
g21960 and n22212_not n22215 ; n22216
g21961 and n21691_not n22216_not ; n22217
g21962 and b[39] n21680_not ; n22218
g21963 and n21674_not n22218 ; n22219
g21964 and n21682_not n22219_not ; n22220
g21965 and n22217_not n22220 ; n22221
g21966 and n21682_not n22221_not ; n22222
g21967 and b[40] n21671_not ; n22223
g21968 and n21665_not n22223 ; n22224
g21969 and n21673_not n22224_not ; n22225
g21970 and n22222_not n22225 ; n22226
g21971 and n21673_not n22226_not ; n22227
g21972 and b[41] n21662_not ; n22228
g21973 and n21656_not n22228 ; n22229
g21974 and n21664_not n22229_not ; n22230
g21975 and n22227_not n22230 ; n22231
g21976 and n21664_not n22231_not ; n22232
g21977 and b[42] n21653_not ; n22233
g21978 and n21647_not n22233 ; n22234
g21979 and n21655_not n22234_not ; n22235
g21980 and n22232_not n22235 ; n22236
g21981 and n21655_not n22236_not ; n22237
g21982 and b[43] n21644_not ; n22238
g21983 and n21638_not n22238 ; n22239
g21984 and n21646_not n22239_not ; n22240
g21985 and n22237_not n22240 ; n22241
g21986 and n21646_not n22241_not ; n22242
g21987 and b[44] n21635_not ; n22243
g21988 and n21629_not n22243 ; n22244
g21989 and n21637_not n22244_not ; n22245
g21990 and n22242_not n22245 ; n22246
g21991 and n21637_not n22246_not ; n22247
g21992 and b[45] n21626_not ; n22248
g21993 and n21620_not n22248 ; n22249
g21994 and n21628_not n22249_not ; n22250
g21995 and n22247_not n22250 ; n22251
g21996 and n21628_not n22251_not ; n22252
g21997 and b[46] n21617_not ; n22253
g21998 and n21611_not n22253 ; n22254
g21999 and n21619_not n22254_not ; n22255
g22000 and n22252_not n22255 ; n22256
g22001 and n21619_not n22256_not ; n22257
g22002 and b[47] n21608_not ; n22258
g22003 and n21602_not n22258 ; n22259
g22004 and n21610_not n22259_not ; n22260
g22005 and n22257_not n22260 ; n22261
g22006 and n21610_not n22261_not ; n22262
g22007 and b[48] n21599_not ; n22263
g22008 and n21593_not n22263 ; n22264
g22009 and n21601_not n22264_not ; n22265
g22010 and n22262_not n22265 ; n22266
g22011 and n21601_not n22266_not ; n22267
g22012 and b[49] n21590_not ; n22268
g22013 and n21584_not n22268 ; n22269
g22014 and n21592_not n22269_not ; n22270
g22015 and n22267_not n22270 ; n22271
g22016 and n21592_not n22271_not ; n22272
g22017 and b[50] n21581_not ; n22273
g22018 and n21575_not n22273 ; n22274
g22019 and n21583_not n22274_not ; n22275
g22020 and n22272_not n22275 ; n22276
g22021 and n21583_not n22276_not ; n22277
g22022 and b[51] n21572_not ; n22278
g22023 and n21566_not n22278 ; n22279
g22024 and n21574_not n22279_not ; n22280
g22025 and n22277_not n22280 ; n22281
g22026 and n21574_not n22281_not ; n22282
g22027 and b[52] n21563_not ; n22283
g22028 and n21557_not n22283 ; n22284
g22029 and n21565_not n22284_not ; n22285
g22030 and n22282_not n22285 ; n22286
g22031 and n21565_not n22286_not ; n22287
g22032 and b[53] n21554_not ; n22288
g22033 and n21548_not n22288 ; n22289
g22034 and n21556_not n22289_not ; n22290
g22035 and n22287_not n22290 ; n22291
g22036 and n21556_not n22291_not ; n22292
g22037 and b[54] n21545_not ; n22293
g22038 and n21539_not n22293 ; n22294
g22039 and n21547_not n22294_not ; n22295
g22040 and n22292_not n22295 ; n22296
g22041 and n21547_not n22296_not ; n22297
g22042 and n20798_not quotient[9]_not ; n22298
g22043 and n20800_not n21533 ; n22299
g22044 and n21529_not n22299 ; n22300
g22045 and n21530_not n21533_not ; n22301
g22046 and n22300_not n22301_not ; n22302
g22047 and quotient[9] n22302_not ; n22303
g22048 and n22298_not n22303_not ; n22304
g22049 and b[55]_not n22304_not ; n22305
g22050 and b[55] n22298_not ; n22306
g22051 and n22303_not n22306 ; n22307
g22052 and n337 n22307_not ; n22308
g22053 and n22305_not n22308 ; n22309
g22054 and n22297_not n22309 ; n22310
g22055 and n21537 n22304_not ; n22311
g22056 and n22310_not n22311_not ; quotient[8]
g22057 and n21556_not n22295 ; n22313
g22058 and n22291_not n22313 ; n22314
g22059 and n22292_not n22295_not ; n22315
g22060 and n22314_not n22315_not ; n22316
g22061 and quotient[8] n22316_not ; n22317
g22062 and n21546_not n22311_not ; n22318
g22063 and n22310_not n22318 ; n22319
g22064 and n22317_not n22319_not ; n22320
g22065 and b[55]_not n22320_not ; n22321
g22066 and n21565_not n22290 ; n22322
g22067 and n22286_not n22322 ; n22323
g22068 and n22287_not n22290_not ; n22324
g22069 and n22323_not n22324_not ; n22325
g22070 and quotient[8] n22325_not ; n22326
g22071 and n21555_not n22311_not ; n22327
g22072 and n22310_not n22327 ; n22328
g22073 and n22326_not n22328_not ; n22329
g22074 and b[54]_not n22329_not ; n22330
g22075 and n21574_not n22285 ; n22331
g22076 and n22281_not n22331 ; n22332
g22077 and n22282_not n22285_not ; n22333
g22078 and n22332_not n22333_not ; n22334
g22079 and quotient[8] n22334_not ; n22335
g22080 and n21564_not n22311_not ; n22336
g22081 and n22310_not n22336 ; n22337
g22082 and n22335_not n22337_not ; n22338
g22083 and b[53]_not n22338_not ; n22339
g22084 and n21583_not n22280 ; n22340
g22085 and n22276_not n22340 ; n22341
g22086 and n22277_not n22280_not ; n22342
g22087 and n22341_not n22342_not ; n22343
g22088 and quotient[8] n22343_not ; n22344
g22089 and n21573_not n22311_not ; n22345
g22090 and n22310_not n22345 ; n22346
g22091 and n22344_not n22346_not ; n22347
g22092 and b[52]_not n22347_not ; n22348
g22093 and n21592_not n22275 ; n22349
g22094 and n22271_not n22349 ; n22350
g22095 and n22272_not n22275_not ; n22351
g22096 and n22350_not n22351_not ; n22352
g22097 and quotient[8] n22352_not ; n22353
g22098 and n21582_not n22311_not ; n22354
g22099 and n22310_not n22354 ; n22355
g22100 and n22353_not n22355_not ; n22356
g22101 and b[51]_not n22356_not ; n22357
g22102 and n21601_not n22270 ; n22358
g22103 and n22266_not n22358 ; n22359
g22104 and n22267_not n22270_not ; n22360
g22105 and n22359_not n22360_not ; n22361
g22106 and quotient[8] n22361_not ; n22362
g22107 and n21591_not n22311_not ; n22363
g22108 and n22310_not n22363 ; n22364
g22109 and n22362_not n22364_not ; n22365
g22110 and b[50]_not n22365_not ; n22366
g22111 and n21610_not n22265 ; n22367
g22112 and n22261_not n22367 ; n22368
g22113 and n22262_not n22265_not ; n22369
g22114 and n22368_not n22369_not ; n22370
g22115 and quotient[8] n22370_not ; n22371
g22116 and n21600_not n22311_not ; n22372
g22117 and n22310_not n22372 ; n22373
g22118 and n22371_not n22373_not ; n22374
g22119 and b[49]_not n22374_not ; n22375
g22120 and n21619_not n22260 ; n22376
g22121 and n22256_not n22376 ; n22377
g22122 and n22257_not n22260_not ; n22378
g22123 and n22377_not n22378_not ; n22379
g22124 and quotient[8] n22379_not ; n22380
g22125 and n21609_not n22311_not ; n22381
g22126 and n22310_not n22381 ; n22382
g22127 and n22380_not n22382_not ; n22383
g22128 and b[48]_not n22383_not ; n22384
g22129 and n21628_not n22255 ; n22385
g22130 and n22251_not n22385 ; n22386
g22131 and n22252_not n22255_not ; n22387
g22132 and n22386_not n22387_not ; n22388
g22133 and quotient[8] n22388_not ; n22389
g22134 and n21618_not n22311_not ; n22390
g22135 and n22310_not n22390 ; n22391
g22136 and n22389_not n22391_not ; n22392
g22137 and b[47]_not n22392_not ; n22393
g22138 and n21637_not n22250 ; n22394
g22139 and n22246_not n22394 ; n22395
g22140 and n22247_not n22250_not ; n22396
g22141 and n22395_not n22396_not ; n22397
g22142 and quotient[8] n22397_not ; n22398
g22143 and n21627_not n22311_not ; n22399
g22144 and n22310_not n22399 ; n22400
g22145 and n22398_not n22400_not ; n22401
g22146 and b[46]_not n22401_not ; n22402
g22147 and n21646_not n22245 ; n22403
g22148 and n22241_not n22403 ; n22404
g22149 and n22242_not n22245_not ; n22405
g22150 and n22404_not n22405_not ; n22406
g22151 and quotient[8] n22406_not ; n22407
g22152 and n21636_not n22311_not ; n22408
g22153 and n22310_not n22408 ; n22409
g22154 and n22407_not n22409_not ; n22410
g22155 and b[45]_not n22410_not ; n22411
g22156 and n21655_not n22240 ; n22412
g22157 and n22236_not n22412 ; n22413
g22158 and n22237_not n22240_not ; n22414
g22159 and n22413_not n22414_not ; n22415
g22160 and quotient[8] n22415_not ; n22416
g22161 and n21645_not n22311_not ; n22417
g22162 and n22310_not n22417 ; n22418
g22163 and n22416_not n22418_not ; n22419
g22164 and b[44]_not n22419_not ; n22420
g22165 and n21664_not n22235 ; n22421
g22166 and n22231_not n22421 ; n22422
g22167 and n22232_not n22235_not ; n22423
g22168 and n22422_not n22423_not ; n22424
g22169 and quotient[8] n22424_not ; n22425
g22170 and n21654_not n22311_not ; n22426
g22171 and n22310_not n22426 ; n22427
g22172 and n22425_not n22427_not ; n22428
g22173 and b[43]_not n22428_not ; n22429
g22174 and n21673_not n22230 ; n22430
g22175 and n22226_not n22430 ; n22431
g22176 and n22227_not n22230_not ; n22432
g22177 and n22431_not n22432_not ; n22433
g22178 and quotient[8] n22433_not ; n22434
g22179 and n21663_not n22311_not ; n22435
g22180 and n22310_not n22435 ; n22436
g22181 and n22434_not n22436_not ; n22437
g22182 and b[42]_not n22437_not ; n22438
g22183 and n21682_not n22225 ; n22439
g22184 and n22221_not n22439 ; n22440
g22185 and n22222_not n22225_not ; n22441
g22186 and n22440_not n22441_not ; n22442
g22187 and quotient[8] n22442_not ; n22443
g22188 and n21672_not n22311_not ; n22444
g22189 and n22310_not n22444 ; n22445
g22190 and n22443_not n22445_not ; n22446
g22191 and b[41]_not n22446_not ; n22447
g22192 and n21691_not n22220 ; n22448
g22193 and n22216_not n22448 ; n22449
g22194 and n22217_not n22220_not ; n22450
g22195 and n22449_not n22450_not ; n22451
g22196 and quotient[8] n22451_not ; n22452
g22197 and n21681_not n22311_not ; n22453
g22198 and n22310_not n22453 ; n22454
g22199 and n22452_not n22454_not ; n22455
g22200 and b[40]_not n22455_not ; n22456
g22201 and n21700_not n22215 ; n22457
g22202 and n22211_not n22457 ; n22458
g22203 and n22212_not n22215_not ; n22459
g22204 and n22458_not n22459_not ; n22460
g22205 and quotient[8] n22460_not ; n22461
g22206 and n21690_not n22311_not ; n22462
g22207 and n22310_not n22462 ; n22463
g22208 and n22461_not n22463_not ; n22464
g22209 and b[39]_not n22464_not ; n22465
g22210 and n21709_not n22210 ; n22466
g22211 and n22206_not n22466 ; n22467
g22212 and n22207_not n22210_not ; n22468
g22213 and n22467_not n22468_not ; n22469
g22214 and quotient[8] n22469_not ; n22470
g22215 and n21699_not n22311_not ; n22471
g22216 and n22310_not n22471 ; n22472
g22217 and n22470_not n22472_not ; n22473
g22218 and b[38]_not n22473_not ; n22474
g22219 and n21718_not n22205 ; n22475
g22220 and n22201_not n22475 ; n22476
g22221 and n22202_not n22205_not ; n22477
g22222 and n22476_not n22477_not ; n22478
g22223 and quotient[8] n22478_not ; n22479
g22224 and n21708_not n22311_not ; n22480
g22225 and n22310_not n22480 ; n22481
g22226 and n22479_not n22481_not ; n22482
g22227 and b[37]_not n22482_not ; n22483
g22228 and n21727_not n22200 ; n22484
g22229 and n22196_not n22484 ; n22485
g22230 and n22197_not n22200_not ; n22486
g22231 and n22485_not n22486_not ; n22487
g22232 and quotient[8] n22487_not ; n22488
g22233 and n21717_not n22311_not ; n22489
g22234 and n22310_not n22489 ; n22490
g22235 and n22488_not n22490_not ; n22491
g22236 and b[36]_not n22491_not ; n22492
g22237 and n21736_not n22195 ; n22493
g22238 and n22191_not n22493 ; n22494
g22239 and n22192_not n22195_not ; n22495
g22240 and n22494_not n22495_not ; n22496
g22241 and quotient[8] n22496_not ; n22497
g22242 and n21726_not n22311_not ; n22498
g22243 and n22310_not n22498 ; n22499
g22244 and n22497_not n22499_not ; n22500
g22245 and b[35]_not n22500_not ; n22501
g22246 and n21745_not n22190 ; n22502
g22247 and n22186_not n22502 ; n22503
g22248 and n22187_not n22190_not ; n22504
g22249 and n22503_not n22504_not ; n22505
g22250 and quotient[8] n22505_not ; n22506
g22251 and n21735_not n22311_not ; n22507
g22252 and n22310_not n22507 ; n22508
g22253 and n22506_not n22508_not ; n22509
g22254 and b[34]_not n22509_not ; n22510
g22255 and n21754_not n22185 ; n22511
g22256 and n22181_not n22511 ; n22512
g22257 and n22182_not n22185_not ; n22513
g22258 and n22512_not n22513_not ; n22514
g22259 and quotient[8] n22514_not ; n22515
g22260 and n21744_not n22311_not ; n22516
g22261 and n22310_not n22516 ; n22517
g22262 and n22515_not n22517_not ; n22518
g22263 and b[33]_not n22518_not ; n22519
g22264 and n21763_not n22180 ; n22520
g22265 and n22176_not n22520 ; n22521
g22266 and n22177_not n22180_not ; n22522
g22267 and n22521_not n22522_not ; n22523
g22268 and quotient[8] n22523_not ; n22524
g22269 and n21753_not n22311_not ; n22525
g22270 and n22310_not n22525 ; n22526
g22271 and n22524_not n22526_not ; n22527
g22272 and b[32]_not n22527_not ; n22528
g22273 and n21772_not n22175 ; n22529
g22274 and n22171_not n22529 ; n22530
g22275 and n22172_not n22175_not ; n22531
g22276 and n22530_not n22531_not ; n22532
g22277 and quotient[8] n22532_not ; n22533
g22278 and n21762_not n22311_not ; n22534
g22279 and n22310_not n22534 ; n22535
g22280 and n22533_not n22535_not ; n22536
g22281 and b[31]_not n22536_not ; n22537
g22282 and n21781_not n22170 ; n22538
g22283 and n22166_not n22538 ; n22539
g22284 and n22167_not n22170_not ; n22540
g22285 and n22539_not n22540_not ; n22541
g22286 and quotient[8] n22541_not ; n22542
g22287 and n21771_not n22311_not ; n22543
g22288 and n22310_not n22543 ; n22544
g22289 and n22542_not n22544_not ; n22545
g22290 and b[30]_not n22545_not ; n22546
g22291 and n21790_not n22165 ; n22547
g22292 and n22161_not n22547 ; n22548
g22293 and n22162_not n22165_not ; n22549
g22294 and n22548_not n22549_not ; n22550
g22295 and quotient[8] n22550_not ; n22551
g22296 and n21780_not n22311_not ; n22552
g22297 and n22310_not n22552 ; n22553
g22298 and n22551_not n22553_not ; n22554
g22299 and b[29]_not n22554_not ; n22555
g22300 and n21799_not n22160 ; n22556
g22301 and n22156_not n22556 ; n22557
g22302 and n22157_not n22160_not ; n22558
g22303 and n22557_not n22558_not ; n22559
g22304 and quotient[8] n22559_not ; n22560
g22305 and n21789_not n22311_not ; n22561
g22306 and n22310_not n22561 ; n22562
g22307 and n22560_not n22562_not ; n22563
g22308 and b[28]_not n22563_not ; n22564
g22309 and n21808_not n22155 ; n22565
g22310 and n22151_not n22565 ; n22566
g22311 and n22152_not n22155_not ; n22567
g22312 and n22566_not n22567_not ; n22568
g22313 and quotient[8] n22568_not ; n22569
g22314 and n21798_not n22311_not ; n22570
g22315 and n22310_not n22570 ; n22571
g22316 and n22569_not n22571_not ; n22572
g22317 and b[27]_not n22572_not ; n22573
g22318 and n21817_not n22150 ; n22574
g22319 and n22146_not n22574 ; n22575
g22320 and n22147_not n22150_not ; n22576
g22321 and n22575_not n22576_not ; n22577
g22322 and quotient[8] n22577_not ; n22578
g22323 and n21807_not n22311_not ; n22579
g22324 and n22310_not n22579 ; n22580
g22325 and n22578_not n22580_not ; n22581
g22326 and b[26]_not n22581_not ; n22582
g22327 and n21826_not n22145 ; n22583
g22328 and n22141_not n22583 ; n22584
g22329 and n22142_not n22145_not ; n22585
g22330 and n22584_not n22585_not ; n22586
g22331 and quotient[8] n22586_not ; n22587
g22332 and n21816_not n22311_not ; n22588
g22333 and n22310_not n22588 ; n22589
g22334 and n22587_not n22589_not ; n22590
g22335 and b[25]_not n22590_not ; n22591
g22336 and n21835_not n22140 ; n22592
g22337 and n22136_not n22592 ; n22593
g22338 and n22137_not n22140_not ; n22594
g22339 and n22593_not n22594_not ; n22595
g22340 and quotient[8] n22595_not ; n22596
g22341 and n21825_not n22311_not ; n22597
g22342 and n22310_not n22597 ; n22598
g22343 and n22596_not n22598_not ; n22599
g22344 and b[24]_not n22599_not ; n22600
g22345 and n21844_not n22135 ; n22601
g22346 and n22131_not n22601 ; n22602
g22347 and n22132_not n22135_not ; n22603
g22348 and n22602_not n22603_not ; n22604
g22349 and quotient[8] n22604_not ; n22605
g22350 and n21834_not n22311_not ; n22606
g22351 and n22310_not n22606 ; n22607
g22352 and n22605_not n22607_not ; n22608
g22353 and b[23]_not n22608_not ; n22609
g22354 and n21853_not n22130 ; n22610
g22355 and n22126_not n22610 ; n22611
g22356 and n22127_not n22130_not ; n22612
g22357 and n22611_not n22612_not ; n22613
g22358 and quotient[8] n22613_not ; n22614
g22359 and n21843_not n22311_not ; n22615
g22360 and n22310_not n22615 ; n22616
g22361 and n22614_not n22616_not ; n22617
g22362 and b[22]_not n22617_not ; n22618
g22363 and n21862_not n22125 ; n22619
g22364 and n22121_not n22619 ; n22620
g22365 and n22122_not n22125_not ; n22621
g22366 and n22620_not n22621_not ; n22622
g22367 and quotient[8] n22622_not ; n22623
g22368 and n21852_not n22311_not ; n22624
g22369 and n22310_not n22624 ; n22625
g22370 and n22623_not n22625_not ; n22626
g22371 and b[21]_not n22626_not ; n22627
g22372 and n21871_not n22120 ; n22628
g22373 and n22116_not n22628 ; n22629
g22374 and n22117_not n22120_not ; n22630
g22375 and n22629_not n22630_not ; n22631
g22376 and quotient[8] n22631_not ; n22632
g22377 and n21861_not n22311_not ; n22633
g22378 and n22310_not n22633 ; n22634
g22379 and n22632_not n22634_not ; n22635
g22380 and b[20]_not n22635_not ; n22636
g22381 and n21880_not n22115 ; n22637
g22382 and n22111_not n22637 ; n22638
g22383 and n22112_not n22115_not ; n22639
g22384 and n22638_not n22639_not ; n22640
g22385 and quotient[8] n22640_not ; n22641
g22386 and n21870_not n22311_not ; n22642
g22387 and n22310_not n22642 ; n22643
g22388 and n22641_not n22643_not ; n22644
g22389 and b[19]_not n22644_not ; n22645
g22390 and n21889_not n22110 ; n22646
g22391 and n22106_not n22646 ; n22647
g22392 and n22107_not n22110_not ; n22648
g22393 and n22647_not n22648_not ; n22649
g22394 and quotient[8] n22649_not ; n22650
g22395 and n21879_not n22311_not ; n22651
g22396 and n22310_not n22651 ; n22652
g22397 and n22650_not n22652_not ; n22653
g22398 and b[18]_not n22653_not ; n22654
g22399 and n21898_not n22105 ; n22655
g22400 and n22101_not n22655 ; n22656
g22401 and n22102_not n22105_not ; n22657
g22402 and n22656_not n22657_not ; n22658
g22403 and quotient[8] n22658_not ; n22659
g22404 and n21888_not n22311_not ; n22660
g22405 and n22310_not n22660 ; n22661
g22406 and n22659_not n22661_not ; n22662
g22407 and b[17]_not n22662_not ; n22663
g22408 and n21907_not n22100 ; n22664
g22409 and n22096_not n22664 ; n22665
g22410 and n22097_not n22100_not ; n22666
g22411 and n22665_not n22666_not ; n22667
g22412 and quotient[8] n22667_not ; n22668
g22413 and n21897_not n22311_not ; n22669
g22414 and n22310_not n22669 ; n22670
g22415 and n22668_not n22670_not ; n22671
g22416 and b[16]_not n22671_not ; n22672
g22417 and n21916_not n22095 ; n22673
g22418 and n22091_not n22673 ; n22674
g22419 and n22092_not n22095_not ; n22675
g22420 and n22674_not n22675_not ; n22676
g22421 and quotient[8] n22676_not ; n22677
g22422 and n21906_not n22311_not ; n22678
g22423 and n22310_not n22678 ; n22679
g22424 and n22677_not n22679_not ; n22680
g22425 and b[15]_not n22680_not ; n22681
g22426 and n21925_not n22090 ; n22682
g22427 and n22086_not n22682 ; n22683
g22428 and n22087_not n22090_not ; n22684
g22429 and n22683_not n22684_not ; n22685
g22430 and quotient[8] n22685_not ; n22686
g22431 and n21915_not n22311_not ; n22687
g22432 and n22310_not n22687 ; n22688
g22433 and n22686_not n22688_not ; n22689
g22434 and b[14]_not n22689_not ; n22690
g22435 and n21934_not n22085 ; n22691
g22436 and n22081_not n22691 ; n22692
g22437 and n22082_not n22085_not ; n22693
g22438 and n22692_not n22693_not ; n22694
g22439 and quotient[8] n22694_not ; n22695
g22440 and n21924_not n22311_not ; n22696
g22441 and n22310_not n22696 ; n22697
g22442 and n22695_not n22697_not ; n22698
g22443 and b[13]_not n22698_not ; n22699
g22444 and n21943_not n22080 ; n22700
g22445 and n22076_not n22700 ; n22701
g22446 and n22077_not n22080_not ; n22702
g22447 and n22701_not n22702_not ; n22703
g22448 and quotient[8] n22703_not ; n22704
g22449 and n21933_not n22311_not ; n22705
g22450 and n22310_not n22705 ; n22706
g22451 and n22704_not n22706_not ; n22707
g22452 and b[12]_not n22707_not ; n22708
g22453 and n21952_not n22075 ; n22709
g22454 and n22071_not n22709 ; n22710
g22455 and n22072_not n22075_not ; n22711
g22456 and n22710_not n22711_not ; n22712
g22457 and quotient[8] n22712_not ; n22713
g22458 and n21942_not n22311_not ; n22714
g22459 and n22310_not n22714 ; n22715
g22460 and n22713_not n22715_not ; n22716
g22461 and b[11]_not n22716_not ; n22717
g22462 and n21961_not n22070 ; n22718
g22463 and n22066_not n22718 ; n22719
g22464 and n22067_not n22070_not ; n22720
g22465 and n22719_not n22720_not ; n22721
g22466 and quotient[8] n22721_not ; n22722
g22467 and n21951_not n22311_not ; n22723
g22468 and n22310_not n22723 ; n22724
g22469 and n22722_not n22724_not ; n22725
g22470 and b[10]_not n22725_not ; n22726
g22471 and n21970_not n22065 ; n22727
g22472 and n22061_not n22727 ; n22728
g22473 and n22062_not n22065_not ; n22729
g22474 and n22728_not n22729_not ; n22730
g22475 and quotient[8] n22730_not ; n22731
g22476 and n21960_not n22311_not ; n22732
g22477 and n22310_not n22732 ; n22733
g22478 and n22731_not n22733_not ; n22734
g22479 and b[9]_not n22734_not ; n22735
g22480 and n21979_not n22060 ; n22736
g22481 and n22056_not n22736 ; n22737
g22482 and n22057_not n22060_not ; n22738
g22483 and n22737_not n22738_not ; n22739
g22484 and quotient[8] n22739_not ; n22740
g22485 and n21969_not n22311_not ; n22741
g22486 and n22310_not n22741 ; n22742
g22487 and n22740_not n22742_not ; n22743
g22488 and b[8]_not n22743_not ; n22744
g22489 and n21988_not n22055 ; n22745
g22490 and n22051_not n22745 ; n22746
g22491 and n22052_not n22055_not ; n22747
g22492 and n22746_not n22747_not ; n22748
g22493 and quotient[8] n22748_not ; n22749
g22494 and n21978_not n22311_not ; n22750
g22495 and n22310_not n22750 ; n22751
g22496 and n22749_not n22751_not ; n22752
g22497 and b[7]_not n22752_not ; n22753
g22498 and n21997_not n22050 ; n22754
g22499 and n22046_not n22754 ; n22755
g22500 and n22047_not n22050_not ; n22756
g22501 and n22755_not n22756_not ; n22757
g22502 and quotient[8] n22757_not ; n22758
g22503 and n21987_not n22311_not ; n22759
g22504 and n22310_not n22759 ; n22760
g22505 and n22758_not n22760_not ; n22761
g22506 and b[6]_not n22761_not ; n22762
g22507 and n22006_not n22045 ; n22763
g22508 and n22041_not n22763 ; n22764
g22509 and n22042_not n22045_not ; n22765
g22510 and n22764_not n22765_not ; n22766
g22511 and quotient[8] n22766_not ; n22767
g22512 and n21996_not n22311_not ; n22768
g22513 and n22310_not n22768 ; n22769
g22514 and n22767_not n22769_not ; n22770
g22515 and b[5]_not n22770_not ; n22771
g22516 and n22014_not n22040 ; n22772
g22517 and n22036_not n22772 ; n22773
g22518 and n22037_not n22040_not ; n22774
g22519 and n22773_not n22774_not ; n22775
g22520 and quotient[8] n22775_not ; n22776
g22521 and n22005_not n22311_not ; n22777
g22522 and n22310_not n22777 ; n22778
g22523 and n22776_not n22778_not ; n22779
g22524 and b[4]_not n22779_not ; n22780
g22525 and n22031_not n22035 ; n22781
g22526 and n22030_not n22781 ; n22782
g22527 and n22032_not n22035_not ; n22783
g22528 and n22782_not n22783_not ; n22784
g22529 and quotient[8] n22784_not ; n22785
g22530 and n22013_not n22311_not ; n22786
g22531 and n22310_not n22786 ; n22787
g22532 and n22785_not n22787_not ; n22788
g22533 and b[3]_not n22788_not ; n22789
g22534 and n22027_not n22029 ; n22790
g22535 and n22025_not n22790 ; n22791
g22536 and n22030_not n22791_not ; n22792
g22537 and quotient[8] n22792 ; n22793
g22538 and n22024_not n22311_not ; n22794
g22539 and n22310_not n22794 ; n22795
g22540 and n22793_not n22795_not ; n22796
g22541 and b[2]_not n22796_not ; n22797
g22542 and b[0] quotient[8] ; n22798
g22543 and a[8] n22798_not ; n22799
g22544 and n22029 quotient[8] ; n22800
g22545 and n22799_not n22800_not ; n22801
g22546 and b[1] n22801_not ; n22802
g22547 and b[1]_not n22800_not ; n22803
g22548 and n22799_not n22803 ; n22804
g22549 and n22802_not n22804_not ; n22805
g22550 and a[7]_not b[0] ; n22806
g22551 and n22805_not n22806_not ; n22807
g22552 and b[1]_not n22801_not ; n22808
g22553 and n22807_not n22808_not ; n22809
g22554 and b[2] n22795_not ; n22810
g22555 and n22793_not n22810 ; n22811
g22556 and n22797_not n22811_not ; n22812
g22557 and n22809_not n22812 ; n22813
g22558 and n22797_not n22813_not ; n22814
g22559 and b[3] n22787_not ; n22815
g22560 and n22785_not n22815 ; n22816
g22561 and n22789_not n22816_not ; n22817
g22562 and n22814_not n22817 ; n22818
g22563 and n22789_not n22818_not ; n22819
g22564 and b[4] n22778_not ; n22820
g22565 and n22776_not n22820 ; n22821
g22566 and n22780_not n22821_not ; n22822
g22567 and n22819_not n22822 ; n22823
g22568 and n22780_not n22823_not ; n22824
g22569 and b[5] n22769_not ; n22825
g22570 and n22767_not n22825 ; n22826
g22571 and n22771_not n22826_not ; n22827
g22572 and n22824_not n22827 ; n22828
g22573 and n22771_not n22828_not ; n22829
g22574 and b[6] n22760_not ; n22830
g22575 and n22758_not n22830 ; n22831
g22576 and n22762_not n22831_not ; n22832
g22577 and n22829_not n22832 ; n22833
g22578 and n22762_not n22833_not ; n22834
g22579 and b[7] n22751_not ; n22835
g22580 and n22749_not n22835 ; n22836
g22581 and n22753_not n22836_not ; n22837
g22582 and n22834_not n22837 ; n22838
g22583 and n22753_not n22838_not ; n22839
g22584 and b[8] n22742_not ; n22840
g22585 and n22740_not n22840 ; n22841
g22586 and n22744_not n22841_not ; n22842
g22587 and n22839_not n22842 ; n22843
g22588 and n22744_not n22843_not ; n22844
g22589 and b[9] n22733_not ; n22845
g22590 and n22731_not n22845 ; n22846
g22591 and n22735_not n22846_not ; n22847
g22592 and n22844_not n22847 ; n22848
g22593 and n22735_not n22848_not ; n22849
g22594 and b[10] n22724_not ; n22850
g22595 and n22722_not n22850 ; n22851
g22596 and n22726_not n22851_not ; n22852
g22597 and n22849_not n22852 ; n22853
g22598 and n22726_not n22853_not ; n22854
g22599 and b[11] n22715_not ; n22855
g22600 and n22713_not n22855 ; n22856
g22601 and n22717_not n22856_not ; n22857
g22602 and n22854_not n22857 ; n22858
g22603 and n22717_not n22858_not ; n22859
g22604 and b[12] n22706_not ; n22860
g22605 and n22704_not n22860 ; n22861
g22606 and n22708_not n22861_not ; n22862
g22607 and n22859_not n22862 ; n22863
g22608 and n22708_not n22863_not ; n22864
g22609 and b[13] n22697_not ; n22865
g22610 and n22695_not n22865 ; n22866
g22611 and n22699_not n22866_not ; n22867
g22612 and n22864_not n22867 ; n22868
g22613 and n22699_not n22868_not ; n22869
g22614 and b[14] n22688_not ; n22870
g22615 and n22686_not n22870 ; n22871
g22616 and n22690_not n22871_not ; n22872
g22617 and n22869_not n22872 ; n22873
g22618 and n22690_not n22873_not ; n22874
g22619 and b[15] n22679_not ; n22875
g22620 and n22677_not n22875 ; n22876
g22621 and n22681_not n22876_not ; n22877
g22622 and n22874_not n22877 ; n22878
g22623 and n22681_not n22878_not ; n22879
g22624 and b[16] n22670_not ; n22880
g22625 and n22668_not n22880 ; n22881
g22626 and n22672_not n22881_not ; n22882
g22627 and n22879_not n22882 ; n22883
g22628 and n22672_not n22883_not ; n22884
g22629 and b[17] n22661_not ; n22885
g22630 and n22659_not n22885 ; n22886
g22631 and n22663_not n22886_not ; n22887
g22632 and n22884_not n22887 ; n22888
g22633 and n22663_not n22888_not ; n22889
g22634 and b[18] n22652_not ; n22890
g22635 and n22650_not n22890 ; n22891
g22636 and n22654_not n22891_not ; n22892
g22637 and n22889_not n22892 ; n22893
g22638 and n22654_not n22893_not ; n22894
g22639 and b[19] n22643_not ; n22895
g22640 and n22641_not n22895 ; n22896
g22641 and n22645_not n22896_not ; n22897
g22642 and n22894_not n22897 ; n22898
g22643 and n22645_not n22898_not ; n22899
g22644 and b[20] n22634_not ; n22900
g22645 and n22632_not n22900 ; n22901
g22646 and n22636_not n22901_not ; n22902
g22647 and n22899_not n22902 ; n22903
g22648 and n22636_not n22903_not ; n22904
g22649 and b[21] n22625_not ; n22905
g22650 and n22623_not n22905 ; n22906
g22651 and n22627_not n22906_not ; n22907
g22652 and n22904_not n22907 ; n22908
g22653 and n22627_not n22908_not ; n22909
g22654 and b[22] n22616_not ; n22910
g22655 and n22614_not n22910 ; n22911
g22656 and n22618_not n22911_not ; n22912
g22657 and n22909_not n22912 ; n22913
g22658 and n22618_not n22913_not ; n22914
g22659 and b[23] n22607_not ; n22915
g22660 and n22605_not n22915 ; n22916
g22661 and n22609_not n22916_not ; n22917
g22662 and n22914_not n22917 ; n22918
g22663 and n22609_not n22918_not ; n22919
g22664 and b[24] n22598_not ; n22920
g22665 and n22596_not n22920 ; n22921
g22666 and n22600_not n22921_not ; n22922
g22667 and n22919_not n22922 ; n22923
g22668 and n22600_not n22923_not ; n22924
g22669 and b[25] n22589_not ; n22925
g22670 and n22587_not n22925 ; n22926
g22671 and n22591_not n22926_not ; n22927
g22672 and n22924_not n22927 ; n22928
g22673 and n22591_not n22928_not ; n22929
g22674 and b[26] n22580_not ; n22930
g22675 and n22578_not n22930 ; n22931
g22676 and n22582_not n22931_not ; n22932
g22677 and n22929_not n22932 ; n22933
g22678 and n22582_not n22933_not ; n22934
g22679 and b[27] n22571_not ; n22935
g22680 and n22569_not n22935 ; n22936
g22681 and n22573_not n22936_not ; n22937
g22682 and n22934_not n22937 ; n22938
g22683 and n22573_not n22938_not ; n22939
g22684 and b[28] n22562_not ; n22940
g22685 and n22560_not n22940 ; n22941
g22686 and n22564_not n22941_not ; n22942
g22687 and n22939_not n22942 ; n22943
g22688 and n22564_not n22943_not ; n22944
g22689 and b[29] n22553_not ; n22945
g22690 and n22551_not n22945 ; n22946
g22691 and n22555_not n22946_not ; n22947
g22692 and n22944_not n22947 ; n22948
g22693 and n22555_not n22948_not ; n22949
g22694 and b[30] n22544_not ; n22950
g22695 and n22542_not n22950 ; n22951
g22696 and n22546_not n22951_not ; n22952
g22697 and n22949_not n22952 ; n22953
g22698 and n22546_not n22953_not ; n22954
g22699 and b[31] n22535_not ; n22955
g22700 and n22533_not n22955 ; n22956
g22701 and n22537_not n22956_not ; n22957
g22702 and n22954_not n22957 ; n22958
g22703 and n22537_not n22958_not ; n22959
g22704 and b[32] n22526_not ; n22960
g22705 and n22524_not n22960 ; n22961
g22706 and n22528_not n22961_not ; n22962
g22707 and n22959_not n22962 ; n22963
g22708 and n22528_not n22963_not ; n22964
g22709 and b[33] n22517_not ; n22965
g22710 and n22515_not n22965 ; n22966
g22711 and n22519_not n22966_not ; n22967
g22712 and n22964_not n22967 ; n22968
g22713 and n22519_not n22968_not ; n22969
g22714 and b[34] n22508_not ; n22970
g22715 and n22506_not n22970 ; n22971
g22716 and n22510_not n22971_not ; n22972
g22717 and n22969_not n22972 ; n22973
g22718 and n22510_not n22973_not ; n22974
g22719 and b[35] n22499_not ; n22975
g22720 and n22497_not n22975 ; n22976
g22721 and n22501_not n22976_not ; n22977
g22722 and n22974_not n22977 ; n22978
g22723 and n22501_not n22978_not ; n22979
g22724 and b[36] n22490_not ; n22980
g22725 and n22488_not n22980 ; n22981
g22726 and n22492_not n22981_not ; n22982
g22727 and n22979_not n22982 ; n22983
g22728 and n22492_not n22983_not ; n22984
g22729 and b[37] n22481_not ; n22985
g22730 and n22479_not n22985 ; n22986
g22731 and n22483_not n22986_not ; n22987
g22732 and n22984_not n22987 ; n22988
g22733 and n22483_not n22988_not ; n22989
g22734 and b[38] n22472_not ; n22990
g22735 and n22470_not n22990 ; n22991
g22736 and n22474_not n22991_not ; n22992
g22737 and n22989_not n22992 ; n22993
g22738 and n22474_not n22993_not ; n22994
g22739 and b[39] n22463_not ; n22995
g22740 and n22461_not n22995 ; n22996
g22741 and n22465_not n22996_not ; n22997
g22742 and n22994_not n22997 ; n22998
g22743 and n22465_not n22998_not ; n22999
g22744 and b[40] n22454_not ; n23000
g22745 and n22452_not n23000 ; n23001
g22746 and n22456_not n23001_not ; n23002
g22747 and n22999_not n23002 ; n23003
g22748 and n22456_not n23003_not ; n23004
g22749 and b[41] n22445_not ; n23005
g22750 and n22443_not n23005 ; n23006
g22751 and n22447_not n23006_not ; n23007
g22752 and n23004_not n23007 ; n23008
g22753 and n22447_not n23008_not ; n23009
g22754 and b[42] n22436_not ; n23010
g22755 and n22434_not n23010 ; n23011
g22756 and n22438_not n23011_not ; n23012
g22757 and n23009_not n23012 ; n23013
g22758 and n22438_not n23013_not ; n23014
g22759 and b[43] n22427_not ; n23015
g22760 and n22425_not n23015 ; n23016
g22761 and n22429_not n23016_not ; n23017
g22762 and n23014_not n23017 ; n23018
g22763 and n22429_not n23018_not ; n23019
g22764 and b[44] n22418_not ; n23020
g22765 and n22416_not n23020 ; n23021
g22766 and n22420_not n23021_not ; n23022
g22767 and n23019_not n23022 ; n23023
g22768 and n22420_not n23023_not ; n23024
g22769 and b[45] n22409_not ; n23025
g22770 and n22407_not n23025 ; n23026
g22771 and n22411_not n23026_not ; n23027
g22772 and n23024_not n23027 ; n23028
g22773 and n22411_not n23028_not ; n23029
g22774 and b[46] n22400_not ; n23030
g22775 and n22398_not n23030 ; n23031
g22776 and n22402_not n23031_not ; n23032
g22777 and n23029_not n23032 ; n23033
g22778 and n22402_not n23033_not ; n23034
g22779 and b[47] n22391_not ; n23035
g22780 and n22389_not n23035 ; n23036
g22781 and n22393_not n23036_not ; n23037
g22782 and n23034_not n23037 ; n23038
g22783 and n22393_not n23038_not ; n23039
g22784 and b[48] n22382_not ; n23040
g22785 and n22380_not n23040 ; n23041
g22786 and n22384_not n23041_not ; n23042
g22787 and n23039_not n23042 ; n23043
g22788 and n22384_not n23043_not ; n23044
g22789 and b[49] n22373_not ; n23045
g22790 and n22371_not n23045 ; n23046
g22791 and n22375_not n23046_not ; n23047
g22792 and n23044_not n23047 ; n23048
g22793 and n22375_not n23048_not ; n23049
g22794 and b[50] n22364_not ; n23050
g22795 and n22362_not n23050 ; n23051
g22796 and n22366_not n23051_not ; n23052
g22797 and n23049_not n23052 ; n23053
g22798 and n22366_not n23053_not ; n23054
g22799 and b[51] n22355_not ; n23055
g22800 and n22353_not n23055 ; n23056
g22801 and n22357_not n23056_not ; n23057
g22802 and n23054_not n23057 ; n23058
g22803 and n22357_not n23058_not ; n23059
g22804 and b[52] n22346_not ; n23060
g22805 and n22344_not n23060 ; n23061
g22806 and n22348_not n23061_not ; n23062
g22807 and n23059_not n23062 ; n23063
g22808 and n22348_not n23063_not ; n23064
g22809 and b[53] n22337_not ; n23065
g22810 and n22335_not n23065 ; n23066
g22811 and n22339_not n23066_not ; n23067
g22812 and n23064_not n23067 ; n23068
g22813 and n22339_not n23068_not ; n23069
g22814 and b[54] n22328_not ; n23070
g22815 and n22326_not n23070 ; n23071
g22816 and n22330_not n23071_not ; n23072
g22817 and n23069_not n23072 ; n23073
g22818 and n22330_not n23073_not ; n23074
g22819 and b[55] n22319_not ; n23075
g22820 and n22317_not n23075 ; n23076
g22821 and n22321_not n23076_not ; n23077
g22822 and n23074_not n23077 ; n23078
g22823 and n22321_not n23078_not ; n23079
g22824 and n21547_not n22307_not ; n23080
g22825 and n22305_not n23080 ; n23081
g22826 and n22296_not n23081 ; n23082
g22827 and n22305_not n22307_not ; n23083
g22828 and n22297_not n23083_not ; n23084
g22829 and n23082_not n23084_not ; n23085
g22830 and quotient[8] n23085_not ; n23086
g22831 and n22304_not n22311_not ; n23087
g22832 and n22310_not n23087 ; n23088
g22833 and n23086_not n23088_not ; n23089
g22834 and b[56]_not n23089_not ; n23090
g22835 and b[56] n23088_not ; n23091
g22836 and n23086_not n23091 ; n23092
g22837 and n407 n23092_not ; n23093
g22838 and n23090_not n23093 ; n23094
g22839 and n23079_not n23094 ; n23095
g22840 and n337 n23089_not ; n23096
g22841 and n23095_not n23096_not ; quotient[7]
g22842 and n22330_not n23077 ; n23098
g22843 and n23073_not n23098 ; n23099
g22844 and n23074_not n23077_not ; n23100
g22845 and n23099_not n23100_not ; n23101
g22846 and quotient[7] n23101_not ; n23102
g22847 and n22320_not n23096_not ; n23103
g22848 and n23095_not n23103 ; n23104
g22849 and n23102_not n23104_not ; n23105
g22850 and n22321_not n23092_not ; n23106
g22851 and n23090_not n23106 ; n23107
g22852 and n23078_not n23107 ; n23108
g22853 and n23090_not n23092_not ; n23109
g22854 and n23079_not n23109_not ; n23110
g22855 and n23108_not n23110_not ; n23111
g22856 and quotient[7] n23111_not ; n23112
g22857 and n23089_not n23096_not ; n23113
g22858 and n23095_not n23113 ; n23114
g22859 and n23112_not n23114_not ; n23115
g22860 and b[57]_not n23115_not ; n23116
g22861 and b[56]_not n23105_not ; n23117
g22862 and n22339_not n23072 ; n23118
g22863 and n23068_not n23118 ; n23119
g22864 and n23069_not n23072_not ; n23120
g22865 and n23119_not n23120_not ; n23121
g22866 and quotient[7] n23121_not ; n23122
g22867 and n22329_not n23096_not ; n23123
g22868 and n23095_not n23123 ; n23124
g22869 and n23122_not n23124_not ; n23125
g22870 and b[55]_not n23125_not ; n23126
g22871 and n22348_not n23067 ; n23127
g22872 and n23063_not n23127 ; n23128
g22873 and n23064_not n23067_not ; n23129
g22874 and n23128_not n23129_not ; n23130
g22875 and quotient[7] n23130_not ; n23131
g22876 and n22338_not n23096_not ; n23132
g22877 and n23095_not n23132 ; n23133
g22878 and n23131_not n23133_not ; n23134
g22879 and b[54]_not n23134_not ; n23135
g22880 and n22357_not n23062 ; n23136
g22881 and n23058_not n23136 ; n23137
g22882 and n23059_not n23062_not ; n23138
g22883 and n23137_not n23138_not ; n23139
g22884 and quotient[7] n23139_not ; n23140
g22885 and n22347_not n23096_not ; n23141
g22886 and n23095_not n23141 ; n23142
g22887 and n23140_not n23142_not ; n23143
g22888 and b[53]_not n23143_not ; n23144
g22889 and n22366_not n23057 ; n23145
g22890 and n23053_not n23145 ; n23146
g22891 and n23054_not n23057_not ; n23147
g22892 and n23146_not n23147_not ; n23148
g22893 and quotient[7] n23148_not ; n23149
g22894 and n22356_not n23096_not ; n23150
g22895 and n23095_not n23150 ; n23151
g22896 and n23149_not n23151_not ; n23152
g22897 and b[52]_not n23152_not ; n23153
g22898 and n22375_not n23052 ; n23154
g22899 and n23048_not n23154 ; n23155
g22900 and n23049_not n23052_not ; n23156
g22901 and n23155_not n23156_not ; n23157
g22902 and quotient[7] n23157_not ; n23158
g22903 and n22365_not n23096_not ; n23159
g22904 and n23095_not n23159 ; n23160
g22905 and n23158_not n23160_not ; n23161
g22906 and b[51]_not n23161_not ; n23162
g22907 and n22384_not n23047 ; n23163
g22908 and n23043_not n23163 ; n23164
g22909 and n23044_not n23047_not ; n23165
g22910 and n23164_not n23165_not ; n23166
g22911 and quotient[7] n23166_not ; n23167
g22912 and n22374_not n23096_not ; n23168
g22913 and n23095_not n23168 ; n23169
g22914 and n23167_not n23169_not ; n23170
g22915 and b[50]_not n23170_not ; n23171
g22916 and n22393_not n23042 ; n23172
g22917 and n23038_not n23172 ; n23173
g22918 and n23039_not n23042_not ; n23174
g22919 and n23173_not n23174_not ; n23175
g22920 and quotient[7] n23175_not ; n23176
g22921 and n22383_not n23096_not ; n23177
g22922 and n23095_not n23177 ; n23178
g22923 and n23176_not n23178_not ; n23179
g22924 and b[49]_not n23179_not ; n23180
g22925 and n22402_not n23037 ; n23181
g22926 and n23033_not n23181 ; n23182
g22927 and n23034_not n23037_not ; n23183
g22928 and n23182_not n23183_not ; n23184
g22929 and quotient[7] n23184_not ; n23185
g22930 and n22392_not n23096_not ; n23186
g22931 and n23095_not n23186 ; n23187
g22932 and n23185_not n23187_not ; n23188
g22933 and b[48]_not n23188_not ; n23189
g22934 and n22411_not n23032 ; n23190
g22935 and n23028_not n23190 ; n23191
g22936 and n23029_not n23032_not ; n23192
g22937 and n23191_not n23192_not ; n23193
g22938 and quotient[7] n23193_not ; n23194
g22939 and n22401_not n23096_not ; n23195
g22940 and n23095_not n23195 ; n23196
g22941 and n23194_not n23196_not ; n23197
g22942 and b[47]_not n23197_not ; n23198
g22943 and n22420_not n23027 ; n23199
g22944 and n23023_not n23199 ; n23200
g22945 and n23024_not n23027_not ; n23201
g22946 and n23200_not n23201_not ; n23202
g22947 and quotient[7] n23202_not ; n23203
g22948 and n22410_not n23096_not ; n23204
g22949 and n23095_not n23204 ; n23205
g22950 and n23203_not n23205_not ; n23206
g22951 and b[46]_not n23206_not ; n23207
g22952 and n22429_not n23022 ; n23208
g22953 and n23018_not n23208 ; n23209
g22954 and n23019_not n23022_not ; n23210
g22955 and n23209_not n23210_not ; n23211
g22956 and quotient[7] n23211_not ; n23212
g22957 and n22419_not n23096_not ; n23213
g22958 and n23095_not n23213 ; n23214
g22959 and n23212_not n23214_not ; n23215
g22960 and b[45]_not n23215_not ; n23216
g22961 and n22438_not n23017 ; n23217
g22962 and n23013_not n23217 ; n23218
g22963 and n23014_not n23017_not ; n23219
g22964 and n23218_not n23219_not ; n23220
g22965 and quotient[7] n23220_not ; n23221
g22966 and n22428_not n23096_not ; n23222
g22967 and n23095_not n23222 ; n23223
g22968 and n23221_not n23223_not ; n23224
g22969 and b[44]_not n23224_not ; n23225
g22970 and n22447_not n23012 ; n23226
g22971 and n23008_not n23226 ; n23227
g22972 and n23009_not n23012_not ; n23228
g22973 and n23227_not n23228_not ; n23229
g22974 and quotient[7] n23229_not ; n23230
g22975 and n22437_not n23096_not ; n23231
g22976 and n23095_not n23231 ; n23232
g22977 and n23230_not n23232_not ; n23233
g22978 and b[43]_not n23233_not ; n23234
g22979 and n22456_not n23007 ; n23235
g22980 and n23003_not n23235 ; n23236
g22981 and n23004_not n23007_not ; n23237
g22982 and n23236_not n23237_not ; n23238
g22983 and quotient[7] n23238_not ; n23239
g22984 and n22446_not n23096_not ; n23240
g22985 and n23095_not n23240 ; n23241
g22986 and n23239_not n23241_not ; n23242
g22987 and b[42]_not n23242_not ; n23243
g22988 and n22465_not n23002 ; n23244
g22989 and n22998_not n23244 ; n23245
g22990 and n22999_not n23002_not ; n23246
g22991 and n23245_not n23246_not ; n23247
g22992 and quotient[7] n23247_not ; n23248
g22993 and n22455_not n23096_not ; n23249
g22994 and n23095_not n23249 ; n23250
g22995 and n23248_not n23250_not ; n23251
g22996 and b[41]_not n23251_not ; n23252
g22997 and n22474_not n22997 ; n23253
g22998 and n22993_not n23253 ; n23254
g22999 and n22994_not n22997_not ; n23255
g23000 and n23254_not n23255_not ; n23256
g23001 and quotient[7] n23256_not ; n23257
g23002 and n22464_not n23096_not ; n23258
g23003 and n23095_not n23258 ; n23259
g23004 and n23257_not n23259_not ; n23260
g23005 and b[40]_not n23260_not ; n23261
g23006 and n22483_not n22992 ; n23262
g23007 and n22988_not n23262 ; n23263
g23008 and n22989_not n22992_not ; n23264
g23009 and n23263_not n23264_not ; n23265
g23010 and quotient[7] n23265_not ; n23266
g23011 and n22473_not n23096_not ; n23267
g23012 and n23095_not n23267 ; n23268
g23013 and n23266_not n23268_not ; n23269
g23014 and b[39]_not n23269_not ; n23270
g23015 and n22492_not n22987 ; n23271
g23016 and n22983_not n23271 ; n23272
g23017 and n22984_not n22987_not ; n23273
g23018 and n23272_not n23273_not ; n23274
g23019 and quotient[7] n23274_not ; n23275
g23020 and n22482_not n23096_not ; n23276
g23021 and n23095_not n23276 ; n23277
g23022 and n23275_not n23277_not ; n23278
g23023 and b[38]_not n23278_not ; n23279
g23024 and n22501_not n22982 ; n23280
g23025 and n22978_not n23280 ; n23281
g23026 and n22979_not n22982_not ; n23282
g23027 and n23281_not n23282_not ; n23283
g23028 and quotient[7] n23283_not ; n23284
g23029 and n22491_not n23096_not ; n23285
g23030 and n23095_not n23285 ; n23286
g23031 and n23284_not n23286_not ; n23287
g23032 and b[37]_not n23287_not ; n23288
g23033 and n22510_not n22977 ; n23289
g23034 and n22973_not n23289 ; n23290
g23035 and n22974_not n22977_not ; n23291
g23036 and n23290_not n23291_not ; n23292
g23037 and quotient[7] n23292_not ; n23293
g23038 and n22500_not n23096_not ; n23294
g23039 and n23095_not n23294 ; n23295
g23040 and n23293_not n23295_not ; n23296
g23041 and b[36]_not n23296_not ; n23297
g23042 and n22519_not n22972 ; n23298
g23043 and n22968_not n23298 ; n23299
g23044 and n22969_not n22972_not ; n23300
g23045 and n23299_not n23300_not ; n23301
g23046 and quotient[7] n23301_not ; n23302
g23047 and n22509_not n23096_not ; n23303
g23048 and n23095_not n23303 ; n23304
g23049 and n23302_not n23304_not ; n23305
g23050 and b[35]_not n23305_not ; n23306
g23051 and n22528_not n22967 ; n23307
g23052 and n22963_not n23307 ; n23308
g23053 and n22964_not n22967_not ; n23309
g23054 and n23308_not n23309_not ; n23310
g23055 and quotient[7] n23310_not ; n23311
g23056 and n22518_not n23096_not ; n23312
g23057 and n23095_not n23312 ; n23313
g23058 and n23311_not n23313_not ; n23314
g23059 and b[34]_not n23314_not ; n23315
g23060 and n22537_not n22962 ; n23316
g23061 and n22958_not n23316 ; n23317
g23062 and n22959_not n22962_not ; n23318
g23063 and n23317_not n23318_not ; n23319
g23064 and quotient[7] n23319_not ; n23320
g23065 and n22527_not n23096_not ; n23321
g23066 and n23095_not n23321 ; n23322
g23067 and n23320_not n23322_not ; n23323
g23068 and b[33]_not n23323_not ; n23324
g23069 and n22546_not n22957 ; n23325
g23070 and n22953_not n23325 ; n23326
g23071 and n22954_not n22957_not ; n23327
g23072 and n23326_not n23327_not ; n23328
g23073 and quotient[7] n23328_not ; n23329
g23074 and n22536_not n23096_not ; n23330
g23075 and n23095_not n23330 ; n23331
g23076 and n23329_not n23331_not ; n23332
g23077 and b[32]_not n23332_not ; n23333
g23078 and n22555_not n22952 ; n23334
g23079 and n22948_not n23334 ; n23335
g23080 and n22949_not n22952_not ; n23336
g23081 and n23335_not n23336_not ; n23337
g23082 and quotient[7] n23337_not ; n23338
g23083 and n22545_not n23096_not ; n23339
g23084 and n23095_not n23339 ; n23340
g23085 and n23338_not n23340_not ; n23341
g23086 and b[31]_not n23341_not ; n23342
g23087 and n22564_not n22947 ; n23343
g23088 and n22943_not n23343 ; n23344
g23089 and n22944_not n22947_not ; n23345
g23090 and n23344_not n23345_not ; n23346
g23091 and quotient[7] n23346_not ; n23347
g23092 and n22554_not n23096_not ; n23348
g23093 and n23095_not n23348 ; n23349
g23094 and n23347_not n23349_not ; n23350
g23095 and b[30]_not n23350_not ; n23351
g23096 and n22573_not n22942 ; n23352
g23097 and n22938_not n23352 ; n23353
g23098 and n22939_not n22942_not ; n23354
g23099 and n23353_not n23354_not ; n23355
g23100 and quotient[7] n23355_not ; n23356
g23101 and n22563_not n23096_not ; n23357
g23102 and n23095_not n23357 ; n23358
g23103 and n23356_not n23358_not ; n23359
g23104 and b[29]_not n23359_not ; n23360
g23105 and n22582_not n22937 ; n23361
g23106 and n22933_not n23361 ; n23362
g23107 and n22934_not n22937_not ; n23363
g23108 and n23362_not n23363_not ; n23364
g23109 and quotient[7] n23364_not ; n23365
g23110 and n22572_not n23096_not ; n23366
g23111 and n23095_not n23366 ; n23367
g23112 and n23365_not n23367_not ; n23368
g23113 and b[28]_not n23368_not ; n23369
g23114 and n22591_not n22932 ; n23370
g23115 and n22928_not n23370 ; n23371
g23116 and n22929_not n22932_not ; n23372
g23117 and n23371_not n23372_not ; n23373
g23118 and quotient[7] n23373_not ; n23374
g23119 and n22581_not n23096_not ; n23375
g23120 and n23095_not n23375 ; n23376
g23121 and n23374_not n23376_not ; n23377
g23122 and b[27]_not n23377_not ; n23378
g23123 and n22600_not n22927 ; n23379
g23124 and n22923_not n23379 ; n23380
g23125 and n22924_not n22927_not ; n23381
g23126 and n23380_not n23381_not ; n23382
g23127 and quotient[7] n23382_not ; n23383
g23128 and n22590_not n23096_not ; n23384
g23129 and n23095_not n23384 ; n23385
g23130 and n23383_not n23385_not ; n23386
g23131 and b[26]_not n23386_not ; n23387
g23132 and n22609_not n22922 ; n23388
g23133 and n22918_not n23388 ; n23389
g23134 and n22919_not n22922_not ; n23390
g23135 and n23389_not n23390_not ; n23391
g23136 and quotient[7] n23391_not ; n23392
g23137 and n22599_not n23096_not ; n23393
g23138 and n23095_not n23393 ; n23394
g23139 and n23392_not n23394_not ; n23395
g23140 and b[25]_not n23395_not ; n23396
g23141 and n22618_not n22917 ; n23397
g23142 and n22913_not n23397 ; n23398
g23143 and n22914_not n22917_not ; n23399
g23144 and n23398_not n23399_not ; n23400
g23145 and quotient[7] n23400_not ; n23401
g23146 and n22608_not n23096_not ; n23402
g23147 and n23095_not n23402 ; n23403
g23148 and n23401_not n23403_not ; n23404
g23149 and b[24]_not n23404_not ; n23405
g23150 and n22627_not n22912 ; n23406
g23151 and n22908_not n23406 ; n23407
g23152 and n22909_not n22912_not ; n23408
g23153 and n23407_not n23408_not ; n23409
g23154 and quotient[7] n23409_not ; n23410
g23155 and n22617_not n23096_not ; n23411
g23156 and n23095_not n23411 ; n23412
g23157 and n23410_not n23412_not ; n23413
g23158 and b[23]_not n23413_not ; n23414
g23159 and n22636_not n22907 ; n23415
g23160 and n22903_not n23415 ; n23416
g23161 and n22904_not n22907_not ; n23417
g23162 and n23416_not n23417_not ; n23418
g23163 and quotient[7] n23418_not ; n23419
g23164 and n22626_not n23096_not ; n23420
g23165 and n23095_not n23420 ; n23421
g23166 and n23419_not n23421_not ; n23422
g23167 and b[22]_not n23422_not ; n23423
g23168 and n22645_not n22902 ; n23424
g23169 and n22898_not n23424 ; n23425
g23170 and n22899_not n22902_not ; n23426
g23171 and n23425_not n23426_not ; n23427
g23172 and quotient[7] n23427_not ; n23428
g23173 and n22635_not n23096_not ; n23429
g23174 and n23095_not n23429 ; n23430
g23175 and n23428_not n23430_not ; n23431
g23176 and b[21]_not n23431_not ; n23432
g23177 and n22654_not n22897 ; n23433
g23178 and n22893_not n23433 ; n23434
g23179 and n22894_not n22897_not ; n23435
g23180 and n23434_not n23435_not ; n23436
g23181 and quotient[7] n23436_not ; n23437
g23182 and n22644_not n23096_not ; n23438
g23183 and n23095_not n23438 ; n23439
g23184 and n23437_not n23439_not ; n23440
g23185 and b[20]_not n23440_not ; n23441
g23186 and n22663_not n22892 ; n23442
g23187 and n22888_not n23442 ; n23443
g23188 and n22889_not n22892_not ; n23444
g23189 and n23443_not n23444_not ; n23445
g23190 and quotient[7] n23445_not ; n23446
g23191 and n22653_not n23096_not ; n23447
g23192 and n23095_not n23447 ; n23448
g23193 and n23446_not n23448_not ; n23449
g23194 and b[19]_not n23449_not ; n23450
g23195 and n22672_not n22887 ; n23451
g23196 and n22883_not n23451 ; n23452
g23197 and n22884_not n22887_not ; n23453
g23198 and n23452_not n23453_not ; n23454
g23199 and quotient[7] n23454_not ; n23455
g23200 and n22662_not n23096_not ; n23456
g23201 and n23095_not n23456 ; n23457
g23202 and n23455_not n23457_not ; n23458
g23203 and b[18]_not n23458_not ; n23459
g23204 and n22681_not n22882 ; n23460
g23205 and n22878_not n23460 ; n23461
g23206 and n22879_not n22882_not ; n23462
g23207 and n23461_not n23462_not ; n23463
g23208 and quotient[7] n23463_not ; n23464
g23209 and n22671_not n23096_not ; n23465
g23210 and n23095_not n23465 ; n23466
g23211 and n23464_not n23466_not ; n23467
g23212 and b[17]_not n23467_not ; n23468
g23213 and n22690_not n22877 ; n23469
g23214 and n22873_not n23469 ; n23470
g23215 and n22874_not n22877_not ; n23471
g23216 and n23470_not n23471_not ; n23472
g23217 and quotient[7] n23472_not ; n23473
g23218 and n22680_not n23096_not ; n23474
g23219 and n23095_not n23474 ; n23475
g23220 and n23473_not n23475_not ; n23476
g23221 and b[16]_not n23476_not ; n23477
g23222 and n22699_not n22872 ; n23478
g23223 and n22868_not n23478 ; n23479
g23224 and n22869_not n22872_not ; n23480
g23225 and n23479_not n23480_not ; n23481
g23226 and quotient[7] n23481_not ; n23482
g23227 and n22689_not n23096_not ; n23483
g23228 and n23095_not n23483 ; n23484
g23229 and n23482_not n23484_not ; n23485
g23230 and b[15]_not n23485_not ; n23486
g23231 and n22708_not n22867 ; n23487
g23232 and n22863_not n23487 ; n23488
g23233 and n22864_not n22867_not ; n23489
g23234 and n23488_not n23489_not ; n23490
g23235 and quotient[7] n23490_not ; n23491
g23236 and n22698_not n23096_not ; n23492
g23237 and n23095_not n23492 ; n23493
g23238 and n23491_not n23493_not ; n23494
g23239 and b[14]_not n23494_not ; n23495
g23240 and n22717_not n22862 ; n23496
g23241 and n22858_not n23496 ; n23497
g23242 and n22859_not n22862_not ; n23498
g23243 and n23497_not n23498_not ; n23499
g23244 and quotient[7] n23499_not ; n23500
g23245 and n22707_not n23096_not ; n23501
g23246 and n23095_not n23501 ; n23502
g23247 and n23500_not n23502_not ; n23503
g23248 and b[13]_not n23503_not ; n23504
g23249 and n22726_not n22857 ; n23505
g23250 and n22853_not n23505 ; n23506
g23251 and n22854_not n22857_not ; n23507
g23252 and n23506_not n23507_not ; n23508
g23253 and quotient[7] n23508_not ; n23509
g23254 and n22716_not n23096_not ; n23510
g23255 and n23095_not n23510 ; n23511
g23256 and n23509_not n23511_not ; n23512
g23257 and b[12]_not n23512_not ; n23513
g23258 and n22735_not n22852 ; n23514
g23259 and n22848_not n23514 ; n23515
g23260 and n22849_not n22852_not ; n23516
g23261 and n23515_not n23516_not ; n23517
g23262 and quotient[7] n23517_not ; n23518
g23263 and n22725_not n23096_not ; n23519
g23264 and n23095_not n23519 ; n23520
g23265 and n23518_not n23520_not ; n23521
g23266 and b[11]_not n23521_not ; n23522
g23267 and n22744_not n22847 ; n23523
g23268 and n22843_not n23523 ; n23524
g23269 and n22844_not n22847_not ; n23525
g23270 and n23524_not n23525_not ; n23526
g23271 and quotient[7] n23526_not ; n23527
g23272 and n22734_not n23096_not ; n23528
g23273 and n23095_not n23528 ; n23529
g23274 and n23527_not n23529_not ; n23530
g23275 and b[10]_not n23530_not ; n23531
g23276 and n22753_not n22842 ; n23532
g23277 and n22838_not n23532 ; n23533
g23278 and n22839_not n22842_not ; n23534
g23279 and n23533_not n23534_not ; n23535
g23280 and quotient[7] n23535_not ; n23536
g23281 and n22743_not n23096_not ; n23537
g23282 and n23095_not n23537 ; n23538
g23283 and n23536_not n23538_not ; n23539
g23284 and b[9]_not n23539_not ; n23540
g23285 and n22762_not n22837 ; n23541
g23286 and n22833_not n23541 ; n23542
g23287 and n22834_not n22837_not ; n23543
g23288 and n23542_not n23543_not ; n23544
g23289 and quotient[7] n23544_not ; n23545
g23290 and n22752_not n23096_not ; n23546
g23291 and n23095_not n23546 ; n23547
g23292 and n23545_not n23547_not ; n23548
g23293 and b[8]_not n23548_not ; n23549
g23294 and n22771_not n22832 ; n23550
g23295 and n22828_not n23550 ; n23551
g23296 and n22829_not n22832_not ; n23552
g23297 and n23551_not n23552_not ; n23553
g23298 and quotient[7] n23553_not ; n23554
g23299 and n22761_not n23096_not ; n23555
g23300 and n23095_not n23555 ; n23556
g23301 and n23554_not n23556_not ; n23557
g23302 and b[7]_not n23557_not ; n23558
g23303 and n22780_not n22827 ; n23559
g23304 and n22823_not n23559 ; n23560
g23305 and n22824_not n22827_not ; n23561
g23306 and n23560_not n23561_not ; n23562
g23307 and quotient[7] n23562_not ; n23563
g23308 and n22770_not n23096_not ; n23564
g23309 and n23095_not n23564 ; n23565
g23310 and n23563_not n23565_not ; n23566
g23311 and b[6]_not n23566_not ; n23567
g23312 and n22789_not n22822 ; n23568
g23313 and n22818_not n23568 ; n23569
g23314 and n22819_not n22822_not ; n23570
g23315 and n23569_not n23570_not ; n23571
g23316 and quotient[7] n23571_not ; n23572
g23317 and n22779_not n23096_not ; n23573
g23318 and n23095_not n23573 ; n23574
g23319 and n23572_not n23574_not ; n23575
g23320 and b[5]_not n23575_not ; n23576
g23321 and n22797_not n22817 ; n23577
g23322 and n22813_not n23577 ; n23578
g23323 and n22814_not n22817_not ; n23579
g23324 and n23578_not n23579_not ; n23580
g23325 and quotient[7] n23580_not ; n23581
g23326 and n22788_not n23096_not ; n23582
g23327 and n23095_not n23582 ; n23583
g23328 and n23581_not n23583_not ; n23584
g23329 and b[4]_not n23584_not ; n23585
g23330 and n22808_not n22812 ; n23586
g23331 and n22807_not n23586 ; n23587
g23332 and n22809_not n22812_not ; n23588
g23333 and n23587_not n23588_not ; n23589
g23334 and quotient[7] n23589_not ; n23590
g23335 and n22796_not n23096_not ; n23591
g23336 and n23095_not n23591 ; n23592
g23337 and n23590_not n23592_not ; n23593
g23338 and b[3]_not n23593_not ; n23594
g23339 and n22804_not n22806 ; n23595
g23340 and n22802_not n23595 ; n23596
g23341 and n22807_not n23596_not ; n23597
g23342 and quotient[7] n23597 ; n23598
g23343 and n22801_not n23096_not ; n23599
g23344 and n23095_not n23599 ; n23600
g23345 and n23598_not n23600_not ; n23601
g23346 and b[2]_not n23601_not ; n23602
g23347 and b[0] quotient[7] ; n23603
g23348 and a[7] n23603_not ; n23604
g23349 and n22806 quotient[7] ; n23605
g23350 and n23604_not n23605_not ; n23606
g23351 and b[1] n23606_not ; n23607
g23352 and b[1]_not n23605_not ; n23608
g23353 and n23604_not n23608 ; n23609
g23354 and n23607_not n23609_not ; n23610
g23355 and a[6]_not b[0] ; n23611
g23356 and n23610_not n23611_not ; n23612
g23357 and b[1]_not n23606_not ; n23613
g23358 and n23612_not n23613_not ; n23614
g23359 and b[2] n23600_not ; n23615
g23360 and n23598_not n23615 ; n23616
g23361 and n23602_not n23616_not ; n23617
g23362 and n23614_not n23617 ; n23618
g23363 and n23602_not n23618_not ; n23619
g23364 and b[3] n23592_not ; n23620
g23365 and n23590_not n23620 ; n23621
g23366 and n23594_not n23621_not ; n23622
g23367 and n23619_not n23622 ; n23623
g23368 and n23594_not n23623_not ; n23624
g23369 and b[4] n23583_not ; n23625
g23370 and n23581_not n23625 ; n23626
g23371 and n23585_not n23626_not ; n23627
g23372 and n23624_not n23627 ; n23628
g23373 and n23585_not n23628_not ; n23629
g23374 and b[5] n23574_not ; n23630
g23375 and n23572_not n23630 ; n23631
g23376 and n23576_not n23631_not ; n23632
g23377 and n23629_not n23632 ; n23633
g23378 and n23576_not n23633_not ; n23634
g23379 and b[6] n23565_not ; n23635
g23380 and n23563_not n23635 ; n23636
g23381 and n23567_not n23636_not ; n23637
g23382 and n23634_not n23637 ; n23638
g23383 and n23567_not n23638_not ; n23639
g23384 and b[7] n23556_not ; n23640
g23385 and n23554_not n23640 ; n23641
g23386 and n23558_not n23641_not ; n23642
g23387 and n23639_not n23642 ; n23643
g23388 and n23558_not n23643_not ; n23644
g23389 and b[8] n23547_not ; n23645
g23390 and n23545_not n23645 ; n23646
g23391 and n23549_not n23646_not ; n23647
g23392 and n23644_not n23647 ; n23648
g23393 and n23549_not n23648_not ; n23649
g23394 and b[9] n23538_not ; n23650
g23395 and n23536_not n23650 ; n23651
g23396 and n23540_not n23651_not ; n23652
g23397 and n23649_not n23652 ; n23653
g23398 and n23540_not n23653_not ; n23654
g23399 and b[10] n23529_not ; n23655
g23400 and n23527_not n23655 ; n23656
g23401 and n23531_not n23656_not ; n23657
g23402 and n23654_not n23657 ; n23658
g23403 and n23531_not n23658_not ; n23659
g23404 and b[11] n23520_not ; n23660
g23405 and n23518_not n23660 ; n23661
g23406 and n23522_not n23661_not ; n23662
g23407 and n23659_not n23662 ; n23663
g23408 and n23522_not n23663_not ; n23664
g23409 and b[12] n23511_not ; n23665
g23410 and n23509_not n23665 ; n23666
g23411 and n23513_not n23666_not ; n23667
g23412 and n23664_not n23667 ; n23668
g23413 and n23513_not n23668_not ; n23669
g23414 and b[13] n23502_not ; n23670
g23415 and n23500_not n23670 ; n23671
g23416 and n23504_not n23671_not ; n23672
g23417 and n23669_not n23672 ; n23673
g23418 and n23504_not n23673_not ; n23674
g23419 and b[14] n23493_not ; n23675
g23420 and n23491_not n23675 ; n23676
g23421 and n23495_not n23676_not ; n23677
g23422 and n23674_not n23677 ; n23678
g23423 and n23495_not n23678_not ; n23679
g23424 and b[15] n23484_not ; n23680
g23425 and n23482_not n23680 ; n23681
g23426 and n23486_not n23681_not ; n23682
g23427 and n23679_not n23682 ; n23683
g23428 and n23486_not n23683_not ; n23684
g23429 and b[16] n23475_not ; n23685
g23430 and n23473_not n23685 ; n23686
g23431 and n23477_not n23686_not ; n23687
g23432 and n23684_not n23687 ; n23688
g23433 and n23477_not n23688_not ; n23689
g23434 and b[17] n23466_not ; n23690
g23435 and n23464_not n23690 ; n23691
g23436 and n23468_not n23691_not ; n23692
g23437 and n23689_not n23692 ; n23693
g23438 and n23468_not n23693_not ; n23694
g23439 and b[18] n23457_not ; n23695
g23440 and n23455_not n23695 ; n23696
g23441 and n23459_not n23696_not ; n23697
g23442 and n23694_not n23697 ; n23698
g23443 and n23459_not n23698_not ; n23699
g23444 and b[19] n23448_not ; n23700
g23445 and n23446_not n23700 ; n23701
g23446 and n23450_not n23701_not ; n23702
g23447 and n23699_not n23702 ; n23703
g23448 and n23450_not n23703_not ; n23704
g23449 and b[20] n23439_not ; n23705
g23450 and n23437_not n23705 ; n23706
g23451 and n23441_not n23706_not ; n23707
g23452 and n23704_not n23707 ; n23708
g23453 and n23441_not n23708_not ; n23709
g23454 and b[21] n23430_not ; n23710
g23455 and n23428_not n23710 ; n23711
g23456 and n23432_not n23711_not ; n23712
g23457 and n23709_not n23712 ; n23713
g23458 and n23432_not n23713_not ; n23714
g23459 and b[22] n23421_not ; n23715
g23460 and n23419_not n23715 ; n23716
g23461 and n23423_not n23716_not ; n23717
g23462 and n23714_not n23717 ; n23718
g23463 and n23423_not n23718_not ; n23719
g23464 and b[23] n23412_not ; n23720
g23465 and n23410_not n23720 ; n23721
g23466 and n23414_not n23721_not ; n23722
g23467 and n23719_not n23722 ; n23723
g23468 and n23414_not n23723_not ; n23724
g23469 and b[24] n23403_not ; n23725
g23470 and n23401_not n23725 ; n23726
g23471 and n23405_not n23726_not ; n23727
g23472 and n23724_not n23727 ; n23728
g23473 and n23405_not n23728_not ; n23729
g23474 and b[25] n23394_not ; n23730
g23475 and n23392_not n23730 ; n23731
g23476 and n23396_not n23731_not ; n23732
g23477 and n23729_not n23732 ; n23733
g23478 and n23396_not n23733_not ; n23734
g23479 and b[26] n23385_not ; n23735
g23480 and n23383_not n23735 ; n23736
g23481 and n23387_not n23736_not ; n23737
g23482 and n23734_not n23737 ; n23738
g23483 and n23387_not n23738_not ; n23739
g23484 and b[27] n23376_not ; n23740
g23485 and n23374_not n23740 ; n23741
g23486 and n23378_not n23741_not ; n23742
g23487 and n23739_not n23742 ; n23743
g23488 and n23378_not n23743_not ; n23744
g23489 and b[28] n23367_not ; n23745
g23490 and n23365_not n23745 ; n23746
g23491 and n23369_not n23746_not ; n23747
g23492 and n23744_not n23747 ; n23748
g23493 and n23369_not n23748_not ; n23749
g23494 and b[29] n23358_not ; n23750
g23495 and n23356_not n23750 ; n23751
g23496 and n23360_not n23751_not ; n23752
g23497 and n23749_not n23752 ; n23753
g23498 and n23360_not n23753_not ; n23754
g23499 and b[30] n23349_not ; n23755
g23500 and n23347_not n23755 ; n23756
g23501 and n23351_not n23756_not ; n23757
g23502 and n23754_not n23757 ; n23758
g23503 and n23351_not n23758_not ; n23759
g23504 and b[31] n23340_not ; n23760
g23505 and n23338_not n23760 ; n23761
g23506 and n23342_not n23761_not ; n23762
g23507 and n23759_not n23762 ; n23763
g23508 and n23342_not n23763_not ; n23764
g23509 and b[32] n23331_not ; n23765
g23510 and n23329_not n23765 ; n23766
g23511 and n23333_not n23766_not ; n23767
g23512 and n23764_not n23767 ; n23768
g23513 and n23333_not n23768_not ; n23769
g23514 and b[33] n23322_not ; n23770
g23515 and n23320_not n23770 ; n23771
g23516 and n23324_not n23771_not ; n23772
g23517 and n23769_not n23772 ; n23773
g23518 and n23324_not n23773_not ; n23774
g23519 and b[34] n23313_not ; n23775
g23520 and n23311_not n23775 ; n23776
g23521 and n23315_not n23776_not ; n23777
g23522 and n23774_not n23777 ; n23778
g23523 and n23315_not n23778_not ; n23779
g23524 and b[35] n23304_not ; n23780
g23525 and n23302_not n23780 ; n23781
g23526 and n23306_not n23781_not ; n23782
g23527 and n23779_not n23782 ; n23783
g23528 and n23306_not n23783_not ; n23784
g23529 and b[36] n23295_not ; n23785
g23530 and n23293_not n23785 ; n23786
g23531 and n23297_not n23786_not ; n23787
g23532 and n23784_not n23787 ; n23788
g23533 and n23297_not n23788_not ; n23789
g23534 and b[37] n23286_not ; n23790
g23535 and n23284_not n23790 ; n23791
g23536 and n23288_not n23791_not ; n23792
g23537 and n23789_not n23792 ; n23793
g23538 and n23288_not n23793_not ; n23794
g23539 and b[38] n23277_not ; n23795
g23540 and n23275_not n23795 ; n23796
g23541 and n23279_not n23796_not ; n23797
g23542 and n23794_not n23797 ; n23798
g23543 and n23279_not n23798_not ; n23799
g23544 and b[39] n23268_not ; n23800
g23545 and n23266_not n23800 ; n23801
g23546 and n23270_not n23801_not ; n23802
g23547 and n23799_not n23802 ; n23803
g23548 and n23270_not n23803_not ; n23804
g23549 and b[40] n23259_not ; n23805
g23550 and n23257_not n23805 ; n23806
g23551 and n23261_not n23806_not ; n23807
g23552 and n23804_not n23807 ; n23808
g23553 and n23261_not n23808_not ; n23809
g23554 and b[41] n23250_not ; n23810
g23555 and n23248_not n23810 ; n23811
g23556 and n23252_not n23811_not ; n23812
g23557 and n23809_not n23812 ; n23813
g23558 and n23252_not n23813_not ; n23814
g23559 and b[42] n23241_not ; n23815
g23560 and n23239_not n23815 ; n23816
g23561 and n23243_not n23816_not ; n23817
g23562 and n23814_not n23817 ; n23818
g23563 and n23243_not n23818_not ; n23819
g23564 and b[43] n23232_not ; n23820
g23565 and n23230_not n23820 ; n23821
g23566 and n23234_not n23821_not ; n23822
g23567 and n23819_not n23822 ; n23823
g23568 and n23234_not n23823_not ; n23824
g23569 and b[44] n23223_not ; n23825
g23570 and n23221_not n23825 ; n23826
g23571 and n23225_not n23826_not ; n23827
g23572 and n23824_not n23827 ; n23828
g23573 and n23225_not n23828_not ; n23829
g23574 and b[45] n23214_not ; n23830
g23575 and n23212_not n23830 ; n23831
g23576 and n23216_not n23831_not ; n23832
g23577 and n23829_not n23832 ; n23833
g23578 and n23216_not n23833_not ; n23834
g23579 and b[46] n23205_not ; n23835
g23580 and n23203_not n23835 ; n23836
g23581 and n23207_not n23836_not ; n23837
g23582 and n23834_not n23837 ; n23838
g23583 and n23207_not n23838_not ; n23839
g23584 and b[47] n23196_not ; n23840
g23585 and n23194_not n23840 ; n23841
g23586 and n23198_not n23841_not ; n23842
g23587 and n23839_not n23842 ; n23843
g23588 and n23198_not n23843_not ; n23844
g23589 and b[48] n23187_not ; n23845
g23590 and n23185_not n23845 ; n23846
g23591 and n23189_not n23846_not ; n23847
g23592 and n23844_not n23847 ; n23848
g23593 and n23189_not n23848_not ; n23849
g23594 and b[49] n23178_not ; n23850
g23595 and n23176_not n23850 ; n23851
g23596 and n23180_not n23851_not ; n23852
g23597 and n23849_not n23852 ; n23853
g23598 and n23180_not n23853_not ; n23854
g23599 and b[50] n23169_not ; n23855
g23600 and n23167_not n23855 ; n23856
g23601 and n23171_not n23856_not ; n23857
g23602 and n23854_not n23857 ; n23858
g23603 and n23171_not n23858_not ; n23859
g23604 and b[51] n23160_not ; n23860
g23605 and n23158_not n23860 ; n23861
g23606 and n23162_not n23861_not ; n23862
g23607 and n23859_not n23862 ; n23863
g23608 and n23162_not n23863_not ; n23864
g23609 and b[52] n23151_not ; n23865
g23610 and n23149_not n23865 ; n23866
g23611 and n23153_not n23866_not ; n23867
g23612 and n23864_not n23867 ; n23868
g23613 and n23153_not n23868_not ; n23869
g23614 and b[53] n23142_not ; n23870
g23615 and n23140_not n23870 ; n23871
g23616 and n23144_not n23871_not ; n23872
g23617 and n23869_not n23872 ; n23873
g23618 and n23144_not n23873_not ; n23874
g23619 and b[54] n23133_not ; n23875
g23620 and n23131_not n23875 ; n23876
g23621 and n23135_not n23876_not ; n23877
g23622 and n23874_not n23877 ; n23878
g23623 and n23135_not n23878_not ; n23879
g23624 and b[55] n23124_not ; n23880
g23625 and n23122_not n23880 ; n23881
g23626 and n23126_not n23881_not ; n23882
g23627 and n23879_not n23882 ; n23883
g23628 and n23126_not n23883_not ; n23884
g23629 and b[56] n23104_not ; n23885
g23630 and n23102_not n23885 ; n23886
g23631 and n23117_not n23886_not ; n23887
g23632 and n23884_not n23887 ; n23888
g23633 and n23117_not n23888_not ; n23889
g23634 and b[57] n23114_not ; n23890
g23635 and n23112_not n23890 ; n23891
g23636 and n23116_not n23891_not ; n23892
g23637 and n23889_not n23892 ; n23893
g23638 and n23116_not n23893_not ; n23894
g23639 and n280 n282 ; n23895
g23640 and n23894_not n23895 ; quotient[6]
g23641 and n23105_not quotient[6]_not ; n23897
g23642 and n23126_not n23887 ; n23898
g23643 and n23883_not n23898 ; n23899
g23644 and n23884_not n23887_not ; n23900
g23645 and n23899_not n23900_not ; n23901
g23646 and n23895 n23901_not ; n23902
g23647 and n23894_not n23902 ; n23903
g23648 and n23897_not n23903_not ; n23904
g23649 and b[57]_not n23904_not ; n23905
g23650 and n23125_not quotient[6]_not ; n23906
g23651 and n23135_not n23882 ; n23907
g23652 and n23878_not n23907 ; n23908
g23653 and n23879_not n23882_not ; n23909
g23654 and n23908_not n23909_not ; n23910
g23655 and n23895 n23910_not ; n23911
g23656 and n23894_not n23911 ; n23912
g23657 and n23906_not n23912_not ; n23913
g23658 and b[56]_not n23913_not ; n23914
g23659 and n23134_not quotient[6]_not ; n23915
g23660 and n23144_not n23877 ; n23916
g23661 and n23873_not n23916 ; n23917
g23662 and n23874_not n23877_not ; n23918
g23663 and n23917_not n23918_not ; n23919
g23664 and n23895 n23919_not ; n23920
g23665 and n23894_not n23920 ; n23921
g23666 and n23915_not n23921_not ; n23922
g23667 and b[55]_not n23922_not ; n23923
g23668 and n23143_not quotient[6]_not ; n23924
g23669 and n23153_not n23872 ; n23925
g23670 and n23868_not n23925 ; n23926
g23671 and n23869_not n23872_not ; n23927
g23672 and n23926_not n23927_not ; n23928
g23673 and n23895 n23928_not ; n23929
g23674 and n23894_not n23929 ; n23930
g23675 and n23924_not n23930_not ; n23931
g23676 and b[54]_not n23931_not ; n23932
g23677 and n23152_not quotient[6]_not ; n23933
g23678 and n23162_not n23867 ; n23934
g23679 and n23863_not n23934 ; n23935
g23680 and n23864_not n23867_not ; n23936
g23681 and n23935_not n23936_not ; n23937
g23682 and n23895 n23937_not ; n23938
g23683 and n23894_not n23938 ; n23939
g23684 and n23933_not n23939_not ; n23940
g23685 and b[53]_not n23940_not ; n23941
g23686 and n23161_not quotient[6]_not ; n23942
g23687 and n23171_not n23862 ; n23943
g23688 and n23858_not n23943 ; n23944
g23689 and n23859_not n23862_not ; n23945
g23690 and n23944_not n23945_not ; n23946
g23691 and n23895 n23946_not ; n23947
g23692 and n23894_not n23947 ; n23948
g23693 and n23942_not n23948_not ; n23949
g23694 and b[52]_not n23949_not ; n23950
g23695 and n23170_not quotient[6]_not ; n23951
g23696 and n23180_not n23857 ; n23952
g23697 and n23853_not n23952 ; n23953
g23698 and n23854_not n23857_not ; n23954
g23699 and n23953_not n23954_not ; n23955
g23700 and n23895 n23955_not ; n23956
g23701 and n23894_not n23956 ; n23957
g23702 and n23951_not n23957_not ; n23958
g23703 and b[51]_not n23958_not ; n23959
g23704 and n23179_not quotient[6]_not ; n23960
g23705 and n23189_not n23852 ; n23961
g23706 and n23848_not n23961 ; n23962
g23707 and n23849_not n23852_not ; n23963
g23708 and n23962_not n23963_not ; n23964
g23709 and n23895 n23964_not ; n23965
g23710 and n23894_not n23965 ; n23966
g23711 and n23960_not n23966_not ; n23967
g23712 and b[50]_not n23967_not ; n23968
g23713 and n23188_not quotient[6]_not ; n23969
g23714 and n23198_not n23847 ; n23970
g23715 and n23843_not n23970 ; n23971
g23716 and n23844_not n23847_not ; n23972
g23717 and n23971_not n23972_not ; n23973
g23718 and n23895 n23973_not ; n23974
g23719 and n23894_not n23974 ; n23975
g23720 and n23969_not n23975_not ; n23976
g23721 and b[49]_not n23976_not ; n23977
g23722 and n23197_not quotient[6]_not ; n23978
g23723 and n23207_not n23842 ; n23979
g23724 and n23838_not n23979 ; n23980
g23725 and n23839_not n23842_not ; n23981
g23726 and n23980_not n23981_not ; n23982
g23727 and n23895 n23982_not ; n23983
g23728 and n23894_not n23983 ; n23984
g23729 and n23978_not n23984_not ; n23985
g23730 and b[48]_not n23985_not ; n23986
g23731 and n23206_not quotient[6]_not ; n23987
g23732 and n23216_not n23837 ; n23988
g23733 and n23833_not n23988 ; n23989
g23734 and n23834_not n23837_not ; n23990
g23735 and n23989_not n23990_not ; n23991
g23736 and n23895 n23991_not ; n23992
g23737 and n23894_not n23992 ; n23993
g23738 and n23987_not n23993_not ; n23994
g23739 and b[47]_not n23994_not ; n23995
g23740 and n23215_not quotient[6]_not ; n23996
g23741 and n23225_not n23832 ; n23997
g23742 and n23828_not n23997 ; n23998
g23743 and n23829_not n23832_not ; n23999
g23744 and n23998_not n23999_not ; n24000
g23745 and n23895 n24000_not ; n24001
g23746 and n23894_not n24001 ; n24002
g23747 and n23996_not n24002_not ; n24003
g23748 and b[46]_not n24003_not ; n24004
g23749 and n23224_not quotient[6]_not ; n24005
g23750 and n23234_not n23827 ; n24006
g23751 and n23823_not n24006 ; n24007
g23752 and n23824_not n23827_not ; n24008
g23753 and n24007_not n24008_not ; n24009
g23754 and n23895 n24009_not ; n24010
g23755 and n23894_not n24010 ; n24011
g23756 and n24005_not n24011_not ; n24012
g23757 and b[45]_not n24012_not ; n24013
g23758 and n23233_not quotient[6]_not ; n24014
g23759 and n23243_not n23822 ; n24015
g23760 and n23818_not n24015 ; n24016
g23761 and n23819_not n23822_not ; n24017
g23762 and n24016_not n24017_not ; n24018
g23763 and n23895 n24018_not ; n24019
g23764 and n23894_not n24019 ; n24020
g23765 and n24014_not n24020_not ; n24021
g23766 and b[44]_not n24021_not ; n24022
g23767 and n23242_not quotient[6]_not ; n24023
g23768 and n23252_not n23817 ; n24024
g23769 and n23813_not n24024 ; n24025
g23770 and n23814_not n23817_not ; n24026
g23771 and n24025_not n24026_not ; n24027
g23772 and n23895 n24027_not ; n24028
g23773 and n23894_not n24028 ; n24029
g23774 and n24023_not n24029_not ; n24030
g23775 and b[43]_not n24030_not ; n24031
g23776 and n23251_not quotient[6]_not ; n24032
g23777 and n23261_not n23812 ; n24033
g23778 and n23808_not n24033 ; n24034
g23779 and n23809_not n23812_not ; n24035
g23780 and n24034_not n24035_not ; n24036
g23781 and n23895 n24036_not ; n24037
g23782 and n23894_not n24037 ; n24038
g23783 and n24032_not n24038_not ; n24039
g23784 and b[42]_not n24039_not ; n24040
g23785 and n23260_not quotient[6]_not ; n24041
g23786 and n23270_not n23807 ; n24042
g23787 and n23803_not n24042 ; n24043
g23788 and n23804_not n23807_not ; n24044
g23789 and n24043_not n24044_not ; n24045
g23790 and n23895 n24045_not ; n24046
g23791 and n23894_not n24046 ; n24047
g23792 and n24041_not n24047_not ; n24048
g23793 and b[41]_not n24048_not ; n24049
g23794 and n23269_not quotient[6]_not ; n24050
g23795 and n23279_not n23802 ; n24051
g23796 and n23798_not n24051 ; n24052
g23797 and n23799_not n23802_not ; n24053
g23798 and n24052_not n24053_not ; n24054
g23799 and n23895 n24054_not ; n24055
g23800 and n23894_not n24055 ; n24056
g23801 and n24050_not n24056_not ; n24057
g23802 and b[40]_not n24057_not ; n24058
g23803 and n23278_not quotient[6]_not ; n24059
g23804 and n23288_not n23797 ; n24060
g23805 and n23793_not n24060 ; n24061
g23806 and n23794_not n23797_not ; n24062
g23807 and n24061_not n24062_not ; n24063
g23808 and n23895 n24063_not ; n24064
g23809 and n23894_not n24064 ; n24065
g23810 and n24059_not n24065_not ; n24066
g23811 and b[39]_not n24066_not ; n24067
g23812 and n23287_not quotient[6]_not ; n24068
g23813 and n23297_not n23792 ; n24069
g23814 and n23788_not n24069 ; n24070
g23815 and n23789_not n23792_not ; n24071
g23816 and n24070_not n24071_not ; n24072
g23817 and n23895 n24072_not ; n24073
g23818 and n23894_not n24073 ; n24074
g23819 and n24068_not n24074_not ; n24075
g23820 and b[38]_not n24075_not ; n24076
g23821 and n23296_not quotient[6]_not ; n24077
g23822 and n23306_not n23787 ; n24078
g23823 and n23783_not n24078 ; n24079
g23824 and n23784_not n23787_not ; n24080
g23825 and n24079_not n24080_not ; n24081
g23826 and n23895 n24081_not ; n24082
g23827 and n23894_not n24082 ; n24083
g23828 and n24077_not n24083_not ; n24084
g23829 and b[37]_not n24084_not ; n24085
g23830 and n23305_not quotient[6]_not ; n24086
g23831 and n23315_not n23782 ; n24087
g23832 and n23778_not n24087 ; n24088
g23833 and n23779_not n23782_not ; n24089
g23834 and n24088_not n24089_not ; n24090
g23835 and n23895 n24090_not ; n24091
g23836 and n23894_not n24091 ; n24092
g23837 and n24086_not n24092_not ; n24093
g23838 and b[36]_not n24093_not ; n24094
g23839 and n23314_not quotient[6]_not ; n24095
g23840 and n23324_not n23777 ; n24096
g23841 and n23773_not n24096 ; n24097
g23842 and n23774_not n23777_not ; n24098
g23843 and n24097_not n24098_not ; n24099
g23844 and n23895 n24099_not ; n24100
g23845 and n23894_not n24100 ; n24101
g23846 and n24095_not n24101_not ; n24102
g23847 and b[35]_not n24102_not ; n24103
g23848 and n23323_not quotient[6]_not ; n24104
g23849 and n23333_not n23772 ; n24105
g23850 and n23768_not n24105 ; n24106
g23851 and n23769_not n23772_not ; n24107
g23852 and n24106_not n24107_not ; n24108
g23853 and n23895 n24108_not ; n24109
g23854 and n23894_not n24109 ; n24110
g23855 and n24104_not n24110_not ; n24111
g23856 and b[34]_not n24111_not ; n24112
g23857 and n23332_not quotient[6]_not ; n24113
g23858 and n23342_not n23767 ; n24114
g23859 and n23763_not n24114 ; n24115
g23860 and n23764_not n23767_not ; n24116
g23861 and n24115_not n24116_not ; n24117
g23862 and n23895 n24117_not ; n24118
g23863 and n23894_not n24118 ; n24119
g23864 and n24113_not n24119_not ; n24120
g23865 and b[33]_not n24120_not ; n24121
g23866 and n23341_not quotient[6]_not ; n24122
g23867 and n23351_not n23762 ; n24123
g23868 and n23758_not n24123 ; n24124
g23869 and n23759_not n23762_not ; n24125
g23870 and n24124_not n24125_not ; n24126
g23871 and n23895 n24126_not ; n24127
g23872 and n23894_not n24127 ; n24128
g23873 and n24122_not n24128_not ; n24129
g23874 and b[32]_not n24129_not ; n24130
g23875 and n23350_not quotient[6]_not ; n24131
g23876 and n23360_not n23757 ; n24132
g23877 and n23753_not n24132 ; n24133
g23878 and n23754_not n23757_not ; n24134
g23879 and n24133_not n24134_not ; n24135
g23880 and n23895 n24135_not ; n24136
g23881 and n23894_not n24136 ; n24137
g23882 and n24131_not n24137_not ; n24138
g23883 and b[31]_not n24138_not ; n24139
g23884 and n23359_not quotient[6]_not ; n24140
g23885 and n23369_not n23752 ; n24141
g23886 and n23748_not n24141 ; n24142
g23887 and n23749_not n23752_not ; n24143
g23888 and n24142_not n24143_not ; n24144
g23889 and n23895 n24144_not ; n24145
g23890 and n23894_not n24145 ; n24146
g23891 and n24140_not n24146_not ; n24147
g23892 and b[30]_not n24147_not ; n24148
g23893 and n23368_not quotient[6]_not ; n24149
g23894 and n23378_not n23747 ; n24150
g23895 and n23743_not n24150 ; n24151
g23896 and n23744_not n23747_not ; n24152
g23897 and n24151_not n24152_not ; n24153
g23898 and n23895 n24153_not ; n24154
g23899 and n23894_not n24154 ; n24155
g23900 and n24149_not n24155_not ; n24156
g23901 and b[29]_not n24156_not ; n24157
g23902 and n23377_not quotient[6]_not ; n24158
g23903 and n23387_not n23742 ; n24159
g23904 and n23738_not n24159 ; n24160
g23905 and n23739_not n23742_not ; n24161
g23906 and n24160_not n24161_not ; n24162
g23907 and n23895 n24162_not ; n24163
g23908 and n23894_not n24163 ; n24164
g23909 and n24158_not n24164_not ; n24165
g23910 and b[28]_not n24165_not ; n24166
g23911 and n23386_not quotient[6]_not ; n24167
g23912 and n23396_not n23737 ; n24168
g23913 and n23733_not n24168 ; n24169
g23914 and n23734_not n23737_not ; n24170
g23915 and n24169_not n24170_not ; n24171
g23916 and n23895 n24171_not ; n24172
g23917 and n23894_not n24172 ; n24173
g23918 and n24167_not n24173_not ; n24174
g23919 and b[27]_not n24174_not ; n24175
g23920 and n23395_not quotient[6]_not ; n24176
g23921 and n23405_not n23732 ; n24177
g23922 and n23728_not n24177 ; n24178
g23923 and n23729_not n23732_not ; n24179
g23924 and n24178_not n24179_not ; n24180
g23925 and n23895 n24180_not ; n24181
g23926 and n23894_not n24181 ; n24182
g23927 and n24176_not n24182_not ; n24183
g23928 and b[26]_not n24183_not ; n24184
g23929 and n23404_not quotient[6]_not ; n24185
g23930 and n23414_not n23727 ; n24186
g23931 and n23723_not n24186 ; n24187
g23932 and n23724_not n23727_not ; n24188
g23933 and n24187_not n24188_not ; n24189
g23934 and n23895 n24189_not ; n24190
g23935 and n23894_not n24190 ; n24191
g23936 and n24185_not n24191_not ; n24192
g23937 and b[25]_not n24192_not ; n24193
g23938 and n23413_not quotient[6]_not ; n24194
g23939 and n23423_not n23722 ; n24195
g23940 and n23718_not n24195 ; n24196
g23941 and n23719_not n23722_not ; n24197
g23942 and n24196_not n24197_not ; n24198
g23943 and n23895 n24198_not ; n24199
g23944 and n23894_not n24199 ; n24200
g23945 and n24194_not n24200_not ; n24201
g23946 and b[24]_not n24201_not ; n24202
g23947 and n23422_not quotient[6]_not ; n24203
g23948 and n23432_not n23717 ; n24204
g23949 and n23713_not n24204 ; n24205
g23950 and n23714_not n23717_not ; n24206
g23951 and n24205_not n24206_not ; n24207
g23952 and n23895 n24207_not ; n24208
g23953 and n23894_not n24208 ; n24209
g23954 and n24203_not n24209_not ; n24210
g23955 and b[23]_not n24210_not ; n24211
g23956 and n23431_not quotient[6]_not ; n24212
g23957 and n23441_not n23712 ; n24213
g23958 and n23708_not n24213 ; n24214
g23959 and n23709_not n23712_not ; n24215
g23960 and n24214_not n24215_not ; n24216
g23961 and n23895 n24216_not ; n24217
g23962 and n23894_not n24217 ; n24218
g23963 and n24212_not n24218_not ; n24219
g23964 and b[22]_not n24219_not ; n24220
g23965 and n23440_not quotient[6]_not ; n24221
g23966 and n23450_not n23707 ; n24222
g23967 and n23703_not n24222 ; n24223
g23968 and n23704_not n23707_not ; n24224
g23969 and n24223_not n24224_not ; n24225
g23970 and n23895 n24225_not ; n24226
g23971 and n23894_not n24226 ; n24227
g23972 and n24221_not n24227_not ; n24228
g23973 and b[21]_not n24228_not ; n24229
g23974 and n23449_not quotient[6]_not ; n24230
g23975 and n23459_not n23702 ; n24231
g23976 and n23698_not n24231 ; n24232
g23977 and n23699_not n23702_not ; n24233
g23978 and n24232_not n24233_not ; n24234
g23979 and n23895 n24234_not ; n24235
g23980 and n23894_not n24235 ; n24236
g23981 and n24230_not n24236_not ; n24237
g23982 and b[20]_not n24237_not ; n24238
g23983 and n23458_not quotient[6]_not ; n24239
g23984 and n23468_not n23697 ; n24240
g23985 and n23693_not n24240 ; n24241
g23986 and n23694_not n23697_not ; n24242
g23987 and n24241_not n24242_not ; n24243
g23988 and n23895 n24243_not ; n24244
g23989 and n23894_not n24244 ; n24245
g23990 and n24239_not n24245_not ; n24246
g23991 and b[19]_not n24246_not ; n24247
g23992 and n23467_not quotient[6]_not ; n24248
g23993 and n23477_not n23692 ; n24249
g23994 and n23688_not n24249 ; n24250
g23995 and n23689_not n23692_not ; n24251
g23996 and n24250_not n24251_not ; n24252
g23997 and n23895 n24252_not ; n24253
g23998 and n23894_not n24253 ; n24254
g23999 and n24248_not n24254_not ; n24255
g24000 and b[18]_not n24255_not ; n24256
g24001 and n23476_not quotient[6]_not ; n24257
g24002 and n23486_not n23687 ; n24258
g24003 and n23683_not n24258 ; n24259
g24004 and n23684_not n23687_not ; n24260
g24005 and n24259_not n24260_not ; n24261
g24006 and n23895 n24261_not ; n24262
g24007 and n23894_not n24262 ; n24263
g24008 and n24257_not n24263_not ; n24264
g24009 and b[17]_not n24264_not ; n24265
g24010 and n23485_not quotient[6]_not ; n24266
g24011 and n23495_not n23682 ; n24267
g24012 and n23678_not n24267 ; n24268
g24013 and n23679_not n23682_not ; n24269
g24014 and n24268_not n24269_not ; n24270
g24015 and n23895 n24270_not ; n24271
g24016 and n23894_not n24271 ; n24272
g24017 and n24266_not n24272_not ; n24273
g24018 and b[16]_not n24273_not ; n24274
g24019 and n23494_not quotient[6]_not ; n24275
g24020 and n23504_not n23677 ; n24276
g24021 and n23673_not n24276 ; n24277
g24022 and n23674_not n23677_not ; n24278
g24023 and n24277_not n24278_not ; n24279
g24024 and n23895 n24279_not ; n24280
g24025 and n23894_not n24280 ; n24281
g24026 and n24275_not n24281_not ; n24282
g24027 and b[15]_not n24282_not ; n24283
g24028 and n23503_not quotient[6]_not ; n24284
g24029 and n23513_not n23672 ; n24285
g24030 and n23668_not n24285 ; n24286
g24031 and n23669_not n23672_not ; n24287
g24032 and n24286_not n24287_not ; n24288
g24033 and n23895 n24288_not ; n24289
g24034 and n23894_not n24289 ; n24290
g24035 and n24284_not n24290_not ; n24291
g24036 and b[14]_not n24291_not ; n24292
g24037 and n23512_not quotient[6]_not ; n24293
g24038 and n23522_not n23667 ; n24294
g24039 and n23663_not n24294 ; n24295
g24040 and n23664_not n23667_not ; n24296
g24041 and n24295_not n24296_not ; n24297
g24042 and n23895 n24297_not ; n24298
g24043 and n23894_not n24298 ; n24299
g24044 and n24293_not n24299_not ; n24300
g24045 and b[13]_not n24300_not ; n24301
g24046 and n23521_not quotient[6]_not ; n24302
g24047 and n23531_not n23662 ; n24303
g24048 and n23658_not n24303 ; n24304
g24049 and n23659_not n23662_not ; n24305
g24050 and n24304_not n24305_not ; n24306
g24051 and n23895 n24306_not ; n24307
g24052 and n23894_not n24307 ; n24308
g24053 and n24302_not n24308_not ; n24309
g24054 and b[12]_not n24309_not ; n24310
g24055 and n23530_not quotient[6]_not ; n24311
g24056 and n23540_not n23657 ; n24312
g24057 and n23653_not n24312 ; n24313
g24058 and n23654_not n23657_not ; n24314
g24059 and n24313_not n24314_not ; n24315
g24060 and n23895 n24315_not ; n24316
g24061 and n23894_not n24316 ; n24317
g24062 and n24311_not n24317_not ; n24318
g24063 and b[11]_not n24318_not ; n24319
g24064 and n23539_not quotient[6]_not ; n24320
g24065 and n23549_not n23652 ; n24321
g24066 and n23648_not n24321 ; n24322
g24067 and n23649_not n23652_not ; n24323
g24068 and n24322_not n24323_not ; n24324
g24069 and n23895 n24324_not ; n24325
g24070 and n23894_not n24325 ; n24326
g24071 and n24320_not n24326_not ; n24327
g24072 and b[10]_not n24327_not ; n24328
g24073 and n23548_not quotient[6]_not ; n24329
g24074 and n23558_not n23647 ; n24330
g24075 and n23643_not n24330 ; n24331
g24076 and n23644_not n23647_not ; n24332
g24077 and n24331_not n24332_not ; n24333
g24078 and n23895 n24333_not ; n24334
g24079 and n23894_not n24334 ; n24335
g24080 and n24329_not n24335_not ; n24336
g24081 and b[9]_not n24336_not ; n24337
g24082 and n23557_not quotient[6]_not ; n24338
g24083 and n23567_not n23642 ; n24339
g24084 and n23638_not n24339 ; n24340
g24085 and n23639_not n23642_not ; n24341
g24086 and n24340_not n24341_not ; n24342
g24087 and n23895 n24342_not ; n24343
g24088 and n23894_not n24343 ; n24344
g24089 and n24338_not n24344_not ; n24345
g24090 and b[8]_not n24345_not ; n24346
g24091 and n23566_not quotient[6]_not ; n24347
g24092 and n23576_not n23637 ; n24348
g24093 and n23633_not n24348 ; n24349
g24094 and n23634_not n23637_not ; n24350
g24095 and n24349_not n24350_not ; n24351
g24096 and n23895 n24351_not ; n24352
g24097 and n23894_not n24352 ; n24353
g24098 and n24347_not n24353_not ; n24354
g24099 and b[7]_not n24354_not ; n24355
g24100 and n23575_not quotient[6]_not ; n24356
g24101 and n23585_not n23632 ; n24357
g24102 and n23628_not n24357 ; n24358
g24103 and n23629_not n23632_not ; n24359
g24104 and n24358_not n24359_not ; n24360
g24105 and n23895 n24360_not ; n24361
g24106 and n23894_not n24361 ; n24362
g24107 and n24356_not n24362_not ; n24363
g24108 and b[6]_not n24363_not ; n24364
g24109 and n23584_not quotient[6]_not ; n24365
g24110 and n23594_not n23627 ; n24366
g24111 and n23623_not n24366 ; n24367
g24112 and n23624_not n23627_not ; n24368
g24113 and n24367_not n24368_not ; n24369
g24114 and n23895 n24369_not ; n24370
g24115 and n23894_not n24370 ; n24371
g24116 and n24365_not n24371_not ; n24372
g24117 and b[5]_not n24372_not ; n24373
g24118 and n23593_not quotient[6]_not ; n24374
g24119 and n23602_not n23622 ; n24375
g24120 and n23618_not n24375 ; n24376
g24121 and n23619_not n23622_not ; n24377
g24122 and n24376_not n24377_not ; n24378
g24123 and n23895 n24378_not ; n24379
g24124 and n23894_not n24379 ; n24380
g24125 and n24374_not n24380_not ; n24381
g24126 and b[4]_not n24381_not ; n24382
g24127 and n23601_not quotient[6]_not ; n24383
g24128 and n23613_not n23617 ; n24384
g24129 and n23612_not n24384 ; n24385
g24130 and n23614_not n23617_not ; n24386
g24131 and n24385_not n24386_not ; n24387
g24132 and n23895 n24387_not ; n24388
g24133 and n23894_not n24388 ; n24389
g24134 and n24383_not n24389_not ; n24390
g24135 and b[3]_not n24390_not ; n24391
g24136 and n23606_not quotient[6]_not ; n24392
g24137 and n23609_not n23611 ; n24393
g24138 and n23607_not n24393 ; n24394
g24139 and n23895 n24394_not ; n24395
g24140 and n23612_not n24395 ; n24396
g24141 and n23894_not n24396 ; n24397
g24142 and n24392_not n24397_not ; n24398
g24143 and b[2]_not n24398_not ; n24399
g24144 and b[0] b[58]_not ; n24400
g24145 and n405 n24400 ; n24401
g24146 and n403 n24401 ; n24402
g24147 and n23894_not n24402 ; n24403
g24148 and a[6] n24403_not ; n24404
g24149 and n282 n23611 ; n24405
g24150 and n280 n24405 ; n24406
g24151 and n23894_not n24406 ; n24407
g24152 and n24404_not n24407_not ; n24408
g24153 and b[1] n24408_not ; n24409
g24154 and b[1]_not n24407_not ; n24410
g24155 and n24404_not n24410 ; n24411
g24156 and n24409_not n24411_not ; n24412
g24157 and a[5]_not b[0] ; n24413
g24158 and n24412_not n24413_not ; n24414
g24159 and b[1]_not n24408_not ; n24415
g24160 and n24414_not n24415_not ; n24416
g24161 and b[2] n24397_not ; n24417
g24162 and n24392_not n24417 ; n24418
g24163 and n24399_not n24418_not ; n24419
g24164 and n24416_not n24419 ; n24420
g24165 and n24399_not n24420_not ; n24421
g24166 and b[3] n24389_not ; n24422
g24167 and n24383_not n24422 ; n24423
g24168 and n24391_not n24423_not ; n24424
g24169 and n24421_not n24424 ; n24425
g24170 and n24391_not n24425_not ; n24426
g24171 and b[4] n24380_not ; n24427
g24172 and n24374_not n24427 ; n24428
g24173 and n24382_not n24428_not ; n24429
g24174 and n24426_not n24429 ; n24430
g24175 and n24382_not n24430_not ; n24431
g24176 and b[5] n24371_not ; n24432
g24177 and n24365_not n24432 ; n24433
g24178 and n24373_not n24433_not ; n24434
g24179 and n24431_not n24434 ; n24435
g24180 and n24373_not n24435_not ; n24436
g24181 and b[6] n24362_not ; n24437
g24182 and n24356_not n24437 ; n24438
g24183 and n24364_not n24438_not ; n24439
g24184 and n24436_not n24439 ; n24440
g24185 and n24364_not n24440_not ; n24441
g24186 and b[7] n24353_not ; n24442
g24187 and n24347_not n24442 ; n24443
g24188 and n24355_not n24443_not ; n24444
g24189 and n24441_not n24444 ; n24445
g24190 and n24355_not n24445_not ; n24446
g24191 and b[8] n24344_not ; n24447
g24192 and n24338_not n24447 ; n24448
g24193 and n24346_not n24448_not ; n24449
g24194 and n24446_not n24449 ; n24450
g24195 and n24346_not n24450_not ; n24451
g24196 and b[9] n24335_not ; n24452
g24197 and n24329_not n24452 ; n24453
g24198 and n24337_not n24453_not ; n24454
g24199 and n24451_not n24454 ; n24455
g24200 and n24337_not n24455_not ; n24456
g24201 and b[10] n24326_not ; n24457
g24202 and n24320_not n24457 ; n24458
g24203 and n24328_not n24458_not ; n24459
g24204 and n24456_not n24459 ; n24460
g24205 and n24328_not n24460_not ; n24461
g24206 and b[11] n24317_not ; n24462
g24207 and n24311_not n24462 ; n24463
g24208 and n24319_not n24463_not ; n24464
g24209 and n24461_not n24464 ; n24465
g24210 and n24319_not n24465_not ; n24466
g24211 and b[12] n24308_not ; n24467
g24212 and n24302_not n24467 ; n24468
g24213 and n24310_not n24468_not ; n24469
g24214 and n24466_not n24469 ; n24470
g24215 and n24310_not n24470_not ; n24471
g24216 and b[13] n24299_not ; n24472
g24217 and n24293_not n24472 ; n24473
g24218 and n24301_not n24473_not ; n24474
g24219 and n24471_not n24474 ; n24475
g24220 and n24301_not n24475_not ; n24476
g24221 and b[14] n24290_not ; n24477
g24222 and n24284_not n24477 ; n24478
g24223 and n24292_not n24478_not ; n24479
g24224 and n24476_not n24479 ; n24480
g24225 and n24292_not n24480_not ; n24481
g24226 and b[15] n24281_not ; n24482
g24227 and n24275_not n24482 ; n24483
g24228 and n24283_not n24483_not ; n24484
g24229 and n24481_not n24484 ; n24485
g24230 and n24283_not n24485_not ; n24486
g24231 and b[16] n24272_not ; n24487
g24232 and n24266_not n24487 ; n24488
g24233 and n24274_not n24488_not ; n24489
g24234 and n24486_not n24489 ; n24490
g24235 and n24274_not n24490_not ; n24491
g24236 and b[17] n24263_not ; n24492
g24237 and n24257_not n24492 ; n24493
g24238 and n24265_not n24493_not ; n24494
g24239 and n24491_not n24494 ; n24495
g24240 and n24265_not n24495_not ; n24496
g24241 and b[18] n24254_not ; n24497
g24242 and n24248_not n24497 ; n24498
g24243 and n24256_not n24498_not ; n24499
g24244 and n24496_not n24499 ; n24500
g24245 and n24256_not n24500_not ; n24501
g24246 and b[19] n24245_not ; n24502
g24247 and n24239_not n24502 ; n24503
g24248 and n24247_not n24503_not ; n24504
g24249 and n24501_not n24504 ; n24505
g24250 and n24247_not n24505_not ; n24506
g24251 and b[20] n24236_not ; n24507
g24252 and n24230_not n24507 ; n24508
g24253 and n24238_not n24508_not ; n24509
g24254 and n24506_not n24509 ; n24510
g24255 and n24238_not n24510_not ; n24511
g24256 and b[21] n24227_not ; n24512
g24257 and n24221_not n24512 ; n24513
g24258 and n24229_not n24513_not ; n24514
g24259 and n24511_not n24514 ; n24515
g24260 and n24229_not n24515_not ; n24516
g24261 and b[22] n24218_not ; n24517
g24262 and n24212_not n24517 ; n24518
g24263 and n24220_not n24518_not ; n24519
g24264 and n24516_not n24519 ; n24520
g24265 and n24220_not n24520_not ; n24521
g24266 and b[23] n24209_not ; n24522
g24267 and n24203_not n24522 ; n24523
g24268 and n24211_not n24523_not ; n24524
g24269 and n24521_not n24524 ; n24525
g24270 and n24211_not n24525_not ; n24526
g24271 and b[24] n24200_not ; n24527
g24272 and n24194_not n24527 ; n24528
g24273 and n24202_not n24528_not ; n24529
g24274 and n24526_not n24529 ; n24530
g24275 and n24202_not n24530_not ; n24531
g24276 and b[25] n24191_not ; n24532
g24277 and n24185_not n24532 ; n24533
g24278 and n24193_not n24533_not ; n24534
g24279 and n24531_not n24534 ; n24535
g24280 and n24193_not n24535_not ; n24536
g24281 and b[26] n24182_not ; n24537
g24282 and n24176_not n24537 ; n24538
g24283 and n24184_not n24538_not ; n24539
g24284 and n24536_not n24539 ; n24540
g24285 and n24184_not n24540_not ; n24541
g24286 and b[27] n24173_not ; n24542
g24287 and n24167_not n24542 ; n24543
g24288 and n24175_not n24543_not ; n24544
g24289 and n24541_not n24544 ; n24545
g24290 and n24175_not n24545_not ; n24546
g24291 and b[28] n24164_not ; n24547
g24292 and n24158_not n24547 ; n24548
g24293 and n24166_not n24548_not ; n24549
g24294 and n24546_not n24549 ; n24550
g24295 and n24166_not n24550_not ; n24551
g24296 and b[29] n24155_not ; n24552
g24297 and n24149_not n24552 ; n24553
g24298 and n24157_not n24553_not ; n24554
g24299 and n24551_not n24554 ; n24555
g24300 and n24157_not n24555_not ; n24556
g24301 and b[30] n24146_not ; n24557
g24302 and n24140_not n24557 ; n24558
g24303 and n24148_not n24558_not ; n24559
g24304 and n24556_not n24559 ; n24560
g24305 and n24148_not n24560_not ; n24561
g24306 and b[31] n24137_not ; n24562
g24307 and n24131_not n24562 ; n24563
g24308 and n24139_not n24563_not ; n24564
g24309 and n24561_not n24564 ; n24565
g24310 and n24139_not n24565_not ; n24566
g24311 and b[32] n24128_not ; n24567
g24312 and n24122_not n24567 ; n24568
g24313 and n24130_not n24568_not ; n24569
g24314 and n24566_not n24569 ; n24570
g24315 and n24130_not n24570_not ; n24571
g24316 and b[33] n24119_not ; n24572
g24317 and n24113_not n24572 ; n24573
g24318 and n24121_not n24573_not ; n24574
g24319 and n24571_not n24574 ; n24575
g24320 and n24121_not n24575_not ; n24576
g24321 and b[34] n24110_not ; n24577
g24322 and n24104_not n24577 ; n24578
g24323 and n24112_not n24578_not ; n24579
g24324 and n24576_not n24579 ; n24580
g24325 and n24112_not n24580_not ; n24581
g24326 and b[35] n24101_not ; n24582
g24327 and n24095_not n24582 ; n24583
g24328 and n24103_not n24583_not ; n24584
g24329 and n24581_not n24584 ; n24585
g24330 and n24103_not n24585_not ; n24586
g24331 and b[36] n24092_not ; n24587
g24332 and n24086_not n24587 ; n24588
g24333 and n24094_not n24588_not ; n24589
g24334 and n24586_not n24589 ; n24590
g24335 and n24094_not n24590_not ; n24591
g24336 and b[37] n24083_not ; n24592
g24337 and n24077_not n24592 ; n24593
g24338 and n24085_not n24593_not ; n24594
g24339 and n24591_not n24594 ; n24595
g24340 and n24085_not n24595_not ; n24596
g24341 and b[38] n24074_not ; n24597
g24342 and n24068_not n24597 ; n24598
g24343 and n24076_not n24598_not ; n24599
g24344 and n24596_not n24599 ; n24600
g24345 and n24076_not n24600_not ; n24601
g24346 and b[39] n24065_not ; n24602
g24347 and n24059_not n24602 ; n24603
g24348 and n24067_not n24603_not ; n24604
g24349 and n24601_not n24604 ; n24605
g24350 and n24067_not n24605_not ; n24606
g24351 and b[40] n24056_not ; n24607
g24352 and n24050_not n24607 ; n24608
g24353 and n24058_not n24608_not ; n24609
g24354 and n24606_not n24609 ; n24610
g24355 and n24058_not n24610_not ; n24611
g24356 and b[41] n24047_not ; n24612
g24357 and n24041_not n24612 ; n24613
g24358 and n24049_not n24613_not ; n24614
g24359 and n24611_not n24614 ; n24615
g24360 and n24049_not n24615_not ; n24616
g24361 and b[42] n24038_not ; n24617
g24362 and n24032_not n24617 ; n24618
g24363 and n24040_not n24618_not ; n24619
g24364 and n24616_not n24619 ; n24620
g24365 and n24040_not n24620_not ; n24621
g24366 and b[43] n24029_not ; n24622
g24367 and n24023_not n24622 ; n24623
g24368 and n24031_not n24623_not ; n24624
g24369 and n24621_not n24624 ; n24625
g24370 and n24031_not n24625_not ; n24626
g24371 and b[44] n24020_not ; n24627
g24372 and n24014_not n24627 ; n24628
g24373 and n24022_not n24628_not ; n24629
g24374 and n24626_not n24629 ; n24630
g24375 and n24022_not n24630_not ; n24631
g24376 and b[45] n24011_not ; n24632
g24377 and n24005_not n24632 ; n24633
g24378 and n24013_not n24633_not ; n24634
g24379 and n24631_not n24634 ; n24635
g24380 and n24013_not n24635_not ; n24636
g24381 and b[46] n24002_not ; n24637
g24382 and n23996_not n24637 ; n24638
g24383 and n24004_not n24638_not ; n24639
g24384 and n24636_not n24639 ; n24640
g24385 and n24004_not n24640_not ; n24641
g24386 and b[47] n23993_not ; n24642
g24387 and n23987_not n24642 ; n24643
g24388 and n23995_not n24643_not ; n24644
g24389 and n24641_not n24644 ; n24645
g24390 and n23995_not n24645_not ; n24646
g24391 and b[48] n23984_not ; n24647
g24392 and n23978_not n24647 ; n24648
g24393 and n23986_not n24648_not ; n24649
g24394 and n24646_not n24649 ; n24650
g24395 and n23986_not n24650_not ; n24651
g24396 and b[49] n23975_not ; n24652
g24397 and n23969_not n24652 ; n24653
g24398 and n23977_not n24653_not ; n24654
g24399 and n24651_not n24654 ; n24655
g24400 and n23977_not n24655_not ; n24656
g24401 and b[50] n23966_not ; n24657
g24402 and n23960_not n24657 ; n24658
g24403 and n23968_not n24658_not ; n24659
g24404 and n24656_not n24659 ; n24660
g24405 and n23968_not n24660_not ; n24661
g24406 and b[51] n23957_not ; n24662
g24407 and n23951_not n24662 ; n24663
g24408 and n23959_not n24663_not ; n24664
g24409 and n24661_not n24664 ; n24665
g24410 and n23959_not n24665_not ; n24666
g24411 and b[52] n23948_not ; n24667
g24412 and n23942_not n24667 ; n24668
g24413 and n23950_not n24668_not ; n24669
g24414 and n24666_not n24669 ; n24670
g24415 and n23950_not n24670_not ; n24671
g24416 and b[53] n23939_not ; n24672
g24417 and n23933_not n24672 ; n24673
g24418 and n23941_not n24673_not ; n24674
g24419 and n24671_not n24674 ; n24675
g24420 and n23941_not n24675_not ; n24676
g24421 and b[54] n23930_not ; n24677
g24422 and n23924_not n24677 ; n24678
g24423 and n23932_not n24678_not ; n24679
g24424 and n24676_not n24679 ; n24680
g24425 and n23932_not n24680_not ; n24681
g24426 and b[55] n23921_not ; n24682
g24427 and n23915_not n24682 ; n24683
g24428 and n23923_not n24683_not ; n24684
g24429 and n24681_not n24684 ; n24685
g24430 and n23923_not n24685_not ; n24686
g24431 and b[56] n23912_not ; n24687
g24432 and n23906_not n24687 ; n24688
g24433 and n23914_not n24688_not ; n24689
g24434 and n24686_not n24689 ; n24690
g24435 and n23914_not n24690_not ; n24691
g24436 and b[57] n23903_not ; n24692
g24437 and n23897_not n24692 ; n24693
g24438 and n23905_not n24693_not ; n24694
g24439 and n24691_not n24694 ; n24695
g24440 and n23905_not n24695_not ; n24696
g24441 and n23115_not quotient[6]_not ; n24697
g24442 and n23117_not n23892 ; n24698
g24443 and n23888_not n24698 ; n24699
g24444 and n23889_not n23892_not ; n24700
g24445 and n24699_not n24700_not ; n24701
g24446 and quotient[6] n24701_not ; n24702
g24447 and n24697_not n24702_not ; n24703
g24448 and b[58]_not n24703_not ; n24704
g24449 and b[58] n24697_not ; n24705
g24450 and n24702_not n24705 ; n24706
g24451 and n403 n405 ; n24707
g24452 and n24706_not n24707 ; n24708
g24453 and n24704_not n24708 ; n24709
g24454 and n24696_not n24709 ; n24710
g24455 and n23895 n24703_not ; n24711
g24456 and n24710_not n24711_not ; quotient[5]
g24457 and n23914_not n24694 ; n24713
g24458 and n24690_not n24713 ; n24714
g24459 and n24691_not n24694_not ; n24715
g24460 and n24714_not n24715_not ; n24716
g24461 and quotient[5] n24716_not ; n24717
g24462 and n23904_not n24711_not ; n24718
g24463 and n24710_not n24718 ; n24719
g24464 and n24717_not n24719_not ; n24720
g24465 and b[58]_not n24720_not ; n24721
g24466 and n23923_not n24689 ; n24722
g24467 and n24685_not n24722 ; n24723
g24468 and n24686_not n24689_not ; n24724
g24469 and n24723_not n24724_not ; n24725
g24470 and quotient[5] n24725_not ; n24726
g24471 and n23913_not n24711_not ; n24727
g24472 and n24710_not n24727 ; n24728
g24473 and n24726_not n24728_not ; n24729
g24474 and b[57]_not n24729_not ; n24730
g24475 and n23932_not n24684 ; n24731
g24476 and n24680_not n24731 ; n24732
g24477 and n24681_not n24684_not ; n24733
g24478 and n24732_not n24733_not ; n24734
g24479 and quotient[5] n24734_not ; n24735
g24480 and n23922_not n24711_not ; n24736
g24481 and n24710_not n24736 ; n24737
g24482 and n24735_not n24737_not ; n24738
g24483 and b[56]_not n24738_not ; n24739
g24484 and n23941_not n24679 ; n24740
g24485 and n24675_not n24740 ; n24741
g24486 and n24676_not n24679_not ; n24742
g24487 and n24741_not n24742_not ; n24743
g24488 and quotient[5] n24743_not ; n24744
g24489 and n23931_not n24711_not ; n24745
g24490 and n24710_not n24745 ; n24746
g24491 and n24744_not n24746_not ; n24747
g24492 and b[55]_not n24747_not ; n24748
g24493 and n23950_not n24674 ; n24749
g24494 and n24670_not n24749 ; n24750
g24495 and n24671_not n24674_not ; n24751
g24496 and n24750_not n24751_not ; n24752
g24497 and quotient[5] n24752_not ; n24753
g24498 and n23940_not n24711_not ; n24754
g24499 and n24710_not n24754 ; n24755
g24500 and n24753_not n24755_not ; n24756
g24501 and b[54]_not n24756_not ; n24757
g24502 and n23959_not n24669 ; n24758
g24503 and n24665_not n24758 ; n24759
g24504 and n24666_not n24669_not ; n24760
g24505 and n24759_not n24760_not ; n24761
g24506 and quotient[5] n24761_not ; n24762
g24507 and n23949_not n24711_not ; n24763
g24508 and n24710_not n24763 ; n24764
g24509 and n24762_not n24764_not ; n24765
g24510 and b[53]_not n24765_not ; n24766
g24511 and n23968_not n24664 ; n24767
g24512 and n24660_not n24767 ; n24768
g24513 and n24661_not n24664_not ; n24769
g24514 and n24768_not n24769_not ; n24770
g24515 and quotient[5] n24770_not ; n24771
g24516 and n23958_not n24711_not ; n24772
g24517 and n24710_not n24772 ; n24773
g24518 and n24771_not n24773_not ; n24774
g24519 and b[52]_not n24774_not ; n24775
g24520 and n23977_not n24659 ; n24776
g24521 and n24655_not n24776 ; n24777
g24522 and n24656_not n24659_not ; n24778
g24523 and n24777_not n24778_not ; n24779
g24524 and quotient[5] n24779_not ; n24780
g24525 and n23967_not n24711_not ; n24781
g24526 and n24710_not n24781 ; n24782
g24527 and n24780_not n24782_not ; n24783
g24528 and b[51]_not n24783_not ; n24784
g24529 and n23986_not n24654 ; n24785
g24530 and n24650_not n24785 ; n24786
g24531 and n24651_not n24654_not ; n24787
g24532 and n24786_not n24787_not ; n24788
g24533 and quotient[5] n24788_not ; n24789
g24534 and n23976_not n24711_not ; n24790
g24535 and n24710_not n24790 ; n24791
g24536 and n24789_not n24791_not ; n24792
g24537 and b[50]_not n24792_not ; n24793
g24538 and n23995_not n24649 ; n24794
g24539 and n24645_not n24794 ; n24795
g24540 and n24646_not n24649_not ; n24796
g24541 and n24795_not n24796_not ; n24797
g24542 and quotient[5] n24797_not ; n24798
g24543 and n23985_not n24711_not ; n24799
g24544 and n24710_not n24799 ; n24800
g24545 and n24798_not n24800_not ; n24801
g24546 and b[49]_not n24801_not ; n24802
g24547 and n24004_not n24644 ; n24803
g24548 and n24640_not n24803 ; n24804
g24549 and n24641_not n24644_not ; n24805
g24550 and n24804_not n24805_not ; n24806
g24551 and quotient[5] n24806_not ; n24807
g24552 and n23994_not n24711_not ; n24808
g24553 and n24710_not n24808 ; n24809
g24554 and n24807_not n24809_not ; n24810
g24555 and b[48]_not n24810_not ; n24811
g24556 and n24013_not n24639 ; n24812
g24557 and n24635_not n24812 ; n24813
g24558 and n24636_not n24639_not ; n24814
g24559 and n24813_not n24814_not ; n24815
g24560 and quotient[5] n24815_not ; n24816
g24561 and n24003_not n24711_not ; n24817
g24562 and n24710_not n24817 ; n24818
g24563 and n24816_not n24818_not ; n24819
g24564 and b[47]_not n24819_not ; n24820
g24565 and n24022_not n24634 ; n24821
g24566 and n24630_not n24821 ; n24822
g24567 and n24631_not n24634_not ; n24823
g24568 and n24822_not n24823_not ; n24824
g24569 and quotient[5] n24824_not ; n24825
g24570 and n24012_not n24711_not ; n24826
g24571 and n24710_not n24826 ; n24827
g24572 and n24825_not n24827_not ; n24828
g24573 and b[46]_not n24828_not ; n24829
g24574 and n24031_not n24629 ; n24830
g24575 and n24625_not n24830 ; n24831
g24576 and n24626_not n24629_not ; n24832
g24577 and n24831_not n24832_not ; n24833
g24578 and quotient[5] n24833_not ; n24834
g24579 and n24021_not n24711_not ; n24835
g24580 and n24710_not n24835 ; n24836
g24581 and n24834_not n24836_not ; n24837
g24582 and b[45]_not n24837_not ; n24838
g24583 and n24040_not n24624 ; n24839
g24584 and n24620_not n24839 ; n24840
g24585 and n24621_not n24624_not ; n24841
g24586 and n24840_not n24841_not ; n24842
g24587 and quotient[5] n24842_not ; n24843
g24588 and n24030_not n24711_not ; n24844
g24589 and n24710_not n24844 ; n24845
g24590 and n24843_not n24845_not ; n24846
g24591 and b[44]_not n24846_not ; n24847
g24592 and n24049_not n24619 ; n24848
g24593 and n24615_not n24848 ; n24849
g24594 and n24616_not n24619_not ; n24850
g24595 and n24849_not n24850_not ; n24851
g24596 and quotient[5] n24851_not ; n24852
g24597 and n24039_not n24711_not ; n24853
g24598 and n24710_not n24853 ; n24854
g24599 and n24852_not n24854_not ; n24855
g24600 and b[43]_not n24855_not ; n24856
g24601 and n24058_not n24614 ; n24857
g24602 and n24610_not n24857 ; n24858
g24603 and n24611_not n24614_not ; n24859
g24604 and n24858_not n24859_not ; n24860
g24605 and quotient[5] n24860_not ; n24861
g24606 and n24048_not n24711_not ; n24862
g24607 and n24710_not n24862 ; n24863
g24608 and n24861_not n24863_not ; n24864
g24609 and b[42]_not n24864_not ; n24865
g24610 and n24067_not n24609 ; n24866
g24611 and n24605_not n24866 ; n24867
g24612 and n24606_not n24609_not ; n24868
g24613 and n24867_not n24868_not ; n24869
g24614 and quotient[5] n24869_not ; n24870
g24615 and n24057_not n24711_not ; n24871
g24616 and n24710_not n24871 ; n24872
g24617 and n24870_not n24872_not ; n24873
g24618 and b[41]_not n24873_not ; n24874
g24619 and n24076_not n24604 ; n24875
g24620 and n24600_not n24875 ; n24876
g24621 and n24601_not n24604_not ; n24877
g24622 and n24876_not n24877_not ; n24878
g24623 and quotient[5] n24878_not ; n24879
g24624 and n24066_not n24711_not ; n24880
g24625 and n24710_not n24880 ; n24881
g24626 and n24879_not n24881_not ; n24882
g24627 and b[40]_not n24882_not ; n24883
g24628 and n24085_not n24599 ; n24884
g24629 and n24595_not n24884 ; n24885
g24630 and n24596_not n24599_not ; n24886
g24631 and n24885_not n24886_not ; n24887
g24632 and quotient[5] n24887_not ; n24888
g24633 and n24075_not n24711_not ; n24889
g24634 and n24710_not n24889 ; n24890
g24635 and n24888_not n24890_not ; n24891
g24636 and b[39]_not n24891_not ; n24892
g24637 and n24094_not n24594 ; n24893
g24638 and n24590_not n24893 ; n24894
g24639 and n24591_not n24594_not ; n24895
g24640 and n24894_not n24895_not ; n24896
g24641 and quotient[5] n24896_not ; n24897
g24642 and n24084_not n24711_not ; n24898
g24643 and n24710_not n24898 ; n24899
g24644 and n24897_not n24899_not ; n24900
g24645 and b[38]_not n24900_not ; n24901
g24646 and n24103_not n24589 ; n24902
g24647 and n24585_not n24902 ; n24903
g24648 and n24586_not n24589_not ; n24904
g24649 and n24903_not n24904_not ; n24905
g24650 and quotient[5] n24905_not ; n24906
g24651 and n24093_not n24711_not ; n24907
g24652 and n24710_not n24907 ; n24908
g24653 and n24906_not n24908_not ; n24909
g24654 and b[37]_not n24909_not ; n24910
g24655 and n24112_not n24584 ; n24911
g24656 and n24580_not n24911 ; n24912
g24657 and n24581_not n24584_not ; n24913
g24658 and n24912_not n24913_not ; n24914
g24659 and quotient[5] n24914_not ; n24915
g24660 and n24102_not n24711_not ; n24916
g24661 and n24710_not n24916 ; n24917
g24662 and n24915_not n24917_not ; n24918
g24663 and b[36]_not n24918_not ; n24919
g24664 and n24121_not n24579 ; n24920
g24665 and n24575_not n24920 ; n24921
g24666 and n24576_not n24579_not ; n24922
g24667 and n24921_not n24922_not ; n24923
g24668 and quotient[5] n24923_not ; n24924
g24669 and n24111_not n24711_not ; n24925
g24670 and n24710_not n24925 ; n24926
g24671 and n24924_not n24926_not ; n24927
g24672 and b[35]_not n24927_not ; n24928
g24673 and n24130_not n24574 ; n24929
g24674 and n24570_not n24929 ; n24930
g24675 and n24571_not n24574_not ; n24931
g24676 and n24930_not n24931_not ; n24932
g24677 and quotient[5] n24932_not ; n24933
g24678 and n24120_not n24711_not ; n24934
g24679 and n24710_not n24934 ; n24935
g24680 and n24933_not n24935_not ; n24936
g24681 and b[34]_not n24936_not ; n24937
g24682 and n24139_not n24569 ; n24938
g24683 and n24565_not n24938 ; n24939
g24684 and n24566_not n24569_not ; n24940
g24685 and n24939_not n24940_not ; n24941
g24686 and quotient[5] n24941_not ; n24942
g24687 and n24129_not n24711_not ; n24943
g24688 and n24710_not n24943 ; n24944
g24689 and n24942_not n24944_not ; n24945
g24690 and b[33]_not n24945_not ; n24946
g24691 and n24148_not n24564 ; n24947
g24692 and n24560_not n24947 ; n24948
g24693 and n24561_not n24564_not ; n24949
g24694 and n24948_not n24949_not ; n24950
g24695 and quotient[5] n24950_not ; n24951
g24696 and n24138_not n24711_not ; n24952
g24697 and n24710_not n24952 ; n24953
g24698 and n24951_not n24953_not ; n24954
g24699 and b[32]_not n24954_not ; n24955
g24700 and n24157_not n24559 ; n24956
g24701 and n24555_not n24956 ; n24957
g24702 and n24556_not n24559_not ; n24958
g24703 and n24957_not n24958_not ; n24959
g24704 and quotient[5] n24959_not ; n24960
g24705 and n24147_not n24711_not ; n24961
g24706 and n24710_not n24961 ; n24962
g24707 and n24960_not n24962_not ; n24963
g24708 and b[31]_not n24963_not ; n24964
g24709 and n24166_not n24554 ; n24965
g24710 and n24550_not n24965 ; n24966
g24711 and n24551_not n24554_not ; n24967
g24712 and n24966_not n24967_not ; n24968
g24713 and quotient[5] n24968_not ; n24969
g24714 and n24156_not n24711_not ; n24970
g24715 and n24710_not n24970 ; n24971
g24716 and n24969_not n24971_not ; n24972
g24717 and b[30]_not n24972_not ; n24973
g24718 and n24175_not n24549 ; n24974
g24719 and n24545_not n24974 ; n24975
g24720 and n24546_not n24549_not ; n24976
g24721 and n24975_not n24976_not ; n24977
g24722 and quotient[5] n24977_not ; n24978
g24723 and n24165_not n24711_not ; n24979
g24724 and n24710_not n24979 ; n24980
g24725 and n24978_not n24980_not ; n24981
g24726 and b[29]_not n24981_not ; n24982
g24727 and n24184_not n24544 ; n24983
g24728 and n24540_not n24983 ; n24984
g24729 and n24541_not n24544_not ; n24985
g24730 and n24984_not n24985_not ; n24986
g24731 and quotient[5] n24986_not ; n24987
g24732 and n24174_not n24711_not ; n24988
g24733 and n24710_not n24988 ; n24989
g24734 and n24987_not n24989_not ; n24990
g24735 and b[28]_not n24990_not ; n24991
g24736 and n24193_not n24539 ; n24992
g24737 and n24535_not n24992 ; n24993
g24738 and n24536_not n24539_not ; n24994
g24739 and n24993_not n24994_not ; n24995
g24740 and quotient[5] n24995_not ; n24996
g24741 and n24183_not n24711_not ; n24997
g24742 and n24710_not n24997 ; n24998
g24743 and n24996_not n24998_not ; n24999
g24744 and b[27]_not n24999_not ; n25000
g24745 and n24202_not n24534 ; n25001
g24746 and n24530_not n25001 ; n25002
g24747 and n24531_not n24534_not ; n25003
g24748 and n25002_not n25003_not ; n25004
g24749 and quotient[5] n25004_not ; n25005
g24750 and n24192_not n24711_not ; n25006
g24751 and n24710_not n25006 ; n25007
g24752 and n25005_not n25007_not ; n25008
g24753 and b[26]_not n25008_not ; n25009
g24754 and n24211_not n24529 ; n25010
g24755 and n24525_not n25010 ; n25011
g24756 and n24526_not n24529_not ; n25012
g24757 and n25011_not n25012_not ; n25013
g24758 and quotient[5] n25013_not ; n25014
g24759 and n24201_not n24711_not ; n25015
g24760 and n24710_not n25015 ; n25016
g24761 and n25014_not n25016_not ; n25017
g24762 and b[25]_not n25017_not ; n25018
g24763 and n24220_not n24524 ; n25019
g24764 and n24520_not n25019 ; n25020
g24765 and n24521_not n24524_not ; n25021
g24766 and n25020_not n25021_not ; n25022
g24767 and quotient[5] n25022_not ; n25023
g24768 and n24210_not n24711_not ; n25024
g24769 and n24710_not n25024 ; n25025
g24770 and n25023_not n25025_not ; n25026
g24771 and b[24]_not n25026_not ; n25027
g24772 and n24229_not n24519 ; n25028
g24773 and n24515_not n25028 ; n25029
g24774 and n24516_not n24519_not ; n25030
g24775 and n25029_not n25030_not ; n25031
g24776 and quotient[5] n25031_not ; n25032
g24777 and n24219_not n24711_not ; n25033
g24778 and n24710_not n25033 ; n25034
g24779 and n25032_not n25034_not ; n25035
g24780 and b[23]_not n25035_not ; n25036
g24781 and n24238_not n24514 ; n25037
g24782 and n24510_not n25037 ; n25038
g24783 and n24511_not n24514_not ; n25039
g24784 and n25038_not n25039_not ; n25040
g24785 and quotient[5] n25040_not ; n25041
g24786 and n24228_not n24711_not ; n25042
g24787 and n24710_not n25042 ; n25043
g24788 and n25041_not n25043_not ; n25044
g24789 and b[22]_not n25044_not ; n25045
g24790 and n24247_not n24509 ; n25046
g24791 and n24505_not n25046 ; n25047
g24792 and n24506_not n24509_not ; n25048
g24793 and n25047_not n25048_not ; n25049
g24794 and quotient[5] n25049_not ; n25050
g24795 and n24237_not n24711_not ; n25051
g24796 and n24710_not n25051 ; n25052
g24797 and n25050_not n25052_not ; n25053
g24798 and b[21]_not n25053_not ; n25054
g24799 and n24256_not n24504 ; n25055
g24800 and n24500_not n25055 ; n25056
g24801 and n24501_not n24504_not ; n25057
g24802 and n25056_not n25057_not ; n25058
g24803 and quotient[5] n25058_not ; n25059
g24804 and n24246_not n24711_not ; n25060
g24805 and n24710_not n25060 ; n25061
g24806 and n25059_not n25061_not ; n25062
g24807 and b[20]_not n25062_not ; n25063
g24808 and n24265_not n24499 ; n25064
g24809 and n24495_not n25064 ; n25065
g24810 and n24496_not n24499_not ; n25066
g24811 and n25065_not n25066_not ; n25067
g24812 and quotient[5] n25067_not ; n25068
g24813 and n24255_not n24711_not ; n25069
g24814 and n24710_not n25069 ; n25070
g24815 and n25068_not n25070_not ; n25071
g24816 and b[19]_not n25071_not ; n25072
g24817 and n24274_not n24494 ; n25073
g24818 and n24490_not n25073 ; n25074
g24819 and n24491_not n24494_not ; n25075
g24820 and n25074_not n25075_not ; n25076
g24821 and quotient[5] n25076_not ; n25077
g24822 and n24264_not n24711_not ; n25078
g24823 and n24710_not n25078 ; n25079
g24824 and n25077_not n25079_not ; n25080
g24825 and b[18]_not n25080_not ; n25081
g24826 and n24283_not n24489 ; n25082
g24827 and n24485_not n25082 ; n25083
g24828 and n24486_not n24489_not ; n25084
g24829 and n25083_not n25084_not ; n25085
g24830 and quotient[5] n25085_not ; n25086
g24831 and n24273_not n24711_not ; n25087
g24832 and n24710_not n25087 ; n25088
g24833 and n25086_not n25088_not ; n25089
g24834 and b[17]_not n25089_not ; n25090
g24835 and n24292_not n24484 ; n25091
g24836 and n24480_not n25091 ; n25092
g24837 and n24481_not n24484_not ; n25093
g24838 and n25092_not n25093_not ; n25094
g24839 and quotient[5] n25094_not ; n25095
g24840 and n24282_not n24711_not ; n25096
g24841 and n24710_not n25096 ; n25097
g24842 and n25095_not n25097_not ; n25098
g24843 and b[16]_not n25098_not ; n25099
g24844 and n24301_not n24479 ; n25100
g24845 and n24475_not n25100 ; n25101
g24846 and n24476_not n24479_not ; n25102
g24847 and n25101_not n25102_not ; n25103
g24848 and quotient[5] n25103_not ; n25104
g24849 and n24291_not n24711_not ; n25105
g24850 and n24710_not n25105 ; n25106
g24851 and n25104_not n25106_not ; n25107
g24852 and b[15]_not n25107_not ; n25108
g24853 and n24310_not n24474 ; n25109
g24854 and n24470_not n25109 ; n25110
g24855 and n24471_not n24474_not ; n25111
g24856 and n25110_not n25111_not ; n25112
g24857 and quotient[5] n25112_not ; n25113
g24858 and n24300_not n24711_not ; n25114
g24859 and n24710_not n25114 ; n25115
g24860 and n25113_not n25115_not ; n25116
g24861 and b[14]_not n25116_not ; n25117
g24862 and n24319_not n24469 ; n25118
g24863 and n24465_not n25118 ; n25119
g24864 and n24466_not n24469_not ; n25120
g24865 and n25119_not n25120_not ; n25121
g24866 and quotient[5] n25121_not ; n25122
g24867 and n24309_not n24711_not ; n25123
g24868 and n24710_not n25123 ; n25124
g24869 and n25122_not n25124_not ; n25125
g24870 and b[13]_not n25125_not ; n25126
g24871 and n24328_not n24464 ; n25127
g24872 and n24460_not n25127 ; n25128
g24873 and n24461_not n24464_not ; n25129
g24874 and n25128_not n25129_not ; n25130
g24875 and quotient[5] n25130_not ; n25131
g24876 and n24318_not n24711_not ; n25132
g24877 and n24710_not n25132 ; n25133
g24878 and n25131_not n25133_not ; n25134
g24879 and b[12]_not n25134_not ; n25135
g24880 and n24337_not n24459 ; n25136
g24881 and n24455_not n25136 ; n25137
g24882 and n24456_not n24459_not ; n25138
g24883 and n25137_not n25138_not ; n25139
g24884 and quotient[5] n25139_not ; n25140
g24885 and n24327_not n24711_not ; n25141
g24886 and n24710_not n25141 ; n25142
g24887 and n25140_not n25142_not ; n25143
g24888 and b[11]_not n25143_not ; n25144
g24889 and n24346_not n24454 ; n25145
g24890 and n24450_not n25145 ; n25146
g24891 and n24451_not n24454_not ; n25147
g24892 and n25146_not n25147_not ; n25148
g24893 and quotient[5] n25148_not ; n25149
g24894 and n24336_not n24711_not ; n25150
g24895 and n24710_not n25150 ; n25151
g24896 and n25149_not n25151_not ; n25152
g24897 and b[10]_not n25152_not ; n25153
g24898 and n24355_not n24449 ; n25154
g24899 and n24445_not n25154 ; n25155
g24900 and n24446_not n24449_not ; n25156
g24901 and n25155_not n25156_not ; n25157
g24902 and quotient[5] n25157_not ; n25158
g24903 and n24345_not n24711_not ; n25159
g24904 and n24710_not n25159 ; n25160
g24905 and n25158_not n25160_not ; n25161
g24906 and b[9]_not n25161_not ; n25162
g24907 and n24364_not n24444 ; n25163
g24908 and n24440_not n25163 ; n25164
g24909 and n24441_not n24444_not ; n25165
g24910 and n25164_not n25165_not ; n25166
g24911 and quotient[5] n25166_not ; n25167
g24912 and n24354_not n24711_not ; n25168
g24913 and n24710_not n25168 ; n25169
g24914 and n25167_not n25169_not ; n25170
g24915 and b[8]_not n25170_not ; n25171
g24916 and n24373_not n24439 ; n25172
g24917 and n24435_not n25172 ; n25173
g24918 and n24436_not n24439_not ; n25174
g24919 and n25173_not n25174_not ; n25175
g24920 and quotient[5] n25175_not ; n25176
g24921 and n24363_not n24711_not ; n25177
g24922 and n24710_not n25177 ; n25178
g24923 and n25176_not n25178_not ; n25179
g24924 and b[7]_not n25179_not ; n25180
g24925 and n24382_not n24434 ; n25181
g24926 and n24430_not n25181 ; n25182
g24927 and n24431_not n24434_not ; n25183
g24928 and n25182_not n25183_not ; n25184
g24929 and quotient[5] n25184_not ; n25185
g24930 and n24372_not n24711_not ; n25186
g24931 and n24710_not n25186 ; n25187
g24932 and n25185_not n25187_not ; n25188
g24933 and b[6]_not n25188_not ; n25189
g24934 and n24391_not n24429 ; n25190
g24935 and n24425_not n25190 ; n25191
g24936 and n24426_not n24429_not ; n25192
g24937 and n25191_not n25192_not ; n25193
g24938 and quotient[5] n25193_not ; n25194
g24939 and n24381_not n24711_not ; n25195
g24940 and n24710_not n25195 ; n25196
g24941 and n25194_not n25196_not ; n25197
g24942 and b[5]_not n25197_not ; n25198
g24943 and n24399_not n24424 ; n25199
g24944 and n24420_not n25199 ; n25200
g24945 and n24421_not n24424_not ; n25201
g24946 and n25200_not n25201_not ; n25202
g24947 and quotient[5] n25202_not ; n25203
g24948 and n24390_not n24711_not ; n25204
g24949 and n24710_not n25204 ; n25205
g24950 and n25203_not n25205_not ; n25206
g24951 and b[4]_not n25206_not ; n25207
g24952 and n24415_not n24419 ; n25208
g24953 and n24414_not n25208 ; n25209
g24954 and n24416_not n24419_not ; n25210
g24955 and n25209_not n25210_not ; n25211
g24956 and quotient[5] n25211_not ; n25212
g24957 and n24398_not n24711_not ; n25213
g24958 and n24710_not n25213 ; n25214
g24959 and n25212_not n25214_not ; n25215
g24960 and b[3]_not n25215_not ; n25216
g24961 and n24411_not n24413 ; n25217
g24962 and n24409_not n25217 ; n25218
g24963 and n24414_not n25218_not ; n25219
g24964 and quotient[5] n25219 ; n25220
g24965 and n24408_not n24711_not ; n25221
g24966 and n24710_not n25221 ; n25222
g24967 and n25220_not n25222_not ; n25223
g24968 and b[2]_not n25223_not ; n25224
g24969 and b[0] quotient[5] ; n25225
g24970 and a[5] n25225_not ; n25226
g24971 and n24413 quotient[5] ; n25227
g24972 and n25226_not n25227_not ; n25228
g24973 and b[1] n25228_not ; n25229
g24974 and b[1]_not n25227_not ; n25230
g24975 and n25226_not n25230 ; n25231
g24976 and n25229_not n25231_not ; n25232
g24977 and a[4]_not b[0] ; n25233
g24978 and n25232_not n25233_not ; n25234
g24979 and b[1]_not n25228_not ; n25235
g24980 and n25234_not n25235_not ; n25236
g24981 and b[2] n25222_not ; n25237
g24982 and n25220_not n25237 ; n25238
g24983 and n25224_not n25238_not ; n25239
g24984 and n25236_not n25239 ; n25240
g24985 and n25224_not n25240_not ; n25241
g24986 and b[3] n25214_not ; n25242
g24987 and n25212_not n25242 ; n25243
g24988 and n25216_not n25243_not ; n25244
g24989 and n25241_not n25244 ; n25245
g24990 and n25216_not n25245_not ; n25246
g24991 and b[4] n25205_not ; n25247
g24992 and n25203_not n25247 ; n25248
g24993 and n25207_not n25248_not ; n25249
g24994 and n25246_not n25249 ; n25250
g24995 and n25207_not n25250_not ; n25251
g24996 and b[5] n25196_not ; n25252
g24997 and n25194_not n25252 ; n25253
g24998 and n25198_not n25253_not ; n25254
g24999 and n25251_not n25254 ; n25255
g25000 and n25198_not n25255_not ; n25256
g25001 and b[6] n25187_not ; n25257
g25002 and n25185_not n25257 ; n25258
g25003 and n25189_not n25258_not ; n25259
g25004 and n25256_not n25259 ; n25260
g25005 and n25189_not n25260_not ; n25261
g25006 and b[7] n25178_not ; n25262
g25007 and n25176_not n25262 ; n25263
g25008 and n25180_not n25263_not ; n25264
g25009 and n25261_not n25264 ; n25265
g25010 and n25180_not n25265_not ; n25266
g25011 and b[8] n25169_not ; n25267
g25012 and n25167_not n25267 ; n25268
g25013 and n25171_not n25268_not ; n25269
g25014 and n25266_not n25269 ; n25270
g25015 and n25171_not n25270_not ; n25271
g25016 and b[9] n25160_not ; n25272
g25017 and n25158_not n25272 ; n25273
g25018 and n25162_not n25273_not ; n25274
g25019 and n25271_not n25274 ; n25275
g25020 and n25162_not n25275_not ; n25276
g25021 and b[10] n25151_not ; n25277
g25022 and n25149_not n25277 ; n25278
g25023 and n25153_not n25278_not ; n25279
g25024 and n25276_not n25279 ; n25280
g25025 and n25153_not n25280_not ; n25281
g25026 and b[11] n25142_not ; n25282
g25027 and n25140_not n25282 ; n25283
g25028 and n25144_not n25283_not ; n25284
g25029 and n25281_not n25284 ; n25285
g25030 and n25144_not n25285_not ; n25286
g25031 and b[12] n25133_not ; n25287
g25032 and n25131_not n25287 ; n25288
g25033 and n25135_not n25288_not ; n25289
g25034 and n25286_not n25289 ; n25290
g25035 and n25135_not n25290_not ; n25291
g25036 and b[13] n25124_not ; n25292
g25037 and n25122_not n25292 ; n25293
g25038 and n25126_not n25293_not ; n25294
g25039 and n25291_not n25294 ; n25295
g25040 and n25126_not n25295_not ; n25296
g25041 and b[14] n25115_not ; n25297
g25042 and n25113_not n25297 ; n25298
g25043 and n25117_not n25298_not ; n25299
g25044 and n25296_not n25299 ; n25300
g25045 and n25117_not n25300_not ; n25301
g25046 and b[15] n25106_not ; n25302
g25047 and n25104_not n25302 ; n25303
g25048 and n25108_not n25303_not ; n25304
g25049 and n25301_not n25304 ; n25305
g25050 and n25108_not n25305_not ; n25306
g25051 and b[16] n25097_not ; n25307
g25052 and n25095_not n25307 ; n25308
g25053 and n25099_not n25308_not ; n25309
g25054 and n25306_not n25309 ; n25310
g25055 and n25099_not n25310_not ; n25311
g25056 and b[17] n25088_not ; n25312
g25057 and n25086_not n25312 ; n25313
g25058 and n25090_not n25313_not ; n25314
g25059 and n25311_not n25314 ; n25315
g25060 and n25090_not n25315_not ; n25316
g25061 and b[18] n25079_not ; n25317
g25062 and n25077_not n25317 ; n25318
g25063 and n25081_not n25318_not ; n25319
g25064 and n25316_not n25319 ; n25320
g25065 and n25081_not n25320_not ; n25321
g25066 and b[19] n25070_not ; n25322
g25067 and n25068_not n25322 ; n25323
g25068 and n25072_not n25323_not ; n25324
g25069 and n25321_not n25324 ; n25325
g25070 and n25072_not n25325_not ; n25326
g25071 and b[20] n25061_not ; n25327
g25072 and n25059_not n25327 ; n25328
g25073 and n25063_not n25328_not ; n25329
g25074 and n25326_not n25329 ; n25330
g25075 and n25063_not n25330_not ; n25331
g25076 and b[21] n25052_not ; n25332
g25077 and n25050_not n25332 ; n25333
g25078 and n25054_not n25333_not ; n25334
g25079 and n25331_not n25334 ; n25335
g25080 and n25054_not n25335_not ; n25336
g25081 and b[22] n25043_not ; n25337
g25082 and n25041_not n25337 ; n25338
g25083 and n25045_not n25338_not ; n25339
g25084 and n25336_not n25339 ; n25340
g25085 and n25045_not n25340_not ; n25341
g25086 and b[23] n25034_not ; n25342
g25087 and n25032_not n25342 ; n25343
g25088 and n25036_not n25343_not ; n25344
g25089 and n25341_not n25344 ; n25345
g25090 and n25036_not n25345_not ; n25346
g25091 and b[24] n25025_not ; n25347
g25092 and n25023_not n25347 ; n25348
g25093 and n25027_not n25348_not ; n25349
g25094 and n25346_not n25349 ; n25350
g25095 and n25027_not n25350_not ; n25351
g25096 and b[25] n25016_not ; n25352
g25097 and n25014_not n25352 ; n25353
g25098 and n25018_not n25353_not ; n25354
g25099 and n25351_not n25354 ; n25355
g25100 and n25018_not n25355_not ; n25356
g25101 and b[26] n25007_not ; n25357
g25102 and n25005_not n25357 ; n25358
g25103 and n25009_not n25358_not ; n25359
g25104 and n25356_not n25359 ; n25360
g25105 and n25009_not n25360_not ; n25361
g25106 and b[27] n24998_not ; n25362
g25107 and n24996_not n25362 ; n25363
g25108 and n25000_not n25363_not ; n25364
g25109 and n25361_not n25364 ; n25365
g25110 and n25000_not n25365_not ; n25366
g25111 and b[28] n24989_not ; n25367
g25112 and n24987_not n25367 ; n25368
g25113 and n24991_not n25368_not ; n25369
g25114 and n25366_not n25369 ; n25370
g25115 and n24991_not n25370_not ; n25371
g25116 and b[29] n24980_not ; n25372
g25117 and n24978_not n25372 ; n25373
g25118 and n24982_not n25373_not ; n25374
g25119 and n25371_not n25374 ; n25375
g25120 and n24982_not n25375_not ; n25376
g25121 and b[30] n24971_not ; n25377
g25122 and n24969_not n25377 ; n25378
g25123 and n24973_not n25378_not ; n25379
g25124 and n25376_not n25379 ; n25380
g25125 and n24973_not n25380_not ; n25381
g25126 and b[31] n24962_not ; n25382
g25127 and n24960_not n25382 ; n25383
g25128 and n24964_not n25383_not ; n25384
g25129 and n25381_not n25384 ; n25385
g25130 and n24964_not n25385_not ; n25386
g25131 and b[32] n24953_not ; n25387
g25132 and n24951_not n25387 ; n25388
g25133 and n24955_not n25388_not ; n25389
g25134 and n25386_not n25389 ; n25390
g25135 and n24955_not n25390_not ; n25391
g25136 and b[33] n24944_not ; n25392
g25137 and n24942_not n25392 ; n25393
g25138 and n24946_not n25393_not ; n25394
g25139 and n25391_not n25394 ; n25395
g25140 and n24946_not n25395_not ; n25396
g25141 and b[34] n24935_not ; n25397
g25142 and n24933_not n25397 ; n25398
g25143 and n24937_not n25398_not ; n25399
g25144 and n25396_not n25399 ; n25400
g25145 and n24937_not n25400_not ; n25401
g25146 and b[35] n24926_not ; n25402
g25147 and n24924_not n25402 ; n25403
g25148 and n24928_not n25403_not ; n25404
g25149 and n25401_not n25404 ; n25405
g25150 and n24928_not n25405_not ; n25406
g25151 and b[36] n24917_not ; n25407
g25152 and n24915_not n25407 ; n25408
g25153 and n24919_not n25408_not ; n25409
g25154 and n25406_not n25409 ; n25410
g25155 and n24919_not n25410_not ; n25411
g25156 and b[37] n24908_not ; n25412
g25157 and n24906_not n25412 ; n25413
g25158 and n24910_not n25413_not ; n25414
g25159 and n25411_not n25414 ; n25415
g25160 and n24910_not n25415_not ; n25416
g25161 and b[38] n24899_not ; n25417
g25162 and n24897_not n25417 ; n25418
g25163 and n24901_not n25418_not ; n25419
g25164 and n25416_not n25419 ; n25420
g25165 and n24901_not n25420_not ; n25421
g25166 and b[39] n24890_not ; n25422
g25167 and n24888_not n25422 ; n25423
g25168 and n24892_not n25423_not ; n25424
g25169 and n25421_not n25424 ; n25425
g25170 and n24892_not n25425_not ; n25426
g25171 and b[40] n24881_not ; n25427
g25172 and n24879_not n25427 ; n25428
g25173 and n24883_not n25428_not ; n25429
g25174 and n25426_not n25429 ; n25430
g25175 and n24883_not n25430_not ; n25431
g25176 and b[41] n24872_not ; n25432
g25177 and n24870_not n25432 ; n25433
g25178 and n24874_not n25433_not ; n25434
g25179 and n25431_not n25434 ; n25435
g25180 and n24874_not n25435_not ; n25436
g25181 and b[42] n24863_not ; n25437
g25182 and n24861_not n25437 ; n25438
g25183 and n24865_not n25438_not ; n25439
g25184 and n25436_not n25439 ; n25440
g25185 and n24865_not n25440_not ; n25441
g25186 and b[43] n24854_not ; n25442
g25187 and n24852_not n25442 ; n25443
g25188 and n24856_not n25443_not ; n25444
g25189 and n25441_not n25444 ; n25445
g25190 and n24856_not n25445_not ; n25446
g25191 and b[44] n24845_not ; n25447
g25192 and n24843_not n25447 ; n25448
g25193 and n24847_not n25448_not ; n25449
g25194 and n25446_not n25449 ; n25450
g25195 and n24847_not n25450_not ; n25451
g25196 and b[45] n24836_not ; n25452
g25197 and n24834_not n25452 ; n25453
g25198 and n24838_not n25453_not ; n25454
g25199 and n25451_not n25454 ; n25455
g25200 and n24838_not n25455_not ; n25456
g25201 and b[46] n24827_not ; n25457
g25202 and n24825_not n25457 ; n25458
g25203 and n24829_not n25458_not ; n25459
g25204 and n25456_not n25459 ; n25460
g25205 and n24829_not n25460_not ; n25461
g25206 and b[47] n24818_not ; n25462
g25207 and n24816_not n25462 ; n25463
g25208 and n24820_not n25463_not ; n25464
g25209 and n25461_not n25464 ; n25465
g25210 and n24820_not n25465_not ; n25466
g25211 and b[48] n24809_not ; n25467
g25212 and n24807_not n25467 ; n25468
g25213 and n24811_not n25468_not ; n25469
g25214 and n25466_not n25469 ; n25470
g25215 and n24811_not n25470_not ; n25471
g25216 and b[49] n24800_not ; n25472
g25217 and n24798_not n25472 ; n25473
g25218 and n24802_not n25473_not ; n25474
g25219 and n25471_not n25474 ; n25475
g25220 and n24802_not n25475_not ; n25476
g25221 and b[50] n24791_not ; n25477
g25222 and n24789_not n25477 ; n25478
g25223 and n24793_not n25478_not ; n25479
g25224 and n25476_not n25479 ; n25480
g25225 and n24793_not n25480_not ; n25481
g25226 and b[51] n24782_not ; n25482
g25227 and n24780_not n25482 ; n25483
g25228 and n24784_not n25483_not ; n25484
g25229 and n25481_not n25484 ; n25485
g25230 and n24784_not n25485_not ; n25486
g25231 and b[52] n24773_not ; n25487
g25232 and n24771_not n25487 ; n25488
g25233 and n24775_not n25488_not ; n25489
g25234 and n25486_not n25489 ; n25490
g25235 and n24775_not n25490_not ; n25491
g25236 and b[53] n24764_not ; n25492
g25237 and n24762_not n25492 ; n25493
g25238 and n24766_not n25493_not ; n25494
g25239 and n25491_not n25494 ; n25495
g25240 and n24766_not n25495_not ; n25496
g25241 and b[54] n24755_not ; n25497
g25242 and n24753_not n25497 ; n25498
g25243 and n24757_not n25498_not ; n25499
g25244 and n25496_not n25499 ; n25500
g25245 and n24757_not n25500_not ; n25501
g25246 and b[55] n24746_not ; n25502
g25247 and n24744_not n25502 ; n25503
g25248 and n24748_not n25503_not ; n25504
g25249 and n25501_not n25504 ; n25505
g25250 and n24748_not n25505_not ; n25506
g25251 and b[56] n24737_not ; n25507
g25252 and n24735_not n25507 ; n25508
g25253 and n24739_not n25508_not ; n25509
g25254 and n25506_not n25509 ; n25510
g25255 and n24739_not n25510_not ; n25511
g25256 and b[57] n24728_not ; n25512
g25257 and n24726_not n25512 ; n25513
g25258 and n24730_not n25513_not ; n25514
g25259 and n25511_not n25514 ; n25515
g25260 and n24730_not n25515_not ; n25516
g25261 and b[58] n24719_not ; n25517
g25262 and n24717_not n25517 ; n25518
g25263 and n24721_not n25518_not ; n25519
g25264 and n25516_not n25519 ; n25520
g25265 and n24721_not n25520_not ; n25521
g25266 and n23905_not n24706_not ; n25522
g25267 and n24704_not n25522 ; n25523
g25268 and n24695_not n25523 ; n25524
g25269 and n24704_not n24706_not ; n25525
g25270 and n24696_not n25525_not ; n25526
g25271 and n25524_not n25526_not ; n25527
g25272 and quotient[5] n25527_not ; n25528
g25273 and n24703_not n24711_not ; n25529
g25274 and n24710_not n25529 ; n25530
g25275 and n25528_not n25530_not ; n25531
g25276 and b[59]_not n25531_not ; n25532
g25277 and b[59] n25530_not ; n25533
g25278 and n25528_not n25533 ; n25534
g25279 and n280 n25534_not ; n25535
g25280 and n25532_not n25535 ; n25536
g25281 and n25521_not n25536 ; n25537
g25282 and n24707 n25531_not ; n25538
g25283 and n25537_not n25538_not ; quotient[4]
g25284 and n24730_not n25519 ; n25540
g25285 and n25515_not n25540 ; n25541
g25286 and n25516_not n25519_not ; n25542
g25287 and n25541_not n25542_not ; n25543
g25288 and quotient[4] n25543_not ; n25544
g25289 and n24720_not n25538_not ; n25545
g25290 and n25537_not n25545 ; n25546
g25291 and n25544_not n25546_not ; n25547
g25292 and b[59]_not n25547_not ; n25548
g25293 and n24739_not n25514 ; n25549
g25294 and n25510_not n25549 ; n25550
g25295 and n25511_not n25514_not ; n25551
g25296 and n25550_not n25551_not ; n25552
g25297 and quotient[4] n25552_not ; n25553
g25298 and n24729_not n25538_not ; n25554
g25299 and n25537_not n25554 ; n25555
g25300 and n25553_not n25555_not ; n25556
g25301 and b[58]_not n25556_not ; n25557
g25302 and n24748_not n25509 ; n25558
g25303 and n25505_not n25558 ; n25559
g25304 and n25506_not n25509_not ; n25560
g25305 and n25559_not n25560_not ; n25561
g25306 and quotient[4] n25561_not ; n25562
g25307 and n24738_not n25538_not ; n25563
g25308 and n25537_not n25563 ; n25564
g25309 and n25562_not n25564_not ; n25565
g25310 and b[57]_not n25565_not ; n25566
g25311 and n24757_not n25504 ; n25567
g25312 and n25500_not n25567 ; n25568
g25313 and n25501_not n25504_not ; n25569
g25314 and n25568_not n25569_not ; n25570
g25315 and quotient[4] n25570_not ; n25571
g25316 and n24747_not n25538_not ; n25572
g25317 and n25537_not n25572 ; n25573
g25318 and n25571_not n25573_not ; n25574
g25319 and b[56]_not n25574_not ; n25575
g25320 and n24766_not n25499 ; n25576
g25321 and n25495_not n25576 ; n25577
g25322 and n25496_not n25499_not ; n25578
g25323 and n25577_not n25578_not ; n25579
g25324 and quotient[4] n25579_not ; n25580
g25325 and n24756_not n25538_not ; n25581
g25326 and n25537_not n25581 ; n25582
g25327 and n25580_not n25582_not ; n25583
g25328 and b[55]_not n25583_not ; n25584
g25329 and n24775_not n25494 ; n25585
g25330 and n25490_not n25585 ; n25586
g25331 and n25491_not n25494_not ; n25587
g25332 and n25586_not n25587_not ; n25588
g25333 and quotient[4] n25588_not ; n25589
g25334 and n24765_not n25538_not ; n25590
g25335 and n25537_not n25590 ; n25591
g25336 and n25589_not n25591_not ; n25592
g25337 and b[54]_not n25592_not ; n25593
g25338 and n24784_not n25489 ; n25594
g25339 and n25485_not n25594 ; n25595
g25340 and n25486_not n25489_not ; n25596
g25341 and n25595_not n25596_not ; n25597
g25342 and quotient[4] n25597_not ; n25598
g25343 and n24774_not n25538_not ; n25599
g25344 and n25537_not n25599 ; n25600
g25345 and n25598_not n25600_not ; n25601
g25346 and b[53]_not n25601_not ; n25602
g25347 and n24793_not n25484 ; n25603
g25348 and n25480_not n25603 ; n25604
g25349 and n25481_not n25484_not ; n25605
g25350 and n25604_not n25605_not ; n25606
g25351 and quotient[4] n25606_not ; n25607
g25352 and n24783_not n25538_not ; n25608
g25353 and n25537_not n25608 ; n25609
g25354 and n25607_not n25609_not ; n25610
g25355 and b[52]_not n25610_not ; n25611
g25356 and n24802_not n25479 ; n25612
g25357 and n25475_not n25612 ; n25613
g25358 and n25476_not n25479_not ; n25614
g25359 and n25613_not n25614_not ; n25615
g25360 and quotient[4] n25615_not ; n25616
g25361 and n24792_not n25538_not ; n25617
g25362 and n25537_not n25617 ; n25618
g25363 and n25616_not n25618_not ; n25619
g25364 and b[51]_not n25619_not ; n25620
g25365 and n24811_not n25474 ; n25621
g25366 and n25470_not n25621 ; n25622
g25367 and n25471_not n25474_not ; n25623
g25368 and n25622_not n25623_not ; n25624
g25369 and quotient[4] n25624_not ; n25625
g25370 and n24801_not n25538_not ; n25626
g25371 and n25537_not n25626 ; n25627
g25372 and n25625_not n25627_not ; n25628
g25373 and b[50]_not n25628_not ; n25629
g25374 and n24820_not n25469 ; n25630
g25375 and n25465_not n25630 ; n25631
g25376 and n25466_not n25469_not ; n25632
g25377 and n25631_not n25632_not ; n25633
g25378 and quotient[4] n25633_not ; n25634
g25379 and n24810_not n25538_not ; n25635
g25380 and n25537_not n25635 ; n25636
g25381 and n25634_not n25636_not ; n25637
g25382 and b[49]_not n25637_not ; n25638
g25383 and n24829_not n25464 ; n25639
g25384 and n25460_not n25639 ; n25640
g25385 and n25461_not n25464_not ; n25641
g25386 and n25640_not n25641_not ; n25642
g25387 and quotient[4] n25642_not ; n25643
g25388 and n24819_not n25538_not ; n25644
g25389 and n25537_not n25644 ; n25645
g25390 and n25643_not n25645_not ; n25646
g25391 and b[48]_not n25646_not ; n25647
g25392 and n24838_not n25459 ; n25648
g25393 and n25455_not n25648 ; n25649
g25394 and n25456_not n25459_not ; n25650
g25395 and n25649_not n25650_not ; n25651
g25396 and quotient[4] n25651_not ; n25652
g25397 and n24828_not n25538_not ; n25653
g25398 and n25537_not n25653 ; n25654
g25399 and n25652_not n25654_not ; n25655
g25400 and b[47]_not n25655_not ; n25656
g25401 and n24847_not n25454 ; n25657
g25402 and n25450_not n25657 ; n25658
g25403 and n25451_not n25454_not ; n25659
g25404 and n25658_not n25659_not ; n25660
g25405 and quotient[4] n25660_not ; n25661
g25406 and n24837_not n25538_not ; n25662
g25407 and n25537_not n25662 ; n25663
g25408 and n25661_not n25663_not ; n25664
g25409 and b[46]_not n25664_not ; n25665
g25410 and n24856_not n25449 ; n25666
g25411 and n25445_not n25666 ; n25667
g25412 and n25446_not n25449_not ; n25668
g25413 and n25667_not n25668_not ; n25669
g25414 and quotient[4] n25669_not ; n25670
g25415 and n24846_not n25538_not ; n25671
g25416 and n25537_not n25671 ; n25672
g25417 and n25670_not n25672_not ; n25673
g25418 and b[45]_not n25673_not ; n25674
g25419 and n24865_not n25444 ; n25675
g25420 and n25440_not n25675 ; n25676
g25421 and n25441_not n25444_not ; n25677
g25422 and n25676_not n25677_not ; n25678
g25423 and quotient[4] n25678_not ; n25679
g25424 and n24855_not n25538_not ; n25680
g25425 and n25537_not n25680 ; n25681
g25426 and n25679_not n25681_not ; n25682
g25427 and b[44]_not n25682_not ; n25683
g25428 and n24874_not n25439 ; n25684
g25429 and n25435_not n25684 ; n25685
g25430 and n25436_not n25439_not ; n25686
g25431 and n25685_not n25686_not ; n25687
g25432 and quotient[4] n25687_not ; n25688
g25433 and n24864_not n25538_not ; n25689
g25434 and n25537_not n25689 ; n25690
g25435 and n25688_not n25690_not ; n25691
g25436 and b[43]_not n25691_not ; n25692
g25437 and n24883_not n25434 ; n25693
g25438 and n25430_not n25693 ; n25694
g25439 and n25431_not n25434_not ; n25695
g25440 and n25694_not n25695_not ; n25696
g25441 and quotient[4] n25696_not ; n25697
g25442 and n24873_not n25538_not ; n25698
g25443 and n25537_not n25698 ; n25699
g25444 and n25697_not n25699_not ; n25700
g25445 and b[42]_not n25700_not ; n25701
g25446 and n24892_not n25429 ; n25702
g25447 and n25425_not n25702 ; n25703
g25448 and n25426_not n25429_not ; n25704
g25449 and n25703_not n25704_not ; n25705
g25450 and quotient[4] n25705_not ; n25706
g25451 and n24882_not n25538_not ; n25707
g25452 and n25537_not n25707 ; n25708
g25453 and n25706_not n25708_not ; n25709
g25454 and b[41]_not n25709_not ; n25710
g25455 and n24901_not n25424 ; n25711
g25456 and n25420_not n25711 ; n25712
g25457 and n25421_not n25424_not ; n25713
g25458 and n25712_not n25713_not ; n25714
g25459 and quotient[4] n25714_not ; n25715
g25460 and n24891_not n25538_not ; n25716
g25461 and n25537_not n25716 ; n25717
g25462 and n25715_not n25717_not ; n25718
g25463 and b[40]_not n25718_not ; n25719
g25464 and n24910_not n25419 ; n25720
g25465 and n25415_not n25720 ; n25721
g25466 and n25416_not n25419_not ; n25722
g25467 and n25721_not n25722_not ; n25723
g25468 and quotient[4] n25723_not ; n25724
g25469 and n24900_not n25538_not ; n25725
g25470 and n25537_not n25725 ; n25726
g25471 and n25724_not n25726_not ; n25727
g25472 and b[39]_not n25727_not ; n25728
g25473 and n24919_not n25414 ; n25729
g25474 and n25410_not n25729 ; n25730
g25475 and n25411_not n25414_not ; n25731
g25476 and n25730_not n25731_not ; n25732
g25477 and quotient[4] n25732_not ; n25733
g25478 and n24909_not n25538_not ; n25734
g25479 and n25537_not n25734 ; n25735
g25480 and n25733_not n25735_not ; n25736
g25481 and b[38]_not n25736_not ; n25737
g25482 and n24928_not n25409 ; n25738
g25483 and n25405_not n25738 ; n25739
g25484 and n25406_not n25409_not ; n25740
g25485 and n25739_not n25740_not ; n25741
g25486 and quotient[4] n25741_not ; n25742
g25487 and n24918_not n25538_not ; n25743
g25488 and n25537_not n25743 ; n25744
g25489 and n25742_not n25744_not ; n25745
g25490 and b[37]_not n25745_not ; n25746
g25491 and n24937_not n25404 ; n25747
g25492 and n25400_not n25747 ; n25748
g25493 and n25401_not n25404_not ; n25749
g25494 and n25748_not n25749_not ; n25750
g25495 and quotient[4] n25750_not ; n25751
g25496 and n24927_not n25538_not ; n25752
g25497 and n25537_not n25752 ; n25753
g25498 and n25751_not n25753_not ; n25754
g25499 and b[36]_not n25754_not ; n25755
g25500 and n24946_not n25399 ; n25756
g25501 and n25395_not n25756 ; n25757
g25502 and n25396_not n25399_not ; n25758
g25503 and n25757_not n25758_not ; n25759
g25504 and quotient[4] n25759_not ; n25760
g25505 and n24936_not n25538_not ; n25761
g25506 and n25537_not n25761 ; n25762
g25507 and n25760_not n25762_not ; n25763
g25508 and b[35]_not n25763_not ; n25764
g25509 and n24955_not n25394 ; n25765
g25510 and n25390_not n25765 ; n25766
g25511 and n25391_not n25394_not ; n25767
g25512 and n25766_not n25767_not ; n25768
g25513 and quotient[4] n25768_not ; n25769
g25514 and n24945_not n25538_not ; n25770
g25515 and n25537_not n25770 ; n25771
g25516 and n25769_not n25771_not ; n25772
g25517 and b[34]_not n25772_not ; n25773
g25518 and n24964_not n25389 ; n25774
g25519 and n25385_not n25774 ; n25775
g25520 and n25386_not n25389_not ; n25776
g25521 and n25775_not n25776_not ; n25777
g25522 and quotient[4] n25777_not ; n25778
g25523 and n24954_not n25538_not ; n25779
g25524 and n25537_not n25779 ; n25780
g25525 and n25778_not n25780_not ; n25781
g25526 and b[33]_not n25781_not ; n25782
g25527 and n24973_not n25384 ; n25783
g25528 and n25380_not n25783 ; n25784
g25529 and n25381_not n25384_not ; n25785
g25530 and n25784_not n25785_not ; n25786
g25531 and quotient[4] n25786_not ; n25787
g25532 and n24963_not n25538_not ; n25788
g25533 and n25537_not n25788 ; n25789
g25534 and n25787_not n25789_not ; n25790
g25535 and b[32]_not n25790_not ; n25791
g25536 and n24982_not n25379 ; n25792
g25537 and n25375_not n25792 ; n25793
g25538 and n25376_not n25379_not ; n25794
g25539 and n25793_not n25794_not ; n25795
g25540 and quotient[4] n25795_not ; n25796
g25541 and n24972_not n25538_not ; n25797
g25542 and n25537_not n25797 ; n25798
g25543 and n25796_not n25798_not ; n25799
g25544 and b[31]_not n25799_not ; n25800
g25545 and n24991_not n25374 ; n25801
g25546 and n25370_not n25801 ; n25802
g25547 and n25371_not n25374_not ; n25803
g25548 and n25802_not n25803_not ; n25804
g25549 and quotient[4] n25804_not ; n25805
g25550 and n24981_not n25538_not ; n25806
g25551 and n25537_not n25806 ; n25807
g25552 and n25805_not n25807_not ; n25808
g25553 and b[30]_not n25808_not ; n25809
g25554 and n25000_not n25369 ; n25810
g25555 and n25365_not n25810 ; n25811
g25556 and n25366_not n25369_not ; n25812
g25557 and n25811_not n25812_not ; n25813
g25558 and quotient[4] n25813_not ; n25814
g25559 and n24990_not n25538_not ; n25815
g25560 and n25537_not n25815 ; n25816
g25561 and n25814_not n25816_not ; n25817
g25562 and b[29]_not n25817_not ; n25818
g25563 and n25009_not n25364 ; n25819
g25564 and n25360_not n25819 ; n25820
g25565 and n25361_not n25364_not ; n25821
g25566 and n25820_not n25821_not ; n25822
g25567 and quotient[4] n25822_not ; n25823
g25568 and n24999_not n25538_not ; n25824
g25569 and n25537_not n25824 ; n25825
g25570 and n25823_not n25825_not ; n25826
g25571 and b[28]_not n25826_not ; n25827
g25572 and n25018_not n25359 ; n25828
g25573 and n25355_not n25828 ; n25829
g25574 and n25356_not n25359_not ; n25830
g25575 and n25829_not n25830_not ; n25831
g25576 and quotient[4] n25831_not ; n25832
g25577 and n25008_not n25538_not ; n25833
g25578 and n25537_not n25833 ; n25834
g25579 and n25832_not n25834_not ; n25835
g25580 and b[27]_not n25835_not ; n25836
g25581 and n25027_not n25354 ; n25837
g25582 and n25350_not n25837 ; n25838
g25583 and n25351_not n25354_not ; n25839
g25584 and n25838_not n25839_not ; n25840
g25585 and quotient[4] n25840_not ; n25841
g25586 and n25017_not n25538_not ; n25842
g25587 and n25537_not n25842 ; n25843
g25588 and n25841_not n25843_not ; n25844
g25589 and b[26]_not n25844_not ; n25845
g25590 and n25036_not n25349 ; n25846
g25591 and n25345_not n25846 ; n25847
g25592 and n25346_not n25349_not ; n25848
g25593 and n25847_not n25848_not ; n25849
g25594 and quotient[4] n25849_not ; n25850
g25595 and n25026_not n25538_not ; n25851
g25596 and n25537_not n25851 ; n25852
g25597 and n25850_not n25852_not ; n25853
g25598 and b[25]_not n25853_not ; n25854
g25599 and n25045_not n25344 ; n25855
g25600 and n25340_not n25855 ; n25856
g25601 and n25341_not n25344_not ; n25857
g25602 and n25856_not n25857_not ; n25858
g25603 and quotient[4] n25858_not ; n25859
g25604 and n25035_not n25538_not ; n25860
g25605 and n25537_not n25860 ; n25861
g25606 and n25859_not n25861_not ; n25862
g25607 and b[24]_not n25862_not ; n25863
g25608 and n25054_not n25339 ; n25864
g25609 and n25335_not n25864 ; n25865
g25610 and n25336_not n25339_not ; n25866
g25611 and n25865_not n25866_not ; n25867
g25612 and quotient[4] n25867_not ; n25868
g25613 and n25044_not n25538_not ; n25869
g25614 and n25537_not n25869 ; n25870
g25615 and n25868_not n25870_not ; n25871
g25616 and b[23]_not n25871_not ; n25872
g25617 and n25063_not n25334 ; n25873
g25618 and n25330_not n25873 ; n25874
g25619 and n25331_not n25334_not ; n25875
g25620 and n25874_not n25875_not ; n25876
g25621 and quotient[4] n25876_not ; n25877
g25622 and n25053_not n25538_not ; n25878
g25623 and n25537_not n25878 ; n25879
g25624 and n25877_not n25879_not ; n25880
g25625 and b[22]_not n25880_not ; n25881
g25626 and n25072_not n25329 ; n25882
g25627 and n25325_not n25882 ; n25883
g25628 and n25326_not n25329_not ; n25884
g25629 and n25883_not n25884_not ; n25885
g25630 and quotient[4] n25885_not ; n25886
g25631 and n25062_not n25538_not ; n25887
g25632 and n25537_not n25887 ; n25888
g25633 and n25886_not n25888_not ; n25889
g25634 and b[21]_not n25889_not ; n25890
g25635 and n25081_not n25324 ; n25891
g25636 and n25320_not n25891 ; n25892
g25637 and n25321_not n25324_not ; n25893
g25638 and n25892_not n25893_not ; n25894
g25639 and quotient[4] n25894_not ; n25895
g25640 and n25071_not n25538_not ; n25896
g25641 and n25537_not n25896 ; n25897
g25642 and n25895_not n25897_not ; n25898
g25643 and b[20]_not n25898_not ; n25899
g25644 and n25090_not n25319 ; n25900
g25645 and n25315_not n25900 ; n25901
g25646 and n25316_not n25319_not ; n25902
g25647 and n25901_not n25902_not ; n25903
g25648 and quotient[4] n25903_not ; n25904
g25649 and n25080_not n25538_not ; n25905
g25650 and n25537_not n25905 ; n25906
g25651 and n25904_not n25906_not ; n25907
g25652 and b[19]_not n25907_not ; n25908
g25653 and n25099_not n25314 ; n25909
g25654 and n25310_not n25909 ; n25910
g25655 and n25311_not n25314_not ; n25911
g25656 and n25910_not n25911_not ; n25912
g25657 and quotient[4] n25912_not ; n25913
g25658 and n25089_not n25538_not ; n25914
g25659 and n25537_not n25914 ; n25915
g25660 and n25913_not n25915_not ; n25916
g25661 and b[18]_not n25916_not ; n25917
g25662 and n25108_not n25309 ; n25918
g25663 and n25305_not n25918 ; n25919
g25664 and n25306_not n25309_not ; n25920
g25665 and n25919_not n25920_not ; n25921
g25666 and quotient[4] n25921_not ; n25922
g25667 and n25098_not n25538_not ; n25923
g25668 and n25537_not n25923 ; n25924
g25669 and n25922_not n25924_not ; n25925
g25670 and b[17]_not n25925_not ; n25926
g25671 and n25117_not n25304 ; n25927
g25672 and n25300_not n25927 ; n25928
g25673 and n25301_not n25304_not ; n25929
g25674 and n25928_not n25929_not ; n25930
g25675 and quotient[4] n25930_not ; n25931
g25676 and n25107_not n25538_not ; n25932
g25677 and n25537_not n25932 ; n25933
g25678 and n25931_not n25933_not ; n25934
g25679 and b[16]_not n25934_not ; n25935
g25680 and n25126_not n25299 ; n25936
g25681 and n25295_not n25936 ; n25937
g25682 and n25296_not n25299_not ; n25938
g25683 and n25937_not n25938_not ; n25939
g25684 and quotient[4] n25939_not ; n25940
g25685 and n25116_not n25538_not ; n25941
g25686 and n25537_not n25941 ; n25942
g25687 and n25940_not n25942_not ; n25943
g25688 and b[15]_not n25943_not ; n25944
g25689 and n25135_not n25294 ; n25945
g25690 and n25290_not n25945 ; n25946
g25691 and n25291_not n25294_not ; n25947
g25692 and n25946_not n25947_not ; n25948
g25693 and quotient[4] n25948_not ; n25949
g25694 and n25125_not n25538_not ; n25950
g25695 and n25537_not n25950 ; n25951
g25696 and n25949_not n25951_not ; n25952
g25697 and b[14]_not n25952_not ; n25953
g25698 and n25144_not n25289 ; n25954
g25699 and n25285_not n25954 ; n25955
g25700 and n25286_not n25289_not ; n25956
g25701 and n25955_not n25956_not ; n25957
g25702 and quotient[4] n25957_not ; n25958
g25703 and n25134_not n25538_not ; n25959
g25704 and n25537_not n25959 ; n25960
g25705 and n25958_not n25960_not ; n25961
g25706 and b[13]_not n25961_not ; n25962
g25707 and n25153_not n25284 ; n25963
g25708 and n25280_not n25963 ; n25964
g25709 and n25281_not n25284_not ; n25965
g25710 and n25964_not n25965_not ; n25966
g25711 and quotient[4] n25966_not ; n25967
g25712 and n25143_not n25538_not ; n25968
g25713 and n25537_not n25968 ; n25969
g25714 and n25967_not n25969_not ; n25970
g25715 and b[12]_not n25970_not ; n25971
g25716 and n25162_not n25279 ; n25972
g25717 and n25275_not n25972 ; n25973
g25718 and n25276_not n25279_not ; n25974
g25719 and n25973_not n25974_not ; n25975
g25720 and quotient[4] n25975_not ; n25976
g25721 and n25152_not n25538_not ; n25977
g25722 and n25537_not n25977 ; n25978
g25723 and n25976_not n25978_not ; n25979
g25724 and b[11]_not n25979_not ; n25980
g25725 and n25171_not n25274 ; n25981
g25726 and n25270_not n25981 ; n25982
g25727 and n25271_not n25274_not ; n25983
g25728 and n25982_not n25983_not ; n25984
g25729 and quotient[4] n25984_not ; n25985
g25730 and n25161_not n25538_not ; n25986
g25731 and n25537_not n25986 ; n25987
g25732 and n25985_not n25987_not ; n25988
g25733 and b[10]_not n25988_not ; n25989
g25734 and n25180_not n25269 ; n25990
g25735 and n25265_not n25990 ; n25991
g25736 and n25266_not n25269_not ; n25992
g25737 and n25991_not n25992_not ; n25993
g25738 and quotient[4] n25993_not ; n25994
g25739 and n25170_not n25538_not ; n25995
g25740 and n25537_not n25995 ; n25996
g25741 and n25994_not n25996_not ; n25997
g25742 and b[9]_not n25997_not ; n25998
g25743 and n25189_not n25264 ; n25999
g25744 and n25260_not n25999 ; n26000
g25745 and n25261_not n25264_not ; n26001
g25746 and n26000_not n26001_not ; n26002
g25747 and quotient[4] n26002_not ; n26003
g25748 and n25179_not n25538_not ; n26004
g25749 and n25537_not n26004 ; n26005
g25750 and n26003_not n26005_not ; n26006
g25751 and b[8]_not n26006_not ; n26007
g25752 and n25198_not n25259 ; n26008
g25753 and n25255_not n26008 ; n26009
g25754 and n25256_not n25259_not ; n26010
g25755 and n26009_not n26010_not ; n26011
g25756 and quotient[4] n26011_not ; n26012
g25757 and n25188_not n25538_not ; n26013
g25758 and n25537_not n26013 ; n26014
g25759 and n26012_not n26014_not ; n26015
g25760 and b[7]_not n26015_not ; n26016
g25761 and n25207_not n25254 ; n26017
g25762 and n25250_not n26017 ; n26018
g25763 and n25251_not n25254_not ; n26019
g25764 and n26018_not n26019_not ; n26020
g25765 and quotient[4] n26020_not ; n26021
g25766 and n25197_not n25538_not ; n26022
g25767 and n25537_not n26022 ; n26023
g25768 and n26021_not n26023_not ; n26024
g25769 and b[6]_not n26024_not ; n26025
g25770 and n25216_not n25249 ; n26026
g25771 and n25245_not n26026 ; n26027
g25772 and n25246_not n25249_not ; n26028
g25773 and n26027_not n26028_not ; n26029
g25774 and quotient[4] n26029_not ; n26030
g25775 and n25206_not n25538_not ; n26031
g25776 and n25537_not n26031 ; n26032
g25777 and n26030_not n26032_not ; n26033
g25778 and b[5]_not n26033_not ; n26034
g25779 and n25224_not n25244 ; n26035
g25780 and n25240_not n26035 ; n26036
g25781 and n25241_not n25244_not ; n26037
g25782 and n26036_not n26037_not ; n26038
g25783 and quotient[4] n26038_not ; n26039
g25784 and n25215_not n25538_not ; n26040
g25785 and n25537_not n26040 ; n26041
g25786 and n26039_not n26041_not ; n26042
g25787 and b[4]_not n26042_not ; n26043
g25788 and n25235_not n25239 ; n26044
g25789 and n25234_not n26044 ; n26045
g25790 and n25236_not n25239_not ; n26046
g25791 and n26045_not n26046_not ; n26047
g25792 and quotient[4] n26047_not ; n26048
g25793 and n25223_not n25538_not ; n26049
g25794 and n25537_not n26049 ; n26050
g25795 and n26048_not n26050_not ; n26051
g25796 and b[3]_not n26051_not ; n26052
g25797 and n25231_not n25233 ; n26053
g25798 and n25229_not n26053 ; n26054
g25799 and n25234_not n26054_not ; n26055
g25800 and quotient[4] n26055 ; n26056
g25801 and n25228_not n25538_not ; n26057
g25802 and n25537_not n26057 ; n26058
g25803 and n26056_not n26058_not ; n26059
g25804 and b[2]_not n26059_not ; n26060
g25805 and b[0] quotient[4] ; n26061
g25806 and a[4] n26061_not ; n26062
g25807 and n25233 quotient[4] ; n26063
g25808 and n26062_not n26063_not ; n26064
g25809 and b[1] n26064_not ; n26065
g25810 and b[1]_not n26063_not ; n26066
g25811 and n26062_not n26066 ; n26067
g25812 and n26065_not n26067_not ; n26068
g25813 and a[3]_not b[0] ; n26069
g25814 and n26068_not n26069_not ; n26070
g25815 and b[1]_not n26064_not ; n26071
g25816 and n26070_not n26071_not ; n26072
g25817 and b[2] n26058_not ; n26073
g25818 and n26056_not n26073 ; n26074
g25819 and n26060_not n26074_not ; n26075
g25820 and n26072_not n26075 ; n26076
g25821 and n26060_not n26076_not ; n26077
g25822 and b[3] n26050_not ; n26078
g25823 and n26048_not n26078 ; n26079
g25824 and n26052_not n26079_not ; n26080
g25825 and n26077_not n26080 ; n26081
g25826 and n26052_not n26081_not ; n26082
g25827 and b[4] n26041_not ; n26083
g25828 and n26039_not n26083 ; n26084
g25829 and n26043_not n26084_not ; n26085
g25830 and n26082_not n26085 ; n26086
g25831 and n26043_not n26086_not ; n26087
g25832 and b[5] n26032_not ; n26088
g25833 and n26030_not n26088 ; n26089
g25834 and n26034_not n26089_not ; n26090
g25835 and n26087_not n26090 ; n26091
g25836 and n26034_not n26091_not ; n26092
g25837 and b[6] n26023_not ; n26093
g25838 and n26021_not n26093 ; n26094
g25839 and n26025_not n26094_not ; n26095
g25840 and n26092_not n26095 ; n26096
g25841 and n26025_not n26096_not ; n26097
g25842 and b[7] n26014_not ; n26098
g25843 and n26012_not n26098 ; n26099
g25844 and n26016_not n26099_not ; n26100
g25845 and n26097_not n26100 ; n26101
g25846 and n26016_not n26101_not ; n26102
g25847 and b[8] n26005_not ; n26103
g25848 and n26003_not n26103 ; n26104
g25849 and n26007_not n26104_not ; n26105
g25850 and n26102_not n26105 ; n26106
g25851 and n26007_not n26106_not ; n26107
g25852 and b[9] n25996_not ; n26108
g25853 and n25994_not n26108 ; n26109
g25854 and n25998_not n26109_not ; n26110
g25855 and n26107_not n26110 ; n26111
g25856 and n25998_not n26111_not ; n26112
g25857 and b[10] n25987_not ; n26113
g25858 and n25985_not n26113 ; n26114
g25859 and n25989_not n26114_not ; n26115
g25860 and n26112_not n26115 ; n26116
g25861 and n25989_not n26116_not ; n26117
g25862 and b[11] n25978_not ; n26118
g25863 and n25976_not n26118 ; n26119
g25864 and n25980_not n26119_not ; n26120
g25865 and n26117_not n26120 ; n26121
g25866 and n25980_not n26121_not ; n26122
g25867 and b[12] n25969_not ; n26123
g25868 and n25967_not n26123 ; n26124
g25869 and n25971_not n26124_not ; n26125
g25870 and n26122_not n26125 ; n26126
g25871 and n25971_not n26126_not ; n26127
g25872 and b[13] n25960_not ; n26128
g25873 and n25958_not n26128 ; n26129
g25874 and n25962_not n26129_not ; n26130
g25875 and n26127_not n26130 ; n26131
g25876 and n25962_not n26131_not ; n26132
g25877 and b[14] n25951_not ; n26133
g25878 and n25949_not n26133 ; n26134
g25879 and n25953_not n26134_not ; n26135
g25880 and n26132_not n26135 ; n26136
g25881 and n25953_not n26136_not ; n26137
g25882 and b[15] n25942_not ; n26138
g25883 and n25940_not n26138 ; n26139
g25884 and n25944_not n26139_not ; n26140
g25885 and n26137_not n26140 ; n26141
g25886 and n25944_not n26141_not ; n26142
g25887 and b[16] n25933_not ; n26143
g25888 and n25931_not n26143 ; n26144
g25889 and n25935_not n26144_not ; n26145
g25890 and n26142_not n26145 ; n26146
g25891 and n25935_not n26146_not ; n26147
g25892 and b[17] n25924_not ; n26148
g25893 and n25922_not n26148 ; n26149
g25894 and n25926_not n26149_not ; n26150
g25895 and n26147_not n26150 ; n26151
g25896 and n25926_not n26151_not ; n26152
g25897 and b[18] n25915_not ; n26153
g25898 and n25913_not n26153 ; n26154
g25899 and n25917_not n26154_not ; n26155
g25900 and n26152_not n26155 ; n26156
g25901 and n25917_not n26156_not ; n26157
g25902 and b[19] n25906_not ; n26158
g25903 and n25904_not n26158 ; n26159
g25904 and n25908_not n26159_not ; n26160
g25905 and n26157_not n26160 ; n26161
g25906 and n25908_not n26161_not ; n26162
g25907 and b[20] n25897_not ; n26163
g25908 and n25895_not n26163 ; n26164
g25909 and n25899_not n26164_not ; n26165
g25910 and n26162_not n26165 ; n26166
g25911 and n25899_not n26166_not ; n26167
g25912 and b[21] n25888_not ; n26168
g25913 and n25886_not n26168 ; n26169
g25914 and n25890_not n26169_not ; n26170
g25915 and n26167_not n26170 ; n26171
g25916 and n25890_not n26171_not ; n26172
g25917 and b[22] n25879_not ; n26173
g25918 and n25877_not n26173 ; n26174
g25919 and n25881_not n26174_not ; n26175
g25920 and n26172_not n26175 ; n26176
g25921 and n25881_not n26176_not ; n26177
g25922 and b[23] n25870_not ; n26178
g25923 and n25868_not n26178 ; n26179
g25924 and n25872_not n26179_not ; n26180
g25925 and n26177_not n26180 ; n26181
g25926 and n25872_not n26181_not ; n26182
g25927 and b[24] n25861_not ; n26183
g25928 and n25859_not n26183 ; n26184
g25929 and n25863_not n26184_not ; n26185
g25930 and n26182_not n26185 ; n26186
g25931 and n25863_not n26186_not ; n26187
g25932 and b[25] n25852_not ; n26188
g25933 and n25850_not n26188 ; n26189
g25934 and n25854_not n26189_not ; n26190
g25935 and n26187_not n26190 ; n26191
g25936 and n25854_not n26191_not ; n26192
g25937 and b[26] n25843_not ; n26193
g25938 and n25841_not n26193 ; n26194
g25939 and n25845_not n26194_not ; n26195
g25940 and n26192_not n26195 ; n26196
g25941 and n25845_not n26196_not ; n26197
g25942 and b[27] n25834_not ; n26198
g25943 and n25832_not n26198 ; n26199
g25944 and n25836_not n26199_not ; n26200
g25945 and n26197_not n26200 ; n26201
g25946 and n25836_not n26201_not ; n26202
g25947 and b[28] n25825_not ; n26203
g25948 and n25823_not n26203 ; n26204
g25949 and n25827_not n26204_not ; n26205
g25950 and n26202_not n26205 ; n26206
g25951 and n25827_not n26206_not ; n26207
g25952 and b[29] n25816_not ; n26208
g25953 and n25814_not n26208 ; n26209
g25954 and n25818_not n26209_not ; n26210
g25955 and n26207_not n26210 ; n26211
g25956 and n25818_not n26211_not ; n26212
g25957 and b[30] n25807_not ; n26213
g25958 and n25805_not n26213 ; n26214
g25959 and n25809_not n26214_not ; n26215
g25960 and n26212_not n26215 ; n26216
g25961 and n25809_not n26216_not ; n26217
g25962 and b[31] n25798_not ; n26218
g25963 and n25796_not n26218 ; n26219
g25964 and n25800_not n26219_not ; n26220
g25965 and n26217_not n26220 ; n26221
g25966 and n25800_not n26221_not ; n26222
g25967 and b[32] n25789_not ; n26223
g25968 and n25787_not n26223 ; n26224
g25969 and n25791_not n26224_not ; n26225
g25970 and n26222_not n26225 ; n26226
g25971 and n25791_not n26226_not ; n26227
g25972 and b[33] n25780_not ; n26228
g25973 and n25778_not n26228 ; n26229
g25974 and n25782_not n26229_not ; n26230
g25975 and n26227_not n26230 ; n26231
g25976 and n25782_not n26231_not ; n26232
g25977 and b[34] n25771_not ; n26233
g25978 and n25769_not n26233 ; n26234
g25979 and n25773_not n26234_not ; n26235
g25980 and n26232_not n26235 ; n26236
g25981 and n25773_not n26236_not ; n26237
g25982 and b[35] n25762_not ; n26238
g25983 and n25760_not n26238 ; n26239
g25984 and n25764_not n26239_not ; n26240
g25985 and n26237_not n26240 ; n26241
g25986 and n25764_not n26241_not ; n26242
g25987 and b[36] n25753_not ; n26243
g25988 and n25751_not n26243 ; n26244
g25989 and n25755_not n26244_not ; n26245
g25990 and n26242_not n26245 ; n26246
g25991 and n25755_not n26246_not ; n26247
g25992 and b[37] n25744_not ; n26248
g25993 and n25742_not n26248 ; n26249
g25994 and n25746_not n26249_not ; n26250
g25995 and n26247_not n26250 ; n26251
g25996 and n25746_not n26251_not ; n26252
g25997 and b[38] n25735_not ; n26253
g25998 and n25733_not n26253 ; n26254
g25999 and n25737_not n26254_not ; n26255
g26000 and n26252_not n26255 ; n26256
g26001 and n25737_not n26256_not ; n26257
g26002 and b[39] n25726_not ; n26258
g26003 and n25724_not n26258 ; n26259
g26004 and n25728_not n26259_not ; n26260
g26005 and n26257_not n26260 ; n26261
g26006 and n25728_not n26261_not ; n26262
g26007 and b[40] n25717_not ; n26263
g26008 and n25715_not n26263 ; n26264
g26009 and n25719_not n26264_not ; n26265
g26010 and n26262_not n26265 ; n26266
g26011 and n25719_not n26266_not ; n26267
g26012 and b[41] n25708_not ; n26268
g26013 and n25706_not n26268 ; n26269
g26014 and n25710_not n26269_not ; n26270
g26015 and n26267_not n26270 ; n26271
g26016 and n25710_not n26271_not ; n26272
g26017 and b[42] n25699_not ; n26273
g26018 and n25697_not n26273 ; n26274
g26019 and n25701_not n26274_not ; n26275
g26020 and n26272_not n26275 ; n26276
g26021 and n25701_not n26276_not ; n26277
g26022 and b[43] n25690_not ; n26278
g26023 and n25688_not n26278 ; n26279
g26024 and n25692_not n26279_not ; n26280
g26025 and n26277_not n26280 ; n26281
g26026 and n25692_not n26281_not ; n26282
g26027 and b[44] n25681_not ; n26283
g26028 and n25679_not n26283 ; n26284
g26029 and n25683_not n26284_not ; n26285
g26030 and n26282_not n26285 ; n26286
g26031 and n25683_not n26286_not ; n26287
g26032 and b[45] n25672_not ; n26288
g26033 and n25670_not n26288 ; n26289
g26034 and n25674_not n26289_not ; n26290
g26035 and n26287_not n26290 ; n26291
g26036 and n25674_not n26291_not ; n26292
g26037 and b[46] n25663_not ; n26293
g26038 and n25661_not n26293 ; n26294
g26039 and n25665_not n26294_not ; n26295
g26040 and n26292_not n26295 ; n26296
g26041 and n25665_not n26296_not ; n26297
g26042 and b[47] n25654_not ; n26298
g26043 and n25652_not n26298 ; n26299
g26044 and n25656_not n26299_not ; n26300
g26045 and n26297_not n26300 ; n26301
g26046 and n25656_not n26301_not ; n26302
g26047 and b[48] n25645_not ; n26303
g26048 and n25643_not n26303 ; n26304
g26049 and n25647_not n26304_not ; n26305
g26050 and n26302_not n26305 ; n26306
g26051 and n25647_not n26306_not ; n26307
g26052 and b[49] n25636_not ; n26308
g26053 and n25634_not n26308 ; n26309
g26054 and n25638_not n26309_not ; n26310
g26055 and n26307_not n26310 ; n26311
g26056 and n25638_not n26311_not ; n26312
g26057 and b[50] n25627_not ; n26313
g26058 and n25625_not n26313 ; n26314
g26059 and n25629_not n26314_not ; n26315
g26060 and n26312_not n26315 ; n26316
g26061 and n25629_not n26316_not ; n26317
g26062 and b[51] n25618_not ; n26318
g26063 and n25616_not n26318 ; n26319
g26064 and n25620_not n26319_not ; n26320
g26065 and n26317_not n26320 ; n26321
g26066 and n25620_not n26321_not ; n26322
g26067 and b[52] n25609_not ; n26323
g26068 and n25607_not n26323 ; n26324
g26069 and n25611_not n26324_not ; n26325
g26070 and n26322_not n26325 ; n26326
g26071 and n25611_not n26326_not ; n26327
g26072 and b[53] n25600_not ; n26328
g26073 and n25598_not n26328 ; n26329
g26074 and n25602_not n26329_not ; n26330
g26075 and n26327_not n26330 ; n26331
g26076 and n25602_not n26331_not ; n26332
g26077 and b[54] n25591_not ; n26333
g26078 and n25589_not n26333 ; n26334
g26079 and n25593_not n26334_not ; n26335
g26080 and n26332_not n26335 ; n26336
g26081 and n25593_not n26336_not ; n26337
g26082 and b[55] n25582_not ; n26338
g26083 and n25580_not n26338 ; n26339
g26084 and n25584_not n26339_not ; n26340
g26085 and n26337_not n26340 ; n26341
g26086 and n25584_not n26341_not ; n26342
g26087 and b[56] n25573_not ; n26343
g26088 and n25571_not n26343 ; n26344
g26089 and n25575_not n26344_not ; n26345
g26090 and n26342_not n26345 ; n26346
g26091 and n25575_not n26346_not ; n26347
g26092 and b[57] n25564_not ; n26348
g26093 and n25562_not n26348 ; n26349
g26094 and n25566_not n26349_not ; n26350
g26095 and n26347_not n26350 ; n26351
g26096 and n25566_not n26351_not ; n26352
g26097 and b[58] n25555_not ; n26353
g26098 and n25553_not n26353 ; n26354
g26099 and n25557_not n26354_not ; n26355
g26100 and n26352_not n26355 ; n26356
g26101 and n25557_not n26356_not ; n26357
g26102 and b[59] n25546_not ; n26358
g26103 and n25544_not n26358 ; n26359
g26104 and n25548_not n26359_not ; n26360
g26105 and n26357_not n26360 ; n26361
g26106 and n25548_not n26361_not ; n26362
g26107 and n24721_not n25534_not ; n26363
g26108 and n25532_not n26363 ; n26364
g26109 and n25520_not n26364 ; n26365
g26110 and n25532_not n25534_not ; n26366
g26111 and n25521_not n26366_not ; n26367
g26112 and n26365_not n26367_not ; n26368
g26113 and quotient[4] n26368_not ; n26369
g26114 and n25531_not n25538_not ; n26370
g26115 and n25537_not n26370 ; n26371
g26116 and n26369_not n26371_not ; n26372
g26117 and b[60]_not n26372_not ; n26373
g26118 and b[60] n26371_not ; n26374
g26119 and n26369_not n26374 ; n26375
g26120 and n403 n26375_not ; n26376
g26121 and n26373_not n26376 ; n26377
g26122 and n26362_not n26377 ; n26378
g26123 and n280 n26372_not ; n26379
g26124 and n26378_not n26379_not ; quotient[3]
g26125 and n25557_not n26360 ; n26381
g26126 and n26356_not n26381 ; n26382
g26127 and n26357_not n26360_not ; n26383
g26128 and n26382_not n26383_not ; n26384
g26129 and quotient[3] n26384_not ; n26385
g26130 and n25547_not n26379_not ; n26386
g26131 and n26378_not n26386 ; n26387
g26132 and n26385_not n26387_not ; n26388
g26133 and b[60]_not n26388_not ; n26389
g26134 and n25566_not n26355 ; n26390
g26135 and n26351_not n26390 ; n26391
g26136 and n26352_not n26355_not ; n26392
g26137 and n26391_not n26392_not ; n26393
g26138 and quotient[3] n26393_not ; n26394
g26139 and n25556_not n26379_not ; n26395
g26140 and n26378_not n26395 ; n26396
g26141 and n26394_not n26396_not ; n26397
g26142 and b[59]_not n26397_not ; n26398
g26143 and n25575_not n26350 ; n26399
g26144 and n26346_not n26399 ; n26400
g26145 and n26347_not n26350_not ; n26401
g26146 and n26400_not n26401_not ; n26402
g26147 and quotient[3] n26402_not ; n26403
g26148 and n25565_not n26379_not ; n26404
g26149 and n26378_not n26404 ; n26405
g26150 and n26403_not n26405_not ; n26406
g26151 and b[58]_not n26406_not ; n26407
g26152 and n25584_not n26345 ; n26408
g26153 and n26341_not n26408 ; n26409
g26154 and n26342_not n26345_not ; n26410
g26155 and n26409_not n26410_not ; n26411
g26156 and quotient[3] n26411_not ; n26412
g26157 and n25574_not n26379_not ; n26413
g26158 and n26378_not n26413 ; n26414
g26159 and n26412_not n26414_not ; n26415
g26160 and b[57]_not n26415_not ; n26416
g26161 and n25593_not n26340 ; n26417
g26162 and n26336_not n26417 ; n26418
g26163 and n26337_not n26340_not ; n26419
g26164 and n26418_not n26419_not ; n26420
g26165 and quotient[3] n26420_not ; n26421
g26166 and n25583_not n26379_not ; n26422
g26167 and n26378_not n26422 ; n26423
g26168 and n26421_not n26423_not ; n26424
g26169 and b[56]_not n26424_not ; n26425
g26170 and n25602_not n26335 ; n26426
g26171 and n26331_not n26426 ; n26427
g26172 and n26332_not n26335_not ; n26428
g26173 and n26427_not n26428_not ; n26429
g26174 and quotient[3] n26429_not ; n26430
g26175 and n25592_not n26379_not ; n26431
g26176 and n26378_not n26431 ; n26432
g26177 and n26430_not n26432_not ; n26433
g26178 and b[55]_not n26433_not ; n26434
g26179 and n25611_not n26330 ; n26435
g26180 and n26326_not n26435 ; n26436
g26181 and n26327_not n26330_not ; n26437
g26182 and n26436_not n26437_not ; n26438
g26183 and quotient[3] n26438_not ; n26439
g26184 and n25601_not n26379_not ; n26440
g26185 and n26378_not n26440 ; n26441
g26186 and n26439_not n26441_not ; n26442
g26187 and b[54]_not n26442_not ; n26443
g26188 and n25620_not n26325 ; n26444
g26189 and n26321_not n26444 ; n26445
g26190 and n26322_not n26325_not ; n26446
g26191 and n26445_not n26446_not ; n26447
g26192 and quotient[3] n26447_not ; n26448
g26193 and n25610_not n26379_not ; n26449
g26194 and n26378_not n26449 ; n26450
g26195 and n26448_not n26450_not ; n26451
g26196 and b[53]_not n26451_not ; n26452
g26197 and n25629_not n26320 ; n26453
g26198 and n26316_not n26453 ; n26454
g26199 and n26317_not n26320_not ; n26455
g26200 and n26454_not n26455_not ; n26456
g26201 and quotient[3] n26456_not ; n26457
g26202 and n25619_not n26379_not ; n26458
g26203 and n26378_not n26458 ; n26459
g26204 and n26457_not n26459_not ; n26460
g26205 and b[52]_not n26460_not ; n26461
g26206 and n25638_not n26315 ; n26462
g26207 and n26311_not n26462 ; n26463
g26208 and n26312_not n26315_not ; n26464
g26209 and n26463_not n26464_not ; n26465
g26210 and quotient[3] n26465_not ; n26466
g26211 and n25628_not n26379_not ; n26467
g26212 and n26378_not n26467 ; n26468
g26213 and n26466_not n26468_not ; n26469
g26214 and b[51]_not n26469_not ; n26470
g26215 and n25647_not n26310 ; n26471
g26216 and n26306_not n26471 ; n26472
g26217 and n26307_not n26310_not ; n26473
g26218 and n26472_not n26473_not ; n26474
g26219 and quotient[3] n26474_not ; n26475
g26220 and n25637_not n26379_not ; n26476
g26221 and n26378_not n26476 ; n26477
g26222 and n26475_not n26477_not ; n26478
g26223 and b[50]_not n26478_not ; n26479
g26224 and n25656_not n26305 ; n26480
g26225 and n26301_not n26480 ; n26481
g26226 and n26302_not n26305_not ; n26482
g26227 and n26481_not n26482_not ; n26483
g26228 and quotient[3] n26483_not ; n26484
g26229 and n25646_not n26379_not ; n26485
g26230 and n26378_not n26485 ; n26486
g26231 and n26484_not n26486_not ; n26487
g26232 and b[49]_not n26487_not ; n26488
g26233 and n25665_not n26300 ; n26489
g26234 and n26296_not n26489 ; n26490
g26235 and n26297_not n26300_not ; n26491
g26236 and n26490_not n26491_not ; n26492
g26237 and quotient[3] n26492_not ; n26493
g26238 and n25655_not n26379_not ; n26494
g26239 and n26378_not n26494 ; n26495
g26240 and n26493_not n26495_not ; n26496
g26241 and b[48]_not n26496_not ; n26497
g26242 and n25674_not n26295 ; n26498
g26243 and n26291_not n26498 ; n26499
g26244 and n26292_not n26295_not ; n26500
g26245 and n26499_not n26500_not ; n26501
g26246 and quotient[3] n26501_not ; n26502
g26247 and n25664_not n26379_not ; n26503
g26248 and n26378_not n26503 ; n26504
g26249 and n26502_not n26504_not ; n26505
g26250 and b[47]_not n26505_not ; n26506
g26251 and n25683_not n26290 ; n26507
g26252 and n26286_not n26507 ; n26508
g26253 and n26287_not n26290_not ; n26509
g26254 and n26508_not n26509_not ; n26510
g26255 and quotient[3] n26510_not ; n26511
g26256 and n25673_not n26379_not ; n26512
g26257 and n26378_not n26512 ; n26513
g26258 and n26511_not n26513_not ; n26514
g26259 and b[46]_not n26514_not ; n26515
g26260 and n25692_not n26285 ; n26516
g26261 and n26281_not n26516 ; n26517
g26262 and n26282_not n26285_not ; n26518
g26263 and n26517_not n26518_not ; n26519
g26264 and quotient[3] n26519_not ; n26520
g26265 and n25682_not n26379_not ; n26521
g26266 and n26378_not n26521 ; n26522
g26267 and n26520_not n26522_not ; n26523
g26268 and b[45]_not n26523_not ; n26524
g26269 and n25701_not n26280 ; n26525
g26270 and n26276_not n26525 ; n26526
g26271 and n26277_not n26280_not ; n26527
g26272 and n26526_not n26527_not ; n26528
g26273 and quotient[3] n26528_not ; n26529
g26274 and n25691_not n26379_not ; n26530
g26275 and n26378_not n26530 ; n26531
g26276 and n26529_not n26531_not ; n26532
g26277 and b[44]_not n26532_not ; n26533
g26278 and n25710_not n26275 ; n26534
g26279 and n26271_not n26534 ; n26535
g26280 and n26272_not n26275_not ; n26536
g26281 and n26535_not n26536_not ; n26537
g26282 and quotient[3] n26537_not ; n26538
g26283 and n25700_not n26379_not ; n26539
g26284 and n26378_not n26539 ; n26540
g26285 and n26538_not n26540_not ; n26541
g26286 and b[43]_not n26541_not ; n26542
g26287 and n25719_not n26270 ; n26543
g26288 and n26266_not n26543 ; n26544
g26289 and n26267_not n26270_not ; n26545
g26290 and n26544_not n26545_not ; n26546
g26291 and quotient[3] n26546_not ; n26547
g26292 and n25709_not n26379_not ; n26548
g26293 and n26378_not n26548 ; n26549
g26294 and n26547_not n26549_not ; n26550
g26295 and b[42]_not n26550_not ; n26551
g26296 and n25728_not n26265 ; n26552
g26297 and n26261_not n26552 ; n26553
g26298 and n26262_not n26265_not ; n26554
g26299 and n26553_not n26554_not ; n26555
g26300 and quotient[3] n26555_not ; n26556
g26301 and n25718_not n26379_not ; n26557
g26302 and n26378_not n26557 ; n26558
g26303 and n26556_not n26558_not ; n26559
g26304 and b[41]_not n26559_not ; n26560
g26305 and n25737_not n26260 ; n26561
g26306 and n26256_not n26561 ; n26562
g26307 and n26257_not n26260_not ; n26563
g26308 and n26562_not n26563_not ; n26564
g26309 and quotient[3] n26564_not ; n26565
g26310 and n25727_not n26379_not ; n26566
g26311 and n26378_not n26566 ; n26567
g26312 and n26565_not n26567_not ; n26568
g26313 and b[40]_not n26568_not ; n26569
g26314 and n25746_not n26255 ; n26570
g26315 and n26251_not n26570 ; n26571
g26316 and n26252_not n26255_not ; n26572
g26317 and n26571_not n26572_not ; n26573
g26318 and quotient[3] n26573_not ; n26574
g26319 and n25736_not n26379_not ; n26575
g26320 and n26378_not n26575 ; n26576
g26321 and n26574_not n26576_not ; n26577
g26322 and b[39]_not n26577_not ; n26578
g26323 and n25755_not n26250 ; n26579
g26324 and n26246_not n26579 ; n26580
g26325 and n26247_not n26250_not ; n26581
g26326 and n26580_not n26581_not ; n26582
g26327 and quotient[3] n26582_not ; n26583
g26328 and n25745_not n26379_not ; n26584
g26329 and n26378_not n26584 ; n26585
g26330 and n26583_not n26585_not ; n26586
g26331 and b[38]_not n26586_not ; n26587
g26332 and n25764_not n26245 ; n26588
g26333 and n26241_not n26588 ; n26589
g26334 and n26242_not n26245_not ; n26590
g26335 and n26589_not n26590_not ; n26591
g26336 and quotient[3] n26591_not ; n26592
g26337 and n25754_not n26379_not ; n26593
g26338 and n26378_not n26593 ; n26594
g26339 and n26592_not n26594_not ; n26595
g26340 and b[37]_not n26595_not ; n26596
g26341 and n25773_not n26240 ; n26597
g26342 and n26236_not n26597 ; n26598
g26343 and n26237_not n26240_not ; n26599
g26344 and n26598_not n26599_not ; n26600
g26345 and quotient[3] n26600_not ; n26601
g26346 and n25763_not n26379_not ; n26602
g26347 and n26378_not n26602 ; n26603
g26348 and n26601_not n26603_not ; n26604
g26349 and b[36]_not n26604_not ; n26605
g26350 and n25782_not n26235 ; n26606
g26351 and n26231_not n26606 ; n26607
g26352 and n26232_not n26235_not ; n26608
g26353 and n26607_not n26608_not ; n26609
g26354 and quotient[3] n26609_not ; n26610
g26355 and n25772_not n26379_not ; n26611
g26356 and n26378_not n26611 ; n26612
g26357 and n26610_not n26612_not ; n26613
g26358 and b[35]_not n26613_not ; n26614
g26359 and n25791_not n26230 ; n26615
g26360 and n26226_not n26615 ; n26616
g26361 and n26227_not n26230_not ; n26617
g26362 and n26616_not n26617_not ; n26618
g26363 and quotient[3] n26618_not ; n26619
g26364 and n25781_not n26379_not ; n26620
g26365 and n26378_not n26620 ; n26621
g26366 and n26619_not n26621_not ; n26622
g26367 and b[34]_not n26622_not ; n26623
g26368 and n25800_not n26225 ; n26624
g26369 and n26221_not n26624 ; n26625
g26370 and n26222_not n26225_not ; n26626
g26371 and n26625_not n26626_not ; n26627
g26372 and quotient[3] n26627_not ; n26628
g26373 and n25790_not n26379_not ; n26629
g26374 and n26378_not n26629 ; n26630
g26375 and n26628_not n26630_not ; n26631
g26376 and b[33]_not n26631_not ; n26632
g26377 and n25809_not n26220 ; n26633
g26378 and n26216_not n26633 ; n26634
g26379 and n26217_not n26220_not ; n26635
g26380 and n26634_not n26635_not ; n26636
g26381 and quotient[3] n26636_not ; n26637
g26382 and n25799_not n26379_not ; n26638
g26383 and n26378_not n26638 ; n26639
g26384 and n26637_not n26639_not ; n26640
g26385 and b[32]_not n26640_not ; n26641
g26386 and n25818_not n26215 ; n26642
g26387 and n26211_not n26642 ; n26643
g26388 and n26212_not n26215_not ; n26644
g26389 and n26643_not n26644_not ; n26645
g26390 and quotient[3] n26645_not ; n26646
g26391 and n25808_not n26379_not ; n26647
g26392 and n26378_not n26647 ; n26648
g26393 and n26646_not n26648_not ; n26649
g26394 and b[31]_not n26649_not ; n26650
g26395 and n25827_not n26210 ; n26651
g26396 and n26206_not n26651 ; n26652
g26397 and n26207_not n26210_not ; n26653
g26398 and n26652_not n26653_not ; n26654
g26399 and quotient[3] n26654_not ; n26655
g26400 and n25817_not n26379_not ; n26656
g26401 and n26378_not n26656 ; n26657
g26402 and n26655_not n26657_not ; n26658
g26403 and b[30]_not n26658_not ; n26659
g26404 and n25836_not n26205 ; n26660
g26405 and n26201_not n26660 ; n26661
g26406 and n26202_not n26205_not ; n26662
g26407 and n26661_not n26662_not ; n26663
g26408 and quotient[3] n26663_not ; n26664
g26409 and n25826_not n26379_not ; n26665
g26410 and n26378_not n26665 ; n26666
g26411 and n26664_not n26666_not ; n26667
g26412 and b[29]_not n26667_not ; n26668
g26413 and n25845_not n26200 ; n26669
g26414 and n26196_not n26669 ; n26670
g26415 and n26197_not n26200_not ; n26671
g26416 and n26670_not n26671_not ; n26672
g26417 and quotient[3] n26672_not ; n26673
g26418 and n25835_not n26379_not ; n26674
g26419 and n26378_not n26674 ; n26675
g26420 and n26673_not n26675_not ; n26676
g26421 and b[28]_not n26676_not ; n26677
g26422 and n25854_not n26195 ; n26678
g26423 and n26191_not n26678 ; n26679
g26424 and n26192_not n26195_not ; n26680
g26425 and n26679_not n26680_not ; n26681
g26426 and quotient[3] n26681_not ; n26682
g26427 and n25844_not n26379_not ; n26683
g26428 and n26378_not n26683 ; n26684
g26429 and n26682_not n26684_not ; n26685
g26430 and b[27]_not n26685_not ; n26686
g26431 and n25863_not n26190 ; n26687
g26432 and n26186_not n26687 ; n26688
g26433 and n26187_not n26190_not ; n26689
g26434 and n26688_not n26689_not ; n26690
g26435 and quotient[3] n26690_not ; n26691
g26436 and n25853_not n26379_not ; n26692
g26437 and n26378_not n26692 ; n26693
g26438 and n26691_not n26693_not ; n26694
g26439 and b[26]_not n26694_not ; n26695
g26440 and n25872_not n26185 ; n26696
g26441 and n26181_not n26696 ; n26697
g26442 and n26182_not n26185_not ; n26698
g26443 and n26697_not n26698_not ; n26699
g26444 and quotient[3] n26699_not ; n26700
g26445 and n25862_not n26379_not ; n26701
g26446 and n26378_not n26701 ; n26702
g26447 and n26700_not n26702_not ; n26703
g26448 and b[25]_not n26703_not ; n26704
g26449 and n25881_not n26180 ; n26705
g26450 and n26176_not n26705 ; n26706
g26451 and n26177_not n26180_not ; n26707
g26452 and n26706_not n26707_not ; n26708
g26453 and quotient[3] n26708_not ; n26709
g26454 and n25871_not n26379_not ; n26710
g26455 and n26378_not n26710 ; n26711
g26456 and n26709_not n26711_not ; n26712
g26457 and b[24]_not n26712_not ; n26713
g26458 and n25890_not n26175 ; n26714
g26459 and n26171_not n26714 ; n26715
g26460 and n26172_not n26175_not ; n26716
g26461 and n26715_not n26716_not ; n26717
g26462 and quotient[3] n26717_not ; n26718
g26463 and n25880_not n26379_not ; n26719
g26464 and n26378_not n26719 ; n26720
g26465 and n26718_not n26720_not ; n26721
g26466 and b[23]_not n26721_not ; n26722
g26467 and n25899_not n26170 ; n26723
g26468 and n26166_not n26723 ; n26724
g26469 and n26167_not n26170_not ; n26725
g26470 and n26724_not n26725_not ; n26726
g26471 and quotient[3] n26726_not ; n26727
g26472 and n25889_not n26379_not ; n26728
g26473 and n26378_not n26728 ; n26729
g26474 and n26727_not n26729_not ; n26730
g26475 and b[22]_not n26730_not ; n26731
g26476 and n25908_not n26165 ; n26732
g26477 and n26161_not n26732 ; n26733
g26478 and n26162_not n26165_not ; n26734
g26479 and n26733_not n26734_not ; n26735
g26480 and quotient[3] n26735_not ; n26736
g26481 and n25898_not n26379_not ; n26737
g26482 and n26378_not n26737 ; n26738
g26483 and n26736_not n26738_not ; n26739
g26484 and b[21]_not n26739_not ; n26740
g26485 and n25917_not n26160 ; n26741
g26486 and n26156_not n26741 ; n26742
g26487 and n26157_not n26160_not ; n26743
g26488 and n26742_not n26743_not ; n26744
g26489 and quotient[3] n26744_not ; n26745
g26490 and n25907_not n26379_not ; n26746
g26491 and n26378_not n26746 ; n26747
g26492 and n26745_not n26747_not ; n26748
g26493 and b[20]_not n26748_not ; n26749
g26494 and n25926_not n26155 ; n26750
g26495 and n26151_not n26750 ; n26751
g26496 and n26152_not n26155_not ; n26752
g26497 and n26751_not n26752_not ; n26753
g26498 and quotient[3] n26753_not ; n26754
g26499 and n25916_not n26379_not ; n26755
g26500 and n26378_not n26755 ; n26756
g26501 and n26754_not n26756_not ; n26757
g26502 and b[19]_not n26757_not ; n26758
g26503 and n25935_not n26150 ; n26759
g26504 and n26146_not n26759 ; n26760
g26505 and n26147_not n26150_not ; n26761
g26506 and n26760_not n26761_not ; n26762
g26507 and quotient[3] n26762_not ; n26763
g26508 and n25925_not n26379_not ; n26764
g26509 and n26378_not n26764 ; n26765
g26510 and n26763_not n26765_not ; n26766
g26511 and b[18]_not n26766_not ; n26767
g26512 and n25944_not n26145 ; n26768
g26513 and n26141_not n26768 ; n26769
g26514 and n26142_not n26145_not ; n26770
g26515 and n26769_not n26770_not ; n26771
g26516 and quotient[3] n26771_not ; n26772
g26517 and n25934_not n26379_not ; n26773
g26518 and n26378_not n26773 ; n26774
g26519 and n26772_not n26774_not ; n26775
g26520 and b[17]_not n26775_not ; n26776
g26521 and n25953_not n26140 ; n26777
g26522 and n26136_not n26777 ; n26778
g26523 and n26137_not n26140_not ; n26779
g26524 and n26778_not n26779_not ; n26780
g26525 and quotient[3] n26780_not ; n26781
g26526 and n25943_not n26379_not ; n26782
g26527 and n26378_not n26782 ; n26783
g26528 and n26781_not n26783_not ; n26784
g26529 and b[16]_not n26784_not ; n26785
g26530 and n25962_not n26135 ; n26786
g26531 and n26131_not n26786 ; n26787
g26532 and n26132_not n26135_not ; n26788
g26533 and n26787_not n26788_not ; n26789
g26534 and quotient[3] n26789_not ; n26790
g26535 and n25952_not n26379_not ; n26791
g26536 and n26378_not n26791 ; n26792
g26537 and n26790_not n26792_not ; n26793
g26538 and b[15]_not n26793_not ; n26794
g26539 and n25971_not n26130 ; n26795
g26540 and n26126_not n26795 ; n26796
g26541 and n26127_not n26130_not ; n26797
g26542 and n26796_not n26797_not ; n26798
g26543 and quotient[3] n26798_not ; n26799
g26544 and n25961_not n26379_not ; n26800
g26545 and n26378_not n26800 ; n26801
g26546 and n26799_not n26801_not ; n26802
g26547 and b[14]_not n26802_not ; n26803
g26548 and n25980_not n26125 ; n26804
g26549 and n26121_not n26804 ; n26805
g26550 and n26122_not n26125_not ; n26806
g26551 and n26805_not n26806_not ; n26807
g26552 and quotient[3] n26807_not ; n26808
g26553 and n25970_not n26379_not ; n26809
g26554 and n26378_not n26809 ; n26810
g26555 and n26808_not n26810_not ; n26811
g26556 and b[13]_not n26811_not ; n26812
g26557 and n25989_not n26120 ; n26813
g26558 and n26116_not n26813 ; n26814
g26559 and n26117_not n26120_not ; n26815
g26560 and n26814_not n26815_not ; n26816
g26561 and quotient[3] n26816_not ; n26817
g26562 and n25979_not n26379_not ; n26818
g26563 and n26378_not n26818 ; n26819
g26564 and n26817_not n26819_not ; n26820
g26565 and b[12]_not n26820_not ; n26821
g26566 and n25998_not n26115 ; n26822
g26567 and n26111_not n26822 ; n26823
g26568 and n26112_not n26115_not ; n26824
g26569 and n26823_not n26824_not ; n26825
g26570 and quotient[3] n26825_not ; n26826
g26571 and n25988_not n26379_not ; n26827
g26572 and n26378_not n26827 ; n26828
g26573 and n26826_not n26828_not ; n26829
g26574 and b[11]_not n26829_not ; n26830
g26575 and n26007_not n26110 ; n26831
g26576 and n26106_not n26831 ; n26832
g26577 and n26107_not n26110_not ; n26833
g26578 and n26832_not n26833_not ; n26834
g26579 and quotient[3] n26834_not ; n26835
g26580 and n25997_not n26379_not ; n26836
g26581 and n26378_not n26836 ; n26837
g26582 and n26835_not n26837_not ; n26838
g26583 and b[10]_not n26838_not ; n26839
g26584 and n26016_not n26105 ; n26840
g26585 and n26101_not n26840 ; n26841
g26586 and n26102_not n26105_not ; n26842
g26587 and n26841_not n26842_not ; n26843
g26588 and quotient[3] n26843_not ; n26844
g26589 and n26006_not n26379_not ; n26845
g26590 and n26378_not n26845 ; n26846
g26591 and n26844_not n26846_not ; n26847
g26592 and b[9]_not n26847_not ; n26848
g26593 and n26025_not n26100 ; n26849
g26594 and n26096_not n26849 ; n26850
g26595 and n26097_not n26100_not ; n26851
g26596 and n26850_not n26851_not ; n26852
g26597 and quotient[3] n26852_not ; n26853
g26598 and n26015_not n26379_not ; n26854
g26599 and n26378_not n26854 ; n26855
g26600 and n26853_not n26855_not ; n26856
g26601 and b[8]_not n26856_not ; n26857
g26602 and n26034_not n26095 ; n26858
g26603 and n26091_not n26858 ; n26859
g26604 and n26092_not n26095_not ; n26860
g26605 and n26859_not n26860_not ; n26861
g26606 and quotient[3] n26861_not ; n26862
g26607 and n26024_not n26379_not ; n26863
g26608 and n26378_not n26863 ; n26864
g26609 and n26862_not n26864_not ; n26865
g26610 and b[7]_not n26865_not ; n26866
g26611 and n26043_not n26090 ; n26867
g26612 and n26086_not n26867 ; n26868
g26613 and n26087_not n26090_not ; n26869
g26614 and n26868_not n26869_not ; n26870
g26615 and quotient[3] n26870_not ; n26871
g26616 and n26033_not n26379_not ; n26872
g26617 and n26378_not n26872 ; n26873
g26618 and n26871_not n26873_not ; n26874
g26619 and b[6]_not n26874_not ; n26875
g26620 and n26052_not n26085 ; n26876
g26621 and n26081_not n26876 ; n26877
g26622 and n26082_not n26085_not ; n26878
g26623 and n26877_not n26878_not ; n26879
g26624 and quotient[3] n26879_not ; n26880
g26625 and n26042_not n26379_not ; n26881
g26626 and n26378_not n26881 ; n26882
g26627 and n26880_not n26882_not ; n26883
g26628 and b[5]_not n26883_not ; n26884
g26629 and n26060_not n26080 ; n26885
g26630 and n26076_not n26885 ; n26886
g26631 and n26077_not n26080_not ; n26887
g26632 and n26886_not n26887_not ; n26888
g26633 and quotient[3] n26888_not ; n26889
g26634 and n26051_not n26379_not ; n26890
g26635 and n26378_not n26890 ; n26891
g26636 and n26889_not n26891_not ; n26892
g26637 and b[4]_not n26892_not ; n26893
g26638 and n26071_not n26075 ; n26894
g26639 and n26070_not n26894 ; n26895
g26640 and n26072_not n26075_not ; n26896
g26641 and n26895_not n26896_not ; n26897
g26642 and quotient[3] n26897_not ; n26898
g26643 and n26059_not n26379_not ; n26899
g26644 and n26378_not n26899 ; n26900
g26645 and n26898_not n26900_not ; n26901
g26646 and b[3]_not n26901_not ; n26902
g26647 and n26067_not n26069 ; n26903
g26648 and n26065_not n26903 ; n26904
g26649 and n26070_not n26904_not ; n26905
g26650 and quotient[3] n26905 ; n26906
g26651 and n26064_not n26379_not ; n26907
g26652 and n26378_not n26907 ; n26908
g26653 and n26906_not n26908_not ; n26909
g26654 and b[2]_not n26909_not ; n26910
g26655 and b[0] quotient[3] ; n26911
g26656 and a[3] n26911_not ; n26912
g26657 and n26069 quotient[3] ; n26913
g26658 and n26912_not n26913_not ; n26914
g26659 and b[1] n26914_not ; n26915
g26660 and b[1]_not n26913_not ; n26916
g26661 and n26912_not n26916 ; n26917
g26662 and n26915_not n26917_not ; n26918
g26663 and a[2]_not b[0] ; n26919
g26664 and n26918_not n26919_not ; n26920
g26665 and b[1]_not n26914_not ; n26921
g26666 and n26920_not n26921_not ; n26922
g26667 and b[2] n26908_not ; n26923
g26668 and n26906_not n26923 ; n26924
g26669 and n26910_not n26924_not ; n26925
g26670 and n26922_not n26925 ; n26926
g26671 and n26910_not n26926_not ; n26927
g26672 and b[3] n26900_not ; n26928
g26673 and n26898_not n26928 ; n26929
g26674 and n26902_not n26929_not ; n26930
g26675 and n26927_not n26930 ; n26931
g26676 and n26902_not n26931_not ; n26932
g26677 and b[4] n26891_not ; n26933
g26678 and n26889_not n26933 ; n26934
g26679 and n26893_not n26934_not ; n26935
g26680 and n26932_not n26935 ; n26936
g26681 and n26893_not n26936_not ; n26937
g26682 and b[5] n26882_not ; n26938
g26683 and n26880_not n26938 ; n26939
g26684 and n26884_not n26939_not ; n26940
g26685 and n26937_not n26940 ; n26941
g26686 and n26884_not n26941_not ; n26942
g26687 and b[6] n26873_not ; n26943
g26688 and n26871_not n26943 ; n26944
g26689 and n26875_not n26944_not ; n26945
g26690 and n26942_not n26945 ; n26946
g26691 and n26875_not n26946_not ; n26947
g26692 and b[7] n26864_not ; n26948
g26693 and n26862_not n26948 ; n26949
g26694 and n26866_not n26949_not ; n26950
g26695 and n26947_not n26950 ; n26951
g26696 and n26866_not n26951_not ; n26952
g26697 and b[8] n26855_not ; n26953
g26698 and n26853_not n26953 ; n26954
g26699 and n26857_not n26954_not ; n26955
g26700 and n26952_not n26955 ; n26956
g26701 and n26857_not n26956_not ; n26957
g26702 and b[9] n26846_not ; n26958
g26703 and n26844_not n26958 ; n26959
g26704 and n26848_not n26959_not ; n26960
g26705 and n26957_not n26960 ; n26961
g26706 and n26848_not n26961_not ; n26962
g26707 and b[10] n26837_not ; n26963
g26708 and n26835_not n26963 ; n26964
g26709 and n26839_not n26964_not ; n26965
g26710 and n26962_not n26965 ; n26966
g26711 and n26839_not n26966_not ; n26967
g26712 and b[11] n26828_not ; n26968
g26713 and n26826_not n26968 ; n26969
g26714 and n26830_not n26969_not ; n26970
g26715 and n26967_not n26970 ; n26971
g26716 and n26830_not n26971_not ; n26972
g26717 and b[12] n26819_not ; n26973
g26718 and n26817_not n26973 ; n26974
g26719 and n26821_not n26974_not ; n26975
g26720 and n26972_not n26975 ; n26976
g26721 and n26821_not n26976_not ; n26977
g26722 and b[13] n26810_not ; n26978
g26723 and n26808_not n26978 ; n26979
g26724 and n26812_not n26979_not ; n26980
g26725 and n26977_not n26980 ; n26981
g26726 and n26812_not n26981_not ; n26982
g26727 and b[14] n26801_not ; n26983
g26728 and n26799_not n26983 ; n26984
g26729 and n26803_not n26984_not ; n26985
g26730 and n26982_not n26985 ; n26986
g26731 and n26803_not n26986_not ; n26987
g26732 and b[15] n26792_not ; n26988
g26733 and n26790_not n26988 ; n26989
g26734 and n26794_not n26989_not ; n26990
g26735 and n26987_not n26990 ; n26991
g26736 and n26794_not n26991_not ; n26992
g26737 and b[16] n26783_not ; n26993
g26738 and n26781_not n26993 ; n26994
g26739 and n26785_not n26994_not ; n26995
g26740 and n26992_not n26995 ; n26996
g26741 and n26785_not n26996_not ; n26997
g26742 and b[17] n26774_not ; n26998
g26743 and n26772_not n26998 ; n26999
g26744 and n26776_not n26999_not ; n27000
g26745 and n26997_not n27000 ; n27001
g26746 and n26776_not n27001_not ; n27002
g26747 and b[18] n26765_not ; n27003
g26748 and n26763_not n27003 ; n27004
g26749 and n26767_not n27004_not ; n27005
g26750 and n27002_not n27005 ; n27006
g26751 and n26767_not n27006_not ; n27007
g26752 and b[19] n26756_not ; n27008
g26753 and n26754_not n27008 ; n27009
g26754 and n26758_not n27009_not ; n27010
g26755 and n27007_not n27010 ; n27011
g26756 and n26758_not n27011_not ; n27012
g26757 and b[20] n26747_not ; n27013
g26758 and n26745_not n27013 ; n27014
g26759 and n26749_not n27014_not ; n27015
g26760 and n27012_not n27015 ; n27016
g26761 and n26749_not n27016_not ; n27017
g26762 and b[21] n26738_not ; n27018
g26763 and n26736_not n27018 ; n27019
g26764 and n26740_not n27019_not ; n27020
g26765 and n27017_not n27020 ; n27021
g26766 and n26740_not n27021_not ; n27022
g26767 and b[22] n26729_not ; n27023
g26768 and n26727_not n27023 ; n27024
g26769 and n26731_not n27024_not ; n27025
g26770 and n27022_not n27025 ; n27026
g26771 and n26731_not n27026_not ; n27027
g26772 and b[23] n26720_not ; n27028
g26773 and n26718_not n27028 ; n27029
g26774 and n26722_not n27029_not ; n27030
g26775 and n27027_not n27030 ; n27031
g26776 and n26722_not n27031_not ; n27032
g26777 and b[24] n26711_not ; n27033
g26778 and n26709_not n27033 ; n27034
g26779 and n26713_not n27034_not ; n27035
g26780 and n27032_not n27035 ; n27036
g26781 and n26713_not n27036_not ; n27037
g26782 and b[25] n26702_not ; n27038
g26783 and n26700_not n27038 ; n27039
g26784 and n26704_not n27039_not ; n27040
g26785 and n27037_not n27040 ; n27041
g26786 and n26704_not n27041_not ; n27042
g26787 and b[26] n26693_not ; n27043
g26788 and n26691_not n27043 ; n27044
g26789 and n26695_not n27044_not ; n27045
g26790 and n27042_not n27045 ; n27046
g26791 and n26695_not n27046_not ; n27047
g26792 and b[27] n26684_not ; n27048
g26793 and n26682_not n27048 ; n27049
g26794 and n26686_not n27049_not ; n27050
g26795 and n27047_not n27050 ; n27051
g26796 and n26686_not n27051_not ; n27052
g26797 and b[28] n26675_not ; n27053
g26798 and n26673_not n27053 ; n27054
g26799 and n26677_not n27054_not ; n27055
g26800 and n27052_not n27055 ; n27056
g26801 and n26677_not n27056_not ; n27057
g26802 and b[29] n26666_not ; n27058
g26803 and n26664_not n27058 ; n27059
g26804 and n26668_not n27059_not ; n27060
g26805 and n27057_not n27060 ; n27061
g26806 and n26668_not n27061_not ; n27062
g26807 and b[30] n26657_not ; n27063
g26808 and n26655_not n27063 ; n27064
g26809 and n26659_not n27064_not ; n27065
g26810 and n27062_not n27065 ; n27066
g26811 and n26659_not n27066_not ; n27067
g26812 and b[31] n26648_not ; n27068
g26813 and n26646_not n27068 ; n27069
g26814 and n26650_not n27069_not ; n27070
g26815 and n27067_not n27070 ; n27071
g26816 and n26650_not n27071_not ; n27072
g26817 and b[32] n26639_not ; n27073
g26818 and n26637_not n27073 ; n27074
g26819 and n26641_not n27074_not ; n27075
g26820 and n27072_not n27075 ; n27076
g26821 and n26641_not n27076_not ; n27077
g26822 and b[33] n26630_not ; n27078
g26823 and n26628_not n27078 ; n27079
g26824 and n26632_not n27079_not ; n27080
g26825 and n27077_not n27080 ; n27081
g26826 and n26632_not n27081_not ; n27082
g26827 and b[34] n26621_not ; n27083
g26828 and n26619_not n27083 ; n27084
g26829 and n26623_not n27084_not ; n27085
g26830 and n27082_not n27085 ; n27086
g26831 and n26623_not n27086_not ; n27087
g26832 and b[35] n26612_not ; n27088
g26833 and n26610_not n27088 ; n27089
g26834 and n26614_not n27089_not ; n27090
g26835 and n27087_not n27090 ; n27091
g26836 and n26614_not n27091_not ; n27092
g26837 and b[36] n26603_not ; n27093
g26838 and n26601_not n27093 ; n27094
g26839 and n26605_not n27094_not ; n27095
g26840 and n27092_not n27095 ; n27096
g26841 and n26605_not n27096_not ; n27097
g26842 and b[37] n26594_not ; n27098
g26843 and n26592_not n27098 ; n27099
g26844 and n26596_not n27099_not ; n27100
g26845 and n27097_not n27100 ; n27101
g26846 and n26596_not n27101_not ; n27102
g26847 and b[38] n26585_not ; n27103
g26848 and n26583_not n27103 ; n27104
g26849 and n26587_not n27104_not ; n27105
g26850 and n27102_not n27105 ; n27106
g26851 and n26587_not n27106_not ; n27107
g26852 and b[39] n26576_not ; n27108
g26853 and n26574_not n27108 ; n27109
g26854 and n26578_not n27109_not ; n27110
g26855 and n27107_not n27110 ; n27111
g26856 and n26578_not n27111_not ; n27112
g26857 and b[40] n26567_not ; n27113
g26858 and n26565_not n27113 ; n27114
g26859 and n26569_not n27114_not ; n27115
g26860 and n27112_not n27115 ; n27116
g26861 and n26569_not n27116_not ; n27117
g26862 and b[41] n26558_not ; n27118
g26863 and n26556_not n27118 ; n27119
g26864 and n26560_not n27119_not ; n27120
g26865 and n27117_not n27120 ; n27121
g26866 and n26560_not n27121_not ; n27122
g26867 and b[42] n26549_not ; n27123
g26868 and n26547_not n27123 ; n27124
g26869 and n26551_not n27124_not ; n27125
g26870 and n27122_not n27125 ; n27126
g26871 and n26551_not n27126_not ; n27127
g26872 and b[43] n26540_not ; n27128
g26873 and n26538_not n27128 ; n27129
g26874 and n26542_not n27129_not ; n27130
g26875 and n27127_not n27130 ; n27131
g26876 and n26542_not n27131_not ; n27132
g26877 and b[44] n26531_not ; n27133
g26878 and n26529_not n27133 ; n27134
g26879 and n26533_not n27134_not ; n27135
g26880 and n27132_not n27135 ; n27136
g26881 and n26533_not n27136_not ; n27137
g26882 and b[45] n26522_not ; n27138
g26883 and n26520_not n27138 ; n27139
g26884 and n26524_not n27139_not ; n27140
g26885 and n27137_not n27140 ; n27141
g26886 and n26524_not n27141_not ; n27142
g26887 and b[46] n26513_not ; n27143
g26888 and n26511_not n27143 ; n27144
g26889 and n26515_not n27144_not ; n27145
g26890 and n27142_not n27145 ; n27146
g26891 and n26515_not n27146_not ; n27147
g26892 and b[47] n26504_not ; n27148
g26893 and n26502_not n27148 ; n27149
g26894 and n26506_not n27149_not ; n27150
g26895 and n27147_not n27150 ; n27151
g26896 and n26506_not n27151_not ; n27152
g26897 and b[48] n26495_not ; n27153
g26898 and n26493_not n27153 ; n27154
g26899 and n26497_not n27154_not ; n27155
g26900 and n27152_not n27155 ; n27156
g26901 and n26497_not n27156_not ; n27157
g26902 and b[49] n26486_not ; n27158
g26903 and n26484_not n27158 ; n27159
g26904 and n26488_not n27159_not ; n27160
g26905 and n27157_not n27160 ; n27161
g26906 and n26488_not n27161_not ; n27162
g26907 and b[50] n26477_not ; n27163
g26908 and n26475_not n27163 ; n27164
g26909 and n26479_not n27164_not ; n27165
g26910 and n27162_not n27165 ; n27166
g26911 and n26479_not n27166_not ; n27167
g26912 and b[51] n26468_not ; n27168
g26913 and n26466_not n27168 ; n27169
g26914 and n26470_not n27169_not ; n27170
g26915 and n27167_not n27170 ; n27171
g26916 and n26470_not n27171_not ; n27172
g26917 and b[52] n26459_not ; n27173
g26918 and n26457_not n27173 ; n27174
g26919 and n26461_not n27174_not ; n27175
g26920 and n27172_not n27175 ; n27176
g26921 and n26461_not n27176_not ; n27177
g26922 and b[53] n26450_not ; n27178
g26923 and n26448_not n27178 ; n27179
g26924 and n26452_not n27179_not ; n27180
g26925 and n27177_not n27180 ; n27181
g26926 and n26452_not n27181_not ; n27182
g26927 and b[54] n26441_not ; n27183
g26928 and n26439_not n27183 ; n27184
g26929 and n26443_not n27184_not ; n27185
g26930 and n27182_not n27185 ; n27186
g26931 and n26443_not n27186_not ; n27187
g26932 and b[55] n26432_not ; n27188
g26933 and n26430_not n27188 ; n27189
g26934 and n26434_not n27189_not ; n27190
g26935 and n27187_not n27190 ; n27191
g26936 and n26434_not n27191_not ; n27192
g26937 and b[56] n26423_not ; n27193
g26938 and n26421_not n27193 ; n27194
g26939 and n26425_not n27194_not ; n27195
g26940 and n27192_not n27195 ; n27196
g26941 and n26425_not n27196_not ; n27197
g26942 and b[57] n26414_not ; n27198
g26943 and n26412_not n27198 ; n27199
g26944 and n26416_not n27199_not ; n27200
g26945 and n27197_not n27200 ; n27201
g26946 and n26416_not n27201_not ; n27202
g26947 and b[58] n26405_not ; n27203
g26948 and n26403_not n27203 ; n27204
g26949 and n26407_not n27204_not ; n27205
g26950 and n27202_not n27205 ; n27206
g26951 and n26407_not n27206_not ; n27207
g26952 and b[59] n26396_not ; n27208
g26953 and n26394_not n27208 ; n27209
g26954 and n26398_not n27209_not ; n27210
g26955 and n27207_not n27210 ; n27211
g26956 and n26398_not n27211_not ; n27212
g26957 and b[60] n26387_not ; n27213
g26958 and n26385_not n27213 ; n27214
g26959 and n26389_not n27214_not ; n27215
g26960 and n27212_not n27215 ; n27216
g26961 and n26389_not n27216_not ; n27217
g26962 and n25548_not n26375_not ; n27218
g26963 and n26373_not n27218 ; n27219
g26964 and n26361_not n27219 ; n27220
g26965 and n26373_not n26375_not ; n27221
g26966 and n26362_not n27221_not ; n27222
g26967 and n27220_not n27222_not ; n27223
g26968 and quotient[3] n27223_not ; n27224
g26969 and n26372_not n26379_not ; n27225
g26970 and n26378_not n27225 ; n27226
g26971 and n27224_not n27226_not ; n27227
g26972 and b[61]_not n27227_not ; n27228
g26973 and b[61] n27226_not ; n27229
g26974 and n27224_not n27229 ; n27230
g26975 and n279 n27230_not ; n27231
g26976 and n27228_not n27231 ; n27232
g26977 and n27217_not n27232 ; n27233
g26978 and n403 n27227_not ; n27234
g26979 and n27233_not n27234_not ; quotient[2]
g26980 and n26398_not n27215 ; n27236
g26981 and n27211_not n27236 ; n27237
g26982 and n27212_not n27215_not ; n27238
g26983 and n27237_not n27238_not ; n27239
g26984 and quotient[2] n27239_not ; n27240
g26985 and n26388_not n27234_not ; n27241
g26986 and n27233_not n27241 ; n27242
g26987 and n27240_not n27242_not ; n27243
g26988 and b[61]_not n27243_not ; n27244
g26989 and n26407_not n27210 ; n27245
g26990 and n27206_not n27245 ; n27246
g26991 and n27207_not n27210_not ; n27247
g26992 and n27246_not n27247_not ; n27248
g26993 and quotient[2] n27248_not ; n27249
g26994 and n26397_not n27234_not ; n27250
g26995 and n27233_not n27250 ; n27251
g26996 and n27249_not n27251_not ; n27252
g26997 and b[60]_not n27252_not ; n27253
g26998 and n26416_not n27205 ; n27254
g26999 and n27201_not n27254 ; n27255
g27000 and n27202_not n27205_not ; n27256
g27001 and n27255_not n27256_not ; n27257
g27002 and quotient[2] n27257_not ; n27258
g27003 and n26406_not n27234_not ; n27259
g27004 and n27233_not n27259 ; n27260
g27005 and n27258_not n27260_not ; n27261
g27006 and b[59]_not n27261_not ; n27262
g27007 and n26425_not n27200 ; n27263
g27008 and n27196_not n27263 ; n27264
g27009 and n27197_not n27200_not ; n27265
g27010 and n27264_not n27265_not ; n27266
g27011 and quotient[2] n27266_not ; n27267
g27012 and n26415_not n27234_not ; n27268
g27013 and n27233_not n27268 ; n27269
g27014 and n27267_not n27269_not ; n27270
g27015 and b[58]_not n27270_not ; n27271
g27016 and n26434_not n27195 ; n27272
g27017 and n27191_not n27272 ; n27273
g27018 and n27192_not n27195_not ; n27274
g27019 and n27273_not n27274_not ; n27275
g27020 and quotient[2] n27275_not ; n27276
g27021 and n26424_not n27234_not ; n27277
g27022 and n27233_not n27277 ; n27278
g27023 and n27276_not n27278_not ; n27279
g27024 and b[57]_not n27279_not ; n27280
g27025 and n26443_not n27190 ; n27281
g27026 and n27186_not n27281 ; n27282
g27027 and n27187_not n27190_not ; n27283
g27028 and n27282_not n27283_not ; n27284
g27029 and quotient[2] n27284_not ; n27285
g27030 and n26433_not n27234_not ; n27286
g27031 and n27233_not n27286 ; n27287
g27032 and n27285_not n27287_not ; n27288
g27033 and b[56]_not n27288_not ; n27289
g27034 and n26452_not n27185 ; n27290
g27035 and n27181_not n27290 ; n27291
g27036 and n27182_not n27185_not ; n27292
g27037 and n27291_not n27292_not ; n27293
g27038 and quotient[2] n27293_not ; n27294
g27039 and n26442_not n27234_not ; n27295
g27040 and n27233_not n27295 ; n27296
g27041 and n27294_not n27296_not ; n27297
g27042 and b[55]_not n27297_not ; n27298
g27043 and n26461_not n27180 ; n27299
g27044 and n27176_not n27299 ; n27300
g27045 and n27177_not n27180_not ; n27301
g27046 and n27300_not n27301_not ; n27302
g27047 and quotient[2] n27302_not ; n27303
g27048 and n26451_not n27234_not ; n27304
g27049 and n27233_not n27304 ; n27305
g27050 and n27303_not n27305_not ; n27306
g27051 and b[54]_not n27306_not ; n27307
g27052 and n26470_not n27175 ; n27308
g27053 and n27171_not n27308 ; n27309
g27054 and n27172_not n27175_not ; n27310
g27055 and n27309_not n27310_not ; n27311
g27056 and quotient[2] n27311_not ; n27312
g27057 and n26460_not n27234_not ; n27313
g27058 and n27233_not n27313 ; n27314
g27059 and n27312_not n27314_not ; n27315
g27060 and b[53]_not n27315_not ; n27316
g27061 and n26479_not n27170 ; n27317
g27062 and n27166_not n27317 ; n27318
g27063 and n27167_not n27170_not ; n27319
g27064 and n27318_not n27319_not ; n27320
g27065 and quotient[2] n27320_not ; n27321
g27066 and n26469_not n27234_not ; n27322
g27067 and n27233_not n27322 ; n27323
g27068 and n27321_not n27323_not ; n27324
g27069 and b[52]_not n27324_not ; n27325
g27070 and n26488_not n27165 ; n27326
g27071 and n27161_not n27326 ; n27327
g27072 and n27162_not n27165_not ; n27328
g27073 and n27327_not n27328_not ; n27329
g27074 and quotient[2] n27329_not ; n27330
g27075 and n26478_not n27234_not ; n27331
g27076 and n27233_not n27331 ; n27332
g27077 and n27330_not n27332_not ; n27333
g27078 and b[51]_not n27333_not ; n27334
g27079 and n26497_not n27160 ; n27335
g27080 and n27156_not n27335 ; n27336
g27081 and n27157_not n27160_not ; n27337
g27082 and n27336_not n27337_not ; n27338
g27083 and quotient[2] n27338_not ; n27339
g27084 and n26487_not n27234_not ; n27340
g27085 and n27233_not n27340 ; n27341
g27086 and n27339_not n27341_not ; n27342
g27087 and b[50]_not n27342_not ; n27343
g27088 and n26506_not n27155 ; n27344
g27089 and n27151_not n27344 ; n27345
g27090 and n27152_not n27155_not ; n27346
g27091 and n27345_not n27346_not ; n27347
g27092 and quotient[2] n27347_not ; n27348
g27093 and n26496_not n27234_not ; n27349
g27094 and n27233_not n27349 ; n27350
g27095 and n27348_not n27350_not ; n27351
g27096 and b[49]_not n27351_not ; n27352
g27097 and n26515_not n27150 ; n27353
g27098 and n27146_not n27353 ; n27354
g27099 and n27147_not n27150_not ; n27355
g27100 and n27354_not n27355_not ; n27356
g27101 and quotient[2] n27356_not ; n27357
g27102 and n26505_not n27234_not ; n27358
g27103 and n27233_not n27358 ; n27359
g27104 and n27357_not n27359_not ; n27360
g27105 and b[48]_not n27360_not ; n27361
g27106 and n26524_not n27145 ; n27362
g27107 and n27141_not n27362 ; n27363
g27108 and n27142_not n27145_not ; n27364
g27109 and n27363_not n27364_not ; n27365
g27110 and quotient[2] n27365_not ; n27366
g27111 and n26514_not n27234_not ; n27367
g27112 and n27233_not n27367 ; n27368
g27113 and n27366_not n27368_not ; n27369
g27114 and b[47]_not n27369_not ; n27370
g27115 and n26533_not n27140 ; n27371
g27116 and n27136_not n27371 ; n27372
g27117 and n27137_not n27140_not ; n27373
g27118 and n27372_not n27373_not ; n27374
g27119 and quotient[2] n27374_not ; n27375
g27120 and n26523_not n27234_not ; n27376
g27121 and n27233_not n27376 ; n27377
g27122 and n27375_not n27377_not ; n27378
g27123 and b[46]_not n27378_not ; n27379
g27124 and n26542_not n27135 ; n27380
g27125 and n27131_not n27380 ; n27381
g27126 and n27132_not n27135_not ; n27382
g27127 and n27381_not n27382_not ; n27383
g27128 and quotient[2] n27383_not ; n27384
g27129 and n26532_not n27234_not ; n27385
g27130 and n27233_not n27385 ; n27386
g27131 and n27384_not n27386_not ; n27387
g27132 and b[45]_not n27387_not ; n27388
g27133 and n26551_not n27130 ; n27389
g27134 and n27126_not n27389 ; n27390
g27135 and n27127_not n27130_not ; n27391
g27136 and n27390_not n27391_not ; n27392
g27137 and quotient[2] n27392_not ; n27393
g27138 and n26541_not n27234_not ; n27394
g27139 and n27233_not n27394 ; n27395
g27140 and n27393_not n27395_not ; n27396
g27141 and b[44]_not n27396_not ; n27397
g27142 and n26560_not n27125 ; n27398
g27143 and n27121_not n27398 ; n27399
g27144 and n27122_not n27125_not ; n27400
g27145 and n27399_not n27400_not ; n27401
g27146 and quotient[2] n27401_not ; n27402
g27147 and n26550_not n27234_not ; n27403
g27148 and n27233_not n27403 ; n27404
g27149 and n27402_not n27404_not ; n27405
g27150 and b[43]_not n27405_not ; n27406
g27151 and n26569_not n27120 ; n27407
g27152 and n27116_not n27407 ; n27408
g27153 and n27117_not n27120_not ; n27409
g27154 and n27408_not n27409_not ; n27410
g27155 and quotient[2] n27410_not ; n27411
g27156 and n26559_not n27234_not ; n27412
g27157 and n27233_not n27412 ; n27413
g27158 and n27411_not n27413_not ; n27414
g27159 and b[42]_not n27414_not ; n27415
g27160 and n26578_not n27115 ; n27416
g27161 and n27111_not n27416 ; n27417
g27162 and n27112_not n27115_not ; n27418
g27163 and n27417_not n27418_not ; n27419
g27164 and quotient[2] n27419_not ; n27420
g27165 and n26568_not n27234_not ; n27421
g27166 and n27233_not n27421 ; n27422
g27167 and n27420_not n27422_not ; n27423
g27168 and b[41]_not n27423_not ; n27424
g27169 and n26587_not n27110 ; n27425
g27170 and n27106_not n27425 ; n27426
g27171 and n27107_not n27110_not ; n27427
g27172 and n27426_not n27427_not ; n27428
g27173 and quotient[2] n27428_not ; n27429
g27174 and n26577_not n27234_not ; n27430
g27175 and n27233_not n27430 ; n27431
g27176 and n27429_not n27431_not ; n27432
g27177 and b[40]_not n27432_not ; n27433
g27178 and n26596_not n27105 ; n27434
g27179 and n27101_not n27434 ; n27435
g27180 and n27102_not n27105_not ; n27436
g27181 and n27435_not n27436_not ; n27437
g27182 and quotient[2] n27437_not ; n27438
g27183 and n26586_not n27234_not ; n27439
g27184 and n27233_not n27439 ; n27440
g27185 and n27438_not n27440_not ; n27441
g27186 and b[39]_not n27441_not ; n27442
g27187 and n26605_not n27100 ; n27443
g27188 and n27096_not n27443 ; n27444
g27189 and n27097_not n27100_not ; n27445
g27190 and n27444_not n27445_not ; n27446
g27191 and quotient[2] n27446_not ; n27447
g27192 and n26595_not n27234_not ; n27448
g27193 and n27233_not n27448 ; n27449
g27194 and n27447_not n27449_not ; n27450
g27195 and b[38]_not n27450_not ; n27451
g27196 and n26614_not n27095 ; n27452
g27197 and n27091_not n27452 ; n27453
g27198 and n27092_not n27095_not ; n27454
g27199 and n27453_not n27454_not ; n27455
g27200 and quotient[2] n27455_not ; n27456
g27201 and n26604_not n27234_not ; n27457
g27202 and n27233_not n27457 ; n27458
g27203 and n27456_not n27458_not ; n27459
g27204 and b[37]_not n27459_not ; n27460
g27205 and n26623_not n27090 ; n27461
g27206 and n27086_not n27461 ; n27462
g27207 and n27087_not n27090_not ; n27463
g27208 and n27462_not n27463_not ; n27464
g27209 and quotient[2] n27464_not ; n27465
g27210 and n26613_not n27234_not ; n27466
g27211 and n27233_not n27466 ; n27467
g27212 and n27465_not n27467_not ; n27468
g27213 and b[36]_not n27468_not ; n27469
g27214 and n26632_not n27085 ; n27470
g27215 and n27081_not n27470 ; n27471
g27216 and n27082_not n27085_not ; n27472
g27217 and n27471_not n27472_not ; n27473
g27218 and quotient[2] n27473_not ; n27474
g27219 and n26622_not n27234_not ; n27475
g27220 and n27233_not n27475 ; n27476
g27221 and n27474_not n27476_not ; n27477
g27222 and b[35]_not n27477_not ; n27478
g27223 and n26641_not n27080 ; n27479
g27224 and n27076_not n27479 ; n27480
g27225 and n27077_not n27080_not ; n27481
g27226 and n27480_not n27481_not ; n27482
g27227 and quotient[2] n27482_not ; n27483
g27228 and n26631_not n27234_not ; n27484
g27229 and n27233_not n27484 ; n27485
g27230 and n27483_not n27485_not ; n27486
g27231 and b[34]_not n27486_not ; n27487
g27232 and n26650_not n27075 ; n27488
g27233 and n27071_not n27488 ; n27489
g27234 and n27072_not n27075_not ; n27490
g27235 and n27489_not n27490_not ; n27491
g27236 and quotient[2] n27491_not ; n27492
g27237 and n26640_not n27234_not ; n27493
g27238 and n27233_not n27493 ; n27494
g27239 and n27492_not n27494_not ; n27495
g27240 and b[33]_not n27495_not ; n27496
g27241 and n26659_not n27070 ; n27497
g27242 and n27066_not n27497 ; n27498
g27243 and n27067_not n27070_not ; n27499
g27244 and n27498_not n27499_not ; n27500
g27245 and quotient[2] n27500_not ; n27501
g27246 and n26649_not n27234_not ; n27502
g27247 and n27233_not n27502 ; n27503
g27248 and n27501_not n27503_not ; n27504
g27249 and b[32]_not n27504_not ; n27505
g27250 and n26668_not n27065 ; n27506
g27251 and n27061_not n27506 ; n27507
g27252 and n27062_not n27065_not ; n27508
g27253 and n27507_not n27508_not ; n27509
g27254 and quotient[2] n27509_not ; n27510
g27255 and n26658_not n27234_not ; n27511
g27256 and n27233_not n27511 ; n27512
g27257 and n27510_not n27512_not ; n27513
g27258 and b[31]_not n27513_not ; n27514
g27259 and n26677_not n27060 ; n27515
g27260 and n27056_not n27515 ; n27516
g27261 and n27057_not n27060_not ; n27517
g27262 and n27516_not n27517_not ; n27518
g27263 and quotient[2] n27518_not ; n27519
g27264 and n26667_not n27234_not ; n27520
g27265 and n27233_not n27520 ; n27521
g27266 and n27519_not n27521_not ; n27522
g27267 and b[30]_not n27522_not ; n27523
g27268 and n26686_not n27055 ; n27524
g27269 and n27051_not n27524 ; n27525
g27270 and n27052_not n27055_not ; n27526
g27271 and n27525_not n27526_not ; n27527
g27272 and quotient[2] n27527_not ; n27528
g27273 and n26676_not n27234_not ; n27529
g27274 and n27233_not n27529 ; n27530
g27275 and n27528_not n27530_not ; n27531
g27276 and b[29]_not n27531_not ; n27532
g27277 and n26695_not n27050 ; n27533
g27278 and n27046_not n27533 ; n27534
g27279 and n27047_not n27050_not ; n27535
g27280 and n27534_not n27535_not ; n27536
g27281 and quotient[2] n27536_not ; n27537
g27282 and n26685_not n27234_not ; n27538
g27283 and n27233_not n27538 ; n27539
g27284 and n27537_not n27539_not ; n27540
g27285 and b[28]_not n27540_not ; n27541
g27286 and n26704_not n27045 ; n27542
g27287 and n27041_not n27542 ; n27543
g27288 and n27042_not n27045_not ; n27544
g27289 and n27543_not n27544_not ; n27545
g27290 and quotient[2] n27545_not ; n27546
g27291 and n26694_not n27234_not ; n27547
g27292 and n27233_not n27547 ; n27548
g27293 and n27546_not n27548_not ; n27549
g27294 and b[27]_not n27549_not ; n27550
g27295 and n26713_not n27040 ; n27551
g27296 and n27036_not n27551 ; n27552
g27297 and n27037_not n27040_not ; n27553
g27298 and n27552_not n27553_not ; n27554
g27299 and quotient[2] n27554_not ; n27555
g27300 and n26703_not n27234_not ; n27556
g27301 and n27233_not n27556 ; n27557
g27302 and n27555_not n27557_not ; n27558
g27303 and b[26]_not n27558_not ; n27559
g27304 and n26722_not n27035 ; n27560
g27305 and n27031_not n27560 ; n27561
g27306 and n27032_not n27035_not ; n27562
g27307 and n27561_not n27562_not ; n27563
g27308 and quotient[2] n27563_not ; n27564
g27309 and n26712_not n27234_not ; n27565
g27310 and n27233_not n27565 ; n27566
g27311 and n27564_not n27566_not ; n27567
g27312 and b[25]_not n27567_not ; n27568
g27313 and n26731_not n27030 ; n27569
g27314 and n27026_not n27569 ; n27570
g27315 and n27027_not n27030_not ; n27571
g27316 and n27570_not n27571_not ; n27572
g27317 and quotient[2] n27572_not ; n27573
g27318 and n26721_not n27234_not ; n27574
g27319 and n27233_not n27574 ; n27575
g27320 and n27573_not n27575_not ; n27576
g27321 and b[24]_not n27576_not ; n27577
g27322 and n26740_not n27025 ; n27578
g27323 and n27021_not n27578 ; n27579
g27324 and n27022_not n27025_not ; n27580
g27325 and n27579_not n27580_not ; n27581
g27326 and quotient[2] n27581_not ; n27582
g27327 and n26730_not n27234_not ; n27583
g27328 and n27233_not n27583 ; n27584
g27329 and n27582_not n27584_not ; n27585
g27330 and b[23]_not n27585_not ; n27586
g27331 and n26749_not n27020 ; n27587
g27332 and n27016_not n27587 ; n27588
g27333 and n27017_not n27020_not ; n27589
g27334 and n27588_not n27589_not ; n27590
g27335 and quotient[2] n27590_not ; n27591
g27336 and n26739_not n27234_not ; n27592
g27337 and n27233_not n27592 ; n27593
g27338 and n27591_not n27593_not ; n27594
g27339 and b[22]_not n27594_not ; n27595
g27340 and n26758_not n27015 ; n27596
g27341 and n27011_not n27596 ; n27597
g27342 and n27012_not n27015_not ; n27598
g27343 and n27597_not n27598_not ; n27599
g27344 and quotient[2] n27599_not ; n27600
g27345 and n26748_not n27234_not ; n27601
g27346 and n27233_not n27601 ; n27602
g27347 and n27600_not n27602_not ; n27603
g27348 and b[21]_not n27603_not ; n27604
g27349 and n26767_not n27010 ; n27605
g27350 and n27006_not n27605 ; n27606
g27351 and n27007_not n27010_not ; n27607
g27352 and n27606_not n27607_not ; n27608
g27353 and quotient[2] n27608_not ; n27609
g27354 and n26757_not n27234_not ; n27610
g27355 and n27233_not n27610 ; n27611
g27356 and n27609_not n27611_not ; n27612
g27357 and b[20]_not n27612_not ; n27613
g27358 and n26776_not n27005 ; n27614
g27359 and n27001_not n27614 ; n27615
g27360 and n27002_not n27005_not ; n27616
g27361 and n27615_not n27616_not ; n27617
g27362 and quotient[2] n27617_not ; n27618
g27363 and n26766_not n27234_not ; n27619
g27364 and n27233_not n27619 ; n27620
g27365 and n27618_not n27620_not ; n27621
g27366 and b[19]_not n27621_not ; n27622
g27367 and n26785_not n27000 ; n27623
g27368 and n26996_not n27623 ; n27624
g27369 and n26997_not n27000_not ; n27625
g27370 and n27624_not n27625_not ; n27626
g27371 and quotient[2] n27626_not ; n27627
g27372 and n26775_not n27234_not ; n27628
g27373 and n27233_not n27628 ; n27629
g27374 and n27627_not n27629_not ; n27630
g27375 and b[18]_not n27630_not ; n27631
g27376 and n26794_not n26995 ; n27632
g27377 and n26991_not n27632 ; n27633
g27378 and n26992_not n26995_not ; n27634
g27379 and n27633_not n27634_not ; n27635
g27380 and quotient[2] n27635_not ; n27636
g27381 and n26784_not n27234_not ; n27637
g27382 and n27233_not n27637 ; n27638
g27383 and n27636_not n27638_not ; n27639
g27384 and b[17]_not n27639_not ; n27640
g27385 and n26803_not n26990 ; n27641
g27386 and n26986_not n27641 ; n27642
g27387 and n26987_not n26990_not ; n27643
g27388 and n27642_not n27643_not ; n27644
g27389 and quotient[2] n27644_not ; n27645
g27390 and n26793_not n27234_not ; n27646
g27391 and n27233_not n27646 ; n27647
g27392 and n27645_not n27647_not ; n27648
g27393 and b[16]_not n27648_not ; n27649
g27394 and n26812_not n26985 ; n27650
g27395 and n26981_not n27650 ; n27651
g27396 and n26982_not n26985_not ; n27652
g27397 and n27651_not n27652_not ; n27653
g27398 and quotient[2] n27653_not ; n27654
g27399 and n26802_not n27234_not ; n27655
g27400 and n27233_not n27655 ; n27656
g27401 and n27654_not n27656_not ; n27657
g27402 and b[15]_not n27657_not ; n27658
g27403 and n26821_not n26980 ; n27659
g27404 and n26976_not n27659 ; n27660
g27405 and n26977_not n26980_not ; n27661
g27406 and n27660_not n27661_not ; n27662
g27407 and quotient[2] n27662_not ; n27663
g27408 and n26811_not n27234_not ; n27664
g27409 and n27233_not n27664 ; n27665
g27410 and n27663_not n27665_not ; n27666
g27411 and b[14]_not n27666_not ; n27667
g27412 and n26830_not n26975 ; n27668
g27413 and n26971_not n27668 ; n27669
g27414 and n26972_not n26975_not ; n27670
g27415 and n27669_not n27670_not ; n27671
g27416 and quotient[2] n27671_not ; n27672
g27417 and n26820_not n27234_not ; n27673
g27418 and n27233_not n27673 ; n27674
g27419 and n27672_not n27674_not ; n27675
g27420 and b[13]_not n27675_not ; n27676
g27421 and n26839_not n26970 ; n27677
g27422 and n26966_not n27677 ; n27678
g27423 and n26967_not n26970_not ; n27679
g27424 and n27678_not n27679_not ; n27680
g27425 and quotient[2] n27680_not ; n27681
g27426 and n26829_not n27234_not ; n27682
g27427 and n27233_not n27682 ; n27683
g27428 and n27681_not n27683_not ; n27684
g27429 and b[12]_not n27684_not ; n27685
g27430 and n26848_not n26965 ; n27686
g27431 and n26961_not n27686 ; n27687
g27432 and n26962_not n26965_not ; n27688
g27433 and n27687_not n27688_not ; n27689
g27434 and quotient[2] n27689_not ; n27690
g27435 and n26838_not n27234_not ; n27691
g27436 and n27233_not n27691 ; n27692
g27437 and n27690_not n27692_not ; n27693
g27438 and b[11]_not n27693_not ; n27694
g27439 and n26857_not n26960 ; n27695
g27440 and n26956_not n27695 ; n27696
g27441 and n26957_not n26960_not ; n27697
g27442 and n27696_not n27697_not ; n27698
g27443 and quotient[2] n27698_not ; n27699
g27444 and n26847_not n27234_not ; n27700
g27445 and n27233_not n27700 ; n27701
g27446 and n27699_not n27701_not ; n27702
g27447 and b[10]_not n27702_not ; n27703
g27448 and n26866_not n26955 ; n27704
g27449 and n26951_not n27704 ; n27705
g27450 and n26952_not n26955_not ; n27706
g27451 and n27705_not n27706_not ; n27707
g27452 and quotient[2] n27707_not ; n27708
g27453 and n26856_not n27234_not ; n27709
g27454 and n27233_not n27709 ; n27710
g27455 and n27708_not n27710_not ; n27711
g27456 and b[9]_not n27711_not ; n27712
g27457 and n26875_not n26950 ; n27713
g27458 and n26946_not n27713 ; n27714
g27459 and n26947_not n26950_not ; n27715
g27460 and n27714_not n27715_not ; n27716
g27461 and quotient[2] n27716_not ; n27717
g27462 and n26865_not n27234_not ; n27718
g27463 and n27233_not n27718 ; n27719
g27464 and n27717_not n27719_not ; n27720
g27465 and b[8]_not n27720_not ; n27721
g27466 and n26884_not n26945 ; n27722
g27467 and n26941_not n27722 ; n27723
g27468 and n26942_not n26945_not ; n27724
g27469 and n27723_not n27724_not ; n27725
g27470 and quotient[2] n27725_not ; n27726
g27471 and n26874_not n27234_not ; n27727
g27472 and n27233_not n27727 ; n27728
g27473 and n27726_not n27728_not ; n27729
g27474 and b[7]_not n27729_not ; n27730
g27475 and n26893_not n26940 ; n27731
g27476 and n26936_not n27731 ; n27732
g27477 and n26937_not n26940_not ; n27733
g27478 and n27732_not n27733_not ; n27734
g27479 and quotient[2] n27734_not ; n27735
g27480 and n26883_not n27234_not ; n27736
g27481 and n27233_not n27736 ; n27737
g27482 and n27735_not n27737_not ; n27738
g27483 and b[6]_not n27738_not ; n27739
g27484 and n26902_not n26935 ; n27740
g27485 and n26931_not n27740 ; n27741
g27486 and n26932_not n26935_not ; n27742
g27487 and n27741_not n27742_not ; n27743
g27488 and quotient[2] n27743_not ; n27744
g27489 and n26892_not n27234_not ; n27745
g27490 and n27233_not n27745 ; n27746
g27491 and n27744_not n27746_not ; n27747
g27492 and b[5]_not n27747_not ; n27748
g27493 and n26910_not n26930 ; n27749
g27494 and n26926_not n27749 ; n27750
g27495 and n26927_not n26930_not ; n27751
g27496 and n27750_not n27751_not ; n27752
g27497 and quotient[2] n27752_not ; n27753
g27498 and n26901_not n27234_not ; n27754
g27499 and n27233_not n27754 ; n27755
g27500 and n27753_not n27755_not ; n27756
g27501 and b[4]_not n27756_not ; n27757
g27502 and n26921_not n26925 ; n27758
g27503 and n26920_not n27758 ; n27759
g27504 and n26922_not n26925_not ; n27760
g27505 and n27759_not n27760_not ; n27761
g27506 and quotient[2] n27761_not ; n27762
g27507 and n26909_not n27234_not ; n27763
g27508 and n27233_not n27763 ; n27764
g27509 and n27762_not n27764_not ; n27765
g27510 and b[3]_not n27765_not ; n27766
g27511 and n26917_not n26919 ; n27767
g27512 and n26915_not n27767 ; n27768
g27513 and n26920_not n27768_not ; n27769
g27514 and quotient[2] n27769 ; n27770
g27515 and n26914_not n27234_not ; n27771
g27516 and n27233_not n27771 ; n27772
g27517 and n27770_not n27772_not ; n27773
g27518 and b[2]_not n27773_not ; n27774
g27519 and b[0] quotient[2] ; n27775
g27520 and a[2] n27775_not ; n27776
g27521 and n26919 quotient[2] ; n27777
g27522 and n27776_not n27777_not ; n27778
g27523 and b[1] n27778_not ; n27779
g27524 and b[1]_not n27777_not ; n27780
g27525 and n27776_not n27780 ; n27781
g27526 and n27779_not n27781_not ; n27782
g27527 and a[1]_not b[0] ; n27783
g27528 and n27782_not n27783_not ; n27784
g27529 and b[1]_not n27778_not ; n27785
g27530 and n27784_not n27785_not ; n27786
g27531 and b[2] n27772_not ; n27787
g27532 and n27770_not n27787 ; n27788
g27533 and n27774_not n27788_not ; n27789
g27534 and n27786_not n27789 ; n27790
g27535 and n27774_not n27790_not ; n27791
g27536 and b[3] n27764_not ; n27792
g27537 and n27762_not n27792 ; n27793
g27538 and n27766_not n27793_not ; n27794
g27539 and n27791_not n27794 ; n27795
g27540 and n27766_not n27795_not ; n27796
g27541 and b[4] n27755_not ; n27797
g27542 and n27753_not n27797 ; n27798
g27543 and n27757_not n27798_not ; n27799
g27544 and n27796_not n27799 ; n27800
g27545 and n27757_not n27800_not ; n27801
g27546 and b[5] n27746_not ; n27802
g27547 and n27744_not n27802 ; n27803
g27548 and n27748_not n27803_not ; n27804
g27549 and n27801_not n27804 ; n27805
g27550 and n27748_not n27805_not ; n27806
g27551 and b[6] n27737_not ; n27807
g27552 and n27735_not n27807 ; n27808
g27553 and n27739_not n27808_not ; n27809
g27554 and n27806_not n27809 ; n27810
g27555 and n27739_not n27810_not ; n27811
g27556 and b[7] n27728_not ; n27812
g27557 and n27726_not n27812 ; n27813
g27558 and n27730_not n27813_not ; n27814
g27559 and n27811_not n27814 ; n27815
g27560 and n27730_not n27815_not ; n27816
g27561 and b[8] n27719_not ; n27817
g27562 and n27717_not n27817 ; n27818
g27563 and n27721_not n27818_not ; n27819
g27564 and n27816_not n27819 ; n27820
g27565 and n27721_not n27820_not ; n27821
g27566 and b[9] n27710_not ; n27822
g27567 and n27708_not n27822 ; n27823
g27568 and n27712_not n27823_not ; n27824
g27569 and n27821_not n27824 ; n27825
g27570 and n27712_not n27825_not ; n27826
g27571 and b[10] n27701_not ; n27827
g27572 and n27699_not n27827 ; n27828
g27573 and n27703_not n27828_not ; n27829
g27574 and n27826_not n27829 ; n27830
g27575 and n27703_not n27830_not ; n27831
g27576 and b[11] n27692_not ; n27832
g27577 and n27690_not n27832 ; n27833
g27578 and n27694_not n27833_not ; n27834
g27579 and n27831_not n27834 ; n27835
g27580 and n27694_not n27835_not ; n27836
g27581 and b[12] n27683_not ; n27837
g27582 and n27681_not n27837 ; n27838
g27583 and n27685_not n27838_not ; n27839
g27584 and n27836_not n27839 ; n27840
g27585 and n27685_not n27840_not ; n27841
g27586 and b[13] n27674_not ; n27842
g27587 and n27672_not n27842 ; n27843
g27588 and n27676_not n27843_not ; n27844
g27589 and n27841_not n27844 ; n27845
g27590 and n27676_not n27845_not ; n27846
g27591 and b[14] n27665_not ; n27847
g27592 and n27663_not n27847 ; n27848
g27593 and n27667_not n27848_not ; n27849
g27594 and n27846_not n27849 ; n27850
g27595 and n27667_not n27850_not ; n27851
g27596 and b[15] n27656_not ; n27852
g27597 and n27654_not n27852 ; n27853
g27598 and n27658_not n27853_not ; n27854
g27599 and n27851_not n27854 ; n27855
g27600 and n27658_not n27855_not ; n27856
g27601 and b[16] n27647_not ; n27857
g27602 and n27645_not n27857 ; n27858
g27603 and n27649_not n27858_not ; n27859
g27604 and n27856_not n27859 ; n27860
g27605 and n27649_not n27860_not ; n27861
g27606 and b[17] n27638_not ; n27862
g27607 and n27636_not n27862 ; n27863
g27608 and n27640_not n27863_not ; n27864
g27609 and n27861_not n27864 ; n27865
g27610 and n27640_not n27865_not ; n27866
g27611 and b[18] n27629_not ; n27867
g27612 and n27627_not n27867 ; n27868
g27613 and n27631_not n27868_not ; n27869
g27614 and n27866_not n27869 ; n27870
g27615 and n27631_not n27870_not ; n27871
g27616 and b[19] n27620_not ; n27872
g27617 and n27618_not n27872 ; n27873
g27618 and n27622_not n27873_not ; n27874
g27619 and n27871_not n27874 ; n27875
g27620 and n27622_not n27875_not ; n27876
g27621 and b[20] n27611_not ; n27877
g27622 and n27609_not n27877 ; n27878
g27623 and n27613_not n27878_not ; n27879
g27624 and n27876_not n27879 ; n27880
g27625 and n27613_not n27880_not ; n27881
g27626 and b[21] n27602_not ; n27882
g27627 and n27600_not n27882 ; n27883
g27628 and n27604_not n27883_not ; n27884
g27629 and n27881_not n27884 ; n27885
g27630 and n27604_not n27885_not ; n27886
g27631 and b[22] n27593_not ; n27887
g27632 and n27591_not n27887 ; n27888
g27633 and n27595_not n27888_not ; n27889
g27634 and n27886_not n27889 ; n27890
g27635 and n27595_not n27890_not ; n27891
g27636 and b[23] n27584_not ; n27892
g27637 and n27582_not n27892 ; n27893
g27638 and n27586_not n27893_not ; n27894
g27639 and n27891_not n27894 ; n27895
g27640 and n27586_not n27895_not ; n27896
g27641 and b[24] n27575_not ; n27897
g27642 and n27573_not n27897 ; n27898
g27643 and n27577_not n27898_not ; n27899
g27644 and n27896_not n27899 ; n27900
g27645 and n27577_not n27900_not ; n27901
g27646 and b[25] n27566_not ; n27902
g27647 and n27564_not n27902 ; n27903
g27648 and n27568_not n27903_not ; n27904
g27649 and n27901_not n27904 ; n27905
g27650 and n27568_not n27905_not ; n27906
g27651 and b[26] n27557_not ; n27907
g27652 and n27555_not n27907 ; n27908
g27653 and n27559_not n27908_not ; n27909
g27654 and n27906_not n27909 ; n27910
g27655 and n27559_not n27910_not ; n27911
g27656 and b[27] n27548_not ; n27912
g27657 and n27546_not n27912 ; n27913
g27658 and n27550_not n27913_not ; n27914
g27659 and n27911_not n27914 ; n27915
g27660 and n27550_not n27915_not ; n27916
g27661 and b[28] n27539_not ; n27917
g27662 and n27537_not n27917 ; n27918
g27663 and n27541_not n27918_not ; n27919
g27664 and n27916_not n27919 ; n27920
g27665 and n27541_not n27920_not ; n27921
g27666 and b[29] n27530_not ; n27922
g27667 and n27528_not n27922 ; n27923
g27668 and n27532_not n27923_not ; n27924
g27669 and n27921_not n27924 ; n27925
g27670 and n27532_not n27925_not ; n27926
g27671 and b[30] n27521_not ; n27927
g27672 and n27519_not n27927 ; n27928
g27673 and n27523_not n27928_not ; n27929
g27674 and n27926_not n27929 ; n27930
g27675 and n27523_not n27930_not ; n27931
g27676 and b[31] n27512_not ; n27932
g27677 and n27510_not n27932 ; n27933
g27678 and n27514_not n27933_not ; n27934
g27679 and n27931_not n27934 ; n27935
g27680 and n27514_not n27935_not ; n27936
g27681 and b[32] n27503_not ; n27937
g27682 and n27501_not n27937 ; n27938
g27683 and n27505_not n27938_not ; n27939
g27684 and n27936_not n27939 ; n27940
g27685 and n27505_not n27940_not ; n27941
g27686 and b[33] n27494_not ; n27942
g27687 and n27492_not n27942 ; n27943
g27688 and n27496_not n27943_not ; n27944
g27689 and n27941_not n27944 ; n27945
g27690 and n27496_not n27945_not ; n27946
g27691 and b[34] n27485_not ; n27947
g27692 and n27483_not n27947 ; n27948
g27693 and n27487_not n27948_not ; n27949
g27694 and n27946_not n27949 ; n27950
g27695 and n27487_not n27950_not ; n27951
g27696 and b[35] n27476_not ; n27952
g27697 and n27474_not n27952 ; n27953
g27698 and n27478_not n27953_not ; n27954
g27699 and n27951_not n27954 ; n27955
g27700 and n27478_not n27955_not ; n27956
g27701 and b[36] n27467_not ; n27957
g27702 and n27465_not n27957 ; n27958
g27703 and n27469_not n27958_not ; n27959
g27704 and n27956_not n27959 ; n27960
g27705 and n27469_not n27960_not ; n27961
g27706 and b[37] n27458_not ; n27962
g27707 and n27456_not n27962 ; n27963
g27708 and n27460_not n27963_not ; n27964
g27709 and n27961_not n27964 ; n27965
g27710 and n27460_not n27965_not ; n27966
g27711 and b[38] n27449_not ; n27967
g27712 and n27447_not n27967 ; n27968
g27713 and n27451_not n27968_not ; n27969
g27714 and n27966_not n27969 ; n27970
g27715 and n27451_not n27970_not ; n27971
g27716 and b[39] n27440_not ; n27972
g27717 and n27438_not n27972 ; n27973
g27718 and n27442_not n27973_not ; n27974
g27719 and n27971_not n27974 ; n27975
g27720 and n27442_not n27975_not ; n27976
g27721 and b[40] n27431_not ; n27977
g27722 and n27429_not n27977 ; n27978
g27723 and n27433_not n27978_not ; n27979
g27724 and n27976_not n27979 ; n27980
g27725 and n27433_not n27980_not ; n27981
g27726 and b[41] n27422_not ; n27982
g27727 and n27420_not n27982 ; n27983
g27728 and n27424_not n27983_not ; n27984
g27729 and n27981_not n27984 ; n27985
g27730 and n27424_not n27985_not ; n27986
g27731 and b[42] n27413_not ; n27987
g27732 and n27411_not n27987 ; n27988
g27733 and n27415_not n27988_not ; n27989
g27734 and n27986_not n27989 ; n27990
g27735 and n27415_not n27990_not ; n27991
g27736 and b[43] n27404_not ; n27992
g27737 and n27402_not n27992 ; n27993
g27738 and n27406_not n27993_not ; n27994
g27739 and n27991_not n27994 ; n27995
g27740 and n27406_not n27995_not ; n27996
g27741 and b[44] n27395_not ; n27997
g27742 and n27393_not n27997 ; n27998
g27743 and n27397_not n27998_not ; n27999
g27744 and n27996_not n27999 ; n28000
g27745 and n27397_not n28000_not ; n28001
g27746 and b[45] n27386_not ; n28002
g27747 and n27384_not n28002 ; n28003
g27748 and n27388_not n28003_not ; n28004
g27749 and n28001_not n28004 ; n28005
g27750 and n27388_not n28005_not ; n28006
g27751 and b[46] n27377_not ; n28007
g27752 and n27375_not n28007 ; n28008
g27753 and n27379_not n28008_not ; n28009
g27754 and n28006_not n28009 ; n28010
g27755 and n27379_not n28010_not ; n28011
g27756 and b[47] n27368_not ; n28012
g27757 and n27366_not n28012 ; n28013
g27758 and n27370_not n28013_not ; n28014
g27759 and n28011_not n28014 ; n28015
g27760 and n27370_not n28015_not ; n28016
g27761 and b[48] n27359_not ; n28017
g27762 and n27357_not n28017 ; n28018
g27763 and n27361_not n28018_not ; n28019
g27764 and n28016_not n28019 ; n28020
g27765 and n27361_not n28020_not ; n28021
g27766 and b[49] n27350_not ; n28022
g27767 and n27348_not n28022 ; n28023
g27768 and n27352_not n28023_not ; n28024
g27769 and n28021_not n28024 ; n28025
g27770 and n27352_not n28025_not ; n28026
g27771 and b[50] n27341_not ; n28027
g27772 and n27339_not n28027 ; n28028
g27773 and n27343_not n28028_not ; n28029
g27774 and n28026_not n28029 ; n28030
g27775 and n27343_not n28030_not ; n28031
g27776 and b[51] n27332_not ; n28032
g27777 and n27330_not n28032 ; n28033
g27778 and n27334_not n28033_not ; n28034
g27779 and n28031_not n28034 ; n28035
g27780 and n27334_not n28035_not ; n28036
g27781 and b[52] n27323_not ; n28037
g27782 and n27321_not n28037 ; n28038
g27783 and n27325_not n28038_not ; n28039
g27784 and n28036_not n28039 ; n28040
g27785 and n27325_not n28040_not ; n28041
g27786 and b[53] n27314_not ; n28042
g27787 and n27312_not n28042 ; n28043
g27788 and n27316_not n28043_not ; n28044
g27789 and n28041_not n28044 ; n28045
g27790 and n27316_not n28045_not ; n28046
g27791 and b[54] n27305_not ; n28047
g27792 and n27303_not n28047 ; n28048
g27793 and n27307_not n28048_not ; n28049
g27794 and n28046_not n28049 ; n28050
g27795 and n27307_not n28050_not ; n28051
g27796 and b[55] n27296_not ; n28052
g27797 and n27294_not n28052 ; n28053
g27798 and n27298_not n28053_not ; n28054
g27799 and n28051_not n28054 ; n28055
g27800 and n27298_not n28055_not ; n28056
g27801 and b[56] n27287_not ; n28057
g27802 and n27285_not n28057 ; n28058
g27803 and n27289_not n28058_not ; n28059
g27804 and n28056_not n28059 ; n28060
g27805 and n27289_not n28060_not ; n28061
g27806 and b[57] n27278_not ; n28062
g27807 and n27276_not n28062 ; n28063
g27808 and n27280_not n28063_not ; n28064
g27809 and n28061_not n28064 ; n28065
g27810 and n27280_not n28065_not ; n28066
g27811 and b[58] n27269_not ; n28067
g27812 and n27267_not n28067 ; n28068
g27813 and n27271_not n28068_not ; n28069
g27814 and n28066_not n28069 ; n28070
g27815 and n27271_not n28070_not ; n28071
g27816 and b[59] n27260_not ; n28072
g27817 and n27258_not n28072 ; n28073
g27818 and n27262_not n28073_not ; n28074
g27819 and n28071_not n28074 ; n28075
g27820 and n27262_not n28075_not ; n28076
g27821 and b[60] n27251_not ; n28077
g27822 and n27249_not n28077 ; n28078
g27823 and n27253_not n28078_not ; n28079
g27824 and n28076_not n28079 ; n28080
g27825 and n27253_not n28080_not ; n28081
g27826 and b[61] n27242_not ; n28082
g27827 and n27240_not n28082 ; n28083
g27828 and n27244_not n28083_not ; n28084
g27829 and n28081_not n28084 ; n28085
g27830 and n27244_not n28085_not ; n28086
g27831 and n26389_not n27230_not ; n28087
g27832 and n27228_not n28087 ; n28088
g27833 and n27216_not n28088 ; n28089
g27834 and n27228_not n27230_not ; n28090
g27835 and n27217_not n28090_not ; n28091
g27836 and n28089_not n28091_not ; n28092
g27837 and quotient[2] n28092_not ; n28093
g27838 and n27227_not n27234_not ; n28094
g27839 and n27233_not n28094 ; n28095
g27840 and n28093_not n28095_not ; n28096
g27841 and b[62]_not n28096_not ; n28097
g27842 and b[62] n28095_not ; n28098
g27843 and n28093_not n28098 ; n28099
g27844 and b[63]_not n28099_not ; n28100
g27845 and n28097_not n28100 ; n28101
g27846 and n28086_not n28101 ; n28102
g27847 and n279 n28096_not ; n28103
g27848 and n28102_not n28103_not ; quotient[1]
g27849 and n27262_not n28079 ; n28105
g27850 and n28075_not n28105 ; n28106
g27851 and n28076_not n28079_not ; n28107
g27852 and n28106_not n28107_not ; n28108
g27853 and quotient[1] n28108_not ; n28109
g27854 and n27252_not n28103_not ; n28110
g27855 and n28102_not n28110 ; n28111
g27856 and n28109_not n28111_not ; n28112
g27857 and n27280_not n28069 ; n28113
g27858 and n28065_not n28113 ; n28114
g27859 and n28066_not n28069_not ; n28115
g27860 and n28114_not n28115_not ; n28116
g27861 and quotient[1] n28116_not ; n28117
g27862 and n27270_not n28103_not ; n28118
g27863 and n28102_not n28118 ; n28119
g27864 and n28117_not n28119_not ; n28120
g27865 and n27298_not n28059 ; n28121
g27866 and n28055_not n28121 ; n28122
g27867 and n28056_not n28059_not ; n28123
g27868 and n28122_not n28123_not ; n28124
g27869 and quotient[1] n28124_not ; n28125
g27870 and n27288_not n28103_not ; n28126
g27871 and n28102_not n28126 ; n28127
g27872 and n28125_not n28127_not ; n28128
g27873 and n27316_not n28049 ; n28129
g27874 and n28045_not n28129 ; n28130
g27875 and n28046_not n28049_not ; n28131
g27876 and n28130_not n28131_not ; n28132
g27877 and quotient[1] n28132_not ; n28133
g27878 and n27306_not n28103_not ; n28134
g27879 and n28102_not n28134 ; n28135
g27880 and n28133_not n28135_not ; n28136
g27881 and n27334_not n28039 ; n28137
g27882 and n28035_not n28137 ; n28138
g27883 and n28036_not n28039_not ; n28139
g27884 and n28138_not n28139_not ; n28140
g27885 and quotient[1] n28140_not ; n28141
g27886 and n27324_not n28103_not ; n28142
g27887 and n28102_not n28142 ; n28143
g27888 and n28141_not n28143_not ; n28144
g27889 and n27352_not n28029 ; n28145
g27890 and n28025_not n28145 ; n28146
g27891 and n28026_not n28029_not ; n28147
g27892 and n28146_not n28147_not ; n28148
g27893 and quotient[1] n28148_not ; n28149
g27894 and n27342_not n28103_not ; n28150
g27895 and n28102_not n28150 ; n28151
g27896 and n28149_not n28151_not ; n28152
g27897 and n27370_not n28019 ; n28153
g27898 and n28015_not n28153 ; n28154
g27899 and n28016_not n28019_not ; n28155
g27900 and n28154_not n28155_not ; n28156
g27901 and quotient[1] n28156_not ; n28157
g27902 and n27360_not n28103_not ; n28158
g27903 and n28102_not n28158 ; n28159
g27904 and n28157_not n28159_not ; n28160
g27905 and n27388_not n28009 ; n28161
g27906 and n28005_not n28161 ; n28162
g27907 and n28006_not n28009_not ; n28163
g27908 and n28162_not n28163_not ; n28164
g27909 and quotient[1] n28164_not ; n28165
g27910 and n27378_not n28103_not ; n28166
g27911 and n28102_not n28166 ; n28167
g27912 and n28165_not n28167_not ; n28168
g27913 and n27406_not n27999 ; n28169
g27914 and n27995_not n28169 ; n28170
g27915 and n27996_not n27999_not ; n28171
g27916 and n28170_not n28171_not ; n28172
g27917 and quotient[1] n28172_not ; n28173
g27918 and n27396_not n28103_not ; n28174
g27919 and n28102_not n28174 ; n28175
g27920 and n28173_not n28175_not ; n28176
g27921 and n27424_not n27989 ; n28177
g27922 and n27985_not n28177 ; n28178
g27923 and n27986_not n27989_not ; n28179
g27924 and n28178_not n28179_not ; n28180
g27925 and quotient[1] n28180_not ; n28181
g27926 and n27414_not n28103_not ; n28182
g27927 and n28102_not n28182 ; n28183
g27928 and n28181_not n28183_not ; n28184
g27929 and n27442_not n27979 ; n28185
g27930 and n27975_not n28185 ; n28186
g27931 and n27976_not n27979_not ; n28187
g27932 and n28186_not n28187_not ; n28188
g27933 and quotient[1] n28188_not ; n28189
g27934 and n27432_not n28103_not ; n28190
g27935 and n28102_not n28190 ; n28191
g27936 and n28189_not n28191_not ; n28192
g27937 and n27460_not n27969 ; n28193
g27938 and n27965_not n28193 ; n28194
g27939 and n27966_not n27969_not ; n28195
g27940 and n28194_not n28195_not ; n28196
g27941 and quotient[1] n28196_not ; n28197
g27942 and n27450_not n28103_not ; n28198
g27943 and n28102_not n28198 ; n28199
g27944 and n28197_not n28199_not ; n28200
g27945 and n27478_not n27959 ; n28201
g27946 and n27955_not n28201 ; n28202
g27947 and n27956_not n27959_not ; n28203
g27948 and n28202_not n28203_not ; n28204
g27949 and quotient[1] n28204_not ; n28205
g27950 and n27468_not n28103_not ; n28206
g27951 and n28102_not n28206 ; n28207
g27952 and n28205_not n28207_not ; n28208
g27953 and n27496_not n27949 ; n28209
g27954 and n27945_not n28209 ; n28210
g27955 and n27946_not n27949_not ; n28211
g27956 and n28210_not n28211_not ; n28212
g27957 and quotient[1] n28212_not ; n28213
g27958 and n27486_not n28103_not ; n28214
g27959 and n28102_not n28214 ; n28215
g27960 and n28213_not n28215_not ; n28216
g27961 and n27514_not n27939 ; n28217
g27962 and n27935_not n28217 ; n28218
g27963 and n27936_not n27939_not ; n28219
g27964 and n28218_not n28219_not ; n28220
g27965 and quotient[1] n28220_not ; n28221
g27966 and n27504_not n28103_not ; n28222
g27967 and n28102_not n28222 ; n28223
g27968 and n28221_not n28223_not ; n28224
g27969 and n27532_not n27929 ; n28225
g27970 and n27925_not n28225 ; n28226
g27971 and n27926_not n27929_not ; n28227
g27972 and n28226_not n28227_not ; n28228
g27973 and quotient[1] n28228_not ; n28229
g27974 and n27522_not n28103_not ; n28230
g27975 and n28102_not n28230 ; n28231
g27976 and n28229_not n28231_not ; n28232
g27977 and n27550_not n27919 ; n28233
g27978 and n27915_not n28233 ; n28234
g27979 and n27916_not n27919_not ; n28235
g27980 and n28234_not n28235_not ; n28236
g27981 and quotient[1] n28236_not ; n28237
g27982 and n27540_not n28103_not ; n28238
g27983 and n28102_not n28238 ; n28239
g27984 and n28237_not n28239_not ; n28240
g27985 and n27568_not n27909 ; n28241
g27986 and n27905_not n28241 ; n28242
g27987 and n27906_not n27909_not ; n28243
g27988 and n28242_not n28243_not ; n28244
g27989 and quotient[1] n28244_not ; n28245
g27990 and n27558_not n28103_not ; n28246
g27991 and n28102_not n28246 ; n28247
g27992 and n28245_not n28247_not ; n28248
g27993 and n27586_not n27899 ; n28249
g27994 and n27895_not n28249 ; n28250
g27995 and n27896_not n27899_not ; n28251
g27996 and n28250_not n28251_not ; n28252
g27997 and quotient[1] n28252_not ; n28253
g27998 and n27576_not n28103_not ; n28254
g27999 and n28102_not n28254 ; n28255
g28000 and n28253_not n28255_not ; n28256
g28001 and n27604_not n27889 ; n28257
g28002 and n27885_not n28257 ; n28258
g28003 and n27886_not n27889_not ; n28259
g28004 and n28258_not n28259_not ; n28260
g28005 and quotient[1] n28260_not ; n28261
g28006 and n27594_not n28103_not ; n28262
g28007 and n28102_not n28262 ; n28263
g28008 and n28261_not n28263_not ; n28264
g28009 and n27622_not n27879 ; n28265
g28010 and n27875_not n28265 ; n28266
g28011 and n27876_not n27879_not ; n28267
g28012 and n28266_not n28267_not ; n28268
g28013 and quotient[1] n28268_not ; n28269
g28014 and n27612_not n28103_not ; n28270
g28015 and n28102_not n28270 ; n28271
g28016 and n28269_not n28271_not ; n28272
g28017 and n27640_not n27869 ; n28273
g28018 and n27865_not n28273 ; n28274
g28019 and n27866_not n27869_not ; n28275
g28020 and n28274_not n28275_not ; n28276
g28021 and quotient[1] n28276_not ; n28277
g28022 and n27630_not n28103_not ; n28278
g28023 and n28102_not n28278 ; n28279
g28024 and n28277_not n28279_not ; n28280
g28025 and n27658_not n27859 ; n28281
g28026 and n27855_not n28281 ; n28282
g28027 and n27856_not n27859_not ; n28283
g28028 and n28282_not n28283_not ; n28284
g28029 and quotient[1] n28284_not ; n28285
g28030 and n27648_not n28103_not ; n28286
g28031 and n28102_not n28286 ; n28287
g28032 and n28285_not n28287_not ; n28288
g28033 and n27676_not n27849 ; n28289
g28034 and n27845_not n28289 ; n28290
g28035 and n27846_not n27849_not ; n28291
g28036 and n28290_not n28291_not ; n28292
g28037 and quotient[1] n28292_not ; n28293
g28038 and n27666_not n28103_not ; n28294
g28039 and n28102_not n28294 ; n28295
g28040 and n28293_not n28295_not ; n28296
g28041 and n27694_not n27839 ; n28297
g28042 and n27835_not n28297 ; n28298
g28043 and n27836_not n27839_not ; n28299
g28044 and n28298_not n28299_not ; n28300
g28045 and quotient[1] n28300_not ; n28301
g28046 and n27684_not n28103_not ; n28302
g28047 and n28102_not n28302 ; n28303
g28048 and n28301_not n28303_not ; n28304
g28049 and n27712_not n27829 ; n28305
g28050 and n27825_not n28305 ; n28306
g28051 and n27826_not n27829_not ; n28307
g28052 and n28306_not n28307_not ; n28308
g28053 and quotient[1] n28308_not ; n28309
g28054 and n27702_not n28103_not ; n28310
g28055 and n28102_not n28310 ; n28311
g28056 and n28309_not n28311_not ; n28312
g28057 and n27730_not n27819 ; n28313
g28058 and n27815_not n28313 ; n28314
g28059 and n27816_not n27819_not ; n28315
g28060 and n28314_not n28315_not ; n28316
g28061 and quotient[1] n28316_not ; n28317
g28062 and n27720_not n28103_not ; n28318
g28063 and n28102_not n28318 ; n28319
g28064 and n28317_not n28319_not ; n28320
g28065 and n27748_not n27809 ; n28321
g28066 and n27805_not n28321 ; n28322
g28067 and n27806_not n27809_not ; n28323
g28068 and n28322_not n28323_not ; n28324
g28069 and quotient[1] n28324_not ; n28325
g28070 and n27738_not n28103_not ; n28326
g28071 and n28102_not n28326 ; n28327
g28072 and n28325_not n28327_not ; n28328
g28073 and n27766_not n27799 ; n28329
g28074 and n27795_not n28329 ; n28330
g28075 and n27796_not n27799_not ; n28331
g28076 and n28330_not n28331_not ; n28332
g28077 and quotient[1] n28332_not ; n28333
g28078 and n27756_not n28103_not ; n28334
g28079 and n28102_not n28334 ; n28335
g28080 and n28333_not n28335_not ; n28336
g28081 and n27785_not n27789 ; n28337
g28082 and n27784_not n28337 ; n28338
g28083 and n27786_not n27789_not ; n28339
g28084 and n28338_not n28339_not ; n28340
g28085 and quotient[1] n28340_not ; n28341
g28086 and n27773_not n28103_not ; n28342
g28087 and n28102_not n28342 ; n28343
g28088 and n28341_not n28343_not ; n28344
g28089 and a[0]_not b[0] ; n28345
g28090 and b[0] quotient[1] ; n28346
g28091 and a[1] n28346_not ; n28347
g28092 and n27783 quotient[1] ; n28348
g28093 and n28347_not n28348_not ; n28349
g28094 and n28345_not n28349_not ; n28350
g28095 and n28345 n28348_not ; n28351
g28096 and n28347_not n28351 ; n28352
g28097 and b[1]_not n28352_not ; n28353
g28098 and n27781_not n27783 ; n28354
g28099 and n27779_not n28354 ; n28355
g28100 and n27784_not n28355_not ; n28356
g28101 and quotient[1] n28356 ; n28357
g28102 and n27778_not n28103_not ; n28358
g28103 and n28102_not n28358 ; n28359
g28104 and n28357_not n28359_not ; n28360
g28105 and n28353_not n28360 ; n28361
g28106 and n28350_not n28361 ; n28362
g28107 and b[2]_not n28362_not ; n28363
g28108 and n28350_not n28353_not ; n28364
g28109 and n28360_not n28364_not ; n28365
g28110 and n28363_not n28365_not ; n28366
g28111 and n28344_not n28366_not ; n28367
g28112 and n28344 n28365_not ; n28368
g28113 and n28363_not n28368 ; n28369
g28114 and b[3]_not n28369_not ; n28370
g28115 and n27774_not n27794 ; n28371
g28116 and n27790_not n28371 ; n28372
g28117 and n27791_not n27794_not ; n28373
g28118 and n28372_not n28373_not ; n28374
g28119 and quotient[1] n28374_not ; n28375
g28120 and n27765_not n28103_not ; n28376
g28121 and n28102_not n28376 ; n28377
g28122 and n28375_not n28377_not ; n28378
g28123 and n28370_not n28378 ; n28379
g28124 and n28367_not n28379 ; n28380
g28125 and b[4]_not n28380_not ; n28381
g28126 and n28367_not n28370_not ; n28382
g28127 and n28378_not n28382_not ; n28383
g28128 and n28381_not n28383_not ; n28384
g28129 and n28336_not n28384_not ; n28385
g28130 and n28336 n28383_not ; n28386
g28131 and n28381_not n28386 ; n28387
g28132 and b[5]_not n28387_not ; n28388
g28133 and n27757_not n27804 ; n28389
g28134 and n27800_not n28389 ; n28390
g28135 and n27801_not n27804_not ; n28391
g28136 and n28390_not n28391_not ; n28392
g28137 and quotient[1] n28392_not ; n28393
g28138 and n27747_not n28103_not ; n28394
g28139 and n28102_not n28394 ; n28395
g28140 and n28393_not n28395_not ; n28396
g28141 and n28388_not n28396 ; n28397
g28142 and n28385_not n28397 ; n28398
g28143 and b[6]_not n28398_not ; n28399
g28144 and n28385_not n28388_not ; n28400
g28145 and n28396_not n28400_not ; n28401
g28146 and n28399_not n28401_not ; n28402
g28147 and n28328_not n28402_not ; n28403
g28148 and n28328 n28401_not ; n28404
g28149 and n28399_not n28404 ; n28405
g28150 and b[7]_not n28405_not ; n28406
g28151 and n27739_not n27814 ; n28407
g28152 and n27810_not n28407 ; n28408
g28153 and n27811_not n27814_not ; n28409
g28154 and n28408_not n28409_not ; n28410
g28155 and quotient[1] n28410_not ; n28411
g28156 and n27729_not n28103_not ; n28412
g28157 and n28102_not n28412 ; n28413
g28158 and n28411_not n28413_not ; n28414
g28159 and n28406_not n28414 ; n28415
g28160 and n28403_not n28415 ; n28416
g28161 and b[8]_not n28416_not ; n28417
g28162 and n28403_not n28406_not ; n28418
g28163 and n28414_not n28418_not ; n28419
g28164 and n28417_not n28419_not ; n28420
g28165 and n28320_not n28420_not ; n28421
g28166 and n28320 n28419_not ; n28422
g28167 and n28417_not n28422 ; n28423
g28168 and b[9]_not n28423_not ; n28424
g28169 and n27721_not n27824 ; n28425
g28170 and n27820_not n28425 ; n28426
g28171 and n27821_not n27824_not ; n28427
g28172 and n28426_not n28427_not ; n28428
g28173 and quotient[1] n28428_not ; n28429
g28174 and n27711_not n28103_not ; n28430
g28175 and n28102_not n28430 ; n28431
g28176 and n28429_not n28431_not ; n28432
g28177 and n28424_not n28432 ; n28433
g28178 and n28421_not n28433 ; n28434
g28179 and b[10]_not n28434_not ; n28435
g28180 and n28421_not n28424_not ; n28436
g28181 and n28432_not n28436_not ; n28437
g28182 and n28435_not n28437_not ; n28438
g28183 and n28312_not n28438_not ; n28439
g28184 and n28312 n28437_not ; n28440
g28185 and n28435_not n28440 ; n28441
g28186 and b[11]_not n28441_not ; n28442
g28187 and n27703_not n27834 ; n28443
g28188 and n27830_not n28443 ; n28444
g28189 and n27831_not n27834_not ; n28445
g28190 and n28444_not n28445_not ; n28446
g28191 and quotient[1] n28446_not ; n28447
g28192 and n27693_not n28103_not ; n28448
g28193 and n28102_not n28448 ; n28449
g28194 and n28447_not n28449_not ; n28450
g28195 and n28442_not n28450 ; n28451
g28196 and n28439_not n28451 ; n28452
g28197 and b[12]_not n28452_not ; n28453
g28198 and n28439_not n28442_not ; n28454
g28199 and n28450_not n28454_not ; n28455
g28200 and n28453_not n28455_not ; n28456
g28201 and n28304_not n28456_not ; n28457
g28202 and n28304 n28455_not ; n28458
g28203 and n28453_not n28458 ; n28459
g28204 and b[13]_not n28459_not ; n28460
g28205 and n27685_not n27844 ; n28461
g28206 and n27840_not n28461 ; n28462
g28207 and n27841_not n27844_not ; n28463
g28208 and n28462_not n28463_not ; n28464
g28209 and quotient[1] n28464_not ; n28465
g28210 and n27675_not n28103_not ; n28466
g28211 and n28102_not n28466 ; n28467
g28212 and n28465_not n28467_not ; n28468
g28213 and n28460_not n28468 ; n28469
g28214 and n28457_not n28469 ; n28470
g28215 and b[14]_not n28470_not ; n28471
g28216 and n28457_not n28460_not ; n28472
g28217 and n28468_not n28472_not ; n28473
g28218 and n28471_not n28473_not ; n28474
g28219 and n28296_not n28474_not ; n28475
g28220 and n28296 n28473_not ; n28476
g28221 and n28471_not n28476 ; n28477
g28222 and b[15]_not n28477_not ; n28478
g28223 and n27667_not n27854 ; n28479
g28224 and n27850_not n28479 ; n28480
g28225 and n27851_not n27854_not ; n28481
g28226 and n28480_not n28481_not ; n28482
g28227 and quotient[1] n28482_not ; n28483
g28228 and n27657_not n28103_not ; n28484
g28229 and n28102_not n28484 ; n28485
g28230 and n28483_not n28485_not ; n28486
g28231 and n28478_not n28486 ; n28487
g28232 and n28475_not n28487 ; n28488
g28233 and b[16]_not n28488_not ; n28489
g28234 and n28475_not n28478_not ; n28490
g28235 and n28486_not n28490_not ; n28491
g28236 and n28489_not n28491_not ; n28492
g28237 and n28288_not n28492_not ; n28493
g28238 and n28288 n28491_not ; n28494
g28239 and n28489_not n28494 ; n28495
g28240 and b[17]_not n28495_not ; n28496
g28241 and n27649_not n27864 ; n28497
g28242 and n27860_not n28497 ; n28498
g28243 and n27861_not n27864_not ; n28499
g28244 and n28498_not n28499_not ; n28500
g28245 and quotient[1] n28500_not ; n28501
g28246 and n27639_not n28103_not ; n28502
g28247 and n28102_not n28502 ; n28503
g28248 and n28501_not n28503_not ; n28504
g28249 and n28496_not n28504 ; n28505
g28250 and n28493_not n28505 ; n28506
g28251 and b[18]_not n28506_not ; n28507
g28252 and n28493_not n28496_not ; n28508
g28253 and n28504_not n28508_not ; n28509
g28254 and n28507_not n28509_not ; n28510
g28255 and n28280_not n28510_not ; n28511
g28256 and n28280 n28509_not ; n28512
g28257 and n28507_not n28512 ; n28513
g28258 and b[19]_not n28513_not ; n28514
g28259 and n27631_not n27874 ; n28515
g28260 and n27870_not n28515 ; n28516
g28261 and n27871_not n27874_not ; n28517
g28262 and n28516_not n28517_not ; n28518
g28263 and quotient[1] n28518_not ; n28519
g28264 and n27621_not n28103_not ; n28520
g28265 and n28102_not n28520 ; n28521
g28266 and n28519_not n28521_not ; n28522
g28267 and n28514_not n28522 ; n28523
g28268 and n28511_not n28523 ; n28524
g28269 and b[20]_not n28524_not ; n28525
g28270 and n28511_not n28514_not ; n28526
g28271 and n28522_not n28526_not ; n28527
g28272 and n28525_not n28527_not ; n28528
g28273 and n28272_not n28528_not ; n28529
g28274 and n28272 n28527_not ; n28530
g28275 and n28525_not n28530 ; n28531
g28276 and b[21]_not n28531_not ; n28532
g28277 and n27613_not n27884 ; n28533
g28278 and n27880_not n28533 ; n28534
g28279 and n27881_not n27884_not ; n28535
g28280 and n28534_not n28535_not ; n28536
g28281 and quotient[1] n28536_not ; n28537
g28282 and n27603_not n28103_not ; n28538
g28283 and n28102_not n28538 ; n28539
g28284 and n28537_not n28539_not ; n28540
g28285 and n28532_not n28540 ; n28541
g28286 and n28529_not n28541 ; n28542
g28287 and b[22]_not n28542_not ; n28543
g28288 and n28529_not n28532_not ; n28544
g28289 and n28540_not n28544_not ; n28545
g28290 and n28543_not n28545_not ; n28546
g28291 and n28264_not n28546_not ; n28547
g28292 and n28264 n28545_not ; n28548
g28293 and n28543_not n28548 ; n28549
g28294 and b[23]_not n28549_not ; n28550
g28295 and n27595_not n27894 ; n28551
g28296 and n27890_not n28551 ; n28552
g28297 and n27891_not n27894_not ; n28553
g28298 and n28552_not n28553_not ; n28554
g28299 and quotient[1] n28554_not ; n28555
g28300 and n27585_not n28103_not ; n28556
g28301 and n28102_not n28556 ; n28557
g28302 and n28555_not n28557_not ; n28558
g28303 and n28550_not n28558 ; n28559
g28304 and n28547_not n28559 ; n28560
g28305 and b[24]_not n28560_not ; n28561
g28306 and n28547_not n28550_not ; n28562
g28307 and n28558_not n28562_not ; n28563
g28308 and n28561_not n28563_not ; n28564
g28309 and n28256_not n28564_not ; n28565
g28310 and n28256 n28563_not ; n28566
g28311 and n28561_not n28566 ; n28567
g28312 and b[25]_not n28567_not ; n28568
g28313 and n27577_not n27904 ; n28569
g28314 and n27900_not n28569 ; n28570
g28315 and n27901_not n27904_not ; n28571
g28316 and n28570_not n28571_not ; n28572
g28317 and quotient[1] n28572_not ; n28573
g28318 and n27567_not n28103_not ; n28574
g28319 and n28102_not n28574 ; n28575
g28320 and n28573_not n28575_not ; n28576
g28321 and n28568_not n28576 ; n28577
g28322 and n28565_not n28577 ; n28578
g28323 and b[26]_not n28578_not ; n28579
g28324 and n28565_not n28568_not ; n28580
g28325 and n28576_not n28580_not ; n28581
g28326 and n28579_not n28581_not ; n28582
g28327 and n28248_not n28582_not ; n28583
g28328 and n28248 n28581_not ; n28584
g28329 and n28579_not n28584 ; n28585
g28330 and b[27]_not n28585_not ; n28586
g28331 and n27559_not n27914 ; n28587
g28332 and n27910_not n28587 ; n28588
g28333 and n27911_not n27914_not ; n28589
g28334 and n28588_not n28589_not ; n28590
g28335 and quotient[1] n28590_not ; n28591
g28336 and n27549_not n28103_not ; n28592
g28337 and n28102_not n28592 ; n28593
g28338 and n28591_not n28593_not ; n28594
g28339 and n28586_not n28594 ; n28595
g28340 and n28583_not n28595 ; n28596
g28341 and b[28]_not n28596_not ; n28597
g28342 and n28583_not n28586_not ; n28598
g28343 and n28594_not n28598_not ; n28599
g28344 and n28597_not n28599_not ; n28600
g28345 and n28240_not n28600_not ; n28601
g28346 and n28240 n28599_not ; n28602
g28347 and n28597_not n28602 ; n28603
g28348 and b[29]_not n28603_not ; n28604
g28349 and n27541_not n27924 ; n28605
g28350 and n27920_not n28605 ; n28606
g28351 and n27921_not n27924_not ; n28607
g28352 and n28606_not n28607_not ; n28608
g28353 and quotient[1] n28608_not ; n28609
g28354 and n27531_not n28103_not ; n28610
g28355 and n28102_not n28610 ; n28611
g28356 and n28609_not n28611_not ; n28612
g28357 and n28604_not n28612 ; n28613
g28358 and n28601_not n28613 ; n28614
g28359 and b[30]_not n28614_not ; n28615
g28360 and n28601_not n28604_not ; n28616
g28361 and n28612_not n28616_not ; n28617
g28362 and n28615_not n28617_not ; n28618
g28363 and n28232_not n28618_not ; n28619
g28364 and n28232 n28617_not ; n28620
g28365 and n28615_not n28620 ; n28621
g28366 and b[31]_not n28621_not ; n28622
g28367 and n27523_not n27934 ; n28623
g28368 and n27930_not n28623 ; n28624
g28369 and n27931_not n27934_not ; n28625
g28370 and n28624_not n28625_not ; n28626
g28371 and quotient[1] n28626_not ; n28627
g28372 and n27513_not n28103_not ; n28628
g28373 and n28102_not n28628 ; n28629
g28374 and n28627_not n28629_not ; n28630
g28375 and n28622_not n28630 ; n28631
g28376 and n28619_not n28631 ; n28632
g28377 and b[32]_not n28632_not ; n28633
g28378 and n28619_not n28622_not ; n28634
g28379 and n28630_not n28634_not ; n28635
g28380 and n28633_not n28635_not ; n28636
g28381 and n28224_not n28636_not ; n28637
g28382 and n28224 n28635_not ; n28638
g28383 and n28633_not n28638 ; n28639
g28384 and b[33]_not n28639_not ; n28640
g28385 and n27505_not n27944 ; n28641
g28386 and n27940_not n28641 ; n28642
g28387 and n27941_not n27944_not ; n28643
g28388 and n28642_not n28643_not ; n28644
g28389 and quotient[1] n28644_not ; n28645
g28390 and n27495_not n28103_not ; n28646
g28391 and n28102_not n28646 ; n28647
g28392 and n28645_not n28647_not ; n28648
g28393 and n28640_not n28648 ; n28649
g28394 and n28637_not n28649 ; n28650
g28395 and b[34]_not n28650_not ; n28651
g28396 and n28637_not n28640_not ; n28652
g28397 and n28648_not n28652_not ; n28653
g28398 and n28651_not n28653_not ; n28654
g28399 and n28216_not n28654_not ; n28655
g28400 and n28216 n28653_not ; n28656
g28401 and n28651_not n28656 ; n28657
g28402 and b[35]_not n28657_not ; n28658
g28403 and n27487_not n27954 ; n28659
g28404 and n27950_not n28659 ; n28660
g28405 and n27951_not n27954_not ; n28661
g28406 and n28660_not n28661_not ; n28662
g28407 and quotient[1] n28662_not ; n28663
g28408 and n27477_not n28103_not ; n28664
g28409 and n28102_not n28664 ; n28665
g28410 and n28663_not n28665_not ; n28666
g28411 and n28658_not n28666 ; n28667
g28412 and n28655_not n28667 ; n28668
g28413 and b[36]_not n28668_not ; n28669
g28414 and n28655_not n28658_not ; n28670
g28415 and n28666_not n28670_not ; n28671
g28416 and n28669_not n28671_not ; n28672
g28417 and n28208_not n28672_not ; n28673
g28418 and n28208 n28671_not ; n28674
g28419 and n28669_not n28674 ; n28675
g28420 and b[37]_not n28675_not ; n28676
g28421 and n27469_not n27964 ; n28677
g28422 and n27960_not n28677 ; n28678
g28423 and n27961_not n27964_not ; n28679
g28424 and n28678_not n28679_not ; n28680
g28425 and quotient[1] n28680_not ; n28681
g28426 and n27459_not n28103_not ; n28682
g28427 and n28102_not n28682 ; n28683
g28428 and n28681_not n28683_not ; n28684
g28429 and n28676_not n28684 ; n28685
g28430 and n28673_not n28685 ; n28686
g28431 and b[38]_not n28686_not ; n28687
g28432 and n28673_not n28676_not ; n28688
g28433 and n28684_not n28688_not ; n28689
g28434 and n28687_not n28689_not ; n28690
g28435 and n28200_not n28690_not ; n28691
g28436 and n28200 n28689_not ; n28692
g28437 and n28687_not n28692 ; n28693
g28438 and b[39]_not n28693_not ; n28694
g28439 and n27451_not n27974 ; n28695
g28440 and n27970_not n28695 ; n28696
g28441 and n27971_not n27974_not ; n28697
g28442 and n28696_not n28697_not ; n28698
g28443 and quotient[1] n28698_not ; n28699
g28444 and n27441_not n28103_not ; n28700
g28445 and n28102_not n28700 ; n28701
g28446 and n28699_not n28701_not ; n28702
g28447 and n28694_not n28702 ; n28703
g28448 and n28691_not n28703 ; n28704
g28449 and b[40]_not n28704_not ; n28705
g28450 and n28691_not n28694_not ; n28706
g28451 and n28702_not n28706_not ; n28707
g28452 and n28705_not n28707_not ; n28708
g28453 and n28192_not n28708_not ; n28709
g28454 and n28192 n28707_not ; n28710
g28455 and n28705_not n28710 ; n28711
g28456 and b[41]_not n28711_not ; n28712
g28457 and n27433_not n27984 ; n28713
g28458 and n27980_not n28713 ; n28714
g28459 and n27981_not n27984_not ; n28715
g28460 and n28714_not n28715_not ; n28716
g28461 and quotient[1] n28716_not ; n28717
g28462 and n27423_not n28103_not ; n28718
g28463 and n28102_not n28718 ; n28719
g28464 and n28717_not n28719_not ; n28720
g28465 and n28712_not n28720 ; n28721
g28466 and n28709_not n28721 ; n28722
g28467 and b[42]_not n28722_not ; n28723
g28468 and n28709_not n28712_not ; n28724
g28469 and n28720_not n28724_not ; n28725
g28470 and n28723_not n28725_not ; n28726
g28471 and n28184_not n28726_not ; n28727
g28472 and n28184 n28725_not ; n28728
g28473 and n28723_not n28728 ; n28729
g28474 and b[43]_not n28729_not ; n28730
g28475 and n27415_not n27994 ; n28731
g28476 and n27990_not n28731 ; n28732
g28477 and n27991_not n27994_not ; n28733
g28478 and n28732_not n28733_not ; n28734
g28479 and quotient[1] n28734_not ; n28735
g28480 and n27405_not n28103_not ; n28736
g28481 and n28102_not n28736 ; n28737
g28482 and n28735_not n28737_not ; n28738
g28483 and n28730_not n28738 ; n28739
g28484 and n28727_not n28739 ; n28740
g28485 and b[44]_not n28740_not ; n28741
g28486 and n28727_not n28730_not ; n28742
g28487 and n28738_not n28742_not ; n28743
g28488 and n28741_not n28743_not ; n28744
g28489 and n28176_not n28744_not ; n28745
g28490 and n28176 n28743_not ; n28746
g28491 and n28741_not n28746 ; n28747
g28492 and b[45]_not n28747_not ; n28748
g28493 and n27397_not n28004 ; n28749
g28494 and n28000_not n28749 ; n28750
g28495 and n28001_not n28004_not ; n28751
g28496 and n28750_not n28751_not ; n28752
g28497 and quotient[1] n28752_not ; n28753
g28498 and n27387_not n28103_not ; n28754
g28499 and n28102_not n28754 ; n28755
g28500 and n28753_not n28755_not ; n28756
g28501 and n28748_not n28756 ; n28757
g28502 and n28745_not n28757 ; n28758
g28503 and b[46]_not n28758_not ; n28759
g28504 and n28745_not n28748_not ; n28760
g28505 and n28756_not n28760_not ; n28761
g28506 and n28759_not n28761_not ; n28762
g28507 and n28168_not n28762_not ; n28763
g28508 and n28168 n28761_not ; n28764
g28509 and n28759_not n28764 ; n28765
g28510 and b[47]_not n28765_not ; n28766
g28511 and n27379_not n28014 ; n28767
g28512 and n28010_not n28767 ; n28768
g28513 and n28011_not n28014_not ; n28769
g28514 and n28768_not n28769_not ; n28770
g28515 and quotient[1] n28770_not ; n28771
g28516 and n27369_not n28103_not ; n28772
g28517 and n28102_not n28772 ; n28773
g28518 and n28771_not n28773_not ; n28774
g28519 and n28766_not n28774 ; n28775
g28520 and n28763_not n28775 ; n28776
g28521 and b[48]_not n28776_not ; n28777
g28522 and n28763_not n28766_not ; n28778
g28523 and n28774_not n28778_not ; n28779
g28524 and n28777_not n28779_not ; n28780
g28525 and n28160_not n28780_not ; n28781
g28526 and n28160 n28779_not ; n28782
g28527 and n28777_not n28782 ; n28783
g28528 and b[49]_not n28783_not ; n28784
g28529 and n27361_not n28024 ; n28785
g28530 and n28020_not n28785 ; n28786
g28531 and n28021_not n28024_not ; n28787
g28532 and n28786_not n28787_not ; n28788
g28533 and quotient[1] n28788_not ; n28789
g28534 and n27351_not n28103_not ; n28790
g28535 and n28102_not n28790 ; n28791
g28536 and n28789_not n28791_not ; n28792
g28537 and n28784_not n28792 ; n28793
g28538 and n28781_not n28793 ; n28794
g28539 and b[50]_not n28794_not ; n28795
g28540 and n28781_not n28784_not ; n28796
g28541 and n28792_not n28796_not ; n28797
g28542 and n28795_not n28797_not ; n28798
g28543 and n28152_not n28798_not ; n28799
g28544 and n28152 n28797_not ; n28800
g28545 and n28795_not n28800 ; n28801
g28546 and b[51]_not n28801_not ; n28802
g28547 and n27343_not n28034 ; n28803
g28548 and n28030_not n28803 ; n28804
g28549 and n28031_not n28034_not ; n28805
g28550 and n28804_not n28805_not ; n28806
g28551 and quotient[1] n28806_not ; n28807
g28552 and n27333_not n28103_not ; n28808
g28553 and n28102_not n28808 ; n28809
g28554 and n28807_not n28809_not ; n28810
g28555 and n28802_not n28810 ; n28811
g28556 and n28799_not n28811 ; n28812
g28557 and b[52]_not n28812_not ; n28813
g28558 and n28799_not n28802_not ; n28814
g28559 and n28810_not n28814_not ; n28815
g28560 and n28813_not n28815_not ; n28816
g28561 and n28144_not n28816_not ; n28817
g28562 and n28144 n28815_not ; n28818
g28563 and n28813_not n28818 ; n28819
g28564 and b[53]_not n28819_not ; n28820
g28565 and n27325_not n28044 ; n28821
g28566 and n28040_not n28821 ; n28822
g28567 and n28041_not n28044_not ; n28823
g28568 and n28822_not n28823_not ; n28824
g28569 and quotient[1] n28824_not ; n28825
g28570 and n27315_not n28103_not ; n28826
g28571 and n28102_not n28826 ; n28827
g28572 and n28825_not n28827_not ; n28828
g28573 and n28820_not n28828 ; n28829
g28574 and n28817_not n28829 ; n28830
g28575 and b[54]_not n28830_not ; n28831
g28576 and n28817_not n28820_not ; n28832
g28577 and n28828_not n28832_not ; n28833
g28578 and n28831_not n28833_not ; n28834
g28579 and n28136_not n28834_not ; n28835
g28580 and n28136 n28833_not ; n28836
g28581 and n28831_not n28836 ; n28837
g28582 and b[55]_not n28837_not ; n28838
g28583 and n27307_not n28054 ; n28839
g28584 and n28050_not n28839 ; n28840
g28585 and n28051_not n28054_not ; n28841
g28586 and n28840_not n28841_not ; n28842
g28587 and quotient[1] n28842_not ; n28843
g28588 and n27297_not n28103_not ; n28844
g28589 and n28102_not n28844 ; n28845
g28590 and n28843_not n28845_not ; n28846
g28591 and n28838_not n28846 ; n28847
g28592 and n28835_not n28847 ; n28848
g28593 and b[56]_not n28848_not ; n28849
g28594 and n28835_not n28838_not ; n28850
g28595 and n28846_not n28850_not ; n28851
g28596 and n28849_not n28851_not ; n28852
g28597 and n28128_not n28852_not ; n28853
g28598 and n28128 n28851_not ; n28854
g28599 and n28849_not n28854 ; n28855
g28600 and b[57]_not n28855_not ; n28856
g28601 and n27289_not n28064 ; n28857
g28602 and n28060_not n28857 ; n28858
g28603 and n28061_not n28064_not ; n28859
g28604 and n28858_not n28859_not ; n28860
g28605 and quotient[1] n28860_not ; n28861
g28606 and n27279_not n28103_not ; n28862
g28607 and n28102_not n28862 ; n28863
g28608 and n28861_not n28863_not ; n28864
g28609 and n28856_not n28864 ; n28865
g28610 and n28853_not n28865 ; n28866
g28611 and b[58]_not n28866_not ; n28867
g28612 and n28853_not n28856_not ; n28868
g28613 and n28864_not n28868_not ; n28869
g28614 and n28867_not n28869_not ; n28870
g28615 and n28120_not n28870_not ; n28871
g28616 and n28120 n28869_not ; n28872
g28617 and n28867_not n28872 ; n28873
g28618 and b[59]_not n28873_not ; n28874
g28619 and n27271_not n28074 ; n28875
g28620 and n28070_not n28875 ; n28876
g28621 and n28071_not n28074_not ; n28877
g28622 and n28876_not n28877_not ; n28878
g28623 and quotient[1] n28878_not ; n28879
g28624 and n27261_not n28103_not ; n28880
g28625 and n28102_not n28880 ; n28881
g28626 and n28879_not n28881_not ; n28882
g28627 and n28874_not n28882 ; n28883
g28628 and n28871_not n28883 ; n28884
g28629 and b[60]_not n28884_not ; n28885
g28630 and n28871_not n28874_not ; n28886
g28631 and n28882_not n28886_not ; n28887
g28632 and n28885_not n28887_not ; n28888
g28633 and n28112_not n28888_not ; n28889
g28634 and n28112 n28887_not ; n28890
g28635 and n28885_not n28890 ; n28891
g28636 and b[61]_not n28891_not ; n28892
g28637 and n27253_not n28084 ; n28893
g28638 and n28080_not n28893 ; n28894
g28639 and n28081_not n28084_not ; n28895
g28640 and n28894_not n28895_not ; n28896
g28641 and quotient[1] n28896_not ; n28897
g28642 and n27243_not n28103_not ; n28898
g28643 and n28102_not n28898 ; n28899
g28644 and n28897_not n28899_not ; n28900
g28645 and n28892_not n28900 ; n28901
g28646 and n28889_not n28901 ; n28902
g28647 and b[62]_not n28902_not ; n28903
g28648 and n28889_not n28892_not ; n28904
g28649 and n28900_not n28904_not ; n28905
g28650 and n27244_not n28099_not ; n28906
g28651 and n28097_not n28906 ; n28907
g28652 and n28085_not n28907 ; n28908
g28653 and n28097_not n28099_not ; n28909
g28654 and n28086_not n28909_not ; n28910
g28655 and n28908_not n28910_not ; n28911
g28656 and quotient[1] n28911_not ; n28912
g28657 and n28096_not n28103_not ; n28913
g28658 and n28102_not n28913 ; n28914
g28659 and n28912_not n28914_not ; n28915
g28660 and n28905_not n28915 ; n28916
g28661 and n28903_not n28916 ; n28917
g28662 and b[63]_not n28917_not ; n28918
g28663 and n28903_not n28905_not ; n28919
g28664 and n28915_not n28919_not ; n28920
g28665 and n28918_not n28920_not ; quotient[0]
g28666 and n583_not n600 ; quotient[59]
g28667 and n334 n344 ; n28923
g28668 and n432 n28923 ; n28924
g28669 and n327_not n28924 ; quotient[62]
g28670 and b[1]_not b[2]_not ; n28926
g28671 and n383 n28926 ; n28927
g28672 and n257_not n28927 ; n28928
g28673 and n592 n28928 ; n28929
g28674 and n643 n28929 ; quotient[63]
g28675 and n260 n267 ; n28931
g28676 and n333 n28931 ; n28932
g28677 and n344 n28932 ; n28933
g28678 and n432 n28933 ; n28934
g28679 and n324 n28934_not ; n28935
g28680 and n326_not n28935_not ; n28936
g28681 and a[63] n28934_not ; n28937
g28682 and n347 n28937_not ; n28938
g28683 and n28936_not n28938 ; n28939
g28684 and n358 n28936_not ; n28940
g28685 and n28937 n28940_not ; n28941
g28686 and n28939_not n28941_not ; n28942
g28687 and n425 n28936_not ; n28943
g28688 and a[62] n28943_not ; n28944
g28689 and n433 n28936_not ; n28945
g28690 and n28944_not n28945_not ; n28946
g28691 and n363_not n28946_not ; n28947
g28692 and n437_not n28947_not ; n28948
g28693 and b[2] n28939_not ; n28949
g28694 and n28941_not n28949 ; n28950
g28695 and b[2]_not n28942_not ; n28951
g28696 and n28950_not n28951_not ; n28952
g28697 and n28948 n28952_not ; n28953
g28698 and b[2]_not n28953_not ; n28954
g28699 and n28948_not n28950_not ; n28955
g28700 and n28951_not n28955_not ; n28956
g28701 and n450 n28956_not ; n28957
g28702 and n28954_not n28957 ; n28958
g28703 and n28942_not n28958_not ; n28959
g28704 and n450 n28955_not ; n28960
g28705 and n28953_not n28960 ; n28961
g28706 and n28956_not n28961 ; n28962
g28707 and b[3] n28962_not ; n28963
g28708 and n28959_not n28963 ; n28964
g28709 and n467 n28956_not ; n28965
g28710 and n28946_not n28965_not ; n28966
g28711 and n476 n28945_not ; n28967
g28712 and n28944_not n28967 ; n28968
g28713 and n28956_not n28968 ; n28969
g28714 and n28966_not n28969_not ; n28970
g28715 and b[2]_not n28970_not ; n28971
g28716 and b[2] n28969_not ; n28972
g28717 and n28966_not n28972 ; n28973
g28718 and n488 n28956_not ; n28974
g28719 and a[61] n28974_not ; n28975
g28720 and n495 n28956_not ; n28976
g28721 and n28975_not n28976_not ; n28977
g28722 and n499_not n28977_not ; n28978
g28723 and n501_not n28978_not ; n28979
g28724 and n28973_not n28979_not ; n28980
g28725 and n28971_not n28980_not ; n28981
g28726 and n28964_not n28981_not ; n28982
g28727 and n28959_not n28962_not ; n28983
g28728 and b[3]_not n28983_not ; n28984
g28729 and n28982_not n28984_not ; n28985
g28730 and n28964_not n28984_not ; n28986
g28731 and n28981_not n28986 ; n28987
g28732 and n28981 n28986_not ; n28988
g28733 and n513 n28988_not ; n28989
g28734 and n28987_not n28989 ; n28990
g28735 and n28985_not n28990 ; n28991
g28736 and n513 n28985_not ; n28992
g28737 and n28983_not n28992_not ; n28993
g28738 and b[4] n28993_not ; n28994
g28739 and n28991_not n28994 ; n28995
g28740 and n28971_not n28973_not ; n28996
g28741 and n28979 n28996_not ; n28997
g28742 and n513 n28980_not ; n28998
g28743 and n28997_not n28998 ; n28999
g28744 and n28985_not n28999 ; n29000
g28745 and b[2]_not n28997_not ; n29001
g28746 and n513 n29001_not ; n29002
g28747 and n28985_not n29002 ; n29003
g28748 and n28970_not n29003_not ; n29004
g28749 and n29000_not n29004_not ; n29005
g28750 and b[3]_not n29005_not ; n29006
g28751 and b[3] n29000_not ; n29007
g28752 and n29004_not n29007 ; n29008
g28753 and n543 n28985_not ; n29009
g28754 and n28977_not n29009_not ; n29010
g28755 and n550 n28976_not ; n29011
g28756 and n28975_not n29011 ; n29012
g28757 and n28985_not n29012 ; n29013
g28758 and n29010_not n29013_not ; n29014
g28759 and b[2]_not n29014_not ; n29015
g28760 and b[2] n29013_not ; n29016
g28761 and n29010_not n29016 ; n29017
g28762 and n564 n28985_not ; n29018
g28763 and a[60] n29018_not ; n29019
g28764 and n570 n28985_not ; n29020
g28765 and n29019_not n29020_not ; n29021
g28766 and n559_not n29021_not ; n29022
g28767 and n574_not n29022_not ; n29023
g28768 and n29017_not n29023_not ; n29024
g28769 and n29015_not n29024_not ; n29025
g28770 and n29008_not n29025_not ; n29026
g28771 and n29006_not n29026_not ; n29027
g28772 and n28995_not n29027_not ; n29028
g28773 and n28991_not n28993_not ; n29029
g28774 and b[4]_not n29029_not ; n29030
g28775 and n29028_not n29030_not ; n29031
g28776 and n29006_not n29008_not ; n29032
g28777 and n29015_not n29032_not ; n29033
g28778 and n29024_not n29033 ; n29034
g28779 and n600 n29034_not ; n29035
g28780 and n29026_not n29035 ; n29036
g28781 and n29031_not n29036 ; n29037
g28782 and b[3]_not n29034_not ; n29038
g28783 and n600 n29038_not ; n29039
g28784 and n29031_not n29039 ; n29040
g28785 and n29005_not n29040_not ; n29041
g28786 and n29037_not n29041_not ; n29042
g28787 and b[4] n29042_not ; n29043
g28788 and b[4]_not n29037_not ; n29044
g28789 and n29041_not n29044 ; n29045
g28790 and n29043_not n29045_not ; n29046
g28791 and n29015_not n29017_not ; n29047
g28792 and n29023 n29047_not ; n29048
g28793 and n600 n29024_not ; n29049
g28794 and n29048_not n29049 ; n29050
g28795 and n29031_not n29050 ; n29051
g28796 and b[2]_not n29048_not ; n29052
g28797 and n600 n29052_not ; n29053
g28798 and n29031_not n29053 ; n29054
g28799 and n29014_not n29054_not ; n29055
g28800 and n29051_not n29055_not ; n29056
g28801 and b[3] n29056_not ; n29057
g28802 and b[3]_not n29051_not ; n29058
g28803 and n29055_not n29058 ; n29059
g28804 and n29057_not n29059_not ; n29060
g28805 and n635 n29031_not ; n29061
g28806 and n29021_not n29061_not ; n29062
g28807 and n644 n29020_not ; n29063
g28808 and n29019_not n29063 ; n29064
g28809 and n29031_not n29064 ; n29065
g28810 and n29062_not n29065_not ; n29066
g28811 and b[2]_not n29066_not ; n29067
g28812 and n655 n29031_not ; n29068
g28813 and a[59] n29068_not ; n29069
g28814 and n661 n29031_not ; n29070
g28815 and n29069_not n29070_not ; n29071
g28816 and b[1] n29071_not ; n29072
g28817 and b[1]_not n29070_not ; n29073
g28818 and n29069_not n29073 ; n29074
g28819 and n29072_not n29074_not ; n29075
g28820 and n668_not n29075_not ; n29076
g28821 and b[1]_not n29071_not ; n29077
g28822 and n29076_not n29077_not ; n29078
g28823 and b[2] n29065_not ; n29079
g28824 and n29062_not n29079 ; n29080
g28825 and n29067_not n29080_not ; n29081
g28826 and n29078_not n29081 ; n29082
g28827 and n29067_not n29082_not ; n29083
g28828 and n29060_not n29083_not ; n29084
g28829 and b[3]_not n29056_not ; n29085
g28830 and n29084_not n29085_not ; n29086
g28831 and n29046_not n29086_not ; n29087
g28832 and b[4]_not n29042_not ; n29088
g28833 and n29087_not n29088_not ; n29089
g28834 and n28995_not n29030_not ; n29090
g28835 and n29006_not n29090_not ; n29091
g28836 and n29026_not n29091 ; n29092
g28837 and n600 n29092_not ; n29093
g28838 and n29028_not n29093 ; n29094
g28839 and n29031_not n29094 ; n29095
g28840 and b[4]_not n29092_not ; n29096
g28841 and n600 n29096_not ; n29097
g28842 and n29031_not n29097 ; n29098
g28843 and n29029_not n29098_not ; n29099
g28844 and n29095_not n29099_not ; n29100
g28845 and b[5] n29100_not ; n29101
g28846 and b[5]_not n29095_not ; n29102
g28847 and n29099_not n29102 ; n29103
g28848 and n29101_not n29103_not ; n29104
g28849 and n701 n29104_not ; n29105
g28850 and n29089_not n29105 ; n29106
g28851 and n600 n29100_not ; n29107
g28852 and n29106_not n29107_not ; n29108
g28853 and n29046 n29085_not ; n29109
g28854 and n29084_not n29109 ; n29110
g28855 and n29087_not n29110_not ; n29111
g28856 and n29108_not n29111 ; n29112
g28857 and n29042_not n29107_not ; n29113
g28858 and n29106_not n29113 ; n29114
g28859 and n29112_not n29114_not ; n29115
g28860 and n29089_not n29104_not ; n29116
g28861 and n29088_not n29104 ; n29117
g28862 and n29087_not n29117 ; n29118
g28863 and n29116_not n29118_not ; n29119
g28864 and n29108_not n29119 ; n29120
g28865 and n29100_not n29107_not ; n29121
g28866 and n29106_not n29121 ; n29122
g28867 and n29120_not n29122_not ; n29123
g28868 and b[6]_not n29123_not ; n29124
g28869 and b[5]_not n29115_not ; n29125
g28870 and n29060 n29067_not ; n29126
g28871 and n29082_not n29126 ; n29127
g28872 and n29084_not n29127_not ; n29128
g28873 and n29108_not n29128 ; n29129
g28874 and n29056_not n29107_not ; n29130
g28875 and n29106_not n29130 ; n29131
g28876 and n29129_not n29131_not ; n29132
g28877 and b[4]_not n29132_not ; n29133
g28878 and n29077_not n29081 ; n29134
g28879 and n29076_not n29134 ; n29135
g28880 and n29078_not n29081_not ; n29136
g28881 and n29135_not n29136_not ; n29137
g28882 and n29108_not n29137_not ; n29138
g28883 and n29066_not n29107_not ; n29139
g28884 and n29106_not n29139 ; n29140
g28885 and n29138_not n29140_not ; n29141
g28886 and b[3]_not n29141_not ; n29142
g28887 and n668 n29074_not ; n29143
g28888 and n29072_not n29143 ; n29144
g28889 and n29076_not n29144_not ; n29145
g28890 and n29108_not n29145 ; n29146
g28891 and n29071_not n29107_not ; n29147
g28892 and n29106_not n29147 ; n29148
g28893 and n29146_not n29148_not ; n29149
g28894 and b[2]_not n29149_not ; n29150
g28895 and b[0] n29108_not ; n29151
g28896 and a[58] n29151_not ; n29152
g28897 and n668 n29108_not ; n29153
g28898 and n29152_not n29153_not ; n29154
g28899 and b[1] n29154_not ; n29155
g28900 and b[1]_not n29153_not ; n29156
g28901 and n29152_not n29156 ; n29157
g28902 and n29155_not n29157_not ; n29158
g28903 and n756_not n29158_not ; n29159
g28904 and b[1]_not n29154_not ; n29160
g28905 and n29159_not n29160_not ; n29161
g28906 and b[2] n29148_not ; n29162
g28907 and n29146_not n29162 ; n29163
g28908 and n29150_not n29163_not ; n29164
g28909 and n29161_not n29164 ; n29165
g28910 and n29150_not n29165_not ; n29166
g28911 and b[3] n29140_not ; n29167
g28912 and n29138_not n29167 ; n29168
g28913 and n29142_not n29168_not ; n29169
g28914 and n29166_not n29169 ; n29170
g28915 and n29142_not n29170_not ; n29171
g28916 and b[4] n29131_not ; n29172
g28917 and n29129_not n29172 ; n29173
g28918 and n29133_not n29173_not ; n29174
g28919 and n29171_not n29174 ; n29175
g28920 and n29133_not n29175_not ; n29176
g28921 and b[5] n29114_not ; n29177
g28922 and n29112_not n29177 ; n29178
g28923 and n29125_not n29178_not ; n29179
g28924 and n29176_not n29179 ; n29180
g28925 and n29125_not n29180_not ; n29181
g28926 and b[6] n29122_not ; n29182
g28927 and n29120_not n29182 ; n29183
g28928 and n29124_not n29183_not ; n29184
g28929 and n29181_not n29184 ; n29185
g28930 and n29124_not n29185_not ; n29186
g28931 and n788 n29186_not ; n29187
g28932 and n29115_not n29187_not ; n29188
g28933 and n29133_not n29179 ; n29189
g28934 and n29175_not n29189 ; n29190
g28935 and n29176_not n29179_not ; n29191
g28936 and n29190_not n29191_not ; n29192
g28937 and n788 n29192_not ; n29193
g28938 and n29186_not n29193 ; n29194
g28939 and n29188_not n29194_not ; n29195
g28940 and n29123_not n29187_not ; n29196
g28941 and n29125_not n29184 ; n29197
g28942 and n29180_not n29197 ; n29198
g28943 and n29181_not n29184_not ; n29199
g28944 and n29198_not n29199_not ; n29200
g28945 and n29187 n29200_not ; n29201
g28946 and n29196_not n29201_not ; n29202
g28947 and b[7]_not n29202_not ; n29203
g28948 and b[6]_not n29195_not ; n29204
g28949 and n29132_not n29187_not ; n29205
g28950 and n29142_not n29174 ; n29206
g28951 and n29170_not n29206 ; n29207
g28952 and n29171_not n29174_not ; n29208
g28953 and n29207_not n29208_not ; n29209
g28954 and n788 n29209_not ; n29210
g28955 and n29186_not n29210 ; n29211
g28956 and n29205_not n29211_not ; n29212
g28957 and b[5]_not n29212_not ; n29213
g28958 and n29141_not n29187_not ; n29214
g28959 and n29150_not n29169 ; n29215
g28960 and n29165_not n29215 ; n29216
g28961 and n29166_not n29169_not ; n29217
g28962 and n29216_not n29217_not ; n29218
g28963 and n788 n29218_not ; n29219
g28964 and n29186_not n29219 ; n29220
g28965 and n29214_not n29220_not ; n29221
g28966 and b[4]_not n29221_not ; n29222
g28967 and n29149_not n29187_not ; n29223
g28968 and n29160_not n29164 ; n29224
g28969 and n29159_not n29224 ; n29225
g28970 and n29161_not n29164_not ; n29226
g28971 and n29225_not n29226_not ; n29227
g28972 and n788 n29227_not ; n29228
g28973 and n29186_not n29228 ; n29229
g28974 and n29223_not n29229_not ; n29230
g28975 and b[3]_not n29230_not ; n29231
g28976 and n29154_not n29187_not ; n29232
g28977 and n756 n29157_not ; n29233
g28978 and n29155_not n29233 ; n29234
g28979 and n788 n29234_not ; n29235
g28980 and n29159_not n29235 ; n29236
g28981 and n29186_not n29236 ; n29237
g28982 and n29232_not n29237_not ; n29238
g28983 and b[2]_not n29238_not ; n29239
g28984 and n846 n29186_not ; n29240
g28985 and a[57] n29240_not ; n29241
g28986 and n853 n29186_not ; n29242
g28987 and n29241_not n29242_not ; n29243
g28988 and b[1] n29243_not ; n29244
g28989 and b[1]_not n29242_not ; n29245
g28990 and n29241_not n29245 ; n29246
g28991 and n29244_not n29246_not ; n29247
g28992 and n860_not n29247_not ; n29248
g28993 and b[1]_not n29243_not ; n29249
g28994 and n29248_not n29249_not ; n29250
g28995 and b[2] n29237_not ; n29251
g28996 and n29232_not n29251 ; n29252
g28997 and n29239_not n29252_not ; n29253
g28998 and n29250_not n29253 ; n29254
g28999 and n29239_not n29254_not ; n29255
g29000 and b[3] n29229_not ; n29256
g29001 and n29223_not n29256 ; n29257
g29002 and n29231_not n29257_not ; n29258
g29003 and n29255_not n29258 ; n29259
g29004 and n29231_not n29259_not ; n29260
g29005 and b[4] n29220_not ; n29261
g29006 and n29214_not n29261 ; n29262
g29007 and n29222_not n29262_not ; n29263
g29008 and n29260_not n29263 ; n29264
g29009 and n29222_not n29264_not ; n29265
g29010 and b[5] n29211_not ; n29266
g29011 and n29205_not n29266 ; n29267
g29012 and n29213_not n29267_not ; n29268
g29013 and n29265_not n29268 ; n29269
g29014 and n29213_not n29269_not ; n29270
g29015 and b[6] n29194_not ; n29271
g29016 and n29188_not n29271 ; n29272
g29017 and n29204_not n29272_not ; n29273
g29018 and n29270_not n29273 ; n29274
g29019 and n29204_not n29274_not ; n29275
g29020 and b[7] n29196_not ; n29276
g29021 and n29201_not n29276 ; n29277
g29022 and n29203_not n29277_not ; n29278
g29023 and n29275_not n29278 ; n29279
g29024 and n29203_not n29279_not ; n29280
g29025 and n895 n29280_not ; n29281
g29026 and n29195_not n29281_not ; n29282
g29027 and n29213_not n29273 ; n29283
g29028 and n29269_not n29283 ; n29284
g29029 and n29270_not n29273_not ; n29285
g29030 and n29284_not n29285_not ; n29286
g29031 and n895 n29286_not ; n29287
g29032 and n29280_not n29287 ; n29288
g29033 and n29282_not n29288_not ; n29289
g29034 and b[7]_not n29289_not ; n29290
g29035 and n29212_not n29281_not ; n29291
g29036 and n29222_not n29268 ; n29292
g29037 and n29264_not n29292 ; n29293
g29038 and n29265_not n29268_not ; n29294
g29039 and n29293_not n29294_not ; n29295
g29040 and n895 n29295_not ; n29296
g29041 and n29280_not n29296 ; n29297
g29042 and n29291_not n29297_not ; n29298
g29043 and b[6]_not n29298_not ; n29299
g29044 and n29221_not n29281_not ; n29300
g29045 and n29231_not n29263 ; n29301
g29046 and n29259_not n29301 ; n29302
g29047 and n29260_not n29263_not ; n29303
g29048 and n29302_not n29303_not ; n29304
g29049 and n895 n29304_not ; n29305
g29050 and n29280_not n29305 ; n29306
g29051 and n29300_not n29306_not ; n29307
g29052 and b[5]_not n29307_not ; n29308
g29053 and n29230_not n29281_not ; n29309
g29054 and n29239_not n29258 ; n29310
g29055 and n29254_not n29310 ; n29311
g29056 and n29255_not n29258_not ; n29312
g29057 and n29311_not n29312_not ; n29313
g29058 and n895 n29313_not ; n29314
g29059 and n29280_not n29314 ; n29315
g29060 and n29309_not n29315_not ; n29316
g29061 and b[4]_not n29316_not ; n29317
g29062 and n29238_not n29281_not ; n29318
g29063 and n29249_not n29253 ; n29319
g29064 and n29248_not n29319 ; n29320
g29065 and n29250_not n29253_not ; n29321
g29066 and n29320_not n29321_not ; n29322
g29067 and n895 n29322_not ; n29323
g29068 and n29280_not n29323 ; n29324
g29069 and n29318_not n29324_not ; n29325
g29070 and b[3]_not n29325_not ; n29326
g29071 and n29243_not n29281_not ; n29327
g29072 and n860 n29246_not ; n29328
g29073 and n29244_not n29328 ; n29329
g29074 and n895 n29329_not ; n29330
g29075 and n29248_not n29330 ; n29331
g29076 and n29280_not n29331 ; n29332
g29077 and n29327_not n29332_not ; n29333
g29078 and b[2]_not n29333_not ; n29334
g29079 and n954 n29280_not ; n29335
g29080 and a[56] n29335_not ; n29336
g29081 and n960 n29280_not ; n29337
g29082 and n29336_not n29337_not ; n29338
g29083 and b[1] n29338_not ; n29339
g29084 and b[1]_not n29337_not ; n29340
g29085 and n29336_not n29340 ; n29341
g29086 and n29339_not n29341_not ; n29342
g29087 and n967_not n29342_not ; n29343
g29088 and b[1]_not n29338_not ; n29344
g29089 and n29343_not n29344_not ; n29345
g29090 and b[2] n29332_not ; n29346
g29091 and n29327_not n29346 ; n29347
g29092 and n29334_not n29347_not ; n29348
g29093 and n29345_not n29348 ; n29349
g29094 and n29334_not n29349_not ; n29350
g29095 and b[3] n29324_not ; n29351
g29096 and n29318_not n29351 ; n29352
g29097 and n29326_not n29352_not ; n29353
g29098 and n29350_not n29353 ; n29354
g29099 and n29326_not n29354_not ; n29355
g29100 and b[4] n29315_not ; n29356
g29101 and n29309_not n29356 ; n29357
g29102 and n29317_not n29357_not ; n29358
g29103 and n29355_not n29358 ; n29359
g29104 and n29317_not n29359_not ; n29360
g29105 and b[5] n29306_not ; n29361
g29106 and n29300_not n29361 ; n29362
g29107 and n29308_not n29362_not ; n29363
g29108 and n29360_not n29363 ; n29364
g29109 and n29308_not n29364_not ; n29365
g29110 and b[6] n29297_not ; n29366
g29111 and n29291_not n29366 ; n29367
g29112 and n29299_not n29367_not ; n29368
g29113 and n29365_not n29368 ; n29369
g29114 and n29299_not n29369_not ; n29370
g29115 and b[7] n29288_not ; n29371
g29116 and n29282_not n29371 ; n29372
g29117 and n29290_not n29372_not ; n29373
g29118 and n29370_not n29373 ; n29374
g29119 and n29290_not n29374_not ; n29375
g29120 and n29202_not n29281_not ; n29376
g29121 and n29204_not n29278 ; n29377
g29122 and n29274_not n29377 ; n29378
g29123 and n29275_not n29278_not ; n29379
g29124 and n29378_not n29379_not ; n29380
g29125 and n29281 n29380_not ; n29381
g29126 and n29376_not n29381_not ; n29382
g29127 and b[8]_not n29382_not ; n29383
g29128 and b[8] n29376_not ; n29384
g29129 and n29381_not n29384 ; n29385
g29130 and n1012 n29385_not ; n29386
g29131 and n29383_not n29386 ; n29387
g29132 and n29375_not n29387 ; n29388
g29133 and n895 n29382_not ; n29389
g29134 and n29388_not n29389_not ; n29390
g29135 and n29299_not n29373 ; n29391
g29136 and n29369_not n29391 ; n29392
g29137 and n29370_not n29373_not ; n29393
g29138 and n29392_not n29393_not ; n29394
g29139 and n29390_not n29394_not ; n29395
g29140 and n29289_not n29389_not ; n29396
g29141 and n29388_not n29396 ; n29397
g29142 and n29395_not n29397_not ; n29398
g29143 and n29290_not n29385_not ; n29399
g29144 and n29383_not n29399 ; n29400
g29145 and n29374_not n29400 ; n29401
g29146 and n29383_not n29385_not ; n29402
g29147 and n29375_not n29402_not ; n29403
g29148 and n29401_not n29403_not ; n29404
g29149 and n29390_not n29404_not ; n29405
g29150 and n29382_not n29389_not ; n29406
g29151 and n29388_not n29406 ; n29407
g29152 and n29405_not n29407_not ; n29408
g29153 and b[9]_not n29408_not ; n29409
g29154 and b[8]_not n29398_not ; n29410
g29155 and n29308_not n29368 ; n29411
g29156 and n29364_not n29411 ; n29412
g29157 and n29365_not n29368_not ; n29413
g29158 and n29412_not n29413_not ; n29414
g29159 and n29390_not n29414_not ; n29415
g29160 and n29298_not n29389_not ; n29416
g29161 and n29388_not n29416 ; n29417
g29162 and n29415_not n29417_not ; n29418
g29163 and b[7]_not n29418_not ; n29419
g29164 and n29317_not n29363 ; n29420
g29165 and n29359_not n29420 ; n29421
g29166 and n29360_not n29363_not ; n29422
g29167 and n29421_not n29422_not ; n29423
g29168 and n29390_not n29423_not ; n29424
g29169 and n29307_not n29389_not ; n29425
g29170 and n29388_not n29425 ; n29426
g29171 and n29424_not n29426_not ; n29427
g29172 and b[6]_not n29427_not ; n29428
g29173 and n29326_not n29358 ; n29429
g29174 and n29354_not n29429 ; n29430
g29175 and n29355_not n29358_not ; n29431
g29176 and n29430_not n29431_not ; n29432
g29177 and n29390_not n29432_not ; n29433
g29178 and n29316_not n29389_not ; n29434
g29179 and n29388_not n29434 ; n29435
g29180 and n29433_not n29435_not ; n29436
g29181 and b[5]_not n29436_not ; n29437
g29182 and n29334_not n29353 ; n29438
g29183 and n29349_not n29438 ; n29439
g29184 and n29350_not n29353_not ; n29440
g29185 and n29439_not n29440_not ; n29441
g29186 and n29390_not n29441_not ; n29442
g29187 and n29325_not n29389_not ; n29443
g29188 and n29388_not n29443 ; n29444
g29189 and n29442_not n29444_not ; n29445
g29190 and b[4]_not n29445_not ; n29446
g29191 and n29344_not n29348 ; n29447
g29192 and n29343_not n29447 ; n29448
g29193 and n29345_not n29348_not ; n29449
g29194 and n29448_not n29449_not ; n29450
g29195 and n29390_not n29450_not ; n29451
g29196 and n29333_not n29389_not ; n29452
g29197 and n29388_not n29452 ; n29453
g29198 and n29451_not n29453_not ; n29454
g29199 and b[3]_not n29454_not ; n29455
g29200 and n967 n29341_not ; n29456
g29201 and n29339_not n29456 ; n29457
g29202 and n29343_not n29457_not ; n29458
g29203 and n29390_not n29458 ; n29459
g29204 and n29338_not n29389_not ; n29460
g29205 and n29388_not n29460 ; n29461
g29206 and n29459_not n29461_not ; n29462
g29207 and b[2]_not n29462_not ; n29463
g29208 and b[0] n29390_not ; n29464
g29209 and a[55] n29464_not ; n29465
g29210 and n967 n29390_not ; n29466
g29211 and n29465_not n29466_not ; n29467
g29212 and b[1] n29467_not ; n29468
g29213 and b[1]_not n29466_not ; n29469
g29214 and n29465_not n29469 ; n29470
g29215 and n29468_not n29470_not ; n29471
g29216 and n1099_not n29471_not ; n29472
g29217 and b[1]_not n29467_not ; n29473
g29218 and n29472_not n29473_not ; n29474
g29219 and b[2] n29461_not ; n29475
g29220 and n29459_not n29475 ; n29476
g29221 and n29463_not n29476_not ; n29477
g29222 and n29474_not n29477 ; n29478
g29223 and n29463_not n29478_not ; n29479
g29224 and b[3] n29453_not ; n29480
g29225 and n29451_not n29480 ; n29481
g29226 and n29455_not n29481_not ; n29482
g29227 and n29479_not n29482 ; n29483
g29228 and n29455_not n29483_not ; n29484
g29229 and b[4] n29444_not ; n29485
g29230 and n29442_not n29485 ; n29486
g29231 and n29446_not n29486_not ; n29487
g29232 and n29484_not n29487 ; n29488
g29233 and n29446_not n29488_not ; n29489
g29234 and b[5] n29435_not ; n29490
g29235 and n29433_not n29490 ; n29491
g29236 and n29437_not n29491_not ; n29492
g29237 and n29489_not n29492 ; n29493
g29238 and n29437_not n29493_not ; n29494
g29239 and b[6] n29426_not ; n29495
g29240 and n29424_not n29495 ; n29496
g29241 and n29428_not n29496_not ; n29497
g29242 and n29494_not n29497 ; n29498
g29243 and n29428_not n29498_not ; n29499
g29244 and b[7] n29417_not ; n29500
g29245 and n29415_not n29500 ; n29501
g29246 and n29419_not n29501_not ; n29502
g29247 and n29499_not n29502 ; n29503
g29248 and n29419_not n29503_not ; n29504
g29249 and b[8] n29397_not ; n29505
g29250 and n29395_not n29505 ; n29506
g29251 and n29410_not n29506_not ; n29507
g29252 and n29504_not n29507 ; n29508
g29253 and n29410_not n29508_not ; n29509
g29254 and b[9] n29407_not ; n29510
g29255 and n29405_not n29510 ; n29511
g29256 and n29409_not n29511_not ; n29512
g29257 and n29509_not n29512 ; n29513
g29258 and n29409_not n29513_not ; n29514
g29259 and n1145 n29514_not ; n29515
g29260 and n29398_not n29515_not ; n29516
g29261 and n29419_not n29507 ; n29517
g29262 and n29503_not n29517 ; n29518
g29263 and n29504_not n29507_not ; n29519
g29264 and n29518_not n29519_not ; n29520
g29265 and n1145 n29520_not ; n29521
g29266 and n29514_not n29521 ; n29522
g29267 and n29516_not n29522_not ; n29523
g29268 and n29408_not n29515_not ; n29524
g29269 and n29410_not n29512 ; n29525
g29270 and n29508_not n29525 ; n29526
g29271 and n29509_not n29512_not ; n29527
g29272 and n29526_not n29527_not ; n29528
g29273 and n29515 n29528_not ; n29529
g29274 and n29524_not n29529_not ; n29530
g29275 and b[10]_not n29530_not ; n29531
g29276 and b[9]_not n29523_not ; n29532
g29277 and n29418_not n29515_not ; n29533
g29278 and n29428_not n29502 ; n29534
g29279 and n29498_not n29534 ; n29535
g29280 and n29499_not n29502_not ; n29536
g29281 and n29535_not n29536_not ; n29537
g29282 and n1145 n29537_not ; n29538
g29283 and n29514_not n29538 ; n29539
g29284 and n29533_not n29539_not ; n29540
g29285 and b[8]_not n29540_not ; n29541
g29286 and n29427_not n29515_not ; n29542
g29287 and n29437_not n29497 ; n29543
g29288 and n29493_not n29543 ; n29544
g29289 and n29494_not n29497_not ; n29545
g29290 and n29544_not n29545_not ; n29546
g29291 and n1145 n29546_not ; n29547
g29292 and n29514_not n29547 ; n29548
g29293 and n29542_not n29548_not ; n29549
g29294 and b[7]_not n29549_not ; n29550
g29295 and n29436_not n29515_not ; n29551
g29296 and n29446_not n29492 ; n29552
g29297 and n29488_not n29552 ; n29553
g29298 and n29489_not n29492_not ; n29554
g29299 and n29553_not n29554_not ; n29555
g29300 and n1145 n29555_not ; n29556
g29301 and n29514_not n29556 ; n29557
g29302 and n29551_not n29557_not ; n29558
g29303 and b[6]_not n29558_not ; n29559
g29304 and n29445_not n29515_not ; n29560
g29305 and n29455_not n29487 ; n29561
g29306 and n29483_not n29561 ; n29562
g29307 and n29484_not n29487_not ; n29563
g29308 and n29562_not n29563_not ; n29564
g29309 and n1145 n29564_not ; n29565
g29310 and n29514_not n29565 ; n29566
g29311 and n29560_not n29566_not ; n29567
g29312 and b[5]_not n29567_not ; n29568
g29313 and n29454_not n29515_not ; n29569
g29314 and n29463_not n29482 ; n29570
g29315 and n29478_not n29570 ; n29571
g29316 and n29479_not n29482_not ; n29572
g29317 and n29571_not n29572_not ; n29573
g29318 and n1145 n29573_not ; n29574
g29319 and n29514_not n29574 ; n29575
g29320 and n29569_not n29575_not ; n29576
g29321 and b[4]_not n29576_not ; n29577
g29322 and n29462_not n29515_not ; n29578
g29323 and n29473_not n29477 ; n29579
g29324 and n29472_not n29579 ; n29580
g29325 and n29474_not n29477_not ; n29581
g29326 and n29580_not n29581_not ; n29582
g29327 and n1145 n29582_not ; n29583
g29328 and n29514_not n29583 ; n29584
g29329 and n29578_not n29584_not ; n29585
g29330 and b[3]_not n29585_not ; n29586
g29331 and n29467_not n29515_not ; n29587
g29332 and n1099 n29470_not ; n29588
g29333 and n29468_not n29588 ; n29589
g29334 and n1145 n29589_not ; n29590
g29335 and n29472_not n29590 ; n29591
g29336 and n29514_not n29591 ; n29592
g29337 and n29587_not n29592_not ; n29593
g29338 and b[2]_not n29593_not ; n29594
g29339 and n1230 n29514_not ; n29595
g29340 and a[54] n29595_not ; n29596
g29341 and n1236 n29514_not ; n29597
g29342 and n29596_not n29597_not ; n29598
g29343 and b[1] n29598_not ; n29599
g29344 and b[1]_not n29597_not ; n29600
g29345 and n29596_not n29600 ; n29601
g29346 and n29599_not n29601_not ; n29602
g29347 and n1243_not n29602_not ; n29603
g29348 and b[1]_not n29598_not ; n29604
g29349 and n29603_not n29604_not ; n29605
g29350 and b[2] n29592_not ; n29606
g29351 and n29587_not n29606 ; n29607
g29352 and n29594_not n29607_not ; n29608
g29353 and n29605_not n29608 ; n29609
g29354 and n29594_not n29609_not ; n29610
g29355 and b[3] n29584_not ; n29611
g29356 and n29578_not n29611 ; n29612
g29357 and n29586_not n29612_not ; n29613
g29358 and n29610_not n29613 ; n29614
g29359 and n29586_not n29614_not ; n29615
g29360 and b[4] n29575_not ; n29616
g29361 and n29569_not n29616 ; n29617
g29362 and n29577_not n29617_not ; n29618
g29363 and n29615_not n29618 ; n29619
g29364 and n29577_not n29619_not ; n29620
g29365 and b[5] n29566_not ; n29621
g29366 and n29560_not n29621 ; n29622
g29367 and n29568_not n29622_not ; n29623
g29368 and n29620_not n29623 ; n29624
g29369 and n29568_not n29624_not ; n29625
g29370 and b[6] n29557_not ; n29626
g29371 and n29551_not n29626 ; n29627
g29372 and n29559_not n29627_not ; n29628
g29373 and n29625_not n29628 ; n29629
g29374 and n29559_not n29629_not ; n29630
g29375 and b[7] n29548_not ; n29631
g29376 and n29542_not n29631 ; n29632
g29377 and n29550_not n29632_not ; n29633
g29378 and n29630_not n29633 ; n29634
g29379 and n29550_not n29634_not ; n29635
g29380 and b[8] n29539_not ; n29636
g29381 and n29533_not n29636 ; n29637
g29382 and n29541_not n29637_not ; n29638
g29383 and n29635_not n29638 ; n29639
g29384 and n29541_not n29639_not ; n29640
g29385 and b[9] n29522_not ; n29641
g29386 and n29516_not n29641 ; n29642
g29387 and n29532_not n29642_not ; n29643
g29388 and n29640_not n29643 ; n29644
g29389 and n29532_not n29644_not ; n29645
g29390 and b[10] n29524_not ; n29646
g29391 and n29529_not n29646 ; n29647
g29392 and n29531_not n29647_not ; n29648
g29393 and n29645_not n29648 ; n29649
g29394 and n29531_not n29649_not ; n29650
g29395 and n1294 n29650_not ; n29651
g29396 and n29523_not n29651_not ; n29652
g29397 and n29541_not n29643 ; n29653
g29398 and n29639_not n29653 ; n29654
g29399 and n29640_not n29643_not ; n29655
g29400 and n29654_not n29655_not ; n29656
g29401 and n1294 n29656_not ; n29657
g29402 and n29650_not n29657 ; n29658
g29403 and n29652_not n29658_not ; n29659
g29404 and b[10]_not n29659_not ; n29660
g29405 and n29540_not n29651_not ; n29661
g29406 and n29550_not n29638 ; n29662
g29407 and n29634_not n29662 ; n29663
g29408 and n29635_not n29638_not ; n29664
g29409 and n29663_not n29664_not ; n29665
g29410 and n1294 n29665_not ; n29666
g29411 and n29650_not n29666 ; n29667
g29412 and n29661_not n29667_not ; n29668
g29413 and b[9]_not n29668_not ; n29669
g29414 and n29549_not n29651_not ; n29670
g29415 and n29559_not n29633 ; n29671
g29416 and n29629_not n29671 ; n29672
g29417 and n29630_not n29633_not ; n29673
g29418 and n29672_not n29673_not ; n29674
g29419 and n1294 n29674_not ; n29675
g29420 and n29650_not n29675 ; n29676
g29421 and n29670_not n29676_not ; n29677
g29422 and b[8]_not n29677_not ; n29678
g29423 and n29558_not n29651_not ; n29679
g29424 and n29568_not n29628 ; n29680
g29425 and n29624_not n29680 ; n29681
g29426 and n29625_not n29628_not ; n29682
g29427 and n29681_not n29682_not ; n29683
g29428 and n1294 n29683_not ; n29684
g29429 and n29650_not n29684 ; n29685
g29430 and n29679_not n29685_not ; n29686
g29431 and b[7]_not n29686_not ; n29687
g29432 and n29567_not n29651_not ; n29688
g29433 and n29577_not n29623 ; n29689
g29434 and n29619_not n29689 ; n29690
g29435 and n29620_not n29623_not ; n29691
g29436 and n29690_not n29691_not ; n29692
g29437 and n1294 n29692_not ; n29693
g29438 and n29650_not n29693 ; n29694
g29439 and n29688_not n29694_not ; n29695
g29440 and b[6]_not n29695_not ; n29696
g29441 and n29576_not n29651_not ; n29697
g29442 and n29586_not n29618 ; n29698
g29443 and n29614_not n29698 ; n29699
g29444 and n29615_not n29618_not ; n29700
g29445 and n29699_not n29700_not ; n29701
g29446 and n1294 n29701_not ; n29702
g29447 and n29650_not n29702 ; n29703
g29448 and n29697_not n29703_not ; n29704
g29449 and b[5]_not n29704_not ; n29705
g29450 and n29585_not n29651_not ; n29706
g29451 and n29594_not n29613 ; n29707
g29452 and n29609_not n29707 ; n29708
g29453 and n29610_not n29613_not ; n29709
g29454 and n29708_not n29709_not ; n29710
g29455 and n1294 n29710_not ; n29711
g29456 and n29650_not n29711 ; n29712
g29457 and n29706_not n29712_not ; n29713
g29458 and b[4]_not n29713_not ; n29714
g29459 and n29593_not n29651_not ; n29715
g29460 and n29604_not n29608 ; n29716
g29461 and n29603_not n29716 ; n29717
g29462 and n29605_not n29608_not ; n29718
g29463 and n29717_not n29718_not ; n29719
g29464 and n1294 n29719_not ; n29720
g29465 and n29650_not n29720 ; n29721
g29466 and n29715_not n29721_not ; n29722
g29467 and b[3]_not n29722_not ; n29723
g29468 and n29598_not n29651_not ; n29724
g29469 and n1243 n29601_not ; n29725
g29470 and n29599_not n29725 ; n29726
g29471 and n1294 n29726_not ; n29727
g29472 and n29603_not n29727 ; n29728
g29473 and n29650_not n29728 ; n29729
g29474 and n29724_not n29729_not ; n29730
g29475 and b[2]_not n29730_not ; n29731
g29476 and n1379 n29650_not ; n29732
g29477 and a[53] n29732_not ; n29733
g29478 and n1385 n29650_not ; n29734
g29479 and n29733_not n29734_not ; n29735
g29480 and b[1] n29735_not ; n29736
g29481 and b[1]_not n29734_not ; n29737
g29482 and n29733_not n29737 ; n29738
g29483 and n29736_not n29738_not ; n29739
g29484 and n1392_not n29739_not ; n29740
g29485 and b[1]_not n29735_not ; n29741
g29486 and n29740_not n29741_not ; n29742
g29487 and b[2] n29729_not ; n29743
g29488 and n29724_not n29743 ; n29744
g29489 and n29731_not n29744_not ; n29745
g29490 and n29742_not n29745 ; n29746
g29491 and n29731_not n29746_not ; n29747
g29492 and b[3] n29721_not ; n29748
g29493 and n29715_not n29748 ; n29749
g29494 and n29723_not n29749_not ; n29750
g29495 and n29747_not n29750 ; n29751
g29496 and n29723_not n29751_not ; n29752
g29497 and b[4] n29712_not ; n29753
g29498 and n29706_not n29753 ; n29754
g29499 and n29714_not n29754_not ; n29755
g29500 and n29752_not n29755 ; n29756
g29501 and n29714_not n29756_not ; n29757
g29502 and b[5] n29703_not ; n29758
g29503 and n29697_not n29758 ; n29759
g29504 and n29705_not n29759_not ; n29760
g29505 and n29757_not n29760 ; n29761
g29506 and n29705_not n29761_not ; n29762
g29507 and b[6] n29694_not ; n29763
g29508 and n29688_not n29763 ; n29764
g29509 and n29696_not n29764_not ; n29765
g29510 and n29762_not n29765 ; n29766
g29511 and n29696_not n29766_not ; n29767
g29512 and b[7] n29685_not ; n29768
g29513 and n29679_not n29768 ; n29769
g29514 and n29687_not n29769_not ; n29770
g29515 and n29767_not n29770 ; n29771
g29516 and n29687_not n29771_not ; n29772
g29517 and b[8] n29676_not ; n29773
g29518 and n29670_not n29773 ; n29774
g29519 and n29678_not n29774_not ; n29775
g29520 and n29772_not n29775 ; n29776
g29521 and n29678_not n29776_not ; n29777
g29522 and b[9] n29667_not ; n29778
g29523 and n29661_not n29778 ; n29779
g29524 and n29669_not n29779_not ; n29780
g29525 and n29777_not n29780 ; n29781
g29526 and n29669_not n29781_not ; n29782
g29527 and b[10] n29658_not ; n29783
g29528 and n29652_not n29783 ; n29784
g29529 and n29660_not n29784_not ; n29785
g29530 and n29782_not n29785 ; n29786
g29531 and n29660_not n29786_not ; n29787
g29532 and n29530_not n29651_not ; n29788
g29533 and n29532_not n29648 ; n29789
g29534 and n29644_not n29789 ; n29790
g29535 and n29645_not n29648_not ; n29791
g29536 and n29790_not n29791_not ; n29792
g29537 and n29651 n29792_not ; n29793
g29538 and n29788_not n29793_not ; n29794
g29539 and b[11]_not n29794_not ; n29795
g29540 and b[11] n29788_not ; n29796
g29541 and n29793_not n29796 ; n29797
g29542 and n1452 n29797_not ; n29798
g29543 and n29795_not n29798 ; n29799
g29544 and n29787_not n29799 ; n29800
g29545 and n1294 n29794_not ; n29801
g29546 and n29800_not n29801_not ; n29802
g29547 and n29669_not n29785 ; n29803
g29548 and n29781_not n29803 ; n29804
g29549 and n29782_not n29785_not ; n29805
g29550 and n29804_not n29805_not ; n29806
g29551 and n29802_not n29806_not ; n29807
g29552 and n29659_not n29801_not ; n29808
g29553 and n29800_not n29808 ; n29809
g29554 and n29807_not n29809_not ; n29810
g29555 and n29660_not n29797_not ; n29811
g29556 and n29795_not n29811 ; n29812
g29557 and n29786_not n29812 ; n29813
g29558 and n29795_not n29797_not ; n29814
g29559 and n29787_not n29814_not ; n29815
g29560 and n29813_not n29815_not ; n29816
g29561 and n29802_not n29816_not ; n29817
g29562 and n29794_not n29801_not ; n29818
g29563 and n29800_not n29818 ; n29819
g29564 and n29817_not n29819_not ; n29820
g29565 and b[12]_not n29820_not ; n29821
g29566 and b[11]_not n29810_not ; n29822
g29567 and n29678_not n29780 ; n29823
g29568 and n29776_not n29823 ; n29824
g29569 and n29777_not n29780_not ; n29825
g29570 and n29824_not n29825_not ; n29826
g29571 and n29802_not n29826_not ; n29827
g29572 and n29668_not n29801_not ; n29828
g29573 and n29800_not n29828 ; n29829
g29574 and n29827_not n29829_not ; n29830
g29575 and b[10]_not n29830_not ; n29831
g29576 and n29687_not n29775 ; n29832
g29577 and n29771_not n29832 ; n29833
g29578 and n29772_not n29775_not ; n29834
g29579 and n29833_not n29834_not ; n29835
g29580 and n29802_not n29835_not ; n29836
g29581 and n29677_not n29801_not ; n29837
g29582 and n29800_not n29837 ; n29838
g29583 and n29836_not n29838_not ; n29839
g29584 and b[9]_not n29839_not ; n29840
g29585 and n29696_not n29770 ; n29841
g29586 and n29766_not n29841 ; n29842
g29587 and n29767_not n29770_not ; n29843
g29588 and n29842_not n29843_not ; n29844
g29589 and n29802_not n29844_not ; n29845
g29590 and n29686_not n29801_not ; n29846
g29591 and n29800_not n29846 ; n29847
g29592 and n29845_not n29847_not ; n29848
g29593 and b[8]_not n29848_not ; n29849
g29594 and n29705_not n29765 ; n29850
g29595 and n29761_not n29850 ; n29851
g29596 and n29762_not n29765_not ; n29852
g29597 and n29851_not n29852_not ; n29853
g29598 and n29802_not n29853_not ; n29854
g29599 and n29695_not n29801_not ; n29855
g29600 and n29800_not n29855 ; n29856
g29601 and n29854_not n29856_not ; n29857
g29602 and b[7]_not n29857_not ; n29858
g29603 and n29714_not n29760 ; n29859
g29604 and n29756_not n29859 ; n29860
g29605 and n29757_not n29760_not ; n29861
g29606 and n29860_not n29861_not ; n29862
g29607 and n29802_not n29862_not ; n29863
g29608 and n29704_not n29801_not ; n29864
g29609 and n29800_not n29864 ; n29865
g29610 and n29863_not n29865_not ; n29866
g29611 and b[6]_not n29866_not ; n29867
g29612 and n29723_not n29755 ; n29868
g29613 and n29751_not n29868 ; n29869
g29614 and n29752_not n29755_not ; n29870
g29615 and n29869_not n29870_not ; n29871
g29616 and n29802_not n29871_not ; n29872
g29617 and n29713_not n29801_not ; n29873
g29618 and n29800_not n29873 ; n29874
g29619 and n29872_not n29874_not ; n29875
g29620 and b[5]_not n29875_not ; n29876
g29621 and n29731_not n29750 ; n29877
g29622 and n29746_not n29877 ; n29878
g29623 and n29747_not n29750_not ; n29879
g29624 and n29878_not n29879_not ; n29880
g29625 and n29802_not n29880_not ; n29881
g29626 and n29722_not n29801_not ; n29882
g29627 and n29800_not n29882 ; n29883
g29628 and n29881_not n29883_not ; n29884
g29629 and b[4]_not n29884_not ; n29885
g29630 and n29741_not n29745 ; n29886
g29631 and n29740_not n29886 ; n29887
g29632 and n29742_not n29745_not ; n29888
g29633 and n29887_not n29888_not ; n29889
g29634 and n29802_not n29889_not ; n29890
g29635 and n29730_not n29801_not ; n29891
g29636 and n29800_not n29891 ; n29892
g29637 and n29890_not n29892_not ; n29893
g29638 and b[3]_not n29893_not ; n29894
g29639 and n1392 n29738_not ; n29895
g29640 and n29736_not n29895 ; n29896
g29641 and n29740_not n29896_not ; n29897
g29642 and n29802_not n29897 ; n29898
g29643 and n29735_not n29801_not ; n29899
g29644 and n29800_not n29899 ; n29900
g29645 and n29898_not n29900_not ; n29901
g29646 and b[2]_not n29901_not ; n29902
g29647 and b[0] n29802_not ; n29903
g29648 and a[52] n29903_not ; n29904
g29649 and n1392 n29802_not ; n29905
g29650 and n29904_not n29905_not ; n29906
g29651 and b[1] n29906_not ; n29907
g29652 and b[1]_not n29905_not ; n29908
g29653 and n29904_not n29908 ; n29909
g29654 and n29907_not n29909_not ; n29910
g29655 and n1566_not n29910_not ; n29911
g29656 and b[1]_not n29906_not ; n29912
g29657 and n29911_not n29912_not ; n29913
g29658 and b[2] n29900_not ; n29914
g29659 and n29898_not n29914 ; n29915
g29660 and n29902_not n29915_not ; n29916
g29661 and n29913_not n29916 ; n29917
g29662 and n29902_not n29917_not ; n29918
g29663 and b[3] n29892_not ; n29919
g29664 and n29890_not n29919 ; n29920
g29665 and n29894_not n29920_not ; n29921
g29666 and n29918_not n29921 ; n29922
g29667 and n29894_not n29922_not ; n29923
g29668 and b[4] n29883_not ; n29924
g29669 and n29881_not n29924 ; n29925
g29670 and n29885_not n29925_not ; n29926
g29671 and n29923_not n29926 ; n29927
g29672 and n29885_not n29927_not ; n29928
g29673 and b[5] n29874_not ; n29929
g29674 and n29872_not n29929 ; n29930
g29675 and n29876_not n29930_not ; n29931
g29676 and n29928_not n29931 ; n29932
g29677 and n29876_not n29932_not ; n29933
g29678 and b[6] n29865_not ; n29934
g29679 and n29863_not n29934 ; n29935
g29680 and n29867_not n29935_not ; n29936
g29681 and n29933_not n29936 ; n29937
g29682 and n29867_not n29937_not ; n29938
g29683 and b[7] n29856_not ; n29939
g29684 and n29854_not n29939 ; n29940
g29685 and n29858_not n29940_not ; n29941
g29686 and n29938_not n29941 ; n29942
g29687 and n29858_not n29942_not ; n29943
g29688 and b[8] n29847_not ; n29944
g29689 and n29845_not n29944 ; n29945
g29690 and n29849_not n29945_not ; n29946
g29691 and n29943_not n29946 ; n29947
g29692 and n29849_not n29947_not ; n29948
g29693 and b[9] n29838_not ; n29949
g29694 and n29836_not n29949 ; n29950
g29695 and n29840_not n29950_not ; n29951
g29696 and n29948_not n29951 ; n29952
g29697 and n29840_not n29952_not ; n29953
g29698 and b[10] n29829_not ; n29954
g29699 and n29827_not n29954 ; n29955
g29700 and n29831_not n29955_not ; n29956
g29701 and n29953_not n29956 ; n29957
g29702 and n29831_not n29957_not ; n29958
g29703 and b[11] n29809_not ; n29959
g29704 and n29807_not n29959 ; n29960
g29705 and n29822_not n29960_not ; n29961
g29706 and n29958_not n29961 ; n29962
g29707 and n29822_not n29962_not ; n29963
g29708 and b[12] n29819_not ; n29964
g29709 and n29817_not n29964 ; n29965
g29710 and n29821_not n29965_not ; n29966
g29711 and n29963_not n29966 ; n29967
g29712 and n29821_not n29967_not ; n29968
g29713 and n1626 n29968_not ; n29969
g29714 and n29810_not n29969_not ; n29970
g29715 and n29831_not n29961 ; n29971
g29716 and n29957_not n29971 ; n29972
g29717 and n29958_not n29961_not ; n29973
g29718 and n29972_not n29973_not ; n29974
g29719 and n1626 n29974_not ; n29975
g29720 and n29968_not n29975 ; n29976
g29721 and n29970_not n29976_not ; n29977
g29722 and n29820_not n29969_not ; n29978
g29723 and n29822_not n29966 ; n29979
g29724 and n29962_not n29979 ; n29980
g29725 and n29963_not n29966_not ; n29981
g29726 and n29980_not n29981_not ; n29982
g29727 and n29969 n29982_not ; n29983
g29728 and n29978_not n29983_not ; n29984
g29729 and b[13]_not n29984_not ; n29985
g29730 and b[12]_not n29977_not ; n29986
g29731 and n29830_not n29969_not ; n29987
g29732 and n29840_not n29956 ; n29988
g29733 and n29952_not n29988 ; n29989
g29734 and n29953_not n29956_not ; n29990
g29735 and n29989_not n29990_not ; n29991
g29736 and n1626 n29991_not ; n29992
g29737 and n29968_not n29992 ; n29993
g29738 and n29987_not n29993_not ; n29994
g29739 and b[11]_not n29994_not ; n29995
g29740 and n29839_not n29969_not ; n29996
g29741 and n29849_not n29951 ; n29997
g29742 and n29947_not n29997 ; n29998
g29743 and n29948_not n29951_not ; n29999
g29744 and n29998_not n29999_not ; n30000
g29745 and n1626 n30000_not ; n30001
g29746 and n29968_not n30001 ; n30002
g29747 and n29996_not n30002_not ; n30003
g29748 and b[10]_not n30003_not ; n30004
g29749 and n29848_not n29969_not ; n30005
g29750 and n29858_not n29946 ; n30006
g29751 and n29942_not n30006 ; n30007
g29752 and n29943_not n29946_not ; n30008
g29753 and n30007_not n30008_not ; n30009
g29754 and n1626 n30009_not ; n30010
g29755 and n29968_not n30010 ; n30011
g29756 and n30005_not n30011_not ; n30012
g29757 and b[9]_not n30012_not ; n30013
g29758 and n29857_not n29969_not ; n30014
g29759 and n29867_not n29941 ; n30015
g29760 and n29937_not n30015 ; n30016
g29761 and n29938_not n29941_not ; n30017
g29762 and n30016_not n30017_not ; n30018
g29763 and n1626 n30018_not ; n30019
g29764 and n29968_not n30019 ; n30020
g29765 and n30014_not n30020_not ; n30021
g29766 and b[8]_not n30021_not ; n30022
g29767 and n29866_not n29969_not ; n30023
g29768 and n29876_not n29936 ; n30024
g29769 and n29932_not n30024 ; n30025
g29770 and n29933_not n29936_not ; n30026
g29771 and n30025_not n30026_not ; n30027
g29772 and n1626 n30027_not ; n30028
g29773 and n29968_not n30028 ; n30029
g29774 and n30023_not n30029_not ; n30030
g29775 and b[7]_not n30030_not ; n30031
g29776 and n29875_not n29969_not ; n30032
g29777 and n29885_not n29931 ; n30033
g29778 and n29927_not n30033 ; n30034
g29779 and n29928_not n29931_not ; n30035
g29780 and n30034_not n30035_not ; n30036
g29781 and n1626 n30036_not ; n30037
g29782 and n29968_not n30037 ; n30038
g29783 and n30032_not n30038_not ; n30039
g29784 and b[6]_not n30039_not ; n30040
g29785 and n29884_not n29969_not ; n30041
g29786 and n29894_not n29926 ; n30042
g29787 and n29922_not n30042 ; n30043
g29788 and n29923_not n29926_not ; n30044
g29789 and n30043_not n30044_not ; n30045
g29790 and n1626 n30045_not ; n30046
g29791 and n29968_not n30046 ; n30047
g29792 and n30041_not n30047_not ; n30048
g29793 and b[5]_not n30048_not ; n30049
g29794 and n29893_not n29969_not ; n30050
g29795 and n29902_not n29921 ; n30051
g29796 and n29917_not n30051 ; n30052
g29797 and n29918_not n29921_not ; n30053
g29798 and n30052_not n30053_not ; n30054
g29799 and n1626 n30054_not ; n30055
g29800 and n29968_not n30055 ; n30056
g29801 and n30050_not n30056_not ; n30057
g29802 and b[4]_not n30057_not ; n30058
g29803 and n29901_not n29969_not ; n30059
g29804 and n29912_not n29916 ; n30060
g29805 and n29911_not n30060 ; n30061
g29806 and n29913_not n29916_not ; n30062
g29807 and n30061_not n30062_not ; n30063
g29808 and n1626 n30063_not ; n30064
g29809 and n29968_not n30064 ; n30065
g29810 and n30059_not n30065_not ; n30066
g29811 and b[3]_not n30066_not ; n30067
g29812 and n29906_not n29969_not ; n30068
g29813 and n1566 n29909_not ; n30069
g29814 and n29907_not n30069 ; n30070
g29815 and n1626 n30070_not ; n30071
g29816 and n29911_not n30071 ; n30072
g29817 and n29968_not n30072 ; n30073
g29818 and n30068_not n30073_not ; n30074
g29819 and b[2]_not n30074_not ; n30075
g29820 and n1738 n29968_not ; n30076
g29821 and a[51] n30076_not ; n30077
g29822 and n1743 n29968_not ; n30078
g29823 and n30077_not n30078_not ; n30079
g29824 and b[1] n30079_not ; n30080
g29825 and b[1]_not n30078_not ; n30081
g29826 and n30077_not n30081 ; n30082
g29827 and n30080_not n30082_not ; n30083
g29828 and n1750_not n30083_not ; n30084
g29829 and b[1]_not n30079_not ; n30085
g29830 and n30084_not n30085_not ; n30086
g29831 and b[2] n30073_not ; n30087
g29832 and n30068_not n30087 ; n30088
g29833 and n30075_not n30088_not ; n30089
g29834 and n30086_not n30089 ; n30090
g29835 and n30075_not n30090_not ; n30091
g29836 and b[3] n30065_not ; n30092
g29837 and n30059_not n30092 ; n30093
g29838 and n30067_not n30093_not ; n30094
g29839 and n30091_not n30094 ; n30095
g29840 and n30067_not n30095_not ; n30096
g29841 and b[4] n30056_not ; n30097
g29842 and n30050_not n30097 ; n30098
g29843 and n30058_not n30098_not ; n30099
g29844 and n30096_not n30099 ; n30100
g29845 and n30058_not n30100_not ; n30101
g29846 and b[5] n30047_not ; n30102
g29847 and n30041_not n30102 ; n30103
g29848 and n30049_not n30103_not ; n30104
g29849 and n30101_not n30104 ; n30105
g29850 and n30049_not n30105_not ; n30106
g29851 and b[6] n30038_not ; n30107
g29852 and n30032_not n30107 ; n30108
g29853 and n30040_not n30108_not ; n30109
g29854 and n30106_not n30109 ; n30110
g29855 and n30040_not n30110_not ; n30111
g29856 and b[7] n30029_not ; n30112
g29857 and n30023_not n30112 ; n30113
g29858 and n30031_not n30113_not ; n30114
g29859 and n30111_not n30114 ; n30115
g29860 and n30031_not n30115_not ; n30116
g29861 and b[8] n30020_not ; n30117
g29862 and n30014_not n30117 ; n30118
g29863 and n30022_not n30118_not ; n30119
g29864 and n30116_not n30119 ; n30120
g29865 and n30022_not n30120_not ; n30121
g29866 and b[9] n30011_not ; n30122
g29867 and n30005_not n30122 ; n30123
g29868 and n30013_not n30123_not ; n30124
g29869 and n30121_not n30124 ; n30125
g29870 and n30013_not n30125_not ; n30126
g29871 and b[10] n30002_not ; n30127
g29872 and n29996_not n30127 ; n30128
g29873 and n30004_not n30128_not ; n30129
g29874 and n30126_not n30129 ; n30130
g29875 and n30004_not n30130_not ; n30131
g29876 and b[11] n29993_not ; n30132
g29877 and n29987_not n30132 ; n30133
g29878 and n29995_not n30133_not ; n30134
g29879 and n30131_not n30134 ; n30135
g29880 and n29995_not n30135_not ; n30136
g29881 and b[12] n29976_not ; n30137
g29882 and n29970_not n30137 ; n30138
g29883 and n29986_not n30138_not ; n30139
g29884 and n30136_not n30139 ; n30140
g29885 and n29986_not n30140_not ; n30141
g29886 and b[13] n29978_not ; n30142
g29887 and n29983_not n30142 ; n30143
g29888 and n29985_not n30143_not ; n30144
g29889 and n30141_not n30144 ; n30145
g29890 and n29985_not n30145_not ; n30146
g29891 and n1816 n30146_not ; n30147
g29892 and n29977_not n30147_not ; n30148
g29893 and n29995_not n30139 ; n30149
g29894 and n30135_not n30149 ; n30150
g29895 and n30136_not n30139_not ; n30151
g29896 and n30150_not n30151_not ; n30152
g29897 and n1816 n30152_not ; n30153
g29898 and n30146_not n30153 ; n30154
g29899 and n30148_not n30154_not ; n30155
g29900 and b[13]_not n30155_not ; n30156
g29901 and n29994_not n30147_not ; n30157
g29902 and n30004_not n30134 ; n30158
g29903 and n30130_not n30158 ; n30159
g29904 and n30131_not n30134_not ; n30160
g29905 and n30159_not n30160_not ; n30161
g29906 and n1816 n30161_not ; n30162
g29907 and n30146_not n30162 ; n30163
g29908 and n30157_not n30163_not ; n30164
g29909 and b[12]_not n30164_not ; n30165
g29910 and n30003_not n30147_not ; n30166
g29911 and n30013_not n30129 ; n30167
g29912 and n30125_not n30167 ; n30168
g29913 and n30126_not n30129_not ; n30169
g29914 and n30168_not n30169_not ; n30170
g29915 and n1816 n30170_not ; n30171
g29916 and n30146_not n30171 ; n30172
g29917 and n30166_not n30172_not ; n30173
g29918 and b[11]_not n30173_not ; n30174
g29919 and n30012_not n30147_not ; n30175
g29920 and n30022_not n30124 ; n30176
g29921 and n30120_not n30176 ; n30177
g29922 and n30121_not n30124_not ; n30178
g29923 and n30177_not n30178_not ; n30179
g29924 and n1816 n30179_not ; n30180
g29925 and n30146_not n30180 ; n30181
g29926 and n30175_not n30181_not ; n30182
g29927 and b[10]_not n30182_not ; n30183
g29928 and n30021_not n30147_not ; n30184
g29929 and n30031_not n30119 ; n30185
g29930 and n30115_not n30185 ; n30186
g29931 and n30116_not n30119_not ; n30187
g29932 and n30186_not n30187_not ; n30188
g29933 and n1816 n30188_not ; n30189
g29934 and n30146_not n30189 ; n30190
g29935 and n30184_not n30190_not ; n30191
g29936 and b[9]_not n30191_not ; n30192
g29937 and n30030_not n30147_not ; n30193
g29938 and n30040_not n30114 ; n30194
g29939 and n30110_not n30194 ; n30195
g29940 and n30111_not n30114_not ; n30196
g29941 and n30195_not n30196_not ; n30197
g29942 and n1816 n30197_not ; n30198
g29943 and n30146_not n30198 ; n30199
g29944 and n30193_not n30199_not ; n30200
g29945 and b[8]_not n30200_not ; n30201
g29946 and n30039_not n30147_not ; n30202
g29947 and n30049_not n30109 ; n30203
g29948 and n30105_not n30203 ; n30204
g29949 and n30106_not n30109_not ; n30205
g29950 and n30204_not n30205_not ; n30206
g29951 and n1816 n30206_not ; n30207
g29952 and n30146_not n30207 ; n30208
g29953 and n30202_not n30208_not ; n30209
g29954 and b[7]_not n30209_not ; n30210
g29955 and n30048_not n30147_not ; n30211
g29956 and n30058_not n30104 ; n30212
g29957 and n30100_not n30212 ; n30213
g29958 and n30101_not n30104_not ; n30214
g29959 and n30213_not n30214_not ; n30215
g29960 and n1816 n30215_not ; n30216
g29961 and n30146_not n30216 ; n30217
g29962 and n30211_not n30217_not ; n30218
g29963 and b[6]_not n30218_not ; n30219
g29964 and n30057_not n30147_not ; n30220
g29965 and n30067_not n30099 ; n30221
g29966 and n30095_not n30221 ; n30222
g29967 and n30096_not n30099_not ; n30223
g29968 and n30222_not n30223_not ; n30224
g29969 and n1816 n30224_not ; n30225
g29970 and n30146_not n30225 ; n30226
g29971 and n30220_not n30226_not ; n30227
g29972 and b[5]_not n30227_not ; n30228
g29973 and n30066_not n30147_not ; n30229
g29974 and n30075_not n30094 ; n30230
g29975 and n30090_not n30230 ; n30231
g29976 and n30091_not n30094_not ; n30232
g29977 and n30231_not n30232_not ; n30233
g29978 and n1816 n30233_not ; n30234
g29979 and n30146_not n30234 ; n30235
g29980 and n30229_not n30235_not ; n30236
g29981 and b[4]_not n30236_not ; n30237
g29982 and n30074_not n30147_not ; n30238
g29983 and n30085_not n30089 ; n30239
g29984 and n30084_not n30239 ; n30240
g29985 and n30086_not n30089_not ; n30241
g29986 and n30240_not n30241_not ; n30242
g29987 and n1816 n30242_not ; n30243
g29988 and n30146_not n30243 ; n30244
g29989 and n30238_not n30244_not ; n30245
g29990 and b[3]_not n30245_not ; n30246
g29991 and n30079_not n30147_not ; n30247
g29992 and n1750 n30082_not ; n30248
g29993 and n30080_not n30248 ; n30249
g29994 and n1816 n30249_not ; n30250
g29995 and n30084_not n30250 ; n30251
g29996 and n30146_not n30251 ; n30252
g29997 and n30247_not n30252_not ; n30253
g29998 and b[2]_not n30253_not ; n30254
g29999 and n1929 n30146_not ; n30255
g30000 and a[50] n30255_not ; n30256
g30001 and n1935 n30146_not ; n30257
g30002 and n30256_not n30257_not ; n30258
g30003 and b[1] n30258_not ; n30259
g30004 and b[1]_not n30257_not ; n30260
g30005 and n30256_not n30260 ; n30261
g30006 and n30259_not n30261_not ; n30262
g30007 and n1942_not n30262_not ; n30263
g30008 and b[1]_not n30258_not ; n30264
g30009 and n30263_not n30264_not ; n30265
g30010 and b[2] n30252_not ; n30266
g30011 and n30247_not n30266 ; n30267
g30012 and n30254_not n30267_not ; n30268
g30013 and n30265_not n30268 ; n30269
g30014 and n30254_not n30269_not ; n30270
g30015 and b[3] n30244_not ; n30271
g30016 and n30238_not n30271 ; n30272
g30017 and n30246_not n30272_not ; n30273
g30018 and n30270_not n30273 ; n30274
g30019 and n30246_not n30274_not ; n30275
g30020 and b[4] n30235_not ; n30276
g30021 and n30229_not n30276 ; n30277
g30022 and n30237_not n30277_not ; n30278
g30023 and n30275_not n30278 ; n30279
g30024 and n30237_not n30279_not ; n30280
g30025 and b[5] n30226_not ; n30281
g30026 and n30220_not n30281 ; n30282
g30027 and n30228_not n30282_not ; n30283
g30028 and n30280_not n30283 ; n30284
g30029 and n30228_not n30284_not ; n30285
g30030 and b[6] n30217_not ; n30286
g30031 and n30211_not n30286 ; n30287
g30032 and n30219_not n30287_not ; n30288
g30033 and n30285_not n30288 ; n30289
g30034 and n30219_not n30289_not ; n30290
g30035 and b[7] n30208_not ; n30291
g30036 and n30202_not n30291 ; n30292
g30037 and n30210_not n30292_not ; n30293
g30038 and n30290_not n30293 ; n30294
g30039 and n30210_not n30294_not ; n30295
g30040 and b[8] n30199_not ; n30296
g30041 and n30193_not n30296 ; n30297
g30042 and n30201_not n30297_not ; n30298
g30043 and n30295_not n30298 ; n30299
g30044 and n30201_not n30299_not ; n30300
g30045 and b[9] n30190_not ; n30301
g30046 and n30184_not n30301 ; n30302
g30047 and n30192_not n30302_not ; n30303
g30048 and n30300_not n30303 ; n30304
g30049 and n30192_not n30304_not ; n30305
g30050 and b[10] n30181_not ; n30306
g30051 and n30175_not n30306 ; n30307
g30052 and n30183_not n30307_not ; n30308
g30053 and n30305_not n30308 ; n30309
g30054 and n30183_not n30309_not ; n30310
g30055 and b[11] n30172_not ; n30311
g30056 and n30166_not n30311 ; n30312
g30057 and n30174_not n30312_not ; n30313
g30058 and n30310_not n30313 ; n30314
g30059 and n30174_not n30314_not ; n30315
g30060 and b[12] n30163_not ; n30316
g30061 and n30157_not n30316 ; n30317
g30062 and n30165_not n30317_not ; n30318
g30063 and n30315_not n30318 ; n30319
g30064 and n30165_not n30319_not ; n30320
g30065 and b[13] n30154_not ; n30321
g30066 and n30148_not n30321 ; n30322
g30067 and n30156_not n30322_not ; n30323
g30068 and n30320_not n30323 ; n30324
g30069 and n30156_not n30324_not ; n30325
g30070 and n29984_not n30147_not ; n30326
g30071 and n29986_not n30144 ; n30327
g30072 and n30140_not n30327 ; n30328
g30073 and n30141_not n30144_not ; n30329
g30074 and n30328_not n30329_not ; n30330
g30075 and n30147 n30330_not ; n30331
g30076 and n30326_not n30331_not ; n30332
g30077 and b[14]_not n30332_not ; n30333
g30078 and b[14] n30326_not ; n30334
g30079 and n30331_not n30334 ; n30335
g30080 and n2018 n30335_not ; n30336
g30081 and n30333_not n30336 ; n30337
g30082 and n30325_not n30337 ; n30338
g30083 and n1816 n30332_not ; n30339
g30084 and n30338_not n30339_not ; n30340
g30085 and n30165_not n30323 ; n30341
g30086 and n30319_not n30341 ; n30342
g30087 and n30320_not n30323_not ; n30343
g30088 and n30342_not n30343_not ; n30344
g30089 and n30340_not n30344_not ; n30345
g30090 and n30155_not n30339_not ; n30346
g30091 and n30338_not n30346 ; n30347
g30092 and n30345_not n30347_not ; n30348
g30093 and n30156_not n30335_not ; n30349
g30094 and n30333_not n30349 ; n30350
g30095 and n30324_not n30350 ; n30351
g30096 and n30333_not n30335_not ; n30352
g30097 and n30325_not n30352_not ; n30353
g30098 and n30351_not n30353_not ; n30354
g30099 and n30340_not n30354_not ; n30355
g30100 and n30332_not n30339_not ; n30356
g30101 and n30338_not n30356 ; n30357
g30102 and n30355_not n30357_not ; n30358
g30103 and b[15]_not n30358_not ; n30359
g30104 and b[14]_not n30348_not ; n30360
g30105 and n30174_not n30318 ; n30361
g30106 and n30314_not n30361 ; n30362
g30107 and n30315_not n30318_not ; n30363
g30108 and n30362_not n30363_not ; n30364
g30109 and n30340_not n30364_not ; n30365
g30110 and n30164_not n30339_not ; n30366
g30111 and n30338_not n30366 ; n30367
g30112 and n30365_not n30367_not ; n30368
g30113 and b[13]_not n30368_not ; n30369
g30114 and n30183_not n30313 ; n30370
g30115 and n30309_not n30370 ; n30371
g30116 and n30310_not n30313_not ; n30372
g30117 and n30371_not n30372_not ; n30373
g30118 and n30340_not n30373_not ; n30374
g30119 and n30173_not n30339_not ; n30375
g30120 and n30338_not n30375 ; n30376
g30121 and n30374_not n30376_not ; n30377
g30122 and b[12]_not n30377_not ; n30378
g30123 and n30192_not n30308 ; n30379
g30124 and n30304_not n30379 ; n30380
g30125 and n30305_not n30308_not ; n30381
g30126 and n30380_not n30381_not ; n30382
g30127 and n30340_not n30382_not ; n30383
g30128 and n30182_not n30339_not ; n30384
g30129 and n30338_not n30384 ; n30385
g30130 and n30383_not n30385_not ; n30386
g30131 and b[11]_not n30386_not ; n30387
g30132 and n30201_not n30303 ; n30388
g30133 and n30299_not n30388 ; n30389
g30134 and n30300_not n30303_not ; n30390
g30135 and n30389_not n30390_not ; n30391
g30136 and n30340_not n30391_not ; n30392
g30137 and n30191_not n30339_not ; n30393
g30138 and n30338_not n30393 ; n30394
g30139 and n30392_not n30394_not ; n30395
g30140 and b[10]_not n30395_not ; n30396
g30141 and n30210_not n30298 ; n30397
g30142 and n30294_not n30397 ; n30398
g30143 and n30295_not n30298_not ; n30399
g30144 and n30398_not n30399_not ; n30400
g30145 and n30340_not n30400_not ; n30401
g30146 and n30200_not n30339_not ; n30402
g30147 and n30338_not n30402 ; n30403
g30148 and n30401_not n30403_not ; n30404
g30149 and b[9]_not n30404_not ; n30405
g30150 and n30219_not n30293 ; n30406
g30151 and n30289_not n30406 ; n30407
g30152 and n30290_not n30293_not ; n30408
g30153 and n30407_not n30408_not ; n30409
g30154 and n30340_not n30409_not ; n30410
g30155 and n30209_not n30339_not ; n30411
g30156 and n30338_not n30411 ; n30412
g30157 and n30410_not n30412_not ; n30413
g30158 and b[8]_not n30413_not ; n30414
g30159 and n30228_not n30288 ; n30415
g30160 and n30284_not n30415 ; n30416
g30161 and n30285_not n30288_not ; n30417
g30162 and n30416_not n30417_not ; n30418
g30163 and n30340_not n30418_not ; n30419
g30164 and n30218_not n30339_not ; n30420
g30165 and n30338_not n30420 ; n30421
g30166 and n30419_not n30421_not ; n30422
g30167 and b[7]_not n30422_not ; n30423
g30168 and n30237_not n30283 ; n30424
g30169 and n30279_not n30424 ; n30425
g30170 and n30280_not n30283_not ; n30426
g30171 and n30425_not n30426_not ; n30427
g30172 and n30340_not n30427_not ; n30428
g30173 and n30227_not n30339_not ; n30429
g30174 and n30338_not n30429 ; n30430
g30175 and n30428_not n30430_not ; n30431
g30176 and b[6]_not n30431_not ; n30432
g30177 and n30246_not n30278 ; n30433
g30178 and n30274_not n30433 ; n30434
g30179 and n30275_not n30278_not ; n30435
g30180 and n30434_not n30435_not ; n30436
g30181 and n30340_not n30436_not ; n30437
g30182 and n30236_not n30339_not ; n30438
g30183 and n30338_not n30438 ; n30439
g30184 and n30437_not n30439_not ; n30440
g30185 and b[5]_not n30440_not ; n30441
g30186 and n30254_not n30273 ; n30442
g30187 and n30269_not n30442 ; n30443
g30188 and n30270_not n30273_not ; n30444
g30189 and n30443_not n30444_not ; n30445
g30190 and n30340_not n30445_not ; n30446
g30191 and n30245_not n30339_not ; n30447
g30192 and n30338_not n30447 ; n30448
g30193 and n30446_not n30448_not ; n30449
g30194 and b[4]_not n30449_not ; n30450
g30195 and n30264_not n30268 ; n30451
g30196 and n30263_not n30451 ; n30452
g30197 and n30265_not n30268_not ; n30453
g30198 and n30452_not n30453_not ; n30454
g30199 and n30340_not n30454_not ; n30455
g30200 and n30253_not n30339_not ; n30456
g30201 and n30338_not n30456 ; n30457
g30202 and n30455_not n30457_not ; n30458
g30203 and b[3]_not n30458_not ; n30459
g30204 and n1942 n30261_not ; n30460
g30205 and n30259_not n30460 ; n30461
g30206 and n30263_not n30461_not ; n30462
g30207 and n30340_not n30462 ; n30463
g30208 and n30258_not n30339_not ; n30464
g30209 and n30338_not n30464 ; n30465
g30210 and n30463_not n30465_not ; n30466
g30211 and b[2]_not n30466_not ; n30467
g30212 and b[0] n30340_not ; n30468
g30213 and a[49] n30468_not ; n30469
g30214 and n1942 n30340_not ; n30470
g30215 and n30469_not n30470_not ; n30471
g30216 and b[1] n30471_not ; n30472
g30217 and b[1]_not n30470_not ; n30473
g30218 and n30469_not n30473 ; n30474
g30219 and n30472_not n30474_not ; n30475
g30220 and n2159_not n30475_not ; n30476
g30221 and b[1]_not n30471_not ; n30477
g30222 and n30476_not n30477_not ; n30478
g30223 and b[2] n30465_not ; n30479
g30224 and n30463_not n30479 ; n30480
g30225 and n30467_not n30480_not ; n30481
g30226 and n30478_not n30481 ; n30482
g30227 and n30467_not n30482_not ; n30483
g30228 and b[3] n30457_not ; n30484
g30229 and n30455_not n30484 ; n30485
g30230 and n30459_not n30485_not ; n30486
g30231 and n30483_not n30486 ; n30487
g30232 and n30459_not n30487_not ; n30488
g30233 and b[4] n30448_not ; n30489
g30234 and n30446_not n30489 ; n30490
g30235 and n30450_not n30490_not ; n30491
g30236 and n30488_not n30491 ; n30492
g30237 and n30450_not n30492_not ; n30493
g30238 and b[5] n30439_not ; n30494
g30239 and n30437_not n30494 ; n30495
g30240 and n30441_not n30495_not ; n30496
g30241 and n30493_not n30496 ; n30497
g30242 and n30441_not n30497_not ; n30498
g30243 and b[6] n30430_not ; n30499
g30244 and n30428_not n30499 ; n30500
g30245 and n30432_not n30500_not ; n30501
g30246 and n30498_not n30501 ; n30502
g30247 and n30432_not n30502_not ; n30503
g30248 and b[7] n30421_not ; n30504
g30249 and n30419_not n30504 ; n30505
g30250 and n30423_not n30505_not ; n30506
g30251 and n30503_not n30506 ; n30507
g30252 and n30423_not n30507_not ; n30508
g30253 and b[8] n30412_not ; n30509
g30254 and n30410_not n30509 ; n30510
g30255 and n30414_not n30510_not ; n30511
g30256 and n30508_not n30511 ; n30512
g30257 and n30414_not n30512_not ; n30513
g30258 and b[9] n30403_not ; n30514
g30259 and n30401_not n30514 ; n30515
g30260 and n30405_not n30515_not ; n30516
g30261 and n30513_not n30516 ; n30517
g30262 and n30405_not n30517_not ; n30518
g30263 and b[10] n30394_not ; n30519
g30264 and n30392_not n30519 ; n30520
g30265 and n30396_not n30520_not ; n30521
g30266 and n30518_not n30521 ; n30522
g30267 and n30396_not n30522_not ; n30523
g30268 and b[11] n30385_not ; n30524
g30269 and n30383_not n30524 ; n30525
g30270 and n30387_not n30525_not ; n30526
g30271 and n30523_not n30526 ; n30527
g30272 and n30387_not n30527_not ; n30528
g30273 and b[12] n30376_not ; n30529
g30274 and n30374_not n30529 ; n30530
g30275 and n30378_not n30530_not ; n30531
g30276 and n30528_not n30531 ; n30532
g30277 and n30378_not n30532_not ; n30533
g30278 and b[13] n30367_not ; n30534
g30279 and n30365_not n30534 ; n30535
g30280 and n30369_not n30535_not ; n30536
g30281 and n30533_not n30536 ; n30537
g30282 and n30369_not n30537_not ; n30538
g30283 and b[14] n30347_not ; n30539
g30284 and n30345_not n30539 ; n30540
g30285 and n30360_not n30540_not ; n30541
g30286 and n30538_not n30541 ; n30542
g30287 and n30360_not n30542_not ; n30543
g30288 and b[15] n30357_not ; n30544
g30289 and n30355_not n30544 ; n30545
g30290 and n30359_not n30545_not ; n30546
g30291 and n30543_not n30546 ; n30547
g30292 and n30359_not n30547_not ; n30548
g30293 and n346 n30548_not ; n30549
g30294 and n30348_not n30549_not ; n30550
g30295 and n30369_not n30541 ; n30551
g30296 and n30537_not n30551 ; n30552
g30297 and n30538_not n30541_not ; n30553
g30298 and n30552_not n30553_not ; n30554
g30299 and n346 n30554_not ; n30555
g30300 and n30548_not n30555 ; n30556
g30301 and n30550_not n30556_not ; n30557
g30302 and n30358_not n30549_not ; n30558
g30303 and n30360_not n30546 ; n30559
g30304 and n30542_not n30559 ; n30560
g30305 and n30543_not n30546_not ; n30561
g30306 and n30560_not n30561_not ; n30562
g30307 and n30549 n30562_not ; n30563
g30308 and n30558_not n30563_not ; n30564
g30309 and b[16]_not n30564_not ; n30565
g30310 and b[15]_not n30557_not ; n30566
g30311 and n30368_not n30549_not ; n30567
g30312 and n30378_not n30536 ; n30568
g30313 and n30532_not n30568 ; n30569
g30314 and n30533_not n30536_not ; n30570
g30315 and n30569_not n30570_not ; n30571
g30316 and n346 n30571_not ; n30572
g30317 and n30548_not n30572 ; n30573
g30318 and n30567_not n30573_not ; n30574
g30319 and b[14]_not n30574_not ; n30575
g30320 and n30377_not n30549_not ; n30576
g30321 and n30387_not n30531 ; n30577
g30322 and n30527_not n30577 ; n30578
g30323 and n30528_not n30531_not ; n30579
g30324 and n30578_not n30579_not ; n30580
g30325 and n346 n30580_not ; n30581
g30326 and n30548_not n30581 ; n30582
g30327 and n30576_not n30582_not ; n30583
g30328 and b[13]_not n30583_not ; n30584
g30329 and n30386_not n30549_not ; n30585
g30330 and n30396_not n30526 ; n30586
g30331 and n30522_not n30586 ; n30587
g30332 and n30523_not n30526_not ; n30588
g30333 and n30587_not n30588_not ; n30589
g30334 and n346 n30589_not ; n30590
g30335 and n30548_not n30590 ; n30591
g30336 and n30585_not n30591_not ; n30592
g30337 and b[12]_not n30592_not ; n30593
g30338 and n30395_not n30549_not ; n30594
g30339 and n30405_not n30521 ; n30595
g30340 and n30517_not n30595 ; n30596
g30341 and n30518_not n30521_not ; n30597
g30342 and n30596_not n30597_not ; n30598
g30343 and n346 n30598_not ; n30599
g30344 and n30548_not n30599 ; n30600
g30345 and n30594_not n30600_not ; n30601
g30346 and b[11]_not n30601_not ; n30602
g30347 and n30404_not n30549_not ; n30603
g30348 and n30414_not n30516 ; n30604
g30349 and n30512_not n30604 ; n30605
g30350 and n30513_not n30516_not ; n30606
g30351 and n30605_not n30606_not ; n30607
g30352 and n346 n30607_not ; n30608
g30353 and n30548_not n30608 ; n30609
g30354 and n30603_not n30609_not ; n30610
g30355 and b[10]_not n30610_not ; n30611
g30356 and n30413_not n30549_not ; n30612
g30357 and n30423_not n30511 ; n30613
g30358 and n30507_not n30613 ; n30614
g30359 and n30508_not n30511_not ; n30615
g30360 and n30614_not n30615_not ; n30616
g30361 and n346 n30616_not ; n30617
g30362 and n30548_not n30617 ; n30618
g30363 and n30612_not n30618_not ; n30619
g30364 and b[9]_not n30619_not ; n30620
g30365 and n30422_not n30549_not ; n30621
g30366 and n30432_not n30506 ; n30622
g30367 and n30502_not n30622 ; n30623
g30368 and n30503_not n30506_not ; n30624
g30369 and n30623_not n30624_not ; n30625
g30370 and n346 n30625_not ; n30626
g30371 and n30548_not n30626 ; n30627
g30372 and n30621_not n30627_not ; n30628
g30373 and b[8]_not n30628_not ; n30629
g30374 and n30431_not n30549_not ; n30630
g30375 and n30441_not n30501 ; n30631
g30376 and n30497_not n30631 ; n30632
g30377 and n30498_not n30501_not ; n30633
g30378 and n30632_not n30633_not ; n30634
g30379 and n346 n30634_not ; n30635
g30380 and n30548_not n30635 ; n30636
g30381 and n30630_not n30636_not ; n30637
g30382 and b[7]_not n30637_not ; n30638
g30383 and n30440_not n30549_not ; n30639
g30384 and n30450_not n30496 ; n30640
g30385 and n30492_not n30640 ; n30641
g30386 and n30493_not n30496_not ; n30642
g30387 and n30641_not n30642_not ; n30643
g30388 and n346 n30643_not ; n30644
g30389 and n30548_not n30644 ; n30645
g30390 and n30639_not n30645_not ; n30646
g30391 and b[6]_not n30646_not ; n30647
g30392 and n30449_not n30549_not ; n30648
g30393 and n30459_not n30491 ; n30649
g30394 and n30487_not n30649 ; n30650
g30395 and n30488_not n30491_not ; n30651
g30396 and n30650_not n30651_not ; n30652
g30397 and n346 n30652_not ; n30653
g30398 and n30548_not n30653 ; n30654
g30399 and n30648_not n30654_not ; n30655
g30400 and b[5]_not n30655_not ; n30656
g30401 and n30458_not n30549_not ; n30657
g30402 and n30467_not n30486 ; n30658
g30403 and n30482_not n30658 ; n30659
g30404 and n30483_not n30486_not ; n30660
g30405 and n30659_not n30660_not ; n30661
g30406 and n346 n30661_not ; n30662
g30407 and n30548_not n30662 ; n30663
g30408 and n30657_not n30663_not ; n30664
g30409 and b[4]_not n30664_not ; n30665
g30410 and n30466_not n30549_not ; n30666
g30411 and n30477_not n30481 ; n30667
g30412 and n30476_not n30667 ; n30668
g30413 and n30478_not n30481_not ; n30669
g30414 and n30668_not n30669_not ; n30670
g30415 and n346 n30670_not ; n30671
g30416 and n30548_not n30671 ; n30672
g30417 and n30666_not n30672_not ; n30673
g30418 and b[3]_not n30673_not ; n30674
g30419 and n30471_not n30549_not ; n30675
g30420 and n2159 n30474_not ; n30676
g30421 and n30472_not n30676 ; n30677
g30422 and n346 n30677_not ; n30678
g30423 and n30476_not n30678 ; n30679
g30424 and n30548_not n30679 ; n30680
g30425 and n30675_not n30680_not ; n30681
g30426 and b[2]_not n30681_not ; n30682
g30427 and n2370 n30548_not ; n30683
g30428 and a[48] n30683_not ; n30684
g30429 and n2375 n30548_not ; n30685
g30430 and n30684_not n30685_not ; n30686
g30431 and b[1] n30686_not ; n30687
g30432 and b[1]_not n30685_not ; n30688
g30433 and n30684_not n30688 ; n30689
g30434 and n30687_not n30689_not ; n30690
g30435 and n2382_not n30690_not ; n30691
g30436 and b[1]_not n30686_not ; n30692
g30437 and n30691_not n30692_not ; n30693
g30438 and b[2] n30680_not ; n30694
g30439 and n30675_not n30694 ; n30695
g30440 and n30682_not n30695_not ; n30696
g30441 and n30693_not n30696 ; n30697
g30442 and n30682_not n30697_not ; n30698
g30443 and b[3] n30672_not ; n30699
g30444 and n30666_not n30699 ; n30700
g30445 and n30674_not n30700_not ; n30701
g30446 and n30698_not n30701 ; n30702
g30447 and n30674_not n30702_not ; n30703
g30448 and b[4] n30663_not ; n30704
g30449 and n30657_not n30704 ; n30705
g30450 and n30665_not n30705_not ; n30706
g30451 and n30703_not n30706 ; n30707
g30452 and n30665_not n30707_not ; n30708
g30453 and b[5] n30654_not ; n30709
g30454 and n30648_not n30709 ; n30710
g30455 and n30656_not n30710_not ; n30711
g30456 and n30708_not n30711 ; n30712
g30457 and n30656_not n30712_not ; n30713
g30458 and b[6] n30645_not ; n30714
g30459 and n30639_not n30714 ; n30715
g30460 and n30647_not n30715_not ; n30716
g30461 and n30713_not n30716 ; n30717
g30462 and n30647_not n30717_not ; n30718
g30463 and b[7] n30636_not ; n30719
g30464 and n30630_not n30719 ; n30720
g30465 and n30638_not n30720_not ; n30721
g30466 and n30718_not n30721 ; n30722
g30467 and n30638_not n30722_not ; n30723
g30468 and b[8] n30627_not ; n30724
g30469 and n30621_not n30724 ; n30725
g30470 and n30629_not n30725_not ; n30726
g30471 and n30723_not n30726 ; n30727
g30472 and n30629_not n30727_not ; n30728
g30473 and b[9] n30618_not ; n30729
g30474 and n30612_not n30729 ; n30730
g30475 and n30620_not n30730_not ; n30731
g30476 and n30728_not n30731 ; n30732
g30477 and n30620_not n30732_not ; n30733
g30478 and b[10] n30609_not ; n30734
g30479 and n30603_not n30734 ; n30735
g30480 and n30611_not n30735_not ; n30736
g30481 and n30733_not n30736 ; n30737
g30482 and n30611_not n30737_not ; n30738
g30483 and b[11] n30600_not ; n30739
g30484 and n30594_not n30739 ; n30740
g30485 and n30602_not n30740_not ; n30741
g30486 and n30738_not n30741 ; n30742
g30487 and n30602_not n30742_not ; n30743
g30488 and b[12] n30591_not ; n30744
g30489 and n30585_not n30744 ; n30745
g30490 and n30593_not n30745_not ; n30746
g30491 and n30743_not n30746 ; n30747
g30492 and n30593_not n30747_not ; n30748
g30493 and b[13] n30582_not ; n30749
g30494 and n30576_not n30749 ; n30750
g30495 and n30584_not n30750_not ; n30751
g30496 and n30748_not n30751 ; n30752
g30497 and n30584_not n30752_not ; n30753
g30498 and b[14] n30573_not ; n30754
g30499 and n30567_not n30754 ; n30755
g30500 and n30575_not n30755_not ; n30756
g30501 and n30753_not n30756 ; n30757
g30502 and n30575_not n30757_not ; n30758
g30503 and b[15] n30556_not ; n30759
g30504 and n30550_not n30759 ; n30760
g30505 and n30566_not n30760_not ; n30761
g30506 and n30758_not n30761 ; n30762
g30507 and n30566_not n30762_not ; n30763
g30508 and b[16] n30558_not ; n30764
g30509 and n30563_not n30764 ; n30765
g30510 and n30565_not n30765_not ; n30766
g30511 and n30763_not n30766 ; n30767
g30512 and n30565_not n30767_not ; n30768
g30513 and n475 n30768_not ; n30769
g30514 and n30557_not n30769_not ; n30770
g30515 and n30575_not n30761 ; n30771
g30516 and n30757_not n30771 ; n30772
g30517 and n30758_not n30761_not ; n30773
g30518 and n30772_not n30773_not ; n30774
g30519 and n475 n30774_not ; n30775
g30520 and n30768_not n30775 ; n30776
g30521 and n30770_not n30776_not ; n30777
g30522 and b[16]_not n30777_not ; n30778
g30523 and n30574_not n30769_not ; n30779
g30524 and n30584_not n30756 ; n30780
g30525 and n30752_not n30780 ; n30781
g30526 and n30753_not n30756_not ; n30782
g30527 and n30781_not n30782_not ; n30783
g30528 and n475 n30783_not ; n30784
g30529 and n30768_not n30784 ; n30785
g30530 and n30779_not n30785_not ; n30786
g30531 and b[15]_not n30786_not ; n30787
g30532 and n30583_not n30769_not ; n30788
g30533 and n30593_not n30751 ; n30789
g30534 and n30747_not n30789 ; n30790
g30535 and n30748_not n30751_not ; n30791
g30536 and n30790_not n30791_not ; n30792
g30537 and n475 n30792_not ; n30793
g30538 and n30768_not n30793 ; n30794
g30539 and n30788_not n30794_not ; n30795
g30540 and b[14]_not n30795_not ; n30796
g30541 and n30592_not n30769_not ; n30797
g30542 and n30602_not n30746 ; n30798
g30543 and n30742_not n30798 ; n30799
g30544 and n30743_not n30746_not ; n30800
g30545 and n30799_not n30800_not ; n30801
g30546 and n475 n30801_not ; n30802
g30547 and n30768_not n30802 ; n30803
g30548 and n30797_not n30803_not ; n30804
g30549 and b[13]_not n30804_not ; n30805
g30550 and n30601_not n30769_not ; n30806
g30551 and n30611_not n30741 ; n30807
g30552 and n30737_not n30807 ; n30808
g30553 and n30738_not n30741_not ; n30809
g30554 and n30808_not n30809_not ; n30810
g30555 and n475 n30810_not ; n30811
g30556 and n30768_not n30811 ; n30812
g30557 and n30806_not n30812_not ; n30813
g30558 and b[12]_not n30813_not ; n30814
g30559 and n30610_not n30769_not ; n30815
g30560 and n30620_not n30736 ; n30816
g30561 and n30732_not n30816 ; n30817
g30562 and n30733_not n30736_not ; n30818
g30563 and n30817_not n30818_not ; n30819
g30564 and n475 n30819_not ; n30820
g30565 and n30768_not n30820 ; n30821
g30566 and n30815_not n30821_not ; n30822
g30567 and b[11]_not n30822_not ; n30823
g30568 and n30619_not n30769_not ; n30824
g30569 and n30629_not n30731 ; n30825
g30570 and n30727_not n30825 ; n30826
g30571 and n30728_not n30731_not ; n30827
g30572 and n30826_not n30827_not ; n30828
g30573 and n475 n30828_not ; n30829
g30574 and n30768_not n30829 ; n30830
g30575 and n30824_not n30830_not ; n30831
g30576 and b[10]_not n30831_not ; n30832
g30577 and n30628_not n30769_not ; n30833
g30578 and n30638_not n30726 ; n30834
g30579 and n30722_not n30834 ; n30835
g30580 and n30723_not n30726_not ; n30836
g30581 and n30835_not n30836_not ; n30837
g30582 and n475 n30837_not ; n30838
g30583 and n30768_not n30838 ; n30839
g30584 and n30833_not n30839_not ; n30840
g30585 and b[9]_not n30840_not ; n30841
g30586 and n30637_not n30769_not ; n30842
g30587 and n30647_not n30721 ; n30843
g30588 and n30717_not n30843 ; n30844
g30589 and n30718_not n30721_not ; n30845
g30590 and n30844_not n30845_not ; n30846
g30591 and n475 n30846_not ; n30847
g30592 and n30768_not n30847 ; n30848
g30593 and n30842_not n30848_not ; n30849
g30594 and b[8]_not n30849_not ; n30850
g30595 and n30646_not n30769_not ; n30851
g30596 and n30656_not n30716 ; n30852
g30597 and n30712_not n30852 ; n30853
g30598 and n30713_not n30716_not ; n30854
g30599 and n30853_not n30854_not ; n30855
g30600 and n475 n30855_not ; n30856
g30601 and n30768_not n30856 ; n30857
g30602 and n30851_not n30857_not ; n30858
g30603 and b[7]_not n30858_not ; n30859
g30604 and n30655_not n30769_not ; n30860
g30605 and n30665_not n30711 ; n30861
g30606 and n30707_not n30861 ; n30862
g30607 and n30708_not n30711_not ; n30863
g30608 and n30862_not n30863_not ; n30864
g30609 and n475 n30864_not ; n30865
g30610 and n30768_not n30865 ; n30866
g30611 and n30860_not n30866_not ; n30867
g30612 and b[6]_not n30867_not ; n30868
g30613 and n30664_not n30769_not ; n30869
g30614 and n30674_not n30706 ; n30870
g30615 and n30702_not n30870 ; n30871
g30616 and n30703_not n30706_not ; n30872
g30617 and n30871_not n30872_not ; n30873
g30618 and n475 n30873_not ; n30874
g30619 and n30768_not n30874 ; n30875
g30620 and n30869_not n30875_not ; n30876
g30621 and b[5]_not n30876_not ; n30877
g30622 and n30673_not n30769_not ; n30878
g30623 and n30682_not n30701 ; n30879
g30624 and n30697_not n30879 ; n30880
g30625 and n30698_not n30701_not ; n30881
g30626 and n30880_not n30881_not ; n30882
g30627 and n475 n30882_not ; n30883
g30628 and n30768_not n30883 ; n30884
g30629 and n30878_not n30884_not ; n30885
g30630 and b[4]_not n30885_not ; n30886
g30631 and n30681_not n30769_not ; n30887
g30632 and n30692_not n30696 ; n30888
g30633 and n30691_not n30888 ; n30889
g30634 and n30693_not n30696_not ; n30890
g30635 and n30889_not n30890_not ; n30891
g30636 and n475 n30891_not ; n30892
g30637 and n30768_not n30892 ; n30893
g30638 and n30887_not n30893_not ; n30894
g30639 and b[3]_not n30894_not ; n30895
g30640 and n30686_not n30769_not ; n30896
g30641 and n2382 n30689_not ; n30897
g30642 and n30687_not n30897 ; n30898
g30643 and n475 n30898_not ; n30899
g30644 and n30691_not n30899 ; n30900
g30645 and n30768_not n30900 ; n30901
g30646 and n30896_not n30901_not ; n30902
g30647 and b[2]_not n30902_not ; n30903
g30648 and n2601 n30768_not ; n30904
g30649 and a[47] n30904_not ; n30905
g30650 and n2606 n30768_not ; n30906
g30651 and n30905_not n30906_not ; n30907
g30652 and b[1] n30907_not ; n30908
g30653 and b[1]_not n30906_not ; n30909
g30654 and n30905_not n30909 ; n30910
g30655 and n30908_not n30910_not ; n30911
g30656 and n2613_not n30911_not ; n30912
g30657 and b[1]_not n30907_not ; n30913
g30658 and n30912_not n30913_not ; n30914
g30659 and b[2] n30901_not ; n30915
g30660 and n30896_not n30915 ; n30916
g30661 and n30903_not n30916_not ; n30917
g30662 and n30914_not n30917 ; n30918
g30663 and n30903_not n30918_not ; n30919
g30664 and b[3] n30893_not ; n30920
g30665 and n30887_not n30920 ; n30921
g30666 and n30895_not n30921_not ; n30922
g30667 and n30919_not n30922 ; n30923
g30668 and n30895_not n30923_not ; n30924
g30669 and b[4] n30884_not ; n30925
g30670 and n30878_not n30925 ; n30926
g30671 and n30886_not n30926_not ; n30927
g30672 and n30924_not n30927 ; n30928
g30673 and n30886_not n30928_not ; n30929
g30674 and b[5] n30875_not ; n30930
g30675 and n30869_not n30930 ; n30931
g30676 and n30877_not n30931_not ; n30932
g30677 and n30929_not n30932 ; n30933
g30678 and n30877_not n30933_not ; n30934
g30679 and b[6] n30866_not ; n30935
g30680 and n30860_not n30935 ; n30936
g30681 and n30868_not n30936_not ; n30937
g30682 and n30934_not n30937 ; n30938
g30683 and n30868_not n30938_not ; n30939
g30684 and b[7] n30857_not ; n30940
g30685 and n30851_not n30940 ; n30941
g30686 and n30859_not n30941_not ; n30942
g30687 and n30939_not n30942 ; n30943
g30688 and n30859_not n30943_not ; n30944
g30689 and b[8] n30848_not ; n30945
g30690 and n30842_not n30945 ; n30946
g30691 and n30850_not n30946_not ; n30947
g30692 and n30944_not n30947 ; n30948
g30693 and n30850_not n30948_not ; n30949
g30694 and b[9] n30839_not ; n30950
g30695 and n30833_not n30950 ; n30951
g30696 and n30841_not n30951_not ; n30952
g30697 and n30949_not n30952 ; n30953
g30698 and n30841_not n30953_not ; n30954
g30699 and b[10] n30830_not ; n30955
g30700 and n30824_not n30955 ; n30956
g30701 and n30832_not n30956_not ; n30957
g30702 and n30954_not n30957 ; n30958
g30703 and n30832_not n30958_not ; n30959
g30704 and b[11] n30821_not ; n30960
g30705 and n30815_not n30960 ; n30961
g30706 and n30823_not n30961_not ; n30962
g30707 and n30959_not n30962 ; n30963
g30708 and n30823_not n30963_not ; n30964
g30709 and b[12] n30812_not ; n30965
g30710 and n30806_not n30965 ; n30966
g30711 and n30814_not n30966_not ; n30967
g30712 and n30964_not n30967 ; n30968
g30713 and n30814_not n30968_not ; n30969
g30714 and b[13] n30803_not ; n30970
g30715 and n30797_not n30970 ; n30971
g30716 and n30805_not n30971_not ; n30972
g30717 and n30969_not n30972 ; n30973
g30718 and n30805_not n30973_not ; n30974
g30719 and b[14] n30794_not ; n30975
g30720 and n30788_not n30975 ; n30976
g30721 and n30796_not n30976_not ; n30977
g30722 and n30974_not n30977 ; n30978
g30723 and n30796_not n30978_not ; n30979
g30724 and b[15] n30785_not ; n30980
g30725 and n30779_not n30980 ; n30981
g30726 and n30787_not n30981_not ; n30982
g30727 and n30979_not n30982 ; n30983
g30728 and n30787_not n30983_not ; n30984
g30729 and b[16] n30776_not ; n30985
g30730 and n30770_not n30985 ; n30986
g30731 and n30778_not n30986_not ; n30987
g30732 and n30984_not n30987 ; n30988
g30733 and n30778_not n30988_not ; n30989
g30734 and n30564_not n30769_not ; n30990
g30735 and n30566_not n30766 ; n30991
g30736 and n30762_not n30991 ; n30992
g30737 and n30763_not n30766_not ; n30993
g30738 and n30992_not n30993_not ; n30994
g30739 and n30769 n30994_not ; n30995
g30740 and n30990_not n30995_not ; n30996
g30741 and b[17]_not n30996_not ; n30997
g30742 and b[17] n30990_not ; n30998
g30743 and n30995_not n30998 ; n30999
g30744 and n2705 n30999_not ; n31000
g30745 and n30997_not n31000 ; n31001
g30746 and n30989_not n31001 ; n31002
g30747 and n475 n30996_not ; n31003
g30748 and n31002_not n31003_not ; n31004
g30749 and n30787_not n30987 ; n31005
g30750 and n30983_not n31005 ; n31006
g30751 and n30984_not n30987_not ; n31007
g30752 and n31006_not n31007_not ; n31008
g30753 and n31004_not n31008_not ; n31009
g30754 and n30777_not n31003_not ; n31010
g30755 and n31002_not n31010 ; n31011
g30756 and n31009_not n31011_not ; n31012
g30757 and n30778_not n30999_not ; n31013
g30758 and n30997_not n31013 ; n31014
g30759 and n30988_not n31014 ; n31015
g30760 and n30997_not n30999_not ; n31016
g30761 and n30989_not n31016_not ; n31017
g30762 and n31015_not n31017_not ; n31018
g30763 and n31004_not n31018_not ; n31019
g30764 and n30996_not n31003_not ; n31020
g30765 and n31002_not n31020 ; n31021
g30766 and n31019_not n31021_not ; n31022
g30767 and b[18]_not n31022_not ; n31023
g30768 and b[17]_not n31012_not ; n31024
g30769 and n30796_not n30982 ; n31025
g30770 and n30978_not n31025 ; n31026
g30771 and n30979_not n30982_not ; n31027
g30772 and n31026_not n31027_not ; n31028
g30773 and n31004_not n31028_not ; n31029
g30774 and n30786_not n31003_not ; n31030
g30775 and n31002_not n31030 ; n31031
g30776 and n31029_not n31031_not ; n31032
g30777 and b[16]_not n31032_not ; n31033
g30778 and n30805_not n30977 ; n31034
g30779 and n30973_not n31034 ; n31035
g30780 and n30974_not n30977_not ; n31036
g30781 and n31035_not n31036_not ; n31037
g30782 and n31004_not n31037_not ; n31038
g30783 and n30795_not n31003_not ; n31039
g30784 and n31002_not n31039 ; n31040
g30785 and n31038_not n31040_not ; n31041
g30786 and b[15]_not n31041_not ; n31042
g30787 and n30814_not n30972 ; n31043
g30788 and n30968_not n31043 ; n31044
g30789 and n30969_not n30972_not ; n31045
g30790 and n31044_not n31045_not ; n31046
g30791 and n31004_not n31046_not ; n31047
g30792 and n30804_not n31003_not ; n31048
g30793 and n31002_not n31048 ; n31049
g30794 and n31047_not n31049_not ; n31050
g30795 and b[14]_not n31050_not ; n31051
g30796 and n30823_not n30967 ; n31052
g30797 and n30963_not n31052 ; n31053
g30798 and n30964_not n30967_not ; n31054
g30799 and n31053_not n31054_not ; n31055
g30800 and n31004_not n31055_not ; n31056
g30801 and n30813_not n31003_not ; n31057
g30802 and n31002_not n31057 ; n31058
g30803 and n31056_not n31058_not ; n31059
g30804 and b[13]_not n31059_not ; n31060
g30805 and n30832_not n30962 ; n31061
g30806 and n30958_not n31061 ; n31062
g30807 and n30959_not n30962_not ; n31063
g30808 and n31062_not n31063_not ; n31064
g30809 and n31004_not n31064_not ; n31065
g30810 and n30822_not n31003_not ; n31066
g30811 and n31002_not n31066 ; n31067
g30812 and n31065_not n31067_not ; n31068
g30813 and b[12]_not n31068_not ; n31069
g30814 and n30841_not n30957 ; n31070
g30815 and n30953_not n31070 ; n31071
g30816 and n30954_not n30957_not ; n31072
g30817 and n31071_not n31072_not ; n31073
g30818 and n31004_not n31073_not ; n31074
g30819 and n30831_not n31003_not ; n31075
g30820 and n31002_not n31075 ; n31076
g30821 and n31074_not n31076_not ; n31077
g30822 and b[11]_not n31077_not ; n31078
g30823 and n30850_not n30952 ; n31079
g30824 and n30948_not n31079 ; n31080
g30825 and n30949_not n30952_not ; n31081
g30826 and n31080_not n31081_not ; n31082
g30827 and n31004_not n31082_not ; n31083
g30828 and n30840_not n31003_not ; n31084
g30829 and n31002_not n31084 ; n31085
g30830 and n31083_not n31085_not ; n31086
g30831 and b[10]_not n31086_not ; n31087
g30832 and n30859_not n30947 ; n31088
g30833 and n30943_not n31088 ; n31089
g30834 and n30944_not n30947_not ; n31090
g30835 and n31089_not n31090_not ; n31091
g30836 and n31004_not n31091_not ; n31092
g30837 and n30849_not n31003_not ; n31093
g30838 and n31002_not n31093 ; n31094
g30839 and n31092_not n31094_not ; n31095
g30840 and b[9]_not n31095_not ; n31096
g30841 and n30868_not n30942 ; n31097
g30842 and n30938_not n31097 ; n31098
g30843 and n30939_not n30942_not ; n31099
g30844 and n31098_not n31099_not ; n31100
g30845 and n31004_not n31100_not ; n31101
g30846 and n30858_not n31003_not ; n31102
g30847 and n31002_not n31102 ; n31103
g30848 and n31101_not n31103_not ; n31104
g30849 and b[8]_not n31104_not ; n31105
g30850 and n30877_not n30937 ; n31106
g30851 and n30933_not n31106 ; n31107
g30852 and n30934_not n30937_not ; n31108
g30853 and n31107_not n31108_not ; n31109
g30854 and n31004_not n31109_not ; n31110
g30855 and n30867_not n31003_not ; n31111
g30856 and n31002_not n31111 ; n31112
g30857 and n31110_not n31112_not ; n31113
g30858 and b[7]_not n31113_not ; n31114
g30859 and n30886_not n30932 ; n31115
g30860 and n30928_not n31115 ; n31116
g30861 and n30929_not n30932_not ; n31117
g30862 and n31116_not n31117_not ; n31118
g30863 and n31004_not n31118_not ; n31119
g30864 and n30876_not n31003_not ; n31120
g30865 and n31002_not n31120 ; n31121
g30866 and n31119_not n31121_not ; n31122
g30867 and b[6]_not n31122_not ; n31123
g30868 and n30895_not n30927 ; n31124
g30869 and n30923_not n31124 ; n31125
g30870 and n30924_not n30927_not ; n31126
g30871 and n31125_not n31126_not ; n31127
g30872 and n31004_not n31127_not ; n31128
g30873 and n30885_not n31003_not ; n31129
g30874 and n31002_not n31129 ; n31130
g30875 and n31128_not n31130_not ; n31131
g30876 and b[5]_not n31131_not ; n31132
g30877 and n30903_not n30922 ; n31133
g30878 and n30918_not n31133 ; n31134
g30879 and n30919_not n30922_not ; n31135
g30880 and n31134_not n31135_not ; n31136
g30881 and n31004_not n31136_not ; n31137
g30882 and n30894_not n31003_not ; n31138
g30883 and n31002_not n31138 ; n31139
g30884 and n31137_not n31139_not ; n31140
g30885 and b[4]_not n31140_not ; n31141
g30886 and n30913_not n30917 ; n31142
g30887 and n30912_not n31142 ; n31143
g30888 and n30914_not n30917_not ; n31144
g30889 and n31143_not n31144_not ; n31145
g30890 and n31004_not n31145_not ; n31146
g30891 and n30902_not n31003_not ; n31147
g30892 and n31002_not n31147 ; n31148
g30893 and n31146_not n31148_not ; n31149
g30894 and b[3]_not n31149_not ; n31150
g30895 and n2613 n30910_not ; n31151
g30896 and n30908_not n31151 ; n31152
g30897 and n30912_not n31152_not ; n31153
g30898 and n31004_not n31153 ; n31154
g30899 and n30907_not n31003_not ; n31155
g30900 and n31002_not n31155 ; n31156
g30901 and n31154_not n31156_not ; n31157
g30902 and b[2]_not n31157_not ; n31158
g30903 and b[0] n31004_not ; n31159
g30904 and a[46] n31159_not ; n31160
g30905 and n2613 n31004_not ; n31161
g30906 and n31160_not n31161_not ; n31162
g30907 and b[1] n31162_not ; n31163
g30908 and b[1]_not n31161_not ; n31164
g30909 and n31160_not n31164 ; n31165
g30910 and n31163_not n31165_not ; n31166
g30911 and n2873_not n31166_not ; n31167
g30912 and b[1]_not n31162_not ; n31168
g30913 and n31167_not n31168_not ; n31169
g30914 and b[2] n31156_not ; n31170
g30915 and n31154_not n31170 ; n31171
g30916 and n31158_not n31171_not ; n31172
g30917 and n31169_not n31172 ; n31173
g30918 and n31158_not n31173_not ; n31174
g30919 and b[3] n31148_not ; n31175
g30920 and n31146_not n31175 ; n31176
g30921 and n31150_not n31176_not ; n31177
g30922 and n31174_not n31177 ; n31178
g30923 and n31150_not n31178_not ; n31179
g30924 and b[4] n31139_not ; n31180
g30925 and n31137_not n31180 ; n31181
g30926 and n31141_not n31181_not ; n31182
g30927 and n31179_not n31182 ; n31183
g30928 and n31141_not n31183_not ; n31184
g30929 and b[5] n31130_not ; n31185
g30930 and n31128_not n31185 ; n31186
g30931 and n31132_not n31186_not ; n31187
g30932 and n31184_not n31187 ; n31188
g30933 and n31132_not n31188_not ; n31189
g30934 and b[6] n31121_not ; n31190
g30935 and n31119_not n31190 ; n31191
g30936 and n31123_not n31191_not ; n31192
g30937 and n31189_not n31192 ; n31193
g30938 and n31123_not n31193_not ; n31194
g30939 and b[7] n31112_not ; n31195
g30940 and n31110_not n31195 ; n31196
g30941 and n31114_not n31196_not ; n31197
g30942 and n31194_not n31197 ; n31198
g30943 and n31114_not n31198_not ; n31199
g30944 and b[8] n31103_not ; n31200
g30945 and n31101_not n31200 ; n31201
g30946 and n31105_not n31201_not ; n31202
g30947 and n31199_not n31202 ; n31203
g30948 and n31105_not n31203_not ; n31204
g30949 and b[9] n31094_not ; n31205
g30950 and n31092_not n31205 ; n31206
g30951 and n31096_not n31206_not ; n31207
g30952 and n31204_not n31207 ; n31208
g30953 and n31096_not n31208_not ; n31209
g30954 and b[10] n31085_not ; n31210
g30955 and n31083_not n31210 ; n31211
g30956 and n31087_not n31211_not ; n31212
g30957 and n31209_not n31212 ; n31213
g30958 and n31087_not n31213_not ; n31214
g30959 and b[11] n31076_not ; n31215
g30960 and n31074_not n31215 ; n31216
g30961 and n31078_not n31216_not ; n31217
g30962 and n31214_not n31217 ; n31218
g30963 and n31078_not n31218_not ; n31219
g30964 and b[12] n31067_not ; n31220
g30965 and n31065_not n31220 ; n31221
g30966 and n31069_not n31221_not ; n31222
g30967 and n31219_not n31222 ; n31223
g30968 and n31069_not n31223_not ; n31224
g30969 and b[13] n31058_not ; n31225
g30970 and n31056_not n31225 ; n31226
g30971 and n31060_not n31226_not ; n31227
g30972 and n31224_not n31227 ; n31228
g30973 and n31060_not n31228_not ; n31229
g30974 and b[14] n31049_not ; n31230
g30975 and n31047_not n31230 ; n31231
g30976 and n31051_not n31231_not ; n31232
g30977 and n31229_not n31232 ; n31233
g30978 and n31051_not n31233_not ; n31234
g30979 and b[15] n31040_not ; n31235
g30980 and n31038_not n31235 ; n31236
g30981 and n31042_not n31236_not ; n31237
g30982 and n31234_not n31237 ; n31238
g30983 and n31042_not n31238_not ; n31239
g30984 and b[16] n31031_not ; n31240
g30985 and n31029_not n31240 ; n31241
g30986 and n31033_not n31241_not ; n31242
g30987 and n31239_not n31242 ; n31243
g30988 and n31033_not n31243_not ; n31244
g30989 and b[17] n31011_not ; n31245
g30990 and n31009_not n31245 ; n31246
g30991 and n31024_not n31246_not ; n31247
g30992 and n31244_not n31247 ; n31248
g30993 and n31024_not n31248_not ; n31249
g30994 and b[18] n31021_not ; n31250
g30995 and n31019_not n31250 ; n31251
g30996 and n31023_not n31251_not ; n31252
g30997 and n31249_not n31252 ; n31253
g30998 and n31023_not n31253_not ; n31254
g30999 and n2965 n31254_not ; n31255
g31000 and n31012_not n31255_not ; n31256
g31001 and n31033_not n31247 ; n31257
g31002 and n31243_not n31257 ; n31258
g31003 and n31244_not n31247_not ; n31259
g31004 and n31258_not n31259_not ; n31260
g31005 and n2965 n31260_not ; n31261
g31006 and n31254_not n31261 ; n31262
g31007 and n31256_not n31262_not ; n31263
g31008 and n31022_not n31255_not ; n31264
g31009 and n31024_not n31252 ; n31265
g31010 and n31248_not n31265 ; n31266
g31011 and n31249_not n31252_not ; n31267
g31012 and n31266_not n31267_not ; n31268
g31013 and n31255 n31268_not ; n31269
g31014 and n31264_not n31269_not ; n31270
g31015 and b[19]_not n31270_not ; n31271
g31016 and b[18]_not n31263_not ; n31272
g31017 and n31032_not n31255_not ; n31273
g31018 and n31042_not n31242 ; n31274
g31019 and n31238_not n31274 ; n31275
g31020 and n31239_not n31242_not ; n31276
g31021 and n31275_not n31276_not ; n31277
g31022 and n2965 n31277_not ; n31278
g31023 and n31254_not n31278 ; n31279
g31024 and n31273_not n31279_not ; n31280
g31025 and b[17]_not n31280_not ; n31281
g31026 and n31041_not n31255_not ; n31282
g31027 and n31051_not n31237 ; n31283
g31028 and n31233_not n31283 ; n31284
g31029 and n31234_not n31237_not ; n31285
g31030 and n31284_not n31285_not ; n31286
g31031 and n2965 n31286_not ; n31287
g31032 and n31254_not n31287 ; n31288
g31033 and n31282_not n31288_not ; n31289
g31034 and b[16]_not n31289_not ; n31290
g31035 and n31050_not n31255_not ; n31291
g31036 and n31060_not n31232 ; n31292
g31037 and n31228_not n31292 ; n31293
g31038 and n31229_not n31232_not ; n31294
g31039 and n31293_not n31294_not ; n31295
g31040 and n2965 n31295_not ; n31296
g31041 and n31254_not n31296 ; n31297
g31042 and n31291_not n31297_not ; n31298
g31043 and b[15]_not n31298_not ; n31299
g31044 and n31059_not n31255_not ; n31300
g31045 and n31069_not n31227 ; n31301
g31046 and n31223_not n31301 ; n31302
g31047 and n31224_not n31227_not ; n31303
g31048 and n31302_not n31303_not ; n31304
g31049 and n2965 n31304_not ; n31305
g31050 and n31254_not n31305 ; n31306
g31051 and n31300_not n31306_not ; n31307
g31052 and b[14]_not n31307_not ; n31308
g31053 and n31068_not n31255_not ; n31309
g31054 and n31078_not n31222 ; n31310
g31055 and n31218_not n31310 ; n31311
g31056 and n31219_not n31222_not ; n31312
g31057 and n31311_not n31312_not ; n31313
g31058 and n2965 n31313_not ; n31314
g31059 and n31254_not n31314 ; n31315
g31060 and n31309_not n31315_not ; n31316
g31061 and b[13]_not n31316_not ; n31317
g31062 and n31077_not n31255_not ; n31318
g31063 and n31087_not n31217 ; n31319
g31064 and n31213_not n31319 ; n31320
g31065 and n31214_not n31217_not ; n31321
g31066 and n31320_not n31321_not ; n31322
g31067 and n2965 n31322_not ; n31323
g31068 and n31254_not n31323 ; n31324
g31069 and n31318_not n31324_not ; n31325
g31070 and b[12]_not n31325_not ; n31326
g31071 and n31086_not n31255_not ; n31327
g31072 and n31096_not n31212 ; n31328
g31073 and n31208_not n31328 ; n31329
g31074 and n31209_not n31212_not ; n31330
g31075 and n31329_not n31330_not ; n31331
g31076 and n2965 n31331_not ; n31332
g31077 and n31254_not n31332 ; n31333
g31078 and n31327_not n31333_not ; n31334
g31079 and b[11]_not n31334_not ; n31335
g31080 and n31095_not n31255_not ; n31336
g31081 and n31105_not n31207 ; n31337
g31082 and n31203_not n31337 ; n31338
g31083 and n31204_not n31207_not ; n31339
g31084 and n31338_not n31339_not ; n31340
g31085 and n2965 n31340_not ; n31341
g31086 and n31254_not n31341 ; n31342
g31087 and n31336_not n31342_not ; n31343
g31088 and b[10]_not n31343_not ; n31344
g31089 and n31104_not n31255_not ; n31345
g31090 and n31114_not n31202 ; n31346
g31091 and n31198_not n31346 ; n31347
g31092 and n31199_not n31202_not ; n31348
g31093 and n31347_not n31348_not ; n31349
g31094 and n2965 n31349_not ; n31350
g31095 and n31254_not n31350 ; n31351
g31096 and n31345_not n31351_not ; n31352
g31097 and b[9]_not n31352_not ; n31353
g31098 and n31113_not n31255_not ; n31354
g31099 and n31123_not n31197 ; n31355
g31100 and n31193_not n31355 ; n31356
g31101 and n31194_not n31197_not ; n31357
g31102 and n31356_not n31357_not ; n31358
g31103 and n2965 n31358_not ; n31359
g31104 and n31254_not n31359 ; n31360
g31105 and n31354_not n31360_not ; n31361
g31106 and b[8]_not n31361_not ; n31362
g31107 and n31122_not n31255_not ; n31363
g31108 and n31132_not n31192 ; n31364
g31109 and n31188_not n31364 ; n31365
g31110 and n31189_not n31192_not ; n31366
g31111 and n31365_not n31366_not ; n31367
g31112 and n2965 n31367_not ; n31368
g31113 and n31254_not n31368 ; n31369
g31114 and n31363_not n31369_not ; n31370
g31115 and b[7]_not n31370_not ; n31371
g31116 and n31131_not n31255_not ; n31372
g31117 and n31141_not n31187 ; n31373
g31118 and n31183_not n31373 ; n31374
g31119 and n31184_not n31187_not ; n31375
g31120 and n31374_not n31375_not ; n31376
g31121 and n2965 n31376_not ; n31377
g31122 and n31254_not n31377 ; n31378
g31123 and n31372_not n31378_not ; n31379
g31124 and b[6]_not n31379_not ; n31380
g31125 and n31140_not n31255_not ; n31381
g31126 and n31150_not n31182 ; n31382
g31127 and n31178_not n31382 ; n31383
g31128 and n31179_not n31182_not ; n31384
g31129 and n31383_not n31384_not ; n31385
g31130 and n2965 n31385_not ; n31386
g31131 and n31254_not n31386 ; n31387
g31132 and n31381_not n31387_not ; n31388
g31133 and b[5]_not n31388_not ; n31389
g31134 and n31149_not n31255_not ; n31390
g31135 and n31158_not n31177 ; n31391
g31136 and n31173_not n31391 ; n31392
g31137 and n31174_not n31177_not ; n31393
g31138 and n31392_not n31393_not ; n31394
g31139 and n2965 n31394_not ; n31395
g31140 and n31254_not n31395 ; n31396
g31141 and n31390_not n31396_not ; n31397
g31142 and b[4]_not n31397_not ; n31398
g31143 and n31157_not n31255_not ; n31399
g31144 and n31168_not n31172 ; n31400
g31145 and n31167_not n31400 ; n31401
g31146 and n31169_not n31172_not ; n31402
g31147 and n31401_not n31402_not ; n31403
g31148 and n2965 n31403_not ; n31404
g31149 and n31254_not n31404 ; n31405
g31150 and n31399_not n31405_not ; n31406
g31151 and b[3]_not n31406_not ; n31407
g31152 and n31162_not n31255_not ; n31408
g31153 and n2873 n31165_not ; n31409
g31154 and n31163_not n31409 ; n31410
g31155 and n2965 n31410_not ; n31411
g31156 and n31167_not n31411 ; n31412
g31157 and n31254_not n31412 ; n31413
g31158 and n31408_not n31413_not ; n31414
g31159 and b[2]_not n31414_not ; n31415
g31160 and n3131 n31254_not ; n31416
g31161 and a[45] n31416_not ; n31417
g31162 and n3138 n31254_not ; n31418
g31163 and n31417_not n31418_not ; n31419
g31164 and b[1] n31419_not ; n31420
g31165 and b[1]_not n31418_not ; n31421
g31166 and n31417_not n31421 ; n31422
g31167 and n31420_not n31422_not ; n31423
g31168 and n3145_not n31423_not ; n31424
g31169 and b[1]_not n31419_not ; n31425
g31170 and n31424_not n31425_not ; n31426
g31171 and b[2] n31413_not ; n31427
g31172 and n31408_not n31427 ; n31428
g31173 and n31415_not n31428_not ; n31429
g31174 and n31426_not n31429 ; n31430
g31175 and n31415_not n31430_not ; n31431
g31176 and b[3] n31405_not ; n31432
g31177 and n31399_not n31432 ; n31433
g31178 and n31407_not n31433_not ; n31434
g31179 and n31431_not n31434 ; n31435
g31180 and n31407_not n31435_not ; n31436
g31181 and b[4] n31396_not ; n31437
g31182 and n31390_not n31437 ; n31438
g31183 and n31398_not n31438_not ; n31439
g31184 and n31436_not n31439 ; n31440
g31185 and n31398_not n31440_not ; n31441
g31186 and b[5] n31387_not ; n31442
g31187 and n31381_not n31442 ; n31443
g31188 and n31389_not n31443_not ; n31444
g31189 and n31441_not n31444 ; n31445
g31190 and n31389_not n31445_not ; n31446
g31191 and b[6] n31378_not ; n31447
g31192 and n31372_not n31447 ; n31448
g31193 and n31380_not n31448_not ; n31449
g31194 and n31446_not n31449 ; n31450
g31195 and n31380_not n31450_not ; n31451
g31196 and b[7] n31369_not ; n31452
g31197 and n31363_not n31452 ; n31453
g31198 and n31371_not n31453_not ; n31454
g31199 and n31451_not n31454 ; n31455
g31200 and n31371_not n31455_not ; n31456
g31201 and b[8] n31360_not ; n31457
g31202 and n31354_not n31457 ; n31458
g31203 and n31362_not n31458_not ; n31459
g31204 and n31456_not n31459 ; n31460
g31205 and n31362_not n31460_not ; n31461
g31206 and b[9] n31351_not ; n31462
g31207 and n31345_not n31462 ; n31463
g31208 and n31353_not n31463_not ; n31464
g31209 and n31461_not n31464 ; n31465
g31210 and n31353_not n31465_not ; n31466
g31211 and b[10] n31342_not ; n31467
g31212 and n31336_not n31467 ; n31468
g31213 and n31344_not n31468_not ; n31469
g31214 and n31466_not n31469 ; n31470
g31215 and n31344_not n31470_not ; n31471
g31216 and b[11] n31333_not ; n31472
g31217 and n31327_not n31472 ; n31473
g31218 and n31335_not n31473_not ; n31474
g31219 and n31471_not n31474 ; n31475
g31220 and n31335_not n31475_not ; n31476
g31221 and b[12] n31324_not ; n31477
g31222 and n31318_not n31477 ; n31478
g31223 and n31326_not n31478_not ; n31479
g31224 and n31476_not n31479 ; n31480
g31225 and n31326_not n31480_not ; n31481
g31226 and b[13] n31315_not ; n31482
g31227 and n31309_not n31482 ; n31483
g31228 and n31317_not n31483_not ; n31484
g31229 and n31481_not n31484 ; n31485
g31230 and n31317_not n31485_not ; n31486
g31231 and b[14] n31306_not ; n31487
g31232 and n31300_not n31487 ; n31488
g31233 and n31308_not n31488_not ; n31489
g31234 and n31486_not n31489 ; n31490
g31235 and n31308_not n31490_not ; n31491
g31236 and b[15] n31297_not ; n31492
g31237 and n31291_not n31492 ; n31493
g31238 and n31299_not n31493_not ; n31494
g31239 and n31491_not n31494 ; n31495
g31240 and n31299_not n31495_not ; n31496
g31241 and b[16] n31288_not ; n31497
g31242 and n31282_not n31497 ; n31498
g31243 and n31290_not n31498_not ; n31499
g31244 and n31496_not n31499 ; n31500
g31245 and n31290_not n31500_not ; n31501
g31246 and b[17] n31279_not ; n31502
g31247 and n31273_not n31502 ; n31503
g31248 and n31281_not n31503_not ; n31504
g31249 and n31501_not n31504 ; n31505
g31250 and n31281_not n31505_not ; n31506
g31251 and b[18] n31262_not ; n31507
g31252 and n31256_not n31507 ; n31508
g31253 and n31272_not n31508_not ; n31509
g31254 and n31506_not n31509 ; n31510
g31255 and n31272_not n31510_not ; n31511
g31256 and b[19] n31264_not ; n31512
g31257 and n31269_not n31512 ; n31513
g31258 and n31271_not n31513_not ; n31514
g31259 and n31511_not n31514 ; n31515
g31260 and n31271_not n31515_not ; n31516
g31261 and n320 n31516_not ; n31517
g31262 and n31263_not n31517_not ; n31518
g31263 and n31281_not n31509 ; n31519
g31264 and n31505_not n31519 ; n31520
g31265 and n31506_not n31509_not ; n31521
g31266 and n31520_not n31521_not ; n31522
g31267 and n320 n31522_not ; n31523
g31268 and n31516_not n31523 ; n31524
g31269 and n31518_not n31524_not ; n31525
g31270 and b[19]_not n31525_not ; n31526
g31271 and n31280_not n31517_not ; n31527
g31272 and n31290_not n31504 ; n31528
g31273 and n31500_not n31528 ; n31529
g31274 and n31501_not n31504_not ; n31530
g31275 and n31529_not n31530_not ; n31531
g31276 and n320 n31531_not ; n31532
g31277 and n31516_not n31532 ; n31533
g31278 and n31527_not n31533_not ; n31534
g31279 and b[18]_not n31534_not ; n31535
g31280 and n31289_not n31517_not ; n31536
g31281 and n31299_not n31499 ; n31537
g31282 and n31495_not n31537 ; n31538
g31283 and n31496_not n31499_not ; n31539
g31284 and n31538_not n31539_not ; n31540
g31285 and n320 n31540_not ; n31541
g31286 and n31516_not n31541 ; n31542
g31287 and n31536_not n31542_not ; n31543
g31288 and b[17]_not n31543_not ; n31544
g31289 and n31298_not n31517_not ; n31545
g31290 and n31308_not n31494 ; n31546
g31291 and n31490_not n31546 ; n31547
g31292 and n31491_not n31494_not ; n31548
g31293 and n31547_not n31548_not ; n31549
g31294 and n320 n31549_not ; n31550
g31295 and n31516_not n31550 ; n31551
g31296 and n31545_not n31551_not ; n31552
g31297 and b[16]_not n31552_not ; n31553
g31298 and n31307_not n31517_not ; n31554
g31299 and n31317_not n31489 ; n31555
g31300 and n31485_not n31555 ; n31556
g31301 and n31486_not n31489_not ; n31557
g31302 and n31556_not n31557_not ; n31558
g31303 and n320 n31558_not ; n31559
g31304 and n31516_not n31559 ; n31560
g31305 and n31554_not n31560_not ; n31561
g31306 and b[15]_not n31561_not ; n31562
g31307 and n31316_not n31517_not ; n31563
g31308 and n31326_not n31484 ; n31564
g31309 and n31480_not n31564 ; n31565
g31310 and n31481_not n31484_not ; n31566
g31311 and n31565_not n31566_not ; n31567
g31312 and n320 n31567_not ; n31568
g31313 and n31516_not n31568 ; n31569
g31314 and n31563_not n31569_not ; n31570
g31315 and b[14]_not n31570_not ; n31571
g31316 and n31325_not n31517_not ; n31572
g31317 and n31335_not n31479 ; n31573
g31318 and n31475_not n31573 ; n31574
g31319 and n31476_not n31479_not ; n31575
g31320 and n31574_not n31575_not ; n31576
g31321 and n320 n31576_not ; n31577
g31322 and n31516_not n31577 ; n31578
g31323 and n31572_not n31578_not ; n31579
g31324 and b[13]_not n31579_not ; n31580
g31325 and n31334_not n31517_not ; n31581
g31326 and n31344_not n31474 ; n31582
g31327 and n31470_not n31582 ; n31583
g31328 and n31471_not n31474_not ; n31584
g31329 and n31583_not n31584_not ; n31585
g31330 and n320 n31585_not ; n31586
g31331 and n31516_not n31586 ; n31587
g31332 and n31581_not n31587_not ; n31588
g31333 and b[12]_not n31588_not ; n31589
g31334 and n31343_not n31517_not ; n31590
g31335 and n31353_not n31469 ; n31591
g31336 and n31465_not n31591 ; n31592
g31337 and n31466_not n31469_not ; n31593
g31338 and n31592_not n31593_not ; n31594
g31339 and n320 n31594_not ; n31595
g31340 and n31516_not n31595 ; n31596
g31341 and n31590_not n31596_not ; n31597
g31342 and b[11]_not n31597_not ; n31598
g31343 and n31352_not n31517_not ; n31599
g31344 and n31362_not n31464 ; n31600
g31345 and n31460_not n31600 ; n31601
g31346 and n31461_not n31464_not ; n31602
g31347 and n31601_not n31602_not ; n31603
g31348 and n320 n31603_not ; n31604
g31349 and n31516_not n31604 ; n31605
g31350 and n31599_not n31605_not ; n31606
g31351 and b[10]_not n31606_not ; n31607
g31352 and n31361_not n31517_not ; n31608
g31353 and n31371_not n31459 ; n31609
g31354 and n31455_not n31609 ; n31610
g31355 and n31456_not n31459_not ; n31611
g31356 and n31610_not n31611_not ; n31612
g31357 and n320 n31612_not ; n31613
g31358 and n31516_not n31613 ; n31614
g31359 and n31608_not n31614_not ; n31615
g31360 and b[9]_not n31615_not ; n31616
g31361 and n31370_not n31517_not ; n31617
g31362 and n31380_not n31454 ; n31618
g31363 and n31450_not n31618 ; n31619
g31364 and n31451_not n31454_not ; n31620
g31365 and n31619_not n31620_not ; n31621
g31366 and n320 n31621_not ; n31622
g31367 and n31516_not n31622 ; n31623
g31368 and n31617_not n31623_not ; n31624
g31369 and b[8]_not n31624_not ; n31625
g31370 and n31379_not n31517_not ; n31626
g31371 and n31389_not n31449 ; n31627
g31372 and n31445_not n31627 ; n31628
g31373 and n31446_not n31449_not ; n31629
g31374 and n31628_not n31629_not ; n31630
g31375 and n320 n31630_not ; n31631
g31376 and n31516_not n31631 ; n31632
g31377 and n31626_not n31632_not ; n31633
g31378 and b[7]_not n31633_not ; n31634
g31379 and n31388_not n31517_not ; n31635
g31380 and n31398_not n31444 ; n31636
g31381 and n31440_not n31636 ; n31637
g31382 and n31441_not n31444_not ; n31638
g31383 and n31637_not n31638_not ; n31639
g31384 and n320 n31639_not ; n31640
g31385 and n31516_not n31640 ; n31641
g31386 and n31635_not n31641_not ; n31642
g31387 and b[6]_not n31642_not ; n31643
g31388 and n31397_not n31517_not ; n31644
g31389 and n31407_not n31439 ; n31645
g31390 and n31435_not n31645 ; n31646
g31391 and n31436_not n31439_not ; n31647
g31392 and n31646_not n31647_not ; n31648
g31393 and n320 n31648_not ; n31649
g31394 and n31516_not n31649 ; n31650
g31395 and n31644_not n31650_not ; n31651
g31396 and b[5]_not n31651_not ; n31652
g31397 and n31406_not n31517_not ; n31653
g31398 and n31415_not n31434 ; n31654
g31399 and n31430_not n31654 ; n31655
g31400 and n31431_not n31434_not ; n31656
g31401 and n31655_not n31656_not ; n31657
g31402 and n320 n31657_not ; n31658
g31403 and n31516_not n31658 ; n31659
g31404 and n31653_not n31659_not ; n31660
g31405 and b[4]_not n31660_not ; n31661
g31406 and n31414_not n31517_not ; n31662
g31407 and n31425_not n31429 ; n31663
g31408 and n31424_not n31663 ; n31664
g31409 and n31426_not n31429_not ; n31665
g31410 and n31664_not n31665_not ; n31666
g31411 and n320 n31666_not ; n31667
g31412 and n31516_not n31667 ; n31668
g31413 and n31662_not n31668_not ; n31669
g31414 and b[3]_not n31669_not ; n31670
g31415 and n31419_not n31517_not ; n31671
g31416 and n3145 n31422_not ; n31672
g31417 and n31420_not n31672 ; n31673
g31418 and n320 n31673_not ; n31674
g31419 and n31424_not n31674 ; n31675
g31420 and n31516_not n31675 ; n31676
g31421 and n31671_not n31676_not ; n31677
g31422 and b[2]_not n31677_not ; n31678
g31423 and n3405 n31516_not ; n31679
g31424 and a[44] n31679_not ; n31680
g31425 and n3411 n31516_not ; n31681
g31426 and n31680_not n31681_not ; n31682
g31427 and b[1] n31682_not ; n31683
g31428 and b[1]_not n31681_not ; n31684
g31429 and n31680_not n31684 ; n31685
g31430 and n31683_not n31685_not ; n31686
g31431 and n3418_not n31686_not ; n31687
g31432 and b[1]_not n31682_not ; n31688
g31433 and n31687_not n31688_not ; n31689
g31434 and b[2] n31676_not ; n31690
g31435 and n31671_not n31690 ; n31691
g31436 and n31678_not n31691_not ; n31692
g31437 and n31689_not n31692 ; n31693
g31438 and n31678_not n31693_not ; n31694
g31439 and b[3] n31668_not ; n31695
g31440 and n31662_not n31695 ; n31696
g31441 and n31670_not n31696_not ; n31697
g31442 and n31694_not n31697 ; n31698
g31443 and n31670_not n31698_not ; n31699
g31444 and b[4] n31659_not ; n31700
g31445 and n31653_not n31700 ; n31701
g31446 and n31661_not n31701_not ; n31702
g31447 and n31699_not n31702 ; n31703
g31448 and n31661_not n31703_not ; n31704
g31449 and b[5] n31650_not ; n31705
g31450 and n31644_not n31705 ; n31706
g31451 and n31652_not n31706_not ; n31707
g31452 and n31704_not n31707 ; n31708
g31453 and n31652_not n31708_not ; n31709
g31454 and b[6] n31641_not ; n31710
g31455 and n31635_not n31710 ; n31711
g31456 and n31643_not n31711_not ; n31712
g31457 and n31709_not n31712 ; n31713
g31458 and n31643_not n31713_not ; n31714
g31459 and b[7] n31632_not ; n31715
g31460 and n31626_not n31715 ; n31716
g31461 and n31634_not n31716_not ; n31717
g31462 and n31714_not n31717 ; n31718
g31463 and n31634_not n31718_not ; n31719
g31464 and b[8] n31623_not ; n31720
g31465 and n31617_not n31720 ; n31721
g31466 and n31625_not n31721_not ; n31722
g31467 and n31719_not n31722 ; n31723
g31468 and n31625_not n31723_not ; n31724
g31469 and b[9] n31614_not ; n31725
g31470 and n31608_not n31725 ; n31726
g31471 and n31616_not n31726_not ; n31727
g31472 and n31724_not n31727 ; n31728
g31473 and n31616_not n31728_not ; n31729
g31474 and b[10] n31605_not ; n31730
g31475 and n31599_not n31730 ; n31731
g31476 and n31607_not n31731_not ; n31732
g31477 and n31729_not n31732 ; n31733
g31478 and n31607_not n31733_not ; n31734
g31479 and b[11] n31596_not ; n31735
g31480 and n31590_not n31735 ; n31736
g31481 and n31598_not n31736_not ; n31737
g31482 and n31734_not n31737 ; n31738
g31483 and n31598_not n31738_not ; n31739
g31484 and b[12] n31587_not ; n31740
g31485 and n31581_not n31740 ; n31741
g31486 and n31589_not n31741_not ; n31742
g31487 and n31739_not n31742 ; n31743
g31488 and n31589_not n31743_not ; n31744
g31489 and b[13] n31578_not ; n31745
g31490 and n31572_not n31745 ; n31746
g31491 and n31580_not n31746_not ; n31747
g31492 and n31744_not n31747 ; n31748
g31493 and n31580_not n31748_not ; n31749
g31494 and b[14] n31569_not ; n31750
g31495 and n31563_not n31750 ; n31751
g31496 and n31571_not n31751_not ; n31752
g31497 and n31749_not n31752 ; n31753
g31498 and n31571_not n31753_not ; n31754
g31499 and b[15] n31560_not ; n31755
g31500 and n31554_not n31755 ; n31756
g31501 and n31562_not n31756_not ; n31757
g31502 and n31754_not n31757 ; n31758
g31503 and n31562_not n31758_not ; n31759
g31504 and b[16] n31551_not ; n31760
g31505 and n31545_not n31760 ; n31761
g31506 and n31553_not n31761_not ; n31762
g31507 and n31759_not n31762 ; n31763
g31508 and n31553_not n31763_not ; n31764
g31509 and b[17] n31542_not ; n31765
g31510 and n31536_not n31765 ; n31766
g31511 and n31544_not n31766_not ; n31767
g31512 and n31764_not n31767 ; n31768
g31513 and n31544_not n31768_not ; n31769
g31514 and b[18] n31533_not ; n31770
g31515 and n31527_not n31770 ; n31771
g31516 and n31535_not n31771_not ; n31772
g31517 and n31769_not n31772 ; n31773
g31518 and n31535_not n31773_not ; n31774
g31519 and b[19] n31524_not ; n31775
g31520 and n31518_not n31775 ; n31776
g31521 and n31526_not n31776_not ; n31777
g31522 and n31774_not n31777 ; n31778
g31523 and n31526_not n31778_not ; n31779
g31524 and n31270_not n31517_not ; n31780
g31525 and n31272_not n31514 ; n31781
g31526 and n31510_not n31781 ; n31782
g31527 and n31511_not n31514_not ; n31783
g31528 and n31782_not n31783_not ; n31784
g31529 and n31517 n31784_not ; n31785
g31530 and n31780_not n31785_not ; n31786
g31531 and b[20]_not n31786_not ; n31787
g31532 and b[20] n31780_not ; n31788
g31533 and n31785_not n31788 ; n31789
g31534 and n643 n31789_not ; n31790
g31535 and n31787_not n31790 ; n31791
g31536 and n31779_not n31791 ; n31792
g31537 and n320 n31786_not ; n31793
g31538 and n31792_not n31793_not ; n31794
g31539 and n31535_not n31777 ; n31795
g31540 and n31773_not n31795 ; n31796
g31541 and n31774_not n31777_not ; n31797
g31542 and n31796_not n31797_not ; n31798
g31543 and n31794_not n31798_not ; n31799
g31544 and n31525_not n31793_not ; n31800
g31545 and n31792_not n31800 ; n31801
g31546 and n31799_not n31801_not ; n31802
g31547 and n31526_not n31789_not ; n31803
g31548 and n31787_not n31803 ; n31804
g31549 and n31778_not n31804 ; n31805
g31550 and n31787_not n31789_not ; n31806
g31551 and n31779_not n31806_not ; n31807
g31552 and n31805_not n31807_not ; n31808
g31553 and n31794_not n31808_not ; n31809
g31554 and n31786_not n31793_not ; n31810
g31555 and n31792_not n31810 ; n31811
g31556 and n31809_not n31811_not ; n31812
g31557 and b[21]_not n31812_not ; n31813
g31558 and b[20]_not n31802_not ; n31814
g31559 and n31544_not n31772 ; n31815
g31560 and n31768_not n31815 ; n31816
g31561 and n31769_not n31772_not ; n31817
g31562 and n31816_not n31817_not ; n31818
g31563 and n31794_not n31818_not ; n31819
g31564 and n31534_not n31793_not ; n31820
g31565 and n31792_not n31820 ; n31821
g31566 and n31819_not n31821_not ; n31822
g31567 and b[19]_not n31822_not ; n31823
g31568 and n31553_not n31767 ; n31824
g31569 and n31763_not n31824 ; n31825
g31570 and n31764_not n31767_not ; n31826
g31571 and n31825_not n31826_not ; n31827
g31572 and n31794_not n31827_not ; n31828
g31573 and n31543_not n31793_not ; n31829
g31574 and n31792_not n31829 ; n31830
g31575 and n31828_not n31830_not ; n31831
g31576 and b[18]_not n31831_not ; n31832
g31577 and n31562_not n31762 ; n31833
g31578 and n31758_not n31833 ; n31834
g31579 and n31759_not n31762_not ; n31835
g31580 and n31834_not n31835_not ; n31836
g31581 and n31794_not n31836_not ; n31837
g31582 and n31552_not n31793_not ; n31838
g31583 and n31792_not n31838 ; n31839
g31584 and n31837_not n31839_not ; n31840
g31585 and b[17]_not n31840_not ; n31841
g31586 and n31571_not n31757 ; n31842
g31587 and n31753_not n31842 ; n31843
g31588 and n31754_not n31757_not ; n31844
g31589 and n31843_not n31844_not ; n31845
g31590 and n31794_not n31845_not ; n31846
g31591 and n31561_not n31793_not ; n31847
g31592 and n31792_not n31847 ; n31848
g31593 and n31846_not n31848_not ; n31849
g31594 and b[16]_not n31849_not ; n31850
g31595 and n31580_not n31752 ; n31851
g31596 and n31748_not n31851 ; n31852
g31597 and n31749_not n31752_not ; n31853
g31598 and n31852_not n31853_not ; n31854
g31599 and n31794_not n31854_not ; n31855
g31600 and n31570_not n31793_not ; n31856
g31601 and n31792_not n31856 ; n31857
g31602 and n31855_not n31857_not ; n31858
g31603 and b[15]_not n31858_not ; n31859
g31604 and n31589_not n31747 ; n31860
g31605 and n31743_not n31860 ; n31861
g31606 and n31744_not n31747_not ; n31862
g31607 and n31861_not n31862_not ; n31863
g31608 and n31794_not n31863_not ; n31864
g31609 and n31579_not n31793_not ; n31865
g31610 and n31792_not n31865 ; n31866
g31611 and n31864_not n31866_not ; n31867
g31612 and b[14]_not n31867_not ; n31868
g31613 and n31598_not n31742 ; n31869
g31614 and n31738_not n31869 ; n31870
g31615 and n31739_not n31742_not ; n31871
g31616 and n31870_not n31871_not ; n31872
g31617 and n31794_not n31872_not ; n31873
g31618 and n31588_not n31793_not ; n31874
g31619 and n31792_not n31874 ; n31875
g31620 and n31873_not n31875_not ; n31876
g31621 and b[13]_not n31876_not ; n31877
g31622 and n31607_not n31737 ; n31878
g31623 and n31733_not n31878 ; n31879
g31624 and n31734_not n31737_not ; n31880
g31625 and n31879_not n31880_not ; n31881
g31626 and n31794_not n31881_not ; n31882
g31627 and n31597_not n31793_not ; n31883
g31628 and n31792_not n31883 ; n31884
g31629 and n31882_not n31884_not ; n31885
g31630 and b[12]_not n31885_not ; n31886
g31631 and n31616_not n31732 ; n31887
g31632 and n31728_not n31887 ; n31888
g31633 and n31729_not n31732_not ; n31889
g31634 and n31888_not n31889_not ; n31890
g31635 and n31794_not n31890_not ; n31891
g31636 and n31606_not n31793_not ; n31892
g31637 and n31792_not n31892 ; n31893
g31638 and n31891_not n31893_not ; n31894
g31639 and b[11]_not n31894_not ; n31895
g31640 and n31625_not n31727 ; n31896
g31641 and n31723_not n31896 ; n31897
g31642 and n31724_not n31727_not ; n31898
g31643 and n31897_not n31898_not ; n31899
g31644 and n31794_not n31899_not ; n31900
g31645 and n31615_not n31793_not ; n31901
g31646 and n31792_not n31901 ; n31902
g31647 and n31900_not n31902_not ; n31903
g31648 and b[10]_not n31903_not ; n31904
g31649 and n31634_not n31722 ; n31905
g31650 and n31718_not n31905 ; n31906
g31651 and n31719_not n31722_not ; n31907
g31652 and n31906_not n31907_not ; n31908
g31653 and n31794_not n31908_not ; n31909
g31654 and n31624_not n31793_not ; n31910
g31655 and n31792_not n31910 ; n31911
g31656 and n31909_not n31911_not ; n31912
g31657 and b[9]_not n31912_not ; n31913
g31658 and n31643_not n31717 ; n31914
g31659 and n31713_not n31914 ; n31915
g31660 and n31714_not n31717_not ; n31916
g31661 and n31915_not n31916_not ; n31917
g31662 and n31794_not n31917_not ; n31918
g31663 and n31633_not n31793_not ; n31919
g31664 and n31792_not n31919 ; n31920
g31665 and n31918_not n31920_not ; n31921
g31666 and b[8]_not n31921_not ; n31922
g31667 and n31652_not n31712 ; n31923
g31668 and n31708_not n31923 ; n31924
g31669 and n31709_not n31712_not ; n31925
g31670 and n31924_not n31925_not ; n31926
g31671 and n31794_not n31926_not ; n31927
g31672 and n31642_not n31793_not ; n31928
g31673 and n31792_not n31928 ; n31929
g31674 and n31927_not n31929_not ; n31930
g31675 and b[7]_not n31930_not ; n31931
g31676 and n31661_not n31707 ; n31932
g31677 and n31703_not n31932 ; n31933
g31678 and n31704_not n31707_not ; n31934
g31679 and n31933_not n31934_not ; n31935
g31680 and n31794_not n31935_not ; n31936
g31681 and n31651_not n31793_not ; n31937
g31682 and n31792_not n31937 ; n31938
g31683 and n31936_not n31938_not ; n31939
g31684 and b[6]_not n31939_not ; n31940
g31685 and n31670_not n31702 ; n31941
g31686 and n31698_not n31941 ; n31942
g31687 and n31699_not n31702_not ; n31943
g31688 and n31942_not n31943_not ; n31944
g31689 and n31794_not n31944_not ; n31945
g31690 and n31660_not n31793_not ; n31946
g31691 and n31792_not n31946 ; n31947
g31692 and n31945_not n31947_not ; n31948
g31693 and b[5]_not n31948_not ; n31949
g31694 and n31678_not n31697 ; n31950
g31695 and n31693_not n31950 ; n31951
g31696 and n31694_not n31697_not ; n31952
g31697 and n31951_not n31952_not ; n31953
g31698 and n31794_not n31953_not ; n31954
g31699 and n31669_not n31793_not ; n31955
g31700 and n31792_not n31955 ; n31956
g31701 and n31954_not n31956_not ; n31957
g31702 and b[4]_not n31957_not ; n31958
g31703 and n31688_not n31692 ; n31959
g31704 and n31687_not n31959 ; n31960
g31705 and n31689_not n31692_not ; n31961
g31706 and n31960_not n31961_not ; n31962
g31707 and n31794_not n31962_not ; n31963
g31708 and n31677_not n31793_not ; n31964
g31709 and n31792_not n31964 ; n31965
g31710 and n31963_not n31965_not ; n31966
g31711 and b[3]_not n31966_not ; n31967
g31712 and n3418 n31685_not ; n31968
g31713 and n31683_not n31968 ; n31969
g31714 and n31687_not n31969_not ; n31970
g31715 and n31794_not n31970 ; n31971
g31716 and n31682_not n31793_not ; n31972
g31717 and n31792_not n31972 ; n31973
g31718 and n31971_not n31973_not ; n31974
g31719 and b[2]_not n31974_not ; n31975
g31720 and b[0] n31794_not ; n31976
g31721 and a[43] n31976_not ; n31977
g31722 and n3418 n31794_not ; n31978
g31723 and n31977_not n31978_not ; n31979
g31724 and b[1] n31979_not ; n31980
g31725 and b[1]_not n31978_not ; n31981
g31726 and n31977_not n31981 ; n31982
g31727 and n31980_not n31982_not ; n31983
g31728 and n3716_not n31983_not ; n31984
g31729 and b[1]_not n31979_not ; n31985
g31730 and n31984_not n31985_not ; n31986
g31731 and b[2] n31973_not ; n31987
g31732 and n31971_not n31987 ; n31988
g31733 and n31975_not n31988_not ; n31989
g31734 and n31986_not n31989 ; n31990
g31735 and n31975_not n31990_not ; n31991
g31736 and b[3] n31965_not ; n31992
g31737 and n31963_not n31992 ; n31993
g31738 and n31967_not n31993_not ; n31994
g31739 and n31991_not n31994 ; n31995
g31740 and n31967_not n31995_not ; n31996
g31741 and b[4] n31956_not ; n31997
g31742 and n31954_not n31997 ; n31998
g31743 and n31958_not n31998_not ; n31999
g31744 and n31996_not n31999 ; n32000
g31745 and n31958_not n32000_not ; n32001
g31746 and b[5] n31947_not ; n32002
g31747 and n31945_not n32002 ; n32003
g31748 and n31949_not n32003_not ; n32004
g31749 and n32001_not n32004 ; n32005
g31750 and n31949_not n32005_not ; n32006
g31751 and b[6] n31938_not ; n32007
g31752 and n31936_not n32007 ; n32008
g31753 and n31940_not n32008_not ; n32009
g31754 and n32006_not n32009 ; n32010
g31755 and n31940_not n32010_not ; n32011
g31756 and b[7] n31929_not ; n32012
g31757 and n31927_not n32012 ; n32013
g31758 and n31931_not n32013_not ; n32014
g31759 and n32011_not n32014 ; n32015
g31760 and n31931_not n32015_not ; n32016
g31761 and b[8] n31920_not ; n32017
g31762 and n31918_not n32017 ; n32018
g31763 and n31922_not n32018_not ; n32019
g31764 and n32016_not n32019 ; n32020
g31765 and n31922_not n32020_not ; n32021
g31766 and b[9] n31911_not ; n32022
g31767 and n31909_not n32022 ; n32023
g31768 and n31913_not n32023_not ; n32024
g31769 and n32021_not n32024 ; n32025
g31770 and n31913_not n32025_not ; n32026
g31771 and b[10] n31902_not ; n32027
g31772 and n31900_not n32027 ; n32028
g31773 and n31904_not n32028_not ; n32029
g31774 and n32026_not n32029 ; n32030
g31775 and n31904_not n32030_not ; n32031
g31776 and b[11] n31893_not ; n32032
g31777 and n31891_not n32032 ; n32033
g31778 and n31895_not n32033_not ; n32034
g31779 and n32031_not n32034 ; n32035
g31780 and n31895_not n32035_not ; n32036
g31781 and b[12] n31884_not ; n32037
g31782 and n31882_not n32037 ; n32038
g31783 and n31886_not n32038_not ; n32039
g31784 and n32036_not n32039 ; n32040
g31785 and n31886_not n32040_not ; n32041
g31786 and b[13] n31875_not ; n32042
g31787 and n31873_not n32042 ; n32043
g31788 and n31877_not n32043_not ; n32044
g31789 and n32041_not n32044 ; n32045
g31790 and n31877_not n32045_not ; n32046
g31791 and b[14] n31866_not ; n32047
g31792 and n31864_not n32047 ; n32048
g31793 and n31868_not n32048_not ; n32049
g31794 and n32046_not n32049 ; n32050
g31795 and n31868_not n32050_not ; n32051
g31796 and b[15] n31857_not ; n32052
g31797 and n31855_not n32052 ; n32053
g31798 and n31859_not n32053_not ; n32054
g31799 and n32051_not n32054 ; n32055
g31800 and n31859_not n32055_not ; n32056
g31801 and b[16] n31848_not ; n32057
g31802 and n31846_not n32057 ; n32058
g31803 and n31850_not n32058_not ; n32059
g31804 and n32056_not n32059 ; n32060
g31805 and n31850_not n32060_not ; n32061
g31806 and b[17] n31839_not ; n32062
g31807 and n31837_not n32062 ; n32063
g31808 and n31841_not n32063_not ; n32064
g31809 and n32061_not n32064 ; n32065
g31810 and n31841_not n32065_not ; n32066
g31811 and b[18] n31830_not ; n32067
g31812 and n31828_not n32067 ; n32068
g31813 and n31832_not n32068_not ; n32069
g31814 and n32066_not n32069 ; n32070
g31815 and n31832_not n32070_not ; n32071
g31816 and b[19] n31821_not ; n32072
g31817 and n31819_not n32072 ; n32073
g31818 and n31823_not n32073_not ; n32074
g31819 and n32071_not n32074 ; n32075
g31820 and n31823_not n32075_not ; n32076
g31821 and b[20] n31801_not ; n32077
g31822 and n31799_not n32077 ; n32078
g31823 and n31814_not n32078_not ; n32079
g31824 and n32076_not n32079 ; n32080
g31825 and n31814_not n32080_not ; n32081
g31826 and b[21] n31811_not ; n32082
g31827 and n31809_not n32082 ; n32083
g31828 and n31813_not n32083_not ; n32084
g31829 and n32081_not n32084 ; n32085
g31830 and n31813_not n32085_not ; n32086
g31831 and n3823 n32086_not ; n32087
g31832 and n31802_not n32087_not ; n32088
g31833 and n31823_not n32079 ; n32089
g31834 and n32075_not n32089 ; n32090
g31835 and n32076_not n32079_not ; n32091
g31836 and n32090_not n32091_not ; n32092
g31837 and n3823 n32092_not ; n32093
g31838 and n32086_not n32093 ; n32094
g31839 and n32088_not n32094_not ; n32095
g31840 and n31812_not n32087_not ; n32096
g31841 and n31814_not n32084 ; n32097
g31842 and n32080_not n32097 ; n32098
g31843 and n32081_not n32084_not ; n32099
g31844 and n32098_not n32099_not ; n32100
g31845 and n32087 n32100_not ; n32101
g31846 and n32096_not n32101_not ; n32102
g31847 and b[22]_not n32102_not ; n32103
g31848 and b[21]_not n32095_not ; n32104
g31849 and n31822_not n32087_not ; n32105
g31850 and n31832_not n32074 ; n32106
g31851 and n32070_not n32106 ; n32107
g31852 and n32071_not n32074_not ; n32108
g31853 and n32107_not n32108_not ; n32109
g31854 and n3823 n32109_not ; n32110
g31855 and n32086_not n32110 ; n32111
g31856 and n32105_not n32111_not ; n32112
g31857 and b[20]_not n32112_not ; n32113
g31858 and n31831_not n32087_not ; n32114
g31859 and n31841_not n32069 ; n32115
g31860 and n32065_not n32115 ; n32116
g31861 and n32066_not n32069_not ; n32117
g31862 and n32116_not n32117_not ; n32118
g31863 and n3823 n32118_not ; n32119
g31864 and n32086_not n32119 ; n32120
g31865 and n32114_not n32120_not ; n32121
g31866 and b[19]_not n32121_not ; n32122
g31867 and n31840_not n32087_not ; n32123
g31868 and n31850_not n32064 ; n32124
g31869 and n32060_not n32124 ; n32125
g31870 and n32061_not n32064_not ; n32126
g31871 and n32125_not n32126_not ; n32127
g31872 and n3823 n32127_not ; n32128
g31873 and n32086_not n32128 ; n32129
g31874 and n32123_not n32129_not ; n32130
g31875 and b[18]_not n32130_not ; n32131
g31876 and n31849_not n32087_not ; n32132
g31877 and n31859_not n32059 ; n32133
g31878 and n32055_not n32133 ; n32134
g31879 and n32056_not n32059_not ; n32135
g31880 and n32134_not n32135_not ; n32136
g31881 and n3823 n32136_not ; n32137
g31882 and n32086_not n32137 ; n32138
g31883 and n32132_not n32138_not ; n32139
g31884 and b[17]_not n32139_not ; n32140
g31885 and n31858_not n32087_not ; n32141
g31886 and n31868_not n32054 ; n32142
g31887 and n32050_not n32142 ; n32143
g31888 and n32051_not n32054_not ; n32144
g31889 and n32143_not n32144_not ; n32145
g31890 and n3823 n32145_not ; n32146
g31891 and n32086_not n32146 ; n32147
g31892 and n32141_not n32147_not ; n32148
g31893 and b[16]_not n32148_not ; n32149
g31894 and n31867_not n32087_not ; n32150
g31895 and n31877_not n32049 ; n32151
g31896 and n32045_not n32151 ; n32152
g31897 and n32046_not n32049_not ; n32153
g31898 and n32152_not n32153_not ; n32154
g31899 and n3823 n32154_not ; n32155
g31900 and n32086_not n32155 ; n32156
g31901 and n32150_not n32156_not ; n32157
g31902 and b[15]_not n32157_not ; n32158
g31903 and n31876_not n32087_not ; n32159
g31904 and n31886_not n32044 ; n32160
g31905 and n32040_not n32160 ; n32161
g31906 and n32041_not n32044_not ; n32162
g31907 and n32161_not n32162_not ; n32163
g31908 and n3823 n32163_not ; n32164
g31909 and n32086_not n32164 ; n32165
g31910 and n32159_not n32165_not ; n32166
g31911 and b[14]_not n32166_not ; n32167
g31912 and n31885_not n32087_not ; n32168
g31913 and n31895_not n32039 ; n32169
g31914 and n32035_not n32169 ; n32170
g31915 and n32036_not n32039_not ; n32171
g31916 and n32170_not n32171_not ; n32172
g31917 and n3823 n32172_not ; n32173
g31918 and n32086_not n32173 ; n32174
g31919 and n32168_not n32174_not ; n32175
g31920 and b[13]_not n32175_not ; n32176
g31921 and n31894_not n32087_not ; n32177
g31922 and n31904_not n32034 ; n32178
g31923 and n32030_not n32178 ; n32179
g31924 and n32031_not n32034_not ; n32180
g31925 and n32179_not n32180_not ; n32181
g31926 and n3823 n32181_not ; n32182
g31927 and n32086_not n32182 ; n32183
g31928 and n32177_not n32183_not ; n32184
g31929 and b[12]_not n32184_not ; n32185
g31930 and n31903_not n32087_not ; n32186
g31931 and n31913_not n32029 ; n32187
g31932 and n32025_not n32187 ; n32188
g31933 and n32026_not n32029_not ; n32189
g31934 and n32188_not n32189_not ; n32190
g31935 and n3823 n32190_not ; n32191
g31936 and n32086_not n32191 ; n32192
g31937 and n32186_not n32192_not ; n32193
g31938 and b[11]_not n32193_not ; n32194
g31939 and n31912_not n32087_not ; n32195
g31940 and n31922_not n32024 ; n32196
g31941 and n32020_not n32196 ; n32197
g31942 and n32021_not n32024_not ; n32198
g31943 and n32197_not n32198_not ; n32199
g31944 and n3823 n32199_not ; n32200
g31945 and n32086_not n32200 ; n32201
g31946 and n32195_not n32201_not ; n32202
g31947 and b[10]_not n32202_not ; n32203
g31948 and n31921_not n32087_not ; n32204
g31949 and n31931_not n32019 ; n32205
g31950 and n32015_not n32205 ; n32206
g31951 and n32016_not n32019_not ; n32207
g31952 and n32206_not n32207_not ; n32208
g31953 and n3823 n32208_not ; n32209
g31954 and n32086_not n32209 ; n32210
g31955 and n32204_not n32210_not ; n32211
g31956 and b[9]_not n32211_not ; n32212
g31957 and n31930_not n32087_not ; n32213
g31958 and n31940_not n32014 ; n32214
g31959 and n32010_not n32214 ; n32215
g31960 and n32011_not n32014_not ; n32216
g31961 and n32215_not n32216_not ; n32217
g31962 and n3823 n32217_not ; n32218
g31963 and n32086_not n32218 ; n32219
g31964 and n32213_not n32219_not ; n32220
g31965 and b[8]_not n32220_not ; n32221
g31966 and n31939_not n32087_not ; n32222
g31967 and n31949_not n32009 ; n32223
g31968 and n32005_not n32223 ; n32224
g31969 and n32006_not n32009_not ; n32225
g31970 and n32224_not n32225_not ; n32226
g31971 and n3823 n32226_not ; n32227
g31972 and n32086_not n32227 ; n32228
g31973 and n32222_not n32228_not ; n32229
g31974 and b[7]_not n32229_not ; n32230
g31975 and n31948_not n32087_not ; n32231
g31976 and n31958_not n32004 ; n32232
g31977 and n32000_not n32232 ; n32233
g31978 and n32001_not n32004_not ; n32234
g31979 and n32233_not n32234_not ; n32235
g31980 and n3823 n32235_not ; n32236
g31981 and n32086_not n32236 ; n32237
g31982 and n32231_not n32237_not ; n32238
g31983 and b[6]_not n32238_not ; n32239
g31984 and n31957_not n32087_not ; n32240
g31985 and n31967_not n31999 ; n32241
g31986 and n31995_not n32241 ; n32242
g31987 and n31996_not n31999_not ; n32243
g31988 and n32242_not n32243_not ; n32244
g31989 and n3823 n32244_not ; n32245
g31990 and n32086_not n32245 ; n32246
g31991 and n32240_not n32246_not ; n32247
g31992 and b[5]_not n32247_not ; n32248
g31993 and n31966_not n32087_not ; n32249
g31994 and n31975_not n31994 ; n32250
g31995 and n31990_not n32250 ; n32251
g31996 and n31991_not n31994_not ; n32252
g31997 and n32251_not n32252_not ; n32253
g31998 and n3823 n32253_not ; n32254
g31999 and n32086_not n32254 ; n32255
g32000 and n32249_not n32255_not ; n32256
g32001 and b[4]_not n32256_not ; n32257
g32002 and n31974_not n32087_not ; n32258
g32003 and n31985_not n31989 ; n32259
g32004 and n31984_not n32259 ; n32260
g32005 and n31986_not n31989_not ; n32261
g32006 and n32260_not n32261_not ; n32262
g32007 and n3823 n32262_not ; n32263
g32008 and n32086_not n32263 ; n32264
g32009 and n32258_not n32264_not ; n32265
g32010 and b[3]_not n32265_not ; n32266
g32011 and n31979_not n32087_not ; n32267
g32012 and n3716 n31982_not ; n32268
g32013 and n31980_not n32268 ; n32269
g32014 and n3823 n32269_not ; n32270
g32015 and n31984_not n32270 ; n32271
g32016 and n32086_not n32271 ; n32272
g32017 and n32267_not n32272_not ; n32273
g32018 and b[2]_not n32273_not ; n32274
g32019 and n4017 n32086_not ; n32275
g32020 and a[42] n32275_not ; n32276
g32021 and n4024 n32086_not ; n32277
g32022 and n32276_not n32277_not ; n32278
g32023 and b[1] n32278_not ; n32279
g32024 and b[1]_not n32277_not ; n32280
g32025 and n32276_not n32280 ; n32281
g32026 and n32279_not n32281_not ; n32282
g32027 and n4031_not n32282_not ; n32283
g32028 and b[1]_not n32278_not ; n32284
g32029 and n32283_not n32284_not ; n32285
g32030 and b[2] n32272_not ; n32286
g32031 and n32267_not n32286 ; n32287
g32032 and n32274_not n32287_not ; n32288
g32033 and n32285_not n32288 ; n32289
g32034 and n32274_not n32289_not ; n32290
g32035 and b[3] n32264_not ; n32291
g32036 and n32258_not n32291 ; n32292
g32037 and n32266_not n32292_not ; n32293
g32038 and n32290_not n32293 ; n32294
g32039 and n32266_not n32294_not ; n32295
g32040 and b[4] n32255_not ; n32296
g32041 and n32249_not n32296 ; n32297
g32042 and n32257_not n32297_not ; n32298
g32043 and n32295_not n32298 ; n32299
g32044 and n32257_not n32299_not ; n32300
g32045 and b[5] n32246_not ; n32301
g32046 and n32240_not n32301 ; n32302
g32047 and n32248_not n32302_not ; n32303
g32048 and n32300_not n32303 ; n32304
g32049 and n32248_not n32304_not ; n32305
g32050 and b[6] n32237_not ; n32306
g32051 and n32231_not n32306 ; n32307
g32052 and n32239_not n32307_not ; n32308
g32053 and n32305_not n32308 ; n32309
g32054 and n32239_not n32309_not ; n32310
g32055 and b[7] n32228_not ; n32311
g32056 and n32222_not n32311 ; n32312
g32057 and n32230_not n32312_not ; n32313
g32058 and n32310_not n32313 ; n32314
g32059 and n32230_not n32314_not ; n32315
g32060 and b[8] n32219_not ; n32316
g32061 and n32213_not n32316 ; n32317
g32062 and n32221_not n32317_not ; n32318
g32063 and n32315_not n32318 ; n32319
g32064 and n32221_not n32319_not ; n32320
g32065 and b[9] n32210_not ; n32321
g32066 and n32204_not n32321 ; n32322
g32067 and n32212_not n32322_not ; n32323
g32068 and n32320_not n32323 ; n32324
g32069 and n32212_not n32324_not ; n32325
g32070 and b[10] n32201_not ; n32326
g32071 and n32195_not n32326 ; n32327
g32072 and n32203_not n32327_not ; n32328
g32073 and n32325_not n32328 ; n32329
g32074 and n32203_not n32329_not ; n32330
g32075 and b[11] n32192_not ; n32331
g32076 and n32186_not n32331 ; n32332
g32077 and n32194_not n32332_not ; n32333
g32078 and n32330_not n32333 ; n32334
g32079 and n32194_not n32334_not ; n32335
g32080 and b[12] n32183_not ; n32336
g32081 and n32177_not n32336 ; n32337
g32082 and n32185_not n32337_not ; n32338
g32083 and n32335_not n32338 ; n32339
g32084 and n32185_not n32339_not ; n32340
g32085 and b[13] n32174_not ; n32341
g32086 and n32168_not n32341 ; n32342
g32087 and n32176_not n32342_not ; n32343
g32088 and n32340_not n32343 ; n32344
g32089 and n32176_not n32344_not ; n32345
g32090 and b[14] n32165_not ; n32346
g32091 and n32159_not n32346 ; n32347
g32092 and n32167_not n32347_not ; n32348
g32093 and n32345_not n32348 ; n32349
g32094 and n32167_not n32349_not ; n32350
g32095 and b[15] n32156_not ; n32351
g32096 and n32150_not n32351 ; n32352
g32097 and n32158_not n32352_not ; n32353
g32098 and n32350_not n32353 ; n32354
g32099 and n32158_not n32354_not ; n32355
g32100 and b[16] n32147_not ; n32356
g32101 and n32141_not n32356 ; n32357
g32102 and n32149_not n32357_not ; n32358
g32103 and n32355_not n32358 ; n32359
g32104 and n32149_not n32359_not ; n32360
g32105 and b[17] n32138_not ; n32361
g32106 and n32132_not n32361 ; n32362
g32107 and n32140_not n32362_not ; n32363
g32108 and n32360_not n32363 ; n32364
g32109 and n32140_not n32364_not ; n32365
g32110 and b[18] n32129_not ; n32366
g32111 and n32123_not n32366 ; n32367
g32112 and n32131_not n32367_not ; n32368
g32113 and n32365_not n32368 ; n32369
g32114 and n32131_not n32369_not ; n32370
g32115 and b[19] n32120_not ; n32371
g32116 and n32114_not n32371 ; n32372
g32117 and n32122_not n32372_not ; n32373
g32118 and n32370_not n32373 ; n32374
g32119 and n32122_not n32374_not ; n32375
g32120 and b[20] n32111_not ; n32376
g32121 and n32105_not n32376 ; n32377
g32122 and n32113_not n32377_not ; n32378
g32123 and n32375_not n32378 ; n32379
g32124 and n32113_not n32379_not ; n32380
g32125 and b[21] n32094_not ; n32381
g32126 and n32088_not n32381 ; n32382
g32127 and n32104_not n32382_not ; n32383
g32128 and n32380_not n32383 ; n32384
g32129 and n32104_not n32384_not ; n32385
g32130 and b[22] n32096_not ; n32386
g32131 and n32101_not n32386 ; n32387
g32132 and n32103_not n32387_not ; n32388
g32133 and n32385_not n32388 ; n32389
g32134 and n32103_not n32389_not ; n32390
g32135 and n4143 n32390_not ; n32391
g32136 and n32095_not n32391_not ; n32392
g32137 and n32113_not n32383 ; n32393
g32138 and n32379_not n32393 ; n32394
g32139 and n32380_not n32383_not ; n32395
g32140 and n32394_not n32395_not ; n32396
g32141 and n4143 n32396_not ; n32397
g32142 and n32390_not n32397 ; n32398
g32143 and n32392_not n32398_not ; n32399
g32144 and b[22]_not n32399_not ; n32400
g32145 and n32112_not n32391_not ; n32401
g32146 and n32122_not n32378 ; n32402
g32147 and n32374_not n32402 ; n32403
g32148 and n32375_not n32378_not ; n32404
g32149 and n32403_not n32404_not ; n32405
g32150 and n4143 n32405_not ; n32406
g32151 and n32390_not n32406 ; n32407
g32152 and n32401_not n32407_not ; n32408
g32153 and b[21]_not n32408_not ; n32409
g32154 and n32121_not n32391_not ; n32410
g32155 and n32131_not n32373 ; n32411
g32156 and n32369_not n32411 ; n32412
g32157 and n32370_not n32373_not ; n32413
g32158 and n32412_not n32413_not ; n32414
g32159 and n4143 n32414_not ; n32415
g32160 and n32390_not n32415 ; n32416
g32161 and n32410_not n32416_not ; n32417
g32162 and b[20]_not n32417_not ; n32418
g32163 and n32130_not n32391_not ; n32419
g32164 and n32140_not n32368 ; n32420
g32165 and n32364_not n32420 ; n32421
g32166 and n32365_not n32368_not ; n32422
g32167 and n32421_not n32422_not ; n32423
g32168 and n4143 n32423_not ; n32424
g32169 and n32390_not n32424 ; n32425
g32170 and n32419_not n32425_not ; n32426
g32171 and b[19]_not n32426_not ; n32427
g32172 and n32139_not n32391_not ; n32428
g32173 and n32149_not n32363 ; n32429
g32174 and n32359_not n32429 ; n32430
g32175 and n32360_not n32363_not ; n32431
g32176 and n32430_not n32431_not ; n32432
g32177 and n4143 n32432_not ; n32433
g32178 and n32390_not n32433 ; n32434
g32179 and n32428_not n32434_not ; n32435
g32180 and b[18]_not n32435_not ; n32436
g32181 and n32148_not n32391_not ; n32437
g32182 and n32158_not n32358 ; n32438
g32183 and n32354_not n32438 ; n32439
g32184 and n32355_not n32358_not ; n32440
g32185 and n32439_not n32440_not ; n32441
g32186 and n4143 n32441_not ; n32442
g32187 and n32390_not n32442 ; n32443
g32188 and n32437_not n32443_not ; n32444
g32189 and b[17]_not n32444_not ; n32445
g32190 and n32157_not n32391_not ; n32446
g32191 and n32167_not n32353 ; n32447
g32192 and n32349_not n32447 ; n32448
g32193 and n32350_not n32353_not ; n32449
g32194 and n32448_not n32449_not ; n32450
g32195 and n4143 n32450_not ; n32451
g32196 and n32390_not n32451 ; n32452
g32197 and n32446_not n32452_not ; n32453
g32198 and b[16]_not n32453_not ; n32454
g32199 and n32166_not n32391_not ; n32455
g32200 and n32176_not n32348 ; n32456
g32201 and n32344_not n32456 ; n32457
g32202 and n32345_not n32348_not ; n32458
g32203 and n32457_not n32458_not ; n32459
g32204 and n4143 n32459_not ; n32460
g32205 and n32390_not n32460 ; n32461
g32206 and n32455_not n32461_not ; n32462
g32207 and b[15]_not n32462_not ; n32463
g32208 and n32175_not n32391_not ; n32464
g32209 and n32185_not n32343 ; n32465
g32210 and n32339_not n32465 ; n32466
g32211 and n32340_not n32343_not ; n32467
g32212 and n32466_not n32467_not ; n32468
g32213 and n4143 n32468_not ; n32469
g32214 and n32390_not n32469 ; n32470
g32215 and n32464_not n32470_not ; n32471
g32216 and b[14]_not n32471_not ; n32472
g32217 and n32184_not n32391_not ; n32473
g32218 and n32194_not n32338 ; n32474
g32219 and n32334_not n32474 ; n32475
g32220 and n32335_not n32338_not ; n32476
g32221 and n32475_not n32476_not ; n32477
g32222 and n4143 n32477_not ; n32478
g32223 and n32390_not n32478 ; n32479
g32224 and n32473_not n32479_not ; n32480
g32225 and b[13]_not n32480_not ; n32481
g32226 and n32193_not n32391_not ; n32482
g32227 and n32203_not n32333 ; n32483
g32228 and n32329_not n32483 ; n32484
g32229 and n32330_not n32333_not ; n32485
g32230 and n32484_not n32485_not ; n32486
g32231 and n4143 n32486_not ; n32487
g32232 and n32390_not n32487 ; n32488
g32233 and n32482_not n32488_not ; n32489
g32234 and b[12]_not n32489_not ; n32490
g32235 and n32202_not n32391_not ; n32491
g32236 and n32212_not n32328 ; n32492
g32237 and n32324_not n32492 ; n32493
g32238 and n32325_not n32328_not ; n32494
g32239 and n32493_not n32494_not ; n32495
g32240 and n4143 n32495_not ; n32496
g32241 and n32390_not n32496 ; n32497
g32242 and n32491_not n32497_not ; n32498
g32243 and b[11]_not n32498_not ; n32499
g32244 and n32211_not n32391_not ; n32500
g32245 and n32221_not n32323 ; n32501
g32246 and n32319_not n32501 ; n32502
g32247 and n32320_not n32323_not ; n32503
g32248 and n32502_not n32503_not ; n32504
g32249 and n4143 n32504_not ; n32505
g32250 and n32390_not n32505 ; n32506
g32251 and n32500_not n32506_not ; n32507
g32252 and b[10]_not n32507_not ; n32508
g32253 and n32220_not n32391_not ; n32509
g32254 and n32230_not n32318 ; n32510
g32255 and n32314_not n32510 ; n32511
g32256 and n32315_not n32318_not ; n32512
g32257 and n32511_not n32512_not ; n32513
g32258 and n4143 n32513_not ; n32514
g32259 and n32390_not n32514 ; n32515
g32260 and n32509_not n32515_not ; n32516
g32261 and b[9]_not n32516_not ; n32517
g32262 and n32229_not n32391_not ; n32518
g32263 and n32239_not n32313 ; n32519
g32264 and n32309_not n32519 ; n32520
g32265 and n32310_not n32313_not ; n32521
g32266 and n32520_not n32521_not ; n32522
g32267 and n4143 n32522_not ; n32523
g32268 and n32390_not n32523 ; n32524
g32269 and n32518_not n32524_not ; n32525
g32270 and b[8]_not n32525_not ; n32526
g32271 and n32238_not n32391_not ; n32527
g32272 and n32248_not n32308 ; n32528
g32273 and n32304_not n32528 ; n32529
g32274 and n32305_not n32308_not ; n32530
g32275 and n32529_not n32530_not ; n32531
g32276 and n4143 n32531_not ; n32532
g32277 and n32390_not n32532 ; n32533
g32278 and n32527_not n32533_not ; n32534
g32279 and b[7]_not n32534_not ; n32535
g32280 and n32247_not n32391_not ; n32536
g32281 and n32257_not n32303 ; n32537
g32282 and n32299_not n32537 ; n32538
g32283 and n32300_not n32303_not ; n32539
g32284 and n32538_not n32539_not ; n32540
g32285 and n4143 n32540_not ; n32541
g32286 and n32390_not n32541 ; n32542
g32287 and n32536_not n32542_not ; n32543
g32288 and b[6]_not n32543_not ; n32544
g32289 and n32256_not n32391_not ; n32545
g32290 and n32266_not n32298 ; n32546
g32291 and n32294_not n32546 ; n32547
g32292 and n32295_not n32298_not ; n32548
g32293 and n32547_not n32548_not ; n32549
g32294 and n4143 n32549_not ; n32550
g32295 and n32390_not n32550 ; n32551
g32296 and n32545_not n32551_not ; n32552
g32297 and b[5]_not n32552_not ; n32553
g32298 and n32265_not n32391_not ; n32554
g32299 and n32274_not n32293 ; n32555
g32300 and n32289_not n32555 ; n32556
g32301 and n32290_not n32293_not ; n32557
g32302 and n32556_not n32557_not ; n32558
g32303 and n4143 n32558_not ; n32559
g32304 and n32390_not n32559 ; n32560
g32305 and n32554_not n32560_not ; n32561
g32306 and b[4]_not n32561_not ; n32562
g32307 and n32273_not n32391_not ; n32563
g32308 and n32284_not n32288 ; n32564
g32309 and n32283_not n32564 ; n32565
g32310 and n32285_not n32288_not ; n32566
g32311 and n32565_not n32566_not ; n32567
g32312 and n4143 n32567_not ; n32568
g32313 and n32390_not n32568 ; n32569
g32314 and n32563_not n32569_not ; n32570
g32315 and b[3]_not n32570_not ; n32571
g32316 and n32278_not n32391_not ; n32572
g32317 and n4031 n32281_not ; n32573
g32318 and n32279_not n32573 ; n32574
g32319 and n4143 n32574_not ; n32575
g32320 and n32283_not n32575 ; n32576
g32321 and n32390_not n32576 ; n32577
g32322 and n32572_not n32577_not ; n32578
g32323 and b[2]_not n32578_not ; n32579
g32324 and n4337 n32390_not ; n32580
g32325 and a[41] n32580_not ; n32581
g32326 and n4344 n32390_not ; n32582
g32327 and n32581_not n32582_not ; n32583
g32328 and b[1] n32583_not ; n32584
g32329 and b[1]_not n32582_not ; n32585
g32330 and n32581_not n32585 ; n32586
g32331 and n32584_not n32586_not ; n32587
g32332 and n4351_not n32587_not ; n32588
g32333 and b[1]_not n32583_not ; n32589
g32334 and n32588_not n32589_not ; n32590
g32335 and b[2] n32577_not ; n32591
g32336 and n32572_not n32591 ; n32592
g32337 and n32579_not n32592_not ; n32593
g32338 and n32590_not n32593 ; n32594
g32339 and n32579_not n32594_not ; n32595
g32340 and b[3] n32569_not ; n32596
g32341 and n32563_not n32596 ; n32597
g32342 and n32571_not n32597_not ; n32598
g32343 and n32595_not n32598 ; n32599
g32344 and n32571_not n32599_not ; n32600
g32345 and b[4] n32560_not ; n32601
g32346 and n32554_not n32601 ; n32602
g32347 and n32562_not n32602_not ; n32603
g32348 and n32600_not n32603 ; n32604
g32349 and n32562_not n32604_not ; n32605
g32350 and b[5] n32551_not ; n32606
g32351 and n32545_not n32606 ; n32607
g32352 and n32553_not n32607_not ; n32608
g32353 and n32605_not n32608 ; n32609
g32354 and n32553_not n32609_not ; n32610
g32355 and b[6] n32542_not ; n32611
g32356 and n32536_not n32611 ; n32612
g32357 and n32544_not n32612_not ; n32613
g32358 and n32610_not n32613 ; n32614
g32359 and n32544_not n32614_not ; n32615
g32360 and b[7] n32533_not ; n32616
g32361 and n32527_not n32616 ; n32617
g32362 and n32535_not n32617_not ; n32618
g32363 and n32615_not n32618 ; n32619
g32364 and n32535_not n32619_not ; n32620
g32365 and b[8] n32524_not ; n32621
g32366 and n32518_not n32621 ; n32622
g32367 and n32526_not n32622_not ; n32623
g32368 and n32620_not n32623 ; n32624
g32369 and n32526_not n32624_not ; n32625
g32370 and b[9] n32515_not ; n32626
g32371 and n32509_not n32626 ; n32627
g32372 and n32517_not n32627_not ; n32628
g32373 and n32625_not n32628 ; n32629
g32374 and n32517_not n32629_not ; n32630
g32375 and b[10] n32506_not ; n32631
g32376 and n32500_not n32631 ; n32632
g32377 and n32508_not n32632_not ; n32633
g32378 and n32630_not n32633 ; n32634
g32379 and n32508_not n32634_not ; n32635
g32380 and b[11] n32497_not ; n32636
g32381 and n32491_not n32636 ; n32637
g32382 and n32499_not n32637_not ; n32638
g32383 and n32635_not n32638 ; n32639
g32384 and n32499_not n32639_not ; n32640
g32385 and b[12] n32488_not ; n32641
g32386 and n32482_not n32641 ; n32642
g32387 and n32490_not n32642_not ; n32643
g32388 and n32640_not n32643 ; n32644
g32389 and n32490_not n32644_not ; n32645
g32390 and b[13] n32479_not ; n32646
g32391 and n32473_not n32646 ; n32647
g32392 and n32481_not n32647_not ; n32648
g32393 and n32645_not n32648 ; n32649
g32394 and n32481_not n32649_not ; n32650
g32395 and b[14] n32470_not ; n32651
g32396 and n32464_not n32651 ; n32652
g32397 and n32472_not n32652_not ; n32653
g32398 and n32650_not n32653 ; n32654
g32399 and n32472_not n32654_not ; n32655
g32400 and b[15] n32461_not ; n32656
g32401 and n32455_not n32656 ; n32657
g32402 and n32463_not n32657_not ; n32658
g32403 and n32655_not n32658 ; n32659
g32404 and n32463_not n32659_not ; n32660
g32405 and b[16] n32452_not ; n32661
g32406 and n32446_not n32661 ; n32662
g32407 and n32454_not n32662_not ; n32663
g32408 and n32660_not n32663 ; n32664
g32409 and n32454_not n32664_not ; n32665
g32410 and b[17] n32443_not ; n32666
g32411 and n32437_not n32666 ; n32667
g32412 and n32445_not n32667_not ; n32668
g32413 and n32665_not n32668 ; n32669
g32414 and n32445_not n32669_not ; n32670
g32415 and b[18] n32434_not ; n32671
g32416 and n32428_not n32671 ; n32672
g32417 and n32436_not n32672_not ; n32673
g32418 and n32670_not n32673 ; n32674
g32419 and n32436_not n32674_not ; n32675
g32420 and b[19] n32425_not ; n32676
g32421 and n32419_not n32676 ; n32677
g32422 and n32427_not n32677_not ; n32678
g32423 and n32675_not n32678 ; n32679
g32424 and n32427_not n32679_not ; n32680
g32425 and b[20] n32416_not ; n32681
g32426 and n32410_not n32681 ; n32682
g32427 and n32418_not n32682_not ; n32683
g32428 and n32680_not n32683 ; n32684
g32429 and n32418_not n32684_not ; n32685
g32430 and b[21] n32407_not ; n32686
g32431 and n32401_not n32686 ; n32687
g32432 and n32409_not n32687_not ; n32688
g32433 and n32685_not n32688 ; n32689
g32434 and n32409_not n32689_not ; n32690
g32435 and b[22] n32398_not ; n32691
g32436 and n32392_not n32691 ; n32692
g32437 and n32400_not n32692_not ; n32693
g32438 and n32690_not n32693 ; n32694
g32439 and n32400_not n32694_not ; n32695
g32440 and n32102_not n32391_not ; n32696
g32441 and n32104_not n32388 ; n32697
g32442 and n32384_not n32697 ; n32698
g32443 and n32385_not n32388_not ; n32699
g32444 and n32698_not n32699_not ; n32700
g32445 and n32391 n32700_not ; n32701
g32446 and n32696_not n32701_not ; n32702
g32447 and b[23]_not n32702_not ; n32703
g32448 and b[23] n32696_not ; n32704
g32449 and n32701_not n32704 ; n32705
g32450 and n4471 n32705_not ; n32706
g32451 and n32703_not n32706 ; n32707
g32452 and n32695_not n32707 ; n32708
g32453 and n4143 n32702_not ; n32709
g32454 and n32708_not n32709_not ; n32710
g32455 and n32409_not n32693 ; n32711
g32456 and n32689_not n32711 ; n32712
g32457 and n32690_not n32693_not ; n32713
g32458 and n32712_not n32713_not ; n32714
g32459 and n32710_not n32714_not ; n32715
g32460 and n32399_not n32709_not ; n32716
g32461 and n32708_not n32716 ; n32717
g32462 and n32715_not n32717_not ; n32718
g32463 and n32400_not n32705_not ; n32719
g32464 and n32703_not n32719 ; n32720
g32465 and n32694_not n32720 ; n32721
g32466 and n32703_not n32705_not ; n32722
g32467 and n32695_not n32722_not ; n32723
g32468 and n32721_not n32723_not ; n32724
g32469 and n32710_not n32724_not ; n32725
g32470 and n32702_not n32709_not ; n32726
g32471 and n32708_not n32726 ; n32727
g32472 and n32725_not n32727_not ; n32728
g32473 and b[24]_not n32728_not ; n32729
g32474 and b[23]_not n32718_not ; n32730
g32475 and n32418_not n32688 ; n32731
g32476 and n32684_not n32731 ; n32732
g32477 and n32685_not n32688_not ; n32733
g32478 and n32732_not n32733_not ; n32734
g32479 and n32710_not n32734_not ; n32735
g32480 and n32408_not n32709_not ; n32736
g32481 and n32708_not n32736 ; n32737
g32482 and n32735_not n32737_not ; n32738
g32483 and b[22]_not n32738_not ; n32739
g32484 and n32427_not n32683 ; n32740
g32485 and n32679_not n32740 ; n32741
g32486 and n32680_not n32683_not ; n32742
g32487 and n32741_not n32742_not ; n32743
g32488 and n32710_not n32743_not ; n32744
g32489 and n32417_not n32709_not ; n32745
g32490 and n32708_not n32745 ; n32746
g32491 and n32744_not n32746_not ; n32747
g32492 and b[21]_not n32747_not ; n32748
g32493 and n32436_not n32678 ; n32749
g32494 and n32674_not n32749 ; n32750
g32495 and n32675_not n32678_not ; n32751
g32496 and n32750_not n32751_not ; n32752
g32497 and n32710_not n32752_not ; n32753
g32498 and n32426_not n32709_not ; n32754
g32499 and n32708_not n32754 ; n32755
g32500 and n32753_not n32755_not ; n32756
g32501 and b[20]_not n32756_not ; n32757
g32502 and n32445_not n32673 ; n32758
g32503 and n32669_not n32758 ; n32759
g32504 and n32670_not n32673_not ; n32760
g32505 and n32759_not n32760_not ; n32761
g32506 and n32710_not n32761_not ; n32762
g32507 and n32435_not n32709_not ; n32763
g32508 and n32708_not n32763 ; n32764
g32509 and n32762_not n32764_not ; n32765
g32510 and b[19]_not n32765_not ; n32766
g32511 and n32454_not n32668 ; n32767
g32512 and n32664_not n32767 ; n32768
g32513 and n32665_not n32668_not ; n32769
g32514 and n32768_not n32769_not ; n32770
g32515 and n32710_not n32770_not ; n32771
g32516 and n32444_not n32709_not ; n32772
g32517 and n32708_not n32772 ; n32773
g32518 and n32771_not n32773_not ; n32774
g32519 and b[18]_not n32774_not ; n32775
g32520 and n32463_not n32663 ; n32776
g32521 and n32659_not n32776 ; n32777
g32522 and n32660_not n32663_not ; n32778
g32523 and n32777_not n32778_not ; n32779
g32524 and n32710_not n32779_not ; n32780
g32525 and n32453_not n32709_not ; n32781
g32526 and n32708_not n32781 ; n32782
g32527 and n32780_not n32782_not ; n32783
g32528 and b[17]_not n32783_not ; n32784
g32529 and n32472_not n32658 ; n32785
g32530 and n32654_not n32785 ; n32786
g32531 and n32655_not n32658_not ; n32787
g32532 and n32786_not n32787_not ; n32788
g32533 and n32710_not n32788_not ; n32789
g32534 and n32462_not n32709_not ; n32790
g32535 and n32708_not n32790 ; n32791
g32536 and n32789_not n32791_not ; n32792
g32537 and b[16]_not n32792_not ; n32793
g32538 and n32481_not n32653 ; n32794
g32539 and n32649_not n32794 ; n32795
g32540 and n32650_not n32653_not ; n32796
g32541 and n32795_not n32796_not ; n32797
g32542 and n32710_not n32797_not ; n32798
g32543 and n32471_not n32709_not ; n32799
g32544 and n32708_not n32799 ; n32800
g32545 and n32798_not n32800_not ; n32801
g32546 and b[15]_not n32801_not ; n32802
g32547 and n32490_not n32648 ; n32803
g32548 and n32644_not n32803 ; n32804
g32549 and n32645_not n32648_not ; n32805
g32550 and n32804_not n32805_not ; n32806
g32551 and n32710_not n32806_not ; n32807
g32552 and n32480_not n32709_not ; n32808
g32553 and n32708_not n32808 ; n32809
g32554 and n32807_not n32809_not ; n32810
g32555 and b[14]_not n32810_not ; n32811
g32556 and n32499_not n32643 ; n32812
g32557 and n32639_not n32812 ; n32813
g32558 and n32640_not n32643_not ; n32814
g32559 and n32813_not n32814_not ; n32815
g32560 and n32710_not n32815_not ; n32816
g32561 and n32489_not n32709_not ; n32817
g32562 and n32708_not n32817 ; n32818
g32563 and n32816_not n32818_not ; n32819
g32564 and b[13]_not n32819_not ; n32820
g32565 and n32508_not n32638 ; n32821
g32566 and n32634_not n32821 ; n32822
g32567 and n32635_not n32638_not ; n32823
g32568 and n32822_not n32823_not ; n32824
g32569 and n32710_not n32824_not ; n32825
g32570 and n32498_not n32709_not ; n32826
g32571 and n32708_not n32826 ; n32827
g32572 and n32825_not n32827_not ; n32828
g32573 and b[12]_not n32828_not ; n32829
g32574 and n32517_not n32633 ; n32830
g32575 and n32629_not n32830 ; n32831
g32576 and n32630_not n32633_not ; n32832
g32577 and n32831_not n32832_not ; n32833
g32578 and n32710_not n32833_not ; n32834
g32579 and n32507_not n32709_not ; n32835
g32580 and n32708_not n32835 ; n32836
g32581 and n32834_not n32836_not ; n32837
g32582 and b[11]_not n32837_not ; n32838
g32583 and n32526_not n32628 ; n32839
g32584 and n32624_not n32839 ; n32840
g32585 and n32625_not n32628_not ; n32841
g32586 and n32840_not n32841_not ; n32842
g32587 and n32710_not n32842_not ; n32843
g32588 and n32516_not n32709_not ; n32844
g32589 and n32708_not n32844 ; n32845
g32590 and n32843_not n32845_not ; n32846
g32591 and b[10]_not n32846_not ; n32847
g32592 and n32535_not n32623 ; n32848
g32593 and n32619_not n32848 ; n32849
g32594 and n32620_not n32623_not ; n32850
g32595 and n32849_not n32850_not ; n32851
g32596 and n32710_not n32851_not ; n32852
g32597 and n32525_not n32709_not ; n32853
g32598 and n32708_not n32853 ; n32854
g32599 and n32852_not n32854_not ; n32855
g32600 and b[9]_not n32855_not ; n32856
g32601 and n32544_not n32618 ; n32857
g32602 and n32614_not n32857 ; n32858
g32603 and n32615_not n32618_not ; n32859
g32604 and n32858_not n32859_not ; n32860
g32605 and n32710_not n32860_not ; n32861
g32606 and n32534_not n32709_not ; n32862
g32607 and n32708_not n32862 ; n32863
g32608 and n32861_not n32863_not ; n32864
g32609 and b[8]_not n32864_not ; n32865
g32610 and n32553_not n32613 ; n32866
g32611 and n32609_not n32866 ; n32867
g32612 and n32610_not n32613_not ; n32868
g32613 and n32867_not n32868_not ; n32869
g32614 and n32710_not n32869_not ; n32870
g32615 and n32543_not n32709_not ; n32871
g32616 and n32708_not n32871 ; n32872
g32617 and n32870_not n32872_not ; n32873
g32618 and b[7]_not n32873_not ; n32874
g32619 and n32562_not n32608 ; n32875
g32620 and n32604_not n32875 ; n32876
g32621 and n32605_not n32608_not ; n32877
g32622 and n32876_not n32877_not ; n32878
g32623 and n32710_not n32878_not ; n32879
g32624 and n32552_not n32709_not ; n32880
g32625 and n32708_not n32880 ; n32881
g32626 and n32879_not n32881_not ; n32882
g32627 and b[6]_not n32882_not ; n32883
g32628 and n32571_not n32603 ; n32884
g32629 and n32599_not n32884 ; n32885
g32630 and n32600_not n32603_not ; n32886
g32631 and n32885_not n32886_not ; n32887
g32632 and n32710_not n32887_not ; n32888
g32633 and n32561_not n32709_not ; n32889
g32634 and n32708_not n32889 ; n32890
g32635 and n32888_not n32890_not ; n32891
g32636 and b[5]_not n32891_not ; n32892
g32637 and n32579_not n32598 ; n32893
g32638 and n32594_not n32893 ; n32894
g32639 and n32595_not n32598_not ; n32895
g32640 and n32894_not n32895_not ; n32896
g32641 and n32710_not n32896_not ; n32897
g32642 and n32570_not n32709_not ; n32898
g32643 and n32708_not n32898 ; n32899
g32644 and n32897_not n32899_not ; n32900
g32645 and b[4]_not n32900_not ; n32901
g32646 and n32589_not n32593 ; n32902
g32647 and n32588_not n32902 ; n32903
g32648 and n32590_not n32593_not ; n32904
g32649 and n32903_not n32904_not ; n32905
g32650 and n32710_not n32905_not ; n32906
g32651 and n32578_not n32709_not ; n32907
g32652 and n32708_not n32907 ; n32908
g32653 and n32906_not n32908_not ; n32909
g32654 and b[3]_not n32909_not ; n32910
g32655 and n4351 n32586_not ; n32911
g32656 and n32584_not n32911 ; n32912
g32657 and n32588_not n32912_not ; n32913
g32658 and n32710_not n32913 ; n32914
g32659 and n32583_not n32709_not ; n32915
g32660 and n32708_not n32915 ; n32916
g32661 and n32914_not n32916_not ; n32917
g32662 and b[2]_not n32917_not ; n32918
g32663 and b[0] n32710_not ; n32919
g32664 and a[40] n32919_not ; n32920
g32665 and n4351 n32710_not ; n32921
g32666 and n32920_not n32921_not ; n32922
g32667 and b[1] n32922_not ; n32923
g32668 and b[1]_not n32921_not ; n32924
g32669 and n32920_not n32924 ; n32925
g32670 and n32923_not n32925_not ; n32926
g32671 and n4693_not n32926_not ; n32927
g32672 and b[1]_not n32922_not ; n32928
g32673 and n32927_not n32928_not ; n32929
g32674 and b[2] n32916_not ; n32930
g32675 and n32914_not n32930 ; n32931
g32676 and n32918_not n32931_not ; n32932
g32677 and n32929_not n32932 ; n32933
g32678 and n32918_not n32933_not ; n32934
g32679 and b[3] n32908_not ; n32935
g32680 and n32906_not n32935 ; n32936
g32681 and n32910_not n32936_not ; n32937
g32682 and n32934_not n32937 ; n32938
g32683 and n32910_not n32938_not ; n32939
g32684 and b[4] n32899_not ; n32940
g32685 and n32897_not n32940 ; n32941
g32686 and n32901_not n32941_not ; n32942
g32687 and n32939_not n32942 ; n32943
g32688 and n32901_not n32943_not ; n32944
g32689 and b[5] n32890_not ; n32945
g32690 and n32888_not n32945 ; n32946
g32691 and n32892_not n32946_not ; n32947
g32692 and n32944_not n32947 ; n32948
g32693 and n32892_not n32948_not ; n32949
g32694 and b[6] n32881_not ; n32950
g32695 and n32879_not n32950 ; n32951
g32696 and n32883_not n32951_not ; n32952
g32697 and n32949_not n32952 ; n32953
g32698 and n32883_not n32953_not ; n32954
g32699 and b[7] n32872_not ; n32955
g32700 and n32870_not n32955 ; n32956
g32701 and n32874_not n32956_not ; n32957
g32702 and n32954_not n32957 ; n32958
g32703 and n32874_not n32958_not ; n32959
g32704 and b[8] n32863_not ; n32960
g32705 and n32861_not n32960 ; n32961
g32706 and n32865_not n32961_not ; n32962
g32707 and n32959_not n32962 ; n32963
g32708 and n32865_not n32963_not ; n32964
g32709 and b[9] n32854_not ; n32965
g32710 and n32852_not n32965 ; n32966
g32711 and n32856_not n32966_not ; n32967
g32712 and n32964_not n32967 ; n32968
g32713 and n32856_not n32968_not ; n32969
g32714 and b[10] n32845_not ; n32970
g32715 and n32843_not n32970 ; n32971
g32716 and n32847_not n32971_not ; n32972
g32717 and n32969_not n32972 ; n32973
g32718 and n32847_not n32973_not ; n32974
g32719 and b[11] n32836_not ; n32975
g32720 and n32834_not n32975 ; n32976
g32721 and n32838_not n32976_not ; n32977
g32722 and n32974_not n32977 ; n32978
g32723 and n32838_not n32978_not ; n32979
g32724 and b[12] n32827_not ; n32980
g32725 and n32825_not n32980 ; n32981
g32726 and n32829_not n32981_not ; n32982
g32727 and n32979_not n32982 ; n32983
g32728 and n32829_not n32983_not ; n32984
g32729 and b[13] n32818_not ; n32985
g32730 and n32816_not n32985 ; n32986
g32731 and n32820_not n32986_not ; n32987
g32732 and n32984_not n32987 ; n32988
g32733 and n32820_not n32988_not ; n32989
g32734 and b[14] n32809_not ; n32990
g32735 and n32807_not n32990 ; n32991
g32736 and n32811_not n32991_not ; n32992
g32737 and n32989_not n32992 ; n32993
g32738 and n32811_not n32993_not ; n32994
g32739 and b[15] n32800_not ; n32995
g32740 and n32798_not n32995 ; n32996
g32741 and n32802_not n32996_not ; n32997
g32742 and n32994_not n32997 ; n32998
g32743 and n32802_not n32998_not ; n32999
g32744 and b[16] n32791_not ; n33000
g32745 and n32789_not n33000 ; n33001
g32746 and n32793_not n33001_not ; n33002
g32747 and n32999_not n33002 ; n33003
g32748 and n32793_not n33003_not ; n33004
g32749 and b[17] n32782_not ; n33005
g32750 and n32780_not n33005 ; n33006
g32751 and n32784_not n33006_not ; n33007
g32752 and n33004_not n33007 ; n33008
g32753 and n32784_not n33008_not ; n33009
g32754 and b[18] n32773_not ; n33010
g32755 and n32771_not n33010 ; n33011
g32756 and n32775_not n33011_not ; n33012
g32757 and n33009_not n33012 ; n33013
g32758 and n32775_not n33013_not ; n33014
g32759 and b[19] n32764_not ; n33015
g32760 and n32762_not n33015 ; n33016
g32761 and n32766_not n33016_not ; n33017
g32762 and n33014_not n33017 ; n33018
g32763 and n32766_not n33018_not ; n33019
g32764 and b[20] n32755_not ; n33020
g32765 and n32753_not n33020 ; n33021
g32766 and n32757_not n33021_not ; n33022
g32767 and n33019_not n33022 ; n33023
g32768 and n32757_not n33023_not ; n33024
g32769 and b[21] n32746_not ; n33025
g32770 and n32744_not n33025 ; n33026
g32771 and n32748_not n33026_not ; n33027
g32772 and n33024_not n33027 ; n33028
g32773 and n32748_not n33028_not ; n33029
g32774 and b[22] n32737_not ; n33030
g32775 and n32735_not n33030 ; n33031
g32776 and n32739_not n33031_not ; n33032
g32777 and n33029_not n33032 ; n33033
g32778 and n32739_not n33033_not ; n33034
g32779 and b[23] n32717_not ; n33035
g32780 and n32715_not n33035 ; n33036
g32781 and n32730_not n33036_not ; n33037
g32782 and n33034_not n33037 ; n33038
g32783 and n32730_not n33038_not ; n33039
g32784 and b[24] n32727_not ; n33040
g32785 and n32725_not n33040 ; n33041
g32786 and n32729_not n33041_not ; n33042
g32787 and n33039_not n33042 ; n33043
g32788 and n32729_not n33043_not ; n33044
g32789 and n4813 n33044_not ; n33045
g32790 and n32718_not n33045_not ; n33046
g32791 and n32739_not n33037 ; n33047
g32792 and n33033_not n33047 ; n33048
g32793 and n33034_not n33037_not ; n33049
g32794 and n33048_not n33049_not ; n33050
g32795 and n4813 n33050_not ; n33051
g32796 and n33044_not n33051 ; n33052
g32797 and n33046_not n33052_not ; n33053
g32798 and n32728_not n33045_not ; n33054
g32799 and n32730_not n33042 ; n33055
g32800 and n33038_not n33055 ; n33056
g32801 and n33039_not n33042_not ; n33057
g32802 and n33056_not n33057_not ; n33058
g32803 and n33045 n33058_not ; n33059
g32804 and n33054_not n33059_not ; n33060
g32805 and b[25]_not n33060_not ; n33061
g32806 and b[24]_not n33053_not ; n33062
g32807 and n32738_not n33045_not ; n33063
g32808 and n32748_not n33032 ; n33064
g32809 and n33028_not n33064 ; n33065
g32810 and n33029_not n33032_not ; n33066
g32811 and n33065_not n33066_not ; n33067
g32812 and n4813 n33067_not ; n33068
g32813 and n33044_not n33068 ; n33069
g32814 and n33063_not n33069_not ; n33070
g32815 and b[23]_not n33070_not ; n33071
g32816 and n32747_not n33045_not ; n33072
g32817 and n32757_not n33027 ; n33073
g32818 and n33023_not n33073 ; n33074
g32819 and n33024_not n33027_not ; n33075
g32820 and n33074_not n33075_not ; n33076
g32821 and n4813 n33076_not ; n33077
g32822 and n33044_not n33077 ; n33078
g32823 and n33072_not n33078_not ; n33079
g32824 and b[22]_not n33079_not ; n33080
g32825 and n32756_not n33045_not ; n33081
g32826 and n32766_not n33022 ; n33082
g32827 and n33018_not n33082 ; n33083
g32828 and n33019_not n33022_not ; n33084
g32829 and n33083_not n33084_not ; n33085
g32830 and n4813 n33085_not ; n33086
g32831 and n33044_not n33086 ; n33087
g32832 and n33081_not n33087_not ; n33088
g32833 and b[21]_not n33088_not ; n33089
g32834 and n32765_not n33045_not ; n33090
g32835 and n32775_not n33017 ; n33091
g32836 and n33013_not n33091 ; n33092
g32837 and n33014_not n33017_not ; n33093
g32838 and n33092_not n33093_not ; n33094
g32839 and n4813 n33094_not ; n33095
g32840 and n33044_not n33095 ; n33096
g32841 and n33090_not n33096_not ; n33097
g32842 and b[20]_not n33097_not ; n33098
g32843 and n32774_not n33045_not ; n33099
g32844 and n32784_not n33012 ; n33100
g32845 and n33008_not n33100 ; n33101
g32846 and n33009_not n33012_not ; n33102
g32847 and n33101_not n33102_not ; n33103
g32848 and n4813 n33103_not ; n33104
g32849 and n33044_not n33104 ; n33105
g32850 and n33099_not n33105_not ; n33106
g32851 and b[19]_not n33106_not ; n33107
g32852 and n32783_not n33045_not ; n33108
g32853 and n32793_not n33007 ; n33109
g32854 and n33003_not n33109 ; n33110
g32855 and n33004_not n33007_not ; n33111
g32856 and n33110_not n33111_not ; n33112
g32857 and n4813 n33112_not ; n33113
g32858 and n33044_not n33113 ; n33114
g32859 and n33108_not n33114_not ; n33115
g32860 and b[18]_not n33115_not ; n33116
g32861 and n32792_not n33045_not ; n33117
g32862 and n32802_not n33002 ; n33118
g32863 and n32998_not n33118 ; n33119
g32864 and n32999_not n33002_not ; n33120
g32865 and n33119_not n33120_not ; n33121
g32866 and n4813 n33121_not ; n33122
g32867 and n33044_not n33122 ; n33123
g32868 and n33117_not n33123_not ; n33124
g32869 and b[17]_not n33124_not ; n33125
g32870 and n32801_not n33045_not ; n33126
g32871 and n32811_not n32997 ; n33127
g32872 and n32993_not n33127 ; n33128
g32873 and n32994_not n32997_not ; n33129
g32874 and n33128_not n33129_not ; n33130
g32875 and n4813 n33130_not ; n33131
g32876 and n33044_not n33131 ; n33132
g32877 and n33126_not n33132_not ; n33133
g32878 and b[16]_not n33133_not ; n33134
g32879 and n32810_not n33045_not ; n33135
g32880 and n32820_not n32992 ; n33136
g32881 and n32988_not n33136 ; n33137
g32882 and n32989_not n32992_not ; n33138
g32883 and n33137_not n33138_not ; n33139
g32884 and n4813 n33139_not ; n33140
g32885 and n33044_not n33140 ; n33141
g32886 and n33135_not n33141_not ; n33142
g32887 and b[15]_not n33142_not ; n33143
g32888 and n32819_not n33045_not ; n33144
g32889 and n32829_not n32987 ; n33145
g32890 and n32983_not n33145 ; n33146
g32891 and n32984_not n32987_not ; n33147
g32892 and n33146_not n33147_not ; n33148
g32893 and n4813 n33148_not ; n33149
g32894 and n33044_not n33149 ; n33150
g32895 and n33144_not n33150_not ; n33151
g32896 and b[14]_not n33151_not ; n33152
g32897 and n32828_not n33045_not ; n33153
g32898 and n32838_not n32982 ; n33154
g32899 and n32978_not n33154 ; n33155
g32900 and n32979_not n32982_not ; n33156
g32901 and n33155_not n33156_not ; n33157
g32902 and n4813 n33157_not ; n33158
g32903 and n33044_not n33158 ; n33159
g32904 and n33153_not n33159_not ; n33160
g32905 and b[13]_not n33160_not ; n33161
g32906 and n32837_not n33045_not ; n33162
g32907 and n32847_not n32977 ; n33163
g32908 and n32973_not n33163 ; n33164
g32909 and n32974_not n32977_not ; n33165
g32910 and n33164_not n33165_not ; n33166
g32911 and n4813 n33166_not ; n33167
g32912 and n33044_not n33167 ; n33168
g32913 and n33162_not n33168_not ; n33169
g32914 and b[12]_not n33169_not ; n33170
g32915 and n32846_not n33045_not ; n33171
g32916 and n32856_not n32972 ; n33172
g32917 and n32968_not n33172 ; n33173
g32918 and n32969_not n32972_not ; n33174
g32919 and n33173_not n33174_not ; n33175
g32920 and n4813 n33175_not ; n33176
g32921 and n33044_not n33176 ; n33177
g32922 and n33171_not n33177_not ; n33178
g32923 and b[11]_not n33178_not ; n33179
g32924 and n32855_not n33045_not ; n33180
g32925 and n32865_not n32967 ; n33181
g32926 and n32963_not n33181 ; n33182
g32927 and n32964_not n32967_not ; n33183
g32928 and n33182_not n33183_not ; n33184
g32929 and n4813 n33184_not ; n33185
g32930 and n33044_not n33185 ; n33186
g32931 and n33180_not n33186_not ; n33187
g32932 and b[10]_not n33187_not ; n33188
g32933 and n32864_not n33045_not ; n33189
g32934 and n32874_not n32962 ; n33190
g32935 and n32958_not n33190 ; n33191
g32936 and n32959_not n32962_not ; n33192
g32937 and n33191_not n33192_not ; n33193
g32938 and n4813 n33193_not ; n33194
g32939 and n33044_not n33194 ; n33195
g32940 and n33189_not n33195_not ; n33196
g32941 and b[9]_not n33196_not ; n33197
g32942 and n32873_not n33045_not ; n33198
g32943 and n32883_not n32957 ; n33199
g32944 and n32953_not n33199 ; n33200
g32945 and n32954_not n32957_not ; n33201
g32946 and n33200_not n33201_not ; n33202
g32947 and n4813 n33202_not ; n33203
g32948 and n33044_not n33203 ; n33204
g32949 and n33198_not n33204_not ; n33205
g32950 and b[8]_not n33205_not ; n33206
g32951 and n32882_not n33045_not ; n33207
g32952 and n32892_not n32952 ; n33208
g32953 and n32948_not n33208 ; n33209
g32954 and n32949_not n32952_not ; n33210
g32955 and n33209_not n33210_not ; n33211
g32956 and n4813 n33211_not ; n33212
g32957 and n33044_not n33212 ; n33213
g32958 and n33207_not n33213_not ; n33214
g32959 and b[7]_not n33214_not ; n33215
g32960 and n32891_not n33045_not ; n33216
g32961 and n32901_not n32947 ; n33217
g32962 and n32943_not n33217 ; n33218
g32963 and n32944_not n32947_not ; n33219
g32964 and n33218_not n33219_not ; n33220
g32965 and n4813 n33220_not ; n33221
g32966 and n33044_not n33221 ; n33222
g32967 and n33216_not n33222_not ; n33223
g32968 and b[6]_not n33223_not ; n33224
g32969 and n32900_not n33045_not ; n33225
g32970 and n32910_not n32942 ; n33226
g32971 and n32938_not n33226 ; n33227
g32972 and n32939_not n32942_not ; n33228
g32973 and n33227_not n33228_not ; n33229
g32974 and n4813 n33229_not ; n33230
g32975 and n33044_not n33230 ; n33231
g32976 and n33225_not n33231_not ; n33232
g32977 and b[5]_not n33232_not ; n33233
g32978 and n32909_not n33045_not ; n33234
g32979 and n32918_not n32937 ; n33235
g32980 and n32933_not n33235 ; n33236
g32981 and n32934_not n32937_not ; n33237
g32982 and n33236_not n33237_not ; n33238
g32983 and n4813 n33238_not ; n33239
g32984 and n33044_not n33239 ; n33240
g32985 and n33234_not n33240_not ; n33241
g32986 and b[4]_not n33241_not ; n33242
g32987 and n32917_not n33045_not ; n33243
g32988 and n32928_not n32932 ; n33244
g32989 and n32927_not n33244 ; n33245
g32990 and n32929_not n32932_not ; n33246
g32991 and n33245_not n33246_not ; n33247
g32992 and n4813 n33247_not ; n33248
g32993 and n33044_not n33248 ; n33249
g32994 and n33243_not n33249_not ; n33250
g32995 and b[3]_not n33250_not ; n33251
g32996 and n32922_not n33045_not ; n33252
g32997 and n4693 n32925_not ; n33253
g32998 and n32923_not n33253 ; n33254
g32999 and n4813 n33254_not ; n33255
g33000 and n32927_not n33255 ; n33256
g33001 and n33044_not n33256 ; n33257
g33002 and n33252_not n33257_not ; n33258
g33003 and b[2]_not n33258_not ; n33259
g33004 and n5033 n33044_not ; n33260
g33005 and a[39] n33260_not ; n33261
g33006 and n5039 n33044_not ; n33262
g33007 and n33261_not n33262_not ; n33263
g33008 and b[1] n33263_not ; n33264
g33009 and b[1]_not n33262_not ; n33265
g33010 and n33261_not n33265 ; n33266
g33011 and n33264_not n33266_not ; n33267
g33012 and n5046_not n33267_not ; n33268
g33013 and b[1]_not n33263_not ; n33269
g33014 and n33268_not n33269_not ; n33270
g33015 and b[2] n33257_not ; n33271
g33016 and n33252_not n33271 ; n33272
g33017 and n33259_not n33272_not ; n33273
g33018 and n33270_not n33273 ; n33274
g33019 and n33259_not n33274_not ; n33275
g33020 and b[3] n33249_not ; n33276
g33021 and n33243_not n33276 ; n33277
g33022 and n33251_not n33277_not ; n33278
g33023 and n33275_not n33278 ; n33279
g33024 and n33251_not n33279_not ; n33280
g33025 and b[4] n33240_not ; n33281
g33026 and n33234_not n33281 ; n33282
g33027 and n33242_not n33282_not ; n33283
g33028 and n33280_not n33283 ; n33284
g33029 and n33242_not n33284_not ; n33285
g33030 and b[5] n33231_not ; n33286
g33031 and n33225_not n33286 ; n33287
g33032 and n33233_not n33287_not ; n33288
g33033 and n33285_not n33288 ; n33289
g33034 and n33233_not n33289_not ; n33290
g33035 and b[6] n33222_not ; n33291
g33036 and n33216_not n33291 ; n33292
g33037 and n33224_not n33292_not ; n33293
g33038 and n33290_not n33293 ; n33294
g33039 and n33224_not n33294_not ; n33295
g33040 and b[7] n33213_not ; n33296
g33041 and n33207_not n33296 ; n33297
g33042 and n33215_not n33297_not ; n33298
g33043 and n33295_not n33298 ; n33299
g33044 and n33215_not n33299_not ; n33300
g33045 and b[8] n33204_not ; n33301
g33046 and n33198_not n33301 ; n33302
g33047 and n33206_not n33302_not ; n33303
g33048 and n33300_not n33303 ; n33304
g33049 and n33206_not n33304_not ; n33305
g33050 and b[9] n33195_not ; n33306
g33051 and n33189_not n33306 ; n33307
g33052 and n33197_not n33307_not ; n33308
g33053 and n33305_not n33308 ; n33309
g33054 and n33197_not n33309_not ; n33310
g33055 and b[10] n33186_not ; n33311
g33056 and n33180_not n33311 ; n33312
g33057 and n33188_not n33312_not ; n33313
g33058 and n33310_not n33313 ; n33314
g33059 and n33188_not n33314_not ; n33315
g33060 and b[11] n33177_not ; n33316
g33061 and n33171_not n33316 ; n33317
g33062 and n33179_not n33317_not ; n33318
g33063 and n33315_not n33318 ; n33319
g33064 and n33179_not n33319_not ; n33320
g33065 and b[12] n33168_not ; n33321
g33066 and n33162_not n33321 ; n33322
g33067 and n33170_not n33322_not ; n33323
g33068 and n33320_not n33323 ; n33324
g33069 and n33170_not n33324_not ; n33325
g33070 and b[13] n33159_not ; n33326
g33071 and n33153_not n33326 ; n33327
g33072 and n33161_not n33327_not ; n33328
g33073 and n33325_not n33328 ; n33329
g33074 and n33161_not n33329_not ; n33330
g33075 and b[14] n33150_not ; n33331
g33076 and n33144_not n33331 ; n33332
g33077 and n33152_not n33332_not ; n33333
g33078 and n33330_not n33333 ; n33334
g33079 and n33152_not n33334_not ; n33335
g33080 and b[15] n33141_not ; n33336
g33081 and n33135_not n33336 ; n33337
g33082 and n33143_not n33337_not ; n33338
g33083 and n33335_not n33338 ; n33339
g33084 and n33143_not n33339_not ; n33340
g33085 and b[16] n33132_not ; n33341
g33086 and n33126_not n33341 ; n33342
g33087 and n33134_not n33342_not ; n33343
g33088 and n33340_not n33343 ; n33344
g33089 and n33134_not n33344_not ; n33345
g33090 and b[17] n33123_not ; n33346
g33091 and n33117_not n33346 ; n33347
g33092 and n33125_not n33347_not ; n33348
g33093 and n33345_not n33348 ; n33349
g33094 and n33125_not n33349_not ; n33350
g33095 and b[18] n33114_not ; n33351
g33096 and n33108_not n33351 ; n33352
g33097 and n33116_not n33352_not ; n33353
g33098 and n33350_not n33353 ; n33354
g33099 and n33116_not n33354_not ; n33355
g33100 and b[19] n33105_not ; n33356
g33101 and n33099_not n33356 ; n33357
g33102 and n33107_not n33357_not ; n33358
g33103 and n33355_not n33358 ; n33359
g33104 and n33107_not n33359_not ; n33360
g33105 and b[20] n33096_not ; n33361
g33106 and n33090_not n33361 ; n33362
g33107 and n33098_not n33362_not ; n33363
g33108 and n33360_not n33363 ; n33364
g33109 and n33098_not n33364_not ; n33365
g33110 and b[21] n33087_not ; n33366
g33111 and n33081_not n33366 ; n33367
g33112 and n33089_not n33367_not ; n33368
g33113 and n33365_not n33368 ; n33369
g33114 and n33089_not n33369_not ; n33370
g33115 and b[22] n33078_not ; n33371
g33116 and n33072_not n33371 ; n33372
g33117 and n33080_not n33372_not ; n33373
g33118 and n33370_not n33373 ; n33374
g33119 and n33080_not n33374_not ; n33375
g33120 and b[23] n33069_not ; n33376
g33121 and n33063_not n33376 ; n33377
g33122 and n33071_not n33377_not ; n33378
g33123 and n33375_not n33378 ; n33379
g33124 and n33071_not n33379_not ; n33380
g33125 and b[24] n33052_not ; n33381
g33126 and n33046_not n33381 ; n33382
g33127 and n33062_not n33382_not ; n33383
g33128 and n33380_not n33383 ; n33384
g33129 and n33062_not n33384_not ; n33385
g33130 and b[25] n33054_not ; n33386
g33131 and n33059_not n33386 ; n33387
g33132 and n33061_not n33387_not ; n33388
g33133 and n33385_not n33388 ; n33389
g33134 and n33061_not n33389_not ; n33390
g33135 and n5172 n33390_not ; n33391
g33136 and n33053_not n33391_not ; n33392
g33137 and n33071_not n33383 ; n33393
g33138 and n33379_not n33393 ; n33394
g33139 and n33380_not n33383_not ; n33395
g33140 and n33394_not n33395_not ; n33396
g33141 and n5172 n33396_not ; n33397
g33142 and n33390_not n33397 ; n33398
g33143 and n33392_not n33398_not ; n33399
g33144 and b[25]_not n33399_not ; n33400
g33145 and n33070_not n33391_not ; n33401
g33146 and n33080_not n33378 ; n33402
g33147 and n33374_not n33402 ; n33403
g33148 and n33375_not n33378_not ; n33404
g33149 and n33403_not n33404_not ; n33405
g33150 and n5172 n33405_not ; n33406
g33151 and n33390_not n33406 ; n33407
g33152 and n33401_not n33407_not ; n33408
g33153 and b[24]_not n33408_not ; n33409
g33154 and n33079_not n33391_not ; n33410
g33155 and n33089_not n33373 ; n33411
g33156 and n33369_not n33411 ; n33412
g33157 and n33370_not n33373_not ; n33413
g33158 and n33412_not n33413_not ; n33414
g33159 and n5172 n33414_not ; n33415
g33160 and n33390_not n33415 ; n33416
g33161 and n33410_not n33416_not ; n33417
g33162 and b[23]_not n33417_not ; n33418
g33163 and n33088_not n33391_not ; n33419
g33164 and n33098_not n33368 ; n33420
g33165 and n33364_not n33420 ; n33421
g33166 and n33365_not n33368_not ; n33422
g33167 and n33421_not n33422_not ; n33423
g33168 and n5172 n33423_not ; n33424
g33169 and n33390_not n33424 ; n33425
g33170 and n33419_not n33425_not ; n33426
g33171 and b[22]_not n33426_not ; n33427
g33172 and n33097_not n33391_not ; n33428
g33173 and n33107_not n33363 ; n33429
g33174 and n33359_not n33429 ; n33430
g33175 and n33360_not n33363_not ; n33431
g33176 and n33430_not n33431_not ; n33432
g33177 and n5172 n33432_not ; n33433
g33178 and n33390_not n33433 ; n33434
g33179 and n33428_not n33434_not ; n33435
g33180 and b[21]_not n33435_not ; n33436
g33181 and n33106_not n33391_not ; n33437
g33182 and n33116_not n33358 ; n33438
g33183 and n33354_not n33438 ; n33439
g33184 and n33355_not n33358_not ; n33440
g33185 and n33439_not n33440_not ; n33441
g33186 and n5172 n33441_not ; n33442
g33187 and n33390_not n33442 ; n33443
g33188 and n33437_not n33443_not ; n33444
g33189 and b[20]_not n33444_not ; n33445
g33190 and n33115_not n33391_not ; n33446
g33191 and n33125_not n33353 ; n33447
g33192 and n33349_not n33447 ; n33448
g33193 and n33350_not n33353_not ; n33449
g33194 and n33448_not n33449_not ; n33450
g33195 and n5172 n33450_not ; n33451
g33196 and n33390_not n33451 ; n33452
g33197 and n33446_not n33452_not ; n33453
g33198 and b[19]_not n33453_not ; n33454
g33199 and n33124_not n33391_not ; n33455
g33200 and n33134_not n33348 ; n33456
g33201 and n33344_not n33456 ; n33457
g33202 and n33345_not n33348_not ; n33458
g33203 and n33457_not n33458_not ; n33459
g33204 and n5172 n33459_not ; n33460
g33205 and n33390_not n33460 ; n33461
g33206 and n33455_not n33461_not ; n33462
g33207 and b[18]_not n33462_not ; n33463
g33208 and n33133_not n33391_not ; n33464
g33209 and n33143_not n33343 ; n33465
g33210 and n33339_not n33465 ; n33466
g33211 and n33340_not n33343_not ; n33467
g33212 and n33466_not n33467_not ; n33468
g33213 and n5172 n33468_not ; n33469
g33214 and n33390_not n33469 ; n33470
g33215 and n33464_not n33470_not ; n33471
g33216 and b[17]_not n33471_not ; n33472
g33217 and n33142_not n33391_not ; n33473
g33218 and n33152_not n33338 ; n33474
g33219 and n33334_not n33474 ; n33475
g33220 and n33335_not n33338_not ; n33476
g33221 and n33475_not n33476_not ; n33477
g33222 and n5172 n33477_not ; n33478
g33223 and n33390_not n33478 ; n33479
g33224 and n33473_not n33479_not ; n33480
g33225 and b[16]_not n33480_not ; n33481
g33226 and n33151_not n33391_not ; n33482
g33227 and n33161_not n33333 ; n33483
g33228 and n33329_not n33483 ; n33484
g33229 and n33330_not n33333_not ; n33485
g33230 and n33484_not n33485_not ; n33486
g33231 and n5172 n33486_not ; n33487
g33232 and n33390_not n33487 ; n33488
g33233 and n33482_not n33488_not ; n33489
g33234 and b[15]_not n33489_not ; n33490
g33235 and n33160_not n33391_not ; n33491
g33236 and n33170_not n33328 ; n33492
g33237 and n33324_not n33492 ; n33493
g33238 and n33325_not n33328_not ; n33494
g33239 and n33493_not n33494_not ; n33495
g33240 and n5172 n33495_not ; n33496
g33241 and n33390_not n33496 ; n33497
g33242 and n33491_not n33497_not ; n33498
g33243 and b[14]_not n33498_not ; n33499
g33244 and n33169_not n33391_not ; n33500
g33245 and n33179_not n33323 ; n33501
g33246 and n33319_not n33501 ; n33502
g33247 and n33320_not n33323_not ; n33503
g33248 and n33502_not n33503_not ; n33504
g33249 and n5172 n33504_not ; n33505
g33250 and n33390_not n33505 ; n33506
g33251 and n33500_not n33506_not ; n33507
g33252 and b[13]_not n33507_not ; n33508
g33253 and n33178_not n33391_not ; n33509
g33254 and n33188_not n33318 ; n33510
g33255 and n33314_not n33510 ; n33511
g33256 and n33315_not n33318_not ; n33512
g33257 and n33511_not n33512_not ; n33513
g33258 and n5172 n33513_not ; n33514
g33259 and n33390_not n33514 ; n33515
g33260 and n33509_not n33515_not ; n33516
g33261 and b[12]_not n33516_not ; n33517
g33262 and n33187_not n33391_not ; n33518
g33263 and n33197_not n33313 ; n33519
g33264 and n33309_not n33519 ; n33520
g33265 and n33310_not n33313_not ; n33521
g33266 and n33520_not n33521_not ; n33522
g33267 and n5172 n33522_not ; n33523
g33268 and n33390_not n33523 ; n33524
g33269 and n33518_not n33524_not ; n33525
g33270 and b[11]_not n33525_not ; n33526
g33271 and n33196_not n33391_not ; n33527
g33272 and n33206_not n33308 ; n33528
g33273 and n33304_not n33528 ; n33529
g33274 and n33305_not n33308_not ; n33530
g33275 and n33529_not n33530_not ; n33531
g33276 and n5172 n33531_not ; n33532
g33277 and n33390_not n33532 ; n33533
g33278 and n33527_not n33533_not ; n33534
g33279 and b[10]_not n33534_not ; n33535
g33280 and n33205_not n33391_not ; n33536
g33281 and n33215_not n33303 ; n33537
g33282 and n33299_not n33537 ; n33538
g33283 and n33300_not n33303_not ; n33539
g33284 and n33538_not n33539_not ; n33540
g33285 and n5172 n33540_not ; n33541
g33286 and n33390_not n33541 ; n33542
g33287 and n33536_not n33542_not ; n33543
g33288 and b[9]_not n33543_not ; n33544
g33289 and n33214_not n33391_not ; n33545
g33290 and n33224_not n33298 ; n33546
g33291 and n33294_not n33546 ; n33547
g33292 and n33295_not n33298_not ; n33548
g33293 and n33547_not n33548_not ; n33549
g33294 and n5172 n33549_not ; n33550
g33295 and n33390_not n33550 ; n33551
g33296 and n33545_not n33551_not ; n33552
g33297 and b[8]_not n33552_not ; n33553
g33298 and n33223_not n33391_not ; n33554
g33299 and n33233_not n33293 ; n33555
g33300 and n33289_not n33555 ; n33556
g33301 and n33290_not n33293_not ; n33557
g33302 and n33556_not n33557_not ; n33558
g33303 and n5172 n33558_not ; n33559
g33304 and n33390_not n33559 ; n33560
g33305 and n33554_not n33560_not ; n33561
g33306 and b[7]_not n33561_not ; n33562
g33307 and n33232_not n33391_not ; n33563
g33308 and n33242_not n33288 ; n33564
g33309 and n33284_not n33564 ; n33565
g33310 and n33285_not n33288_not ; n33566
g33311 and n33565_not n33566_not ; n33567
g33312 and n5172 n33567_not ; n33568
g33313 and n33390_not n33568 ; n33569
g33314 and n33563_not n33569_not ; n33570
g33315 and b[6]_not n33570_not ; n33571
g33316 and n33241_not n33391_not ; n33572
g33317 and n33251_not n33283 ; n33573
g33318 and n33279_not n33573 ; n33574
g33319 and n33280_not n33283_not ; n33575
g33320 and n33574_not n33575_not ; n33576
g33321 and n5172 n33576_not ; n33577
g33322 and n33390_not n33577 ; n33578
g33323 and n33572_not n33578_not ; n33579
g33324 and b[5]_not n33579_not ; n33580
g33325 and n33250_not n33391_not ; n33581
g33326 and n33259_not n33278 ; n33582
g33327 and n33274_not n33582 ; n33583
g33328 and n33275_not n33278_not ; n33584
g33329 and n33583_not n33584_not ; n33585
g33330 and n5172 n33585_not ; n33586
g33331 and n33390_not n33586 ; n33587
g33332 and n33581_not n33587_not ; n33588
g33333 and b[4]_not n33588_not ; n33589
g33334 and n33258_not n33391_not ; n33590
g33335 and n33269_not n33273 ; n33591
g33336 and n33268_not n33591 ; n33592
g33337 and n33270_not n33273_not ; n33593
g33338 and n33592_not n33593_not ; n33594
g33339 and n5172 n33594_not ; n33595
g33340 and n33390_not n33595 ; n33596
g33341 and n33590_not n33596_not ; n33597
g33342 and b[3]_not n33597_not ; n33598
g33343 and n33263_not n33391_not ; n33599
g33344 and n5046 n33266_not ; n33600
g33345 and n33264_not n33600 ; n33601
g33346 and n5172 n33601_not ; n33602
g33347 and n33268_not n33602 ; n33603
g33348 and n33390_not n33603 ; n33604
g33349 and n33599_not n33604_not ; n33605
g33350 and b[2]_not n33605_not ; n33606
g33351 and n5393 n33390_not ; n33607
g33352 and a[38] n33607_not ; n33608
g33353 and n5399 n33390_not ; n33609
g33354 and n33608_not n33609_not ; n33610
g33355 and b[1] n33610_not ; n33611
g33356 and b[1]_not n33609_not ; n33612
g33357 and n33608_not n33612 ; n33613
g33358 and n33611_not n33613_not ; n33614
g33359 and n5406_not n33614_not ; n33615
g33360 and b[1]_not n33610_not ; n33616
g33361 and n33615_not n33616_not ; n33617
g33362 and b[2] n33604_not ; n33618
g33363 and n33599_not n33618 ; n33619
g33364 and n33606_not n33619_not ; n33620
g33365 and n33617_not n33620 ; n33621
g33366 and n33606_not n33621_not ; n33622
g33367 and b[3] n33596_not ; n33623
g33368 and n33590_not n33623 ; n33624
g33369 and n33598_not n33624_not ; n33625
g33370 and n33622_not n33625 ; n33626
g33371 and n33598_not n33626_not ; n33627
g33372 and b[4] n33587_not ; n33628
g33373 and n33581_not n33628 ; n33629
g33374 and n33589_not n33629_not ; n33630
g33375 and n33627_not n33630 ; n33631
g33376 and n33589_not n33631_not ; n33632
g33377 and b[5] n33578_not ; n33633
g33378 and n33572_not n33633 ; n33634
g33379 and n33580_not n33634_not ; n33635
g33380 and n33632_not n33635 ; n33636
g33381 and n33580_not n33636_not ; n33637
g33382 and b[6] n33569_not ; n33638
g33383 and n33563_not n33638 ; n33639
g33384 and n33571_not n33639_not ; n33640
g33385 and n33637_not n33640 ; n33641
g33386 and n33571_not n33641_not ; n33642
g33387 and b[7] n33560_not ; n33643
g33388 and n33554_not n33643 ; n33644
g33389 and n33562_not n33644_not ; n33645
g33390 and n33642_not n33645 ; n33646
g33391 and n33562_not n33646_not ; n33647
g33392 and b[8] n33551_not ; n33648
g33393 and n33545_not n33648 ; n33649
g33394 and n33553_not n33649_not ; n33650
g33395 and n33647_not n33650 ; n33651
g33396 and n33553_not n33651_not ; n33652
g33397 and b[9] n33542_not ; n33653
g33398 and n33536_not n33653 ; n33654
g33399 and n33544_not n33654_not ; n33655
g33400 and n33652_not n33655 ; n33656
g33401 and n33544_not n33656_not ; n33657
g33402 and b[10] n33533_not ; n33658
g33403 and n33527_not n33658 ; n33659
g33404 and n33535_not n33659_not ; n33660
g33405 and n33657_not n33660 ; n33661
g33406 and n33535_not n33661_not ; n33662
g33407 and b[11] n33524_not ; n33663
g33408 and n33518_not n33663 ; n33664
g33409 and n33526_not n33664_not ; n33665
g33410 and n33662_not n33665 ; n33666
g33411 and n33526_not n33666_not ; n33667
g33412 and b[12] n33515_not ; n33668
g33413 and n33509_not n33668 ; n33669
g33414 and n33517_not n33669_not ; n33670
g33415 and n33667_not n33670 ; n33671
g33416 and n33517_not n33671_not ; n33672
g33417 and b[13] n33506_not ; n33673
g33418 and n33500_not n33673 ; n33674
g33419 and n33508_not n33674_not ; n33675
g33420 and n33672_not n33675 ; n33676
g33421 and n33508_not n33676_not ; n33677
g33422 and b[14] n33497_not ; n33678
g33423 and n33491_not n33678 ; n33679
g33424 and n33499_not n33679_not ; n33680
g33425 and n33677_not n33680 ; n33681
g33426 and n33499_not n33681_not ; n33682
g33427 and b[15] n33488_not ; n33683
g33428 and n33482_not n33683 ; n33684
g33429 and n33490_not n33684_not ; n33685
g33430 and n33682_not n33685 ; n33686
g33431 and n33490_not n33686_not ; n33687
g33432 and b[16] n33479_not ; n33688
g33433 and n33473_not n33688 ; n33689
g33434 and n33481_not n33689_not ; n33690
g33435 and n33687_not n33690 ; n33691
g33436 and n33481_not n33691_not ; n33692
g33437 and b[17] n33470_not ; n33693
g33438 and n33464_not n33693 ; n33694
g33439 and n33472_not n33694_not ; n33695
g33440 and n33692_not n33695 ; n33696
g33441 and n33472_not n33696_not ; n33697
g33442 and b[18] n33461_not ; n33698
g33443 and n33455_not n33698 ; n33699
g33444 and n33463_not n33699_not ; n33700
g33445 and n33697_not n33700 ; n33701
g33446 and n33463_not n33701_not ; n33702
g33447 and b[19] n33452_not ; n33703
g33448 and n33446_not n33703 ; n33704
g33449 and n33454_not n33704_not ; n33705
g33450 and n33702_not n33705 ; n33706
g33451 and n33454_not n33706_not ; n33707
g33452 and b[20] n33443_not ; n33708
g33453 and n33437_not n33708 ; n33709
g33454 and n33445_not n33709_not ; n33710
g33455 and n33707_not n33710 ; n33711
g33456 and n33445_not n33711_not ; n33712
g33457 and b[21] n33434_not ; n33713
g33458 and n33428_not n33713 ; n33714
g33459 and n33436_not n33714_not ; n33715
g33460 and n33712_not n33715 ; n33716
g33461 and n33436_not n33716_not ; n33717
g33462 and b[22] n33425_not ; n33718
g33463 and n33419_not n33718 ; n33719
g33464 and n33427_not n33719_not ; n33720
g33465 and n33717_not n33720 ; n33721
g33466 and n33427_not n33721_not ; n33722
g33467 and b[23] n33416_not ; n33723
g33468 and n33410_not n33723 ; n33724
g33469 and n33418_not n33724_not ; n33725
g33470 and n33722_not n33725 ; n33726
g33471 and n33418_not n33726_not ; n33727
g33472 and b[24] n33407_not ; n33728
g33473 and n33401_not n33728 ; n33729
g33474 and n33409_not n33729_not ; n33730
g33475 and n33727_not n33730 ; n33731
g33476 and n33409_not n33731_not ; n33732
g33477 and b[25] n33398_not ; n33733
g33478 and n33392_not n33733 ; n33734
g33479 and n33400_not n33734_not ; n33735
g33480 and n33732_not n33735 ; n33736
g33481 and n33400_not n33736_not ; n33737
g33482 and n33060_not n33391_not ; n33738
g33483 and n33062_not n33388 ; n33739
g33484 and n33384_not n33739 ; n33740
g33485 and n33385_not n33388_not ; n33741
g33486 and n33740_not n33741_not ; n33742
g33487 and n33391 n33742_not ; n33743
g33488 and n33738_not n33743_not ; n33744
g33489 and b[26]_not n33744_not ; n33745
g33490 and b[26] n33738_not ; n33746
g33491 and n33743_not n33746 ; n33747
g33492 and n5542 n33747_not ; n33748
g33493 and n33745_not n33748 ; n33749
g33494 and n33737_not n33749 ; n33750
g33495 and n5172 n33744_not ; n33751
g33496 and n33750_not n33751_not ; n33752
g33497 and n33409_not n33735 ; n33753
g33498 and n33731_not n33753 ; n33754
g33499 and n33732_not n33735_not ; n33755
g33500 and n33754_not n33755_not ; n33756
g33501 and n33752_not n33756_not ; n33757
g33502 and n33399_not n33751_not ; n33758
g33503 and n33750_not n33758 ; n33759
g33504 and n33757_not n33759_not ; n33760
g33505 and n33400_not n33747_not ; n33761
g33506 and n33745_not n33761 ; n33762
g33507 and n33736_not n33762 ; n33763
g33508 and n33745_not n33747_not ; n33764
g33509 and n33737_not n33764_not ; n33765
g33510 and n33763_not n33765_not ; n33766
g33511 and n33752_not n33766_not ; n33767
g33512 and n33744_not n33751_not ; n33768
g33513 and n33750_not n33768 ; n33769
g33514 and n33767_not n33769_not ; n33770
g33515 and b[27]_not n33770_not ; n33771
g33516 and b[26]_not n33760_not ; n33772
g33517 and n33418_not n33730 ; n33773
g33518 and n33726_not n33773 ; n33774
g33519 and n33727_not n33730_not ; n33775
g33520 and n33774_not n33775_not ; n33776
g33521 and n33752_not n33776_not ; n33777
g33522 and n33408_not n33751_not ; n33778
g33523 and n33750_not n33778 ; n33779
g33524 and n33777_not n33779_not ; n33780
g33525 and b[25]_not n33780_not ; n33781
g33526 and n33427_not n33725 ; n33782
g33527 and n33721_not n33782 ; n33783
g33528 and n33722_not n33725_not ; n33784
g33529 and n33783_not n33784_not ; n33785
g33530 and n33752_not n33785_not ; n33786
g33531 and n33417_not n33751_not ; n33787
g33532 and n33750_not n33787 ; n33788
g33533 and n33786_not n33788_not ; n33789
g33534 and b[24]_not n33789_not ; n33790
g33535 and n33436_not n33720 ; n33791
g33536 and n33716_not n33791 ; n33792
g33537 and n33717_not n33720_not ; n33793
g33538 and n33792_not n33793_not ; n33794
g33539 and n33752_not n33794_not ; n33795
g33540 and n33426_not n33751_not ; n33796
g33541 and n33750_not n33796 ; n33797
g33542 and n33795_not n33797_not ; n33798
g33543 and b[23]_not n33798_not ; n33799
g33544 and n33445_not n33715 ; n33800
g33545 and n33711_not n33800 ; n33801
g33546 and n33712_not n33715_not ; n33802
g33547 and n33801_not n33802_not ; n33803
g33548 and n33752_not n33803_not ; n33804
g33549 and n33435_not n33751_not ; n33805
g33550 and n33750_not n33805 ; n33806
g33551 and n33804_not n33806_not ; n33807
g33552 and b[22]_not n33807_not ; n33808
g33553 and n33454_not n33710 ; n33809
g33554 and n33706_not n33809 ; n33810
g33555 and n33707_not n33710_not ; n33811
g33556 and n33810_not n33811_not ; n33812
g33557 and n33752_not n33812_not ; n33813
g33558 and n33444_not n33751_not ; n33814
g33559 and n33750_not n33814 ; n33815
g33560 and n33813_not n33815_not ; n33816
g33561 and b[21]_not n33816_not ; n33817
g33562 and n33463_not n33705 ; n33818
g33563 and n33701_not n33818 ; n33819
g33564 and n33702_not n33705_not ; n33820
g33565 and n33819_not n33820_not ; n33821
g33566 and n33752_not n33821_not ; n33822
g33567 and n33453_not n33751_not ; n33823
g33568 and n33750_not n33823 ; n33824
g33569 and n33822_not n33824_not ; n33825
g33570 and b[20]_not n33825_not ; n33826
g33571 and n33472_not n33700 ; n33827
g33572 and n33696_not n33827 ; n33828
g33573 and n33697_not n33700_not ; n33829
g33574 and n33828_not n33829_not ; n33830
g33575 and n33752_not n33830_not ; n33831
g33576 and n33462_not n33751_not ; n33832
g33577 and n33750_not n33832 ; n33833
g33578 and n33831_not n33833_not ; n33834
g33579 and b[19]_not n33834_not ; n33835
g33580 and n33481_not n33695 ; n33836
g33581 and n33691_not n33836 ; n33837
g33582 and n33692_not n33695_not ; n33838
g33583 and n33837_not n33838_not ; n33839
g33584 and n33752_not n33839_not ; n33840
g33585 and n33471_not n33751_not ; n33841
g33586 and n33750_not n33841 ; n33842
g33587 and n33840_not n33842_not ; n33843
g33588 and b[18]_not n33843_not ; n33844
g33589 and n33490_not n33690 ; n33845
g33590 and n33686_not n33845 ; n33846
g33591 and n33687_not n33690_not ; n33847
g33592 and n33846_not n33847_not ; n33848
g33593 and n33752_not n33848_not ; n33849
g33594 and n33480_not n33751_not ; n33850
g33595 and n33750_not n33850 ; n33851
g33596 and n33849_not n33851_not ; n33852
g33597 and b[17]_not n33852_not ; n33853
g33598 and n33499_not n33685 ; n33854
g33599 and n33681_not n33854 ; n33855
g33600 and n33682_not n33685_not ; n33856
g33601 and n33855_not n33856_not ; n33857
g33602 and n33752_not n33857_not ; n33858
g33603 and n33489_not n33751_not ; n33859
g33604 and n33750_not n33859 ; n33860
g33605 and n33858_not n33860_not ; n33861
g33606 and b[16]_not n33861_not ; n33862
g33607 and n33508_not n33680 ; n33863
g33608 and n33676_not n33863 ; n33864
g33609 and n33677_not n33680_not ; n33865
g33610 and n33864_not n33865_not ; n33866
g33611 and n33752_not n33866_not ; n33867
g33612 and n33498_not n33751_not ; n33868
g33613 and n33750_not n33868 ; n33869
g33614 and n33867_not n33869_not ; n33870
g33615 and b[15]_not n33870_not ; n33871
g33616 and n33517_not n33675 ; n33872
g33617 and n33671_not n33872 ; n33873
g33618 and n33672_not n33675_not ; n33874
g33619 and n33873_not n33874_not ; n33875
g33620 and n33752_not n33875_not ; n33876
g33621 and n33507_not n33751_not ; n33877
g33622 and n33750_not n33877 ; n33878
g33623 and n33876_not n33878_not ; n33879
g33624 and b[14]_not n33879_not ; n33880
g33625 and n33526_not n33670 ; n33881
g33626 and n33666_not n33881 ; n33882
g33627 and n33667_not n33670_not ; n33883
g33628 and n33882_not n33883_not ; n33884
g33629 and n33752_not n33884_not ; n33885
g33630 and n33516_not n33751_not ; n33886
g33631 and n33750_not n33886 ; n33887
g33632 and n33885_not n33887_not ; n33888
g33633 and b[13]_not n33888_not ; n33889
g33634 and n33535_not n33665 ; n33890
g33635 and n33661_not n33890 ; n33891
g33636 and n33662_not n33665_not ; n33892
g33637 and n33891_not n33892_not ; n33893
g33638 and n33752_not n33893_not ; n33894
g33639 and n33525_not n33751_not ; n33895
g33640 and n33750_not n33895 ; n33896
g33641 and n33894_not n33896_not ; n33897
g33642 and b[12]_not n33897_not ; n33898
g33643 and n33544_not n33660 ; n33899
g33644 and n33656_not n33899 ; n33900
g33645 and n33657_not n33660_not ; n33901
g33646 and n33900_not n33901_not ; n33902
g33647 and n33752_not n33902_not ; n33903
g33648 and n33534_not n33751_not ; n33904
g33649 and n33750_not n33904 ; n33905
g33650 and n33903_not n33905_not ; n33906
g33651 and b[11]_not n33906_not ; n33907
g33652 and n33553_not n33655 ; n33908
g33653 and n33651_not n33908 ; n33909
g33654 and n33652_not n33655_not ; n33910
g33655 and n33909_not n33910_not ; n33911
g33656 and n33752_not n33911_not ; n33912
g33657 and n33543_not n33751_not ; n33913
g33658 and n33750_not n33913 ; n33914
g33659 and n33912_not n33914_not ; n33915
g33660 and b[10]_not n33915_not ; n33916
g33661 and n33562_not n33650 ; n33917
g33662 and n33646_not n33917 ; n33918
g33663 and n33647_not n33650_not ; n33919
g33664 and n33918_not n33919_not ; n33920
g33665 and n33752_not n33920_not ; n33921
g33666 and n33552_not n33751_not ; n33922
g33667 and n33750_not n33922 ; n33923
g33668 and n33921_not n33923_not ; n33924
g33669 and b[9]_not n33924_not ; n33925
g33670 and n33571_not n33645 ; n33926
g33671 and n33641_not n33926 ; n33927
g33672 and n33642_not n33645_not ; n33928
g33673 and n33927_not n33928_not ; n33929
g33674 and n33752_not n33929_not ; n33930
g33675 and n33561_not n33751_not ; n33931
g33676 and n33750_not n33931 ; n33932
g33677 and n33930_not n33932_not ; n33933
g33678 and b[8]_not n33933_not ; n33934
g33679 and n33580_not n33640 ; n33935
g33680 and n33636_not n33935 ; n33936
g33681 and n33637_not n33640_not ; n33937
g33682 and n33936_not n33937_not ; n33938
g33683 and n33752_not n33938_not ; n33939
g33684 and n33570_not n33751_not ; n33940
g33685 and n33750_not n33940 ; n33941
g33686 and n33939_not n33941_not ; n33942
g33687 and b[7]_not n33942_not ; n33943
g33688 and n33589_not n33635 ; n33944
g33689 and n33631_not n33944 ; n33945
g33690 and n33632_not n33635_not ; n33946
g33691 and n33945_not n33946_not ; n33947
g33692 and n33752_not n33947_not ; n33948
g33693 and n33579_not n33751_not ; n33949
g33694 and n33750_not n33949 ; n33950
g33695 and n33948_not n33950_not ; n33951
g33696 and b[6]_not n33951_not ; n33952
g33697 and n33598_not n33630 ; n33953
g33698 and n33626_not n33953 ; n33954
g33699 and n33627_not n33630_not ; n33955
g33700 and n33954_not n33955_not ; n33956
g33701 and n33752_not n33956_not ; n33957
g33702 and n33588_not n33751_not ; n33958
g33703 and n33750_not n33958 ; n33959
g33704 and n33957_not n33959_not ; n33960
g33705 and b[5]_not n33960_not ; n33961
g33706 and n33606_not n33625 ; n33962
g33707 and n33621_not n33962 ; n33963
g33708 and n33622_not n33625_not ; n33964
g33709 and n33963_not n33964_not ; n33965
g33710 and n33752_not n33965_not ; n33966
g33711 and n33597_not n33751_not ; n33967
g33712 and n33750_not n33967 ; n33968
g33713 and n33966_not n33968_not ; n33969
g33714 and b[4]_not n33969_not ; n33970
g33715 and n33616_not n33620 ; n33971
g33716 and n33615_not n33971 ; n33972
g33717 and n33617_not n33620_not ; n33973
g33718 and n33972_not n33973_not ; n33974
g33719 and n33752_not n33974_not ; n33975
g33720 and n33605_not n33751_not ; n33976
g33721 and n33750_not n33976 ; n33977
g33722 and n33975_not n33977_not ; n33978
g33723 and b[3]_not n33978_not ; n33979
g33724 and n5406 n33613_not ; n33980
g33725 and n33611_not n33980 ; n33981
g33726 and n33615_not n33981_not ; n33982
g33727 and n33752_not n33982 ; n33983
g33728 and n33610_not n33751_not ; n33984
g33729 and n33750_not n33984 ; n33985
g33730 and n33983_not n33985_not ; n33986
g33731 and b[2]_not n33986_not ; n33987
g33732 and b[0] n33752_not ; n33988
g33733 and a[37] n33988_not ; n33989
g33734 and n5406 n33752_not ; n33990
g33735 and n33989_not n33990_not ; n33991
g33736 and b[1] n33991_not ; n33992
g33737 and b[1]_not n33990_not ; n33993
g33738 and n33989_not n33993 ; n33994
g33739 and n33992_not n33994_not ; n33995
g33740 and n5791_not n33995_not ; n33996
g33741 and b[1]_not n33991_not ; n33997
g33742 and n33996_not n33997_not ; n33998
g33743 and b[2] n33985_not ; n33999
g33744 and n33983_not n33999 ; n34000
g33745 and n33987_not n34000_not ; n34001
g33746 and n33998_not n34001 ; n34002
g33747 and n33987_not n34002_not ; n34003
g33748 and b[3] n33977_not ; n34004
g33749 and n33975_not n34004 ; n34005
g33750 and n33979_not n34005_not ; n34006
g33751 and n34003_not n34006 ; n34007
g33752 and n33979_not n34007_not ; n34008
g33753 and b[4] n33968_not ; n34009
g33754 and n33966_not n34009 ; n34010
g33755 and n33970_not n34010_not ; n34011
g33756 and n34008_not n34011 ; n34012
g33757 and n33970_not n34012_not ; n34013
g33758 and b[5] n33959_not ; n34014
g33759 and n33957_not n34014 ; n34015
g33760 and n33961_not n34015_not ; n34016
g33761 and n34013_not n34016 ; n34017
g33762 and n33961_not n34017_not ; n34018
g33763 and b[6] n33950_not ; n34019
g33764 and n33948_not n34019 ; n34020
g33765 and n33952_not n34020_not ; n34021
g33766 and n34018_not n34021 ; n34022
g33767 and n33952_not n34022_not ; n34023
g33768 and b[7] n33941_not ; n34024
g33769 and n33939_not n34024 ; n34025
g33770 and n33943_not n34025_not ; n34026
g33771 and n34023_not n34026 ; n34027
g33772 and n33943_not n34027_not ; n34028
g33773 and b[8] n33932_not ; n34029
g33774 and n33930_not n34029 ; n34030
g33775 and n33934_not n34030_not ; n34031
g33776 and n34028_not n34031 ; n34032
g33777 and n33934_not n34032_not ; n34033
g33778 and b[9] n33923_not ; n34034
g33779 and n33921_not n34034 ; n34035
g33780 and n33925_not n34035_not ; n34036
g33781 and n34033_not n34036 ; n34037
g33782 and n33925_not n34037_not ; n34038
g33783 and b[10] n33914_not ; n34039
g33784 and n33912_not n34039 ; n34040
g33785 and n33916_not n34040_not ; n34041
g33786 and n34038_not n34041 ; n34042
g33787 and n33916_not n34042_not ; n34043
g33788 and b[11] n33905_not ; n34044
g33789 and n33903_not n34044 ; n34045
g33790 and n33907_not n34045_not ; n34046
g33791 and n34043_not n34046 ; n34047
g33792 and n33907_not n34047_not ; n34048
g33793 and b[12] n33896_not ; n34049
g33794 and n33894_not n34049 ; n34050
g33795 and n33898_not n34050_not ; n34051
g33796 and n34048_not n34051 ; n34052
g33797 and n33898_not n34052_not ; n34053
g33798 and b[13] n33887_not ; n34054
g33799 and n33885_not n34054 ; n34055
g33800 and n33889_not n34055_not ; n34056
g33801 and n34053_not n34056 ; n34057
g33802 and n33889_not n34057_not ; n34058
g33803 and b[14] n33878_not ; n34059
g33804 and n33876_not n34059 ; n34060
g33805 and n33880_not n34060_not ; n34061
g33806 and n34058_not n34061 ; n34062
g33807 and n33880_not n34062_not ; n34063
g33808 and b[15] n33869_not ; n34064
g33809 and n33867_not n34064 ; n34065
g33810 and n33871_not n34065_not ; n34066
g33811 and n34063_not n34066 ; n34067
g33812 and n33871_not n34067_not ; n34068
g33813 and b[16] n33860_not ; n34069
g33814 and n33858_not n34069 ; n34070
g33815 and n33862_not n34070_not ; n34071
g33816 and n34068_not n34071 ; n34072
g33817 and n33862_not n34072_not ; n34073
g33818 and b[17] n33851_not ; n34074
g33819 and n33849_not n34074 ; n34075
g33820 and n33853_not n34075_not ; n34076
g33821 and n34073_not n34076 ; n34077
g33822 and n33853_not n34077_not ; n34078
g33823 and b[18] n33842_not ; n34079
g33824 and n33840_not n34079 ; n34080
g33825 and n33844_not n34080_not ; n34081
g33826 and n34078_not n34081 ; n34082
g33827 and n33844_not n34082_not ; n34083
g33828 and b[19] n33833_not ; n34084
g33829 and n33831_not n34084 ; n34085
g33830 and n33835_not n34085_not ; n34086
g33831 and n34083_not n34086 ; n34087
g33832 and n33835_not n34087_not ; n34088
g33833 and b[20] n33824_not ; n34089
g33834 and n33822_not n34089 ; n34090
g33835 and n33826_not n34090_not ; n34091
g33836 and n34088_not n34091 ; n34092
g33837 and n33826_not n34092_not ; n34093
g33838 and b[21] n33815_not ; n34094
g33839 and n33813_not n34094 ; n34095
g33840 and n33817_not n34095_not ; n34096
g33841 and n34093_not n34096 ; n34097
g33842 and n33817_not n34097_not ; n34098
g33843 and b[22] n33806_not ; n34099
g33844 and n33804_not n34099 ; n34100
g33845 and n33808_not n34100_not ; n34101
g33846 and n34098_not n34101 ; n34102
g33847 and n33808_not n34102_not ; n34103
g33848 and b[23] n33797_not ; n34104
g33849 and n33795_not n34104 ; n34105
g33850 and n33799_not n34105_not ; n34106
g33851 and n34103_not n34106 ; n34107
g33852 and n33799_not n34107_not ; n34108
g33853 and b[24] n33788_not ; n34109
g33854 and n33786_not n34109 ; n34110
g33855 and n33790_not n34110_not ; n34111
g33856 and n34108_not n34111 ; n34112
g33857 and n33790_not n34112_not ; n34113
g33858 and b[25] n33779_not ; n34114
g33859 and n33777_not n34114 ; n34115
g33860 and n33781_not n34115_not ; n34116
g33861 and n34113_not n34116 ; n34117
g33862 and n33781_not n34117_not ; n34118
g33863 and b[26] n33759_not ; n34119
g33864 and n33757_not n34119 ; n34120
g33865 and n33772_not n34120_not ; n34121
g33866 and n34118_not n34121 ; n34122
g33867 and n33772_not n34122_not ; n34123
g33868 and b[27] n33769_not ; n34124
g33869 and n33767_not n34124 ; n34125
g33870 and n33771_not n34125_not ; n34126
g33871 and n34123_not n34126 ; n34127
g33872 and n33771_not n34127_not ; n34128
g33873 and n5926 n34128_not ; n34129
g33874 and n33760_not n34129_not ; n34130
g33875 and n33781_not n34121 ; n34131
g33876 and n34117_not n34131 ; n34132
g33877 and n34118_not n34121_not ; n34133
g33878 and n34132_not n34133_not ; n34134
g33879 and n5926 n34134_not ; n34135
g33880 and n34128_not n34135 ; n34136
g33881 and n34130_not n34136_not ; n34137
g33882 and n33770_not n34129_not ; n34138
g33883 and n33772_not n34126 ; n34139
g33884 and n34122_not n34139 ; n34140
g33885 and n34123_not n34126_not ; n34141
g33886 and n34140_not n34141_not ; n34142
g33887 and n34129 n34142_not ; n34143
g33888 and n34138_not n34143_not ; n34144
g33889 and b[28]_not n34144_not ; n34145
g33890 and b[27]_not n34137_not ; n34146
g33891 and n33780_not n34129_not ; n34147
g33892 and n33790_not n34116 ; n34148
g33893 and n34112_not n34148 ; n34149
g33894 and n34113_not n34116_not ; n34150
g33895 and n34149_not n34150_not ; n34151
g33896 and n5926 n34151_not ; n34152
g33897 and n34128_not n34152 ; n34153
g33898 and n34147_not n34153_not ; n34154
g33899 and b[26]_not n34154_not ; n34155
g33900 and n33789_not n34129_not ; n34156
g33901 and n33799_not n34111 ; n34157
g33902 and n34107_not n34157 ; n34158
g33903 and n34108_not n34111_not ; n34159
g33904 and n34158_not n34159_not ; n34160
g33905 and n5926 n34160_not ; n34161
g33906 and n34128_not n34161 ; n34162
g33907 and n34156_not n34162_not ; n34163
g33908 and b[25]_not n34163_not ; n34164
g33909 and n33798_not n34129_not ; n34165
g33910 and n33808_not n34106 ; n34166
g33911 and n34102_not n34166 ; n34167
g33912 and n34103_not n34106_not ; n34168
g33913 and n34167_not n34168_not ; n34169
g33914 and n5926 n34169_not ; n34170
g33915 and n34128_not n34170 ; n34171
g33916 and n34165_not n34171_not ; n34172
g33917 and b[24]_not n34172_not ; n34173
g33918 and n33807_not n34129_not ; n34174
g33919 and n33817_not n34101 ; n34175
g33920 and n34097_not n34175 ; n34176
g33921 and n34098_not n34101_not ; n34177
g33922 and n34176_not n34177_not ; n34178
g33923 and n5926 n34178_not ; n34179
g33924 and n34128_not n34179 ; n34180
g33925 and n34174_not n34180_not ; n34181
g33926 and b[23]_not n34181_not ; n34182
g33927 and n33816_not n34129_not ; n34183
g33928 and n33826_not n34096 ; n34184
g33929 and n34092_not n34184 ; n34185
g33930 and n34093_not n34096_not ; n34186
g33931 and n34185_not n34186_not ; n34187
g33932 and n5926 n34187_not ; n34188
g33933 and n34128_not n34188 ; n34189
g33934 and n34183_not n34189_not ; n34190
g33935 and b[22]_not n34190_not ; n34191
g33936 and n33825_not n34129_not ; n34192
g33937 and n33835_not n34091 ; n34193
g33938 and n34087_not n34193 ; n34194
g33939 and n34088_not n34091_not ; n34195
g33940 and n34194_not n34195_not ; n34196
g33941 and n5926 n34196_not ; n34197
g33942 and n34128_not n34197 ; n34198
g33943 and n34192_not n34198_not ; n34199
g33944 and b[21]_not n34199_not ; n34200
g33945 and n33834_not n34129_not ; n34201
g33946 and n33844_not n34086 ; n34202
g33947 and n34082_not n34202 ; n34203
g33948 and n34083_not n34086_not ; n34204
g33949 and n34203_not n34204_not ; n34205
g33950 and n5926 n34205_not ; n34206
g33951 and n34128_not n34206 ; n34207
g33952 and n34201_not n34207_not ; n34208
g33953 and b[20]_not n34208_not ; n34209
g33954 and n33843_not n34129_not ; n34210
g33955 and n33853_not n34081 ; n34211
g33956 and n34077_not n34211 ; n34212
g33957 and n34078_not n34081_not ; n34213
g33958 and n34212_not n34213_not ; n34214
g33959 and n5926 n34214_not ; n34215
g33960 and n34128_not n34215 ; n34216
g33961 and n34210_not n34216_not ; n34217
g33962 and b[19]_not n34217_not ; n34218
g33963 and n33852_not n34129_not ; n34219
g33964 and n33862_not n34076 ; n34220
g33965 and n34072_not n34220 ; n34221
g33966 and n34073_not n34076_not ; n34222
g33967 and n34221_not n34222_not ; n34223
g33968 and n5926 n34223_not ; n34224
g33969 and n34128_not n34224 ; n34225
g33970 and n34219_not n34225_not ; n34226
g33971 and b[18]_not n34226_not ; n34227
g33972 and n33861_not n34129_not ; n34228
g33973 and n33871_not n34071 ; n34229
g33974 and n34067_not n34229 ; n34230
g33975 and n34068_not n34071_not ; n34231
g33976 and n34230_not n34231_not ; n34232
g33977 and n5926 n34232_not ; n34233
g33978 and n34128_not n34233 ; n34234
g33979 and n34228_not n34234_not ; n34235
g33980 and b[17]_not n34235_not ; n34236
g33981 and n33870_not n34129_not ; n34237
g33982 and n33880_not n34066 ; n34238
g33983 and n34062_not n34238 ; n34239
g33984 and n34063_not n34066_not ; n34240
g33985 and n34239_not n34240_not ; n34241
g33986 and n5926 n34241_not ; n34242
g33987 and n34128_not n34242 ; n34243
g33988 and n34237_not n34243_not ; n34244
g33989 and b[16]_not n34244_not ; n34245
g33990 and n33879_not n34129_not ; n34246
g33991 and n33889_not n34061 ; n34247
g33992 and n34057_not n34247 ; n34248
g33993 and n34058_not n34061_not ; n34249
g33994 and n34248_not n34249_not ; n34250
g33995 and n5926 n34250_not ; n34251
g33996 and n34128_not n34251 ; n34252
g33997 and n34246_not n34252_not ; n34253
g33998 and b[15]_not n34253_not ; n34254
g33999 and n33888_not n34129_not ; n34255
g34000 and n33898_not n34056 ; n34256
g34001 and n34052_not n34256 ; n34257
g34002 and n34053_not n34056_not ; n34258
g34003 and n34257_not n34258_not ; n34259
g34004 and n5926 n34259_not ; n34260
g34005 and n34128_not n34260 ; n34261
g34006 and n34255_not n34261_not ; n34262
g34007 and b[14]_not n34262_not ; n34263
g34008 and n33897_not n34129_not ; n34264
g34009 and n33907_not n34051 ; n34265
g34010 and n34047_not n34265 ; n34266
g34011 and n34048_not n34051_not ; n34267
g34012 and n34266_not n34267_not ; n34268
g34013 and n5926 n34268_not ; n34269
g34014 and n34128_not n34269 ; n34270
g34015 and n34264_not n34270_not ; n34271
g34016 and b[13]_not n34271_not ; n34272
g34017 and n33906_not n34129_not ; n34273
g34018 and n33916_not n34046 ; n34274
g34019 and n34042_not n34274 ; n34275
g34020 and n34043_not n34046_not ; n34276
g34021 and n34275_not n34276_not ; n34277
g34022 and n5926 n34277_not ; n34278
g34023 and n34128_not n34278 ; n34279
g34024 and n34273_not n34279_not ; n34280
g34025 and b[12]_not n34280_not ; n34281
g34026 and n33915_not n34129_not ; n34282
g34027 and n33925_not n34041 ; n34283
g34028 and n34037_not n34283 ; n34284
g34029 and n34038_not n34041_not ; n34285
g34030 and n34284_not n34285_not ; n34286
g34031 and n5926 n34286_not ; n34287
g34032 and n34128_not n34287 ; n34288
g34033 and n34282_not n34288_not ; n34289
g34034 and b[11]_not n34289_not ; n34290
g34035 and n33924_not n34129_not ; n34291
g34036 and n33934_not n34036 ; n34292
g34037 and n34032_not n34292 ; n34293
g34038 and n34033_not n34036_not ; n34294
g34039 and n34293_not n34294_not ; n34295
g34040 and n5926 n34295_not ; n34296
g34041 and n34128_not n34296 ; n34297
g34042 and n34291_not n34297_not ; n34298
g34043 and b[10]_not n34298_not ; n34299
g34044 and n33933_not n34129_not ; n34300
g34045 and n33943_not n34031 ; n34301
g34046 and n34027_not n34301 ; n34302
g34047 and n34028_not n34031_not ; n34303
g34048 and n34302_not n34303_not ; n34304
g34049 and n5926 n34304_not ; n34305
g34050 and n34128_not n34305 ; n34306
g34051 and n34300_not n34306_not ; n34307
g34052 and b[9]_not n34307_not ; n34308
g34053 and n33942_not n34129_not ; n34309
g34054 and n33952_not n34026 ; n34310
g34055 and n34022_not n34310 ; n34311
g34056 and n34023_not n34026_not ; n34312
g34057 and n34311_not n34312_not ; n34313
g34058 and n5926 n34313_not ; n34314
g34059 and n34128_not n34314 ; n34315
g34060 and n34309_not n34315_not ; n34316
g34061 and b[8]_not n34316_not ; n34317
g34062 and n33951_not n34129_not ; n34318
g34063 and n33961_not n34021 ; n34319
g34064 and n34017_not n34319 ; n34320
g34065 and n34018_not n34021_not ; n34321
g34066 and n34320_not n34321_not ; n34322
g34067 and n5926 n34322_not ; n34323
g34068 and n34128_not n34323 ; n34324
g34069 and n34318_not n34324_not ; n34325
g34070 and b[7]_not n34325_not ; n34326
g34071 and n33960_not n34129_not ; n34327
g34072 and n33970_not n34016 ; n34328
g34073 and n34012_not n34328 ; n34329
g34074 and n34013_not n34016_not ; n34330
g34075 and n34329_not n34330_not ; n34331
g34076 and n5926 n34331_not ; n34332
g34077 and n34128_not n34332 ; n34333
g34078 and n34327_not n34333_not ; n34334
g34079 and b[6]_not n34334_not ; n34335
g34080 and n33969_not n34129_not ; n34336
g34081 and n33979_not n34011 ; n34337
g34082 and n34007_not n34337 ; n34338
g34083 and n34008_not n34011_not ; n34339
g34084 and n34338_not n34339_not ; n34340
g34085 and n5926 n34340_not ; n34341
g34086 and n34128_not n34341 ; n34342
g34087 and n34336_not n34342_not ; n34343
g34088 and b[5]_not n34343_not ; n34344
g34089 and n33978_not n34129_not ; n34345
g34090 and n33987_not n34006 ; n34346
g34091 and n34002_not n34346 ; n34347
g34092 and n34003_not n34006_not ; n34348
g34093 and n34347_not n34348_not ; n34349
g34094 and n5926 n34349_not ; n34350
g34095 and n34128_not n34350 ; n34351
g34096 and n34345_not n34351_not ; n34352
g34097 and b[4]_not n34352_not ; n34353
g34098 and n33986_not n34129_not ; n34354
g34099 and n33997_not n34001 ; n34355
g34100 and n33996_not n34355 ; n34356
g34101 and n33998_not n34001_not ; n34357
g34102 and n34356_not n34357_not ; n34358
g34103 and n5926 n34358_not ; n34359
g34104 and n34128_not n34359 ; n34360
g34105 and n34354_not n34360_not ; n34361
g34106 and b[3]_not n34361_not ; n34362
g34107 and n33991_not n34129_not ; n34363
g34108 and n5791 n33994_not ; n34364
g34109 and n33992_not n34364 ; n34365
g34110 and n5926 n34365_not ; n34366
g34111 and n33996_not n34366 ; n34367
g34112 and n34128_not n34367 ; n34368
g34113 and n34363_not n34368_not ; n34369
g34114 and b[2]_not n34369_not ; n34370
g34115 and n6172 n34128_not ; n34371
g34116 and a[36] n34371_not ; n34372
g34117 and n6177 n34128_not ; n34373
g34118 and n34372_not n34373_not ; n34374
g34119 and b[1] n34374_not ; n34375
g34120 and b[1]_not n34373_not ; n34376
g34121 and n34372_not n34376 ; n34377
g34122 and n34375_not n34377_not ; n34378
g34123 and n6184_not n34378_not ; n34379
g34124 and b[1]_not n34374_not ; n34380
g34125 and n34379_not n34380_not ; n34381
g34126 and b[2] n34368_not ; n34382
g34127 and n34363_not n34382 ; n34383
g34128 and n34370_not n34383_not ; n34384
g34129 and n34381_not n34384 ; n34385
g34130 and n34370_not n34385_not ; n34386
g34131 and b[3] n34360_not ; n34387
g34132 and n34354_not n34387 ; n34388
g34133 and n34362_not n34388_not ; n34389
g34134 and n34386_not n34389 ; n34390
g34135 and n34362_not n34390_not ; n34391
g34136 and b[4] n34351_not ; n34392
g34137 and n34345_not n34392 ; n34393
g34138 and n34353_not n34393_not ; n34394
g34139 and n34391_not n34394 ; n34395
g34140 and n34353_not n34395_not ; n34396
g34141 and b[5] n34342_not ; n34397
g34142 and n34336_not n34397 ; n34398
g34143 and n34344_not n34398_not ; n34399
g34144 and n34396_not n34399 ; n34400
g34145 and n34344_not n34400_not ; n34401
g34146 and b[6] n34333_not ; n34402
g34147 and n34327_not n34402 ; n34403
g34148 and n34335_not n34403_not ; n34404
g34149 and n34401_not n34404 ; n34405
g34150 and n34335_not n34405_not ; n34406
g34151 and b[7] n34324_not ; n34407
g34152 and n34318_not n34407 ; n34408
g34153 and n34326_not n34408_not ; n34409
g34154 and n34406_not n34409 ; n34410
g34155 and n34326_not n34410_not ; n34411
g34156 and b[8] n34315_not ; n34412
g34157 and n34309_not n34412 ; n34413
g34158 and n34317_not n34413_not ; n34414
g34159 and n34411_not n34414 ; n34415
g34160 and n34317_not n34415_not ; n34416
g34161 and b[9] n34306_not ; n34417
g34162 and n34300_not n34417 ; n34418
g34163 and n34308_not n34418_not ; n34419
g34164 and n34416_not n34419 ; n34420
g34165 and n34308_not n34420_not ; n34421
g34166 and b[10] n34297_not ; n34422
g34167 and n34291_not n34422 ; n34423
g34168 and n34299_not n34423_not ; n34424
g34169 and n34421_not n34424 ; n34425
g34170 and n34299_not n34425_not ; n34426
g34171 and b[11] n34288_not ; n34427
g34172 and n34282_not n34427 ; n34428
g34173 and n34290_not n34428_not ; n34429
g34174 and n34426_not n34429 ; n34430
g34175 and n34290_not n34430_not ; n34431
g34176 and b[12] n34279_not ; n34432
g34177 and n34273_not n34432 ; n34433
g34178 and n34281_not n34433_not ; n34434
g34179 and n34431_not n34434 ; n34435
g34180 and n34281_not n34435_not ; n34436
g34181 and b[13] n34270_not ; n34437
g34182 and n34264_not n34437 ; n34438
g34183 and n34272_not n34438_not ; n34439
g34184 and n34436_not n34439 ; n34440
g34185 and n34272_not n34440_not ; n34441
g34186 and b[14] n34261_not ; n34442
g34187 and n34255_not n34442 ; n34443
g34188 and n34263_not n34443_not ; n34444
g34189 and n34441_not n34444 ; n34445
g34190 and n34263_not n34445_not ; n34446
g34191 and b[15] n34252_not ; n34447
g34192 and n34246_not n34447 ; n34448
g34193 and n34254_not n34448_not ; n34449
g34194 and n34446_not n34449 ; n34450
g34195 and n34254_not n34450_not ; n34451
g34196 and b[16] n34243_not ; n34452
g34197 and n34237_not n34452 ; n34453
g34198 and n34245_not n34453_not ; n34454
g34199 and n34451_not n34454 ; n34455
g34200 and n34245_not n34455_not ; n34456
g34201 and b[17] n34234_not ; n34457
g34202 and n34228_not n34457 ; n34458
g34203 and n34236_not n34458_not ; n34459
g34204 and n34456_not n34459 ; n34460
g34205 and n34236_not n34460_not ; n34461
g34206 and b[18] n34225_not ; n34462
g34207 and n34219_not n34462 ; n34463
g34208 and n34227_not n34463_not ; n34464
g34209 and n34461_not n34464 ; n34465
g34210 and n34227_not n34465_not ; n34466
g34211 and b[19] n34216_not ; n34467
g34212 and n34210_not n34467 ; n34468
g34213 and n34218_not n34468_not ; n34469
g34214 and n34466_not n34469 ; n34470
g34215 and n34218_not n34470_not ; n34471
g34216 and b[20] n34207_not ; n34472
g34217 and n34201_not n34472 ; n34473
g34218 and n34209_not n34473_not ; n34474
g34219 and n34471_not n34474 ; n34475
g34220 and n34209_not n34475_not ; n34476
g34221 and b[21] n34198_not ; n34477
g34222 and n34192_not n34477 ; n34478
g34223 and n34200_not n34478_not ; n34479
g34224 and n34476_not n34479 ; n34480
g34225 and n34200_not n34480_not ; n34481
g34226 and b[22] n34189_not ; n34482
g34227 and n34183_not n34482 ; n34483
g34228 and n34191_not n34483_not ; n34484
g34229 and n34481_not n34484 ; n34485
g34230 and n34191_not n34485_not ; n34486
g34231 and b[23] n34180_not ; n34487
g34232 and n34174_not n34487 ; n34488
g34233 and n34182_not n34488_not ; n34489
g34234 and n34486_not n34489 ; n34490
g34235 and n34182_not n34490_not ; n34491
g34236 and b[24] n34171_not ; n34492
g34237 and n34165_not n34492 ; n34493
g34238 and n34173_not n34493_not ; n34494
g34239 and n34491_not n34494 ; n34495
g34240 and n34173_not n34495_not ; n34496
g34241 and b[25] n34162_not ; n34497
g34242 and n34156_not n34497 ; n34498
g34243 and n34164_not n34498_not ; n34499
g34244 and n34496_not n34499 ; n34500
g34245 and n34164_not n34500_not ; n34501
g34246 and b[26] n34153_not ; n34502
g34247 and n34147_not n34502 ; n34503
g34248 and n34155_not n34503_not ; n34504
g34249 and n34501_not n34504 ; n34505
g34250 and n34155_not n34505_not ; n34506
g34251 and b[27] n34136_not ; n34507
g34252 and n34130_not n34507 ; n34508
g34253 and n34146_not n34508_not ; n34509
g34254 and n34506_not n34509 ; n34510
g34255 and n34146_not n34510_not ; n34511
g34256 and b[28] n34138_not ; n34512
g34257 and n34143_not n34512 ; n34513
g34258 and n34145_not n34513_not ; n34514
g34259 and n34511_not n34514 ; n34515
g34260 and n34145_not n34515_not ; n34516
g34261 and n6324 n34516_not ; n34517
g34262 and n34137_not n34517_not ; n34518
g34263 and n34155_not n34509 ; n34519
g34264 and n34505_not n34519 ; n34520
g34265 and n34506_not n34509_not ; n34521
g34266 and n34520_not n34521_not ; n34522
g34267 and n6324 n34522_not ; n34523
g34268 and n34516_not n34523 ; n34524
g34269 and n34518_not n34524_not ; n34525
g34270 and b[28]_not n34525_not ; n34526
g34271 and n34154_not n34517_not ; n34527
g34272 and n34164_not n34504 ; n34528
g34273 and n34500_not n34528 ; n34529
g34274 and n34501_not n34504_not ; n34530
g34275 and n34529_not n34530_not ; n34531
g34276 and n6324 n34531_not ; n34532
g34277 and n34516_not n34532 ; n34533
g34278 and n34527_not n34533_not ; n34534
g34279 and b[27]_not n34534_not ; n34535
g34280 and n34163_not n34517_not ; n34536
g34281 and n34173_not n34499 ; n34537
g34282 and n34495_not n34537 ; n34538
g34283 and n34496_not n34499_not ; n34539
g34284 and n34538_not n34539_not ; n34540
g34285 and n6324 n34540_not ; n34541
g34286 and n34516_not n34541 ; n34542
g34287 and n34536_not n34542_not ; n34543
g34288 and b[26]_not n34543_not ; n34544
g34289 and n34172_not n34517_not ; n34545
g34290 and n34182_not n34494 ; n34546
g34291 and n34490_not n34546 ; n34547
g34292 and n34491_not n34494_not ; n34548
g34293 and n34547_not n34548_not ; n34549
g34294 and n6324 n34549_not ; n34550
g34295 and n34516_not n34550 ; n34551
g34296 and n34545_not n34551_not ; n34552
g34297 and b[25]_not n34552_not ; n34553
g34298 and n34181_not n34517_not ; n34554
g34299 and n34191_not n34489 ; n34555
g34300 and n34485_not n34555 ; n34556
g34301 and n34486_not n34489_not ; n34557
g34302 and n34556_not n34557_not ; n34558
g34303 and n6324 n34558_not ; n34559
g34304 and n34516_not n34559 ; n34560
g34305 and n34554_not n34560_not ; n34561
g34306 and b[24]_not n34561_not ; n34562
g34307 and n34190_not n34517_not ; n34563
g34308 and n34200_not n34484 ; n34564
g34309 and n34480_not n34564 ; n34565
g34310 and n34481_not n34484_not ; n34566
g34311 and n34565_not n34566_not ; n34567
g34312 and n6324 n34567_not ; n34568
g34313 and n34516_not n34568 ; n34569
g34314 and n34563_not n34569_not ; n34570
g34315 and b[23]_not n34570_not ; n34571
g34316 and n34199_not n34517_not ; n34572
g34317 and n34209_not n34479 ; n34573
g34318 and n34475_not n34573 ; n34574
g34319 and n34476_not n34479_not ; n34575
g34320 and n34574_not n34575_not ; n34576
g34321 and n6324 n34576_not ; n34577
g34322 and n34516_not n34577 ; n34578
g34323 and n34572_not n34578_not ; n34579
g34324 and b[22]_not n34579_not ; n34580
g34325 and n34208_not n34517_not ; n34581
g34326 and n34218_not n34474 ; n34582
g34327 and n34470_not n34582 ; n34583
g34328 and n34471_not n34474_not ; n34584
g34329 and n34583_not n34584_not ; n34585
g34330 and n6324 n34585_not ; n34586
g34331 and n34516_not n34586 ; n34587
g34332 and n34581_not n34587_not ; n34588
g34333 and b[21]_not n34588_not ; n34589
g34334 and n34217_not n34517_not ; n34590
g34335 and n34227_not n34469 ; n34591
g34336 and n34465_not n34591 ; n34592
g34337 and n34466_not n34469_not ; n34593
g34338 and n34592_not n34593_not ; n34594
g34339 and n6324 n34594_not ; n34595
g34340 and n34516_not n34595 ; n34596
g34341 and n34590_not n34596_not ; n34597
g34342 and b[20]_not n34597_not ; n34598
g34343 and n34226_not n34517_not ; n34599
g34344 and n34236_not n34464 ; n34600
g34345 and n34460_not n34600 ; n34601
g34346 and n34461_not n34464_not ; n34602
g34347 and n34601_not n34602_not ; n34603
g34348 and n6324 n34603_not ; n34604
g34349 and n34516_not n34604 ; n34605
g34350 and n34599_not n34605_not ; n34606
g34351 and b[19]_not n34606_not ; n34607
g34352 and n34235_not n34517_not ; n34608
g34353 and n34245_not n34459 ; n34609
g34354 and n34455_not n34609 ; n34610
g34355 and n34456_not n34459_not ; n34611
g34356 and n34610_not n34611_not ; n34612
g34357 and n6324 n34612_not ; n34613
g34358 and n34516_not n34613 ; n34614
g34359 and n34608_not n34614_not ; n34615
g34360 and b[18]_not n34615_not ; n34616
g34361 and n34244_not n34517_not ; n34617
g34362 and n34254_not n34454 ; n34618
g34363 and n34450_not n34618 ; n34619
g34364 and n34451_not n34454_not ; n34620
g34365 and n34619_not n34620_not ; n34621
g34366 and n6324 n34621_not ; n34622
g34367 and n34516_not n34622 ; n34623
g34368 and n34617_not n34623_not ; n34624
g34369 and b[17]_not n34624_not ; n34625
g34370 and n34253_not n34517_not ; n34626
g34371 and n34263_not n34449 ; n34627
g34372 and n34445_not n34627 ; n34628
g34373 and n34446_not n34449_not ; n34629
g34374 and n34628_not n34629_not ; n34630
g34375 and n6324 n34630_not ; n34631
g34376 and n34516_not n34631 ; n34632
g34377 and n34626_not n34632_not ; n34633
g34378 and b[16]_not n34633_not ; n34634
g34379 and n34262_not n34517_not ; n34635
g34380 and n34272_not n34444 ; n34636
g34381 and n34440_not n34636 ; n34637
g34382 and n34441_not n34444_not ; n34638
g34383 and n34637_not n34638_not ; n34639
g34384 and n6324 n34639_not ; n34640
g34385 and n34516_not n34640 ; n34641
g34386 and n34635_not n34641_not ; n34642
g34387 and b[15]_not n34642_not ; n34643
g34388 and n34271_not n34517_not ; n34644
g34389 and n34281_not n34439 ; n34645
g34390 and n34435_not n34645 ; n34646
g34391 and n34436_not n34439_not ; n34647
g34392 and n34646_not n34647_not ; n34648
g34393 and n6324 n34648_not ; n34649
g34394 and n34516_not n34649 ; n34650
g34395 and n34644_not n34650_not ; n34651
g34396 and b[14]_not n34651_not ; n34652
g34397 and n34280_not n34517_not ; n34653
g34398 and n34290_not n34434 ; n34654
g34399 and n34430_not n34654 ; n34655
g34400 and n34431_not n34434_not ; n34656
g34401 and n34655_not n34656_not ; n34657
g34402 and n6324 n34657_not ; n34658
g34403 and n34516_not n34658 ; n34659
g34404 and n34653_not n34659_not ; n34660
g34405 and b[13]_not n34660_not ; n34661
g34406 and n34289_not n34517_not ; n34662
g34407 and n34299_not n34429 ; n34663
g34408 and n34425_not n34663 ; n34664
g34409 and n34426_not n34429_not ; n34665
g34410 and n34664_not n34665_not ; n34666
g34411 and n6324 n34666_not ; n34667
g34412 and n34516_not n34667 ; n34668
g34413 and n34662_not n34668_not ; n34669
g34414 and b[12]_not n34669_not ; n34670
g34415 and n34298_not n34517_not ; n34671
g34416 and n34308_not n34424 ; n34672
g34417 and n34420_not n34672 ; n34673
g34418 and n34421_not n34424_not ; n34674
g34419 and n34673_not n34674_not ; n34675
g34420 and n6324 n34675_not ; n34676
g34421 and n34516_not n34676 ; n34677
g34422 and n34671_not n34677_not ; n34678
g34423 and b[11]_not n34678_not ; n34679
g34424 and n34307_not n34517_not ; n34680
g34425 and n34317_not n34419 ; n34681
g34426 and n34415_not n34681 ; n34682
g34427 and n34416_not n34419_not ; n34683
g34428 and n34682_not n34683_not ; n34684
g34429 and n6324 n34684_not ; n34685
g34430 and n34516_not n34685 ; n34686
g34431 and n34680_not n34686_not ; n34687
g34432 and b[10]_not n34687_not ; n34688
g34433 and n34316_not n34517_not ; n34689
g34434 and n34326_not n34414 ; n34690
g34435 and n34410_not n34690 ; n34691
g34436 and n34411_not n34414_not ; n34692
g34437 and n34691_not n34692_not ; n34693
g34438 and n6324 n34693_not ; n34694
g34439 and n34516_not n34694 ; n34695
g34440 and n34689_not n34695_not ; n34696
g34441 and b[9]_not n34696_not ; n34697
g34442 and n34325_not n34517_not ; n34698
g34443 and n34335_not n34409 ; n34699
g34444 and n34405_not n34699 ; n34700
g34445 and n34406_not n34409_not ; n34701
g34446 and n34700_not n34701_not ; n34702
g34447 and n6324 n34702_not ; n34703
g34448 and n34516_not n34703 ; n34704
g34449 and n34698_not n34704_not ; n34705
g34450 and b[8]_not n34705_not ; n34706
g34451 and n34334_not n34517_not ; n34707
g34452 and n34344_not n34404 ; n34708
g34453 and n34400_not n34708 ; n34709
g34454 and n34401_not n34404_not ; n34710
g34455 and n34709_not n34710_not ; n34711
g34456 and n6324 n34711_not ; n34712
g34457 and n34516_not n34712 ; n34713
g34458 and n34707_not n34713_not ; n34714
g34459 and b[7]_not n34714_not ; n34715
g34460 and n34343_not n34517_not ; n34716
g34461 and n34353_not n34399 ; n34717
g34462 and n34395_not n34717 ; n34718
g34463 and n34396_not n34399_not ; n34719
g34464 and n34718_not n34719_not ; n34720
g34465 and n6324 n34720_not ; n34721
g34466 and n34516_not n34721 ; n34722
g34467 and n34716_not n34722_not ; n34723
g34468 and b[6]_not n34723_not ; n34724
g34469 and n34352_not n34517_not ; n34725
g34470 and n34362_not n34394 ; n34726
g34471 and n34390_not n34726 ; n34727
g34472 and n34391_not n34394_not ; n34728
g34473 and n34727_not n34728_not ; n34729
g34474 and n6324 n34729_not ; n34730
g34475 and n34516_not n34730 ; n34731
g34476 and n34725_not n34731_not ; n34732
g34477 and b[5]_not n34732_not ; n34733
g34478 and n34361_not n34517_not ; n34734
g34479 and n34370_not n34389 ; n34735
g34480 and n34385_not n34735 ; n34736
g34481 and n34386_not n34389_not ; n34737
g34482 and n34736_not n34737_not ; n34738
g34483 and n6324 n34738_not ; n34739
g34484 and n34516_not n34739 ; n34740
g34485 and n34734_not n34740_not ; n34741
g34486 and b[4]_not n34741_not ; n34742
g34487 and n34369_not n34517_not ; n34743
g34488 and n34380_not n34384 ; n34744
g34489 and n34379_not n34744 ; n34745
g34490 and n34381_not n34384_not ; n34746
g34491 and n34745_not n34746_not ; n34747
g34492 and n6324 n34747_not ; n34748
g34493 and n34516_not n34748 ; n34749
g34494 and n34743_not n34749_not ; n34750
g34495 and b[3]_not n34750_not ; n34751
g34496 and n34374_not n34517_not ; n34752
g34497 and n6184 n34377_not ; n34753
g34498 and n34375_not n34753 ; n34754
g34499 and n6324 n34754_not ; n34755
g34500 and n34379_not n34755 ; n34756
g34501 and n34516_not n34756 ; n34757
g34502 and n34752_not n34757_not ; n34758
g34503 and b[2]_not n34758_not ; n34759
g34504 and n6572 n34516_not ; n34760
g34505 and a[35] n34760_not ; n34761
g34506 and n6577 n34516_not ; n34762
g34507 and n34761_not n34762_not ; n34763
g34508 and b[1] n34763_not ; n34764
g34509 and b[1]_not n34762_not ; n34765
g34510 and n34761_not n34765 ; n34766
g34511 and n34764_not n34766_not ; n34767
g34512 and n6584_not n34767_not ; n34768
g34513 and b[1]_not n34763_not ; n34769
g34514 and n34768_not n34769_not ; n34770
g34515 and b[2] n34757_not ; n34771
g34516 and n34752_not n34771 ; n34772
g34517 and n34759_not n34772_not ; n34773
g34518 and n34770_not n34773 ; n34774
g34519 and n34759_not n34774_not ; n34775
g34520 and b[3] n34749_not ; n34776
g34521 and n34743_not n34776 ; n34777
g34522 and n34751_not n34777_not ; n34778
g34523 and n34775_not n34778 ; n34779
g34524 and n34751_not n34779_not ; n34780
g34525 and b[4] n34740_not ; n34781
g34526 and n34734_not n34781 ; n34782
g34527 and n34742_not n34782_not ; n34783
g34528 and n34780_not n34783 ; n34784
g34529 and n34742_not n34784_not ; n34785
g34530 and b[5] n34731_not ; n34786
g34531 and n34725_not n34786 ; n34787
g34532 and n34733_not n34787_not ; n34788
g34533 and n34785_not n34788 ; n34789
g34534 and n34733_not n34789_not ; n34790
g34535 and b[6] n34722_not ; n34791
g34536 and n34716_not n34791 ; n34792
g34537 and n34724_not n34792_not ; n34793
g34538 and n34790_not n34793 ; n34794
g34539 and n34724_not n34794_not ; n34795
g34540 and b[7] n34713_not ; n34796
g34541 and n34707_not n34796 ; n34797
g34542 and n34715_not n34797_not ; n34798
g34543 and n34795_not n34798 ; n34799
g34544 and n34715_not n34799_not ; n34800
g34545 and b[8] n34704_not ; n34801
g34546 and n34698_not n34801 ; n34802
g34547 and n34706_not n34802_not ; n34803
g34548 and n34800_not n34803 ; n34804
g34549 and n34706_not n34804_not ; n34805
g34550 and b[9] n34695_not ; n34806
g34551 and n34689_not n34806 ; n34807
g34552 and n34697_not n34807_not ; n34808
g34553 and n34805_not n34808 ; n34809
g34554 and n34697_not n34809_not ; n34810
g34555 and b[10] n34686_not ; n34811
g34556 and n34680_not n34811 ; n34812
g34557 and n34688_not n34812_not ; n34813
g34558 and n34810_not n34813 ; n34814
g34559 and n34688_not n34814_not ; n34815
g34560 and b[11] n34677_not ; n34816
g34561 and n34671_not n34816 ; n34817
g34562 and n34679_not n34817_not ; n34818
g34563 and n34815_not n34818 ; n34819
g34564 and n34679_not n34819_not ; n34820
g34565 and b[12] n34668_not ; n34821
g34566 and n34662_not n34821 ; n34822
g34567 and n34670_not n34822_not ; n34823
g34568 and n34820_not n34823 ; n34824
g34569 and n34670_not n34824_not ; n34825
g34570 and b[13] n34659_not ; n34826
g34571 and n34653_not n34826 ; n34827
g34572 and n34661_not n34827_not ; n34828
g34573 and n34825_not n34828 ; n34829
g34574 and n34661_not n34829_not ; n34830
g34575 and b[14] n34650_not ; n34831
g34576 and n34644_not n34831 ; n34832
g34577 and n34652_not n34832_not ; n34833
g34578 and n34830_not n34833 ; n34834
g34579 and n34652_not n34834_not ; n34835
g34580 and b[15] n34641_not ; n34836
g34581 and n34635_not n34836 ; n34837
g34582 and n34643_not n34837_not ; n34838
g34583 and n34835_not n34838 ; n34839
g34584 and n34643_not n34839_not ; n34840
g34585 and b[16] n34632_not ; n34841
g34586 and n34626_not n34841 ; n34842
g34587 and n34634_not n34842_not ; n34843
g34588 and n34840_not n34843 ; n34844
g34589 and n34634_not n34844_not ; n34845
g34590 and b[17] n34623_not ; n34846
g34591 and n34617_not n34846 ; n34847
g34592 and n34625_not n34847_not ; n34848
g34593 and n34845_not n34848 ; n34849
g34594 and n34625_not n34849_not ; n34850
g34595 and b[18] n34614_not ; n34851
g34596 and n34608_not n34851 ; n34852
g34597 and n34616_not n34852_not ; n34853
g34598 and n34850_not n34853 ; n34854
g34599 and n34616_not n34854_not ; n34855
g34600 and b[19] n34605_not ; n34856
g34601 and n34599_not n34856 ; n34857
g34602 and n34607_not n34857_not ; n34858
g34603 and n34855_not n34858 ; n34859
g34604 and n34607_not n34859_not ; n34860
g34605 and b[20] n34596_not ; n34861
g34606 and n34590_not n34861 ; n34862
g34607 and n34598_not n34862_not ; n34863
g34608 and n34860_not n34863 ; n34864
g34609 and n34598_not n34864_not ; n34865
g34610 and b[21] n34587_not ; n34866
g34611 and n34581_not n34866 ; n34867
g34612 and n34589_not n34867_not ; n34868
g34613 and n34865_not n34868 ; n34869
g34614 and n34589_not n34869_not ; n34870
g34615 and b[22] n34578_not ; n34871
g34616 and n34572_not n34871 ; n34872
g34617 and n34580_not n34872_not ; n34873
g34618 and n34870_not n34873 ; n34874
g34619 and n34580_not n34874_not ; n34875
g34620 and b[23] n34569_not ; n34876
g34621 and n34563_not n34876 ; n34877
g34622 and n34571_not n34877_not ; n34878
g34623 and n34875_not n34878 ; n34879
g34624 and n34571_not n34879_not ; n34880
g34625 and b[24] n34560_not ; n34881
g34626 and n34554_not n34881 ; n34882
g34627 and n34562_not n34882_not ; n34883
g34628 and n34880_not n34883 ; n34884
g34629 and n34562_not n34884_not ; n34885
g34630 and b[25] n34551_not ; n34886
g34631 and n34545_not n34886 ; n34887
g34632 and n34553_not n34887_not ; n34888
g34633 and n34885_not n34888 ; n34889
g34634 and n34553_not n34889_not ; n34890
g34635 and b[26] n34542_not ; n34891
g34636 and n34536_not n34891 ; n34892
g34637 and n34544_not n34892_not ; n34893
g34638 and n34890_not n34893 ; n34894
g34639 and n34544_not n34894_not ; n34895
g34640 and b[27] n34533_not ; n34896
g34641 and n34527_not n34896 ; n34897
g34642 and n34535_not n34897_not ; n34898
g34643 and n34895_not n34898 ; n34899
g34644 and n34535_not n34899_not ; n34900
g34645 and b[28] n34524_not ; n34901
g34646 and n34518_not n34901 ; n34902
g34647 and n34526_not n34902_not ; n34903
g34648 and n34900_not n34903 ; n34904
g34649 and n34526_not n34904_not ; n34905
g34650 and n34144_not n34517_not ; n34906
g34651 and n34146_not n34514 ; n34907
g34652 and n34510_not n34907 ; n34908
g34653 and n34511_not n34514_not ; n34909
g34654 and n34908_not n34909_not ; n34910
g34655 and n34517 n34910_not ; n34911
g34656 and n34906_not n34911_not ; n34912
g34657 and b[29]_not n34912_not ; n34913
g34658 and b[29] n34906_not ; n34914
g34659 and n34911_not n34914 ; n34915
g34660 and n6735 n34915_not ; n34916
g34661 and n34913_not n34916 ; n34917
g34662 and n34905_not n34917 ; n34918
g34663 and n6324 n34912_not ; n34919
g34664 and n34918_not n34919_not ; n34920
g34665 and n34535_not n34903 ; n34921
g34666 and n34899_not n34921 ; n34922
g34667 and n34900_not n34903_not ; n34923
g34668 and n34922_not n34923_not ; n34924
g34669 and n34920_not n34924_not ; n34925
g34670 and n34525_not n34919_not ; n34926
g34671 and n34918_not n34926 ; n34927
g34672 and n34925_not n34927_not ; n34928
g34673 and n34526_not n34915_not ; n34929
g34674 and n34913_not n34929 ; n34930
g34675 and n34904_not n34930 ; n34931
g34676 and n34913_not n34915_not ; n34932
g34677 and n34905_not n34932_not ; n34933
g34678 and n34931_not n34933_not ; n34934
g34679 and n34920_not n34934_not ; n34935
g34680 and n34912_not n34919_not ; n34936
g34681 and n34918_not n34936 ; n34937
g34682 and n34935_not n34937_not ; n34938
g34683 and b[30]_not n34938_not ; n34939
g34684 and b[29]_not n34928_not ; n34940
g34685 and n34544_not n34898 ; n34941
g34686 and n34894_not n34941 ; n34942
g34687 and n34895_not n34898_not ; n34943
g34688 and n34942_not n34943_not ; n34944
g34689 and n34920_not n34944_not ; n34945
g34690 and n34534_not n34919_not ; n34946
g34691 and n34918_not n34946 ; n34947
g34692 and n34945_not n34947_not ; n34948
g34693 and b[28]_not n34948_not ; n34949
g34694 and n34553_not n34893 ; n34950
g34695 and n34889_not n34950 ; n34951
g34696 and n34890_not n34893_not ; n34952
g34697 and n34951_not n34952_not ; n34953
g34698 and n34920_not n34953_not ; n34954
g34699 and n34543_not n34919_not ; n34955
g34700 and n34918_not n34955 ; n34956
g34701 and n34954_not n34956_not ; n34957
g34702 and b[27]_not n34957_not ; n34958
g34703 and n34562_not n34888 ; n34959
g34704 and n34884_not n34959 ; n34960
g34705 and n34885_not n34888_not ; n34961
g34706 and n34960_not n34961_not ; n34962
g34707 and n34920_not n34962_not ; n34963
g34708 and n34552_not n34919_not ; n34964
g34709 and n34918_not n34964 ; n34965
g34710 and n34963_not n34965_not ; n34966
g34711 and b[26]_not n34966_not ; n34967
g34712 and n34571_not n34883 ; n34968
g34713 and n34879_not n34968 ; n34969
g34714 and n34880_not n34883_not ; n34970
g34715 and n34969_not n34970_not ; n34971
g34716 and n34920_not n34971_not ; n34972
g34717 and n34561_not n34919_not ; n34973
g34718 and n34918_not n34973 ; n34974
g34719 and n34972_not n34974_not ; n34975
g34720 and b[25]_not n34975_not ; n34976
g34721 and n34580_not n34878 ; n34977
g34722 and n34874_not n34977 ; n34978
g34723 and n34875_not n34878_not ; n34979
g34724 and n34978_not n34979_not ; n34980
g34725 and n34920_not n34980_not ; n34981
g34726 and n34570_not n34919_not ; n34982
g34727 and n34918_not n34982 ; n34983
g34728 and n34981_not n34983_not ; n34984
g34729 and b[24]_not n34984_not ; n34985
g34730 and n34589_not n34873 ; n34986
g34731 and n34869_not n34986 ; n34987
g34732 and n34870_not n34873_not ; n34988
g34733 and n34987_not n34988_not ; n34989
g34734 and n34920_not n34989_not ; n34990
g34735 and n34579_not n34919_not ; n34991
g34736 and n34918_not n34991 ; n34992
g34737 and n34990_not n34992_not ; n34993
g34738 and b[23]_not n34993_not ; n34994
g34739 and n34598_not n34868 ; n34995
g34740 and n34864_not n34995 ; n34996
g34741 and n34865_not n34868_not ; n34997
g34742 and n34996_not n34997_not ; n34998
g34743 and n34920_not n34998_not ; n34999
g34744 and n34588_not n34919_not ; n35000
g34745 and n34918_not n35000 ; n35001
g34746 and n34999_not n35001_not ; n35002
g34747 and b[22]_not n35002_not ; n35003
g34748 and n34607_not n34863 ; n35004
g34749 and n34859_not n35004 ; n35005
g34750 and n34860_not n34863_not ; n35006
g34751 and n35005_not n35006_not ; n35007
g34752 and n34920_not n35007_not ; n35008
g34753 and n34597_not n34919_not ; n35009
g34754 and n34918_not n35009 ; n35010
g34755 and n35008_not n35010_not ; n35011
g34756 and b[21]_not n35011_not ; n35012
g34757 and n34616_not n34858 ; n35013
g34758 and n34854_not n35013 ; n35014
g34759 and n34855_not n34858_not ; n35015
g34760 and n35014_not n35015_not ; n35016
g34761 and n34920_not n35016_not ; n35017
g34762 and n34606_not n34919_not ; n35018
g34763 and n34918_not n35018 ; n35019
g34764 and n35017_not n35019_not ; n35020
g34765 and b[20]_not n35020_not ; n35021
g34766 and n34625_not n34853 ; n35022
g34767 and n34849_not n35022 ; n35023
g34768 and n34850_not n34853_not ; n35024
g34769 and n35023_not n35024_not ; n35025
g34770 and n34920_not n35025_not ; n35026
g34771 and n34615_not n34919_not ; n35027
g34772 and n34918_not n35027 ; n35028
g34773 and n35026_not n35028_not ; n35029
g34774 and b[19]_not n35029_not ; n35030
g34775 and n34634_not n34848 ; n35031
g34776 and n34844_not n35031 ; n35032
g34777 and n34845_not n34848_not ; n35033
g34778 and n35032_not n35033_not ; n35034
g34779 and n34920_not n35034_not ; n35035
g34780 and n34624_not n34919_not ; n35036
g34781 and n34918_not n35036 ; n35037
g34782 and n35035_not n35037_not ; n35038
g34783 and b[18]_not n35038_not ; n35039
g34784 and n34643_not n34843 ; n35040
g34785 and n34839_not n35040 ; n35041
g34786 and n34840_not n34843_not ; n35042
g34787 and n35041_not n35042_not ; n35043
g34788 and n34920_not n35043_not ; n35044
g34789 and n34633_not n34919_not ; n35045
g34790 and n34918_not n35045 ; n35046
g34791 and n35044_not n35046_not ; n35047
g34792 and b[17]_not n35047_not ; n35048
g34793 and n34652_not n34838 ; n35049
g34794 and n34834_not n35049 ; n35050
g34795 and n34835_not n34838_not ; n35051
g34796 and n35050_not n35051_not ; n35052
g34797 and n34920_not n35052_not ; n35053
g34798 and n34642_not n34919_not ; n35054
g34799 and n34918_not n35054 ; n35055
g34800 and n35053_not n35055_not ; n35056
g34801 and b[16]_not n35056_not ; n35057
g34802 and n34661_not n34833 ; n35058
g34803 and n34829_not n35058 ; n35059
g34804 and n34830_not n34833_not ; n35060
g34805 and n35059_not n35060_not ; n35061
g34806 and n34920_not n35061_not ; n35062
g34807 and n34651_not n34919_not ; n35063
g34808 and n34918_not n35063 ; n35064
g34809 and n35062_not n35064_not ; n35065
g34810 and b[15]_not n35065_not ; n35066
g34811 and n34670_not n34828 ; n35067
g34812 and n34824_not n35067 ; n35068
g34813 and n34825_not n34828_not ; n35069
g34814 and n35068_not n35069_not ; n35070
g34815 and n34920_not n35070_not ; n35071
g34816 and n34660_not n34919_not ; n35072
g34817 and n34918_not n35072 ; n35073
g34818 and n35071_not n35073_not ; n35074
g34819 and b[14]_not n35074_not ; n35075
g34820 and n34679_not n34823 ; n35076
g34821 and n34819_not n35076 ; n35077
g34822 and n34820_not n34823_not ; n35078
g34823 and n35077_not n35078_not ; n35079
g34824 and n34920_not n35079_not ; n35080
g34825 and n34669_not n34919_not ; n35081
g34826 and n34918_not n35081 ; n35082
g34827 and n35080_not n35082_not ; n35083
g34828 and b[13]_not n35083_not ; n35084
g34829 and n34688_not n34818 ; n35085
g34830 and n34814_not n35085 ; n35086
g34831 and n34815_not n34818_not ; n35087
g34832 and n35086_not n35087_not ; n35088
g34833 and n34920_not n35088_not ; n35089
g34834 and n34678_not n34919_not ; n35090
g34835 and n34918_not n35090 ; n35091
g34836 and n35089_not n35091_not ; n35092
g34837 and b[12]_not n35092_not ; n35093
g34838 and n34697_not n34813 ; n35094
g34839 and n34809_not n35094 ; n35095
g34840 and n34810_not n34813_not ; n35096
g34841 and n35095_not n35096_not ; n35097
g34842 and n34920_not n35097_not ; n35098
g34843 and n34687_not n34919_not ; n35099
g34844 and n34918_not n35099 ; n35100
g34845 and n35098_not n35100_not ; n35101
g34846 and b[11]_not n35101_not ; n35102
g34847 and n34706_not n34808 ; n35103
g34848 and n34804_not n35103 ; n35104
g34849 and n34805_not n34808_not ; n35105
g34850 and n35104_not n35105_not ; n35106
g34851 and n34920_not n35106_not ; n35107
g34852 and n34696_not n34919_not ; n35108
g34853 and n34918_not n35108 ; n35109
g34854 and n35107_not n35109_not ; n35110
g34855 and b[10]_not n35110_not ; n35111
g34856 and n34715_not n34803 ; n35112
g34857 and n34799_not n35112 ; n35113
g34858 and n34800_not n34803_not ; n35114
g34859 and n35113_not n35114_not ; n35115
g34860 and n34920_not n35115_not ; n35116
g34861 and n34705_not n34919_not ; n35117
g34862 and n34918_not n35117 ; n35118
g34863 and n35116_not n35118_not ; n35119
g34864 and b[9]_not n35119_not ; n35120
g34865 and n34724_not n34798 ; n35121
g34866 and n34794_not n35121 ; n35122
g34867 and n34795_not n34798_not ; n35123
g34868 and n35122_not n35123_not ; n35124
g34869 and n34920_not n35124_not ; n35125
g34870 and n34714_not n34919_not ; n35126
g34871 and n34918_not n35126 ; n35127
g34872 and n35125_not n35127_not ; n35128
g34873 and b[8]_not n35128_not ; n35129
g34874 and n34733_not n34793 ; n35130
g34875 and n34789_not n35130 ; n35131
g34876 and n34790_not n34793_not ; n35132
g34877 and n35131_not n35132_not ; n35133
g34878 and n34920_not n35133_not ; n35134
g34879 and n34723_not n34919_not ; n35135
g34880 and n34918_not n35135 ; n35136
g34881 and n35134_not n35136_not ; n35137
g34882 and b[7]_not n35137_not ; n35138
g34883 and n34742_not n34788 ; n35139
g34884 and n34784_not n35139 ; n35140
g34885 and n34785_not n34788_not ; n35141
g34886 and n35140_not n35141_not ; n35142
g34887 and n34920_not n35142_not ; n35143
g34888 and n34732_not n34919_not ; n35144
g34889 and n34918_not n35144 ; n35145
g34890 and n35143_not n35145_not ; n35146
g34891 and b[6]_not n35146_not ; n35147
g34892 and n34751_not n34783 ; n35148
g34893 and n34779_not n35148 ; n35149
g34894 and n34780_not n34783_not ; n35150
g34895 and n35149_not n35150_not ; n35151
g34896 and n34920_not n35151_not ; n35152
g34897 and n34741_not n34919_not ; n35153
g34898 and n34918_not n35153 ; n35154
g34899 and n35152_not n35154_not ; n35155
g34900 and b[5]_not n35155_not ; n35156
g34901 and n34759_not n34778 ; n35157
g34902 and n34774_not n35157 ; n35158
g34903 and n34775_not n34778_not ; n35159
g34904 and n35158_not n35159_not ; n35160
g34905 and n34920_not n35160_not ; n35161
g34906 and n34750_not n34919_not ; n35162
g34907 and n34918_not n35162 ; n35163
g34908 and n35161_not n35163_not ; n35164
g34909 and b[4]_not n35164_not ; n35165
g34910 and n34769_not n34773 ; n35166
g34911 and n34768_not n35166 ; n35167
g34912 and n34770_not n34773_not ; n35168
g34913 and n35167_not n35168_not ; n35169
g34914 and n34920_not n35169_not ; n35170
g34915 and n34758_not n34919_not ; n35171
g34916 and n34918_not n35171 ; n35172
g34917 and n35170_not n35172_not ; n35173
g34918 and b[3]_not n35173_not ; n35174
g34919 and n6584 n34766_not ; n35175
g34920 and n34764_not n35175 ; n35176
g34921 and n34768_not n35176_not ; n35177
g34922 and n34920_not n35177 ; n35178
g34923 and n34763_not n34919_not ; n35179
g34924 and n34918_not n35179 ; n35180
g34925 and n35178_not n35180_not ; n35181
g34926 and b[2]_not n35181_not ; n35182
g34927 and b[0] n34920_not ; n35183
g34928 and a[34] n35183_not ; n35184
g34929 and n6584 n34920_not ; n35185
g34930 and n35184_not n35185_not ; n35186
g34931 and b[1] n35186_not ; n35187
g34932 and b[1]_not n35185_not ; n35188
g34933 and n35184_not n35188 ; n35189
g34934 and n35187_not n35189_not ; n35190
g34935 and n7011_not n35190_not ; n35191
g34936 and b[1]_not n35186_not ; n35192
g34937 and n35191_not n35192_not ; n35193
g34938 and b[2] n35180_not ; n35194
g34939 and n35178_not n35194 ; n35195
g34940 and n35182_not n35195_not ; n35196
g34941 and n35193_not n35196 ; n35197
g34942 and n35182_not n35197_not ; n35198
g34943 and b[3] n35172_not ; n35199
g34944 and n35170_not n35199 ; n35200
g34945 and n35174_not n35200_not ; n35201
g34946 and n35198_not n35201 ; n35202
g34947 and n35174_not n35202_not ; n35203
g34948 and b[4] n35163_not ; n35204
g34949 and n35161_not n35204 ; n35205
g34950 and n35165_not n35205_not ; n35206
g34951 and n35203_not n35206 ; n35207
g34952 and n35165_not n35207_not ; n35208
g34953 and b[5] n35154_not ; n35209
g34954 and n35152_not n35209 ; n35210
g34955 and n35156_not n35210_not ; n35211
g34956 and n35208_not n35211 ; n35212
g34957 and n35156_not n35212_not ; n35213
g34958 and b[6] n35145_not ; n35214
g34959 and n35143_not n35214 ; n35215
g34960 and n35147_not n35215_not ; n35216
g34961 and n35213_not n35216 ; n35217
g34962 and n35147_not n35217_not ; n35218
g34963 and b[7] n35136_not ; n35219
g34964 and n35134_not n35219 ; n35220
g34965 and n35138_not n35220_not ; n35221
g34966 and n35218_not n35221 ; n35222
g34967 and n35138_not n35222_not ; n35223
g34968 and b[8] n35127_not ; n35224
g34969 and n35125_not n35224 ; n35225
g34970 and n35129_not n35225_not ; n35226
g34971 and n35223_not n35226 ; n35227
g34972 and n35129_not n35227_not ; n35228
g34973 and b[9] n35118_not ; n35229
g34974 and n35116_not n35229 ; n35230
g34975 and n35120_not n35230_not ; n35231
g34976 and n35228_not n35231 ; n35232
g34977 and n35120_not n35232_not ; n35233
g34978 and b[10] n35109_not ; n35234
g34979 and n35107_not n35234 ; n35235
g34980 and n35111_not n35235_not ; n35236
g34981 and n35233_not n35236 ; n35237
g34982 and n35111_not n35237_not ; n35238
g34983 and b[11] n35100_not ; n35239
g34984 and n35098_not n35239 ; n35240
g34985 and n35102_not n35240_not ; n35241
g34986 and n35238_not n35241 ; n35242
g34987 and n35102_not n35242_not ; n35243
g34988 and b[12] n35091_not ; n35244
g34989 and n35089_not n35244 ; n35245
g34990 and n35093_not n35245_not ; n35246
g34991 and n35243_not n35246 ; n35247
g34992 and n35093_not n35247_not ; n35248
g34993 and b[13] n35082_not ; n35249
g34994 and n35080_not n35249 ; n35250
g34995 and n35084_not n35250_not ; n35251
g34996 and n35248_not n35251 ; n35252
g34997 and n35084_not n35252_not ; n35253
g34998 and b[14] n35073_not ; n35254
g34999 and n35071_not n35254 ; n35255
g35000 and n35075_not n35255_not ; n35256
g35001 and n35253_not n35256 ; n35257
g35002 and n35075_not n35257_not ; n35258
g35003 and b[15] n35064_not ; n35259
g35004 and n35062_not n35259 ; n35260
g35005 and n35066_not n35260_not ; n35261
g35006 and n35258_not n35261 ; n35262
g35007 and n35066_not n35262_not ; n35263
g35008 and b[16] n35055_not ; n35264
g35009 and n35053_not n35264 ; n35265
g35010 and n35057_not n35265_not ; n35266
g35011 and n35263_not n35266 ; n35267
g35012 and n35057_not n35267_not ; n35268
g35013 and b[17] n35046_not ; n35269
g35014 and n35044_not n35269 ; n35270
g35015 and n35048_not n35270_not ; n35271
g35016 and n35268_not n35271 ; n35272
g35017 and n35048_not n35272_not ; n35273
g35018 and b[18] n35037_not ; n35274
g35019 and n35035_not n35274 ; n35275
g35020 and n35039_not n35275_not ; n35276
g35021 and n35273_not n35276 ; n35277
g35022 and n35039_not n35277_not ; n35278
g35023 and b[19] n35028_not ; n35279
g35024 and n35026_not n35279 ; n35280
g35025 and n35030_not n35280_not ; n35281
g35026 and n35278_not n35281 ; n35282
g35027 and n35030_not n35282_not ; n35283
g35028 and b[20] n35019_not ; n35284
g35029 and n35017_not n35284 ; n35285
g35030 and n35021_not n35285_not ; n35286
g35031 and n35283_not n35286 ; n35287
g35032 and n35021_not n35287_not ; n35288
g35033 and b[21] n35010_not ; n35289
g35034 and n35008_not n35289 ; n35290
g35035 and n35012_not n35290_not ; n35291
g35036 and n35288_not n35291 ; n35292
g35037 and n35012_not n35292_not ; n35293
g35038 and b[22] n35001_not ; n35294
g35039 and n34999_not n35294 ; n35295
g35040 and n35003_not n35295_not ; n35296
g35041 and n35293_not n35296 ; n35297
g35042 and n35003_not n35297_not ; n35298
g35043 and b[23] n34992_not ; n35299
g35044 and n34990_not n35299 ; n35300
g35045 and n34994_not n35300_not ; n35301
g35046 and n35298_not n35301 ; n35302
g35047 and n34994_not n35302_not ; n35303
g35048 and b[24] n34983_not ; n35304
g35049 and n34981_not n35304 ; n35305
g35050 and n34985_not n35305_not ; n35306
g35051 and n35303_not n35306 ; n35307
g35052 and n34985_not n35307_not ; n35308
g35053 and b[25] n34974_not ; n35309
g35054 and n34972_not n35309 ; n35310
g35055 and n34976_not n35310_not ; n35311
g35056 and n35308_not n35311 ; n35312
g35057 and n34976_not n35312_not ; n35313
g35058 and b[26] n34965_not ; n35314
g35059 and n34963_not n35314 ; n35315
g35060 and n34967_not n35315_not ; n35316
g35061 and n35313_not n35316 ; n35317
g35062 and n34967_not n35317_not ; n35318
g35063 and b[27] n34956_not ; n35319
g35064 and n34954_not n35319 ; n35320
g35065 and n34958_not n35320_not ; n35321
g35066 and n35318_not n35321 ; n35322
g35067 and n34958_not n35322_not ; n35323
g35068 and b[28] n34947_not ; n35324
g35069 and n34945_not n35324 ; n35325
g35070 and n34949_not n35325_not ; n35326
g35071 and n35323_not n35326 ; n35327
g35072 and n34949_not n35327_not ; n35328
g35073 and b[29] n34927_not ; n35329
g35074 and n34925_not n35329 ; n35330
g35075 and n34940_not n35330_not ; n35331
g35076 and n35328_not n35331 ; n35332
g35077 and n34940_not n35332_not ; n35333
g35078 and b[30] n34937_not ; n35334
g35079 and n34935_not n35334 ; n35335
g35080 and n34939_not n35335_not ; n35336
g35081 and n35333_not n35336 ; n35337
g35082 and n34939_not n35337_not ; n35338
g35083 and n7162 n35338_not ; n35339
g35084 and n34928_not n35339_not ; n35340
g35085 and n34949_not n35331 ; n35341
g35086 and n35327_not n35341 ; n35342
g35087 and n35328_not n35331_not ; n35343
g35088 and n35342_not n35343_not ; n35344
g35089 and n7162 n35344_not ; n35345
g35090 and n35338_not n35345 ; n35346
g35091 and n35340_not n35346_not ; n35347
g35092 and n34938_not n35339_not ; n35348
g35093 and n34940_not n35336 ; n35349
g35094 and n35332_not n35349 ; n35350
g35095 and n35333_not n35336_not ; n35351
g35096 and n35350_not n35351_not ; n35352
g35097 and n35339 n35352_not ; n35353
g35098 and n35348_not n35353_not ; n35354
g35099 and b[31]_not n35354_not ; n35355
g35100 and b[30]_not n35347_not ; n35356
g35101 and n34948_not n35339_not ; n35357
g35102 and n34958_not n35326 ; n35358
g35103 and n35322_not n35358 ; n35359
g35104 and n35323_not n35326_not ; n35360
g35105 and n35359_not n35360_not ; n35361
g35106 and n7162 n35361_not ; n35362
g35107 and n35338_not n35362 ; n35363
g35108 and n35357_not n35363_not ; n35364
g35109 and b[29]_not n35364_not ; n35365
g35110 and n34957_not n35339_not ; n35366
g35111 and n34967_not n35321 ; n35367
g35112 and n35317_not n35367 ; n35368
g35113 and n35318_not n35321_not ; n35369
g35114 and n35368_not n35369_not ; n35370
g35115 and n7162 n35370_not ; n35371
g35116 and n35338_not n35371 ; n35372
g35117 and n35366_not n35372_not ; n35373
g35118 and b[28]_not n35373_not ; n35374
g35119 and n34966_not n35339_not ; n35375
g35120 and n34976_not n35316 ; n35376
g35121 and n35312_not n35376 ; n35377
g35122 and n35313_not n35316_not ; n35378
g35123 and n35377_not n35378_not ; n35379
g35124 and n7162 n35379_not ; n35380
g35125 and n35338_not n35380 ; n35381
g35126 and n35375_not n35381_not ; n35382
g35127 and b[27]_not n35382_not ; n35383
g35128 and n34975_not n35339_not ; n35384
g35129 and n34985_not n35311 ; n35385
g35130 and n35307_not n35385 ; n35386
g35131 and n35308_not n35311_not ; n35387
g35132 and n35386_not n35387_not ; n35388
g35133 and n7162 n35388_not ; n35389
g35134 and n35338_not n35389 ; n35390
g35135 and n35384_not n35390_not ; n35391
g35136 and b[26]_not n35391_not ; n35392
g35137 and n34984_not n35339_not ; n35393
g35138 and n34994_not n35306 ; n35394
g35139 and n35302_not n35394 ; n35395
g35140 and n35303_not n35306_not ; n35396
g35141 and n35395_not n35396_not ; n35397
g35142 and n7162 n35397_not ; n35398
g35143 and n35338_not n35398 ; n35399
g35144 and n35393_not n35399_not ; n35400
g35145 and b[25]_not n35400_not ; n35401
g35146 and n34993_not n35339_not ; n35402
g35147 and n35003_not n35301 ; n35403
g35148 and n35297_not n35403 ; n35404
g35149 and n35298_not n35301_not ; n35405
g35150 and n35404_not n35405_not ; n35406
g35151 and n7162 n35406_not ; n35407
g35152 and n35338_not n35407 ; n35408
g35153 and n35402_not n35408_not ; n35409
g35154 and b[24]_not n35409_not ; n35410
g35155 and n35002_not n35339_not ; n35411
g35156 and n35012_not n35296 ; n35412
g35157 and n35292_not n35412 ; n35413
g35158 and n35293_not n35296_not ; n35414
g35159 and n35413_not n35414_not ; n35415
g35160 and n7162 n35415_not ; n35416
g35161 and n35338_not n35416 ; n35417
g35162 and n35411_not n35417_not ; n35418
g35163 and b[23]_not n35418_not ; n35419
g35164 and n35011_not n35339_not ; n35420
g35165 and n35021_not n35291 ; n35421
g35166 and n35287_not n35421 ; n35422
g35167 and n35288_not n35291_not ; n35423
g35168 and n35422_not n35423_not ; n35424
g35169 and n7162 n35424_not ; n35425
g35170 and n35338_not n35425 ; n35426
g35171 and n35420_not n35426_not ; n35427
g35172 and b[22]_not n35427_not ; n35428
g35173 and n35020_not n35339_not ; n35429
g35174 and n35030_not n35286 ; n35430
g35175 and n35282_not n35430 ; n35431
g35176 and n35283_not n35286_not ; n35432
g35177 and n35431_not n35432_not ; n35433
g35178 and n7162 n35433_not ; n35434
g35179 and n35338_not n35434 ; n35435
g35180 and n35429_not n35435_not ; n35436
g35181 and b[21]_not n35436_not ; n35437
g35182 and n35029_not n35339_not ; n35438
g35183 and n35039_not n35281 ; n35439
g35184 and n35277_not n35439 ; n35440
g35185 and n35278_not n35281_not ; n35441
g35186 and n35440_not n35441_not ; n35442
g35187 and n7162 n35442_not ; n35443
g35188 and n35338_not n35443 ; n35444
g35189 and n35438_not n35444_not ; n35445
g35190 and b[20]_not n35445_not ; n35446
g35191 and n35038_not n35339_not ; n35447
g35192 and n35048_not n35276 ; n35448
g35193 and n35272_not n35448 ; n35449
g35194 and n35273_not n35276_not ; n35450
g35195 and n35449_not n35450_not ; n35451
g35196 and n7162 n35451_not ; n35452
g35197 and n35338_not n35452 ; n35453
g35198 and n35447_not n35453_not ; n35454
g35199 and b[19]_not n35454_not ; n35455
g35200 and n35047_not n35339_not ; n35456
g35201 and n35057_not n35271 ; n35457
g35202 and n35267_not n35457 ; n35458
g35203 and n35268_not n35271_not ; n35459
g35204 and n35458_not n35459_not ; n35460
g35205 and n7162 n35460_not ; n35461
g35206 and n35338_not n35461 ; n35462
g35207 and n35456_not n35462_not ; n35463
g35208 and b[18]_not n35463_not ; n35464
g35209 and n35056_not n35339_not ; n35465
g35210 and n35066_not n35266 ; n35466
g35211 and n35262_not n35466 ; n35467
g35212 and n35263_not n35266_not ; n35468
g35213 and n35467_not n35468_not ; n35469
g35214 and n7162 n35469_not ; n35470
g35215 and n35338_not n35470 ; n35471
g35216 and n35465_not n35471_not ; n35472
g35217 and b[17]_not n35472_not ; n35473
g35218 and n35065_not n35339_not ; n35474
g35219 and n35075_not n35261 ; n35475
g35220 and n35257_not n35475 ; n35476
g35221 and n35258_not n35261_not ; n35477
g35222 and n35476_not n35477_not ; n35478
g35223 and n7162 n35478_not ; n35479
g35224 and n35338_not n35479 ; n35480
g35225 and n35474_not n35480_not ; n35481
g35226 and b[16]_not n35481_not ; n35482
g35227 and n35074_not n35339_not ; n35483
g35228 and n35084_not n35256 ; n35484
g35229 and n35252_not n35484 ; n35485
g35230 and n35253_not n35256_not ; n35486
g35231 and n35485_not n35486_not ; n35487
g35232 and n7162 n35487_not ; n35488
g35233 and n35338_not n35488 ; n35489
g35234 and n35483_not n35489_not ; n35490
g35235 and b[15]_not n35490_not ; n35491
g35236 and n35083_not n35339_not ; n35492
g35237 and n35093_not n35251 ; n35493
g35238 and n35247_not n35493 ; n35494
g35239 and n35248_not n35251_not ; n35495
g35240 and n35494_not n35495_not ; n35496
g35241 and n7162 n35496_not ; n35497
g35242 and n35338_not n35497 ; n35498
g35243 and n35492_not n35498_not ; n35499
g35244 and b[14]_not n35499_not ; n35500
g35245 and n35092_not n35339_not ; n35501
g35246 and n35102_not n35246 ; n35502
g35247 and n35242_not n35502 ; n35503
g35248 and n35243_not n35246_not ; n35504
g35249 and n35503_not n35504_not ; n35505
g35250 and n7162 n35505_not ; n35506
g35251 and n35338_not n35506 ; n35507
g35252 and n35501_not n35507_not ; n35508
g35253 and b[13]_not n35508_not ; n35509
g35254 and n35101_not n35339_not ; n35510
g35255 and n35111_not n35241 ; n35511
g35256 and n35237_not n35511 ; n35512
g35257 and n35238_not n35241_not ; n35513
g35258 and n35512_not n35513_not ; n35514
g35259 and n7162 n35514_not ; n35515
g35260 and n35338_not n35515 ; n35516
g35261 and n35510_not n35516_not ; n35517
g35262 and b[12]_not n35517_not ; n35518
g35263 and n35110_not n35339_not ; n35519
g35264 and n35120_not n35236 ; n35520
g35265 and n35232_not n35520 ; n35521
g35266 and n35233_not n35236_not ; n35522
g35267 and n35521_not n35522_not ; n35523
g35268 and n7162 n35523_not ; n35524
g35269 and n35338_not n35524 ; n35525
g35270 and n35519_not n35525_not ; n35526
g35271 and b[11]_not n35526_not ; n35527
g35272 and n35119_not n35339_not ; n35528
g35273 and n35129_not n35231 ; n35529
g35274 and n35227_not n35529 ; n35530
g35275 and n35228_not n35231_not ; n35531
g35276 and n35530_not n35531_not ; n35532
g35277 and n7162 n35532_not ; n35533
g35278 and n35338_not n35533 ; n35534
g35279 and n35528_not n35534_not ; n35535
g35280 and b[10]_not n35535_not ; n35536
g35281 and n35128_not n35339_not ; n35537
g35282 and n35138_not n35226 ; n35538
g35283 and n35222_not n35538 ; n35539
g35284 and n35223_not n35226_not ; n35540
g35285 and n35539_not n35540_not ; n35541
g35286 and n7162 n35541_not ; n35542
g35287 and n35338_not n35542 ; n35543
g35288 and n35537_not n35543_not ; n35544
g35289 and b[9]_not n35544_not ; n35545
g35290 and n35137_not n35339_not ; n35546
g35291 and n35147_not n35221 ; n35547
g35292 and n35217_not n35547 ; n35548
g35293 and n35218_not n35221_not ; n35549
g35294 and n35548_not n35549_not ; n35550
g35295 and n7162 n35550_not ; n35551
g35296 and n35338_not n35551 ; n35552
g35297 and n35546_not n35552_not ; n35553
g35298 and b[8]_not n35553_not ; n35554
g35299 and n35146_not n35339_not ; n35555
g35300 and n35156_not n35216 ; n35556
g35301 and n35212_not n35556 ; n35557
g35302 and n35213_not n35216_not ; n35558
g35303 and n35557_not n35558_not ; n35559
g35304 and n7162 n35559_not ; n35560
g35305 and n35338_not n35560 ; n35561
g35306 and n35555_not n35561_not ; n35562
g35307 and b[7]_not n35562_not ; n35563
g35308 and n35155_not n35339_not ; n35564
g35309 and n35165_not n35211 ; n35565
g35310 and n35207_not n35565 ; n35566
g35311 and n35208_not n35211_not ; n35567
g35312 and n35566_not n35567_not ; n35568
g35313 and n7162 n35568_not ; n35569
g35314 and n35338_not n35569 ; n35570
g35315 and n35564_not n35570_not ; n35571
g35316 and b[6]_not n35571_not ; n35572
g35317 and n35164_not n35339_not ; n35573
g35318 and n35174_not n35206 ; n35574
g35319 and n35202_not n35574 ; n35575
g35320 and n35203_not n35206_not ; n35576
g35321 and n35575_not n35576_not ; n35577
g35322 and n7162 n35577_not ; n35578
g35323 and n35338_not n35578 ; n35579
g35324 and n35573_not n35579_not ; n35580
g35325 and b[5]_not n35580_not ; n35581
g35326 and n35173_not n35339_not ; n35582
g35327 and n35182_not n35201 ; n35583
g35328 and n35197_not n35583 ; n35584
g35329 and n35198_not n35201_not ; n35585
g35330 and n35584_not n35585_not ; n35586
g35331 and n7162 n35586_not ; n35587
g35332 and n35338_not n35587 ; n35588
g35333 and n35582_not n35588_not ; n35589
g35334 and b[4]_not n35589_not ; n35590
g35335 and n35181_not n35339_not ; n35591
g35336 and n35192_not n35196 ; n35592
g35337 and n35191_not n35592 ; n35593
g35338 and n35193_not n35196_not ; n35594
g35339 and n35593_not n35594_not ; n35595
g35340 and n7162 n35595_not ; n35596
g35341 and n35338_not n35596 ; n35597
g35342 and n35591_not n35597_not ; n35598
g35343 and b[3]_not n35598_not ; n35599
g35344 and n35186_not n35339_not ; n35600
g35345 and n7011 n35189_not ; n35601
g35346 and n35187_not n35601 ; n35602
g35347 and n7162 n35602_not ; n35603
g35348 and n35191_not n35603 ; n35604
g35349 and n35338_not n35604 ; n35605
g35350 and n35600_not n35605_not ; n35606
g35351 and b[2]_not n35606_not ; n35607
g35352 and n7435 n35338_not ; n35608
g35353 and a[33] n35608_not ; n35609
g35354 and n7441 n35338_not ; n35610
g35355 and n35609_not n35610_not ; n35611
g35356 and b[1] n35611_not ; n35612
g35357 and b[1]_not n35610_not ; n35613
g35358 and n35609_not n35613 ; n35614
g35359 and n35612_not n35614_not ; n35615
g35360 and n7448_not n35615_not ; n35616
g35361 and b[1]_not n35611_not ; n35617
g35362 and n35616_not n35617_not ; n35618
g35363 and b[2] n35605_not ; n35619
g35364 and n35600_not n35619 ; n35620
g35365 and n35607_not n35620_not ; n35621
g35366 and n35618_not n35621 ; n35622
g35367 and n35607_not n35622_not ; n35623
g35368 and b[3] n35597_not ; n35624
g35369 and n35591_not n35624 ; n35625
g35370 and n35599_not n35625_not ; n35626
g35371 and n35623_not n35626 ; n35627
g35372 and n35599_not n35627_not ; n35628
g35373 and b[4] n35588_not ; n35629
g35374 and n35582_not n35629 ; n35630
g35375 and n35590_not n35630_not ; n35631
g35376 and n35628_not n35631 ; n35632
g35377 and n35590_not n35632_not ; n35633
g35378 and b[5] n35579_not ; n35634
g35379 and n35573_not n35634 ; n35635
g35380 and n35581_not n35635_not ; n35636
g35381 and n35633_not n35636 ; n35637
g35382 and n35581_not n35637_not ; n35638
g35383 and b[6] n35570_not ; n35639
g35384 and n35564_not n35639 ; n35640
g35385 and n35572_not n35640_not ; n35641
g35386 and n35638_not n35641 ; n35642
g35387 and n35572_not n35642_not ; n35643
g35388 and b[7] n35561_not ; n35644
g35389 and n35555_not n35644 ; n35645
g35390 and n35563_not n35645_not ; n35646
g35391 and n35643_not n35646 ; n35647
g35392 and n35563_not n35647_not ; n35648
g35393 and b[8] n35552_not ; n35649
g35394 and n35546_not n35649 ; n35650
g35395 and n35554_not n35650_not ; n35651
g35396 and n35648_not n35651 ; n35652
g35397 and n35554_not n35652_not ; n35653
g35398 and b[9] n35543_not ; n35654
g35399 and n35537_not n35654 ; n35655
g35400 and n35545_not n35655_not ; n35656
g35401 and n35653_not n35656 ; n35657
g35402 and n35545_not n35657_not ; n35658
g35403 and b[10] n35534_not ; n35659
g35404 and n35528_not n35659 ; n35660
g35405 and n35536_not n35660_not ; n35661
g35406 and n35658_not n35661 ; n35662
g35407 and n35536_not n35662_not ; n35663
g35408 and b[11] n35525_not ; n35664
g35409 and n35519_not n35664 ; n35665
g35410 and n35527_not n35665_not ; n35666
g35411 and n35663_not n35666 ; n35667
g35412 and n35527_not n35667_not ; n35668
g35413 and b[12] n35516_not ; n35669
g35414 and n35510_not n35669 ; n35670
g35415 and n35518_not n35670_not ; n35671
g35416 and n35668_not n35671 ; n35672
g35417 and n35518_not n35672_not ; n35673
g35418 and b[13] n35507_not ; n35674
g35419 and n35501_not n35674 ; n35675
g35420 and n35509_not n35675_not ; n35676
g35421 and n35673_not n35676 ; n35677
g35422 and n35509_not n35677_not ; n35678
g35423 and b[14] n35498_not ; n35679
g35424 and n35492_not n35679 ; n35680
g35425 and n35500_not n35680_not ; n35681
g35426 and n35678_not n35681 ; n35682
g35427 and n35500_not n35682_not ; n35683
g35428 and b[15] n35489_not ; n35684
g35429 and n35483_not n35684 ; n35685
g35430 and n35491_not n35685_not ; n35686
g35431 and n35683_not n35686 ; n35687
g35432 and n35491_not n35687_not ; n35688
g35433 and b[16] n35480_not ; n35689
g35434 and n35474_not n35689 ; n35690
g35435 and n35482_not n35690_not ; n35691
g35436 and n35688_not n35691 ; n35692
g35437 and n35482_not n35692_not ; n35693
g35438 and b[17] n35471_not ; n35694
g35439 and n35465_not n35694 ; n35695
g35440 and n35473_not n35695_not ; n35696
g35441 and n35693_not n35696 ; n35697
g35442 and n35473_not n35697_not ; n35698
g35443 and b[18] n35462_not ; n35699
g35444 and n35456_not n35699 ; n35700
g35445 and n35464_not n35700_not ; n35701
g35446 and n35698_not n35701 ; n35702
g35447 and n35464_not n35702_not ; n35703
g35448 and b[19] n35453_not ; n35704
g35449 and n35447_not n35704 ; n35705
g35450 and n35455_not n35705_not ; n35706
g35451 and n35703_not n35706 ; n35707
g35452 and n35455_not n35707_not ; n35708
g35453 and b[20] n35444_not ; n35709
g35454 and n35438_not n35709 ; n35710
g35455 and n35446_not n35710_not ; n35711
g35456 and n35708_not n35711 ; n35712
g35457 and n35446_not n35712_not ; n35713
g35458 and b[21] n35435_not ; n35714
g35459 and n35429_not n35714 ; n35715
g35460 and n35437_not n35715_not ; n35716
g35461 and n35713_not n35716 ; n35717
g35462 and n35437_not n35717_not ; n35718
g35463 and b[22] n35426_not ; n35719
g35464 and n35420_not n35719 ; n35720
g35465 and n35428_not n35720_not ; n35721
g35466 and n35718_not n35721 ; n35722
g35467 and n35428_not n35722_not ; n35723
g35468 and b[23] n35417_not ; n35724
g35469 and n35411_not n35724 ; n35725
g35470 and n35419_not n35725_not ; n35726
g35471 and n35723_not n35726 ; n35727
g35472 and n35419_not n35727_not ; n35728
g35473 and b[24] n35408_not ; n35729
g35474 and n35402_not n35729 ; n35730
g35475 and n35410_not n35730_not ; n35731
g35476 and n35728_not n35731 ; n35732
g35477 and n35410_not n35732_not ; n35733
g35478 and b[25] n35399_not ; n35734
g35479 and n35393_not n35734 ; n35735
g35480 and n35401_not n35735_not ; n35736
g35481 and n35733_not n35736 ; n35737
g35482 and n35401_not n35737_not ; n35738
g35483 and b[26] n35390_not ; n35739
g35484 and n35384_not n35739 ; n35740
g35485 and n35392_not n35740_not ; n35741
g35486 and n35738_not n35741 ; n35742
g35487 and n35392_not n35742_not ; n35743
g35488 and b[27] n35381_not ; n35744
g35489 and n35375_not n35744 ; n35745
g35490 and n35383_not n35745_not ; n35746
g35491 and n35743_not n35746 ; n35747
g35492 and n35383_not n35747_not ; n35748
g35493 and b[28] n35372_not ; n35749
g35494 and n35366_not n35749 ; n35750
g35495 and n35374_not n35750_not ; n35751
g35496 and n35748_not n35751 ; n35752
g35497 and n35374_not n35752_not ; n35753
g35498 and b[29] n35363_not ; n35754
g35499 and n35357_not n35754 ; n35755
g35500 and n35365_not n35755_not ; n35756
g35501 and n35753_not n35756 ; n35757
g35502 and n35365_not n35757_not ; n35758
g35503 and b[30] n35346_not ; n35759
g35504 and n35340_not n35759 ; n35760
g35505 and n35356_not n35760_not ; n35761
g35506 and n35758_not n35761 ; n35762
g35507 and n35356_not n35762_not ; n35763
g35508 and b[31] n35348_not ; n35764
g35509 and n35353_not n35764 ; n35765
g35510 and n35355_not n35765_not ; n35766
g35511 and n35763_not n35766 ; n35767
g35512 and n35355_not n35767_not ; n35768
g35513 and n432 n35768_not ; n35769
g35514 and n35347_not n35769_not ; n35770
g35515 and n35365_not n35761 ; n35771
g35516 and n35757_not n35771 ; n35772
g35517 and n35758_not n35761_not ; n35773
g35518 and n35772_not n35773_not ; n35774
g35519 and n432 n35774_not ; n35775
g35520 and n35768_not n35775 ; n35776
g35521 and n35770_not n35776_not ; n35777
g35522 and b[31]_not n35777_not ; n35778
g35523 and n35364_not n35769_not ; n35779
g35524 and n35374_not n35756 ; n35780
g35525 and n35752_not n35780 ; n35781
g35526 and n35753_not n35756_not ; n35782
g35527 and n35781_not n35782_not ; n35783
g35528 and n432 n35783_not ; n35784
g35529 and n35768_not n35784 ; n35785
g35530 and n35779_not n35785_not ; n35786
g35531 and b[30]_not n35786_not ; n35787
g35532 and n35373_not n35769_not ; n35788
g35533 and n35383_not n35751 ; n35789
g35534 and n35747_not n35789 ; n35790
g35535 and n35748_not n35751_not ; n35791
g35536 and n35790_not n35791_not ; n35792
g35537 and n432 n35792_not ; n35793
g35538 and n35768_not n35793 ; n35794
g35539 and n35788_not n35794_not ; n35795
g35540 and b[29]_not n35795_not ; n35796
g35541 and n35382_not n35769_not ; n35797
g35542 and n35392_not n35746 ; n35798
g35543 and n35742_not n35798 ; n35799
g35544 and n35743_not n35746_not ; n35800
g35545 and n35799_not n35800_not ; n35801
g35546 and n432 n35801_not ; n35802
g35547 and n35768_not n35802 ; n35803
g35548 and n35797_not n35803_not ; n35804
g35549 and b[28]_not n35804_not ; n35805
g35550 and n35391_not n35769_not ; n35806
g35551 and n35401_not n35741 ; n35807
g35552 and n35737_not n35807 ; n35808
g35553 and n35738_not n35741_not ; n35809
g35554 and n35808_not n35809_not ; n35810
g35555 and n432 n35810_not ; n35811
g35556 and n35768_not n35811 ; n35812
g35557 and n35806_not n35812_not ; n35813
g35558 and b[27]_not n35813_not ; n35814
g35559 and n35400_not n35769_not ; n35815
g35560 and n35410_not n35736 ; n35816
g35561 and n35732_not n35816 ; n35817
g35562 and n35733_not n35736_not ; n35818
g35563 and n35817_not n35818_not ; n35819
g35564 and n432 n35819_not ; n35820
g35565 and n35768_not n35820 ; n35821
g35566 and n35815_not n35821_not ; n35822
g35567 and b[26]_not n35822_not ; n35823
g35568 and n35409_not n35769_not ; n35824
g35569 and n35419_not n35731 ; n35825
g35570 and n35727_not n35825 ; n35826
g35571 and n35728_not n35731_not ; n35827
g35572 and n35826_not n35827_not ; n35828
g35573 and n432 n35828_not ; n35829
g35574 and n35768_not n35829 ; n35830
g35575 and n35824_not n35830_not ; n35831
g35576 and b[25]_not n35831_not ; n35832
g35577 and n35418_not n35769_not ; n35833
g35578 and n35428_not n35726 ; n35834
g35579 and n35722_not n35834 ; n35835
g35580 and n35723_not n35726_not ; n35836
g35581 and n35835_not n35836_not ; n35837
g35582 and n432 n35837_not ; n35838
g35583 and n35768_not n35838 ; n35839
g35584 and n35833_not n35839_not ; n35840
g35585 and b[24]_not n35840_not ; n35841
g35586 and n35427_not n35769_not ; n35842
g35587 and n35437_not n35721 ; n35843
g35588 and n35717_not n35843 ; n35844
g35589 and n35718_not n35721_not ; n35845
g35590 and n35844_not n35845_not ; n35846
g35591 and n432 n35846_not ; n35847
g35592 and n35768_not n35847 ; n35848
g35593 and n35842_not n35848_not ; n35849
g35594 and b[23]_not n35849_not ; n35850
g35595 and n35436_not n35769_not ; n35851
g35596 and n35446_not n35716 ; n35852
g35597 and n35712_not n35852 ; n35853
g35598 and n35713_not n35716_not ; n35854
g35599 and n35853_not n35854_not ; n35855
g35600 and n432 n35855_not ; n35856
g35601 and n35768_not n35856 ; n35857
g35602 and n35851_not n35857_not ; n35858
g35603 and b[22]_not n35858_not ; n35859
g35604 and n35445_not n35769_not ; n35860
g35605 and n35455_not n35711 ; n35861
g35606 and n35707_not n35861 ; n35862
g35607 and n35708_not n35711_not ; n35863
g35608 and n35862_not n35863_not ; n35864
g35609 and n432 n35864_not ; n35865
g35610 and n35768_not n35865 ; n35866
g35611 and n35860_not n35866_not ; n35867
g35612 and b[21]_not n35867_not ; n35868
g35613 and n35454_not n35769_not ; n35869
g35614 and n35464_not n35706 ; n35870
g35615 and n35702_not n35870 ; n35871
g35616 and n35703_not n35706_not ; n35872
g35617 and n35871_not n35872_not ; n35873
g35618 and n432 n35873_not ; n35874
g35619 and n35768_not n35874 ; n35875
g35620 and n35869_not n35875_not ; n35876
g35621 and b[20]_not n35876_not ; n35877
g35622 and n35463_not n35769_not ; n35878
g35623 and n35473_not n35701 ; n35879
g35624 and n35697_not n35879 ; n35880
g35625 and n35698_not n35701_not ; n35881
g35626 and n35880_not n35881_not ; n35882
g35627 and n432 n35882_not ; n35883
g35628 and n35768_not n35883 ; n35884
g35629 and n35878_not n35884_not ; n35885
g35630 and b[19]_not n35885_not ; n35886
g35631 and n35472_not n35769_not ; n35887
g35632 and n35482_not n35696 ; n35888
g35633 and n35692_not n35888 ; n35889
g35634 and n35693_not n35696_not ; n35890
g35635 and n35889_not n35890_not ; n35891
g35636 and n432 n35891_not ; n35892
g35637 and n35768_not n35892 ; n35893
g35638 and n35887_not n35893_not ; n35894
g35639 and b[18]_not n35894_not ; n35895
g35640 and n35481_not n35769_not ; n35896
g35641 and n35491_not n35691 ; n35897
g35642 and n35687_not n35897 ; n35898
g35643 and n35688_not n35691_not ; n35899
g35644 and n35898_not n35899_not ; n35900
g35645 and n432 n35900_not ; n35901
g35646 and n35768_not n35901 ; n35902
g35647 and n35896_not n35902_not ; n35903
g35648 and b[17]_not n35903_not ; n35904
g35649 and n35490_not n35769_not ; n35905
g35650 and n35500_not n35686 ; n35906
g35651 and n35682_not n35906 ; n35907
g35652 and n35683_not n35686_not ; n35908
g35653 and n35907_not n35908_not ; n35909
g35654 and n432 n35909_not ; n35910
g35655 and n35768_not n35910 ; n35911
g35656 and n35905_not n35911_not ; n35912
g35657 and b[16]_not n35912_not ; n35913
g35658 and n35499_not n35769_not ; n35914
g35659 and n35509_not n35681 ; n35915
g35660 and n35677_not n35915 ; n35916
g35661 and n35678_not n35681_not ; n35917
g35662 and n35916_not n35917_not ; n35918
g35663 and n432 n35918_not ; n35919
g35664 and n35768_not n35919 ; n35920
g35665 and n35914_not n35920_not ; n35921
g35666 and b[15]_not n35921_not ; n35922
g35667 and n35508_not n35769_not ; n35923
g35668 and n35518_not n35676 ; n35924
g35669 and n35672_not n35924 ; n35925
g35670 and n35673_not n35676_not ; n35926
g35671 and n35925_not n35926_not ; n35927
g35672 and n432 n35927_not ; n35928
g35673 and n35768_not n35928 ; n35929
g35674 and n35923_not n35929_not ; n35930
g35675 and b[14]_not n35930_not ; n35931
g35676 and n35517_not n35769_not ; n35932
g35677 and n35527_not n35671 ; n35933
g35678 and n35667_not n35933 ; n35934
g35679 and n35668_not n35671_not ; n35935
g35680 and n35934_not n35935_not ; n35936
g35681 and n432 n35936_not ; n35937
g35682 and n35768_not n35937 ; n35938
g35683 and n35932_not n35938_not ; n35939
g35684 and b[13]_not n35939_not ; n35940
g35685 and n35526_not n35769_not ; n35941
g35686 and n35536_not n35666 ; n35942
g35687 and n35662_not n35942 ; n35943
g35688 and n35663_not n35666_not ; n35944
g35689 and n35943_not n35944_not ; n35945
g35690 and n432 n35945_not ; n35946
g35691 and n35768_not n35946 ; n35947
g35692 and n35941_not n35947_not ; n35948
g35693 and b[12]_not n35948_not ; n35949
g35694 and n35535_not n35769_not ; n35950
g35695 and n35545_not n35661 ; n35951
g35696 and n35657_not n35951 ; n35952
g35697 and n35658_not n35661_not ; n35953
g35698 and n35952_not n35953_not ; n35954
g35699 and n432 n35954_not ; n35955
g35700 and n35768_not n35955 ; n35956
g35701 and n35950_not n35956_not ; n35957
g35702 and b[11]_not n35957_not ; n35958
g35703 and n35544_not n35769_not ; n35959
g35704 and n35554_not n35656 ; n35960
g35705 and n35652_not n35960 ; n35961
g35706 and n35653_not n35656_not ; n35962
g35707 and n35961_not n35962_not ; n35963
g35708 and n432 n35963_not ; n35964
g35709 and n35768_not n35964 ; n35965
g35710 and n35959_not n35965_not ; n35966
g35711 and b[10]_not n35966_not ; n35967
g35712 and n35553_not n35769_not ; n35968
g35713 and n35563_not n35651 ; n35969
g35714 and n35647_not n35969 ; n35970
g35715 and n35648_not n35651_not ; n35971
g35716 and n35970_not n35971_not ; n35972
g35717 and n432 n35972_not ; n35973
g35718 and n35768_not n35973 ; n35974
g35719 and n35968_not n35974_not ; n35975
g35720 and b[9]_not n35975_not ; n35976
g35721 and n35562_not n35769_not ; n35977
g35722 and n35572_not n35646 ; n35978
g35723 and n35642_not n35978 ; n35979
g35724 and n35643_not n35646_not ; n35980
g35725 and n35979_not n35980_not ; n35981
g35726 and n432 n35981_not ; n35982
g35727 and n35768_not n35982 ; n35983
g35728 and n35977_not n35983_not ; n35984
g35729 and b[8]_not n35984_not ; n35985
g35730 and n35571_not n35769_not ; n35986
g35731 and n35581_not n35641 ; n35987
g35732 and n35637_not n35987 ; n35988
g35733 and n35638_not n35641_not ; n35989
g35734 and n35988_not n35989_not ; n35990
g35735 and n432 n35990_not ; n35991
g35736 and n35768_not n35991 ; n35992
g35737 and n35986_not n35992_not ; n35993
g35738 and b[7]_not n35993_not ; n35994
g35739 and n35580_not n35769_not ; n35995
g35740 and n35590_not n35636 ; n35996
g35741 and n35632_not n35996 ; n35997
g35742 and n35633_not n35636_not ; n35998
g35743 and n35997_not n35998_not ; n35999
g35744 and n432 n35999_not ; n36000
g35745 and n35768_not n36000 ; n36001
g35746 and n35995_not n36001_not ; n36002
g35747 and b[6]_not n36002_not ; n36003
g35748 and n35589_not n35769_not ; n36004
g35749 and n35599_not n35631 ; n36005
g35750 and n35627_not n36005 ; n36006
g35751 and n35628_not n35631_not ; n36007
g35752 and n36006_not n36007_not ; n36008
g35753 and n432 n36008_not ; n36009
g35754 and n35768_not n36009 ; n36010
g35755 and n36004_not n36010_not ; n36011
g35756 and b[5]_not n36011_not ; n36012
g35757 and n35598_not n35769_not ; n36013
g35758 and n35607_not n35626 ; n36014
g35759 and n35622_not n36014 ; n36015
g35760 and n35623_not n35626_not ; n36016
g35761 and n36015_not n36016_not ; n36017
g35762 and n432 n36017_not ; n36018
g35763 and n35768_not n36018 ; n36019
g35764 and n36013_not n36019_not ; n36020
g35765 and b[4]_not n36020_not ; n36021
g35766 and n35606_not n35769_not ; n36022
g35767 and n35617_not n35621 ; n36023
g35768 and n35616_not n36023 ; n36024
g35769 and n35618_not n35621_not ; n36025
g35770 and n36024_not n36025_not ; n36026
g35771 and n432 n36026_not ; n36027
g35772 and n35768_not n36027 ; n36028
g35773 and n36022_not n36028_not ; n36029
g35774 and b[3]_not n36029_not ; n36030
g35775 and n35611_not n35769_not ; n36031
g35776 and n7448 n35614_not ; n36032
g35777 and n35612_not n36032 ; n36033
g35778 and n432 n36033_not ; n36034
g35779 and n35616_not n36034 ; n36035
g35780 and n35768_not n36035 ; n36036
g35781 and n36031_not n36036_not ; n36037
g35782 and b[2]_not n36037_not ; n36038
g35783 and n7875 n35768_not ; n36039
g35784 and a[32] n36039_not ; n36040
g35785 and n7880 n35768_not ; n36041
g35786 and n36040_not n36041_not ; n36042
g35787 and b[1] n36042_not ; n36043
g35788 and b[1]_not n36041_not ; n36044
g35789 and n36040_not n36044 ; n36045
g35790 and n36043_not n36045_not ; n36046
g35791 and n7887_not n36046_not ; n36047
g35792 and b[1]_not n36042_not ; n36048
g35793 and n36047_not n36048_not ; n36049
g35794 and b[2] n36036_not ; n36050
g35795 and n36031_not n36050 ; n36051
g35796 and n36038_not n36051_not ; n36052
g35797 and n36049_not n36052 ; n36053
g35798 and n36038_not n36053_not ; n36054
g35799 and b[3] n36028_not ; n36055
g35800 and n36022_not n36055 ; n36056
g35801 and n36030_not n36056_not ; n36057
g35802 and n36054_not n36057 ; n36058
g35803 and n36030_not n36058_not ; n36059
g35804 and b[4] n36019_not ; n36060
g35805 and n36013_not n36060 ; n36061
g35806 and n36021_not n36061_not ; n36062
g35807 and n36059_not n36062 ; n36063
g35808 and n36021_not n36063_not ; n36064
g35809 and b[5] n36010_not ; n36065
g35810 and n36004_not n36065 ; n36066
g35811 and n36012_not n36066_not ; n36067
g35812 and n36064_not n36067 ; n36068
g35813 and n36012_not n36068_not ; n36069
g35814 and b[6] n36001_not ; n36070
g35815 and n35995_not n36070 ; n36071
g35816 and n36003_not n36071_not ; n36072
g35817 and n36069_not n36072 ; n36073
g35818 and n36003_not n36073_not ; n36074
g35819 and b[7] n35992_not ; n36075
g35820 and n35986_not n36075 ; n36076
g35821 and n35994_not n36076_not ; n36077
g35822 and n36074_not n36077 ; n36078
g35823 and n35994_not n36078_not ; n36079
g35824 and b[8] n35983_not ; n36080
g35825 and n35977_not n36080 ; n36081
g35826 and n35985_not n36081_not ; n36082
g35827 and n36079_not n36082 ; n36083
g35828 and n35985_not n36083_not ; n36084
g35829 and b[9] n35974_not ; n36085
g35830 and n35968_not n36085 ; n36086
g35831 and n35976_not n36086_not ; n36087
g35832 and n36084_not n36087 ; n36088
g35833 and n35976_not n36088_not ; n36089
g35834 and b[10] n35965_not ; n36090
g35835 and n35959_not n36090 ; n36091
g35836 and n35967_not n36091_not ; n36092
g35837 and n36089_not n36092 ; n36093
g35838 and n35967_not n36093_not ; n36094
g35839 and b[11] n35956_not ; n36095
g35840 and n35950_not n36095 ; n36096
g35841 and n35958_not n36096_not ; n36097
g35842 and n36094_not n36097 ; n36098
g35843 and n35958_not n36098_not ; n36099
g35844 and b[12] n35947_not ; n36100
g35845 and n35941_not n36100 ; n36101
g35846 and n35949_not n36101_not ; n36102
g35847 and n36099_not n36102 ; n36103
g35848 and n35949_not n36103_not ; n36104
g35849 and b[13] n35938_not ; n36105
g35850 and n35932_not n36105 ; n36106
g35851 and n35940_not n36106_not ; n36107
g35852 and n36104_not n36107 ; n36108
g35853 and n35940_not n36108_not ; n36109
g35854 and b[14] n35929_not ; n36110
g35855 and n35923_not n36110 ; n36111
g35856 and n35931_not n36111_not ; n36112
g35857 and n36109_not n36112 ; n36113
g35858 and n35931_not n36113_not ; n36114
g35859 and b[15] n35920_not ; n36115
g35860 and n35914_not n36115 ; n36116
g35861 and n35922_not n36116_not ; n36117
g35862 and n36114_not n36117 ; n36118
g35863 and n35922_not n36118_not ; n36119
g35864 and b[16] n35911_not ; n36120
g35865 and n35905_not n36120 ; n36121
g35866 and n35913_not n36121_not ; n36122
g35867 and n36119_not n36122 ; n36123
g35868 and n35913_not n36123_not ; n36124
g35869 and b[17] n35902_not ; n36125
g35870 and n35896_not n36125 ; n36126
g35871 and n35904_not n36126_not ; n36127
g35872 and n36124_not n36127 ; n36128
g35873 and n35904_not n36128_not ; n36129
g35874 and b[18] n35893_not ; n36130
g35875 and n35887_not n36130 ; n36131
g35876 and n35895_not n36131_not ; n36132
g35877 and n36129_not n36132 ; n36133
g35878 and n35895_not n36133_not ; n36134
g35879 and b[19] n35884_not ; n36135
g35880 and n35878_not n36135 ; n36136
g35881 and n35886_not n36136_not ; n36137
g35882 and n36134_not n36137 ; n36138
g35883 and n35886_not n36138_not ; n36139
g35884 and b[20] n35875_not ; n36140
g35885 and n35869_not n36140 ; n36141
g35886 and n35877_not n36141_not ; n36142
g35887 and n36139_not n36142 ; n36143
g35888 and n35877_not n36143_not ; n36144
g35889 and b[21] n35866_not ; n36145
g35890 and n35860_not n36145 ; n36146
g35891 and n35868_not n36146_not ; n36147
g35892 and n36144_not n36147 ; n36148
g35893 and n35868_not n36148_not ; n36149
g35894 and b[22] n35857_not ; n36150
g35895 and n35851_not n36150 ; n36151
g35896 and n35859_not n36151_not ; n36152
g35897 and n36149_not n36152 ; n36153
g35898 and n35859_not n36153_not ; n36154
g35899 and b[23] n35848_not ; n36155
g35900 and n35842_not n36155 ; n36156
g35901 and n35850_not n36156_not ; n36157
g35902 and n36154_not n36157 ; n36158
g35903 and n35850_not n36158_not ; n36159
g35904 and b[24] n35839_not ; n36160
g35905 and n35833_not n36160 ; n36161
g35906 and n35841_not n36161_not ; n36162
g35907 and n36159_not n36162 ; n36163
g35908 and n35841_not n36163_not ; n36164
g35909 and b[25] n35830_not ; n36165
g35910 and n35824_not n36165 ; n36166
g35911 and n35832_not n36166_not ; n36167
g35912 and n36164_not n36167 ; n36168
g35913 and n35832_not n36168_not ; n36169
g35914 and b[26] n35821_not ; n36170
g35915 and n35815_not n36170 ; n36171
g35916 and n35823_not n36171_not ; n36172
g35917 and n36169_not n36172 ; n36173
g35918 and n35823_not n36173_not ; n36174
g35919 and b[27] n35812_not ; n36175
g35920 and n35806_not n36175 ; n36176
g35921 and n35814_not n36176_not ; n36177
g35922 and n36174_not n36177 ; n36178
g35923 and n35814_not n36178_not ; n36179
g35924 and b[28] n35803_not ; n36180
g35925 and n35797_not n36180 ; n36181
g35926 and n35805_not n36181_not ; n36182
g35927 and n36179_not n36182 ; n36183
g35928 and n35805_not n36183_not ; n36184
g35929 and b[29] n35794_not ; n36185
g35930 and n35788_not n36185 ; n36186
g35931 and n35796_not n36186_not ; n36187
g35932 and n36184_not n36187 ; n36188
g35933 and n35796_not n36188_not ; n36189
g35934 and b[30] n35785_not ; n36190
g35935 and n35779_not n36190 ; n36191
g35936 and n35787_not n36191_not ; n36192
g35937 and n36189_not n36192 ; n36193
g35938 and n35787_not n36193_not ; n36194
g35939 and b[31] n35776_not ; n36195
g35940 and n35770_not n36195 ; n36196
g35941 and n35778_not n36196_not ; n36197
g35942 and n36194_not n36197 ; n36198
g35943 and n35778_not n36198_not ; n36199
g35944 and n35354_not n35769_not ; n36200
g35945 and n35356_not n35766 ; n36201
g35946 and n35762_not n36201 ; n36202
g35947 and n35763_not n35766_not ; n36203
g35948 and n36202_not n36203_not ; n36204
g35949 and n35769 n36204_not ; n36205
g35950 and n36200_not n36205_not ; n36206
g35951 and b[32]_not n36206_not ; n36207
g35952 and b[32] n36200_not ; n36208
g35953 and n36205_not n36208 ; n36209
g35954 and n424 n36209_not ; n36210
g35955 and n36207_not n36210 ; n36211
g35956 and n36199_not n36211 ; n36212
g35957 and n432 n36206_not ; n36213
g35958 and n36212_not n36213_not ; n36214
g35959 and n35787_not n36197 ; n36215
g35960 and n36193_not n36215 ; n36216
g35961 and n36194_not n36197_not ; n36217
g35962 and n36216_not n36217_not ; n36218
g35963 and n36214_not n36218_not ; n36219
g35964 and n35777_not n36213_not ; n36220
g35965 and n36212_not n36220 ; n36221
g35966 and n36219_not n36221_not ; n36222
g35967 and n35778_not n36209_not ; n36223
g35968 and n36207_not n36223 ; n36224
g35969 and n36198_not n36224 ; n36225
g35970 and n36207_not n36209_not ; n36226
g35971 and n36199_not n36226_not ; n36227
g35972 and n36225_not n36227_not ; n36228
g35973 and n36214_not n36228_not ; n36229
g35974 and n36206_not n36213_not ; n36230
g35975 and n36212_not n36230 ; n36231
g35976 and n36229_not n36231_not ; n36232
g35977 and b[33]_not n36232_not ; n36233
g35978 and b[32]_not n36222_not ; n36234
g35979 and n35796_not n36192 ; n36235
g35980 and n36188_not n36235 ; n36236
g35981 and n36189_not n36192_not ; n36237
g35982 and n36236_not n36237_not ; n36238
g35983 and n36214_not n36238_not ; n36239
g35984 and n35786_not n36213_not ; n36240
g35985 and n36212_not n36240 ; n36241
g35986 and n36239_not n36241_not ; n36242
g35987 and b[31]_not n36242_not ; n36243
g35988 and n35805_not n36187 ; n36244
g35989 and n36183_not n36244 ; n36245
g35990 and n36184_not n36187_not ; n36246
g35991 and n36245_not n36246_not ; n36247
g35992 and n36214_not n36247_not ; n36248
g35993 and n35795_not n36213_not ; n36249
g35994 and n36212_not n36249 ; n36250
g35995 and n36248_not n36250_not ; n36251
g35996 and b[30]_not n36251_not ; n36252
g35997 and n35814_not n36182 ; n36253
g35998 and n36178_not n36253 ; n36254
g35999 and n36179_not n36182_not ; n36255
g36000 and n36254_not n36255_not ; n36256
g36001 and n36214_not n36256_not ; n36257
g36002 and n35804_not n36213_not ; n36258
g36003 and n36212_not n36258 ; n36259
g36004 and n36257_not n36259_not ; n36260
g36005 and b[29]_not n36260_not ; n36261
g36006 and n35823_not n36177 ; n36262
g36007 and n36173_not n36262 ; n36263
g36008 and n36174_not n36177_not ; n36264
g36009 and n36263_not n36264_not ; n36265
g36010 and n36214_not n36265_not ; n36266
g36011 and n35813_not n36213_not ; n36267
g36012 and n36212_not n36267 ; n36268
g36013 and n36266_not n36268_not ; n36269
g36014 and b[28]_not n36269_not ; n36270
g36015 and n35832_not n36172 ; n36271
g36016 and n36168_not n36271 ; n36272
g36017 and n36169_not n36172_not ; n36273
g36018 and n36272_not n36273_not ; n36274
g36019 and n36214_not n36274_not ; n36275
g36020 and n35822_not n36213_not ; n36276
g36021 and n36212_not n36276 ; n36277
g36022 and n36275_not n36277_not ; n36278
g36023 and b[27]_not n36278_not ; n36279
g36024 and n35841_not n36167 ; n36280
g36025 and n36163_not n36280 ; n36281
g36026 and n36164_not n36167_not ; n36282
g36027 and n36281_not n36282_not ; n36283
g36028 and n36214_not n36283_not ; n36284
g36029 and n35831_not n36213_not ; n36285
g36030 and n36212_not n36285 ; n36286
g36031 and n36284_not n36286_not ; n36287
g36032 and b[26]_not n36287_not ; n36288
g36033 and n35850_not n36162 ; n36289
g36034 and n36158_not n36289 ; n36290
g36035 and n36159_not n36162_not ; n36291
g36036 and n36290_not n36291_not ; n36292
g36037 and n36214_not n36292_not ; n36293
g36038 and n35840_not n36213_not ; n36294
g36039 and n36212_not n36294 ; n36295
g36040 and n36293_not n36295_not ; n36296
g36041 and b[25]_not n36296_not ; n36297
g36042 and n35859_not n36157 ; n36298
g36043 and n36153_not n36298 ; n36299
g36044 and n36154_not n36157_not ; n36300
g36045 and n36299_not n36300_not ; n36301
g36046 and n36214_not n36301_not ; n36302
g36047 and n35849_not n36213_not ; n36303
g36048 and n36212_not n36303 ; n36304
g36049 and n36302_not n36304_not ; n36305
g36050 and b[24]_not n36305_not ; n36306
g36051 and n35868_not n36152 ; n36307
g36052 and n36148_not n36307 ; n36308
g36053 and n36149_not n36152_not ; n36309
g36054 and n36308_not n36309_not ; n36310
g36055 and n36214_not n36310_not ; n36311
g36056 and n35858_not n36213_not ; n36312
g36057 and n36212_not n36312 ; n36313
g36058 and n36311_not n36313_not ; n36314
g36059 and b[23]_not n36314_not ; n36315
g36060 and n35877_not n36147 ; n36316
g36061 and n36143_not n36316 ; n36317
g36062 and n36144_not n36147_not ; n36318
g36063 and n36317_not n36318_not ; n36319
g36064 and n36214_not n36319_not ; n36320
g36065 and n35867_not n36213_not ; n36321
g36066 and n36212_not n36321 ; n36322
g36067 and n36320_not n36322_not ; n36323
g36068 and b[22]_not n36323_not ; n36324
g36069 and n35886_not n36142 ; n36325
g36070 and n36138_not n36325 ; n36326
g36071 and n36139_not n36142_not ; n36327
g36072 and n36326_not n36327_not ; n36328
g36073 and n36214_not n36328_not ; n36329
g36074 and n35876_not n36213_not ; n36330
g36075 and n36212_not n36330 ; n36331
g36076 and n36329_not n36331_not ; n36332
g36077 and b[21]_not n36332_not ; n36333
g36078 and n35895_not n36137 ; n36334
g36079 and n36133_not n36334 ; n36335
g36080 and n36134_not n36137_not ; n36336
g36081 and n36335_not n36336_not ; n36337
g36082 and n36214_not n36337_not ; n36338
g36083 and n35885_not n36213_not ; n36339
g36084 and n36212_not n36339 ; n36340
g36085 and n36338_not n36340_not ; n36341
g36086 and b[20]_not n36341_not ; n36342
g36087 and n35904_not n36132 ; n36343
g36088 and n36128_not n36343 ; n36344
g36089 and n36129_not n36132_not ; n36345
g36090 and n36344_not n36345_not ; n36346
g36091 and n36214_not n36346_not ; n36347
g36092 and n35894_not n36213_not ; n36348
g36093 and n36212_not n36348 ; n36349
g36094 and n36347_not n36349_not ; n36350
g36095 and b[19]_not n36350_not ; n36351
g36096 and n35913_not n36127 ; n36352
g36097 and n36123_not n36352 ; n36353
g36098 and n36124_not n36127_not ; n36354
g36099 and n36353_not n36354_not ; n36355
g36100 and n36214_not n36355_not ; n36356
g36101 and n35903_not n36213_not ; n36357
g36102 and n36212_not n36357 ; n36358
g36103 and n36356_not n36358_not ; n36359
g36104 and b[18]_not n36359_not ; n36360
g36105 and n35922_not n36122 ; n36361
g36106 and n36118_not n36361 ; n36362
g36107 and n36119_not n36122_not ; n36363
g36108 and n36362_not n36363_not ; n36364
g36109 and n36214_not n36364_not ; n36365
g36110 and n35912_not n36213_not ; n36366
g36111 and n36212_not n36366 ; n36367
g36112 and n36365_not n36367_not ; n36368
g36113 and b[17]_not n36368_not ; n36369
g36114 and n35931_not n36117 ; n36370
g36115 and n36113_not n36370 ; n36371
g36116 and n36114_not n36117_not ; n36372
g36117 and n36371_not n36372_not ; n36373
g36118 and n36214_not n36373_not ; n36374
g36119 and n35921_not n36213_not ; n36375
g36120 and n36212_not n36375 ; n36376
g36121 and n36374_not n36376_not ; n36377
g36122 and b[16]_not n36377_not ; n36378
g36123 and n35940_not n36112 ; n36379
g36124 and n36108_not n36379 ; n36380
g36125 and n36109_not n36112_not ; n36381
g36126 and n36380_not n36381_not ; n36382
g36127 and n36214_not n36382_not ; n36383
g36128 and n35930_not n36213_not ; n36384
g36129 and n36212_not n36384 ; n36385
g36130 and n36383_not n36385_not ; n36386
g36131 and b[15]_not n36386_not ; n36387
g36132 and n35949_not n36107 ; n36388
g36133 and n36103_not n36388 ; n36389
g36134 and n36104_not n36107_not ; n36390
g36135 and n36389_not n36390_not ; n36391
g36136 and n36214_not n36391_not ; n36392
g36137 and n35939_not n36213_not ; n36393
g36138 and n36212_not n36393 ; n36394
g36139 and n36392_not n36394_not ; n36395
g36140 and b[14]_not n36395_not ; n36396
g36141 and n35958_not n36102 ; n36397
g36142 and n36098_not n36397 ; n36398
g36143 and n36099_not n36102_not ; n36399
g36144 and n36398_not n36399_not ; n36400
g36145 and n36214_not n36400_not ; n36401
g36146 and n35948_not n36213_not ; n36402
g36147 and n36212_not n36402 ; n36403
g36148 and n36401_not n36403_not ; n36404
g36149 and b[13]_not n36404_not ; n36405
g36150 and n35967_not n36097 ; n36406
g36151 and n36093_not n36406 ; n36407
g36152 and n36094_not n36097_not ; n36408
g36153 and n36407_not n36408_not ; n36409
g36154 and n36214_not n36409_not ; n36410
g36155 and n35957_not n36213_not ; n36411
g36156 and n36212_not n36411 ; n36412
g36157 and n36410_not n36412_not ; n36413
g36158 and b[12]_not n36413_not ; n36414
g36159 and n35976_not n36092 ; n36415
g36160 and n36088_not n36415 ; n36416
g36161 and n36089_not n36092_not ; n36417
g36162 and n36416_not n36417_not ; n36418
g36163 and n36214_not n36418_not ; n36419
g36164 and n35966_not n36213_not ; n36420
g36165 and n36212_not n36420 ; n36421
g36166 and n36419_not n36421_not ; n36422
g36167 and b[11]_not n36422_not ; n36423
g36168 and n35985_not n36087 ; n36424
g36169 and n36083_not n36424 ; n36425
g36170 and n36084_not n36087_not ; n36426
g36171 and n36425_not n36426_not ; n36427
g36172 and n36214_not n36427_not ; n36428
g36173 and n35975_not n36213_not ; n36429
g36174 and n36212_not n36429 ; n36430
g36175 and n36428_not n36430_not ; n36431
g36176 and b[10]_not n36431_not ; n36432
g36177 and n35994_not n36082 ; n36433
g36178 and n36078_not n36433 ; n36434
g36179 and n36079_not n36082_not ; n36435
g36180 and n36434_not n36435_not ; n36436
g36181 and n36214_not n36436_not ; n36437
g36182 and n35984_not n36213_not ; n36438
g36183 and n36212_not n36438 ; n36439
g36184 and n36437_not n36439_not ; n36440
g36185 and b[9]_not n36440_not ; n36441
g36186 and n36003_not n36077 ; n36442
g36187 and n36073_not n36442 ; n36443
g36188 and n36074_not n36077_not ; n36444
g36189 and n36443_not n36444_not ; n36445
g36190 and n36214_not n36445_not ; n36446
g36191 and n35993_not n36213_not ; n36447
g36192 and n36212_not n36447 ; n36448
g36193 and n36446_not n36448_not ; n36449
g36194 and b[8]_not n36449_not ; n36450
g36195 and n36012_not n36072 ; n36451
g36196 and n36068_not n36451 ; n36452
g36197 and n36069_not n36072_not ; n36453
g36198 and n36452_not n36453_not ; n36454
g36199 and n36214_not n36454_not ; n36455
g36200 and n36002_not n36213_not ; n36456
g36201 and n36212_not n36456 ; n36457
g36202 and n36455_not n36457_not ; n36458
g36203 and b[7]_not n36458_not ; n36459
g36204 and n36021_not n36067 ; n36460
g36205 and n36063_not n36460 ; n36461
g36206 and n36064_not n36067_not ; n36462
g36207 and n36461_not n36462_not ; n36463
g36208 and n36214_not n36463_not ; n36464
g36209 and n36011_not n36213_not ; n36465
g36210 and n36212_not n36465 ; n36466
g36211 and n36464_not n36466_not ; n36467
g36212 and b[6]_not n36467_not ; n36468
g36213 and n36030_not n36062 ; n36469
g36214 and n36058_not n36469 ; n36470
g36215 and n36059_not n36062_not ; n36471
g36216 and n36470_not n36471_not ; n36472
g36217 and n36214_not n36472_not ; n36473
g36218 and n36020_not n36213_not ; n36474
g36219 and n36212_not n36474 ; n36475
g36220 and n36473_not n36475_not ; n36476
g36221 and b[5]_not n36476_not ; n36477
g36222 and n36038_not n36057 ; n36478
g36223 and n36053_not n36478 ; n36479
g36224 and n36054_not n36057_not ; n36480
g36225 and n36479_not n36480_not ; n36481
g36226 and n36214_not n36481_not ; n36482
g36227 and n36029_not n36213_not ; n36483
g36228 and n36212_not n36483 ; n36484
g36229 and n36482_not n36484_not ; n36485
g36230 and b[4]_not n36485_not ; n36486
g36231 and n36048_not n36052 ; n36487
g36232 and n36047_not n36487 ; n36488
g36233 and n36049_not n36052_not ; n36489
g36234 and n36488_not n36489_not ; n36490
g36235 and n36214_not n36490_not ; n36491
g36236 and n36037_not n36213_not ; n36492
g36237 and n36212_not n36492 ; n36493
g36238 and n36491_not n36493_not ; n36494
g36239 and b[3]_not n36494_not ; n36495
g36240 and n7887 n36045_not ; n36496
g36241 and n36043_not n36496 ; n36497
g36242 and n36047_not n36497_not ; n36498
g36243 and n36214_not n36498 ; n36499
g36244 and n36042_not n36213_not ; n36500
g36245 and n36212_not n36500 ; n36501
g36246 and n36499_not n36501_not ; n36502
g36247 and b[2]_not n36502_not ; n36503
g36248 and b[0] n36214_not ; n36504
g36249 and a[31] n36504_not ; n36505
g36250 and n7887 n36214_not ; n36506
g36251 and n36505_not n36506_not ; n36507
g36252 and b[1] n36507_not ; n36508
g36253 and b[1]_not n36506_not ; n36509
g36254 and n36505_not n36509 ; n36510
g36255 and n36508_not n36510_not ; n36511
g36256 and n8353_not n36511_not ; n36512
g36257 and b[1]_not n36507_not ; n36513
g36258 and n36512_not n36513_not ; n36514
g36259 and b[2] n36501_not ; n36515
g36260 and n36499_not n36515 ; n36516
g36261 and n36503_not n36516_not ; n36517
g36262 and n36514_not n36517 ; n36518
g36263 and n36503_not n36518_not ; n36519
g36264 and b[3] n36493_not ; n36520
g36265 and n36491_not n36520 ; n36521
g36266 and n36495_not n36521_not ; n36522
g36267 and n36519_not n36522 ; n36523
g36268 and n36495_not n36523_not ; n36524
g36269 and b[4] n36484_not ; n36525
g36270 and n36482_not n36525 ; n36526
g36271 and n36486_not n36526_not ; n36527
g36272 and n36524_not n36527 ; n36528
g36273 and n36486_not n36528_not ; n36529
g36274 and b[5] n36475_not ; n36530
g36275 and n36473_not n36530 ; n36531
g36276 and n36477_not n36531_not ; n36532
g36277 and n36529_not n36532 ; n36533
g36278 and n36477_not n36533_not ; n36534
g36279 and b[6] n36466_not ; n36535
g36280 and n36464_not n36535 ; n36536
g36281 and n36468_not n36536_not ; n36537
g36282 and n36534_not n36537 ; n36538
g36283 and n36468_not n36538_not ; n36539
g36284 and b[7] n36457_not ; n36540
g36285 and n36455_not n36540 ; n36541
g36286 and n36459_not n36541_not ; n36542
g36287 and n36539_not n36542 ; n36543
g36288 and n36459_not n36543_not ; n36544
g36289 and b[8] n36448_not ; n36545
g36290 and n36446_not n36545 ; n36546
g36291 and n36450_not n36546_not ; n36547
g36292 and n36544_not n36547 ; n36548
g36293 and n36450_not n36548_not ; n36549
g36294 and b[9] n36439_not ; n36550
g36295 and n36437_not n36550 ; n36551
g36296 and n36441_not n36551_not ; n36552
g36297 and n36549_not n36552 ; n36553
g36298 and n36441_not n36553_not ; n36554
g36299 and b[10] n36430_not ; n36555
g36300 and n36428_not n36555 ; n36556
g36301 and n36432_not n36556_not ; n36557
g36302 and n36554_not n36557 ; n36558
g36303 and n36432_not n36558_not ; n36559
g36304 and b[11] n36421_not ; n36560
g36305 and n36419_not n36560 ; n36561
g36306 and n36423_not n36561_not ; n36562
g36307 and n36559_not n36562 ; n36563
g36308 and n36423_not n36563_not ; n36564
g36309 and b[12] n36412_not ; n36565
g36310 and n36410_not n36565 ; n36566
g36311 and n36414_not n36566_not ; n36567
g36312 and n36564_not n36567 ; n36568
g36313 and n36414_not n36568_not ; n36569
g36314 and b[13] n36403_not ; n36570
g36315 and n36401_not n36570 ; n36571
g36316 and n36405_not n36571_not ; n36572
g36317 and n36569_not n36572 ; n36573
g36318 and n36405_not n36573_not ; n36574
g36319 and b[14] n36394_not ; n36575
g36320 and n36392_not n36575 ; n36576
g36321 and n36396_not n36576_not ; n36577
g36322 and n36574_not n36577 ; n36578
g36323 and n36396_not n36578_not ; n36579
g36324 and b[15] n36385_not ; n36580
g36325 and n36383_not n36580 ; n36581
g36326 and n36387_not n36581_not ; n36582
g36327 and n36579_not n36582 ; n36583
g36328 and n36387_not n36583_not ; n36584
g36329 and b[16] n36376_not ; n36585
g36330 and n36374_not n36585 ; n36586
g36331 and n36378_not n36586_not ; n36587
g36332 and n36584_not n36587 ; n36588
g36333 and n36378_not n36588_not ; n36589
g36334 and b[17] n36367_not ; n36590
g36335 and n36365_not n36590 ; n36591
g36336 and n36369_not n36591_not ; n36592
g36337 and n36589_not n36592 ; n36593
g36338 and n36369_not n36593_not ; n36594
g36339 and b[18] n36358_not ; n36595
g36340 and n36356_not n36595 ; n36596
g36341 and n36360_not n36596_not ; n36597
g36342 and n36594_not n36597 ; n36598
g36343 and n36360_not n36598_not ; n36599
g36344 and b[19] n36349_not ; n36600
g36345 and n36347_not n36600 ; n36601
g36346 and n36351_not n36601_not ; n36602
g36347 and n36599_not n36602 ; n36603
g36348 and n36351_not n36603_not ; n36604
g36349 and b[20] n36340_not ; n36605
g36350 and n36338_not n36605 ; n36606
g36351 and n36342_not n36606_not ; n36607
g36352 and n36604_not n36607 ; n36608
g36353 and n36342_not n36608_not ; n36609
g36354 and b[21] n36331_not ; n36610
g36355 and n36329_not n36610 ; n36611
g36356 and n36333_not n36611_not ; n36612
g36357 and n36609_not n36612 ; n36613
g36358 and n36333_not n36613_not ; n36614
g36359 and b[22] n36322_not ; n36615
g36360 and n36320_not n36615 ; n36616
g36361 and n36324_not n36616_not ; n36617
g36362 and n36614_not n36617 ; n36618
g36363 and n36324_not n36618_not ; n36619
g36364 and b[23] n36313_not ; n36620
g36365 and n36311_not n36620 ; n36621
g36366 and n36315_not n36621_not ; n36622
g36367 and n36619_not n36622 ; n36623
g36368 and n36315_not n36623_not ; n36624
g36369 and b[24] n36304_not ; n36625
g36370 and n36302_not n36625 ; n36626
g36371 and n36306_not n36626_not ; n36627
g36372 and n36624_not n36627 ; n36628
g36373 and n36306_not n36628_not ; n36629
g36374 and b[25] n36295_not ; n36630
g36375 and n36293_not n36630 ; n36631
g36376 and n36297_not n36631_not ; n36632
g36377 and n36629_not n36632 ; n36633
g36378 and n36297_not n36633_not ; n36634
g36379 and b[26] n36286_not ; n36635
g36380 and n36284_not n36635 ; n36636
g36381 and n36288_not n36636_not ; n36637
g36382 and n36634_not n36637 ; n36638
g36383 and n36288_not n36638_not ; n36639
g36384 and b[27] n36277_not ; n36640
g36385 and n36275_not n36640 ; n36641
g36386 and n36279_not n36641_not ; n36642
g36387 and n36639_not n36642 ; n36643
g36388 and n36279_not n36643_not ; n36644
g36389 and b[28] n36268_not ; n36645
g36390 and n36266_not n36645 ; n36646
g36391 and n36270_not n36646_not ; n36647
g36392 and n36644_not n36647 ; n36648
g36393 and n36270_not n36648_not ; n36649
g36394 and b[29] n36259_not ; n36650
g36395 and n36257_not n36650 ; n36651
g36396 and n36261_not n36651_not ; n36652
g36397 and n36649_not n36652 ; n36653
g36398 and n36261_not n36653_not ; n36654
g36399 and b[30] n36250_not ; n36655
g36400 and n36248_not n36655 ; n36656
g36401 and n36252_not n36656_not ; n36657
g36402 and n36654_not n36657 ; n36658
g36403 and n36252_not n36658_not ; n36659
g36404 and b[31] n36241_not ; n36660
g36405 and n36239_not n36660 ; n36661
g36406 and n36243_not n36661_not ; n36662
g36407 and n36659_not n36662 ; n36663
g36408 and n36243_not n36663_not ; n36664
g36409 and b[32] n36221_not ; n36665
g36410 and n36219_not n36665 ; n36666
g36411 and n36234_not n36666_not ; n36667
g36412 and n36664_not n36667 ; n36668
g36413 and n36234_not n36668_not ; n36669
g36414 and b[33] n36231_not ; n36670
g36415 and n36229_not n36670 ; n36671
g36416 and n36233_not n36671_not ; n36672
g36417 and n36669_not n36672 ; n36673
g36418 and n36233_not n36673_not ; n36674
g36419 and n8519 n36674_not ; n36675
g36420 and n36222_not n36675_not ; n36676
g36421 and n36243_not n36667 ; n36677
g36422 and n36663_not n36677 ; n36678
g36423 and n36664_not n36667_not ; n36679
g36424 and n36678_not n36679_not ; n36680
g36425 and n8519 n36680_not ; n36681
g36426 and n36674_not n36681 ; n36682
g36427 and n36676_not n36682_not ; n36683
g36428 and n36232_not n36675_not ; n36684
g36429 and n36234_not n36672 ; n36685
g36430 and n36668_not n36685 ; n36686
g36431 and n36669_not n36672_not ; n36687
g36432 and n36686_not n36687_not ; n36688
g36433 and n36675 n36688_not ; n36689
g36434 and n36684_not n36689_not ; n36690
g36435 and b[34]_not n36690_not ; n36691
g36436 and b[33]_not n36683_not ; n36692
g36437 and n36242_not n36675_not ; n36693
g36438 and n36252_not n36662 ; n36694
g36439 and n36658_not n36694 ; n36695
g36440 and n36659_not n36662_not ; n36696
g36441 and n36695_not n36696_not ; n36697
g36442 and n8519 n36697_not ; n36698
g36443 and n36674_not n36698 ; n36699
g36444 and n36693_not n36699_not ; n36700
g36445 and b[32]_not n36700_not ; n36701
g36446 and n36251_not n36675_not ; n36702
g36447 and n36261_not n36657 ; n36703
g36448 and n36653_not n36703 ; n36704
g36449 and n36654_not n36657_not ; n36705
g36450 and n36704_not n36705_not ; n36706
g36451 and n8519 n36706_not ; n36707
g36452 and n36674_not n36707 ; n36708
g36453 and n36702_not n36708_not ; n36709
g36454 and b[31]_not n36709_not ; n36710
g36455 and n36260_not n36675_not ; n36711
g36456 and n36270_not n36652 ; n36712
g36457 and n36648_not n36712 ; n36713
g36458 and n36649_not n36652_not ; n36714
g36459 and n36713_not n36714_not ; n36715
g36460 and n8519 n36715_not ; n36716
g36461 and n36674_not n36716 ; n36717
g36462 and n36711_not n36717_not ; n36718
g36463 and b[30]_not n36718_not ; n36719
g36464 and n36269_not n36675_not ; n36720
g36465 and n36279_not n36647 ; n36721
g36466 and n36643_not n36721 ; n36722
g36467 and n36644_not n36647_not ; n36723
g36468 and n36722_not n36723_not ; n36724
g36469 and n8519 n36724_not ; n36725
g36470 and n36674_not n36725 ; n36726
g36471 and n36720_not n36726_not ; n36727
g36472 and b[29]_not n36727_not ; n36728
g36473 and n36278_not n36675_not ; n36729
g36474 and n36288_not n36642 ; n36730
g36475 and n36638_not n36730 ; n36731
g36476 and n36639_not n36642_not ; n36732
g36477 and n36731_not n36732_not ; n36733
g36478 and n8519 n36733_not ; n36734
g36479 and n36674_not n36734 ; n36735
g36480 and n36729_not n36735_not ; n36736
g36481 and b[28]_not n36736_not ; n36737
g36482 and n36287_not n36675_not ; n36738
g36483 and n36297_not n36637 ; n36739
g36484 and n36633_not n36739 ; n36740
g36485 and n36634_not n36637_not ; n36741
g36486 and n36740_not n36741_not ; n36742
g36487 and n8519 n36742_not ; n36743
g36488 and n36674_not n36743 ; n36744
g36489 and n36738_not n36744_not ; n36745
g36490 and b[27]_not n36745_not ; n36746
g36491 and n36296_not n36675_not ; n36747
g36492 and n36306_not n36632 ; n36748
g36493 and n36628_not n36748 ; n36749
g36494 and n36629_not n36632_not ; n36750
g36495 and n36749_not n36750_not ; n36751
g36496 and n8519 n36751_not ; n36752
g36497 and n36674_not n36752 ; n36753
g36498 and n36747_not n36753_not ; n36754
g36499 and b[26]_not n36754_not ; n36755
g36500 and n36305_not n36675_not ; n36756
g36501 and n36315_not n36627 ; n36757
g36502 and n36623_not n36757 ; n36758
g36503 and n36624_not n36627_not ; n36759
g36504 and n36758_not n36759_not ; n36760
g36505 and n8519 n36760_not ; n36761
g36506 and n36674_not n36761 ; n36762
g36507 and n36756_not n36762_not ; n36763
g36508 and b[25]_not n36763_not ; n36764
g36509 and n36314_not n36675_not ; n36765
g36510 and n36324_not n36622 ; n36766
g36511 and n36618_not n36766 ; n36767
g36512 and n36619_not n36622_not ; n36768
g36513 and n36767_not n36768_not ; n36769
g36514 and n8519 n36769_not ; n36770
g36515 and n36674_not n36770 ; n36771
g36516 and n36765_not n36771_not ; n36772
g36517 and b[24]_not n36772_not ; n36773
g36518 and n36323_not n36675_not ; n36774
g36519 and n36333_not n36617 ; n36775
g36520 and n36613_not n36775 ; n36776
g36521 and n36614_not n36617_not ; n36777
g36522 and n36776_not n36777_not ; n36778
g36523 and n8519 n36778_not ; n36779
g36524 and n36674_not n36779 ; n36780
g36525 and n36774_not n36780_not ; n36781
g36526 and b[23]_not n36781_not ; n36782
g36527 and n36332_not n36675_not ; n36783
g36528 and n36342_not n36612 ; n36784
g36529 and n36608_not n36784 ; n36785
g36530 and n36609_not n36612_not ; n36786
g36531 and n36785_not n36786_not ; n36787
g36532 and n8519 n36787_not ; n36788
g36533 and n36674_not n36788 ; n36789
g36534 and n36783_not n36789_not ; n36790
g36535 and b[22]_not n36790_not ; n36791
g36536 and n36341_not n36675_not ; n36792
g36537 and n36351_not n36607 ; n36793
g36538 and n36603_not n36793 ; n36794
g36539 and n36604_not n36607_not ; n36795
g36540 and n36794_not n36795_not ; n36796
g36541 and n8519 n36796_not ; n36797
g36542 and n36674_not n36797 ; n36798
g36543 and n36792_not n36798_not ; n36799
g36544 and b[21]_not n36799_not ; n36800
g36545 and n36350_not n36675_not ; n36801
g36546 and n36360_not n36602 ; n36802
g36547 and n36598_not n36802 ; n36803
g36548 and n36599_not n36602_not ; n36804
g36549 and n36803_not n36804_not ; n36805
g36550 and n8519 n36805_not ; n36806
g36551 and n36674_not n36806 ; n36807
g36552 and n36801_not n36807_not ; n36808
g36553 and b[20]_not n36808_not ; n36809
g36554 and n36359_not n36675_not ; n36810
g36555 and n36369_not n36597 ; n36811
g36556 and n36593_not n36811 ; n36812
g36557 and n36594_not n36597_not ; n36813
g36558 and n36812_not n36813_not ; n36814
g36559 and n8519 n36814_not ; n36815
g36560 and n36674_not n36815 ; n36816
g36561 and n36810_not n36816_not ; n36817
g36562 and b[19]_not n36817_not ; n36818
g36563 and n36368_not n36675_not ; n36819
g36564 and n36378_not n36592 ; n36820
g36565 and n36588_not n36820 ; n36821
g36566 and n36589_not n36592_not ; n36822
g36567 and n36821_not n36822_not ; n36823
g36568 and n8519 n36823_not ; n36824
g36569 and n36674_not n36824 ; n36825
g36570 and n36819_not n36825_not ; n36826
g36571 and b[18]_not n36826_not ; n36827
g36572 and n36377_not n36675_not ; n36828
g36573 and n36387_not n36587 ; n36829
g36574 and n36583_not n36829 ; n36830
g36575 and n36584_not n36587_not ; n36831
g36576 and n36830_not n36831_not ; n36832
g36577 and n8519 n36832_not ; n36833
g36578 and n36674_not n36833 ; n36834
g36579 and n36828_not n36834_not ; n36835
g36580 and b[17]_not n36835_not ; n36836
g36581 and n36386_not n36675_not ; n36837
g36582 and n36396_not n36582 ; n36838
g36583 and n36578_not n36838 ; n36839
g36584 and n36579_not n36582_not ; n36840
g36585 and n36839_not n36840_not ; n36841
g36586 and n8519 n36841_not ; n36842
g36587 and n36674_not n36842 ; n36843
g36588 and n36837_not n36843_not ; n36844
g36589 and b[16]_not n36844_not ; n36845
g36590 and n36395_not n36675_not ; n36846
g36591 and n36405_not n36577 ; n36847
g36592 and n36573_not n36847 ; n36848
g36593 and n36574_not n36577_not ; n36849
g36594 and n36848_not n36849_not ; n36850
g36595 and n8519 n36850_not ; n36851
g36596 and n36674_not n36851 ; n36852
g36597 and n36846_not n36852_not ; n36853
g36598 and b[15]_not n36853_not ; n36854
g36599 and n36404_not n36675_not ; n36855
g36600 and n36414_not n36572 ; n36856
g36601 and n36568_not n36856 ; n36857
g36602 and n36569_not n36572_not ; n36858
g36603 and n36857_not n36858_not ; n36859
g36604 and n8519 n36859_not ; n36860
g36605 and n36674_not n36860 ; n36861
g36606 and n36855_not n36861_not ; n36862
g36607 and b[14]_not n36862_not ; n36863
g36608 and n36413_not n36675_not ; n36864
g36609 and n36423_not n36567 ; n36865
g36610 and n36563_not n36865 ; n36866
g36611 and n36564_not n36567_not ; n36867
g36612 and n36866_not n36867_not ; n36868
g36613 and n8519 n36868_not ; n36869
g36614 and n36674_not n36869 ; n36870
g36615 and n36864_not n36870_not ; n36871
g36616 and b[13]_not n36871_not ; n36872
g36617 and n36422_not n36675_not ; n36873
g36618 and n36432_not n36562 ; n36874
g36619 and n36558_not n36874 ; n36875
g36620 and n36559_not n36562_not ; n36876
g36621 and n36875_not n36876_not ; n36877
g36622 and n8519 n36877_not ; n36878
g36623 and n36674_not n36878 ; n36879
g36624 and n36873_not n36879_not ; n36880
g36625 and b[12]_not n36880_not ; n36881
g36626 and n36431_not n36675_not ; n36882
g36627 and n36441_not n36557 ; n36883
g36628 and n36553_not n36883 ; n36884
g36629 and n36554_not n36557_not ; n36885
g36630 and n36884_not n36885_not ; n36886
g36631 and n8519 n36886_not ; n36887
g36632 and n36674_not n36887 ; n36888
g36633 and n36882_not n36888_not ; n36889
g36634 and b[11]_not n36889_not ; n36890
g36635 and n36440_not n36675_not ; n36891
g36636 and n36450_not n36552 ; n36892
g36637 and n36548_not n36892 ; n36893
g36638 and n36549_not n36552_not ; n36894
g36639 and n36893_not n36894_not ; n36895
g36640 and n8519 n36895_not ; n36896
g36641 and n36674_not n36896 ; n36897
g36642 and n36891_not n36897_not ; n36898
g36643 and b[10]_not n36898_not ; n36899
g36644 and n36449_not n36675_not ; n36900
g36645 and n36459_not n36547 ; n36901
g36646 and n36543_not n36901 ; n36902
g36647 and n36544_not n36547_not ; n36903
g36648 and n36902_not n36903_not ; n36904
g36649 and n8519 n36904_not ; n36905
g36650 and n36674_not n36905 ; n36906
g36651 and n36900_not n36906_not ; n36907
g36652 and b[9]_not n36907_not ; n36908
g36653 and n36458_not n36675_not ; n36909
g36654 and n36468_not n36542 ; n36910
g36655 and n36538_not n36910 ; n36911
g36656 and n36539_not n36542_not ; n36912
g36657 and n36911_not n36912_not ; n36913
g36658 and n8519 n36913_not ; n36914
g36659 and n36674_not n36914 ; n36915
g36660 and n36909_not n36915_not ; n36916
g36661 and b[8]_not n36916_not ; n36917
g36662 and n36467_not n36675_not ; n36918
g36663 and n36477_not n36537 ; n36919
g36664 and n36533_not n36919 ; n36920
g36665 and n36534_not n36537_not ; n36921
g36666 and n36920_not n36921_not ; n36922
g36667 and n8519 n36922_not ; n36923
g36668 and n36674_not n36923 ; n36924
g36669 and n36918_not n36924_not ; n36925
g36670 and b[7]_not n36925_not ; n36926
g36671 and n36476_not n36675_not ; n36927
g36672 and n36486_not n36532 ; n36928
g36673 and n36528_not n36928 ; n36929
g36674 and n36529_not n36532_not ; n36930
g36675 and n36929_not n36930_not ; n36931
g36676 and n8519 n36931_not ; n36932
g36677 and n36674_not n36932 ; n36933
g36678 and n36927_not n36933_not ; n36934
g36679 and b[6]_not n36934_not ; n36935
g36680 and n36485_not n36675_not ; n36936
g36681 and n36495_not n36527 ; n36937
g36682 and n36523_not n36937 ; n36938
g36683 and n36524_not n36527_not ; n36939
g36684 and n36938_not n36939_not ; n36940
g36685 and n8519 n36940_not ; n36941
g36686 and n36674_not n36941 ; n36942
g36687 and n36936_not n36942_not ; n36943
g36688 and b[5]_not n36943_not ; n36944
g36689 and n36494_not n36675_not ; n36945
g36690 and n36503_not n36522 ; n36946
g36691 and n36518_not n36946 ; n36947
g36692 and n36519_not n36522_not ; n36948
g36693 and n36947_not n36948_not ; n36949
g36694 and n8519 n36949_not ; n36950
g36695 and n36674_not n36950 ; n36951
g36696 and n36945_not n36951_not ; n36952
g36697 and b[4]_not n36952_not ; n36953
g36698 and n36502_not n36675_not ; n36954
g36699 and n36513_not n36517 ; n36955
g36700 and n36512_not n36955 ; n36956
g36701 and n36514_not n36517_not ; n36957
g36702 and n36956_not n36957_not ; n36958
g36703 and n8519 n36958_not ; n36959
g36704 and n36674_not n36959 ; n36960
g36705 and n36954_not n36960_not ; n36961
g36706 and b[3]_not n36961_not ; n36962
g36707 and n36507_not n36675_not ; n36963
g36708 and n8353 n36510_not ; n36964
g36709 and n36508_not n36964 ; n36965
g36710 and n8519 n36965_not ; n36966
g36711 and n36512_not n36966 ; n36967
g36712 and n36674_not n36967 ; n36968
g36713 and n36963_not n36968_not ; n36969
g36714 and b[2]_not n36969_not ; n36970
g36715 and n8820 n36674_not ; n36971
g36716 and a[30] n36971_not ; n36972
g36717 and n8826 n36674_not ; n36973
g36718 and n36972_not n36973_not ; n36974
g36719 and b[1] n36974_not ; n36975
g36720 and b[1]_not n36973_not ; n36976
g36721 and n36972_not n36976 ; n36977
g36722 and n36975_not n36977_not ; n36978
g36723 and n8833_not n36978_not ; n36979
g36724 and b[1]_not n36974_not ; n36980
g36725 and n36979_not n36980_not ; n36981
g36726 and b[2] n36968_not ; n36982
g36727 and n36963_not n36982 ; n36983
g36728 and n36970_not n36983_not ; n36984
g36729 and n36981_not n36984 ; n36985
g36730 and n36970_not n36985_not ; n36986
g36731 and b[3] n36960_not ; n36987
g36732 and n36954_not n36987 ; n36988
g36733 and n36962_not n36988_not ; n36989
g36734 and n36986_not n36989 ; n36990
g36735 and n36962_not n36990_not ; n36991
g36736 and b[4] n36951_not ; n36992
g36737 and n36945_not n36992 ; n36993
g36738 and n36953_not n36993_not ; n36994
g36739 and n36991_not n36994 ; n36995
g36740 and n36953_not n36995_not ; n36996
g36741 and b[5] n36942_not ; n36997
g36742 and n36936_not n36997 ; n36998
g36743 and n36944_not n36998_not ; n36999
g36744 and n36996_not n36999 ; n37000
g36745 and n36944_not n37000_not ; n37001
g36746 and b[6] n36933_not ; n37002
g36747 and n36927_not n37002 ; n37003
g36748 and n36935_not n37003_not ; n37004
g36749 and n37001_not n37004 ; n37005
g36750 and n36935_not n37005_not ; n37006
g36751 and b[7] n36924_not ; n37007
g36752 and n36918_not n37007 ; n37008
g36753 and n36926_not n37008_not ; n37009
g36754 and n37006_not n37009 ; n37010
g36755 and n36926_not n37010_not ; n37011
g36756 and b[8] n36915_not ; n37012
g36757 and n36909_not n37012 ; n37013
g36758 and n36917_not n37013_not ; n37014
g36759 and n37011_not n37014 ; n37015
g36760 and n36917_not n37015_not ; n37016
g36761 and b[9] n36906_not ; n37017
g36762 and n36900_not n37017 ; n37018
g36763 and n36908_not n37018_not ; n37019
g36764 and n37016_not n37019 ; n37020
g36765 and n36908_not n37020_not ; n37021
g36766 and b[10] n36897_not ; n37022
g36767 and n36891_not n37022 ; n37023
g36768 and n36899_not n37023_not ; n37024
g36769 and n37021_not n37024 ; n37025
g36770 and n36899_not n37025_not ; n37026
g36771 and b[11] n36888_not ; n37027
g36772 and n36882_not n37027 ; n37028
g36773 and n36890_not n37028_not ; n37029
g36774 and n37026_not n37029 ; n37030
g36775 and n36890_not n37030_not ; n37031
g36776 and b[12] n36879_not ; n37032
g36777 and n36873_not n37032 ; n37033
g36778 and n36881_not n37033_not ; n37034
g36779 and n37031_not n37034 ; n37035
g36780 and n36881_not n37035_not ; n37036
g36781 and b[13] n36870_not ; n37037
g36782 and n36864_not n37037 ; n37038
g36783 and n36872_not n37038_not ; n37039
g36784 and n37036_not n37039 ; n37040
g36785 and n36872_not n37040_not ; n37041
g36786 and b[14] n36861_not ; n37042
g36787 and n36855_not n37042 ; n37043
g36788 and n36863_not n37043_not ; n37044
g36789 and n37041_not n37044 ; n37045
g36790 and n36863_not n37045_not ; n37046
g36791 and b[15] n36852_not ; n37047
g36792 and n36846_not n37047 ; n37048
g36793 and n36854_not n37048_not ; n37049
g36794 and n37046_not n37049 ; n37050
g36795 and n36854_not n37050_not ; n37051
g36796 and b[16] n36843_not ; n37052
g36797 and n36837_not n37052 ; n37053
g36798 and n36845_not n37053_not ; n37054
g36799 and n37051_not n37054 ; n37055
g36800 and n36845_not n37055_not ; n37056
g36801 and b[17] n36834_not ; n37057
g36802 and n36828_not n37057 ; n37058
g36803 and n36836_not n37058_not ; n37059
g36804 and n37056_not n37059 ; n37060
g36805 and n36836_not n37060_not ; n37061
g36806 and b[18] n36825_not ; n37062
g36807 and n36819_not n37062 ; n37063
g36808 and n36827_not n37063_not ; n37064
g36809 and n37061_not n37064 ; n37065
g36810 and n36827_not n37065_not ; n37066
g36811 and b[19] n36816_not ; n37067
g36812 and n36810_not n37067 ; n37068
g36813 and n36818_not n37068_not ; n37069
g36814 and n37066_not n37069 ; n37070
g36815 and n36818_not n37070_not ; n37071
g36816 and b[20] n36807_not ; n37072
g36817 and n36801_not n37072 ; n37073
g36818 and n36809_not n37073_not ; n37074
g36819 and n37071_not n37074 ; n37075
g36820 and n36809_not n37075_not ; n37076
g36821 and b[21] n36798_not ; n37077
g36822 and n36792_not n37077 ; n37078
g36823 and n36800_not n37078_not ; n37079
g36824 and n37076_not n37079 ; n37080
g36825 and n36800_not n37080_not ; n37081
g36826 and b[22] n36789_not ; n37082
g36827 and n36783_not n37082 ; n37083
g36828 and n36791_not n37083_not ; n37084
g36829 and n37081_not n37084 ; n37085
g36830 and n36791_not n37085_not ; n37086
g36831 and b[23] n36780_not ; n37087
g36832 and n36774_not n37087 ; n37088
g36833 and n36782_not n37088_not ; n37089
g36834 and n37086_not n37089 ; n37090
g36835 and n36782_not n37090_not ; n37091
g36836 and b[24] n36771_not ; n37092
g36837 and n36765_not n37092 ; n37093
g36838 and n36773_not n37093_not ; n37094
g36839 and n37091_not n37094 ; n37095
g36840 and n36773_not n37095_not ; n37096
g36841 and b[25] n36762_not ; n37097
g36842 and n36756_not n37097 ; n37098
g36843 and n36764_not n37098_not ; n37099
g36844 and n37096_not n37099 ; n37100
g36845 and n36764_not n37100_not ; n37101
g36846 and b[26] n36753_not ; n37102
g36847 and n36747_not n37102 ; n37103
g36848 and n36755_not n37103_not ; n37104
g36849 and n37101_not n37104 ; n37105
g36850 and n36755_not n37105_not ; n37106
g36851 and b[27] n36744_not ; n37107
g36852 and n36738_not n37107 ; n37108
g36853 and n36746_not n37108_not ; n37109
g36854 and n37106_not n37109 ; n37110
g36855 and n36746_not n37110_not ; n37111
g36856 and b[28] n36735_not ; n37112
g36857 and n36729_not n37112 ; n37113
g36858 and n36737_not n37113_not ; n37114
g36859 and n37111_not n37114 ; n37115
g36860 and n36737_not n37115_not ; n37116
g36861 and b[29] n36726_not ; n37117
g36862 and n36720_not n37117 ; n37118
g36863 and n36728_not n37118_not ; n37119
g36864 and n37116_not n37119 ; n37120
g36865 and n36728_not n37120_not ; n37121
g36866 and b[30] n36717_not ; n37122
g36867 and n36711_not n37122 ; n37123
g36868 and n36719_not n37123_not ; n37124
g36869 and n37121_not n37124 ; n37125
g36870 and n36719_not n37125_not ; n37126
g36871 and b[31] n36708_not ; n37127
g36872 and n36702_not n37127 ; n37128
g36873 and n36710_not n37128_not ; n37129
g36874 and n37126_not n37129 ; n37130
g36875 and n36710_not n37130_not ; n37131
g36876 and b[32] n36699_not ; n37132
g36877 and n36693_not n37132 ; n37133
g36878 and n36701_not n37133_not ; n37134
g36879 and n37131_not n37134 ; n37135
g36880 and n36701_not n37135_not ; n37136
g36881 and b[33] n36682_not ; n37137
g36882 and n36676_not n37137 ; n37138
g36883 and n36692_not n37138_not ; n37139
g36884 and n37136_not n37139 ; n37140
g36885 and n36692_not n37140_not ; n37141
g36886 and b[34] n36684_not ; n37142
g36887 and n36689_not n37142 ; n37143
g36888 and n36691_not n37143_not ; n37144
g36889 and n37141_not n37144 ; n37145
g36890 and n36691_not n37145_not ; n37146
g36891 and n9004 n37146_not ; n37147
g36892 and n36683_not n37147_not ; n37148
g36893 and n36701_not n37139 ; n37149
g36894 and n37135_not n37149 ; n37150
g36895 and n37136_not n37139_not ; n37151
g36896 and n37150_not n37151_not ; n37152
g36897 and n9004 n37152_not ; n37153
g36898 and n37146_not n37153 ; n37154
g36899 and n37148_not n37154_not ; n37155
g36900 and b[34]_not n37155_not ; n37156
g36901 and n36700_not n37147_not ; n37157
g36902 and n36710_not n37134 ; n37158
g36903 and n37130_not n37158 ; n37159
g36904 and n37131_not n37134_not ; n37160
g36905 and n37159_not n37160_not ; n37161
g36906 and n9004 n37161_not ; n37162
g36907 and n37146_not n37162 ; n37163
g36908 and n37157_not n37163_not ; n37164
g36909 and b[33]_not n37164_not ; n37165
g36910 and n36709_not n37147_not ; n37166
g36911 and n36719_not n37129 ; n37167
g36912 and n37125_not n37167 ; n37168
g36913 and n37126_not n37129_not ; n37169
g36914 and n37168_not n37169_not ; n37170
g36915 and n9004 n37170_not ; n37171
g36916 and n37146_not n37171 ; n37172
g36917 and n37166_not n37172_not ; n37173
g36918 and b[32]_not n37173_not ; n37174
g36919 and n36718_not n37147_not ; n37175
g36920 and n36728_not n37124 ; n37176
g36921 and n37120_not n37176 ; n37177
g36922 and n37121_not n37124_not ; n37178
g36923 and n37177_not n37178_not ; n37179
g36924 and n9004 n37179_not ; n37180
g36925 and n37146_not n37180 ; n37181
g36926 and n37175_not n37181_not ; n37182
g36927 and b[31]_not n37182_not ; n37183
g36928 and n36727_not n37147_not ; n37184
g36929 and n36737_not n37119 ; n37185
g36930 and n37115_not n37185 ; n37186
g36931 and n37116_not n37119_not ; n37187
g36932 and n37186_not n37187_not ; n37188
g36933 and n9004 n37188_not ; n37189
g36934 and n37146_not n37189 ; n37190
g36935 and n37184_not n37190_not ; n37191
g36936 and b[30]_not n37191_not ; n37192
g36937 and n36736_not n37147_not ; n37193
g36938 and n36746_not n37114 ; n37194
g36939 and n37110_not n37194 ; n37195
g36940 and n37111_not n37114_not ; n37196
g36941 and n37195_not n37196_not ; n37197
g36942 and n9004 n37197_not ; n37198
g36943 and n37146_not n37198 ; n37199
g36944 and n37193_not n37199_not ; n37200
g36945 and b[29]_not n37200_not ; n37201
g36946 and n36745_not n37147_not ; n37202
g36947 and n36755_not n37109 ; n37203
g36948 and n37105_not n37203 ; n37204
g36949 and n37106_not n37109_not ; n37205
g36950 and n37204_not n37205_not ; n37206
g36951 and n9004 n37206_not ; n37207
g36952 and n37146_not n37207 ; n37208
g36953 and n37202_not n37208_not ; n37209
g36954 and b[28]_not n37209_not ; n37210
g36955 and n36754_not n37147_not ; n37211
g36956 and n36764_not n37104 ; n37212
g36957 and n37100_not n37212 ; n37213
g36958 and n37101_not n37104_not ; n37214
g36959 and n37213_not n37214_not ; n37215
g36960 and n9004 n37215_not ; n37216
g36961 and n37146_not n37216 ; n37217
g36962 and n37211_not n37217_not ; n37218
g36963 and b[27]_not n37218_not ; n37219
g36964 and n36763_not n37147_not ; n37220
g36965 and n36773_not n37099 ; n37221
g36966 and n37095_not n37221 ; n37222
g36967 and n37096_not n37099_not ; n37223
g36968 and n37222_not n37223_not ; n37224
g36969 and n9004 n37224_not ; n37225
g36970 and n37146_not n37225 ; n37226
g36971 and n37220_not n37226_not ; n37227
g36972 and b[26]_not n37227_not ; n37228
g36973 and n36772_not n37147_not ; n37229
g36974 and n36782_not n37094 ; n37230
g36975 and n37090_not n37230 ; n37231
g36976 and n37091_not n37094_not ; n37232
g36977 and n37231_not n37232_not ; n37233
g36978 and n9004 n37233_not ; n37234
g36979 and n37146_not n37234 ; n37235
g36980 and n37229_not n37235_not ; n37236
g36981 and b[25]_not n37236_not ; n37237
g36982 and n36781_not n37147_not ; n37238
g36983 and n36791_not n37089 ; n37239
g36984 and n37085_not n37239 ; n37240
g36985 and n37086_not n37089_not ; n37241
g36986 and n37240_not n37241_not ; n37242
g36987 and n9004 n37242_not ; n37243
g36988 and n37146_not n37243 ; n37244
g36989 and n37238_not n37244_not ; n37245
g36990 and b[24]_not n37245_not ; n37246
g36991 and n36790_not n37147_not ; n37247
g36992 and n36800_not n37084 ; n37248
g36993 and n37080_not n37248 ; n37249
g36994 and n37081_not n37084_not ; n37250
g36995 and n37249_not n37250_not ; n37251
g36996 and n9004 n37251_not ; n37252
g36997 and n37146_not n37252 ; n37253
g36998 and n37247_not n37253_not ; n37254
g36999 and b[23]_not n37254_not ; n37255
g37000 and n36799_not n37147_not ; n37256
g37001 and n36809_not n37079 ; n37257
g37002 and n37075_not n37257 ; n37258
g37003 and n37076_not n37079_not ; n37259
g37004 and n37258_not n37259_not ; n37260
g37005 and n9004 n37260_not ; n37261
g37006 and n37146_not n37261 ; n37262
g37007 and n37256_not n37262_not ; n37263
g37008 and b[22]_not n37263_not ; n37264
g37009 and n36808_not n37147_not ; n37265
g37010 and n36818_not n37074 ; n37266
g37011 and n37070_not n37266 ; n37267
g37012 and n37071_not n37074_not ; n37268
g37013 and n37267_not n37268_not ; n37269
g37014 and n9004 n37269_not ; n37270
g37015 and n37146_not n37270 ; n37271
g37016 and n37265_not n37271_not ; n37272
g37017 and b[21]_not n37272_not ; n37273
g37018 and n36817_not n37147_not ; n37274
g37019 and n36827_not n37069 ; n37275
g37020 and n37065_not n37275 ; n37276
g37021 and n37066_not n37069_not ; n37277
g37022 and n37276_not n37277_not ; n37278
g37023 and n9004 n37278_not ; n37279
g37024 and n37146_not n37279 ; n37280
g37025 and n37274_not n37280_not ; n37281
g37026 and b[20]_not n37281_not ; n37282
g37027 and n36826_not n37147_not ; n37283
g37028 and n36836_not n37064 ; n37284
g37029 and n37060_not n37284 ; n37285
g37030 and n37061_not n37064_not ; n37286
g37031 and n37285_not n37286_not ; n37287
g37032 and n9004 n37287_not ; n37288
g37033 and n37146_not n37288 ; n37289
g37034 and n37283_not n37289_not ; n37290
g37035 and b[19]_not n37290_not ; n37291
g37036 and n36835_not n37147_not ; n37292
g37037 and n36845_not n37059 ; n37293
g37038 and n37055_not n37293 ; n37294
g37039 and n37056_not n37059_not ; n37295
g37040 and n37294_not n37295_not ; n37296
g37041 and n9004 n37296_not ; n37297
g37042 and n37146_not n37297 ; n37298
g37043 and n37292_not n37298_not ; n37299
g37044 and b[18]_not n37299_not ; n37300
g37045 and n36844_not n37147_not ; n37301
g37046 and n36854_not n37054 ; n37302
g37047 and n37050_not n37302 ; n37303
g37048 and n37051_not n37054_not ; n37304
g37049 and n37303_not n37304_not ; n37305
g37050 and n9004 n37305_not ; n37306
g37051 and n37146_not n37306 ; n37307
g37052 and n37301_not n37307_not ; n37308
g37053 and b[17]_not n37308_not ; n37309
g37054 and n36853_not n37147_not ; n37310
g37055 and n36863_not n37049 ; n37311
g37056 and n37045_not n37311 ; n37312
g37057 and n37046_not n37049_not ; n37313
g37058 and n37312_not n37313_not ; n37314
g37059 and n9004 n37314_not ; n37315
g37060 and n37146_not n37315 ; n37316
g37061 and n37310_not n37316_not ; n37317
g37062 and b[16]_not n37317_not ; n37318
g37063 and n36862_not n37147_not ; n37319
g37064 and n36872_not n37044 ; n37320
g37065 and n37040_not n37320 ; n37321
g37066 and n37041_not n37044_not ; n37322
g37067 and n37321_not n37322_not ; n37323
g37068 and n9004 n37323_not ; n37324
g37069 and n37146_not n37324 ; n37325
g37070 and n37319_not n37325_not ; n37326
g37071 and b[15]_not n37326_not ; n37327
g37072 and n36871_not n37147_not ; n37328
g37073 and n36881_not n37039 ; n37329
g37074 and n37035_not n37329 ; n37330
g37075 and n37036_not n37039_not ; n37331
g37076 and n37330_not n37331_not ; n37332
g37077 and n9004 n37332_not ; n37333
g37078 and n37146_not n37333 ; n37334
g37079 and n37328_not n37334_not ; n37335
g37080 and b[14]_not n37335_not ; n37336
g37081 and n36880_not n37147_not ; n37337
g37082 and n36890_not n37034 ; n37338
g37083 and n37030_not n37338 ; n37339
g37084 and n37031_not n37034_not ; n37340
g37085 and n37339_not n37340_not ; n37341
g37086 and n9004 n37341_not ; n37342
g37087 and n37146_not n37342 ; n37343
g37088 and n37337_not n37343_not ; n37344
g37089 and b[13]_not n37344_not ; n37345
g37090 and n36889_not n37147_not ; n37346
g37091 and n36899_not n37029 ; n37347
g37092 and n37025_not n37347 ; n37348
g37093 and n37026_not n37029_not ; n37349
g37094 and n37348_not n37349_not ; n37350
g37095 and n9004 n37350_not ; n37351
g37096 and n37146_not n37351 ; n37352
g37097 and n37346_not n37352_not ; n37353
g37098 and b[12]_not n37353_not ; n37354
g37099 and n36898_not n37147_not ; n37355
g37100 and n36908_not n37024 ; n37356
g37101 and n37020_not n37356 ; n37357
g37102 and n37021_not n37024_not ; n37358
g37103 and n37357_not n37358_not ; n37359
g37104 and n9004 n37359_not ; n37360
g37105 and n37146_not n37360 ; n37361
g37106 and n37355_not n37361_not ; n37362
g37107 and b[11]_not n37362_not ; n37363
g37108 and n36907_not n37147_not ; n37364
g37109 and n36917_not n37019 ; n37365
g37110 and n37015_not n37365 ; n37366
g37111 and n37016_not n37019_not ; n37367
g37112 and n37366_not n37367_not ; n37368
g37113 and n9004 n37368_not ; n37369
g37114 and n37146_not n37369 ; n37370
g37115 and n37364_not n37370_not ; n37371
g37116 and b[10]_not n37371_not ; n37372
g37117 and n36916_not n37147_not ; n37373
g37118 and n36926_not n37014 ; n37374
g37119 and n37010_not n37374 ; n37375
g37120 and n37011_not n37014_not ; n37376
g37121 and n37375_not n37376_not ; n37377
g37122 and n9004 n37377_not ; n37378
g37123 and n37146_not n37378 ; n37379
g37124 and n37373_not n37379_not ; n37380
g37125 and b[9]_not n37380_not ; n37381
g37126 and n36925_not n37147_not ; n37382
g37127 and n36935_not n37009 ; n37383
g37128 and n37005_not n37383 ; n37384
g37129 and n37006_not n37009_not ; n37385
g37130 and n37384_not n37385_not ; n37386
g37131 and n9004 n37386_not ; n37387
g37132 and n37146_not n37387 ; n37388
g37133 and n37382_not n37388_not ; n37389
g37134 and b[8]_not n37389_not ; n37390
g37135 and n36934_not n37147_not ; n37391
g37136 and n36944_not n37004 ; n37392
g37137 and n37000_not n37392 ; n37393
g37138 and n37001_not n37004_not ; n37394
g37139 and n37393_not n37394_not ; n37395
g37140 and n9004 n37395_not ; n37396
g37141 and n37146_not n37396 ; n37397
g37142 and n37391_not n37397_not ; n37398
g37143 and b[7]_not n37398_not ; n37399
g37144 and n36943_not n37147_not ; n37400
g37145 and n36953_not n36999 ; n37401
g37146 and n36995_not n37401 ; n37402
g37147 and n36996_not n36999_not ; n37403
g37148 and n37402_not n37403_not ; n37404
g37149 and n9004 n37404_not ; n37405
g37150 and n37146_not n37405 ; n37406
g37151 and n37400_not n37406_not ; n37407
g37152 and b[6]_not n37407_not ; n37408
g37153 and n36952_not n37147_not ; n37409
g37154 and n36962_not n36994 ; n37410
g37155 and n36990_not n37410 ; n37411
g37156 and n36991_not n36994_not ; n37412
g37157 and n37411_not n37412_not ; n37413
g37158 and n9004 n37413_not ; n37414
g37159 and n37146_not n37414 ; n37415
g37160 and n37409_not n37415_not ; n37416
g37161 and b[5]_not n37416_not ; n37417
g37162 and n36961_not n37147_not ; n37418
g37163 and n36970_not n36989 ; n37419
g37164 and n36985_not n37419 ; n37420
g37165 and n36986_not n36989_not ; n37421
g37166 and n37420_not n37421_not ; n37422
g37167 and n9004 n37422_not ; n37423
g37168 and n37146_not n37423 ; n37424
g37169 and n37418_not n37424_not ; n37425
g37170 and b[4]_not n37425_not ; n37426
g37171 and n36969_not n37147_not ; n37427
g37172 and n36980_not n36984 ; n37428
g37173 and n36979_not n37428 ; n37429
g37174 and n36981_not n36984_not ; n37430
g37175 and n37429_not n37430_not ; n37431
g37176 and n9004 n37431_not ; n37432
g37177 and n37146_not n37432 ; n37433
g37178 and n37427_not n37433_not ; n37434
g37179 and b[3]_not n37434_not ; n37435
g37180 and n36974_not n37147_not ; n37436
g37181 and n8833 n36977_not ; n37437
g37182 and n36975_not n37437 ; n37438
g37183 and n9004 n37438_not ; n37439
g37184 and n36979_not n37439 ; n37440
g37185 and n37146_not n37440 ; n37441
g37186 and n37436_not n37441_not ; n37442
g37187 and b[2]_not n37442_not ; n37443
g37188 and n9305 n37146_not ; n37444
g37189 and a[29] n37444_not ; n37445
g37190 and n9311 n37146_not ; n37446
g37191 and n37445_not n37446_not ; n37447
g37192 and b[1] n37447_not ; n37448
g37193 and b[1]_not n37446_not ; n37449
g37194 and n37445_not n37449 ; n37450
g37195 and n37448_not n37450_not ; n37451
g37196 and n9318_not n37451_not ; n37452
g37197 and b[1]_not n37447_not ; n37453
g37198 and n37452_not n37453_not ; n37454
g37199 and b[2] n37441_not ; n37455
g37200 and n37436_not n37455 ; n37456
g37201 and n37443_not n37456_not ; n37457
g37202 and n37454_not n37457 ; n37458
g37203 and n37443_not n37458_not ; n37459
g37204 and b[3] n37433_not ; n37460
g37205 and n37427_not n37460 ; n37461
g37206 and n37435_not n37461_not ; n37462
g37207 and n37459_not n37462 ; n37463
g37208 and n37435_not n37463_not ; n37464
g37209 and b[4] n37424_not ; n37465
g37210 and n37418_not n37465 ; n37466
g37211 and n37426_not n37466_not ; n37467
g37212 and n37464_not n37467 ; n37468
g37213 and n37426_not n37468_not ; n37469
g37214 and b[5] n37415_not ; n37470
g37215 and n37409_not n37470 ; n37471
g37216 and n37417_not n37471_not ; n37472
g37217 and n37469_not n37472 ; n37473
g37218 and n37417_not n37473_not ; n37474
g37219 and b[6] n37406_not ; n37475
g37220 and n37400_not n37475 ; n37476
g37221 and n37408_not n37476_not ; n37477
g37222 and n37474_not n37477 ; n37478
g37223 and n37408_not n37478_not ; n37479
g37224 and b[7] n37397_not ; n37480
g37225 and n37391_not n37480 ; n37481
g37226 and n37399_not n37481_not ; n37482
g37227 and n37479_not n37482 ; n37483
g37228 and n37399_not n37483_not ; n37484
g37229 and b[8] n37388_not ; n37485
g37230 and n37382_not n37485 ; n37486
g37231 and n37390_not n37486_not ; n37487
g37232 and n37484_not n37487 ; n37488
g37233 and n37390_not n37488_not ; n37489
g37234 and b[9] n37379_not ; n37490
g37235 and n37373_not n37490 ; n37491
g37236 and n37381_not n37491_not ; n37492
g37237 and n37489_not n37492 ; n37493
g37238 and n37381_not n37493_not ; n37494
g37239 and b[10] n37370_not ; n37495
g37240 and n37364_not n37495 ; n37496
g37241 and n37372_not n37496_not ; n37497
g37242 and n37494_not n37497 ; n37498
g37243 and n37372_not n37498_not ; n37499
g37244 and b[11] n37361_not ; n37500
g37245 and n37355_not n37500 ; n37501
g37246 and n37363_not n37501_not ; n37502
g37247 and n37499_not n37502 ; n37503
g37248 and n37363_not n37503_not ; n37504
g37249 and b[12] n37352_not ; n37505
g37250 and n37346_not n37505 ; n37506
g37251 and n37354_not n37506_not ; n37507
g37252 and n37504_not n37507 ; n37508
g37253 and n37354_not n37508_not ; n37509
g37254 and b[13] n37343_not ; n37510
g37255 and n37337_not n37510 ; n37511
g37256 and n37345_not n37511_not ; n37512
g37257 and n37509_not n37512 ; n37513
g37258 and n37345_not n37513_not ; n37514
g37259 and b[14] n37334_not ; n37515
g37260 and n37328_not n37515 ; n37516
g37261 and n37336_not n37516_not ; n37517
g37262 and n37514_not n37517 ; n37518
g37263 and n37336_not n37518_not ; n37519
g37264 and b[15] n37325_not ; n37520
g37265 and n37319_not n37520 ; n37521
g37266 and n37327_not n37521_not ; n37522
g37267 and n37519_not n37522 ; n37523
g37268 and n37327_not n37523_not ; n37524
g37269 and b[16] n37316_not ; n37525
g37270 and n37310_not n37525 ; n37526
g37271 and n37318_not n37526_not ; n37527
g37272 and n37524_not n37527 ; n37528
g37273 and n37318_not n37528_not ; n37529
g37274 and b[17] n37307_not ; n37530
g37275 and n37301_not n37530 ; n37531
g37276 and n37309_not n37531_not ; n37532
g37277 and n37529_not n37532 ; n37533
g37278 and n37309_not n37533_not ; n37534
g37279 and b[18] n37298_not ; n37535
g37280 and n37292_not n37535 ; n37536
g37281 and n37300_not n37536_not ; n37537
g37282 and n37534_not n37537 ; n37538
g37283 and n37300_not n37538_not ; n37539
g37284 and b[19] n37289_not ; n37540
g37285 and n37283_not n37540 ; n37541
g37286 and n37291_not n37541_not ; n37542
g37287 and n37539_not n37542 ; n37543
g37288 and n37291_not n37543_not ; n37544
g37289 and b[20] n37280_not ; n37545
g37290 and n37274_not n37545 ; n37546
g37291 and n37282_not n37546_not ; n37547
g37292 and n37544_not n37547 ; n37548
g37293 and n37282_not n37548_not ; n37549
g37294 and b[21] n37271_not ; n37550
g37295 and n37265_not n37550 ; n37551
g37296 and n37273_not n37551_not ; n37552
g37297 and n37549_not n37552 ; n37553
g37298 and n37273_not n37553_not ; n37554
g37299 and b[22] n37262_not ; n37555
g37300 and n37256_not n37555 ; n37556
g37301 and n37264_not n37556_not ; n37557
g37302 and n37554_not n37557 ; n37558
g37303 and n37264_not n37558_not ; n37559
g37304 and b[23] n37253_not ; n37560
g37305 and n37247_not n37560 ; n37561
g37306 and n37255_not n37561_not ; n37562
g37307 and n37559_not n37562 ; n37563
g37308 and n37255_not n37563_not ; n37564
g37309 and b[24] n37244_not ; n37565
g37310 and n37238_not n37565 ; n37566
g37311 and n37246_not n37566_not ; n37567
g37312 and n37564_not n37567 ; n37568
g37313 and n37246_not n37568_not ; n37569
g37314 and b[25] n37235_not ; n37570
g37315 and n37229_not n37570 ; n37571
g37316 and n37237_not n37571_not ; n37572
g37317 and n37569_not n37572 ; n37573
g37318 and n37237_not n37573_not ; n37574
g37319 and b[26] n37226_not ; n37575
g37320 and n37220_not n37575 ; n37576
g37321 and n37228_not n37576_not ; n37577
g37322 and n37574_not n37577 ; n37578
g37323 and n37228_not n37578_not ; n37579
g37324 and b[27] n37217_not ; n37580
g37325 and n37211_not n37580 ; n37581
g37326 and n37219_not n37581_not ; n37582
g37327 and n37579_not n37582 ; n37583
g37328 and n37219_not n37583_not ; n37584
g37329 and b[28] n37208_not ; n37585
g37330 and n37202_not n37585 ; n37586
g37331 and n37210_not n37586_not ; n37587
g37332 and n37584_not n37587 ; n37588
g37333 and n37210_not n37588_not ; n37589
g37334 and b[29] n37199_not ; n37590
g37335 and n37193_not n37590 ; n37591
g37336 and n37201_not n37591_not ; n37592
g37337 and n37589_not n37592 ; n37593
g37338 and n37201_not n37593_not ; n37594
g37339 and b[30] n37190_not ; n37595
g37340 and n37184_not n37595 ; n37596
g37341 and n37192_not n37596_not ; n37597
g37342 and n37594_not n37597 ; n37598
g37343 and n37192_not n37598_not ; n37599
g37344 and b[31] n37181_not ; n37600
g37345 and n37175_not n37600 ; n37601
g37346 and n37183_not n37601_not ; n37602
g37347 and n37599_not n37602 ; n37603
g37348 and n37183_not n37603_not ; n37604
g37349 and b[32] n37172_not ; n37605
g37350 and n37166_not n37605 ; n37606
g37351 and n37174_not n37606_not ; n37607
g37352 and n37604_not n37607 ; n37608
g37353 and n37174_not n37608_not ; n37609
g37354 and b[33] n37163_not ; n37610
g37355 and n37157_not n37610 ; n37611
g37356 and n37165_not n37611_not ; n37612
g37357 and n37609_not n37612 ; n37613
g37358 and n37165_not n37613_not ; n37614
g37359 and b[34] n37154_not ; n37615
g37360 and n37148_not n37615 ; n37616
g37361 and n37156_not n37616_not ; n37617
g37362 and n37614_not n37617 ; n37618
g37363 and n37156_not n37618_not ; n37619
g37364 and n36690_not n37147_not ; n37620
g37365 and n36692_not n37144 ; n37621
g37366 and n37140_not n37621 ; n37622
g37367 and n37141_not n37144_not ; n37623
g37368 and n37622_not n37623_not ; n37624
g37369 and n37147 n37624_not ; n37625
g37370 and n37620_not n37625_not ; n37626
g37371 and b[35]_not n37626_not ; n37627
g37372 and b[35] n37620_not ; n37628
g37373 and n37625_not n37628 ; n37629
g37374 and n512 n37629_not ; n37630
g37375 and n37627_not n37630 ; n37631
g37376 and n37619_not n37631 ; n37632
g37377 and n9004 n37626_not ; n37633
g37378 and n37632_not n37633_not ; n37634
g37379 and n37165_not n37617 ; n37635
g37380 and n37613_not n37635 ; n37636
g37381 and n37614_not n37617_not ; n37637
g37382 and n37636_not n37637_not ; n37638
g37383 and n37634_not n37638_not ; n37639
g37384 and n37155_not n37633_not ; n37640
g37385 and n37632_not n37640 ; n37641
g37386 and n37639_not n37641_not ; n37642
g37387 and n37156_not n37629_not ; n37643
g37388 and n37627_not n37643 ; n37644
g37389 and n37618_not n37644 ; n37645
g37390 and n37627_not n37629_not ; n37646
g37391 and n37619_not n37646_not ; n37647
g37392 and n37645_not n37647_not ; n37648
g37393 and n37634_not n37648_not ; n37649
g37394 and n37626_not n37633_not ; n37650
g37395 and n37632_not n37650 ; n37651
g37396 and n37649_not n37651_not ; n37652
g37397 and b[36]_not n37652_not ; n37653
g37398 and b[35]_not n37642_not ; n37654
g37399 and n37174_not n37612 ; n37655
g37400 and n37608_not n37655 ; n37656
g37401 and n37609_not n37612_not ; n37657
g37402 and n37656_not n37657_not ; n37658
g37403 and n37634_not n37658_not ; n37659
g37404 and n37164_not n37633_not ; n37660
g37405 and n37632_not n37660 ; n37661
g37406 and n37659_not n37661_not ; n37662
g37407 and b[34]_not n37662_not ; n37663
g37408 and n37183_not n37607 ; n37664
g37409 and n37603_not n37664 ; n37665
g37410 and n37604_not n37607_not ; n37666
g37411 and n37665_not n37666_not ; n37667
g37412 and n37634_not n37667_not ; n37668
g37413 and n37173_not n37633_not ; n37669
g37414 and n37632_not n37669 ; n37670
g37415 and n37668_not n37670_not ; n37671
g37416 and b[33]_not n37671_not ; n37672
g37417 and n37192_not n37602 ; n37673
g37418 and n37598_not n37673 ; n37674
g37419 and n37599_not n37602_not ; n37675
g37420 and n37674_not n37675_not ; n37676
g37421 and n37634_not n37676_not ; n37677
g37422 and n37182_not n37633_not ; n37678
g37423 and n37632_not n37678 ; n37679
g37424 and n37677_not n37679_not ; n37680
g37425 and b[32]_not n37680_not ; n37681
g37426 and n37201_not n37597 ; n37682
g37427 and n37593_not n37682 ; n37683
g37428 and n37594_not n37597_not ; n37684
g37429 and n37683_not n37684_not ; n37685
g37430 and n37634_not n37685_not ; n37686
g37431 and n37191_not n37633_not ; n37687
g37432 and n37632_not n37687 ; n37688
g37433 and n37686_not n37688_not ; n37689
g37434 and b[31]_not n37689_not ; n37690
g37435 and n37210_not n37592 ; n37691
g37436 and n37588_not n37691 ; n37692
g37437 and n37589_not n37592_not ; n37693
g37438 and n37692_not n37693_not ; n37694
g37439 and n37634_not n37694_not ; n37695
g37440 and n37200_not n37633_not ; n37696
g37441 and n37632_not n37696 ; n37697
g37442 and n37695_not n37697_not ; n37698
g37443 and b[30]_not n37698_not ; n37699
g37444 and n37219_not n37587 ; n37700
g37445 and n37583_not n37700 ; n37701
g37446 and n37584_not n37587_not ; n37702
g37447 and n37701_not n37702_not ; n37703
g37448 and n37634_not n37703_not ; n37704
g37449 and n37209_not n37633_not ; n37705
g37450 and n37632_not n37705 ; n37706
g37451 and n37704_not n37706_not ; n37707
g37452 and b[29]_not n37707_not ; n37708
g37453 and n37228_not n37582 ; n37709
g37454 and n37578_not n37709 ; n37710
g37455 and n37579_not n37582_not ; n37711
g37456 and n37710_not n37711_not ; n37712
g37457 and n37634_not n37712_not ; n37713
g37458 and n37218_not n37633_not ; n37714
g37459 and n37632_not n37714 ; n37715
g37460 and n37713_not n37715_not ; n37716
g37461 and b[28]_not n37716_not ; n37717
g37462 and n37237_not n37577 ; n37718
g37463 and n37573_not n37718 ; n37719
g37464 and n37574_not n37577_not ; n37720
g37465 and n37719_not n37720_not ; n37721
g37466 and n37634_not n37721_not ; n37722
g37467 and n37227_not n37633_not ; n37723
g37468 and n37632_not n37723 ; n37724
g37469 and n37722_not n37724_not ; n37725
g37470 and b[27]_not n37725_not ; n37726
g37471 and n37246_not n37572 ; n37727
g37472 and n37568_not n37727 ; n37728
g37473 and n37569_not n37572_not ; n37729
g37474 and n37728_not n37729_not ; n37730
g37475 and n37634_not n37730_not ; n37731
g37476 and n37236_not n37633_not ; n37732
g37477 and n37632_not n37732 ; n37733
g37478 and n37731_not n37733_not ; n37734
g37479 and b[26]_not n37734_not ; n37735
g37480 and n37255_not n37567 ; n37736
g37481 and n37563_not n37736 ; n37737
g37482 and n37564_not n37567_not ; n37738
g37483 and n37737_not n37738_not ; n37739
g37484 and n37634_not n37739_not ; n37740
g37485 and n37245_not n37633_not ; n37741
g37486 and n37632_not n37741 ; n37742
g37487 and n37740_not n37742_not ; n37743
g37488 and b[25]_not n37743_not ; n37744
g37489 and n37264_not n37562 ; n37745
g37490 and n37558_not n37745 ; n37746
g37491 and n37559_not n37562_not ; n37747
g37492 and n37746_not n37747_not ; n37748
g37493 and n37634_not n37748_not ; n37749
g37494 and n37254_not n37633_not ; n37750
g37495 and n37632_not n37750 ; n37751
g37496 and n37749_not n37751_not ; n37752
g37497 and b[24]_not n37752_not ; n37753
g37498 and n37273_not n37557 ; n37754
g37499 and n37553_not n37754 ; n37755
g37500 and n37554_not n37557_not ; n37756
g37501 and n37755_not n37756_not ; n37757
g37502 and n37634_not n37757_not ; n37758
g37503 and n37263_not n37633_not ; n37759
g37504 and n37632_not n37759 ; n37760
g37505 and n37758_not n37760_not ; n37761
g37506 and b[23]_not n37761_not ; n37762
g37507 and n37282_not n37552 ; n37763
g37508 and n37548_not n37763 ; n37764
g37509 and n37549_not n37552_not ; n37765
g37510 and n37764_not n37765_not ; n37766
g37511 and n37634_not n37766_not ; n37767
g37512 and n37272_not n37633_not ; n37768
g37513 and n37632_not n37768 ; n37769
g37514 and n37767_not n37769_not ; n37770
g37515 and b[22]_not n37770_not ; n37771
g37516 and n37291_not n37547 ; n37772
g37517 and n37543_not n37772 ; n37773
g37518 and n37544_not n37547_not ; n37774
g37519 and n37773_not n37774_not ; n37775
g37520 and n37634_not n37775_not ; n37776
g37521 and n37281_not n37633_not ; n37777
g37522 and n37632_not n37777 ; n37778
g37523 and n37776_not n37778_not ; n37779
g37524 and b[21]_not n37779_not ; n37780
g37525 and n37300_not n37542 ; n37781
g37526 and n37538_not n37781 ; n37782
g37527 and n37539_not n37542_not ; n37783
g37528 and n37782_not n37783_not ; n37784
g37529 and n37634_not n37784_not ; n37785
g37530 and n37290_not n37633_not ; n37786
g37531 and n37632_not n37786 ; n37787
g37532 and n37785_not n37787_not ; n37788
g37533 and b[20]_not n37788_not ; n37789
g37534 and n37309_not n37537 ; n37790
g37535 and n37533_not n37790 ; n37791
g37536 and n37534_not n37537_not ; n37792
g37537 and n37791_not n37792_not ; n37793
g37538 and n37634_not n37793_not ; n37794
g37539 and n37299_not n37633_not ; n37795
g37540 and n37632_not n37795 ; n37796
g37541 and n37794_not n37796_not ; n37797
g37542 and b[19]_not n37797_not ; n37798
g37543 and n37318_not n37532 ; n37799
g37544 and n37528_not n37799 ; n37800
g37545 and n37529_not n37532_not ; n37801
g37546 and n37800_not n37801_not ; n37802
g37547 and n37634_not n37802_not ; n37803
g37548 and n37308_not n37633_not ; n37804
g37549 and n37632_not n37804 ; n37805
g37550 and n37803_not n37805_not ; n37806
g37551 and b[18]_not n37806_not ; n37807
g37552 and n37327_not n37527 ; n37808
g37553 and n37523_not n37808 ; n37809
g37554 and n37524_not n37527_not ; n37810
g37555 and n37809_not n37810_not ; n37811
g37556 and n37634_not n37811_not ; n37812
g37557 and n37317_not n37633_not ; n37813
g37558 and n37632_not n37813 ; n37814
g37559 and n37812_not n37814_not ; n37815
g37560 and b[17]_not n37815_not ; n37816
g37561 and n37336_not n37522 ; n37817
g37562 and n37518_not n37817 ; n37818
g37563 and n37519_not n37522_not ; n37819
g37564 and n37818_not n37819_not ; n37820
g37565 and n37634_not n37820_not ; n37821
g37566 and n37326_not n37633_not ; n37822
g37567 and n37632_not n37822 ; n37823
g37568 and n37821_not n37823_not ; n37824
g37569 and b[16]_not n37824_not ; n37825
g37570 and n37345_not n37517 ; n37826
g37571 and n37513_not n37826 ; n37827
g37572 and n37514_not n37517_not ; n37828
g37573 and n37827_not n37828_not ; n37829
g37574 and n37634_not n37829_not ; n37830
g37575 and n37335_not n37633_not ; n37831
g37576 and n37632_not n37831 ; n37832
g37577 and n37830_not n37832_not ; n37833
g37578 and b[15]_not n37833_not ; n37834
g37579 and n37354_not n37512 ; n37835
g37580 and n37508_not n37835 ; n37836
g37581 and n37509_not n37512_not ; n37837
g37582 and n37836_not n37837_not ; n37838
g37583 and n37634_not n37838_not ; n37839
g37584 and n37344_not n37633_not ; n37840
g37585 and n37632_not n37840 ; n37841
g37586 and n37839_not n37841_not ; n37842
g37587 and b[14]_not n37842_not ; n37843
g37588 and n37363_not n37507 ; n37844
g37589 and n37503_not n37844 ; n37845
g37590 and n37504_not n37507_not ; n37846
g37591 and n37845_not n37846_not ; n37847
g37592 and n37634_not n37847_not ; n37848
g37593 and n37353_not n37633_not ; n37849
g37594 and n37632_not n37849 ; n37850
g37595 and n37848_not n37850_not ; n37851
g37596 and b[13]_not n37851_not ; n37852
g37597 and n37372_not n37502 ; n37853
g37598 and n37498_not n37853 ; n37854
g37599 and n37499_not n37502_not ; n37855
g37600 and n37854_not n37855_not ; n37856
g37601 and n37634_not n37856_not ; n37857
g37602 and n37362_not n37633_not ; n37858
g37603 and n37632_not n37858 ; n37859
g37604 and n37857_not n37859_not ; n37860
g37605 and b[12]_not n37860_not ; n37861
g37606 and n37381_not n37497 ; n37862
g37607 and n37493_not n37862 ; n37863
g37608 and n37494_not n37497_not ; n37864
g37609 and n37863_not n37864_not ; n37865
g37610 and n37634_not n37865_not ; n37866
g37611 and n37371_not n37633_not ; n37867
g37612 and n37632_not n37867 ; n37868
g37613 and n37866_not n37868_not ; n37869
g37614 and b[11]_not n37869_not ; n37870
g37615 and n37390_not n37492 ; n37871
g37616 and n37488_not n37871 ; n37872
g37617 and n37489_not n37492_not ; n37873
g37618 and n37872_not n37873_not ; n37874
g37619 and n37634_not n37874_not ; n37875
g37620 and n37380_not n37633_not ; n37876
g37621 and n37632_not n37876 ; n37877
g37622 and n37875_not n37877_not ; n37878
g37623 and b[10]_not n37878_not ; n37879
g37624 and n37399_not n37487 ; n37880
g37625 and n37483_not n37880 ; n37881
g37626 and n37484_not n37487_not ; n37882
g37627 and n37881_not n37882_not ; n37883
g37628 and n37634_not n37883_not ; n37884
g37629 and n37389_not n37633_not ; n37885
g37630 and n37632_not n37885 ; n37886
g37631 and n37884_not n37886_not ; n37887
g37632 and b[9]_not n37887_not ; n37888
g37633 and n37408_not n37482 ; n37889
g37634 and n37478_not n37889 ; n37890
g37635 and n37479_not n37482_not ; n37891
g37636 and n37890_not n37891_not ; n37892
g37637 and n37634_not n37892_not ; n37893
g37638 and n37398_not n37633_not ; n37894
g37639 and n37632_not n37894 ; n37895
g37640 and n37893_not n37895_not ; n37896
g37641 and b[8]_not n37896_not ; n37897
g37642 and n37417_not n37477 ; n37898
g37643 and n37473_not n37898 ; n37899
g37644 and n37474_not n37477_not ; n37900
g37645 and n37899_not n37900_not ; n37901
g37646 and n37634_not n37901_not ; n37902
g37647 and n37407_not n37633_not ; n37903
g37648 and n37632_not n37903 ; n37904
g37649 and n37902_not n37904_not ; n37905
g37650 and b[7]_not n37905_not ; n37906
g37651 and n37426_not n37472 ; n37907
g37652 and n37468_not n37907 ; n37908
g37653 and n37469_not n37472_not ; n37909
g37654 and n37908_not n37909_not ; n37910
g37655 and n37634_not n37910_not ; n37911
g37656 and n37416_not n37633_not ; n37912
g37657 and n37632_not n37912 ; n37913
g37658 and n37911_not n37913_not ; n37914
g37659 and b[6]_not n37914_not ; n37915
g37660 and n37435_not n37467 ; n37916
g37661 and n37463_not n37916 ; n37917
g37662 and n37464_not n37467_not ; n37918
g37663 and n37917_not n37918_not ; n37919
g37664 and n37634_not n37919_not ; n37920
g37665 and n37425_not n37633_not ; n37921
g37666 and n37632_not n37921 ; n37922
g37667 and n37920_not n37922_not ; n37923
g37668 and b[5]_not n37923_not ; n37924
g37669 and n37443_not n37462 ; n37925
g37670 and n37458_not n37925 ; n37926
g37671 and n37459_not n37462_not ; n37927
g37672 and n37926_not n37927_not ; n37928
g37673 and n37634_not n37928_not ; n37929
g37674 and n37434_not n37633_not ; n37930
g37675 and n37632_not n37930 ; n37931
g37676 and n37929_not n37931_not ; n37932
g37677 and b[4]_not n37932_not ; n37933
g37678 and n37453_not n37457 ; n37934
g37679 and n37452_not n37934 ; n37935
g37680 and n37454_not n37457_not ; n37936
g37681 and n37935_not n37936_not ; n37937
g37682 and n37634_not n37937_not ; n37938
g37683 and n37442_not n37633_not ; n37939
g37684 and n37632_not n37939 ; n37940
g37685 and n37938_not n37940_not ; n37941
g37686 and b[3]_not n37941_not ; n37942
g37687 and n9318 n37450_not ; n37943
g37688 and n37448_not n37943 ; n37944
g37689 and n37452_not n37944_not ; n37945
g37690 and n37634_not n37945 ; n37946
g37691 and n37447_not n37633_not ; n37947
g37692 and n37632_not n37947 ; n37948
g37693 and n37946_not n37948_not ; n37949
g37694 and b[2]_not n37949_not ; n37950
g37695 and b[0] n37634_not ; n37951
g37696 and a[28] n37951_not ; n37952
g37697 and n9318 n37634_not ; n37953
g37698 and n37952_not n37953_not ; n37954
g37699 and b[1] n37954_not ; n37955
g37700 and b[1]_not n37953_not ; n37956
g37701 and n37952_not n37956 ; n37957
g37702 and n37955_not n37957_not ; n37958
g37703 and n9826_not n37958_not ; n37959
g37704 and b[1]_not n37954_not ; n37960
g37705 and n37959_not n37960_not ; n37961
g37706 and b[2] n37948_not ; n37962
g37707 and n37946_not n37962 ; n37963
g37708 and n37950_not n37963_not ; n37964
g37709 and n37961_not n37964 ; n37965
g37710 and n37950_not n37965_not ; n37966
g37711 and b[3] n37940_not ; n37967
g37712 and n37938_not n37967 ; n37968
g37713 and n37942_not n37968_not ; n37969
g37714 and n37966_not n37969 ; n37970
g37715 and n37942_not n37970_not ; n37971
g37716 and b[4] n37931_not ; n37972
g37717 and n37929_not n37972 ; n37973
g37718 and n37933_not n37973_not ; n37974
g37719 and n37971_not n37974 ; n37975
g37720 and n37933_not n37975_not ; n37976
g37721 and b[5] n37922_not ; n37977
g37722 and n37920_not n37977 ; n37978
g37723 and n37924_not n37978_not ; n37979
g37724 and n37976_not n37979 ; n37980
g37725 and n37924_not n37980_not ; n37981
g37726 and b[6] n37913_not ; n37982
g37727 and n37911_not n37982 ; n37983
g37728 and n37915_not n37983_not ; n37984
g37729 and n37981_not n37984 ; n37985
g37730 and n37915_not n37985_not ; n37986
g37731 and b[7] n37904_not ; n37987
g37732 and n37902_not n37987 ; n37988
g37733 and n37906_not n37988_not ; n37989
g37734 and n37986_not n37989 ; n37990
g37735 and n37906_not n37990_not ; n37991
g37736 and b[8] n37895_not ; n37992
g37737 and n37893_not n37992 ; n37993
g37738 and n37897_not n37993_not ; n37994
g37739 and n37991_not n37994 ; n37995
g37740 and n37897_not n37995_not ; n37996
g37741 and b[9] n37886_not ; n37997
g37742 and n37884_not n37997 ; n37998
g37743 and n37888_not n37998_not ; n37999
g37744 and n37996_not n37999 ; n38000
g37745 and n37888_not n38000_not ; n38001
g37746 and b[10] n37877_not ; n38002
g37747 and n37875_not n38002 ; n38003
g37748 and n37879_not n38003_not ; n38004
g37749 and n38001_not n38004 ; n38005
g37750 and n37879_not n38005_not ; n38006
g37751 and b[11] n37868_not ; n38007
g37752 and n37866_not n38007 ; n38008
g37753 and n37870_not n38008_not ; n38009
g37754 and n38006_not n38009 ; n38010
g37755 and n37870_not n38010_not ; n38011
g37756 and b[12] n37859_not ; n38012
g37757 and n37857_not n38012 ; n38013
g37758 and n37861_not n38013_not ; n38014
g37759 and n38011_not n38014 ; n38015
g37760 and n37861_not n38015_not ; n38016
g37761 and b[13] n37850_not ; n38017
g37762 and n37848_not n38017 ; n38018
g37763 and n37852_not n38018_not ; n38019
g37764 and n38016_not n38019 ; n38020
g37765 and n37852_not n38020_not ; n38021
g37766 and b[14] n37841_not ; n38022
g37767 and n37839_not n38022 ; n38023
g37768 and n37843_not n38023_not ; n38024
g37769 and n38021_not n38024 ; n38025
g37770 and n37843_not n38025_not ; n38026
g37771 and b[15] n37832_not ; n38027
g37772 and n37830_not n38027 ; n38028
g37773 and n37834_not n38028_not ; n38029
g37774 and n38026_not n38029 ; n38030
g37775 and n37834_not n38030_not ; n38031
g37776 and b[16] n37823_not ; n38032
g37777 and n37821_not n38032 ; n38033
g37778 and n37825_not n38033_not ; n38034
g37779 and n38031_not n38034 ; n38035
g37780 and n37825_not n38035_not ; n38036
g37781 and b[17] n37814_not ; n38037
g37782 and n37812_not n38037 ; n38038
g37783 and n37816_not n38038_not ; n38039
g37784 and n38036_not n38039 ; n38040
g37785 and n37816_not n38040_not ; n38041
g37786 and b[18] n37805_not ; n38042
g37787 and n37803_not n38042 ; n38043
g37788 and n37807_not n38043_not ; n38044
g37789 and n38041_not n38044 ; n38045
g37790 and n37807_not n38045_not ; n38046
g37791 and b[19] n37796_not ; n38047
g37792 and n37794_not n38047 ; n38048
g37793 and n37798_not n38048_not ; n38049
g37794 and n38046_not n38049 ; n38050
g37795 and n37798_not n38050_not ; n38051
g37796 and b[20] n37787_not ; n38052
g37797 and n37785_not n38052 ; n38053
g37798 and n37789_not n38053_not ; n38054
g37799 and n38051_not n38054 ; n38055
g37800 and n37789_not n38055_not ; n38056
g37801 and b[21] n37778_not ; n38057
g37802 and n37776_not n38057 ; n38058
g37803 and n37780_not n38058_not ; n38059
g37804 and n38056_not n38059 ; n38060
g37805 and n37780_not n38060_not ; n38061
g37806 and b[22] n37769_not ; n38062
g37807 and n37767_not n38062 ; n38063
g37808 and n37771_not n38063_not ; n38064
g37809 and n38061_not n38064 ; n38065
g37810 and n37771_not n38065_not ; n38066
g37811 and b[23] n37760_not ; n38067
g37812 and n37758_not n38067 ; n38068
g37813 and n37762_not n38068_not ; n38069
g37814 and n38066_not n38069 ; n38070
g37815 and n37762_not n38070_not ; n38071
g37816 and b[24] n37751_not ; n38072
g37817 and n37749_not n38072 ; n38073
g37818 and n37753_not n38073_not ; n38074
g37819 and n38071_not n38074 ; n38075
g37820 and n37753_not n38075_not ; n38076
g37821 and b[25] n37742_not ; n38077
g37822 and n37740_not n38077 ; n38078
g37823 and n37744_not n38078_not ; n38079
g37824 and n38076_not n38079 ; n38080
g37825 and n37744_not n38080_not ; n38081
g37826 and b[26] n37733_not ; n38082
g37827 and n37731_not n38082 ; n38083
g37828 and n37735_not n38083_not ; n38084
g37829 and n38081_not n38084 ; n38085
g37830 and n37735_not n38085_not ; n38086
g37831 and b[27] n37724_not ; n38087
g37832 and n37722_not n38087 ; n38088
g37833 and n37726_not n38088_not ; n38089
g37834 and n38086_not n38089 ; n38090
g37835 and n37726_not n38090_not ; n38091
g37836 and b[28] n37715_not ; n38092
g37837 and n37713_not n38092 ; n38093
g37838 and n37717_not n38093_not ; n38094
g37839 and n38091_not n38094 ; n38095
g37840 and n37717_not n38095_not ; n38096
g37841 and b[29] n37706_not ; n38097
g37842 and n37704_not n38097 ; n38098
g37843 and n37708_not n38098_not ; n38099
g37844 and n38096_not n38099 ; n38100
g37845 and n37708_not n38100_not ; n38101
g37846 and b[30] n37697_not ; n38102
g37847 and n37695_not n38102 ; n38103
g37848 and n37699_not n38103_not ; n38104
g37849 and n38101_not n38104 ; n38105
g37850 and n37699_not n38105_not ; n38106
g37851 and b[31] n37688_not ; n38107
g37852 and n37686_not n38107 ; n38108
g37853 and n37690_not n38108_not ; n38109
g37854 and n38106_not n38109 ; n38110
g37855 and n37690_not n38110_not ; n38111
g37856 and b[32] n37679_not ; n38112
g37857 and n37677_not n38112 ; n38113
g37858 and n37681_not n38113_not ; n38114
g37859 and n38111_not n38114 ; n38115
g37860 and n37681_not n38115_not ; n38116
g37861 and b[33] n37670_not ; n38117
g37862 and n37668_not n38117 ; n38118
g37863 and n37672_not n38118_not ; n38119
g37864 and n38116_not n38119 ; n38120
g37865 and n37672_not n38120_not ; n38121
g37866 and b[34] n37661_not ; n38122
g37867 and n37659_not n38122 ; n38123
g37868 and n37663_not n38123_not ; n38124
g37869 and n38121_not n38124 ; n38125
g37870 and n37663_not n38125_not ; n38126
g37871 and b[35] n37641_not ; n38127
g37872 and n37639_not n38127 ; n38128
g37873 and n37654_not n38128_not ; n38129
g37874 and n38126_not n38129 ; n38130
g37875 and n37654_not n38130_not ; n38131
g37876 and b[36] n37651_not ; n38132
g37877 and n37649_not n38132 ; n38133
g37878 and n37653_not n38133_not ; n38134
g37879 and n38131_not n38134 ; n38135
g37880 and n37653_not n38135_not ; n38136
g37881 and n599 n38136_not ; n38137
g37882 and n37642_not n38137_not ; n38138
g37883 and n37663_not n38129 ; n38139
g37884 and n38125_not n38139 ; n38140
g37885 and n38126_not n38129_not ; n38141
g37886 and n38140_not n38141_not ; n38142
g37887 and n599 n38142_not ; n38143
g37888 and n38136_not n38143 ; n38144
g37889 and n38138_not n38144_not ; n38145
g37890 and n37652_not n38137_not ; n38146
g37891 and n37654_not n38134 ; n38147
g37892 and n38130_not n38147 ; n38148
g37893 and n38131_not n38134_not ; n38149
g37894 and n38148_not n38149_not ; n38150
g37895 and n38137 n38150_not ; n38151
g37896 and n38146_not n38151_not ; n38152
g37897 and b[37]_not n38152_not ; n38153
g37898 and b[36]_not n38145_not ; n38154
g37899 and n37662_not n38137_not ; n38155
g37900 and n37672_not n38124 ; n38156
g37901 and n38120_not n38156 ; n38157
g37902 and n38121_not n38124_not ; n38158
g37903 and n38157_not n38158_not ; n38159
g37904 and n599 n38159_not ; n38160
g37905 and n38136_not n38160 ; n38161
g37906 and n38155_not n38161_not ; n38162
g37907 and b[35]_not n38162_not ; n38163
g37908 and n37671_not n38137_not ; n38164
g37909 and n37681_not n38119 ; n38165
g37910 and n38115_not n38165 ; n38166
g37911 and n38116_not n38119_not ; n38167
g37912 and n38166_not n38167_not ; n38168
g37913 and n599 n38168_not ; n38169
g37914 and n38136_not n38169 ; n38170
g37915 and n38164_not n38170_not ; n38171
g37916 and b[34]_not n38171_not ; n38172
g37917 and n37680_not n38137_not ; n38173
g37918 and n37690_not n38114 ; n38174
g37919 and n38110_not n38174 ; n38175
g37920 and n38111_not n38114_not ; n38176
g37921 and n38175_not n38176_not ; n38177
g37922 and n599 n38177_not ; n38178
g37923 and n38136_not n38178 ; n38179
g37924 and n38173_not n38179_not ; n38180
g37925 and b[33]_not n38180_not ; n38181
g37926 and n37689_not n38137_not ; n38182
g37927 and n37699_not n38109 ; n38183
g37928 and n38105_not n38183 ; n38184
g37929 and n38106_not n38109_not ; n38185
g37930 and n38184_not n38185_not ; n38186
g37931 and n599 n38186_not ; n38187
g37932 and n38136_not n38187 ; n38188
g37933 and n38182_not n38188_not ; n38189
g37934 and b[32]_not n38189_not ; n38190
g37935 and n37698_not n38137_not ; n38191
g37936 and n37708_not n38104 ; n38192
g37937 and n38100_not n38192 ; n38193
g37938 and n38101_not n38104_not ; n38194
g37939 and n38193_not n38194_not ; n38195
g37940 and n599 n38195_not ; n38196
g37941 and n38136_not n38196 ; n38197
g37942 and n38191_not n38197_not ; n38198
g37943 and b[31]_not n38198_not ; n38199
g37944 and n37707_not n38137_not ; n38200
g37945 and n37717_not n38099 ; n38201
g37946 and n38095_not n38201 ; n38202
g37947 and n38096_not n38099_not ; n38203
g37948 and n38202_not n38203_not ; n38204
g37949 and n599 n38204_not ; n38205
g37950 and n38136_not n38205 ; n38206
g37951 and n38200_not n38206_not ; n38207
g37952 and b[30]_not n38207_not ; n38208
g37953 and n37716_not n38137_not ; n38209
g37954 and n37726_not n38094 ; n38210
g37955 and n38090_not n38210 ; n38211
g37956 and n38091_not n38094_not ; n38212
g37957 and n38211_not n38212_not ; n38213
g37958 and n599 n38213_not ; n38214
g37959 and n38136_not n38214 ; n38215
g37960 and n38209_not n38215_not ; n38216
g37961 and b[29]_not n38216_not ; n38217
g37962 and n37725_not n38137_not ; n38218
g37963 and n37735_not n38089 ; n38219
g37964 and n38085_not n38219 ; n38220
g37965 and n38086_not n38089_not ; n38221
g37966 and n38220_not n38221_not ; n38222
g37967 and n599 n38222_not ; n38223
g37968 and n38136_not n38223 ; n38224
g37969 and n38218_not n38224_not ; n38225
g37970 and b[28]_not n38225_not ; n38226
g37971 and n37734_not n38137_not ; n38227
g37972 and n37744_not n38084 ; n38228
g37973 and n38080_not n38228 ; n38229
g37974 and n38081_not n38084_not ; n38230
g37975 and n38229_not n38230_not ; n38231
g37976 and n599 n38231_not ; n38232
g37977 and n38136_not n38232 ; n38233
g37978 and n38227_not n38233_not ; n38234
g37979 and b[27]_not n38234_not ; n38235
g37980 and n37743_not n38137_not ; n38236
g37981 and n37753_not n38079 ; n38237
g37982 and n38075_not n38237 ; n38238
g37983 and n38076_not n38079_not ; n38239
g37984 and n38238_not n38239_not ; n38240
g37985 and n599 n38240_not ; n38241
g37986 and n38136_not n38241 ; n38242
g37987 and n38236_not n38242_not ; n38243
g37988 and b[26]_not n38243_not ; n38244
g37989 and n37752_not n38137_not ; n38245
g37990 and n37762_not n38074 ; n38246
g37991 and n38070_not n38246 ; n38247
g37992 and n38071_not n38074_not ; n38248
g37993 and n38247_not n38248_not ; n38249
g37994 and n599 n38249_not ; n38250
g37995 and n38136_not n38250 ; n38251
g37996 and n38245_not n38251_not ; n38252
g37997 and b[25]_not n38252_not ; n38253
g37998 and n37761_not n38137_not ; n38254
g37999 and n37771_not n38069 ; n38255
g38000 and n38065_not n38255 ; n38256
g38001 and n38066_not n38069_not ; n38257
g38002 and n38256_not n38257_not ; n38258
g38003 and n599 n38258_not ; n38259
g38004 and n38136_not n38259 ; n38260
g38005 and n38254_not n38260_not ; n38261
g38006 and b[24]_not n38261_not ; n38262
g38007 and n37770_not n38137_not ; n38263
g38008 and n37780_not n38064 ; n38264
g38009 and n38060_not n38264 ; n38265
g38010 and n38061_not n38064_not ; n38266
g38011 and n38265_not n38266_not ; n38267
g38012 and n599 n38267_not ; n38268
g38013 and n38136_not n38268 ; n38269
g38014 and n38263_not n38269_not ; n38270
g38015 and b[23]_not n38270_not ; n38271
g38016 and n37779_not n38137_not ; n38272
g38017 and n37789_not n38059 ; n38273
g38018 and n38055_not n38273 ; n38274
g38019 and n38056_not n38059_not ; n38275
g38020 and n38274_not n38275_not ; n38276
g38021 and n599 n38276_not ; n38277
g38022 and n38136_not n38277 ; n38278
g38023 and n38272_not n38278_not ; n38279
g38024 and b[22]_not n38279_not ; n38280
g38025 and n37788_not n38137_not ; n38281
g38026 and n37798_not n38054 ; n38282
g38027 and n38050_not n38282 ; n38283
g38028 and n38051_not n38054_not ; n38284
g38029 and n38283_not n38284_not ; n38285
g38030 and n599 n38285_not ; n38286
g38031 and n38136_not n38286 ; n38287
g38032 and n38281_not n38287_not ; n38288
g38033 and b[21]_not n38288_not ; n38289
g38034 and n37797_not n38137_not ; n38290
g38035 and n37807_not n38049 ; n38291
g38036 and n38045_not n38291 ; n38292
g38037 and n38046_not n38049_not ; n38293
g38038 and n38292_not n38293_not ; n38294
g38039 and n599 n38294_not ; n38295
g38040 and n38136_not n38295 ; n38296
g38041 and n38290_not n38296_not ; n38297
g38042 and b[20]_not n38297_not ; n38298
g38043 and n37806_not n38137_not ; n38299
g38044 and n37816_not n38044 ; n38300
g38045 and n38040_not n38300 ; n38301
g38046 and n38041_not n38044_not ; n38302
g38047 and n38301_not n38302_not ; n38303
g38048 and n599 n38303_not ; n38304
g38049 and n38136_not n38304 ; n38305
g38050 and n38299_not n38305_not ; n38306
g38051 and b[19]_not n38306_not ; n38307
g38052 and n37815_not n38137_not ; n38308
g38053 and n37825_not n38039 ; n38309
g38054 and n38035_not n38309 ; n38310
g38055 and n38036_not n38039_not ; n38311
g38056 and n38310_not n38311_not ; n38312
g38057 and n599 n38312_not ; n38313
g38058 and n38136_not n38313 ; n38314
g38059 and n38308_not n38314_not ; n38315
g38060 and b[18]_not n38315_not ; n38316
g38061 and n37824_not n38137_not ; n38317
g38062 and n37834_not n38034 ; n38318
g38063 and n38030_not n38318 ; n38319
g38064 and n38031_not n38034_not ; n38320
g38065 and n38319_not n38320_not ; n38321
g38066 and n599 n38321_not ; n38322
g38067 and n38136_not n38322 ; n38323
g38068 and n38317_not n38323_not ; n38324
g38069 and b[17]_not n38324_not ; n38325
g38070 and n37833_not n38137_not ; n38326
g38071 and n37843_not n38029 ; n38327
g38072 and n38025_not n38327 ; n38328
g38073 and n38026_not n38029_not ; n38329
g38074 and n38328_not n38329_not ; n38330
g38075 and n599 n38330_not ; n38331
g38076 and n38136_not n38331 ; n38332
g38077 and n38326_not n38332_not ; n38333
g38078 and b[16]_not n38333_not ; n38334
g38079 and n37842_not n38137_not ; n38335
g38080 and n37852_not n38024 ; n38336
g38081 and n38020_not n38336 ; n38337
g38082 and n38021_not n38024_not ; n38338
g38083 and n38337_not n38338_not ; n38339
g38084 and n599 n38339_not ; n38340
g38085 and n38136_not n38340 ; n38341
g38086 and n38335_not n38341_not ; n38342
g38087 and b[15]_not n38342_not ; n38343
g38088 and n37851_not n38137_not ; n38344
g38089 and n37861_not n38019 ; n38345
g38090 and n38015_not n38345 ; n38346
g38091 and n38016_not n38019_not ; n38347
g38092 and n38346_not n38347_not ; n38348
g38093 and n599 n38348_not ; n38349
g38094 and n38136_not n38349 ; n38350
g38095 and n38344_not n38350_not ; n38351
g38096 and b[14]_not n38351_not ; n38352
g38097 and n37860_not n38137_not ; n38353
g38098 and n37870_not n38014 ; n38354
g38099 and n38010_not n38354 ; n38355
g38100 and n38011_not n38014_not ; n38356
g38101 and n38355_not n38356_not ; n38357
g38102 and n599 n38357_not ; n38358
g38103 and n38136_not n38358 ; n38359
g38104 and n38353_not n38359_not ; n38360
g38105 and b[13]_not n38360_not ; n38361
g38106 and n37869_not n38137_not ; n38362
g38107 and n37879_not n38009 ; n38363
g38108 and n38005_not n38363 ; n38364
g38109 and n38006_not n38009_not ; n38365
g38110 and n38364_not n38365_not ; n38366
g38111 and n599 n38366_not ; n38367
g38112 and n38136_not n38367 ; n38368
g38113 and n38362_not n38368_not ; n38369
g38114 and b[12]_not n38369_not ; n38370
g38115 and n37878_not n38137_not ; n38371
g38116 and n37888_not n38004 ; n38372
g38117 and n38000_not n38372 ; n38373
g38118 and n38001_not n38004_not ; n38374
g38119 and n38373_not n38374_not ; n38375
g38120 and n599 n38375_not ; n38376
g38121 and n38136_not n38376 ; n38377
g38122 and n38371_not n38377_not ; n38378
g38123 and b[11]_not n38378_not ; n38379
g38124 and n37887_not n38137_not ; n38380
g38125 and n37897_not n37999 ; n38381
g38126 and n37995_not n38381 ; n38382
g38127 and n37996_not n37999_not ; n38383
g38128 and n38382_not n38383_not ; n38384
g38129 and n599 n38384_not ; n38385
g38130 and n38136_not n38385 ; n38386
g38131 and n38380_not n38386_not ; n38387
g38132 and b[10]_not n38387_not ; n38388
g38133 and n37896_not n38137_not ; n38389
g38134 and n37906_not n37994 ; n38390
g38135 and n37990_not n38390 ; n38391
g38136 and n37991_not n37994_not ; n38392
g38137 and n38391_not n38392_not ; n38393
g38138 and n599 n38393_not ; n38394
g38139 and n38136_not n38394 ; n38395
g38140 and n38389_not n38395_not ; n38396
g38141 and b[9]_not n38396_not ; n38397
g38142 and n37905_not n38137_not ; n38398
g38143 and n37915_not n37989 ; n38399
g38144 and n37985_not n38399 ; n38400
g38145 and n37986_not n37989_not ; n38401
g38146 and n38400_not n38401_not ; n38402
g38147 and n599 n38402_not ; n38403
g38148 and n38136_not n38403 ; n38404
g38149 and n38398_not n38404_not ; n38405
g38150 and b[8]_not n38405_not ; n38406
g38151 and n37914_not n38137_not ; n38407
g38152 and n37924_not n37984 ; n38408
g38153 and n37980_not n38408 ; n38409
g38154 and n37981_not n37984_not ; n38410
g38155 and n38409_not n38410_not ; n38411
g38156 and n599 n38411_not ; n38412
g38157 and n38136_not n38412 ; n38413
g38158 and n38407_not n38413_not ; n38414
g38159 and b[7]_not n38414_not ; n38415
g38160 and n37923_not n38137_not ; n38416
g38161 and n37933_not n37979 ; n38417
g38162 and n37975_not n38417 ; n38418
g38163 and n37976_not n37979_not ; n38419
g38164 and n38418_not n38419_not ; n38420
g38165 and n599 n38420_not ; n38421
g38166 and n38136_not n38421 ; n38422
g38167 and n38416_not n38422_not ; n38423
g38168 and b[6]_not n38423_not ; n38424
g38169 and n37932_not n38137_not ; n38425
g38170 and n37942_not n37974 ; n38426
g38171 and n37970_not n38426 ; n38427
g38172 and n37971_not n37974_not ; n38428
g38173 and n38427_not n38428_not ; n38429
g38174 and n599 n38429_not ; n38430
g38175 and n38136_not n38430 ; n38431
g38176 and n38425_not n38431_not ; n38432
g38177 and b[5]_not n38432_not ; n38433
g38178 and n37941_not n38137_not ; n38434
g38179 and n37950_not n37969 ; n38435
g38180 and n37965_not n38435 ; n38436
g38181 and n37966_not n37969_not ; n38437
g38182 and n38436_not n38437_not ; n38438
g38183 and n599 n38438_not ; n38439
g38184 and n38136_not n38439 ; n38440
g38185 and n38434_not n38440_not ; n38441
g38186 and b[4]_not n38441_not ; n38442
g38187 and n37949_not n38137_not ; n38443
g38188 and n37960_not n37964 ; n38444
g38189 and n37959_not n38444 ; n38445
g38190 and n37961_not n37964_not ; n38446
g38191 and n38445_not n38446_not ; n38447
g38192 and n599 n38447_not ; n38448
g38193 and n38136_not n38448 ; n38449
g38194 and n38443_not n38449_not ; n38450
g38195 and b[3]_not n38450_not ; n38451
g38196 and n37954_not n38137_not ; n38452
g38197 and n9826 n37957_not ; n38453
g38198 and n37955_not n38453 ; n38454
g38199 and n599 n38454_not ; n38455
g38200 and n37959_not n38455 ; n38456
g38201 and n38136_not n38456 ; n38457
g38202 and n38452_not n38457_not ; n38458
g38203 and b[2]_not n38458_not ; n38459
g38204 and n10332 n38136_not ; n38460
g38205 and a[27] n38460_not ; n38461
g38206 and n10337 n38136_not ; n38462
g38207 and n38461_not n38462_not ; n38463
g38208 and b[1] n38463_not ; n38464
g38209 and b[1]_not n38462_not ; n38465
g38210 and n38461_not n38465 ; n38466
g38211 and n38464_not n38466_not ; n38467
g38212 and n10344_not n38467_not ; n38468
g38213 and b[1]_not n38463_not ; n38469
g38214 and n38468_not n38469_not ; n38470
g38215 and b[2] n38457_not ; n38471
g38216 and n38452_not n38471 ; n38472
g38217 and n38459_not n38472_not ; n38473
g38218 and n38470_not n38473 ; n38474
g38219 and n38459_not n38474_not ; n38475
g38220 and b[3] n38449_not ; n38476
g38221 and n38443_not n38476 ; n38477
g38222 and n38451_not n38477_not ; n38478
g38223 and n38475_not n38478 ; n38479
g38224 and n38451_not n38479_not ; n38480
g38225 and b[4] n38440_not ; n38481
g38226 and n38434_not n38481 ; n38482
g38227 and n38442_not n38482_not ; n38483
g38228 and n38480_not n38483 ; n38484
g38229 and n38442_not n38484_not ; n38485
g38230 and b[5] n38431_not ; n38486
g38231 and n38425_not n38486 ; n38487
g38232 and n38433_not n38487_not ; n38488
g38233 and n38485_not n38488 ; n38489
g38234 and n38433_not n38489_not ; n38490
g38235 and b[6] n38422_not ; n38491
g38236 and n38416_not n38491 ; n38492
g38237 and n38424_not n38492_not ; n38493
g38238 and n38490_not n38493 ; n38494
g38239 and n38424_not n38494_not ; n38495
g38240 and b[7] n38413_not ; n38496
g38241 and n38407_not n38496 ; n38497
g38242 and n38415_not n38497_not ; n38498
g38243 and n38495_not n38498 ; n38499
g38244 and n38415_not n38499_not ; n38500
g38245 and b[8] n38404_not ; n38501
g38246 and n38398_not n38501 ; n38502
g38247 and n38406_not n38502_not ; n38503
g38248 and n38500_not n38503 ; n38504
g38249 and n38406_not n38504_not ; n38505
g38250 and b[9] n38395_not ; n38506
g38251 and n38389_not n38506 ; n38507
g38252 and n38397_not n38507_not ; n38508
g38253 and n38505_not n38508 ; n38509
g38254 and n38397_not n38509_not ; n38510
g38255 and b[10] n38386_not ; n38511
g38256 and n38380_not n38511 ; n38512
g38257 and n38388_not n38512_not ; n38513
g38258 and n38510_not n38513 ; n38514
g38259 and n38388_not n38514_not ; n38515
g38260 and b[11] n38377_not ; n38516
g38261 and n38371_not n38516 ; n38517
g38262 and n38379_not n38517_not ; n38518
g38263 and n38515_not n38518 ; n38519
g38264 and n38379_not n38519_not ; n38520
g38265 and b[12] n38368_not ; n38521
g38266 and n38362_not n38521 ; n38522
g38267 and n38370_not n38522_not ; n38523
g38268 and n38520_not n38523 ; n38524
g38269 and n38370_not n38524_not ; n38525
g38270 and b[13] n38359_not ; n38526
g38271 and n38353_not n38526 ; n38527
g38272 and n38361_not n38527_not ; n38528
g38273 and n38525_not n38528 ; n38529
g38274 and n38361_not n38529_not ; n38530
g38275 and b[14] n38350_not ; n38531
g38276 and n38344_not n38531 ; n38532
g38277 and n38352_not n38532_not ; n38533
g38278 and n38530_not n38533 ; n38534
g38279 and n38352_not n38534_not ; n38535
g38280 and b[15] n38341_not ; n38536
g38281 and n38335_not n38536 ; n38537
g38282 and n38343_not n38537_not ; n38538
g38283 and n38535_not n38538 ; n38539
g38284 and n38343_not n38539_not ; n38540
g38285 and b[16] n38332_not ; n38541
g38286 and n38326_not n38541 ; n38542
g38287 and n38334_not n38542_not ; n38543
g38288 and n38540_not n38543 ; n38544
g38289 and n38334_not n38544_not ; n38545
g38290 and b[17] n38323_not ; n38546
g38291 and n38317_not n38546 ; n38547
g38292 and n38325_not n38547_not ; n38548
g38293 and n38545_not n38548 ; n38549
g38294 and n38325_not n38549_not ; n38550
g38295 and b[18] n38314_not ; n38551
g38296 and n38308_not n38551 ; n38552
g38297 and n38316_not n38552_not ; n38553
g38298 and n38550_not n38553 ; n38554
g38299 and n38316_not n38554_not ; n38555
g38300 and b[19] n38305_not ; n38556
g38301 and n38299_not n38556 ; n38557
g38302 and n38307_not n38557_not ; n38558
g38303 and n38555_not n38558 ; n38559
g38304 and n38307_not n38559_not ; n38560
g38305 and b[20] n38296_not ; n38561
g38306 and n38290_not n38561 ; n38562
g38307 and n38298_not n38562_not ; n38563
g38308 and n38560_not n38563 ; n38564
g38309 and n38298_not n38564_not ; n38565
g38310 and b[21] n38287_not ; n38566
g38311 and n38281_not n38566 ; n38567
g38312 and n38289_not n38567_not ; n38568
g38313 and n38565_not n38568 ; n38569
g38314 and n38289_not n38569_not ; n38570
g38315 and b[22] n38278_not ; n38571
g38316 and n38272_not n38571 ; n38572
g38317 and n38280_not n38572_not ; n38573
g38318 and n38570_not n38573 ; n38574
g38319 and n38280_not n38574_not ; n38575
g38320 and b[23] n38269_not ; n38576
g38321 and n38263_not n38576 ; n38577
g38322 and n38271_not n38577_not ; n38578
g38323 and n38575_not n38578 ; n38579
g38324 and n38271_not n38579_not ; n38580
g38325 and b[24] n38260_not ; n38581
g38326 and n38254_not n38581 ; n38582
g38327 and n38262_not n38582_not ; n38583
g38328 and n38580_not n38583 ; n38584
g38329 and n38262_not n38584_not ; n38585
g38330 and b[25] n38251_not ; n38586
g38331 and n38245_not n38586 ; n38587
g38332 and n38253_not n38587_not ; n38588
g38333 and n38585_not n38588 ; n38589
g38334 and n38253_not n38589_not ; n38590
g38335 and b[26] n38242_not ; n38591
g38336 and n38236_not n38591 ; n38592
g38337 and n38244_not n38592_not ; n38593
g38338 and n38590_not n38593 ; n38594
g38339 and n38244_not n38594_not ; n38595
g38340 and b[27] n38233_not ; n38596
g38341 and n38227_not n38596 ; n38597
g38342 and n38235_not n38597_not ; n38598
g38343 and n38595_not n38598 ; n38599
g38344 and n38235_not n38599_not ; n38600
g38345 and b[28] n38224_not ; n38601
g38346 and n38218_not n38601 ; n38602
g38347 and n38226_not n38602_not ; n38603
g38348 and n38600_not n38603 ; n38604
g38349 and n38226_not n38604_not ; n38605
g38350 and b[29] n38215_not ; n38606
g38351 and n38209_not n38606 ; n38607
g38352 and n38217_not n38607_not ; n38608
g38353 and n38605_not n38608 ; n38609
g38354 and n38217_not n38609_not ; n38610
g38355 and b[30] n38206_not ; n38611
g38356 and n38200_not n38611 ; n38612
g38357 and n38208_not n38612_not ; n38613
g38358 and n38610_not n38613 ; n38614
g38359 and n38208_not n38614_not ; n38615
g38360 and b[31] n38197_not ; n38616
g38361 and n38191_not n38616 ; n38617
g38362 and n38199_not n38617_not ; n38618
g38363 and n38615_not n38618 ; n38619
g38364 and n38199_not n38619_not ; n38620
g38365 and b[32] n38188_not ; n38621
g38366 and n38182_not n38621 ; n38622
g38367 and n38190_not n38622_not ; n38623
g38368 and n38620_not n38623 ; n38624
g38369 and n38190_not n38624_not ; n38625
g38370 and b[33] n38179_not ; n38626
g38371 and n38173_not n38626 ; n38627
g38372 and n38181_not n38627_not ; n38628
g38373 and n38625_not n38628 ; n38629
g38374 and n38181_not n38629_not ; n38630
g38375 and b[34] n38170_not ; n38631
g38376 and n38164_not n38631 ; n38632
g38377 and n38172_not n38632_not ; n38633
g38378 and n38630_not n38633 ; n38634
g38379 and n38172_not n38634_not ; n38635
g38380 and b[35] n38161_not ; n38636
g38381 and n38155_not n38636 ; n38637
g38382 and n38163_not n38637_not ; n38638
g38383 and n38635_not n38638 ; n38639
g38384 and n38163_not n38639_not ; n38640
g38385 and b[36] n38144_not ; n38641
g38386 and n38138_not n38641 ; n38642
g38387 and n38154_not n38642_not ; n38643
g38388 and n38640_not n38643 ; n38644
g38389 and n38154_not n38644_not ; n38645
g38390 and b[37] n38146_not ; n38646
g38391 and n38151_not n38646 ; n38647
g38392 and n38153_not n38647_not ; n38648
g38393 and n38645_not n38648 ; n38649
g38394 and n38153_not n38649_not ; n38650
g38395 and n10530 n38650_not ; n38651
g38396 and n38145_not n38651_not ; n38652
g38397 and n38163_not n38643 ; n38653
g38398 and n38639_not n38653 ; n38654
g38399 and n38640_not n38643_not ; n38655
g38400 and n38654_not n38655_not ; n38656
g38401 and n10530 n38656_not ; n38657
g38402 and n38650_not n38657 ; n38658
g38403 and n38652_not n38658_not ; n38659
g38404 and b[37]_not n38659_not ; n38660
g38405 and n38162_not n38651_not ; n38661
g38406 and n38172_not n38638 ; n38662
g38407 and n38634_not n38662 ; n38663
g38408 and n38635_not n38638_not ; n38664
g38409 and n38663_not n38664_not ; n38665
g38410 and n10530 n38665_not ; n38666
g38411 and n38650_not n38666 ; n38667
g38412 and n38661_not n38667_not ; n38668
g38413 and b[36]_not n38668_not ; n38669
g38414 and n38171_not n38651_not ; n38670
g38415 and n38181_not n38633 ; n38671
g38416 and n38629_not n38671 ; n38672
g38417 and n38630_not n38633_not ; n38673
g38418 and n38672_not n38673_not ; n38674
g38419 and n10530 n38674_not ; n38675
g38420 and n38650_not n38675 ; n38676
g38421 and n38670_not n38676_not ; n38677
g38422 and b[35]_not n38677_not ; n38678
g38423 and n38180_not n38651_not ; n38679
g38424 and n38190_not n38628 ; n38680
g38425 and n38624_not n38680 ; n38681
g38426 and n38625_not n38628_not ; n38682
g38427 and n38681_not n38682_not ; n38683
g38428 and n10530 n38683_not ; n38684
g38429 and n38650_not n38684 ; n38685
g38430 and n38679_not n38685_not ; n38686
g38431 and b[34]_not n38686_not ; n38687
g38432 and n38189_not n38651_not ; n38688
g38433 and n38199_not n38623 ; n38689
g38434 and n38619_not n38689 ; n38690
g38435 and n38620_not n38623_not ; n38691
g38436 and n38690_not n38691_not ; n38692
g38437 and n10530 n38692_not ; n38693
g38438 and n38650_not n38693 ; n38694
g38439 and n38688_not n38694_not ; n38695
g38440 and b[33]_not n38695_not ; n38696
g38441 and n38198_not n38651_not ; n38697
g38442 and n38208_not n38618 ; n38698
g38443 and n38614_not n38698 ; n38699
g38444 and n38615_not n38618_not ; n38700
g38445 and n38699_not n38700_not ; n38701
g38446 and n10530 n38701_not ; n38702
g38447 and n38650_not n38702 ; n38703
g38448 and n38697_not n38703_not ; n38704
g38449 and b[32]_not n38704_not ; n38705
g38450 and n38207_not n38651_not ; n38706
g38451 and n38217_not n38613 ; n38707
g38452 and n38609_not n38707 ; n38708
g38453 and n38610_not n38613_not ; n38709
g38454 and n38708_not n38709_not ; n38710
g38455 and n10530 n38710_not ; n38711
g38456 and n38650_not n38711 ; n38712
g38457 and n38706_not n38712_not ; n38713
g38458 and b[31]_not n38713_not ; n38714
g38459 and n38216_not n38651_not ; n38715
g38460 and n38226_not n38608 ; n38716
g38461 and n38604_not n38716 ; n38717
g38462 and n38605_not n38608_not ; n38718
g38463 and n38717_not n38718_not ; n38719
g38464 and n10530 n38719_not ; n38720
g38465 and n38650_not n38720 ; n38721
g38466 and n38715_not n38721_not ; n38722
g38467 and b[30]_not n38722_not ; n38723
g38468 and n38225_not n38651_not ; n38724
g38469 and n38235_not n38603 ; n38725
g38470 and n38599_not n38725 ; n38726
g38471 and n38600_not n38603_not ; n38727
g38472 and n38726_not n38727_not ; n38728
g38473 and n10530 n38728_not ; n38729
g38474 and n38650_not n38729 ; n38730
g38475 and n38724_not n38730_not ; n38731
g38476 and b[29]_not n38731_not ; n38732
g38477 and n38234_not n38651_not ; n38733
g38478 and n38244_not n38598 ; n38734
g38479 and n38594_not n38734 ; n38735
g38480 and n38595_not n38598_not ; n38736
g38481 and n38735_not n38736_not ; n38737
g38482 and n10530 n38737_not ; n38738
g38483 and n38650_not n38738 ; n38739
g38484 and n38733_not n38739_not ; n38740
g38485 and b[28]_not n38740_not ; n38741
g38486 and n38243_not n38651_not ; n38742
g38487 and n38253_not n38593 ; n38743
g38488 and n38589_not n38743 ; n38744
g38489 and n38590_not n38593_not ; n38745
g38490 and n38744_not n38745_not ; n38746
g38491 and n10530 n38746_not ; n38747
g38492 and n38650_not n38747 ; n38748
g38493 and n38742_not n38748_not ; n38749
g38494 and b[27]_not n38749_not ; n38750
g38495 and n38252_not n38651_not ; n38751
g38496 and n38262_not n38588 ; n38752
g38497 and n38584_not n38752 ; n38753
g38498 and n38585_not n38588_not ; n38754
g38499 and n38753_not n38754_not ; n38755
g38500 and n10530 n38755_not ; n38756
g38501 and n38650_not n38756 ; n38757
g38502 and n38751_not n38757_not ; n38758
g38503 and b[26]_not n38758_not ; n38759
g38504 and n38261_not n38651_not ; n38760
g38505 and n38271_not n38583 ; n38761
g38506 and n38579_not n38761 ; n38762
g38507 and n38580_not n38583_not ; n38763
g38508 and n38762_not n38763_not ; n38764
g38509 and n10530 n38764_not ; n38765
g38510 and n38650_not n38765 ; n38766
g38511 and n38760_not n38766_not ; n38767
g38512 and b[25]_not n38767_not ; n38768
g38513 and n38270_not n38651_not ; n38769
g38514 and n38280_not n38578 ; n38770
g38515 and n38574_not n38770 ; n38771
g38516 and n38575_not n38578_not ; n38772
g38517 and n38771_not n38772_not ; n38773
g38518 and n10530 n38773_not ; n38774
g38519 and n38650_not n38774 ; n38775
g38520 and n38769_not n38775_not ; n38776
g38521 and b[24]_not n38776_not ; n38777
g38522 and n38279_not n38651_not ; n38778
g38523 and n38289_not n38573 ; n38779
g38524 and n38569_not n38779 ; n38780
g38525 and n38570_not n38573_not ; n38781
g38526 and n38780_not n38781_not ; n38782
g38527 and n10530 n38782_not ; n38783
g38528 and n38650_not n38783 ; n38784
g38529 and n38778_not n38784_not ; n38785
g38530 and b[23]_not n38785_not ; n38786
g38531 and n38288_not n38651_not ; n38787
g38532 and n38298_not n38568 ; n38788
g38533 and n38564_not n38788 ; n38789
g38534 and n38565_not n38568_not ; n38790
g38535 and n38789_not n38790_not ; n38791
g38536 and n10530 n38791_not ; n38792
g38537 and n38650_not n38792 ; n38793
g38538 and n38787_not n38793_not ; n38794
g38539 and b[22]_not n38794_not ; n38795
g38540 and n38297_not n38651_not ; n38796
g38541 and n38307_not n38563 ; n38797
g38542 and n38559_not n38797 ; n38798
g38543 and n38560_not n38563_not ; n38799
g38544 and n38798_not n38799_not ; n38800
g38545 and n10530 n38800_not ; n38801
g38546 and n38650_not n38801 ; n38802
g38547 and n38796_not n38802_not ; n38803
g38548 and b[21]_not n38803_not ; n38804
g38549 and n38306_not n38651_not ; n38805
g38550 and n38316_not n38558 ; n38806
g38551 and n38554_not n38806 ; n38807
g38552 and n38555_not n38558_not ; n38808
g38553 and n38807_not n38808_not ; n38809
g38554 and n10530 n38809_not ; n38810
g38555 and n38650_not n38810 ; n38811
g38556 and n38805_not n38811_not ; n38812
g38557 and b[20]_not n38812_not ; n38813
g38558 and n38315_not n38651_not ; n38814
g38559 and n38325_not n38553 ; n38815
g38560 and n38549_not n38815 ; n38816
g38561 and n38550_not n38553_not ; n38817
g38562 and n38816_not n38817_not ; n38818
g38563 and n10530 n38818_not ; n38819
g38564 and n38650_not n38819 ; n38820
g38565 and n38814_not n38820_not ; n38821
g38566 and b[19]_not n38821_not ; n38822
g38567 and n38324_not n38651_not ; n38823
g38568 and n38334_not n38548 ; n38824
g38569 and n38544_not n38824 ; n38825
g38570 and n38545_not n38548_not ; n38826
g38571 and n38825_not n38826_not ; n38827
g38572 and n10530 n38827_not ; n38828
g38573 and n38650_not n38828 ; n38829
g38574 and n38823_not n38829_not ; n38830
g38575 and b[18]_not n38830_not ; n38831
g38576 and n38333_not n38651_not ; n38832
g38577 and n38343_not n38543 ; n38833
g38578 and n38539_not n38833 ; n38834
g38579 and n38540_not n38543_not ; n38835
g38580 and n38834_not n38835_not ; n38836
g38581 and n10530 n38836_not ; n38837
g38582 and n38650_not n38837 ; n38838
g38583 and n38832_not n38838_not ; n38839
g38584 and b[17]_not n38839_not ; n38840
g38585 and n38342_not n38651_not ; n38841
g38586 and n38352_not n38538 ; n38842
g38587 and n38534_not n38842 ; n38843
g38588 and n38535_not n38538_not ; n38844
g38589 and n38843_not n38844_not ; n38845
g38590 and n10530 n38845_not ; n38846
g38591 and n38650_not n38846 ; n38847
g38592 and n38841_not n38847_not ; n38848
g38593 and b[16]_not n38848_not ; n38849
g38594 and n38351_not n38651_not ; n38850
g38595 and n38361_not n38533 ; n38851
g38596 and n38529_not n38851 ; n38852
g38597 and n38530_not n38533_not ; n38853
g38598 and n38852_not n38853_not ; n38854
g38599 and n10530 n38854_not ; n38855
g38600 and n38650_not n38855 ; n38856
g38601 and n38850_not n38856_not ; n38857
g38602 and b[15]_not n38857_not ; n38858
g38603 and n38360_not n38651_not ; n38859
g38604 and n38370_not n38528 ; n38860
g38605 and n38524_not n38860 ; n38861
g38606 and n38525_not n38528_not ; n38862
g38607 and n38861_not n38862_not ; n38863
g38608 and n10530 n38863_not ; n38864
g38609 and n38650_not n38864 ; n38865
g38610 and n38859_not n38865_not ; n38866
g38611 and b[14]_not n38866_not ; n38867
g38612 and n38369_not n38651_not ; n38868
g38613 and n38379_not n38523 ; n38869
g38614 and n38519_not n38869 ; n38870
g38615 and n38520_not n38523_not ; n38871
g38616 and n38870_not n38871_not ; n38872
g38617 and n10530 n38872_not ; n38873
g38618 and n38650_not n38873 ; n38874
g38619 and n38868_not n38874_not ; n38875
g38620 and b[13]_not n38875_not ; n38876
g38621 and n38378_not n38651_not ; n38877
g38622 and n38388_not n38518 ; n38878
g38623 and n38514_not n38878 ; n38879
g38624 and n38515_not n38518_not ; n38880
g38625 and n38879_not n38880_not ; n38881
g38626 and n10530 n38881_not ; n38882
g38627 and n38650_not n38882 ; n38883
g38628 and n38877_not n38883_not ; n38884
g38629 and b[12]_not n38884_not ; n38885
g38630 and n38387_not n38651_not ; n38886
g38631 and n38397_not n38513 ; n38887
g38632 and n38509_not n38887 ; n38888
g38633 and n38510_not n38513_not ; n38889
g38634 and n38888_not n38889_not ; n38890
g38635 and n10530 n38890_not ; n38891
g38636 and n38650_not n38891 ; n38892
g38637 and n38886_not n38892_not ; n38893
g38638 and b[11]_not n38893_not ; n38894
g38639 and n38396_not n38651_not ; n38895
g38640 and n38406_not n38508 ; n38896
g38641 and n38504_not n38896 ; n38897
g38642 and n38505_not n38508_not ; n38898
g38643 and n38897_not n38898_not ; n38899
g38644 and n10530 n38899_not ; n38900
g38645 and n38650_not n38900 ; n38901
g38646 and n38895_not n38901_not ; n38902
g38647 and b[10]_not n38902_not ; n38903
g38648 and n38405_not n38651_not ; n38904
g38649 and n38415_not n38503 ; n38905
g38650 and n38499_not n38905 ; n38906
g38651 and n38500_not n38503_not ; n38907
g38652 and n38906_not n38907_not ; n38908
g38653 and n10530 n38908_not ; n38909
g38654 and n38650_not n38909 ; n38910
g38655 and n38904_not n38910_not ; n38911
g38656 and b[9]_not n38911_not ; n38912
g38657 and n38414_not n38651_not ; n38913
g38658 and n38424_not n38498 ; n38914
g38659 and n38494_not n38914 ; n38915
g38660 and n38495_not n38498_not ; n38916
g38661 and n38915_not n38916_not ; n38917
g38662 and n10530 n38917_not ; n38918
g38663 and n38650_not n38918 ; n38919
g38664 and n38913_not n38919_not ; n38920
g38665 and b[8]_not n38920_not ; n38921
g38666 and n38423_not n38651_not ; n38922
g38667 and n38433_not n38493 ; n38923
g38668 and n38489_not n38923 ; n38924
g38669 and n38490_not n38493_not ; n38925
g38670 and n38924_not n38925_not ; n38926
g38671 and n10530 n38926_not ; n38927
g38672 and n38650_not n38927 ; n38928
g38673 and n38922_not n38928_not ; n38929
g38674 and b[7]_not n38929_not ; n38930
g38675 and n38432_not n38651_not ; n38931
g38676 and n38442_not n38488 ; n38932
g38677 and n38484_not n38932 ; n38933
g38678 and n38485_not n38488_not ; n38934
g38679 and n38933_not n38934_not ; n38935
g38680 and n10530 n38935_not ; n38936
g38681 and n38650_not n38936 ; n38937
g38682 and n38931_not n38937_not ; n38938
g38683 and b[6]_not n38938_not ; n38939
g38684 and n38441_not n38651_not ; n38940
g38685 and n38451_not n38483 ; n38941
g38686 and n38479_not n38941 ; n38942
g38687 and n38480_not n38483_not ; n38943
g38688 and n38942_not n38943_not ; n38944
g38689 and n10530 n38944_not ; n38945
g38690 and n38650_not n38945 ; n38946
g38691 and n38940_not n38946_not ; n38947
g38692 and b[5]_not n38947_not ; n38948
g38693 and n38450_not n38651_not ; n38949
g38694 and n38459_not n38478 ; n38950
g38695 and n38474_not n38950 ; n38951
g38696 and n38475_not n38478_not ; n38952
g38697 and n38951_not n38952_not ; n38953
g38698 and n10530 n38953_not ; n38954
g38699 and n38650_not n38954 ; n38955
g38700 and n38949_not n38955_not ; n38956
g38701 and b[4]_not n38956_not ; n38957
g38702 and n38458_not n38651_not ; n38958
g38703 and n38469_not n38473 ; n38959
g38704 and n38468_not n38959 ; n38960
g38705 and n38470_not n38473_not ; n38961
g38706 and n38960_not n38961_not ; n38962
g38707 and n10530 n38962_not ; n38963
g38708 and n38650_not n38963 ; n38964
g38709 and n38958_not n38964_not ; n38965
g38710 and b[3]_not n38965_not ; n38966
g38711 and n38463_not n38651_not ; n38967
g38712 and n10344 n38466_not ; n38968
g38713 and n38464_not n38968 ; n38969
g38714 and n10530 n38969_not ; n38970
g38715 and n38468_not n38970 ; n38971
g38716 and n38650_not n38971 ; n38972
g38717 and n38967_not n38972_not ; n38973
g38718 and b[2]_not n38973_not ; n38974
g38719 and n10859 n38650_not ; n38975
g38720 and a[26] n38975_not ; n38976
g38721 and n10865 n38650_not ; n38977
g38722 and n38976_not n38977_not ; n38978
g38723 and b[1] n38978_not ; n38979
g38724 and b[1]_not n38977_not ; n38980
g38725 and n38976_not n38980 ; n38981
g38726 and n38979_not n38981_not ; n38982
g38727 and n10872_not n38982_not ; n38983
g38728 and b[1]_not n38978_not ; n38984
g38729 and n38983_not n38984_not ; n38985
g38730 and b[2] n38972_not ; n38986
g38731 and n38967_not n38986 ; n38987
g38732 and n38974_not n38987_not ; n38988
g38733 and n38985_not n38988 ; n38989
g38734 and n38974_not n38989_not ; n38990
g38735 and b[3] n38964_not ; n38991
g38736 and n38958_not n38991 ; n38992
g38737 and n38966_not n38992_not ; n38993
g38738 and n38990_not n38993 ; n38994
g38739 and n38966_not n38994_not ; n38995
g38740 and b[4] n38955_not ; n38996
g38741 and n38949_not n38996 ; n38997
g38742 and n38957_not n38997_not ; n38998
g38743 and n38995_not n38998 ; n38999
g38744 and n38957_not n38999_not ; n39000
g38745 and b[5] n38946_not ; n39001
g38746 and n38940_not n39001 ; n39002
g38747 and n38948_not n39002_not ; n39003
g38748 and n39000_not n39003 ; n39004
g38749 and n38948_not n39004_not ; n39005
g38750 and b[6] n38937_not ; n39006
g38751 and n38931_not n39006 ; n39007
g38752 and n38939_not n39007_not ; n39008
g38753 and n39005_not n39008 ; n39009
g38754 and n38939_not n39009_not ; n39010
g38755 and b[7] n38928_not ; n39011
g38756 and n38922_not n39011 ; n39012
g38757 and n38930_not n39012_not ; n39013
g38758 and n39010_not n39013 ; n39014
g38759 and n38930_not n39014_not ; n39015
g38760 and b[8] n38919_not ; n39016
g38761 and n38913_not n39016 ; n39017
g38762 and n38921_not n39017_not ; n39018
g38763 and n39015_not n39018 ; n39019
g38764 and n38921_not n39019_not ; n39020
g38765 and b[9] n38910_not ; n39021
g38766 and n38904_not n39021 ; n39022
g38767 and n38912_not n39022_not ; n39023
g38768 and n39020_not n39023 ; n39024
g38769 and n38912_not n39024_not ; n39025
g38770 and b[10] n38901_not ; n39026
g38771 and n38895_not n39026 ; n39027
g38772 and n38903_not n39027_not ; n39028
g38773 and n39025_not n39028 ; n39029
g38774 and n38903_not n39029_not ; n39030
g38775 and b[11] n38892_not ; n39031
g38776 and n38886_not n39031 ; n39032
g38777 and n38894_not n39032_not ; n39033
g38778 and n39030_not n39033 ; n39034
g38779 and n38894_not n39034_not ; n39035
g38780 and b[12] n38883_not ; n39036
g38781 and n38877_not n39036 ; n39037
g38782 and n38885_not n39037_not ; n39038
g38783 and n39035_not n39038 ; n39039
g38784 and n38885_not n39039_not ; n39040
g38785 and b[13] n38874_not ; n39041
g38786 and n38868_not n39041 ; n39042
g38787 and n38876_not n39042_not ; n39043
g38788 and n39040_not n39043 ; n39044
g38789 and n38876_not n39044_not ; n39045
g38790 and b[14] n38865_not ; n39046
g38791 and n38859_not n39046 ; n39047
g38792 and n38867_not n39047_not ; n39048
g38793 and n39045_not n39048 ; n39049
g38794 and n38867_not n39049_not ; n39050
g38795 and b[15] n38856_not ; n39051
g38796 and n38850_not n39051 ; n39052
g38797 and n38858_not n39052_not ; n39053
g38798 and n39050_not n39053 ; n39054
g38799 and n38858_not n39054_not ; n39055
g38800 and b[16] n38847_not ; n39056
g38801 and n38841_not n39056 ; n39057
g38802 and n38849_not n39057_not ; n39058
g38803 and n39055_not n39058 ; n39059
g38804 and n38849_not n39059_not ; n39060
g38805 and b[17] n38838_not ; n39061
g38806 and n38832_not n39061 ; n39062
g38807 and n38840_not n39062_not ; n39063
g38808 and n39060_not n39063 ; n39064
g38809 and n38840_not n39064_not ; n39065
g38810 and b[18] n38829_not ; n39066
g38811 and n38823_not n39066 ; n39067
g38812 and n38831_not n39067_not ; n39068
g38813 and n39065_not n39068 ; n39069
g38814 and n38831_not n39069_not ; n39070
g38815 and b[19] n38820_not ; n39071
g38816 and n38814_not n39071 ; n39072
g38817 and n38822_not n39072_not ; n39073
g38818 and n39070_not n39073 ; n39074
g38819 and n38822_not n39074_not ; n39075
g38820 and b[20] n38811_not ; n39076
g38821 and n38805_not n39076 ; n39077
g38822 and n38813_not n39077_not ; n39078
g38823 and n39075_not n39078 ; n39079
g38824 and n38813_not n39079_not ; n39080
g38825 and b[21] n38802_not ; n39081
g38826 and n38796_not n39081 ; n39082
g38827 and n38804_not n39082_not ; n39083
g38828 and n39080_not n39083 ; n39084
g38829 and n38804_not n39084_not ; n39085
g38830 and b[22] n38793_not ; n39086
g38831 and n38787_not n39086 ; n39087
g38832 and n38795_not n39087_not ; n39088
g38833 and n39085_not n39088 ; n39089
g38834 and n38795_not n39089_not ; n39090
g38835 and b[23] n38784_not ; n39091
g38836 and n38778_not n39091 ; n39092
g38837 and n38786_not n39092_not ; n39093
g38838 and n39090_not n39093 ; n39094
g38839 and n38786_not n39094_not ; n39095
g38840 and b[24] n38775_not ; n39096
g38841 and n38769_not n39096 ; n39097
g38842 and n38777_not n39097_not ; n39098
g38843 and n39095_not n39098 ; n39099
g38844 and n38777_not n39099_not ; n39100
g38845 and b[25] n38766_not ; n39101
g38846 and n38760_not n39101 ; n39102
g38847 and n38768_not n39102_not ; n39103
g38848 and n39100_not n39103 ; n39104
g38849 and n38768_not n39104_not ; n39105
g38850 and b[26] n38757_not ; n39106
g38851 and n38751_not n39106 ; n39107
g38852 and n38759_not n39107_not ; n39108
g38853 and n39105_not n39108 ; n39109
g38854 and n38759_not n39109_not ; n39110
g38855 and b[27] n38748_not ; n39111
g38856 and n38742_not n39111 ; n39112
g38857 and n38750_not n39112_not ; n39113
g38858 and n39110_not n39113 ; n39114
g38859 and n38750_not n39114_not ; n39115
g38860 and b[28] n38739_not ; n39116
g38861 and n38733_not n39116 ; n39117
g38862 and n38741_not n39117_not ; n39118
g38863 and n39115_not n39118 ; n39119
g38864 and n38741_not n39119_not ; n39120
g38865 and b[29] n38730_not ; n39121
g38866 and n38724_not n39121 ; n39122
g38867 and n38732_not n39122_not ; n39123
g38868 and n39120_not n39123 ; n39124
g38869 and n38732_not n39124_not ; n39125
g38870 and b[30] n38721_not ; n39126
g38871 and n38715_not n39126 ; n39127
g38872 and n38723_not n39127_not ; n39128
g38873 and n39125_not n39128 ; n39129
g38874 and n38723_not n39129_not ; n39130
g38875 and b[31] n38712_not ; n39131
g38876 and n38706_not n39131 ; n39132
g38877 and n38714_not n39132_not ; n39133
g38878 and n39130_not n39133 ; n39134
g38879 and n38714_not n39134_not ; n39135
g38880 and b[32] n38703_not ; n39136
g38881 and n38697_not n39136 ; n39137
g38882 and n38705_not n39137_not ; n39138
g38883 and n39135_not n39138 ; n39139
g38884 and n38705_not n39139_not ; n39140
g38885 and b[33] n38694_not ; n39141
g38886 and n38688_not n39141 ; n39142
g38887 and n38696_not n39142_not ; n39143
g38888 and n39140_not n39143 ; n39144
g38889 and n38696_not n39144_not ; n39145
g38890 and b[34] n38685_not ; n39146
g38891 and n38679_not n39146 ; n39147
g38892 and n38687_not n39147_not ; n39148
g38893 and n39145_not n39148 ; n39149
g38894 and n38687_not n39149_not ; n39150
g38895 and b[35] n38676_not ; n39151
g38896 and n38670_not n39151 ; n39152
g38897 and n38678_not n39152_not ; n39153
g38898 and n39150_not n39153 ; n39154
g38899 and n38678_not n39154_not ; n39155
g38900 and b[36] n38667_not ; n39156
g38901 and n38661_not n39156 ; n39157
g38902 and n38669_not n39157_not ; n39158
g38903 and n39155_not n39158 ; n39159
g38904 and n38669_not n39159_not ; n39160
g38905 and b[37] n38658_not ; n39161
g38906 and n38652_not n39161 ; n39162
g38907 and n38660_not n39162_not ; n39163
g38908 and n39160_not n39163 ; n39164
g38909 and n38660_not n39164_not ; n39165
g38910 and n38152_not n38651_not ; n39166
g38911 and n38154_not n38648 ; n39167
g38912 and n38644_not n39167 ; n39168
g38913 and n38645_not n38648_not ; n39169
g38914 and n39168_not n39169_not ; n39170
g38915 and n38651 n39170_not ; n39171
g38916 and n39166_not n39171_not ; n39172
g38917 and b[38]_not n39172_not ; n39173
g38918 and b[38] n39166_not ; n39174
g38919 and n39171_not n39174 ; n39175
g38920 and n11068 n39175_not ; n39176
g38921 and n39173_not n39176 ; n39177
g38922 and n39165_not n39177 ; n39178
g38923 and n10530 n39172_not ; n39179
g38924 and n39178_not n39179_not ; n39180
g38925 and n38669_not n39163 ; n39181
g38926 and n39159_not n39181 ; n39182
g38927 and n39160_not n39163_not ; n39183
g38928 and n39182_not n39183_not ; n39184
g38929 and n39180_not n39184_not ; n39185
g38930 and n38659_not n39179_not ; n39186
g38931 and n39178_not n39186 ; n39187
g38932 and n39185_not n39187_not ; n39188
g38933 and n38660_not n39175_not ; n39189
g38934 and n39173_not n39189 ; n39190
g38935 and n39164_not n39190 ; n39191
g38936 and n39173_not n39175_not ; n39192
g38937 and n39165_not n39192_not ; n39193
g38938 and n39191_not n39193_not ; n39194
g38939 and n39180_not n39194_not ; n39195
g38940 and n39172_not n39179_not ; n39196
g38941 and n39178_not n39196 ; n39197
g38942 and n39195_not n39197_not ; n39198
g38943 and b[39]_not n39198_not ; n39199
g38944 and b[38]_not n39188_not ; n39200
g38945 and n38678_not n39158 ; n39201
g38946 and n39154_not n39201 ; n39202
g38947 and n39155_not n39158_not ; n39203
g38948 and n39202_not n39203_not ; n39204
g38949 and n39180_not n39204_not ; n39205
g38950 and n38668_not n39179_not ; n39206
g38951 and n39178_not n39206 ; n39207
g38952 and n39205_not n39207_not ; n39208
g38953 and b[37]_not n39208_not ; n39209
g38954 and n38687_not n39153 ; n39210
g38955 and n39149_not n39210 ; n39211
g38956 and n39150_not n39153_not ; n39212
g38957 and n39211_not n39212_not ; n39213
g38958 and n39180_not n39213_not ; n39214
g38959 and n38677_not n39179_not ; n39215
g38960 and n39178_not n39215 ; n39216
g38961 and n39214_not n39216_not ; n39217
g38962 and b[36]_not n39217_not ; n39218
g38963 and n38696_not n39148 ; n39219
g38964 and n39144_not n39219 ; n39220
g38965 and n39145_not n39148_not ; n39221
g38966 and n39220_not n39221_not ; n39222
g38967 and n39180_not n39222_not ; n39223
g38968 and n38686_not n39179_not ; n39224
g38969 and n39178_not n39224 ; n39225
g38970 and n39223_not n39225_not ; n39226
g38971 and b[35]_not n39226_not ; n39227
g38972 and n38705_not n39143 ; n39228
g38973 and n39139_not n39228 ; n39229
g38974 and n39140_not n39143_not ; n39230
g38975 and n39229_not n39230_not ; n39231
g38976 and n39180_not n39231_not ; n39232
g38977 and n38695_not n39179_not ; n39233
g38978 and n39178_not n39233 ; n39234
g38979 and n39232_not n39234_not ; n39235
g38980 and b[34]_not n39235_not ; n39236
g38981 and n38714_not n39138 ; n39237
g38982 and n39134_not n39237 ; n39238
g38983 and n39135_not n39138_not ; n39239
g38984 and n39238_not n39239_not ; n39240
g38985 and n39180_not n39240_not ; n39241
g38986 and n38704_not n39179_not ; n39242
g38987 and n39178_not n39242 ; n39243
g38988 and n39241_not n39243_not ; n39244
g38989 and b[33]_not n39244_not ; n39245
g38990 and n38723_not n39133 ; n39246
g38991 and n39129_not n39246 ; n39247
g38992 and n39130_not n39133_not ; n39248
g38993 and n39247_not n39248_not ; n39249
g38994 and n39180_not n39249_not ; n39250
g38995 and n38713_not n39179_not ; n39251
g38996 and n39178_not n39251 ; n39252
g38997 and n39250_not n39252_not ; n39253
g38998 and b[32]_not n39253_not ; n39254
g38999 and n38732_not n39128 ; n39255
g39000 and n39124_not n39255 ; n39256
g39001 and n39125_not n39128_not ; n39257
g39002 and n39256_not n39257_not ; n39258
g39003 and n39180_not n39258_not ; n39259
g39004 and n38722_not n39179_not ; n39260
g39005 and n39178_not n39260 ; n39261
g39006 and n39259_not n39261_not ; n39262
g39007 and b[31]_not n39262_not ; n39263
g39008 and n38741_not n39123 ; n39264
g39009 and n39119_not n39264 ; n39265
g39010 and n39120_not n39123_not ; n39266
g39011 and n39265_not n39266_not ; n39267
g39012 and n39180_not n39267_not ; n39268
g39013 and n38731_not n39179_not ; n39269
g39014 and n39178_not n39269 ; n39270
g39015 and n39268_not n39270_not ; n39271
g39016 and b[30]_not n39271_not ; n39272
g39017 and n38750_not n39118 ; n39273
g39018 and n39114_not n39273 ; n39274
g39019 and n39115_not n39118_not ; n39275
g39020 and n39274_not n39275_not ; n39276
g39021 and n39180_not n39276_not ; n39277
g39022 and n38740_not n39179_not ; n39278
g39023 and n39178_not n39278 ; n39279
g39024 and n39277_not n39279_not ; n39280
g39025 and b[29]_not n39280_not ; n39281
g39026 and n38759_not n39113 ; n39282
g39027 and n39109_not n39282 ; n39283
g39028 and n39110_not n39113_not ; n39284
g39029 and n39283_not n39284_not ; n39285
g39030 and n39180_not n39285_not ; n39286
g39031 and n38749_not n39179_not ; n39287
g39032 and n39178_not n39287 ; n39288
g39033 and n39286_not n39288_not ; n39289
g39034 and b[28]_not n39289_not ; n39290
g39035 and n38768_not n39108 ; n39291
g39036 and n39104_not n39291 ; n39292
g39037 and n39105_not n39108_not ; n39293
g39038 and n39292_not n39293_not ; n39294
g39039 and n39180_not n39294_not ; n39295
g39040 and n38758_not n39179_not ; n39296
g39041 and n39178_not n39296 ; n39297
g39042 and n39295_not n39297_not ; n39298
g39043 and b[27]_not n39298_not ; n39299
g39044 and n38777_not n39103 ; n39300
g39045 and n39099_not n39300 ; n39301
g39046 and n39100_not n39103_not ; n39302
g39047 and n39301_not n39302_not ; n39303
g39048 and n39180_not n39303_not ; n39304
g39049 and n38767_not n39179_not ; n39305
g39050 and n39178_not n39305 ; n39306
g39051 and n39304_not n39306_not ; n39307
g39052 and b[26]_not n39307_not ; n39308
g39053 and n38786_not n39098 ; n39309
g39054 and n39094_not n39309 ; n39310
g39055 and n39095_not n39098_not ; n39311
g39056 and n39310_not n39311_not ; n39312
g39057 and n39180_not n39312_not ; n39313
g39058 and n38776_not n39179_not ; n39314
g39059 and n39178_not n39314 ; n39315
g39060 and n39313_not n39315_not ; n39316
g39061 and b[25]_not n39316_not ; n39317
g39062 and n38795_not n39093 ; n39318
g39063 and n39089_not n39318 ; n39319
g39064 and n39090_not n39093_not ; n39320
g39065 and n39319_not n39320_not ; n39321
g39066 and n39180_not n39321_not ; n39322
g39067 and n38785_not n39179_not ; n39323
g39068 and n39178_not n39323 ; n39324
g39069 and n39322_not n39324_not ; n39325
g39070 and b[24]_not n39325_not ; n39326
g39071 and n38804_not n39088 ; n39327
g39072 and n39084_not n39327 ; n39328
g39073 and n39085_not n39088_not ; n39329
g39074 and n39328_not n39329_not ; n39330
g39075 and n39180_not n39330_not ; n39331
g39076 and n38794_not n39179_not ; n39332
g39077 and n39178_not n39332 ; n39333
g39078 and n39331_not n39333_not ; n39334
g39079 and b[23]_not n39334_not ; n39335
g39080 and n38813_not n39083 ; n39336
g39081 and n39079_not n39336 ; n39337
g39082 and n39080_not n39083_not ; n39338
g39083 and n39337_not n39338_not ; n39339
g39084 and n39180_not n39339_not ; n39340
g39085 and n38803_not n39179_not ; n39341
g39086 and n39178_not n39341 ; n39342
g39087 and n39340_not n39342_not ; n39343
g39088 and b[22]_not n39343_not ; n39344
g39089 and n38822_not n39078 ; n39345
g39090 and n39074_not n39345 ; n39346
g39091 and n39075_not n39078_not ; n39347
g39092 and n39346_not n39347_not ; n39348
g39093 and n39180_not n39348_not ; n39349
g39094 and n38812_not n39179_not ; n39350
g39095 and n39178_not n39350 ; n39351
g39096 and n39349_not n39351_not ; n39352
g39097 and b[21]_not n39352_not ; n39353
g39098 and n38831_not n39073 ; n39354
g39099 and n39069_not n39354 ; n39355
g39100 and n39070_not n39073_not ; n39356
g39101 and n39355_not n39356_not ; n39357
g39102 and n39180_not n39357_not ; n39358
g39103 and n38821_not n39179_not ; n39359
g39104 and n39178_not n39359 ; n39360
g39105 and n39358_not n39360_not ; n39361
g39106 and b[20]_not n39361_not ; n39362
g39107 and n38840_not n39068 ; n39363
g39108 and n39064_not n39363 ; n39364
g39109 and n39065_not n39068_not ; n39365
g39110 and n39364_not n39365_not ; n39366
g39111 and n39180_not n39366_not ; n39367
g39112 and n38830_not n39179_not ; n39368
g39113 and n39178_not n39368 ; n39369
g39114 and n39367_not n39369_not ; n39370
g39115 and b[19]_not n39370_not ; n39371
g39116 and n38849_not n39063 ; n39372
g39117 and n39059_not n39372 ; n39373
g39118 and n39060_not n39063_not ; n39374
g39119 and n39373_not n39374_not ; n39375
g39120 and n39180_not n39375_not ; n39376
g39121 and n38839_not n39179_not ; n39377
g39122 and n39178_not n39377 ; n39378
g39123 and n39376_not n39378_not ; n39379
g39124 and b[18]_not n39379_not ; n39380
g39125 and n38858_not n39058 ; n39381
g39126 and n39054_not n39381 ; n39382
g39127 and n39055_not n39058_not ; n39383
g39128 and n39382_not n39383_not ; n39384
g39129 and n39180_not n39384_not ; n39385
g39130 and n38848_not n39179_not ; n39386
g39131 and n39178_not n39386 ; n39387
g39132 and n39385_not n39387_not ; n39388
g39133 and b[17]_not n39388_not ; n39389
g39134 and n38867_not n39053 ; n39390
g39135 and n39049_not n39390 ; n39391
g39136 and n39050_not n39053_not ; n39392
g39137 and n39391_not n39392_not ; n39393
g39138 and n39180_not n39393_not ; n39394
g39139 and n38857_not n39179_not ; n39395
g39140 and n39178_not n39395 ; n39396
g39141 and n39394_not n39396_not ; n39397
g39142 and b[16]_not n39397_not ; n39398
g39143 and n38876_not n39048 ; n39399
g39144 and n39044_not n39399 ; n39400
g39145 and n39045_not n39048_not ; n39401
g39146 and n39400_not n39401_not ; n39402
g39147 and n39180_not n39402_not ; n39403
g39148 and n38866_not n39179_not ; n39404
g39149 and n39178_not n39404 ; n39405
g39150 and n39403_not n39405_not ; n39406
g39151 and b[15]_not n39406_not ; n39407
g39152 and n38885_not n39043 ; n39408
g39153 and n39039_not n39408 ; n39409
g39154 and n39040_not n39043_not ; n39410
g39155 and n39409_not n39410_not ; n39411
g39156 and n39180_not n39411_not ; n39412
g39157 and n38875_not n39179_not ; n39413
g39158 and n39178_not n39413 ; n39414
g39159 and n39412_not n39414_not ; n39415
g39160 and b[14]_not n39415_not ; n39416
g39161 and n38894_not n39038 ; n39417
g39162 and n39034_not n39417 ; n39418
g39163 and n39035_not n39038_not ; n39419
g39164 and n39418_not n39419_not ; n39420
g39165 and n39180_not n39420_not ; n39421
g39166 and n38884_not n39179_not ; n39422
g39167 and n39178_not n39422 ; n39423
g39168 and n39421_not n39423_not ; n39424
g39169 and b[13]_not n39424_not ; n39425
g39170 and n38903_not n39033 ; n39426
g39171 and n39029_not n39426 ; n39427
g39172 and n39030_not n39033_not ; n39428
g39173 and n39427_not n39428_not ; n39429
g39174 and n39180_not n39429_not ; n39430
g39175 and n38893_not n39179_not ; n39431
g39176 and n39178_not n39431 ; n39432
g39177 and n39430_not n39432_not ; n39433
g39178 and b[12]_not n39433_not ; n39434
g39179 and n38912_not n39028 ; n39435
g39180 and n39024_not n39435 ; n39436
g39181 and n39025_not n39028_not ; n39437
g39182 and n39436_not n39437_not ; n39438
g39183 and n39180_not n39438_not ; n39439
g39184 and n38902_not n39179_not ; n39440
g39185 and n39178_not n39440 ; n39441
g39186 and n39439_not n39441_not ; n39442
g39187 and b[11]_not n39442_not ; n39443
g39188 and n38921_not n39023 ; n39444
g39189 and n39019_not n39444 ; n39445
g39190 and n39020_not n39023_not ; n39446
g39191 and n39445_not n39446_not ; n39447
g39192 and n39180_not n39447_not ; n39448
g39193 and n38911_not n39179_not ; n39449
g39194 and n39178_not n39449 ; n39450
g39195 and n39448_not n39450_not ; n39451
g39196 and b[10]_not n39451_not ; n39452
g39197 and n38930_not n39018 ; n39453
g39198 and n39014_not n39453 ; n39454
g39199 and n39015_not n39018_not ; n39455
g39200 and n39454_not n39455_not ; n39456
g39201 and n39180_not n39456_not ; n39457
g39202 and n38920_not n39179_not ; n39458
g39203 and n39178_not n39458 ; n39459
g39204 and n39457_not n39459_not ; n39460
g39205 and b[9]_not n39460_not ; n39461
g39206 and n38939_not n39013 ; n39462
g39207 and n39009_not n39462 ; n39463
g39208 and n39010_not n39013_not ; n39464
g39209 and n39463_not n39464_not ; n39465
g39210 and n39180_not n39465_not ; n39466
g39211 and n38929_not n39179_not ; n39467
g39212 and n39178_not n39467 ; n39468
g39213 and n39466_not n39468_not ; n39469
g39214 and b[8]_not n39469_not ; n39470
g39215 and n38948_not n39008 ; n39471
g39216 and n39004_not n39471 ; n39472
g39217 and n39005_not n39008_not ; n39473
g39218 and n39472_not n39473_not ; n39474
g39219 and n39180_not n39474_not ; n39475
g39220 and n38938_not n39179_not ; n39476
g39221 and n39178_not n39476 ; n39477
g39222 and n39475_not n39477_not ; n39478
g39223 and b[7]_not n39478_not ; n39479
g39224 and n38957_not n39003 ; n39480
g39225 and n38999_not n39480 ; n39481
g39226 and n39000_not n39003_not ; n39482
g39227 and n39481_not n39482_not ; n39483
g39228 and n39180_not n39483_not ; n39484
g39229 and n38947_not n39179_not ; n39485
g39230 and n39178_not n39485 ; n39486
g39231 and n39484_not n39486_not ; n39487
g39232 and b[6]_not n39487_not ; n39488
g39233 and n38966_not n38998 ; n39489
g39234 and n38994_not n39489 ; n39490
g39235 and n38995_not n38998_not ; n39491
g39236 and n39490_not n39491_not ; n39492
g39237 and n39180_not n39492_not ; n39493
g39238 and n38956_not n39179_not ; n39494
g39239 and n39178_not n39494 ; n39495
g39240 and n39493_not n39495_not ; n39496
g39241 and b[5]_not n39496_not ; n39497
g39242 and n38974_not n38993 ; n39498
g39243 and n38989_not n39498 ; n39499
g39244 and n38990_not n38993_not ; n39500
g39245 and n39499_not n39500_not ; n39501
g39246 and n39180_not n39501_not ; n39502
g39247 and n38965_not n39179_not ; n39503
g39248 and n39178_not n39503 ; n39504
g39249 and n39502_not n39504_not ; n39505
g39250 and b[4]_not n39505_not ; n39506
g39251 and n38984_not n38988 ; n39507
g39252 and n38983_not n39507 ; n39508
g39253 and n38985_not n38988_not ; n39509
g39254 and n39508_not n39509_not ; n39510
g39255 and n39180_not n39510_not ; n39511
g39256 and n38973_not n39179_not ; n39512
g39257 and n39178_not n39512 ; n39513
g39258 and n39511_not n39513_not ; n39514
g39259 and b[3]_not n39514_not ; n39515
g39260 and n10872 n38981_not ; n39516
g39261 and n38979_not n39516 ; n39517
g39262 and n38983_not n39517_not ; n39518
g39263 and n39180_not n39518 ; n39519
g39264 and n38978_not n39179_not ; n39520
g39265 and n39178_not n39520 ; n39521
g39266 and n39519_not n39521_not ; n39522
g39267 and b[2]_not n39522_not ; n39523
g39268 and b[0] n39180_not ; n39524
g39269 and a[25] n39524_not ; n39525
g39270 and n10872 n39180_not ; n39526
g39271 and n39525_not n39526_not ; n39527
g39272 and b[1] n39527_not ; n39528
g39273 and b[1]_not n39526_not ; n39529
g39274 and n39525_not n39529 ; n39530
g39275 and n39528_not n39530_not ; n39531
g39276 and n11425_not n39531_not ; n39532
g39277 and b[1]_not n39527_not ; n39533
g39278 and n39532_not n39533_not ; n39534
g39279 and b[2] n39521_not ; n39535
g39280 and n39519_not n39535 ; n39536
g39281 and n39523_not n39536_not ; n39537
g39282 and n39534_not n39537 ; n39538
g39283 and n39523_not n39538_not ; n39539
g39284 and b[3] n39513_not ; n39540
g39285 and n39511_not n39540 ; n39541
g39286 and n39515_not n39541_not ; n39542
g39287 and n39539_not n39542 ; n39543
g39288 and n39515_not n39543_not ; n39544
g39289 and b[4] n39504_not ; n39545
g39290 and n39502_not n39545 ; n39546
g39291 and n39506_not n39546_not ; n39547
g39292 and n39544_not n39547 ; n39548
g39293 and n39506_not n39548_not ; n39549
g39294 and b[5] n39495_not ; n39550
g39295 and n39493_not n39550 ; n39551
g39296 and n39497_not n39551_not ; n39552
g39297 and n39549_not n39552 ; n39553
g39298 and n39497_not n39553_not ; n39554
g39299 and b[6] n39486_not ; n39555
g39300 and n39484_not n39555 ; n39556
g39301 and n39488_not n39556_not ; n39557
g39302 and n39554_not n39557 ; n39558
g39303 and n39488_not n39558_not ; n39559
g39304 and b[7] n39477_not ; n39560
g39305 and n39475_not n39560 ; n39561
g39306 and n39479_not n39561_not ; n39562
g39307 and n39559_not n39562 ; n39563
g39308 and n39479_not n39563_not ; n39564
g39309 and b[8] n39468_not ; n39565
g39310 and n39466_not n39565 ; n39566
g39311 and n39470_not n39566_not ; n39567
g39312 and n39564_not n39567 ; n39568
g39313 and n39470_not n39568_not ; n39569
g39314 and b[9] n39459_not ; n39570
g39315 and n39457_not n39570 ; n39571
g39316 and n39461_not n39571_not ; n39572
g39317 and n39569_not n39572 ; n39573
g39318 and n39461_not n39573_not ; n39574
g39319 and b[10] n39450_not ; n39575
g39320 and n39448_not n39575 ; n39576
g39321 and n39452_not n39576_not ; n39577
g39322 and n39574_not n39577 ; n39578
g39323 and n39452_not n39578_not ; n39579
g39324 and b[11] n39441_not ; n39580
g39325 and n39439_not n39580 ; n39581
g39326 and n39443_not n39581_not ; n39582
g39327 and n39579_not n39582 ; n39583
g39328 and n39443_not n39583_not ; n39584
g39329 and b[12] n39432_not ; n39585
g39330 and n39430_not n39585 ; n39586
g39331 and n39434_not n39586_not ; n39587
g39332 and n39584_not n39587 ; n39588
g39333 and n39434_not n39588_not ; n39589
g39334 and b[13] n39423_not ; n39590
g39335 and n39421_not n39590 ; n39591
g39336 and n39425_not n39591_not ; n39592
g39337 and n39589_not n39592 ; n39593
g39338 and n39425_not n39593_not ; n39594
g39339 and b[14] n39414_not ; n39595
g39340 and n39412_not n39595 ; n39596
g39341 and n39416_not n39596_not ; n39597
g39342 and n39594_not n39597 ; n39598
g39343 and n39416_not n39598_not ; n39599
g39344 and b[15] n39405_not ; n39600
g39345 and n39403_not n39600 ; n39601
g39346 and n39407_not n39601_not ; n39602
g39347 and n39599_not n39602 ; n39603
g39348 and n39407_not n39603_not ; n39604
g39349 and b[16] n39396_not ; n39605
g39350 and n39394_not n39605 ; n39606
g39351 and n39398_not n39606_not ; n39607
g39352 and n39604_not n39607 ; n39608
g39353 and n39398_not n39608_not ; n39609
g39354 and b[17] n39387_not ; n39610
g39355 and n39385_not n39610 ; n39611
g39356 and n39389_not n39611_not ; n39612
g39357 and n39609_not n39612 ; n39613
g39358 and n39389_not n39613_not ; n39614
g39359 and b[18] n39378_not ; n39615
g39360 and n39376_not n39615 ; n39616
g39361 and n39380_not n39616_not ; n39617
g39362 and n39614_not n39617 ; n39618
g39363 and n39380_not n39618_not ; n39619
g39364 and b[19] n39369_not ; n39620
g39365 and n39367_not n39620 ; n39621
g39366 and n39371_not n39621_not ; n39622
g39367 and n39619_not n39622 ; n39623
g39368 and n39371_not n39623_not ; n39624
g39369 and b[20] n39360_not ; n39625
g39370 and n39358_not n39625 ; n39626
g39371 and n39362_not n39626_not ; n39627
g39372 and n39624_not n39627 ; n39628
g39373 and n39362_not n39628_not ; n39629
g39374 and b[21] n39351_not ; n39630
g39375 and n39349_not n39630 ; n39631
g39376 and n39353_not n39631_not ; n39632
g39377 and n39629_not n39632 ; n39633
g39378 and n39353_not n39633_not ; n39634
g39379 and b[22] n39342_not ; n39635
g39380 and n39340_not n39635 ; n39636
g39381 and n39344_not n39636_not ; n39637
g39382 and n39634_not n39637 ; n39638
g39383 and n39344_not n39638_not ; n39639
g39384 and b[23] n39333_not ; n39640
g39385 and n39331_not n39640 ; n39641
g39386 and n39335_not n39641_not ; n39642
g39387 and n39639_not n39642 ; n39643
g39388 and n39335_not n39643_not ; n39644
g39389 and b[24] n39324_not ; n39645
g39390 and n39322_not n39645 ; n39646
g39391 and n39326_not n39646_not ; n39647
g39392 and n39644_not n39647 ; n39648
g39393 and n39326_not n39648_not ; n39649
g39394 and b[25] n39315_not ; n39650
g39395 and n39313_not n39650 ; n39651
g39396 and n39317_not n39651_not ; n39652
g39397 and n39649_not n39652 ; n39653
g39398 and n39317_not n39653_not ; n39654
g39399 and b[26] n39306_not ; n39655
g39400 and n39304_not n39655 ; n39656
g39401 and n39308_not n39656_not ; n39657
g39402 and n39654_not n39657 ; n39658
g39403 and n39308_not n39658_not ; n39659
g39404 and b[27] n39297_not ; n39660
g39405 and n39295_not n39660 ; n39661
g39406 and n39299_not n39661_not ; n39662
g39407 and n39659_not n39662 ; n39663
g39408 and n39299_not n39663_not ; n39664
g39409 and b[28] n39288_not ; n39665
g39410 and n39286_not n39665 ; n39666
g39411 and n39290_not n39666_not ; n39667
g39412 and n39664_not n39667 ; n39668
g39413 and n39290_not n39668_not ; n39669
g39414 and b[29] n39279_not ; n39670
g39415 and n39277_not n39670 ; n39671
g39416 and n39281_not n39671_not ; n39672
g39417 and n39669_not n39672 ; n39673
g39418 and n39281_not n39673_not ; n39674
g39419 and b[30] n39270_not ; n39675
g39420 and n39268_not n39675 ; n39676
g39421 and n39272_not n39676_not ; n39677
g39422 and n39674_not n39677 ; n39678
g39423 and n39272_not n39678_not ; n39679
g39424 and b[31] n39261_not ; n39680
g39425 and n39259_not n39680 ; n39681
g39426 and n39263_not n39681_not ; n39682
g39427 and n39679_not n39682 ; n39683
g39428 and n39263_not n39683_not ; n39684
g39429 and b[32] n39252_not ; n39685
g39430 and n39250_not n39685 ; n39686
g39431 and n39254_not n39686_not ; n39687
g39432 and n39684_not n39687 ; n39688
g39433 and n39254_not n39688_not ; n39689
g39434 and b[33] n39243_not ; n39690
g39435 and n39241_not n39690 ; n39691
g39436 and n39245_not n39691_not ; n39692
g39437 and n39689_not n39692 ; n39693
g39438 and n39245_not n39693_not ; n39694
g39439 and b[34] n39234_not ; n39695
g39440 and n39232_not n39695 ; n39696
g39441 and n39236_not n39696_not ; n39697
g39442 and n39694_not n39697 ; n39698
g39443 and n39236_not n39698_not ; n39699
g39444 and b[35] n39225_not ; n39700
g39445 and n39223_not n39700 ; n39701
g39446 and n39227_not n39701_not ; n39702
g39447 and n39699_not n39702 ; n39703
g39448 and n39227_not n39703_not ; n39704
g39449 and b[36] n39216_not ; n39705
g39450 and n39214_not n39705 ; n39706
g39451 and n39218_not n39706_not ; n39707
g39452 and n39704_not n39707 ; n39708
g39453 and n39218_not n39708_not ; n39709
g39454 and b[37] n39207_not ; n39710
g39455 and n39205_not n39710 ; n39711
g39456 and n39209_not n39711_not ; n39712
g39457 and n39709_not n39712 ; n39713
g39458 and n39209_not n39713_not ; n39714
g39459 and b[38] n39187_not ; n39715
g39460 and n39185_not n39715 ; n39716
g39461 and n39200_not n39716_not ; n39717
g39462 and n39714_not n39717 ; n39718
g39463 and n39200_not n39718_not ; n39719
g39464 and b[39] n39197_not ; n39720
g39465 and n39195_not n39720 ; n39721
g39466 and n39199_not n39721_not ; n39722
g39467 and n39719_not n39722 ; n39723
g39468 and n39199_not n39723_not ; n39724
g39469 and n11619 n39724_not ; n39725
g39470 and n39188_not n39725_not ; n39726
g39471 and n39209_not n39717 ; n39727
g39472 and n39713_not n39727 ; n39728
g39473 and n39714_not n39717_not ; n39729
g39474 and n39728_not n39729_not ; n39730
g39475 and n11619 n39730_not ; n39731
g39476 and n39724_not n39731 ; n39732
g39477 and n39726_not n39732_not ; n39733
g39478 and n39198_not n39725_not ; n39734
g39479 and n39200_not n39722 ; n39735
g39480 and n39718_not n39735 ; n39736
g39481 and n39719_not n39722_not ; n39737
g39482 and n39736_not n39737_not ; n39738
g39483 and n39725 n39738_not ; n39739
g39484 and n39734_not n39739_not ; n39740
g39485 and b[40]_not n39740_not ; n39741
g39486 and b[39]_not n39733_not ; n39742
g39487 and n39208_not n39725_not ; n39743
g39488 and n39218_not n39712 ; n39744
g39489 and n39708_not n39744 ; n39745
g39490 and n39709_not n39712_not ; n39746
g39491 and n39745_not n39746_not ; n39747
g39492 and n11619 n39747_not ; n39748
g39493 and n39724_not n39748 ; n39749
g39494 and n39743_not n39749_not ; n39750
g39495 and b[38]_not n39750_not ; n39751
g39496 and n39217_not n39725_not ; n39752
g39497 and n39227_not n39707 ; n39753
g39498 and n39703_not n39753 ; n39754
g39499 and n39704_not n39707_not ; n39755
g39500 and n39754_not n39755_not ; n39756
g39501 and n11619 n39756_not ; n39757
g39502 and n39724_not n39757 ; n39758
g39503 and n39752_not n39758_not ; n39759
g39504 and b[37]_not n39759_not ; n39760
g39505 and n39226_not n39725_not ; n39761
g39506 and n39236_not n39702 ; n39762
g39507 and n39698_not n39762 ; n39763
g39508 and n39699_not n39702_not ; n39764
g39509 and n39763_not n39764_not ; n39765
g39510 and n11619 n39765_not ; n39766
g39511 and n39724_not n39766 ; n39767
g39512 and n39761_not n39767_not ; n39768
g39513 and b[36]_not n39768_not ; n39769
g39514 and n39235_not n39725_not ; n39770
g39515 and n39245_not n39697 ; n39771
g39516 and n39693_not n39771 ; n39772
g39517 and n39694_not n39697_not ; n39773
g39518 and n39772_not n39773_not ; n39774
g39519 and n11619 n39774_not ; n39775
g39520 and n39724_not n39775 ; n39776
g39521 and n39770_not n39776_not ; n39777
g39522 and b[35]_not n39777_not ; n39778
g39523 and n39244_not n39725_not ; n39779
g39524 and n39254_not n39692 ; n39780
g39525 and n39688_not n39780 ; n39781
g39526 and n39689_not n39692_not ; n39782
g39527 and n39781_not n39782_not ; n39783
g39528 and n11619 n39783_not ; n39784
g39529 and n39724_not n39784 ; n39785
g39530 and n39779_not n39785_not ; n39786
g39531 and b[34]_not n39786_not ; n39787
g39532 and n39253_not n39725_not ; n39788
g39533 and n39263_not n39687 ; n39789
g39534 and n39683_not n39789 ; n39790
g39535 and n39684_not n39687_not ; n39791
g39536 and n39790_not n39791_not ; n39792
g39537 and n11619 n39792_not ; n39793
g39538 and n39724_not n39793 ; n39794
g39539 and n39788_not n39794_not ; n39795
g39540 and b[33]_not n39795_not ; n39796
g39541 and n39262_not n39725_not ; n39797
g39542 and n39272_not n39682 ; n39798
g39543 and n39678_not n39798 ; n39799
g39544 and n39679_not n39682_not ; n39800
g39545 and n39799_not n39800_not ; n39801
g39546 and n11619 n39801_not ; n39802
g39547 and n39724_not n39802 ; n39803
g39548 and n39797_not n39803_not ; n39804
g39549 and b[32]_not n39804_not ; n39805
g39550 and n39271_not n39725_not ; n39806
g39551 and n39281_not n39677 ; n39807
g39552 and n39673_not n39807 ; n39808
g39553 and n39674_not n39677_not ; n39809
g39554 and n39808_not n39809_not ; n39810
g39555 and n11619 n39810_not ; n39811
g39556 and n39724_not n39811 ; n39812
g39557 and n39806_not n39812_not ; n39813
g39558 and b[31]_not n39813_not ; n39814
g39559 and n39280_not n39725_not ; n39815
g39560 and n39290_not n39672 ; n39816
g39561 and n39668_not n39816 ; n39817
g39562 and n39669_not n39672_not ; n39818
g39563 and n39817_not n39818_not ; n39819
g39564 and n11619 n39819_not ; n39820
g39565 and n39724_not n39820 ; n39821
g39566 and n39815_not n39821_not ; n39822
g39567 and b[30]_not n39822_not ; n39823
g39568 and n39289_not n39725_not ; n39824
g39569 and n39299_not n39667 ; n39825
g39570 and n39663_not n39825 ; n39826
g39571 and n39664_not n39667_not ; n39827
g39572 and n39826_not n39827_not ; n39828
g39573 and n11619 n39828_not ; n39829
g39574 and n39724_not n39829 ; n39830
g39575 and n39824_not n39830_not ; n39831
g39576 and b[29]_not n39831_not ; n39832
g39577 and n39298_not n39725_not ; n39833
g39578 and n39308_not n39662 ; n39834
g39579 and n39658_not n39834 ; n39835
g39580 and n39659_not n39662_not ; n39836
g39581 and n39835_not n39836_not ; n39837
g39582 and n11619 n39837_not ; n39838
g39583 and n39724_not n39838 ; n39839
g39584 and n39833_not n39839_not ; n39840
g39585 and b[28]_not n39840_not ; n39841
g39586 and n39307_not n39725_not ; n39842
g39587 and n39317_not n39657 ; n39843
g39588 and n39653_not n39843 ; n39844
g39589 and n39654_not n39657_not ; n39845
g39590 and n39844_not n39845_not ; n39846
g39591 and n11619 n39846_not ; n39847
g39592 and n39724_not n39847 ; n39848
g39593 and n39842_not n39848_not ; n39849
g39594 and b[27]_not n39849_not ; n39850
g39595 and n39316_not n39725_not ; n39851
g39596 and n39326_not n39652 ; n39852
g39597 and n39648_not n39852 ; n39853
g39598 and n39649_not n39652_not ; n39854
g39599 and n39853_not n39854_not ; n39855
g39600 and n11619 n39855_not ; n39856
g39601 and n39724_not n39856 ; n39857
g39602 and n39851_not n39857_not ; n39858
g39603 and b[26]_not n39858_not ; n39859
g39604 and n39325_not n39725_not ; n39860
g39605 and n39335_not n39647 ; n39861
g39606 and n39643_not n39861 ; n39862
g39607 and n39644_not n39647_not ; n39863
g39608 and n39862_not n39863_not ; n39864
g39609 and n11619 n39864_not ; n39865
g39610 and n39724_not n39865 ; n39866
g39611 and n39860_not n39866_not ; n39867
g39612 and b[25]_not n39867_not ; n39868
g39613 and n39334_not n39725_not ; n39869
g39614 and n39344_not n39642 ; n39870
g39615 and n39638_not n39870 ; n39871
g39616 and n39639_not n39642_not ; n39872
g39617 and n39871_not n39872_not ; n39873
g39618 and n11619 n39873_not ; n39874
g39619 and n39724_not n39874 ; n39875
g39620 and n39869_not n39875_not ; n39876
g39621 and b[24]_not n39876_not ; n39877
g39622 and n39343_not n39725_not ; n39878
g39623 and n39353_not n39637 ; n39879
g39624 and n39633_not n39879 ; n39880
g39625 and n39634_not n39637_not ; n39881
g39626 and n39880_not n39881_not ; n39882
g39627 and n11619 n39882_not ; n39883
g39628 and n39724_not n39883 ; n39884
g39629 and n39878_not n39884_not ; n39885
g39630 and b[23]_not n39885_not ; n39886
g39631 and n39352_not n39725_not ; n39887
g39632 and n39362_not n39632 ; n39888
g39633 and n39628_not n39888 ; n39889
g39634 and n39629_not n39632_not ; n39890
g39635 and n39889_not n39890_not ; n39891
g39636 and n11619 n39891_not ; n39892
g39637 and n39724_not n39892 ; n39893
g39638 and n39887_not n39893_not ; n39894
g39639 and b[22]_not n39894_not ; n39895
g39640 and n39361_not n39725_not ; n39896
g39641 and n39371_not n39627 ; n39897
g39642 and n39623_not n39897 ; n39898
g39643 and n39624_not n39627_not ; n39899
g39644 and n39898_not n39899_not ; n39900
g39645 and n11619 n39900_not ; n39901
g39646 and n39724_not n39901 ; n39902
g39647 and n39896_not n39902_not ; n39903
g39648 and b[21]_not n39903_not ; n39904
g39649 and n39370_not n39725_not ; n39905
g39650 and n39380_not n39622 ; n39906
g39651 and n39618_not n39906 ; n39907
g39652 and n39619_not n39622_not ; n39908
g39653 and n39907_not n39908_not ; n39909
g39654 and n11619 n39909_not ; n39910
g39655 and n39724_not n39910 ; n39911
g39656 and n39905_not n39911_not ; n39912
g39657 and b[20]_not n39912_not ; n39913
g39658 and n39379_not n39725_not ; n39914
g39659 and n39389_not n39617 ; n39915
g39660 and n39613_not n39915 ; n39916
g39661 and n39614_not n39617_not ; n39917
g39662 and n39916_not n39917_not ; n39918
g39663 and n11619 n39918_not ; n39919
g39664 and n39724_not n39919 ; n39920
g39665 and n39914_not n39920_not ; n39921
g39666 and b[19]_not n39921_not ; n39922
g39667 and n39388_not n39725_not ; n39923
g39668 and n39398_not n39612 ; n39924
g39669 and n39608_not n39924 ; n39925
g39670 and n39609_not n39612_not ; n39926
g39671 and n39925_not n39926_not ; n39927
g39672 and n11619 n39927_not ; n39928
g39673 and n39724_not n39928 ; n39929
g39674 and n39923_not n39929_not ; n39930
g39675 and b[18]_not n39930_not ; n39931
g39676 and n39397_not n39725_not ; n39932
g39677 and n39407_not n39607 ; n39933
g39678 and n39603_not n39933 ; n39934
g39679 and n39604_not n39607_not ; n39935
g39680 and n39934_not n39935_not ; n39936
g39681 and n11619 n39936_not ; n39937
g39682 and n39724_not n39937 ; n39938
g39683 and n39932_not n39938_not ; n39939
g39684 and b[17]_not n39939_not ; n39940
g39685 and n39406_not n39725_not ; n39941
g39686 and n39416_not n39602 ; n39942
g39687 and n39598_not n39942 ; n39943
g39688 and n39599_not n39602_not ; n39944
g39689 and n39943_not n39944_not ; n39945
g39690 and n11619 n39945_not ; n39946
g39691 and n39724_not n39946 ; n39947
g39692 and n39941_not n39947_not ; n39948
g39693 and b[16]_not n39948_not ; n39949
g39694 and n39415_not n39725_not ; n39950
g39695 and n39425_not n39597 ; n39951
g39696 and n39593_not n39951 ; n39952
g39697 and n39594_not n39597_not ; n39953
g39698 and n39952_not n39953_not ; n39954
g39699 and n11619 n39954_not ; n39955
g39700 and n39724_not n39955 ; n39956
g39701 and n39950_not n39956_not ; n39957
g39702 and b[15]_not n39957_not ; n39958
g39703 and n39424_not n39725_not ; n39959
g39704 and n39434_not n39592 ; n39960
g39705 and n39588_not n39960 ; n39961
g39706 and n39589_not n39592_not ; n39962
g39707 and n39961_not n39962_not ; n39963
g39708 and n11619 n39963_not ; n39964
g39709 and n39724_not n39964 ; n39965
g39710 and n39959_not n39965_not ; n39966
g39711 and b[14]_not n39966_not ; n39967
g39712 and n39433_not n39725_not ; n39968
g39713 and n39443_not n39587 ; n39969
g39714 and n39583_not n39969 ; n39970
g39715 and n39584_not n39587_not ; n39971
g39716 and n39970_not n39971_not ; n39972
g39717 and n11619 n39972_not ; n39973
g39718 and n39724_not n39973 ; n39974
g39719 and n39968_not n39974_not ; n39975
g39720 and b[13]_not n39975_not ; n39976
g39721 and n39442_not n39725_not ; n39977
g39722 and n39452_not n39582 ; n39978
g39723 and n39578_not n39978 ; n39979
g39724 and n39579_not n39582_not ; n39980
g39725 and n39979_not n39980_not ; n39981
g39726 and n11619 n39981_not ; n39982
g39727 and n39724_not n39982 ; n39983
g39728 and n39977_not n39983_not ; n39984
g39729 and b[12]_not n39984_not ; n39985
g39730 and n39451_not n39725_not ; n39986
g39731 and n39461_not n39577 ; n39987
g39732 and n39573_not n39987 ; n39988
g39733 and n39574_not n39577_not ; n39989
g39734 and n39988_not n39989_not ; n39990
g39735 and n11619 n39990_not ; n39991
g39736 and n39724_not n39991 ; n39992
g39737 and n39986_not n39992_not ; n39993
g39738 and b[11]_not n39993_not ; n39994
g39739 and n39460_not n39725_not ; n39995
g39740 and n39470_not n39572 ; n39996
g39741 and n39568_not n39996 ; n39997
g39742 and n39569_not n39572_not ; n39998
g39743 and n39997_not n39998_not ; n39999
g39744 and n11619 n39999_not ; n40000
g39745 and n39724_not n40000 ; n40001
g39746 and n39995_not n40001_not ; n40002
g39747 and b[10]_not n40002_not ; n40003
g39748 and n39469_not n39725_not ; n40004
g39749 and n39479_not n39567 ; n40005
g39750 and n39563_not n40005 ; n40006
g39751 and n39564_not n39567_not ; n40007
g39752 and n40006_not n40007_not ; n40008
g39753 and n11619 n40008_not ; n40009
g39754 and n39724_not n40009 ; n40010
g39755 and n40004_not n40010_not ; n40011
g39756 and b[9]_not n40011_not ; n40012
g39757 and n39478_not n39725_not ; n40013
g39758 and n39488_not n39562 ; n40014
g39759 and n39558_not n40014 ; n40015
g39760 and n39559_not n39562_not ; n40016
g39761 and n40015_not n40016_not ; n40017
g39762 and n11619 n40017_not ; n40018
g39763 and n39724_not n40018 ; n40019
g39764 and n40013_not n40019_not ; n40020
g39765 and b[8]_not n40020_not ; n40021
g39766 and n39487_not n39725_not ; n40022
g39767 and n39497_not n39557 ; n40023
g39768 and n39553_not n40023 ; n40024
g39769 and n39554_not n39557_not ; n40025
g39770 and n40024_not n40025_not ; n40026
g39771 and n11619 n40026_not ; n40027
g39772 and n39724_not n40027 ; n40028
g39773 and n40022_not n40028_not ; n40029
g39774 and b[7]_not n40029_not ; n40030
g39775 and n39496_not n39725_not ; n40031
g39776 and n39506_not n39552 ; n40032
g39777 and n39548_not n40032 ; n40033
g39778 and n39549_not n39552_not ; n40034
g39779 and n40033_not n40034_not ; n40035
g39780 and n11619 n40035_not ; n40036
g39781 and n39724_not n40036 ; n40037
g39782 and n40031_not n40037_not ; n40038
g39783 and b[6]_not n40038_not ; n40039
g39784 and n39505_not n39725_not ; n40040
g39785 and n39515_not n39547 ; n40041
g39786 and n39543_not n40041 ; n40042
g39787 and n39544_not n39547_not ; n40043
g39788 and n40042_not n40043_not ; n40044
g39789 and n11619 n40044_not ; n40045
g39790 and n39724_not n40045 ; n40046
g39791 and n40040_not n40046_not ; n40047
g39792 and b[5]_not n40047_not ; n40048
g39793 and n39514_not n39725_not ; n40049
g39794 and n39523_not n39542 ; n40050
g39795 and n39538_not n40050 ; n40051
g39796 and n39539_not n39542_not ; n40052
g39797 and n40051_not n40052_not ; n40053
g39798 and n11619 n40053_not ; n40054
g39799 and n39724_not n40054 ; n40055
g39800 and n40049_not n40055_not ; n40056
g39801 and b[4]_not n40056_not ; n40057
g39802 and n39522_not n39725_not ; n40058
g39803 and n39533_not n39537 ; n40059
g39804 and n39532_not n40059 ; n40060
g39805 and n39534_not n39537_not ; n40061
g39806 and n40060_not n40061_not ; n40062
g39807 and n11619 n40062_not ; n40063
g39808 and n39724_not n40063 ; n40064
g39809 and n40058_not n40064_not ; n40065
g39810 and b[3]_not n40065_not ; n40066
g39811 and n39527_not n39725_not ; n40067
g39812 and n11425 n39530_not ; n40068
g39813 and n39528_not n40068 ; n40069
g39814 and n11619 n40069_not ; n40070
g39815 and n39532_not n40070 ; n40071
g39816 and n39724_not n40071 ; n40072
g39817 and n40067_not n40072_not ; n40073
g39818 and b[2]_not n40073_not ; n40074
g39819 and n11973 n39724_not ; n40075
g39820 and a[24] n40075_not ; n40076
g39821 and n11978 n39724_not ; n40077
g39822 and n40076_not n40077_not ; n40078
g39823 and b[1] n40078_not ; n40079
g39824 and b[1]_not n40077_not ; n40080
g39825 and n40076_not n40080 ; n40081
g39826 and n40079_not n40081_not ; n40082
g39827 and n11985_not n40082_not ; n40083
g39828 and b[1]_not n40078_not ; n40084
g39829 and n40083_not n40084_not ; n40085
g39830 and b[2] n40072_not ; n40086
g39831 and n40067_not n40086 ; n40087
g39832 and n40074_not n40087_not ; n40088
g39833 and n40085_not n40088 ; n40089
g39834 and n40074_not n40089_not ; n40090
g39835 and b[3] n40064_not ; n40091
g39836 and n40058_not n40091 ; n40092
g39837 and n40066_not n40092_not ; n40093
g39838 and n40090_not n40093 ; n40094
g39839 and n40066_not n40094_not ; n40095
g39840 and b[4] n40055_not ; n40096
g39841 and n40049_not n40096 ; n40097
g39842 and n40057_not n40097_not ; n40098
g39843 and n40095_not n40098 ; n40099
g39844 and n40057_not n40099_not ; n40100
g39845 and b[5] n40046_not ; n40101
g39846 and n40040_not n40101 ; n40102
g39847 and n40048_not n40102_not ; n40103
g39848 and n40100_not n40103 ; n40104
g39849 and n40048_not n40104_not ; n40105
g39850 and b[6] n40037_not ; n40106
g39851 and n40031_not n40106 ; n40107
g39852 and n40039_not n40107_not ; n40108
g39853 and n40105_not n40108 ; n40109
g39854 and n40039_not n40109_not ; n40110
g39855 and b[7] n40028_not ; n40111
g39856 and n40022_not n40111 ; n40112
g39857 and n40030_not n40112_not ; n40113
g39858 and n40110_not n40113 ; n40114
g39859 and n40030_not n40114_not ; n40115
g39860 and b[8] n40019_not ; n40116
g39861 and n40013_not n40116 ; n40117
g39862 and n40021_not n40117_not ; n40118
g39863 and n40115_not n40118 ; n40119
g39864 and n40021_not n40119_not ; n40120
g39865 and b[9] n40010_not ; n40121
g39866 and n40004_not n40121 ; n40122
g39867 and n40012_not n40122_not ; n40123
g39868 and n40120_not n40123 ; n40124
g39869 and n40012_not n40124_not ; n40125
g39870 and b[10] n40001_not ; n40126
g39871 and n39995_not n40126 ; n40127
g39872 and n40003_not n40127_not ; n40128
g39873 and n40125_not n40128 ; n40129
g39874 and n40003_not n40129_not ; n40130
g39875 and b[11] n39992_not ; n40131
g39876 and n39986_not n40131 ; n40132
g39877 and n39994_not n40132_not ; n40133
g39878 and n40130_not n40133 ; n40134
g39879 and n39994_not n40134_not ; n40135
g39880 and b[12] n39983_not ; n40136
g39881 and n39977_not n40136 ; n40137
g39882 and n39985_not n40137_not ; n40138
g39883 and n40135_not n40138 ; n40139
g39884 and n39985_not n40139_not ; n40140
g39885 and b[13] n39974_not ; n40141
g39886 and n39968_not n40141 ; n40142
g39887 and n39976_not n40142_not ; n40143
g39888 and n40140_not n40143 ; n40144
g39889 and n39976_not n40144_not ; n40145
g39890 and b[14] n39965_not ; n40146
g39891 and n39959_not n40146 ; n40147
g39892 and n39967_not n40147_not ; n40148
g39893 and n40145_not n40148 ; n40149
g39894 and n39967_not n40149_not ; n40150
g39895 and b[15] n39956_not ; n40151
g39896 and n39950_not n40151 ; n40152
g39897 and n39958_not n40152_not ; n40153
g39898 and n40150_not n40153 ; n40154
g39899 and n39958_not n40154_not ; n40155
g39900 and b[16] n39947_not ; n40156
g39901 and n39941_not n40156 ; n40157
g39902 and n39949_not n40157_not ; n40158
g39903 and n40155_not n40158 ; n40159
g39904 and n39949_not n40159_not ; n40160
g39905 and b[17] n39938_not ; n40161
g39906 and n39932_not n40161 ; n40162
g39907 and n39940_not n40162_not ; n40163
g39908 and n40160_not n40163 ; n40164
g39909 and n39940_not n40164_not ; n40165
g39910 and b[18] n39929_not ; n40166
g39911 and n39923_not n40166 ; n40167
g39912 and n39931_not n40167_not ; n40168
g39913 and n40165_not n40168 ; n40169
g39914 and n39931_not n40169_not ; n40170
g39915 and b[19] n39920_not ; n40171
g39916 and n39914_not n40171 ; n40172
g39917 and n39922_not n40172_not ; n40173
g39918 and n40170_not n40173 ; n40174
g39919 and n39922_not n40174_not ; n40175
g39920 and b[20] n39911_not ; n40176
g39921 and n39905_not n40176 ; n40177
g39922 and n39913_not n40177_not ; n40178
g39923 and n40175_not n40178 ; n40179
g39924 and n39913_not n40179_not ; n40180
g39925 and b[21] n39902_not ; n40181
g39926 and n39896_not n40181 ; n40182
g39927 and n39904_not n40182_not ; n40183
g39928 and n40180_not n40183 ; n40184
g39929 and n39904_not n40184_not ; n40185
g39930 and b[22] n39893_not ; n40186
g39931 and n39887_not n40186 ; n40187
g39932 and n39895_not n40187_not ; n40188
g39933 and n40185_not n40188 ; n40189
g39934 and n39895_not n40189_not ; n40190
g39935 and b[23] n39884_not ; n40191
g39936 and n39878_not n40191 ; n40192
g39937 and n39886_not n40192_not ; n40193
g39938 and n40190_not n40193 ; n40194
g39939 and n39886_not n40194_not ; n40195
g39940 and b[24] n39875_not ; n40196
g39941 and n39869_not n40196 ; n40197
g39942 and n39877_not n40197_not ; n40198
g39943 and n40195_not n40198 ; n40199
g39944 and n39877_not n40199_not ; n40200
g39945 and b[25] n39866_not ; n40201
g39946 and n39860_not n40201 ; n40202
g39947 and n39868_not n40202_not ; n40203
g39948 and n40200_not n40203 ; n40204
g39949 and n39868_not n40204_not ; n40205
g39950 and b[26] n39857_not ; n40206
g39951 and n39851_not n40206 ; n40207
g39952 and n39859_not n40207_not ; n40208
g39953 and n40205_not n40208 ; n40209
g39954 and n39859_not n40209_not ; n40210
g39955 and b[27] n39848_not ; n40211
g39956 and n39842_not n40211 ; n40212
g39957 and n39850_not n40212_not ; n40213
g39958 and n40210_not n40213 ; n40214
g39959 and n39850_not n40214_not ; n40215
g39960 and b[28] n39839_not ; n40216
g39961 and n39833_not n40216 ; n40217
g39962 and n39841_not n40217_not ; n40218
g39963 and n40215_not n40218 ; n40219
g39964 and n39841_not n40219_not ; n40220
g39965 and b[29] n39830_not ; n40221
g39966 and n39824_not n40221 ; n40222
g39967 and n39832_not n40222_not ; n40223
g39968 and n40220_not n40223 ; n40224
g39969 and n39832_not n40224_not ; n40225
g39970 and b[30] n39821_not ; n40226
g39971 and n39815_not n40226 ; n40227
g39972 and n39823_not n40227_not ; n40228
g39973 and n40225_not n40228 ; n40229
g39974 and n39823_not n40229_not ; n40230
g39975 and b[31] n39812_not ; n40231
g39976 and n39806_not n40231 ; n40232
g39977 and n39814_not n40232_not ; n40233
g39978 and n40230_not n40233 ; n40234
g39979 and n39814_not n40234_not ; n40235
g39980 and b[32] n39803_not ; n40236
g39981 and n39797_not n40236 ; n40237
g39982 and n39805_not n40237_not ; n40238
g39983 and n40235_not n40238 ; n40239
g39984 and n39805_not n40239_not ; n40240
g39985 and b[33] n39794_not ; n40241
g39986 and n39788_not n40241 ; n40242
g39987 and n39796_not n40242_not ; n40243
g39988 and n40240_not n40243 ; n40244
g39989 and n39796_not n40244_not ; n40245
g39990 and b[34] n39785_not ; n40246
g39991 and n39779_not n40246 ; n40247
g39992 and n39787_not n40247_not ; n40248
g39993 and n40245_not n40248 ; n40249
g39994 and n39787_not n40249_not ; n40250
g39995 and b[35] n39776_not ; n40251
g39996 and n39770_not n40251 ; n40252
g39997 and n39778_not n40252_not ; n40253
g39998 and n40250_not n40253 ; n40254
g39999 and n39778_not n40254_not ; n40255
g40000 and b[36] n39767_not ; n40256
g40001 and n39761_not n40256 ; n40257
g40002 and n39769_not n40257_not ; n40258
g40003 and n40255_not n40258 ; n40259
g40004 and n39769_not n40259_not ; n40260
g40005 and b[37] n39758_not ; n40261
g40006 and n39752_not n40261 ; n40262
g40007 and n39760_not n40262_not ; n40263
g40008 and n40260_not n40263 ; n40264
g40009 and n39760_not n40264_not ; n40265
g40010 and b[38] n39749_not ; n40266
g40011 and n39743_not n40266 ; n40267
g40012 and n39751_not n40267_not ; n40268
g40013 and n40265_not n40268 ; n40269
g40014 and n39751_not n40269_not ; n40270
g40015 and b[39] n39732_not ; n40271
g40016 and n39726_not n40271 ; n40272
g40017 and n39742_not n40272_not ; n40273
g40018 and n40270_not n40273 ; n40274
g40019 and n39742_not n40274_not ; n40275
g40020 and b[40] n39734_not ; n40276
g40021 and n39739_not n40276 ; n40277
g40022 and n39741_not n40277_not ; n40278
g40023 and n40275_not n40278 ; n40279
g40024 and n39741_not n40279_not ; n40280
g40025 and n12184 n40280_not ; n40281
g40026 and n39733_not n40281_not ; n40282
g40027 and n39751_not n40273 ; n40283
g40028 and n40269_not n40283 ; n40284
g40029 and n40270_not n40273_not ; n40285
g40030 and n40284_not n40285_not ; n40286
g40031 and n12184 n40286_not ; n40287
g40032 and n40280_not n40287 ; n40288
g40033 and n40282_not n40288_not ; n40289
g40034 and b[40]_not n40289_not ; n40290
g40035 and n39750_not n40281_not ; n40291
g40036 and n39760_not n40268 ; n40292
g40037 and n40264_not n40292 ; n40293
g40038 and n40265_not n40268_not ; n40294
g40039 and n40293_not n40294_not ; n40295
g40040 and n12184 n40295_not ; n40296
g40041 and n40280_not n40296 ; n40297
g40042 and n40291_not n40297_not ; n40298
g40043 and b[39]_not n40298_not ; n40299
g40044 and n39759_not n40281_not ; n40300
g40045 and n39769_not n40263 ; n40301
g40046 and n40259_not n40301 ; n40302
g40047 and n40260_not n40263_not ; n40303
g40048 and n40302_not n40303_not ; n40304
g40049 and n12184 n40304_not ; n40305
g40050 and n40280_not n40305 ; n40306
g40051 and n40300_not n40306_not ; n40307
g40052 and b[38]_not n40307_not ; n40308
g40053 and n39768_not n40281_not ; n40309
g40054 and n39778_not n40258 ; n40310
g40055 and n40254_not n40310 ; n40311
g40056 and n40255_not n40258_not ; n40312
g40057 and n40311_not n40312_not ; n40313
g40058 and n12184 n40313_not ; n40314
g40059 and n40280_not n40314 ; n40315
g40060 and n40309_not n40315_not ; n40316
g40061 and b[37]_not n40316_not ; n40317
g40062 and n39777_not n40281_not ; n40318
g40063 and n39787_not n40253 ; n40319
g40064 and n40249_not n40319 ; n40320
g40065 and n40250_not n40253_not ; n40321
g40066 and n40320_not n40321_not ; n40322
g40067 and n12184 n40322_not ; n40323
g40068 and n40280_not n40323 ; n40324
g40069 and n40318_not n40324_not ; n40325
g40070 and b[36]_not n40325_not ; n40326
g40071 and n39786_not n40281_not ; n40327
g40072 and n39796_not n40248 ; n40328
g40073 and n40244_not n40328 ; n40329
g40074 and n40245_not n40248_not ; n40330
g40075 and n40329_not n40330_not ; n40331
g40076 and n12184 n40331_not ; n40332
g40077 and n40280_not n40332 ; n40333
g40078 and n40327_not n40333_not ; n40334
g40079 and b[35]_not n40334_not ; n40335
g40080 and n39795_not n40281_not ; n40336
g40081 and n39805_not n40243 ; n40337
g40082 and n40239_not n40337 ; n40338
g40083 and n40240_not n40243_not ; n40339
g40084 and n40338_not n40339_not ; n40340
g40085 and n12184 n40340_not ; n40341
g40086 and n40280_not n40341 ; n40342
g40087 and n40336_not n40342_not ; n40343
g40088 and b[34]_not n40343_not ; n40344
g40089 and n39804_not n40281_not ; n40345
g40090 and n39814_not n40238 ; n40346
g40091 and n40234_not n40346 ; n40347
g40092 and n40235_not n40238_not ; n40348
g40093 and n40347_not n40348_not ; n40349
g40094 and n12184 n40349_not ; n40350
g40095 and n40280_not n40350 ; n40351
g40096 and n40345_not n40351_not ; n40352
g40097 and b[33]_not n40352_not ; n40353
g40098 and n39813_not n40281_not ; n40354
g40099 and n39823_not n40233 ; n40355
g40100 and n40229_not n40355 ; n40356
g40101 and n40230_not n40233_not ; n40357
g40102 and n40356_not n40357_not ; n40358
g40103 and n12184 n40358_not ; n40359
g40104 and n40280_not n40359 ; n40360
g40105 and n40354_not n40360_not ; n40361
g40106 and b[32]_not n40361_not ; n40362
g40107 and n39822_not n40281_not ; n40363
g40108 and n39832_not n40228 ; n40364
g40109 and n40224_not n40364 ; n40365
g40110 and n40225_not n40228_not ; n40366
g40111 and n40365_not n40366_not ; n40367
g40112 and n12184 n40367_not ; n40368
g40113 and n40280_not n40368 ; n40369
g40114 and n40363_not n40369_not ; n40370
g40115 and b[31]_not n40370_not ; n40371
g40116 and n39831_not n40281_not ; n40372
g40117 and n39841_not n40223 ; n40373
g40118 and n40219_not n40373 ; n40374
g40119 and n40220_not n40223_not ; n40375
g40120 and n40374_not n40375_not ; n40376
g40121 and n12184 n40376_not ; n40377
g40122 and n40280_not n40377 ; n40378
g40123 and n40372_not n40378_not ; n40379
g40124 and b[30]_not n40379_not ; n40380
g40125 and n39840_not n40281_not ; n40381
g40126 and n39850_not n40218 ; n40382
g40127 and n40214_not n40382 ; n40383
g40128 and n40215_not n40218_not ; n40384
g40129 and n40383_not n40384_not ; n40385
g40130 and n12184 n40385_not ; n40386
g40131 and n40280_not n40386 ; n40387
g40132 and n40381_not n40387_not ; n40388
g40133 and b[29]_not n40388_not ; n40389
g40134 and n39849_not n40281_not ; n40390
g40135 and n39859_not n40213 ; n40391
g40136 and n40209_not n40391 ; n40392
g40137 and n40210_not n40213_not ; n40393
g40138 and n40392_not n40393_not ; n40394
g40139 and n12184 n40394_not ; n40395
g40140 and n40280_not n40395 ; n40396
g40141 and n40390_not n40396_not ; n40397
g40142 and b[28]_not n40397_not ; n40398
g40143 and n39858_not n40281_not ; n40399
g40144 and n39868_not n40208 ; n40400
g40145 and n40204_not n40400 ; n40401
g40146 and n40205_not n40208_not ; n40402
g40147 and n40401_not n40402_not ; n40403
g40148 and n12184 n40403_not ; n40404
g40149 and n40280_not n40404 ; n40405
g40150 and n40399_not n40405_not ; n40406
g40151 and b[27]_not n40406_not ; n40407
g40152 and n39867_not n40281_not ; n40408
g40153 and n39877_not n40203 ; n40409
g40154 and n40199_not n40409 ; n40410
g40155 and n40200_not n40203_not ; n40411
g40156 and n40410_not n40411_not ; n40412
g40157 and n12184 n40412_not ; n40413
g40158 and n40280_not n40413 ; n40414
g40159 and n40408_not n40414_not ; n40415
g40160 and b[26]_not n40415_not ; n40416
g40161 and n39876_not n40281_not ; n40417
g40162 and n39886_not n40198 ; n40418
g40163 and n40194_not n40418 ; n40419
g40164 and n40195_not n40198_not ; n40420
g40165 and n40419_not n40420_not ; n40421
g40166 and n12184 n40421_not ; n40422
g40167 and n40280_not n40422 ; n40423
g40168 and n40417_not n40423_not ; n40424
g40169 and b[25]_not n40424_not ; n40425
g40170 and n39885_not n40281_not ; n40426
g40171 and n39895_not n40193 ; n40427
g40172 and n40189_not n40427 ; n40428
g40173 and n40190_not n40193_not ; n40429
g40174 and n40428_not n40429_not ; n40430
g40175 and n12184 n40430_not ; n40431
g40176 and n40280_not n40431 ; n40432
g40177 and n40426_not n40432_not ; n40433
g40178 and b[24]_not n40433_not ; n40434
g40179 and n39894_not n40281_not ; n40435
g40180 and n39904_not n40188 ; n40436
g40181 and n40184_not n40436 ; n40437
g40182 and n40185_not n40188_not ; n40438
g40183 and n40437_not n40438_not ; n40439
g40184 and n12184 n40439_not ; n40440
g40185 and n40280_not n40440 ; n40441
g40186 and n40435_not n40441_not ; n40442
g40187 and b[23]_not n40442_not ; n40443
g40188 and n39903_not n40281_not ; n40444
g40189 and n39913_not n40183 ; n40445
g40190 and n40179_not n40445 ; n40446
g40191 and n40180_not n40183_not ; n40447
g40192 and n40446_not n40447_not ; n40448
g40193 and n12184 n40448_not ; n40449
g40194 and n40280_not n40449 ; n40450
g40195 and n40444_not n40450_not ; n40451
g40196 and b[22]_not n40451_not ; n40452
g40197 and n39912_not n40281_not ; n40453
g40198 and n39922_not n40178 ; n40454
g40199 and n40174_not n40454 ; n40455
g40200 and n40175_not n40178_not ; n40456
g40201 and n40455_not n40456_not ; n40457
g40202 and n12184 n40457_not ; n40458
g40203 and n40280_not n40458 ; n40459
g40204 and n40453_not n40459_not ; n40460
g40205 and b[21]_not n40460_not ; n40461
g40206 and n39921_not n40281_not ; n40462
g40207 and n39931_not n40173 ; n40463
g40208 and n40169_not n40463 ; n40464
g40209 and n40170_not n40173_not ; n40465
g40210 and n40464_not n40465_not ; n40466
g40211 and n12184 n40466_not ; n40467
g40212 and n40280_not n40467 ; n40468
g40213 and n40462_not n40468_not ; n40469
g40214 and b[20]_not n40469_not ; n40470
g40215 and n39930_not n40281_not ; n40471
g40216 and n39940_not n40168 ; n40472
g40217 and n40164_not n40472 ; n40473
g40218 and n40165_not n40168_not ; n40474
g40219 and n40473_not n40474_not ; n40475
g40220 and n12184 n40475_not ; n40476
g40221 and n40280_not n40476 ; n40477
g40222 and n40471_not n40477_not ; n40478
g40223 and b[19]_not n40478_not ; n40479
g40224 and n39939_not n40281_not ; n40480
g40225 and n39949_not n40163 ; n40481
g40226 and n40159_not n40481 ; n40482
g40227 and n40160_not n40163_not ; n40483
g40228 and n40482_not n40483_not ; n40484
g40229 and n12184 n40484_not ; n40485
g40230 and n40280_not n40485 ; n40486
g40231 and n40480_not n40486_not ; n40487
g40232 and b[18]_not n40487_not ; n40488
g40233 and n39948_not n40281_not ; n40489
g40234 and n39958_not n40158 ; n40490
g40235 and n40154_not n40490 ; n40491
g40236 and n40155_not n40158_not ; n40492
g40237 and n40491_not n40492_not ; n40493
g40238 and n12184 n40493_not ; n40494
g40239 and n40280_not n40494 ; n40495
g40240 and n40489_not n40495_not ; n40496
g40241 and b[17]_not n40496_not ; n40497
g40242 and n39957_not n40281_not ; n40498
g40243 and n39967_not n40153 ; n40499
g40244 and n40149_not n40499 ; n40500
g40245 and n40150_not n40153_not ; n40501
g40246 and n40500_not n40501_not ; n40502
g40247 and n12184 n40502_not ; n40503
g40248 and n40280_not n40503 ; n40504
g40249 and n40498_not n40504_not ; n40505
g40250 and b[16]_not n40505_not ; n40506
g40251 and n39966_not n40281_not ; n40507
g40252 and n39976_not n40148 ; n40508
g40253 and n40144_not n40508 ; n40509
g40254 and n40145_not n40148_not ; n40510
g40255 and n40509_not n40510_not ; n40511
g40256 and n12184 n40511_not ; n40512
g40257 and n40280_not n40512 ; n40513
g40258 and n40507_not n40513_not ; n40514
g40259 and b[15]_not n40514_not ; n40515
g40260 and n39975_not n40281_not ; n40516
g40261 and n39985_not n40143 ; n40517
g40262 and n40139_not n40517 ; n40518
g40263 and n40140_not n40143_not ; n40519
g40264 and n40518_not n40519_not ; n40520
g40265 and n12184 n40520_not ; n40521
g40266 and n40280_not n40521 ; n40522
g40267 and n40516_not n40522_not ; n40523
g40268 and b[14]_not n40523_not ; n40524
g40269 and n39984_not n40281_not ; n40525
g40270 and n39994_not n40138 ; n40526
g40271 and n40134_not n40526 ; n40527
g40272 and n40135_not n40138_not ; n40528
g40273 and n40527_not n40528_not ; n40529
g40274 and n12184 n40529_not ; n40530
g40275 and n40280_not n40530 ; n40531
g40276 and n40525_not n40531_not ; n40532
g40277 and b[13]_not n40532_not ; n40533
g40278 and n39993_not n40281_not ; n40534
g40279 and n40003_not n40133 ; n40535
g40280 and n40129_not n40535 ; n40536
g40281 and n40130_not n40133_not ; n40537
g40282 and n40536_not n40537_not ; n40538
g40283 and n12184 n40538_not ; n40539
g40284 and n40280_not n40539 ; n40540
g40285 and n40534_not n40540_not ; n40541
g40286 and b[12]_not n40541_not ; n40542
g40287 and n40002_not n40281_not ; n40543
g40288 and n40012_not n40128 ; n40544
g40289 and n40124_not n40544 ; n40545
g40290 and n40125_not n40128_not ; n40546
g40291 and n40545_not n40546_not ; n40547
g40292 and n12184 n40547_not ; n40548
g40293 and n40280_not n40548 ; n40549
g40294 and n40543_not n40549_not ; n40550
g40295 and b[11]_not n40550_not ; n40551
g40296 and n40011_not n40281_not ; n40552
g40297 and n40021_not n40123 ; n40553
g40298 and n40119_not n40553 ; n40554
g40299 and n40120_not n40123_not ; n40555
g40300 and n40554_not n40555_not ; n40556
g40301 and n12184 n40556_not ; n40557
g40302 and n40280_not n40557 ; n40558
g40303 and n40552_not n40558_not ; n40559
g40304 and b[10]_not n40559_not ; n40560
g40305 and n40020_not n40281_not ; n40561
g40306 and n40030_not n40118 ; n40562
g40307 and n40114_not n40562 ; n40563
g40308 and n40115_not n40118_not ; n40564
g40309 and n40563_not n40564_not ; n40565
g40310 and n12184 n40565_not ; n40566
g40311 and n40280_not n40566 ; n40567
g40312 and n40561_not n40567_not ; n40568
g40313 and b[9]_not n40568_not ; n40569
g40314 and n40029_not n40281_not ; n40570
g40315 and n40039_not n40113 ; n40571
g40316 and n40109_not n40571 ; n40572
g40317 and n40110_not n40113_not ; n40573
g40318 and n40572_not n40573_not ; n40574
g40319 and n12184 n40574_not ; n40575
g40320 and n40280_not n40575 ; n40576
g40321 and n40570_not n40576_not ; n40577
g40322 and b[8]_not n40577_not ; n40578
g40323 and n40038_not n40281_not ; n40579
g40324 and n40048_not n40108 ; n40580
g40325 and n40104_not n40580 ; n40581
g40326 and n40105_not n40108_not ; n40582
g40327 and n40581_not n40582_not ; n40583
g40328 and n12184 n40583_not ; n40584
g40329 and n40280_not n40584 ; n40585
g40330 and n40579_not n40585_not ; n40586
g40331 and b[7]_not n40586_not ; n40587
g40332 and n40047_not n40281_not ; n40588
g40333 and n40057_not n40103 ; n40589
g40334 and n40099_not n40589 ; n40590
g40335 and n40100_not n40103_not ; n40591
g40336 and n40590_not n40591_not ; n40592
g40337 and n12184 n40592_not ; n40593
g40338 and n40280_not n40593 ; n40594
g40339 and n40588_not n40594_not ; n40595
g40340 and b[6]_not n40595_not ; n40596
g40341 and n40056_not n40281_not ; n40597
g40342 and n40066_not n40098 ; n40598
g40343 and n40094_not n40598 ; n40599
g40344 and n40095_not n40098_not ; n40600
g40345 and n40599_not n40600_not ; n40601
g40346 and n12184 n40601_not ; n40602
g40347 and n40280_not n40602 ; n40603
g40348 and n40597_not n40603_not ; n40604
g40349 and b[5]_not n40604_not ; n40605
g40350 and n40065_not n40281_not ; n40606
g40351 and n40074_not n40093 ; n40607
g40352 and n40089_not n40607 ; n40608
g40353 and n40090_not n40093_not ; n40609
g40354 and n40608_not n40609_not ; n40610
g40355 and n12184 n40610_not ; n40611
g40356 and n40280_not n40611 ; n40612
g40357 and n40606_not n40612_not ; n40613
g40358 and b[4]_not n40613_not ; n40614
g40359 and n40073_not n40281_not ; n40615
g40360 and n40084_not n40088 ; n40616
g40361 and n40083_not n40616 ; n40617
g40362 and n40085_not n40088_not ; n40618
g40363 and n40617_not n40618_not ; n40619
g40364 and n12184 n40619_not ; n40620
g40365 and n40280_not n40620 ; n40621
g40366 and n40615_not n40621_not ; n40622
g40367 and b[3]_not n40622_not ; n40623
g40368 and n40078_not n40281_not ; n40624
g40369 and n11985 n40081_not ; n40625
g40370 and n40079_not n40625 ; n40626
g40371 and n12184 n40626_not ; n40627
g40372 and n40083_not n40627 ; n40628
g40373 and n40280_not n40628 ; n40629
g40374 and n40624_not n40629_not ; n40630
g40375 and b[2]_not n40630_not ; n40631
g40376 and n12539 n40280_not ; n40632
g40377 and a[23] n40632_not ; n40633
g40378 and n12544 n40280_not ; n40634
g40379 and n40633_not n40634_not ; n40635
g40380 and b[1] n40635_not ; n40636
g40381 and b[1]_not n40634_not ; n40637
g40382 and n40633_not n40637 ; n40638
g40383 and n40636_not n40638_not ; n40639
g40384 and n12551_not n40639_not ; n40640
g40385 and b[1]_not n40635_not ; n40641
g40386 and n40640_not n40641_not ; n40642
g40387 and b[2] n40629_not ; n40643
g40388 and n40624_not n40643 ; n40644
g40389 and n40631_not n40644_not ; n40645
g40390 and n40642_not n40645 ; n40646
g40391 and n40631_not n40646_not ; n40647
g40392 and b[3] n40621_not ; n40648
g40393 and n40615_not n40648 ; n40649
g40394 and n40623_not n40649_not ; n40650
g40395 and n40647_not n40650 ; n40651
g40396 and n40623_not n40651_not ; n40652
g40397 and b[4] n40612_not ; n40653
g40398 and n40606_not n40653 ; n40654
g40399 and n40614_not n40654_not ; n40655
g40400 and n40652_not n40655 ; n40656
g40401 and n40614_not n40656_not ; n40657
g40402 and b[5] n40603_not ; n40658
g40403 and n40597_not n40658 ; n40659
g40404 and n40605_not n40659_not ; n40660
g40405 and n40657_not n40660 ; n40661
g40406 and n40605_not n40661_not ; n40662
g40407 and b[6] n40594_not ; n40663
g40408 and n40588_not n40663 ; n40664
g40409 and n40596_not n40664_not ; n40665
g40410 and n40662_not n40665 ; n40666
g40411 and n40596_not n40666_not ; n40667
g40412 and b[7] n40585_not ; n40668
g40413 and n40579_not n40668 ; n40669
g40414 and n40587_not n40669_not ; n40670
g40415 and n40667_not n40670 ; n40671
g40416 and n40587_not n40671_not ; n40672
g40417 and b[8] n40576_not ; n40673
g40418 and n40570_not n40673 ; n40674
g40419 and n40578_not n40674_not ; n40675
g40420 and n40672_not n40675 ; n40676
g40421 and n40578_not n40676_not ; n40677
g40422 and b[9] n40567_not ; n40678
g40423 and n40561_not n40678 ; n40679
g40424 and n40569_not n40679_not ; n40680
g40425 and n40677_not n40680 ; n40681
g40426 and n40569_not n40681_not ; n40682
g40427 and b[10] n40558_not ; n40683
g40428 and n40552_not n40683 ; n40684
g40429 and n40560_not n40684_not ; n40685
g40430 and n40682_not n40685 ; n40686
g40431 and n40560_not n40686_not ; n40687
g40432 and b[11] n40549_not ; n40688
g40433 and n40543_not n40688 ; n40689
g40434 and n40551_not n40689_not ; n40690
g40435 and n40687_not n40690 ; n40691
g40436 and n40551_not n40691_not ; n40692
g40437 and b[12] n40540_not ; n40693
g40438 and n40534_not n40693 ; n40694
g40439 and n40542_not n40694_not ; n40695
g40440 and n40692_not n40695 ; n40696
g40441 and n40542_not n40696_not ; n40697
g40442 and b[13] n40531_not ; n40698
g40443 and n40525_not n40698 ; n40699
g40444 and n40533_not n40699_not ; n40700
g40445 and n40697_not n40700 ; n40701
g40446 and n40533_not n40701_not ; n40702
g40447 and b[14] n40522_not ; n40703
g40448 and n40516_not n40703 ; n40704
g40449 and n40524_not n40704_not ; n40705
g40450 and n40702_not n40705 ; n40706
g40451 and n40524_not n40706_not ; n40707
g40452 and b[15] n40513_not ; n40708
g40453 and n40507_not n40708 ; n40709
g40454 and n40515_not n40709_not ; n40710
g40455 and n40707_not n40710 ; n40711
g40456 and n40515_not n40711_not ; n40712
g40457 and b[16] n40504_not ; n40713
g40458 and n40498_not n40713 ; n40714
g40459 and n40506_not n40714_not ; n40715
g40460 and n40712_not n40715 ; n40716
g40461 and n40506_not n40716_not ; n40717
g40462 and b[17] n40495_not ; n40718
g40463 and n40489_not n40718 ; n40719
g40464 and n40497_not n40719_not ; n40720
g40465 and n40717_not n40720 ; n40721
g40466 and n40497_not n40721_not ; n40722
g40467 and b[18] n40486_not ; n40723
g40468 and n40480_not n40723 ; n40724
g40469 and n40488_not n40724_not ; n40725
g40470 and n40722_not n40725 ; n40726
g40471 and n40488_not n40726_not ; n40727
g40472 and b[19] n40477_not ; n40728
g40473 and n40471_not n40728 ; n40729
g40474 and n40479_not n40729_not ; n40730
g40475 and n40727_not n40730 ; n40731
g40476 and n40479_not n40731_not ; n40732
g40477 and b[20] n40468_not ; n40733
g40478 and n40462_not n40733 ; n40734
g40479 and n40470_not n40734_not ; n40735
g40480 and n40732_not n40735 ; n40736
g40481 and n40470_not n40736_not ; n40737
g40482 and b[21] n40459_not ; n40738
g40483 and n40453_not n40738 ; n40739
g40484 and n40461_not n40739_not ; n40740
g40485 and n40737_not n40740 ; n40741
g40486 and n40461_not n40741_not ; n40742
g40487 and b[22] n40450_not ; n40743
g40488 and n40444_not n40743 ; n40744
g40489 and n40452_not n40744_not ; n40745
g40490 and n40742_not n40745 ; n40746
g40491 and n40452_not n40746_not ; n40747
g40492 and b[23] n40441_not ; n40748
g40493 and n40435_not n40748 ; n40749
g40494 and n40443_not n40749_not ; n40750
g40495 and n40747_not n40750 ; n40751
g40496 and n40443_not n40751_not ; n40752
g40497 and b[24] n40432_not ; n40753
g40498 and n40426_not n40753 ; n40754
g40499 and n40434_not n40754_not ; n40755
g40500 and n40752_not n40755 ; n40756
g40501 and n40434_not n40756_not ; n40757
g40502 and b[25] n40423_not ; n40758
g40503 and n40417_not n40758 ; n40759
g40504 and n40425_not n40759_not ; n40760
g40505 and n40757_not n40760 ; n40761
g40506 and n40425_not n40761_not ; n40762
g40507 and b[26] n40414_not ; n40763
g40508 and n40408_not n40763 ; n40764
g40509 and n40416_not n40764_not ; n40765
g40510 and n40762_not n40765 ; n40766
g40511 and n40416_not n40766_not ; n40767
g40512 and b[27] n40405_not ; n40768
g40513 and n40399_not n40768 ; n40769
g40514 and n40407_not n40769_not ; n40770
g40515 and n40767_not n40770 ; n40771
g40516 and n40407_not n40771_not ; n40772
g40517 and b[28] n40396_not ; n40773
g40518 and n40390_not n40773 ; n40774
g40519 and n40398_not n40774_not ; n40775
g40520 and n40772_not n40775 ; n40776
g40521 and n40398_not n40776_not ; n40777
g40522 and b[29] n40387_not ; n40778
g40523 and n40381_not n40778 ; n40779
g40524 and n40389_not n40779_not ; n40780
g40525 and n40777_not n40780 ; n40781
g40526 and n40389_not n40781_not ; n40782
g40527 and b[30] n40378_not ; n40783
g40528 and n40372_not n40783 ; n40784
g40529 and n40380_not n40784_not ; n40785
g40530 and n40782_not n40785 ; n40786
g40531 and n40380_not n40786_not ; n40787
g40532 and b[31] n40369_not ; n40788
g40533 and n40363_not n40788 ; n40789
g40534 and n40371_not n40789_not ; n40790
g40535 and n40787_not n40790 ; n40791
g40536 and n40371_not n40791_not ; n40792
g40537 and b[32] n40360_not ; n40793
g40538 and n40354_not n40793 ; n40794
g40539 and n40362_not n40794_not ; n40795
g40540 and n40792_not n40795 ; n40796
g40541 and n40362_not n40796_not ; n40797
g40542 and b[33] n40351_not ; n40798
g40543 and n40345_not n40798 ; n40799
g40544 and n40353_not n40799_not ; n40800
g40545 and n40797_not n40800 ; n40801
g40546 and n40353_not n40801_not ; n40802
g40547 and b[34] n40342_not ; n40803
g40548 and n40336_not n40803 ; n40804
g40549 and n40344_not n40804_not ; n40805
g40550 and n40802_not n40805 ; n40806
g40551 and n40344_not n40806_not ; n40807
g40552 and b[35] n40333_not ; n40808
g40553 and n40327_not n40808 ; n40809
g40554 and n40335_not n40809_not ; n40810
g40555 and n40807_not n40810 ; n40811
g40556 and n40335_not n40811_not ; n40812
g40557 and b[36] n40324_not ; n40813
g40558 and n40318_not n40813 ; n40814
g40559 and n40326_not n40814_not ; n40815
g40560 and n40812_not n40815 ; n40816
g40561 and n40326_not n40816_not ; n40817
g40562 and b[37] n40315_not ; n40818
g40563 and n40309_not n40818 ; n40819
g40564 and n40317_not n40819_not ; n40820
g40565 and n40817_not n40820 ; n40821
g40566 and n40317_not n40821_not ; n40822
g40567 and b[38] n40306_not ; n40823
g40568 and n40300_not n40823 ; n40824
g40569 and n40308_not n40824_not ; n40825
g40570 and n40822_not n40825 ; n40826
g40571 and n40308_not n40826_not ; n40827
g40572 and b[39] n40297_not ; n40828
g40573 and n40291_not n40828 ; n40829
g40574 and n40299_not n40829_not ; n40830
g40575 and n40827_not n40830 ; n40831
g40576 and n40299_not n40831_not ; n40832
g40577 and b[40] n40288_not ; n40833
g40578 and n40282_not n40833 ; n40834
g40579 and n40290_not n40834_not ; n40835
g40580 and n40832_not n40835 ; n40836
g40581 and n40290_not n40836_not ; n40837
g40582 and n39740_not n40281_not ; n40838
g40583 and n39742_not n40278 ; n40839
g40584 and n40274_not n40839 ; n40840
g40585 and n40275_not n40278_not ; n40841
g40586 and n40840_not n40841_not ; n40842
g40587 and n40281 n40842_not ; n40843
g40588 and n40838_not n40843_not ; n40844
g40589 and b[41]_not n40844_not ; n40845
g40590 and b[41] n40838_not ; n40846
g40591 and n40843_not n40846 ; n40847
g40592 and n12761 n40847_not ; n40848
g40593 and n40845_not n40848 ; n40849
g40594 and n40837_not n40849 ; n40850
g40595 and n12184 n40844_not ; n40851
g40596 and n40850_not n40851_not ; n40852
g40597 and n40299_not n40835 ; n40853
g40598 and n40831_not n40853 ; n40854
g40599 and n40832_not n40835_not ; n40855
g40600 and n40854_not n40855_not ; n40856
g40601 and n40852_not n40856_not ; n40857
g40602 and n40289_not n40851_not ; n40858
g40603 and n40850_not n40858 ; n40859
g40604 and n40857_not n40859_not ; n40860
g40605 and n40290_not n40847_not ; n40861
g40606 and n40845_not n40861 ; n40862
g40607 and n40836_not n40862 ; n40863
g40608 and n40845_not n40847_not ; n40864
g40609 and n40837_not n40864_not ; n40865
g40610 and n40863_not n40865_not ; n40866
g40611 and n40852_not n40866_not ; n40867
g40612 and n40844_not n40851_not ; n40868
g40613 and n40850_not n40868 ; n40869
g40614 and n40867_not n40869_not ; n40870
g40615 and b[42]_not n40870_not ; n40871
g40616 and b[41]_not n40860_not ; n40872
g40617 and n40308_not n40830 ; n40873
g40618 and n40826_not n40873 ; n40874
g40619 and n40827_not n40830_not ; n40875
g40620 and n40874_not n40875_not ; n40876
g40621 and n40852_not n40876_not ; n40877
g40622 and n40298_not n40851_not ; n40878
g40623 and n40850_not n40878 ; n40879
g40624 and n40877_not n40879_not ; n40880
g40625 and b[40]_not n40880_not ; n40881
g40626 and n40317_not n40825 ; n40882
g40627 and n40821_not n40882 ; n40883
g40628 and n40822_not n40825_not ; n40884
g40629 and n40883_not n40884_not ; n40885
g40630 and n40852_not n40885_not ; n40886
g40631 and n40307_not n40851_not ; n40887
g40632 and n40850_not n40887 ; n40888
g40633 and n40886_not n40888_not ; n40889
g40634 and b[39]_not n40889_not ; n40890
g40635 and n40326_not n40820 ; n40891
g40636 and n40816_not n40891 ; n40892
g40637 and n40817_not n40820_not ; n40893
g40638 and n40892_not n40893_not ; n40894
g40639 and n40852_not n40894_not ; n40895
g40640 and n40316_not n40851_not ; n40896
g40641 and n40850_not n40896 ; n40897
g40642 and n40895_not n40897_not ; n40898
g40643 and b[38]_not n40898_not ; n40899
g40644 and n40335_not n40815 ; n40900
g40645 and n40811_not n40900 ; n40901
g40646 and n40812_not n40815_not ; n40902
g40647 and n40901_not n40902_not ; n40903
g40648 and n40852_not n40903_not ; n40904
g40649 and n40325_not n40851_not ; n40905
g40650 and n40850_not n40905 ; n40906
g40651 and n40904_not n40906_not ; n40907
g40652 and b[37]_not n40907_not ; n40908
g40653 and n40344_not n40810 ; n40909
g40654 and n40806_not n40909 ; n40910
g40655 and n40807_not n40810_not ; n40911
g40656 and n40910_not n40911_not ; n40912
g40657 and n40852_not n40912_not ; n40913
g40658 and n40334_not n40851_not ; n40914
g40659 and n40850_not n40914 ; n40915
g40660 and n40913_not n40915_not ; n40916
g40661 and b[36]_not n40916_not ; n40917
g40662 and n40353_not n40805 ; n40918
g40663 and n40801_not n40918 ; n40919
g40664 and n40802_not n40805_not ; n40920
g40665 and n40919_not n40920_not ; n40921
g40666 and n40852_not n40921_not ; n40922
g40667 and n40343_not n40851_not ; n40923
g40668 and n40850_not n40923 ; n40924
g40669 and n40922_not n40924_not ; n40925
g40670 and b[35]_not n40925_not ; n40926
g40671 and n40362_not n40800 ; n40927
g40672 and n40796_not n40927 ; n40928
g40673 and n40797_not n40800_not ; n40929
g40674 and n40928_not n40929_not ; n40930
g40675 and n40852_not n40930_not ; n40931
g40676 and n40352_not n40851_not ; n40932
g40677 and n40850_not n40932 ; n40933
g40678 and n40931_not n40933_not ; n40934
g40679 and b[34]_not n40934_not ; n40935
g40680 and n40371_not n40795 ; n40936
g40681 and n40791_not n40936 ; n40937
g40682 and n40792_not n40795_not ; n40938
g40683 and n40937_not n40938_not ; n40939
g40684 and n40852_not n40939_not ; n40940
g40685 and n40361_not n40851_not ; n40941
g40686 and n40850_not n40941 ; n40942
g40687 and n40940_not n40942_not ; n40943
g40688 and b[33]_not n40943_not ; n40944
g40689 and n40380_not n40790 ; n40945
g40690 and n40786_not n40945 ; n40946
g40691 and n40787_not n40790_not ; n40947
g40692 and n40946_not n40947_not ; n40948
g40693 and n40852_not n40948_not ; n40949
g40694 and n40370_not n40851_not ; n40950
g40695 and n40850_not n40950 ; n40951
g40696 and n40949_not n40951_not ; n40952
g40697 and b[32]_not n40952_not ; n40953
g40698 and n40389_not n40785 ; n40954
g40699 and n40781_not n40954 ; n40955
g40700 and n40782_not n40785_not ; n40956
g40701 and n40955_not n40956_not ; n40957
g40702 and n40852_not n40957_not ; n40958
g40703 and n40379_not n40851_not ; n40959
g40704 and n40850_not n40959 ; n40960
g40705 and n40958_not n40960_not ; n40961
g40706 and b[31]_not n40961_not ; n40962
g40707 and n40398_not n40780 ; n40963
g40708 and n40776_not n40963 ; n40964
g40709 and n40777_not n40780_not ; n40965
g40710 and n40964_not n40965_not ; n40966
g40711 and n40852_not n40966_not ; n40967
g40712 and n40388_not n40851_not ; n40968
g40713 and n40850_not n40968 ; n40969
g40714 and n40967_not n40969_not ; n40970
g40715 and b[30]_not n40970_not ; n40971
g40716 and n40407_not n40775 ; n40972
g40717 and n40771_not n40972 ; n40973
g40718 and n40772_not n40775_not ; n40974
g40719 and n40973_not n40974_not ; n40975
g40720 and n40852_not n40975_not ; n40976
g40721 and n40397_not n40851_not ; n40977
g40722 and n40850_not n40977 ; n40978
g40723 and n40976_not n40978_not ; n40979
g40724 and b[29]_not n40979_not ; n40980
g40725 and n40416_not n40770 ; n40981
g40726 and n40766_not n40981 ; n40982
g40727 and n40767_not n40770_not ; n40983
g40728 and n40982_not n40983_not ; n40984
g40729 and n40852_not n40984_not ; n40985
g40730 and n40406_not n40851_not ; n40986
g40731 and n40850_not n40986 ; n40987
g40732 and n40985_not n40987_not ; n40988
g40733 and b[28]_not n40988_not ; n40989
g40734 and n40425_not n40765 ; n40990
g40735 and n40761_not n40990 ; n40991
g40736 and n40762_not n40765_not ; n40992
g40737 and n40991_not n40992_not ; n40993
g40738 and n40852_not n40993_not ; n40994
g40739 and n40415_not n40851_not ; n40995
g40740 and n40850_not n40995 ; n40996
g40741 and n40994_not n40996_not ; n40997
g40742 and b[27]_not n40997_not ; n40998
g40743 and n40434_not n40760 ; n40999
g40744 and n40756_not n40999 ; n41000
g40745 and n40757_not n40760_not ; n41001
g40746 and n41000_not n41001_not ; n41002
g40747 and n40852_not n41002_not ; n41003
g40748 and n40424_not n40851_not ; n41004
g40749 and n40850_not n41004 ; n41005
g40750 and n41003_not n41005_not ; n41006
g40751 and b[26]_not n41006_not ; n41007
g40752 and n40443_not n40755 ; n41008
g40753 and n40751_not n41008 ; n41009
g40754 and n40752_not n40755_not ; n41010
g40755 and n41009_not n41010_not ; n41011
g40756 and n40852_not n41011_not ; n41012
g40757 and n40433_not n40851_not ; n41013
g40758 and n40850_not n41013 ; n41014
g40759 and n41012_not n41014_not ; n41015
g40760 and b[25]_not n41015_not ; n41016
g40761 and n40452_not n40750 ; n41017
g40762 and n40746_not n41017 ; n41018
g40763 and n40747_not n40750_not ; n41019
g40764 and n41018_not n41019_not ; n41020
g40765 and n40852_not n41020_not ; n41021
g40766 and n40442_not n40851_not ; n41022
g40767 and n40850_not n41022 ; n41023
g40768 and n41021_not n41023_not ; n41024
g40769 and b[24]_not n41024_not ; n41025
g40770 and n40461_not n40745 ; n41026
g40771 and n40741_not n41026 ; n41027
g40772 and n40742_not n40745_not ; n41028
g40773 and n41027_not n41028_not ; n41029
g40774 and n40852_not n41029_not ; n41030
g40775 and n40451_not n40851_not ; n41031
g40776 and n40850_not n41031 ; n41032
g40777 and n41030_not n41032_not ; n41033
g40778 and b[23]_not n41033_not ; n41034
g40779 and n40470_not n40740 ; n41035
g40780 and n40736_not n41035 ; n41036
g40781 and n40737_not n40740_not ; n41037
g40782 and n41036_not n41037_not ; n41038
g40783 and n40852_not n41038_not ; n41039
g40784 and n40460_not n40851_not ; n41040
g40785 and n40850_not n41040 ; n41041
g40786 and n41039_not n41041_not ; n41042
g40787 and b[22]_not n41042_not ; n41043
g40788 and n40479_not n40735 ; n41044
g40789 and n40731_not n41044 ; n41045
g40790 and n40732_not n40735_not ; n41046
g40791 and n41045_not n41046_not ; n41047
g40792 and n40852_not n41047_not ; n41048
g40793 and n40469_not n40851_not ; n41049
g40794 and n40850_not n41049 ; n41050
g40795 and n41048_not n41050_not ; n41051
g40796 and b[21]_not n41051_not ; n41052
g40797 and n40488_not n40730 ; n41053
g40798 and n40726_not n41053 ; n41054
g40799 and n40727_not n40730_not ; n41055
g40800 and n41054_not n41055_not ; n41056
g40801 and n40852_not n41056_not ; n41057
g40802 and n40478_not n40851_not ; n41058
g40803 and n40850_not n41058 ; n41059
g40804 and n41057_not n41059_not ; n41060
g40805 and b[20]_not n41060_not ; n41061
g40806 and n40497_not n40725 ; n41062
g40807 and n40721_not n41062 ; n41063
g40808 and n40722_not n40725_not ; n41064
g40809 and n41063_not n41064_not ; n41065
g40810 and n40852_not n41065_not ; n41066
g40811 and n40487_not n40851_not ; n41067
g40812 and n40850_not n41067 ; n41068
g40813 and n41066_not n41068_not ; n41069
g40814 and b[19]_not n41069_not ; n41070
g40815 and n40506_not n40720 ; n41071
g40816 and n40716_not n41071 ; n41072
g40817 and n40717_not n40720_not ; n41073
g40818 and n41072_not n41073_not ; n41074
g40819 and n40852_not n41074_not ; n41075
g40820 and n40496_not n40851_not ; n41076
g40821 and n40850_not n41076 ; n41077
g40822 and n41075_not n41077_not ; n41078
g40823 and b[18]_not n41078_not ; n41079
g40824 and n40515_not n40715 ; n41080
g40825 and n40711_not n41080 ; n41081
g40826 and n40712_not n40715_not ; n41082
g40827 and n41081_not n41082_not ; n41083
g40828 and n40852_not n41083_not ; n41084
g40829 and n40505_not n40851_not ; n41085
g40830 and n40850_not n41085 ; n41086
g40831 and n41084_not n41086_not ; n41087
g40832 and b[17]_not n41087_not ; n41088
g40833 and n40524_not n40710 ; n41089
g40834 and n40706_not n41089 ; n41090
g40835 and n40707_not n40710_not ; n41091
g40836 and n41090_not n41091_not ; n41092
g40837 and n40852_not n41092_not ; n41093
g40838 and n40514_not n40851_not ; n41094
g40839 and n40850_not n41094 ; n41095
g40840 and n41093_not n41095_not ; n41096
g40841 and b[16]_not n41096_not ; n41097
g40842 and n40533_not n40705 ; n41098
g40843 and n40701_not n41098 ; n41099
g40844 and n40702_not n40705_not ; n41100
g40845 and n41099_not n41100_not ; n41101
g40846 and n40852_not n41101_not ; n41102
g40847 and n40523_not n40851_not ; n41103
g40848 and n40850_not n41103 ; n41104
g40849 and n41102_not n41104_not ; n41105
g40850 and b[15]_not n41105_not ; n41106
g40851 and n40542_not n40700 ; n41107
g40852 and n40696_not n41107 ; n41108
g40853 and n40697_not n40700_not ; n41109
g40854 and n41108_not n41109_not ; n41110
g40855 and n40852_not n41110_not ; n41111
g40856 and n40532_not n40851_not ; n41112
g40857 and n40850_not n41112 ; n41113
g40858 and n41111_not n41113_not ; n41114
g40859 and b[14]_not n41114_not ; n41115
g40860 and n40551_not n40695 ; n41116
g40861 and n40691_not n41116 ; n41117
g40862 and n40692_not n40695_not ; n41118
g40863 and n41117_not n41118_not ; n41119
g40864 and n40852_not n41119_not ; n41120
g40865 and n40541_not n40851_not ; n41121
g40866 and n40850_not n41121 ; n41122
g40867 and n41120_not n41122_not ; n41123
g40868 and b[13]_not n41123_not ; n41124
g40869 and n40560_not n40690 ; n41125
g40870 and n40686_not n41125 ; n41126
g40871 and n40687_not n40690_not ; n41127
g40872 and n41126_not n41127_not ; n41128
g40873 and n40852_not n41128_not ; n41129
g40874 and n40550_not n40851_not ; n41130
g40875 and n40850_not n41130 ; n41131
g40876 and n41129_not n41131_not ; n41132
g40877 and b[12]_not n41132_not ; n41133
g40878 and n40569_not n40685 ; n41134
g40879 and n40681_not n41134 ; n41135
g40880 and n40682_not n40685_not ; n41136
g40881 and n41135_not n41136_not ; n41137
g40882 and n40852_not n41137_not ; n41138
g40883 and n40559_not n40851_not ; n41139
g40884 and n40850_not n41139 ; n41140
g40885 and n41138_not n41140_not ; n41141
g40886 and b[11]_not n41141_not ; n41142
g40887 and n40578_not n40680 ; n41143
g40888 and n40676_not n41143 ; n41144
g40889 and n40677_not n40680_not ; n41145
g40890 and n41144_not n41145_not ; n41146
g40891 and n40852_not n41146_not ; n41147
g40892 and n40568_not n40851_not ; n41148
g40893 and n40850_not n41148 ; n41149
g40894 and n41147_not n41149_not ; n41150
g40895 and b[10]_not n41150_not ; n41151
g40896 and n40587_not n40675 ; n41152
g40897 and n40671_not n41152 ; n41153
g40898 and n40672_not n40675_not ; n41154
g40899 and n41153_not n41154_not ; n41155
g40900 and n40852_not n41155_not ; n41156
g40901 and n40577_not n40851_not ; n41157
g40902 and n40850_not n41157 ; n41158
g40903 and n41156_not n41158_not ; n41159
g40904 and b[9]_not n41159_not ; n41160
g40905 and n40596_not n40670 ; n41161
g40906 and n40666_not n41161 ; n41162
g40907 and n40667_not n40670_not ; n41163
g40908 and n41162_not n41163_not ; n41164
g40909 and n40852_not n41164_not ; n41165
g40910 and n40586_not n40851_not ; n41166
g40911 and n40850_not n41166 ; n41167
g40912 and n41165_not n41167_not ; n41168
g40913 and b[8]_not n41168_not ; n41169
g40914 and n40605_not n40665 ; n41170
g40915 and n40661_not n41170 ; n41171
g40916 and n40662_not n40665_not ; n41172
g40917 and n41171_not n41172_not ; n41173
g40918 and n40852_not n41173_not ; n41174
g40919 and n40595_not n40851_not ; n41175
g40920 and n40850_not n41175 ; n41176
g40921 and n41174_not n41176_not ; n41177
g40922 and b[7]_not n41177_not ; n41178
g40923 and n40614_not n40660 ; n41179
g40924 and n40656_not n41179 ; n41180
g40925 and n40657_not n40660_not ; n41181
g40926 and n41180_not n41181_not ; n41182
g40927 and n40852_not n41182_not ; n41183
g40928 and n40604_not n40851_not ; n41184
g40929 and n40850_not n41184 ; n41185
g40930 and n41183_not n41185_not ; n41186
g40931 and b[6]_not n41186_not ; n41187
g40932 and n40623_not n40655 ; n41188
g40933 and n40651_not n41188 ; n41189
g40934 and n40652_not n40655_not ; n41190
g40935 and n41189_not n41190_not ; n41191
g40936 and n40852_not n41191_not ; n41192
g40937 and n40613_not n40851_not ; n41193
g40938 and n40850_not n41193 ; n41194
g40939 and n41192_not n41194_not ; n41195
g40940 and b[5]_not n41195_not ; n41196
g40941 and n40631_not n40650 ; n41197
g40942 and n40646_not n41197 ; n41198
g40943 and n40647_not n40650_not ; n41199
g40944 and n41198_not n41199_not ; n41200
g40945 and n40852_not n41200_not ; n41201
g40946 and n40622_not n40851_not ; n41202
g40947 and n40850_not n41202 ; n41203
g40948 and n41201_not n41203_not ; n41204
g40949 and b[4]_not n41204_not ; n41205
g40950 and n40641_not n40645 ; n41206
g40951 and n40640_not n41206 ; n41207
g40952 and n40642_not n40645_not ; n41208
g40953 and n41207_not n41208_not ; n41209
g40954 and n40852_not n41209_not ; n41210
g40955 and n40630_not n40851_not ; n41211
g40956 and n40850_not n41211 ; n41212
g40957 and n41210_not n41212_not ; n41213
g40958 and b[3]_not n41213_not ; n41214
g40959 and n12551 n40638_not ; n41215
g40960 and n40636_not n41215 ; n41216
g40961 and n40640_not n41216_not ; n41217
g40962 and n40852_not n41217 ; n41218
g40963 and n40635_not n40851_not ; n41219
g40964 and n40850_not n41219 ; n41220
g40965 and n41218_not n41220_not ; n41221
g40966 and b[2]_not n41221_not ; n41222
g40967 and b[0] n40852_not ; n41223
g40968 and a[22] n41223_not ; n41224
g40969 and n12551 n40852_not ; n41225
g40970 and n41224_not n41225_not ; n41226
g40971 and b[1] n41226_not ; n41227
g40972 and b[1]_not n41225_not ; n41228
g40973 and n41224_not n41228 ; n41229
g40974 and n41227_not n41229_not ; n41230
g40975 and n13145_not n41230_not ; n41231
g40976 and b[1]_not n41226_not ; n41232
g40977 and n41231_not n41232_not ; n41233
g40978 and b[2] n41220_not ; n41234
g40979 and n41218_not n41234 ; n41235
g40980 and n41222_not n41235_not ; n41236
g40981 and n41233_not n41236 ; n41237
g40982 and n41222_not n41237_not ; n41238
g40983 and b[3] n41212_not ; n41239
g40984 and n41210_not n41239 ; n41240
g40985 and n41214_not n41240_not ; n41241
g40986 and n41238_not n41241 ; n41242
g40987 and n41214_not n41242_not ; n41243
g40988 and b[4] n41203_not ; n41244
g40989 and n41201_not n41244 ; n41245
g40990 and n41205_not n41245_not ; n41246
g40991 and n41243_not n41246 ; n41247
g40992 and n41205_not n41247_not ; n41248
g40993 and b[5] n41194_not ; n41249
g40994 and n41192_not n41249 ; n41250
g40995 and n41196_not n41250_not ; n41251
g40996 and n41248_not n41251 ; n41252
g40997 and n41196_not n41252_not ; n41253
g40998 and b[6] n41185_not ; n41254
g40999 and n41183_not n41254 ; n41255
g41000 and n41187_not n41255_not ; n41256
g41001 and n41253_not n41256 ; n41257
g41002 and n41187_not n41257_not ; n41258
g41003 and b[7] n41176_not ; n41259
g41004 and n41174_not n41259 ; n41260
g41005 and n41178_not n41260_not ; n41261
g41006 and n41258_not n41261 ; n41262
g41007 and n41178_not n41262_not ; n41263
g41008 and b[8] n41167_not ; n41264
g41009 and n41165_not n41264 ; n41265
g41010 and n41169_not n41265_not ; n41266
g41011 and n41263_not n41266 ; n41267
g41012 and n41169_not n41267_not ; n41268
g41013 and b[9] n41158_not ; n41269
g41014 and n41156_not n41269 ; n41270
g41015 and n41160_not n41270_not ; n41271
g41016 and n41268_not n41271 ; n41272
g41017 and n41160_not n41272_not ; n41273
g41018 and b[10] n41149_not ; n41274
g41019 and n41147_not n41274 ; n41275
g41020 and n41151_not n41275_not ; n41276
g41021 and n41273_not n41276 ; n41277
g41022 and n41151_not n41277_not ; n41278
g41023 and b[11] n41140_not ; n41279
g41024 and n41138_not n41279 ; n41280
g41025 and n41142_not n41280_not ; n41281
g41026 and n41278_not n41281 ; n41282
g41027 and n41142_not n41282_not ; n41283
g41028 and b[12] n41131_not ; n41284
g41029 and n41129_not n41284 ; n41285
g41030 and n41133_not n41285_not ; n41286
g41031 and n41283_not n41286 ; n41287
g41032 and n41133_not n41287_not ; n41288
g41033 and b[13] n41122_not ; n41289
g41034 and n41120_not n41289 ; n41290
g41035 and n41124_not n41290_not ; n41291
g41036 and n41288_not n41291 ; n41292
g41037 and n41124_not n41292_not ; n41293
g41038 and b[14] n41113_not ; n41294
g41039 and n41111_not n41294 ; n41295
g41040 and n41115_not n41295_not ; n41296
g41041 and n41293_not n41296 ; n41297
g41042 and n41115_not n41297_not ; n41298
g41043 and b[15] n41104_not ; n41299
g41044 and n41102_not n41299 ; n41300
g41045 and n41106_not n41300_not ; n41301
g41046 and n41298_not n41301 ; n41302
g41047 and n41106_not n41302_not ; n41303
g41048 and b[16] n41095_not ; n41304
g41049 and n41093_not n41304 ; n41305
g41050 and n41097_not n41305_not ; n41306
g41051 and n41303_not n41306 ; n41307
g41052 and n41097_not n41307_not ; n41308
g41053 and b[17] n41086_not ; n41309
g41054 and n41084_not n41309 ; n41310
g41055 and n41088_not n41310_not ; n41311
g41056 and n41308_not n41311 ; n41312
g41057 and n41088_not n41312_not ; n41313
g41058 and b[18] n41077_not ; n41314
g41059 and n41075_not n41314 ; n41315
g41060 and n41079_not n41315_not ; n41316
g41061 and n41313_not n41316 ; n41317
g41062 and n41079_not n41317_not ; n41318
g41063 and b[19] n41068_not ; n41319
g41064 and n41066_not n41319 ; n41320
g41065 and n41070_not n41320_not ; n41321
g41066 and n41318_not n41321 ; n41322
g41067 and n41070_not n41322_not ; n41323
g41068 and b[20] n41059_not ; n41324
g41069 and n41057_not n41324 ; n41325
g41070 and n41061_not n41325_not ; n41326
g41071 and n41323_not n41326 ; n41327
g41072 and n41061_not n41327_not ; n41328
g41073 and b[21] n41050_not ; n41329
g41074 and n41048_not n41329 ; n41330
g41075 and n41052_not n41330_not ; n41331
g41076 and n41328_not n41331 ; n41332
g41077 and n41052_not n41332_not ; n41333
g41078 and b[22] n41041_not ; n41334
g41079 and n41039_not n41334 ; n41335
g41080 and n41043_not n41335_not ; n41336
g41081 and n41333_not n41336 ; n41337
g41082 and n41043_not n41337_not ; n41338
g41083 and b[23] n41032_not ; n41339
g41084 and n41030_not n41339 ; n41340
g41085 and n41034_not n41340_not ; n41341
g41086 and n41338_not n41341 ; n41342
g41087 and n41034_not n41342_not ; n41343
g41088 and b[24] n41023_not ; n41344
g41089 and n41021_not n41344 ; n41345
g41090 and n41025_not n41345_not ; n41346
g41091 and n41343_not n41346 ; n41347
g41092 and n41025_not n41347_not ; n41348
g41093 and b[25] n41014_not ; n41349
g41094 and n41012_not n41349 ; n41350
g41095 and n41016_not n41350_not ; n41351
g41096 and n41348_not n41351 ; n41352
g41097 and n41016_not n41352_not ; n41353
g41098 and b[26] n41005_not ; n41354
g41099 and n41003_not n41354 ; n41355
g41100 and n41007_not n41355_not ; n41356
g41101 and n41353_not n41356 ; n41357
g41102 and n41007_not n41357_not ; n41358
g41103 and b[27] n40996_not ; n41359
g41104 and n40994_not n41359 ; n41360
g41105 and n40998_not n41360_not ; n41361
g41106 and n41358_not n41361 ; n41362
g41107 and n40998_not n41362_not ; n41363
g41108 and b[28] n40987_not ; n41364
g41109 and n40985_not n41364 ; n41365
g41110 and n40989_not n41365_not ; n41366
g41111 and n41363_not n41366 ; n41367
g41112 and n40989_not n41367_not ; n41368
g41113 and b[29] n40978_not ; n41369
g41114 and n40976_not n41369 ; n41370
g41115 and n40980_not n41370_not ; n41371
g41116 and n41368_not n41371 ; n41372
g41117 and n40980_not n41372_not ; n41373
g41118 and b[30] n40969_not ; n41374
g41119 and n40967_not n41374 ; n41375
g41120 and n40971_not n41375_not ; n41376
g41121 and n41373_not n41376 ; n41377
g41122 and n40971_not n41377_not ; n41378
g41123 and b[31] n40960_not ; n41379
g41124 and n40958_not n41379 ; n41380
g41125 and n40962_not n41380_not ; n41381
g41126 and n41378_not n41381 ; n41382
g41127 and n40962_not n41382_not ; n41383
g41128 and b[32] n40951_not ; n41384
g41129 and n40949_not n41384 ; n41385
g41130 and n40953_not n41385_not ; n41386
g41131 and n41383_not n41386 ; n41387
g41132 and n40953_not n41387_not ; n41388
g41133 and b[33] n40942_not ; n41389
g41134 and n40940_not n41389 ; n41390
g41135 and n40944_not n41390_not ; n41391
g41136 and n41388_not n41391 ; n41392
g41137 and n40944_not n41392_not ; n41393
g41138 and b[34] n40933_not ; n41394
g41139 and n40931_not n41394 ; n41395
g41140 and n40935_not n41395_not ; n41396
g41141 and n41393_not n41396 ; n41397
g41142 and n40935_not n41397_not ; n41398
g41143 and b[35] n40924_not ; n41399
g41144 and n40922_not n41399 ; n41400
g41145 and n40926_not n41400_not ; n41401
g41146 and n41398_not n41401 ; n41402
g41147 and n40926_not n41402_not ; n41403
g41148 and b[36] n40915_not ; n41404
g41149 and n40913_not n41404 ; n41405
g41150 and n40917_not n41405_not ; n41406
g41151 and n41403_not n41406 ; n41407
g41152 and n40917_not n41407_not ; n41408
g41153 and b[37] n40906_not ; n41409
g41154 and n40904_not n41409 ; n41410
g41155 and n40908_not n41410_not ; n41411
g41156 and n41408_not n41411 ; n41412
g41157 and n40908_not n41412_not ; n41413
g41158 and b[38] n40897_not ; n41414
g41159 and n40895_not n41414 ; n41415
g41160 and n40899_not n41415_not ; n41416
g41161 and n41413_not n41416 ; n41417
g41162 and n40899_not n41417_not ; n41418
g41163 and b[39] n40888_not ; n41419
g41164 and n40886_not n41419 ; n41420
g41165 and n40890_not n41420_not ; n41421
g41166 and n41418_not n41421 ; n41422
g41167 and n40890_not n41422_not ; n41423
g41168 and b[40] n40879_not ; n41424
g41169 and n40877_not n41424 ; n41425
g41170 and n40881_not n41425_not ; n41426
g41171 and n41423_not n41426 ; n41427
g41172 and n40881_not n41427_not ; n41428
g41173 and b[41] n40859_not ; n41429
g41174 and n40857_not n41429 ; n41430
g41175 and n40872_not n41430_not ; n41431
g41176 and n41428_not n41431 ; n41432
g41177 and n40872_not n41432_not ; n41433
g41178 and b[42] n40869_not ; n41434
g41179 and n40867_not n41434 ; n41435
g41180 and n40871_not n41435_not ; n41436
g41181 and n41433_not n41436 ; n41437
g41182 and n40871_not n41437_not ; n41438
g41183 and n13355 n41438_not ; n41439
g41184 and n40860_not n41439_not ; n41440
g41185 and n40881_not n41431 ; n41441
g41186 and n41427_not n41441 ; n41442
g41187 and n41428_not n41431_not ; n41443
g41188 and n41442_not n41443_not ; n41444
g41189 and n13355 n41444_not ; n41445
g41190 and n41438_not n41445 ; n41446
g41191 and n41440_not n41446_not ; n41447
g41192 and b[42]_not n41447_not ; n41448
g41193 and n40880_not n41439_not ; n41449
g41194 and n40890_not n41426 ; n41450
g41195 and n41422_not n41450 ; n41451
g41196 and n41423_not n41426_not ; n41452
g41197 and n41451_not n41452_not ; n41453
g41198 and n13355 n41453_not ; n41454
g41199 and n41438_not n41454 ; n41455
g41200 and n41449_not n41455_not ; n41456
g41201 and b[41]_not n41456_not ; n41457
g41202 and n40889_not n41439_not ; n41458
g41203 and n40899_not n41421 ; n41459
g41204 and n41417_not n41459 ; n41460
g41205 and n41418_not n41421_not ; n41461
g41206 and n41460_not n41461_not ; n41462
g41207 and n13355 n41462_not ; n41463
g41208 and n41438_not n41463 ; n41464
g41209 and n41458_not n41464_not ; n41465
g41210 and b[40]_not n41465_not ; n41466
g41211 and n40898_not n41439_not ; n41467
g41212 and n40908_not n41416 ; n41468
g41213 and n41412_not n41468 ; n41469
g41214 and n41413_not n41416_not ; n41470
g41215 and n41469_not n41470_not ; n41471
g41216 and n13355 n41471_not ; n41472
g41217 and n41438_not n41472 ; n41473
g41218 and n41467_not n41473_not ; n41474
g41219 and b[39]_not n41474_not ; n41475
g41220 and n40907_not n41439_not ; n41476
g41221 and n40917_not n41411 ; n41477
g41222 and n41407_not n41477 ; n41478
g41223 and n41408_not n41411_not ; n41479
g41224 and n41478_not n41479_not ; n41480
g41225 and n13355 n41480_not ; n41481
g41226 and n41438_not n41481 ; n41482
g41227 and n41476_not n41482_not ; n41483
g41228 and b[38]_not n41483_not ; n41484
g41229 and n40916_not n41439_not ; n41485
g41230 and n40926_not n41406 ; n41486
g41231 and n41402_not n41486 ; n41487
g41232 and n41403_not n41406_not ; n41488
g41233 and n41487_not n41488_not ; n41489
g41234 and n13355 n41489_not ; n41490
g41235 and n41438_not n41490 ; n41491
g41236 and n41485_not n41491_not ; n41492
g41237 and b[37]_not n41492_not ; n41493
g41238 and n40925_not n41439_not ; n41494
g41239 and n40935_not n41401 ; n41495
g41240 and n41397_not n41495 ; n41496
g41241 and n41398_not n41401_not ; n41497
g41242 and n41496_not n41497_not ; n41498
g41243 and n13355 n41498_not ; n41499
g41244 and n41438_not n41499 ; n41500
g41245 and n41494_not n41500_not ; n41501
g41246 and b[36]_not n41501_not ; n41502
g41247 and n40934_not n41439_not ; n41503
g41248 and n40944_not n41396 ; n41504
g41249 and n41392_not n41504 ; n41505
g41250 and n41393_not n41396_not ; n41506
g41251 and n41505_not n41506_not ; n41507
g41252 and n13355 n41507_not ; n41508
g41253 and n41438_not n41508 ; n41509
g41254 and n41503_not n41509_not ; n41510
g41255 and b[35]_not n41510_not ; n41511
g41256 and n40943_not n41439_not ; n41512
g41257 and n40953_not n41391 ; n41513
g41258 and n41387_not n41513 ; n41514
g41259 and n41388_not n41391_not ; n41515
g41260 and n41514_not n41515_not ; n41516
g41261 and n13355 n41516_not ; n41517
g41262 and n41438_not n41517 ; n41518
g41263 and n41512_not n41518_not ; n41519
g41264 and b[34]_not n41519_not ; n41520
g41265 and n40952_not n41439_not ; n41521
g41266 and n40962_not n41386 ; n41522
g41267 and n41382_not n41522 ; n41523
g41268 and n41383_not n41386_not ; n41524
g41269 and n41523_not n41524_not ; n41525
g41270 and n13355 n41525_not ; n41526
g41271 and n41438_not n41526 ; n41527
g41272 and n41521_not n41527_not ; n41528
g41273 and b[33]_not n41528_not ; n41529
g41274 and n40961_not n41439_not ; n41530
g41275 and n40971_not n41381 ; n41531
g41276 and n41377_not n41531 ; n41532
g41277 and n41378_not n41381_not ; n41533
g41278 and n41532_not n41533_not ; n41534
g41279 and n13355 n41534_not ; n41535
g41280 and n41438_not n41535 ; n41536
g41281 and n41530_not n41536_not ; n41537
g41282 and b[32]_not n41537_not ; n41538
g41283 and n40970_not n41439_not ; n41539
g41284 and n40980_not n41376 ; n41540
g41285 and n41372_not n41540 ; n41541
g41286 and n41373_not n41376_not ; n41542
g41287 and n41541_not n41542_not ; n41543
g41288 and n13355 n41543_not ; n41544
g41289 and n41438_not n41544 ; n41545
g41290 and n41539_not n41545_not ; n41546
g41291 and b[31]_not n41546_not ; n41547
g41292 and n40979_not n41439_not ; n41548
g41293 and n40989_not n41371 ; n41549
g41294 and n41367_not n41549 ; n41550
g41295 and n41368_not n41371_not ; n41551
g41296 and n41550_not n41551_not ; n41552
g41297 and n13355 n41552_not ; n41553
g41298 and n41438_not n41553 ; n41554
g41299 and n41548_not n41554_not ; n41555
g41300 and b[30]_not n41555_not ; n41556
g41301 and n40988_not n41439_not ; n41557
g41302 and n40998_not n41366 ; n41558
g41303 and n41362_not n41558 ; n41559
g41304 and n41363_not n41366_not ; n41560
g41305 and n41559_not n41560_not ; n41561
g41306 and n13355 n41561_not ; n41562
g41307 and n41438_not n41562 ; n41563
g41308 and n41557_not n41563_not ; n41564
g41309 and b[29]_not n41564_not ; n41565
g41310 and n40997_not n41439_not ; n41566
g41311 and n41007_not n41361 ; n41567
g41312 and n41357_not n41567 ; n41568
g41313 and n41358_not n41361_not ; n41569
g41314 and n41568_not n41569_not ; n41570
g41315 and n13355 n41570_not ; n41571
g41316 and n41438_not n41571 ; n41572
g41317 and n41566_not n41572_not ; n41573
g41318 and b[28]_not n41573_not ; n41574
g41319 and n41006_not n41439_not ; n41575
g41320 and n41016_not n41356 ; n41576
g41321 and n41352_not n41576 ; n41577
g41322 and n41353_not n41356_not ; n41578
g41323 and n41577_not n41578_not ; n41579
g41324 and n13355 n41579_not ; n41580
g41325 and n41438_not n41580 ; n41581
g41326 and n41575_not n41581_not ; n41582
g41327 and b[27]_not n41582_not ; n41583
g41328 and n41015_not n41439_not ; n41584
g41329 and n41025_not n41351 ; n41585
g41330 and n41347_not n41585 ; n41586
g41331 and n41348_not n41351_not ; n41587
g41332 and n41586_not n41587_not ; n41588
g41333 and n13355 n41588_not ; n41589
g41334 and n41438_not n41589 ; n41590
g41335 and n41584_not n41590_not ; n41591
g41336 and b[26]_not n41591_not ; n41592
g41337 and n41024_not n41439_not ; n41593
g41338 and n41034_not n41346 ; n41594
g41339 and n41342_not n41594 ; n41595
g41340 and n41343_not n41346_not ; n41596
g41341 and n41595_not n41596_not ; n41597
g41342 and n13355 n41597_not ; n41598
g41343 and n41438_not n41598 ; n41599
g41344 and n41593_not n41599_not ; n41600
g41345 and b[25]_not n41600_not ; n41601
g41346 and n41033_not n41439_not ; n41602
g41347 and n41043_not n41341 ; n41603
g41348 and n41337_not n41603 ; n41604
g41349 and n41338_not n41341_not ; n41605
g41350 and n41604_not n41605_not ; n41606
g41351 and n13355 n41606_not ; n41607
g41352 and n41438_not n41607 ; n41608
g41353 and n41602_not n41608_not ; n41609
g41354 and b[24]_not n41609_not ; n41610
g41355 and n41042_not n41439_not ; n41611
g41356 and n41052_not n41336 ; n41612
g41357 and n41332_not n41612 ; n41613
g41358 and n41333_not n41336_not ; n41614
g41359 and n41613_not n41614_not ; n41615
g41360 and n13355 n41615_not ; n41616
g41361 and n41438_not n41616 ; n41617
g41362 and n41611_not n41617_not ; n41618
g41363 and b[23]_not n41618_not ; n41619
g41364 and n41051_not n41439_not ; n41620
g41365 and n41061_not n41331 ; n41621
g41366 and n41327_not n41621 ; n41622
g41367 and n41328_not n41331_not ; n41623
g41368 and n41622_not n41623_not ; n41624
g41369 and n13355 n41624_not ; n41625
g41370 and n41438_not n41625 ; n41626
g41371 and n41620_not n41626_not ; n41627
g41372 and b[22]_not n41627_not ; n41628
g41373 and n41060_not n41439_not ; n41629
g41374 and n41070_not n41326 ; n41630
g41375 and n41322_not n41630 ; n41631
g41376 and n41323_not n41326_not ; n41632
g41377 and n41631_not n41632_not ; n41633
g41378 and n13355 n41633_not ; n41634
g41379 and n41438_not n41634 ; n41635
g41380 and n41629_not n41635_not ; n41636
g41381 and b[21]_not n41636_not ; n41637
g41382 and n41069_not n41439_not ; n41638
g41383 and n41079_not n41321 ; n41639
g41384 and n41317_not n41639 ; n41640
g41385 and n41318_not n41321_not ; n41641
g41386 and n41640_not n41641_not ; n41642
g41387 and n13355 n41642_not ; n41643
g41388 and n41438_not n41643 ; n41644
g41389 and n41638_not n41644_not ; n41645
g41390 and b[20]_not n41645_not ; n41646
g41391 and n41078_not n41439_not ; n41647
g41392 and n41088_not n41316 ; n41648
g41393 and n41312_not n41648 ; n41649
g41394 and n41313_not n41316_not ; n41650
g41395 and n41649_not n41650_not ; n41651
g41396 and n13355 n41651_not ; n41652
g41397 and n41438_not n41652 ; n41653
g41398 and n41647_not n41653_not ; n41654
g41399 and b[19]_not n41654_not ; n41655
g41400 and n41087_not n41439_not ; n41656
g41401 and n41097_not n41311 ; n41657
g41402 and n41307_not n41657 ; n41658
g41403 and n41308_not n41311_not ; n41659
g41404 and n41658_not n41659_not ; n41660
g41405 and n13355 n41660_not ; n41661
g41406 and n41438_not n41661 ; n41662
g41407 and n41656_not n41662_not ; n41663
g41408 and b[18]_not n41663_not ; n41664
g41409 and n41096_not n41439_not ; n41665
g41410 and n41106_not n41306 ; n41666
g41411 and n41302_not n41666 ; n41667
g41412 and n41303_not n41306_not ; n41668
g41413 and n41667_not n41668_not ; n41669
g41414 and n13355 n41669_not ; n41670
g41415 and n41438_not n41670 ; n41671
g41416 and n41665_not n41671_not ; n41672
g41417 and b[17]_not n41672_not ; n41673
g41418 and n41105_not n41439_not ; n41674
g41419 and n41115_not n41301 ; n41675
g41420 and n41297_not n41675 ; n41676
g41421 and n41298_not n41301_not ; n41677
g41422 and n41676_not n41677_not ; n41678
g41423 and n13355 n41678_not ; n41679
g41424 and n41438_not n41679 ; n41680
g41425 and n41674_not n41680_not ; n41681
g41426 and b[16]_not n41681_not ; n41682
g41427 and n41114_not n41439_not ; n41683
g41428 and n41124_not n41296 ; n41684
g41429 and n41292_not n41684 ; n41685
g41430 and n41293_not n41296_not ; n41686
g41431 and n41685_not n41686_not ; n41687
g41432 and n13355 n41687_not ; n41688
g41433 and n41438_not n41688 ; n41689
g41434 and n41683_not n41689_not ; n41690
g41435 and b[15]_not n41690_not ; n41691
g41436 and n41123_not n41439_not ; n41692
g41437 and n41133_not n41291 ; n41693
g41438 and n41287_not n41693 ; n41694
g41439 and n41288_not n41291_not ; n41695
g41440 and n41694_not n41695_not ; n41696
g41441 and n13355 n41696_not ; n41697
g41442 and n41438_not n41697 ; n41698
g41443 and n41692_not n41698_not ; n41699
g41444 and b[14]_not n41699_not ; n41700
g41445 and n41132_not n41439_not ; n41701
g41446 and n41142_not n41286 ; n41702
g41447 and n41282_not n41702 ; n41703
g41448 and n41283_not n41286_not ; n41704
g41449 and n41703_not n41704_not ; n41705
g41450 and n13355 n41705_not ; n41706
g41451 and n41438_not n41706 ; n41707
g41452 and n41701_not n41707_not ; n41708
g41453 and b[13]_not n41708_not ; n41709
g41454 and n41141_not n41439_not ; n41710
g41455 and n41151_not n41281 ; n41711
g41456 and n41277_not n41711 ; n41712
g41457 and n41278_not n41281_not ; n41713
g41458 and n41712_not n41713_not ; n41714
g41459 and n13355 n41714_not ; n41715
g41460 and n41438_not n41715 ; n41716
g41461 and n41710_not n41716_not ; n41717
g41462 and b[12]_not n41717_not ; n41718
g41463 and n41150_not n41439_not ; n41719
g41464 and n41160_not n41276 ; n41720
g41465 and n41272_not n41720 ; n41721
g41466 and n41273_not n41276_not ; n41722
g41467 and n41721_not n41722_not ; n41723
g41468 and n13355 n41723_not ; n41724
g41469 and n41438_not n41724 ; n41725
g41470 and n41719_not n41725_not ; n41726
g41471 and b[11]_not n41726_not ; n41727
g41472 and n41159_not n41439_not ; n41728
g41473 and n41169_not n41271 ; n41729
g41474 and n41267_not n41729 ; n41730
g41475 and n41268_not n41271_not ; n41731
g41476 and n41730_not n41731_not ; n41732
g41477 and n13355 n41732_not ; n41733
g41478 and n41438_not n41733 ; n41734
g41479 and n41728_not n41734_not ; n41735
g41480 and b[10]_not n41735_not ; n41736
g41481 and n41168_not n41439_not ; n41737
g41482 and n41178_not n41266 ; n41738
g41483 and n41262_not n41738 ; n41739
g41484 and n41263_not n41266_not ; n41740
g41485 and n41739_not n41740_not ; n41741
g41486 and n13355 n41741_not ; n41742
g41487 and n41438_not n41742 ; n41743
g41488 and n41737_not n41743_not ; n41744
g41489 and b[9]_not n41744_not ; n41745
g41490 and n41177_not n41439_not ; n41746
g41491 and n41187_not n41261 ; n41747
g41492 and n41257_not n41747 ; n41748
g41493 and n41258_not n41261_not ; n41749
g41494 and n41748_not n41749_not ; n41750
g41495 and n13355 n41750_not ; n41751
g41496 and n41438_not n41751 ; n41752
g41497 and n41746_not n41752_not ; n41753
g41498 and b[8]_not n41753_not ; n41754
g41499 and n41186_not n41439_not ; n41755
g41500 and n41196_not n41256 ; n41756
g41501 and n41252_not n41756 ; n41757
g41502 and n41253_not n41256_not ; n41758
g41503 and n41757_not n41758_not ; n41759
g41504 and n13355 n41759_not ; n41760
g41505 and n41438_not n41760 ; n41761
g41506 and n41755_not n41761_not ; n41762
g41507 and b[7]_not n41762_not ; n41763
g41508 and n41195_not n41439_not ; n41764
g41509 and n41205_not n41251 ; n41765
g41510 and n41247_not n41765 ; n41766
g41511 and n41248_not n41251_not ; n41767
g41512 and n41766_not n41767_not ; n41768
g41513 and n13355 n41768_not ; n41769
g41514 and n41438_not n41769 ; n41770
g41515 and n41764_not n41770_not ; n41771
g41516 and b[6]_not n41771_not ; n41772
g41517 and n41204_not n41439_not ; n41773
g41518 and n41214_not n41246 ; n41774
g41519 and n41242_not n41774 ; n41775
g41520 and n41243_not n41246_not ; n41776
g41521 and n41775_not n41776_not ; n41777
g41522 and n13355 n41777_not ; n41778
g41523 and n41438_not n41778 ; n41779
g41524 and n41773_not n41779_not ; n41780
g41525 and b[5]_not n41780_not ; n41781
g41526 and n41213_not n41439_not ; n41782
g41527 and n41222_not n41241 ; n41783
g41528 and n41237_not n41783 ; n41784
g41529 and n41238_not n41241_not ; n41785
g41530 and n41784_not n41785_not ; n41786
g41531 and n13355 n41786_not ; n41787
g41532 and n41438_not n41787 ; n41788
g41533 and n41782_not n41788_not ; n41789
g41534 and b[4]_not n41789_not ; n41790
g41535 and n41221_not n41439_not ; n41791
g41536 and n41232_not n41236 ; n41792
g41537 and n41231_not n41792 ; n41793
g41538 and n41233_not n41236_not ; n41794
g41539 and n41793_not n41794_not ; n41795
g41540 and n13355 n41795_not ; n41796
g41541 and n41438_not n41796 ; n41797
g41542 and n41791_not n41797_not ; n41798
g41543 and b[3]_not n41798_not ; n41799
g41544 and n41226_not n41439_not ; n41800
g41545 and n13145 n41229_not ; n41801
g41546 and n41227_not n41801 ; n41802
g41547 and n13355 n41802_not ; n41803
g41548 and n41231_not n41803 ; n41804
g41549 and n41438_not n41804 ; n41805
g41550 and n41800_not n41805_not ; n41806
g41551 and b[2]_not n41806_not ; n41807
g41552 and n13727 n41438_not ; n41808
g41553 and a[21] n41808_not ; n41809
g41554 and n13732 n41438_not ; n41810
g41555 and n41809_not n41810_not ; n41811
g41556 and b[1] n41811_not ; n41812
g41557 and b[1]_not n41810_not ; n41813
g41558 and n41809_not n41813 ; n41814
g41559 and n41812_not n41814_not ; n41815
g41560 and n13739_not n41815_not ; n41816
g41561 and b[1]_not n41811_not ; n41817
g41562 and n41816_not n41817_not ; n41818
g41563 and b[2] n41805_not ; n41819
g41564 and n41800_not n41819 ; n41820
g41565 and n41807_not n41820_not ; n41821
g41566 and n41818_not n41821 ; n41822
g41567 and n41807_not n41822_not ; n41823
g41568 and b[3] n41797_not ; n41824
g41569 and n41791_not n41824 ; n41825
g41570 and n41799_not n41825_not ; n41826
g41571 and n41823_not n41826 ; n41827
g41572 and n41799_not n41827_not ; n41828
g41573 and b[4] n41788_not ; n41829
g41574 and n41782_not n41829 ; n41830
g41575 and n41790_not n41830_not ; n41831
g41576 and n41828_not n41831 ; n41832
g41577 and n41790_not n41832_not ; n41833
g41578 and b[5] n41779_not ; n41834
g41579 and n41773_not n41834 ; n41835
g41580 and n41781_not n41835_not ; n41836
g41581 and n41833_not n41836 ; n41837
g41582 and n41781_not n41837_not ; n41838
g41583 and b[6] n41770_not ; n41839
g41584 and n41764_not n41839 ; n41840
g41585 and n41772_not n41840_not ; n41841
g41586 and n41838_not n41841 ; n41842
g41587 and n41772_not n41842_not ; n41843
g41588 and b[7] n41761_not ; n41844
g41589 and n41755_not n41844 ; n41845
g41590 and n41763_not n41845_not ; n41846
g41591 and n41843_not n41846 ; n41847
g41592 and n41763_not n41847_not ; n41848
g41593 and b[8] n41752_not ; n41849
g41594 and n41746_not n41849 ; n41850
g41595 and n41754_not n41850_not ; n41851
g41596 and n41848_not n41851 ; n41852
g41597 and n41754_not n41852_not ; n41853
g41598 and b[9] n41743_not ; n41854
g41599 and n41737_not n41854 ; n41855
g41600 and n41745_not n41855_not ; n41856
g41601 and n41853_not n41856 ; n41857
g41602 and n41745_not n41857_not ; n41858
g41603 and b[10] n41734_not ; n41859
g41604 and n41728_not n41859 ; n41860
g41605 and n41736_not n41860_not ; n41861
g41606 and n41858_not n41861 ; n41862
g41607 and n41736_not n41862_not ; n41863
g41608 and b[11] n41725_not ; n41864
g41609 and n41719_not n41864 ; n41865
g41610 and n41727_not n41865_not ; n41866
g41611 and n41863_not n41866 ; n41867
g41612 and n41727_not n41867_not ; n41868
g41613 and b[12] n41716_not ; n41869
g41614 and n41710_not n41869 ; n41870
g41615 and n41718_not n41870_not ; n41871
g41616 and n41868_not n41871 ; n41872
g41617 and n41718_not n41872_not ; n41873
g41618 and b[13] n41707_not ; n41874
g41619 and n41701_not n41874 ; n41875
g41620 and n41709_not n41875_not ; n41876
g41621 and n41873_not n41876 ; n41877
g41622 and n41709_not n41877_not ; n41878
g41623 and b[14] n41698_not ; n41879
g41624 and n41692_not n41879 ; n41880
g41625 and n41700_not n41880_not ; n41881
g41626 and n41878_not n41881 ; n41882
g41627 and n41700_not n41882_not ; n41883
g41628 and b[15] n41689_not ; n41884
g41629 and n41683_not n41884 ; n41885
g41630 and n41691_not n41885_not ; n41886
g41631 and n41883_not n41886 ; n41887
g41632 and n41691_not n41887_not ; n41888
g41633 and b[16] n41680_not ; n41889
g41634 and n41674_not n41889 ; n41890
g41635 and n41682_not n41890_not ; n41891
g41636 and n41888_not n41891 ; n41892
g41637 and n41682_not n41892_not ; n41893
g41638 and b[17] n41671_not ; n41894
g41639 and n41665_not n41894 ; n41895
g41640 and n41673_not n41895_not ; n41896
g41641 and n41893_not n41896 ; n41897
g41642 and n41673_not n41897_not ; n41898
g41643 and b[18] n41662_not ; n41899
g41644 and n41656_not n41899 ; n41900
g41645 and n41664_not n41900_not ; n41901
g41646 and n41898_not n41901 ; n41902
g41647 and n41664_not n41902_not ; n41903
g41648 and b[19] n41653_not ; n41904
g41649 and n41647_not n41904 ; n41905
g41650 and n41655_not n41905_not ; n41906
g41651 and n41903_not n41906 ; n41907
g41652 and n41655_not n41907_not ; n41908
g41653 and b[20] n41644_not ; n41909
g41654 and n41638_not n41909 ; n41910
g41655 and n41646_not n41910_not ; n41911
g41656 and n41908_not n41911 ; n41912
g41657 and n41646_not n41912_not ; n41913
g41658 and b[21] n41635_not ; n41914
g41659 and n41629_not n41914 ; n41915
g41660 and n41637_not n41915_not ; n41916
g41661 and n41913_not n41916 ; n41917
g41662 and n41637_not n41917_not ; n41918
g41663 and b[22] n41626_not ; n41919
g41664 and n41620_not n41919 ; n41920
g41665 and n41628_not n41920_not ; n41921
g41666 and n41918_not n41921 ; n41922
g41667 and n41628_not n41922_not ; n41923
g41668 and b[23] n41617_not ; n41924
g41669 and n41611_not n41924 ; n41925
g41670 and n41619_not n41925_not ; n41926
g41671 and n41923_not n41926 ; n41927
g41672 and n41619_not n41927_not ; n41928
g41673 and b[24] n41608_not ; n41929
g41674 and n41602_not n41929 ; n41930
g41675 and n41610_not n41930_not ; n41931
g41676 and n41928_not n41931 ; n41932
g41677 and n41610_not n41932_not ; n41933
g41678 and b[25] n41599_not ; n41934
g41679 and n41593_not n41934 ; n41935
g41680 and n41601_not n41935_not ; n41936
g41681 and n41933_not n41936 ; n41937
g41682 and n41601_not n41937_not ; n41938
g41683 and b[26] n41590_not ; n41939
g41684 and n41584_not n41939 ; n41940
g41685 and n41592_not n41940_not ; n41941
g41686 and n41938_not n41941 ; n41942
g41687 and n41592_not n41942_not ; n41943
g41688 and b[27] n41581_not ; n41944
g41689 and n41575_not n41944 ; n41945
g41690 and n41583_not n41945_not ; n41946
g41691 and n41943_not n41946 ; n41947
g41692 and n41583_not n41947_not ; n41948
g41693 and b[28] n41572_not ; n41949
g41694 and n41566_not n41949 ; n41950
g41695 and n41574_not n41950_not ; n41951
g41696 and n41948_not n41951 ; n41952
g41697 and n41574_not n41952_not ; n41953
g41698 and b[29] n41563_not ; n41954
g41699 and n41557_not n41954 ; n41955
g41700 and n41565_not n41955_not ; n41956
g41701 and n41953_not n41956 ; n41957
g41702 and n41565_not n41957_not ; n41958
g41703 and b[30] n41554_not ; n41959
g41704 and n41548_not n41959 ; n41960
g41705 and n41556_not n41960_not ; n41961
g41706 and n41958_not n41961 ; n41962
g41707 and n41556_not n41962_not ; n41963
g41708 and b[31] n41545_not ; n41964
g41709 and n41539_not n41964 ; n41965
g41710 and n41547_not n41965_not ; n41966
g41711 and n41963_not n41966 ; n41967
g41712 and n41547_not n41967_not ; n41968
g41713 and b[32] n41536_not ; n41969
g41714 and n41530_not n41969 ; n41970
g41715 and n41538_not n41970_not ; n41971
g41716 and n41968_not n41971 ; n41972
g41717 and n41538_not n41972_not ; n41973
g41718 and b[33] n41527_not ; n41974
g41719 and n41521_not n41974 ; n41975
g41720 and n41529_not n41975_not ; n41976
g41721 and n41973_not n41976 ; n41977
g41722 and n41529_not n41977_not ; n41978
g41723 and b[34] n41518_not ; n41979
g41724 and n41512_not n41979 ; n41980
g41725 and n41520_not n41980_not ; n41981
g41726 and n41978_not n41981 ; n41982
g41727 and n41520_not n41982_not ; n41983
g41728 and b[35] n41509_not ; n41984
g41729 and n41503_not n41984 ; n41985
g41730 and n41511_not n41985_not ; n41986
g41731 and n41983_not n41986 ; n41987
g41732 and n41511_not n41987_not ; n41988
g41733 and b[36] n41500_not ; n41989
g41734 and n41494_not n41989 ; n41990
g41735 and n41502_not n41990_not ; n41991
g41736 and n41988_not n41991 ; n41992
g41737 and n41502_not n41992_not ; n41993
g41738 and b[37] n41491_not ; n41994
g41739 and n41485_not n41994 ; n41995
g41740 and n41493_not n41995_not ; n41996
g41741 and n41993_not n41996 ; n41997
g41742 and n41493_not n41997_not ; n41998
g41743 and b[38] n41482_not ; n41999
g41744 and n41476_not n41999 ; n42000
g41745 and n41484_not n42000_not ; n42001
g41746 and n41998_not n42001 ; n42002
g41747 and n41484_not n42002_not ; n42003
g41748 and b[39] n41473_not ; n42004
g41749 and n41467_not n42004 ; n42005
g41750 and n41475_not n42005_not ; n42006
g41751 and n42003_not n42006 ; n42007
g41752 and n41475_not n42007_not ; n42008
g41753 and b[40] n41464_not ; n42009
g41754 and n41458_not n42009 ; n42010
g41755 and n41466_not n42010_not ; n42011
g41756 and n42008_not n42011 ; n42012
g41757 and n41466_not n42012_not ; n42013
g41758 and b[41] n41455_not ; n42014
g41759 and n41449_not n42014 ; n42015
g41760 and n41457_not n42015_not ; n42016
g41761 and n42013_not n42016 ; n42017
g41762 and n41457_not n42017_not ; n42018
g41763 and b[42] n41446_not ; n42019
g41764 and n41440_not n42019 ; n42020
g41765 and n41448_not n42020_not ; n42021
g41766 and n42018_not n42021 ; n42022
g41767 and n41448_not n42022_not ; n42023
g41768 and n40870_not n41439_not ; n42024
g41769 and n40872_not n41436 ; n42025
g41770 and n41432_not n42025 ; n42026
g41771 and n41433_not n41436_not ; n42027
g41772 and n42026_not n42027_not ; n42028
g41773 and n41439 n42028_not ; n42029
g41774 and n42024_not n42029_not ; n42030
g41775 and b[43]_not n42030_not ; n42031
g41776 and b[43] n42024_not ; n42032
g41777 and n42029_not n42032 ; n42033
g41778 and n13958 n42033_not ; n42034
g41779 and n42031_not n42034 ; n42035
g41780 and n42023_not n42035 ; n42036
g41781 and n13355 n42030_not ; n42037
g41782 and n42036_not n42037_not ; n42038
g41783 and n41457_not n42021 ; n42039
g41784 and n42017_not n42039 ; n42040
g41785 and n42018_not n42021_not ; n42041
g41786 and n42040_not n42041_not ; n42042
g41787 and n42038_not n42042_not ; n42043
g41788 and n41447_not n42037_not ; n42044
g41789 and n42036_not n42044 ; n42045
g41790 and n42043_not n42045_not ; n42046
g41791 and b[43]_not n42046_not ; n42047
g41792 and n41466_not n42016 ; n42048
g41793 and n42012_not n42048 ; n42049
g41794 and n42013_not n42016_not ; n42050
g41795 and n42049_not n42050_not ; n42051
g41796 and n42038_not n42051_not ; n42052
g41797 and n41456_not n42037_not ; n42053
g41798 and n42036_not n42053 ; n42054
g41799 and n42052_not n42054_not ; n42055
g41800 and b[42]_not n42055_not ; n42056
g41801 and n41475_not n42011 ; n42057
g41802 and n42007_not n42057 ; n42058
g41803 and n42008_not n42011_not ; n42059
g41804 and n42058_not n42059_not ; n42060
g41805 and n42038_not n42060_not ; n42061
g41806 and n41465_not n42037_not ; n42062
g41807 and n42036_not n42062 ; n42063
g41808 and n42061_not n42063_not ; n42064
g41809 and b[41]_not n42064_not ; n42065
g41810 and n41484_not n42006 ; n42066
g41811 and n42002_not n42066 ; n42067
g41812 and n42003_not n42006_not ; n42068
g41813 and n42067_not n42068_not ; n42069
g41814 and n42038_not n42069_not ; n42070
g41815 and n41474_not n42037_not ; n42071
g41816 and n42036_not n42071 ; n42072
g41817 and n42070_not n42072_not ; n42073
g41818 and b[40]_not n42073_not ; n42074
g41819 and n41493_not n42001 ; n42075
g41820 and n41997_not n42075 ; n42076
g41821 and n41998_not n42001_not ; n42077
g41822 and n42076_not n42077_not ; n42078
g41823 and n42038_not n42078_not ; n42079
g41824 and n41483_not n42037_not ; n42080
g41825 and n42036_not n42080 ; n42081
g41826 and n42079_not n42081_not ; n42082
g41827 and b[39]_not n42082_not ; n42083
g41828 and n41502_not n41996 ; n42084
g41829 and n41992_not n42084 ; n42085
g41830 and n41993_not n41996_not ; n42086
g41831 and n42085_not n42086_not ; n42087
g41832 and n42038_not n42087_not ; n42088
g41833 and n41492_not n42037_not ; n42089
g41834 and n42036_not n42089 ; n42090
g41835 and n42088_not n42090_not ; n42091
g41836 and b[38]_not n42091_not ; n42092
g41837 and n41511_not n41991 ; n42093
g41838 and n41987_not n42093 ; n42094
g41839 and n41988_not n41991_not ; n42095
g41840 and n42094_not n42095_not ; n42096
g41841 and n42038_not n42096_not ; n42097
g41842 and n41501_not n42037_not ; n42098
g41843 and n42036_not n42098 ; n42099
g41844 and n42097_not n42099_not ; n42100
g41845 and b[37]_not n42100_not ; n42101
g41846 and n41520_not n41986 ; n42102
g41847 and n41982_not n42102 ; n42103
g41848 and n41983_not n41986_not ; n42104
g41849 and n42103_not n42104_not ; n42105
g41850 and n42038_not n42105_not ; n42106
g41851 and n41510_not n42037_not ; n42107
g41852 and n42036_not n42107 ; n42108
g41853 and n42106_not n42108_not ; n42109
g41854 and b[36]_not n42109_not ; n42110
g41855 and n41529_not n41981 ; n42111
g41856 and n41977_not n42111 ; n42112
g41857 and n41978_not n41981_not ; n42113
g41858 and n42112_not n42113_not ; n42114
g41859 and n42038_not n42114_not ; n42115
g41860 and n41519_not n42037_not ; n42116
g41861 and n42036_not n42116 ; n42117
g41862 and n42115_not n42117_not ; n42118
g41863 and b[35]_not n42118_not ; n42119
g41864 and n41538_not n41976 ; n42120
g41865 and n41972_not n42120 ; n42121
g41866 and n41973_not n41976_not ; n42122
g41867 and n42121_not n42122_not ; n42123
g41868 and n42038_not n42123_not ; n42124
g41869 and n41528_not n42037_not ; n42125
g41870 and n42036_not n42125 ; n42126
g41871 and n42124_not n42126_not ; n42127
g41872 and b[34]_not n42127_not ; n42128
g41873 and n41547_not n41971 ; n42129
g41874 and n41967_not n42129 ; n42130
g41875 and n41968_not n41971_not ; n42131
g41876 and n42130_not n42131_not ; n42132
g41877 and n42038_not n42132_not ; n42133
g41878 and n41537_not n42037_not ; n42134
g41879 and n42036_not n42134 ; n42135
g41880 and n42133_not n42135_not ; n42136
g41881 and b[33]_not n42136_not ; n42137
g41882 and n41556_not n41966 ; n42138
g41883 and n41962_not n42138 ; n42139
g41884 and n41963_not n41966_not ; n42140
g41885 and n42139_not n42140_not ; n42141
g41886 and n42038_not n42141_not ; n42142
g41887 and n41546_not n42037_not ; n42143
g41888 and n42036_not n42143 ; n42144
g41889 and n42142_not n42144_not ; n42145
g41890 and b[32]_not n42145_not ; n42146
g41891 and n41565_not n41961 ; n42147
g41892 and n41957_not n42147 ; n42148
g41893 and n41958_not n41961_not ; n42149
g41894 and n42148_not n42149_not ; n42150
g41895 and n42038_not n42150_not ; n42151
g41896 and n41555_not n42037_not ; n42152
g41897 and n42036_not n42152 ; n42153
g41898 and n42151_not n42153_not ; n42154
g41899 and b[31]_not n42154_not ; n42155
g41900 and n41574_not n41956 ; n42156
g41901 and n41952_not n42156 ; n42157
g41902 and n41953_not n41956_not ; n42158
g41903 and n42157_not n42158_not ; n42159
g41904 and n42038_not n42159_not ; n42160
g41905 and n41564_not n42037_not ; n42161
g41906 and n42036_not n42161 ; n42162
g41907 and n42160_not n42162_not ; n42163
g41908 and b[30]_not n42163_not ; n42164
g41909 and n41583_not n41951 ; n42165
g41910 and n41947_not n42165 ; n42166
g41911 and n41948_not n41951_not ; n42167
g41912 and n42166_not n42167_not ; n42168
g41913 and n42038_not n42168_not ; n42169
g41914 and n41573_not n42037_not ; n42170
g41915 and n42036_not n42170 ; n42171
g41916 and n42169_not n42171_not ; n42172
g41917 and b[29]_not n42172_not ; n42173
g41918 and n41592_not n41946 ; n42174
g41919 and n41942_not n42174 ; n42175
g41920 and n41943_not n41946_not ; n42176
g41921 and n42175_not n42176_not ; n42177
g41922 and n42038_not n42177_not ; n42178
g41923 and n41582_not n42037_not ; n42179
g41924 and n42036_not n42179 ; n42180
g41925 and n42178_not n42180_not ; n42181
g41926 and b[28]_not n42181_not ; n42182
g41927 and n41601_not n41941 ; n42183
g41928 and n41937_not n42183 ; n42184
g41929 and n41938_not n41941_not ; n42185
g41930 and n42184_not n42185_not ; n42186
g41931 and n42038_not n42186_not ; n42187
g41932 and n41591_not n42037_not ; n42188
g41933 and n42036_not n42188 ; n42189
g41934 and n42187_not n42189_not ; n42190
g41935 and b[27]_not n42190_not ; n42191
g41936 and n41610_not n41936 ; n42192
g41937 and n41932_not n42192 ; n42193
g41938 and n41933_not n41936_not ; n42194
g41939 and n42193_not n42194_not ; n42195
g41940 and n42038_not n42195_not ; n42196
g41941 and n41600_not n42037_not ; n42197
g41942 and n42036_not n42197 ; n42198
g41943 and n42196_not n42198_not ; n42199
g41944 and b[26]_not n42199_not ; n42200
g41945 and n41619_not n41931 ; n42201
g41946 and n41927_not n42201 ; n42202
g41947 and n41928_not n41931_not ; n42203
g41948 and n42202_not n42203_not ; n42204
g41949 and n42038_not n42204_not ; n42205
g41950 and n41609_not n42037_not ; n42206
g41951 and n42036_not n42206 ; n42207
g41952 and n42205_not n42207_not ; n42208
g41953 and b[25]_not n42208_not ; n42209
g41954 and n41628_not n41926 ; n42210
g41955 and n41922_not n42210 ; n42211
g41956 and n41923_not n41926_not ; n42212
g41957 and n42211_not n42212_not ; n42213
g41958 and n42038_not n42213_not ; n42214
g41959 and n41618_not n42037_not ; n42215
g41960 and n42036_not n42215 ; n42216
g41961 and n42214_not n42216_not ; n42217
g41962 and b[24]_not n42217_not ; n42218
g41963 and n41637_not n41921 ; n42219
g41964 and n41917_not n42219 ; n42220
g41965 and n41918_not n41921_not ; n42221
g41966 and n42220_not n42221_not ; n42222
g41967 and n42038_not n42222_not ; n42223
g41968 and n41627_not n42037_not ; n42224
g41969 and n42036_not n42224 ; n42225
g41970 and n42223_not n42225_not ; n42226
g41971 and b[23]_not n42226_not ; n42227
g41972 and n41646_not n41916 ; n42228
g41973 and n41912_not n42228 ; n42229
g41974 and n41913_not n41916_not ; n42230
g41975 and n42229_not n42230_not ; n42231
g41976 and n42038_not n42231_not ; n42232
g41977 and n41636_not n42037_not ; n42233
g41978 and n42036_not n42233 ; n42234
g41979 and n42232_not n42234_not ; n42235
g41980 and b[22]_not n42235_not ; n42236
g41981 and n41655_not n41911 ; n42237
g41982 and n41907_not n42237 ; n42238
g41983 and n41908_not n41911_not ; n42239
g41984 and n42238_not n42239_not ; n42240
g41985 and n42038_not n42240_not ; n42241
g41986 and n41645_not n42037_not ; n42242
g41987 and n42036_not n42242 ; n42243
g41988 and n42241_not n42243_not ; n42244
g41989 and b[21]_not n42244_not ; n42245
g41990 and n41664_not n41906 ; n42246
g41991 and n41902_not n42246 ; n42247
g41992 and n41903_not n41906_not ; n42248
g41993 and n42247_not n42248_not ; n42249
g41994 and n42038_not n42249_not ; n42250
g41995 and n41654_not n42037_not ; n42251
g41996 and n42036_not n42251 ; n42252
g41997 and n42250_not n42252_not ; n42253
g41998 and b[20]_not n42253_not ; n42254
g41999 and n41673_not n41901 ; n42255
g42000 and n41897_not n42255 ; n42256
g42001 and n41898_not n41901_not ; n42257
g42002 and n42256_not n42257_not ; n42258
g42003 and n42038_not n42258_not ; n42259
g42004 and n41663_not n42037_not ; n42260
g42005 and n42036_not n42260 ; n42261
g42006 and n42259_not n42261_not ; n42262
g42007 and b[19]_not n42262_not ; n42263
g42008 and n41682_not n41896 ; n42264
g42009 and n41892_not n42264 ; n42265
g42010 and n41893_not n41896_not ; n42266
g42011 and n42265_not n42266_not ; n42267
g42012 and n42038_not n42267_not ; n42268
g42013 and n41672_not n42037_not ; n42269
g42014 and n42036_not n42269 ; n42270
g42015 and n42268_not n42270_not ; n42271
g42016 and b[18]_not n42271_not ; n42272
g42017 and n41691_not n41891 ; n42273
g42018 and n41887_not n42273 ; n42274
g42019 and n41888_not n41891_not ; n42275
g42020 and n42274_not n42275_not ; n42276
g42021 and n42038_not n42276_not ; n42277
g42022 and n41681_not n42037_not ; n42278
g42023 and n42036_not n42278 ; n42279
g42024 and n42277_not n42279_not ; n42280
g42025 and b[17]_not n42280_not ; n42281
g42026 and n41700_not n41886 ; n42282
g42027 and n41882_not n42282 ; n42283
g42028 and n41883_not n41886_not ; n42284
g42029 and n42283_not n42284_not ; n42285
g42030 and n42038_not n42285_not ; n42286
g42031 and n41690_not n42037_not ; n42287
g42032 and n42036_not n42287 ; n42288
g42033 and n42286_not n42288_not ; n42289
g42034 and b[16]_not n42289_not ; n42290
g42035 and n41709_not n41881 ; n42291
g42036 and n41877_not n42291 ; n42292
g42037 and n41878_not n41881_not ; n42293
g42038 and n42292_not n42293_not ; n42294
g42039 and n42038_not n42294_not ; n42295
g42040 and n41699_not n42037_not ; n42296
g42041 and n42036_not n42296 ; n42297
g42042 and n42295_not n42297_not ; n42298
g42043 and b[15]_not n42298_not ; n42299
g42044 and n41718_not n41876 ; n42300
g42045 and n41872_not n42300 ; n42301
g42046 and n41873_not n41876_not ; n42302
g42047 and n42301_not n42302_not ; n42303
g42048 and n42038_not n42303_not ; n42304
g42049 and n41708_not n42037_not ; n42305
g42050 and n42036_not n42305 ; n42306
g42051 and n42304_not n42306_not ; n42307
g42052 and b[14]_not n42307_not ; n42308
g42053 and n41727_not n41871 ; n42309
g42054 and n41867_not n42309 ; n42310
g42055 and n41868_not n41871_not ; n42311
g42056 and n42310_not n42311_not ; n42312
g42057 and n42038_not n42312_not ; n42313
g42058 and n41717_not n42037_not ; n42314
g42059 and n42036_not n42314 ; n42315
g42060 and n42313_not n42315_not ; n42316
g42061 and b[13]_not n42316_not ; n42317
g42062 and n41736_not n41866 ; n42318
g42063 and n41862_not n42318 ; n42319
g42064 and n41863_not n41866_not ; n42320
g42065 and n42319_not n42320_not ; n42321
g42066 and n42038_not n42321_not ; n42322
g42067 and n41726_not n42037_not ; n42323
g42068 and n42036_not n42323 ; n42324
g42069 and n42322_not n42324_not ; n42325
g42070 and b[12]_not n42325_not ; n42326
g42071 and n41745_not n41861 ; n42327
g42072 and n41857_not n42327 ; n42328
g42073 and n41858_not n41861_not ; n42329
g42074 and n42328_not n42329_not ; n42330
g42075 and n42038_not n42330_not ; n42331
g42076 and n41735_not n42037_not ; n42332
g42077 and n42036_not n42332 ; n42333
g42078 and n42331_not n42333_not ; n42334
g42079 and b[11]_not n42334_not ; n42335
g42080 and n41754_not n41856 ; n42336
g42081 and n41852_not n42336 ; n42337
g42082 and n41853_not n41856_not ; n42338
g42083 and n42337_not n42338_not ; n42339
g42084 and n42038_not n42339_not ; n42340
g42085 and n41744_not n42037_not ; n42341
g42086 and n42036_not n42341 ; n42342
g42087 and n42340_not n42342_not ; n42343
g42088 and b[10]_not n42343_not ; n42344
g42089 and n41763_not n41851 ; n42345
g42090 and n41847_not n42345 ; n42346
g42091 and n41848_not n41851_not ; n42347
g42092 and n42346_not n42347_not ; n42348
g42093 and n42038_not n42348_not ; n42349
g42094 and n41753_not n42037_not ; n42350
g42095 and n42036_not n42350 ; n42351
g42096 and n42349_not n42351_not ; n42352
g42097 and b[9]_not n42352_not ; n42353
g42098 and n41772_not n41846 ; n42354
g42099 and n41842_not n42354 ; n42355
g42100 and n41843_not n41846_not ; n42356
g42101 and n42355_not n42356_not ; n42357
g42102 and n42038_not n42357_not ; n42358
g42103 and n41762_not n42037_not ; n42359
g42104 and n42036_not n42359 ; n42360
g42105 and n42358_not n42360_not ; n42361
g42106 and b[8]_not n42361_not ; n42362
g42107 and n41781_not n41841 ; n42363
g42108 and n41837_not n42363 ; n42364
g42109 and n41838_not n41841_not ; n42365
g42110 and n42364_not n42365_not ; n42366
g42111 and n42038_not n42366_not ; n42367
g42112 and n41771_not n42037_not ; n42368
g42113 and n42036_not n42368 ; n42369
g42114 and n42367_not n42369_not ; n42370
g42115 and b[7]_not n42370_not ; n42371
g42116 and n41790_not n41836 ; n42372
g42117 and n41832_not n42372 ; n42373
g42118 and n41833_not n41836_not ; n42374
g42119 and n42373_not n42374_not ; n42375
g42120 and n42038_not n42375_not ; n42376
g42121 and n41780_not n42037_not ; n42377
g42122 and n42036_not n42377 ; n42378
g42123 and n42376_not n42378_not ; n42379
g42124 and b[6]_not n42379_not ; n42380
g42125 and n41799_not n41831 ; n42381
g42126 and n41827_not n42381 ; n42382
g42127 and n41828_not n41831_not ; n42383
g42128 and n42382_not n42383_not ; n42384
g42129 and n42038_not n42384_not ; n42385
g42130 and n41789_not n42037_not ; n42386
g42131 and n42036_not n42386 ; n42387
g42132 and n42385_not n42387_not ; n42388
g42133 and b[5]_not n42388_not ; n42389
g42134 and n41807_not n41826 ; n42390
g42135 and n41822_not n42390 ; n42391
g42136 and n41823_not n41826_not ; n42392
g42137 and n42391_not n42392_not ; n42393
g42138 and n42038_not n42393_not ; n42394
g42139 and n41798_not n42037_not ; n42395
g42140 and n42036_not n42395 ; n42396
g42141 and n42394_not n42396_not ; n42397
g42142 and b[4]_not n42397_not ; n42398
g42143 and n41817_not n41821 ; n42399
g42144 and n41816_not n42399 ; n42400
g42145 and n41818_not n41821_not ; n42401
g42146 and n42400_not n42401_not ; n42402
g42147 and n42038_not n42402_not ; n42403
g42148 and n41806_not n42037_not ; n42404
g42149 and n42036_not n42404 ; n42405
g42150 and n42403_not n42405_not ; n42406
g42151 and b[3]_not n42406_not ; n42407
g42152 and n13739 n41814_not ; n42408
g42153 and n41812_not n42408 ; n42409
g42154 and n41816_not n42409_not ; n42410
g42155 and n42038_not n42410 ; n42411
g42156 and n41811_not n42037_not ; n42412
g42157 and n42036_not n42412 ; n42413
g42158 and n42411_not n42413_not ; n42414
g42159 and b[2]_not n42414_not ; n42415
g42160 and b[0] n42038_not ; n42416
g42161 and a[20] n42416_not ; n42417
g42162 and n13739 n42038_not ; n42418
g42163 and n42417_not n42418_not ; n42419
g42164 and b[1] n42419_not ; n42420
g42165 and b[1]_not n42418_not ; n42421
g42166 and n42417_not n42421 ; n42422
g42167 and n42420_not n42422_not ; n42423
g42168 and n14349_not n42423_not ; n42424
g42169 and b[1]_not n42419_not ; n42425
g42170 and n42424_not n42425_not ; n42426
g42171 and b[2] n42413_not ; n42427
g42172 and n42411_not n42427 ; n42428
g42173 and n42415_not n42428_not ; n42429
g42174 and n42426_not n42429 ; n42430
g42175 and n42415_not n42430_not ; n42431
g42176 and b[3] n42405_not ; n42432
g42177 and n42403_not n42432 ; n42433
g42178 and n42407_not n42433_not ; n42434
g42179 and n42431_not n42434 ; n42435
g42180 and n42407_not n42435_not ; n42436
g42181 and b[4] n42396_not ; n42437
g42182 and n42394_not n42437 ; n42438
g42183 and n42398_not n42438_not ; n42439
g42184 and n42436_not n42439 ; n42440
g42185 and n42398_not n42440_not ; n42441
g42186 and b[5] n42387_not ; n42442
g42187 and n42385_not n42442 ; n42443
g42188 and n42389_not n42443_not ; n42444
g42189 and n42441_not n42444 ; n42445
g42190 and n42389_not n42445_not ; n42446
g42191 and b[6] n42378_not ; n42447
g42192 and n42376_not n42447 ; n42448
g42193 and n42380_not n42448_not ; n42449
g42194 and n42446_not n42449 ; n42450
g42195 and n42380_not n42450_not ; n42451
g42196 and b[7] n42369_not ; n42452
g42197 and n42367_not n42452 ; n42453
g42198 and n42371_not n42453_not ; n42454
g42199 and n42451_not n42454 ; n42455
g42200 and n42371_not n42455_not ; n42456
g42201 and b[8] n42360_not ; n42457
g42202 and n42358_not n42457 ; n42458
g42203 and n42362_not n42458_not ; n42459
g42204 and n42456_not n42459 ; n42460
g42205 and n42362_not n42460_not ; n42461
g42206 and b[9] n42351_not ; n42462
g42207 and n42349_not n42462 ; n42463
g42208 and n42353_not n42463_not ; n42464
g42209 and n42461_not n42464 ; n42465
g42210 and n42353_not n42465_not ; n42466
g42211 and b[10] n42342_not ; n42467
g42212 and n42340_not n42467 ; n42468
g42213 and n42344_not n42468_not ; n42469
g42214 and n42466_not n42469 ; n42470
g42215 and n42344_not n42470_not ; n42471
g42216 and b[11] n42333_not ; n42472
g42217 and n42331_not n42472 ; n42473
g42218 and n42335_not n42473_not ; n42474
g42219 and n42471_not n42474 ; n42475
g42220 and n42335_not n42475_not ; n42476
g42221 and b[12] n42324_not ; n42477
g42222 and n42322_not n42477 ; n42478
g42223 and n42326_not n42478_not ; n42479
g42224 and n42476_not n42479 ; n42480
g42225 and n42326_not n42480_not ; n42481
g42226 and b[13] n42315_not ; n42482
g42227 and n42313_not n42482 ; n42483
g42228 and n42317_not n42483_not ; n42484
g42229 and n42481_not n42484 ; n42485
g42230 and n42317_not n42485_not ; n42486
g42231 and b[14] n42306_not ; n42487
g42232 and n42304_not n42487 ; n42488
g42233 and n42308_not n42488_not ; n42489
g42234 and n42486_not n42489 ; n42490
g42235 and n42308_not n42490_not ; n42491
g42236 and b[15] n42297_not ; n42492
g42237 and n42295_not n42492 ; n42493
g42238 and n42299_not n42493_not ; n42494
g42239 and n42491_not n42494 ; n42495
g42240 and n42299_not n42495_not ; n42496
g42241 and b[16] n42288_not ; n42497
g42242 and n42286_not n42497 ; n42498
g42243 and n42290_not n42498_not ; n42499
g42244 and n42496_not n42499 ; n42500
g42245 and n42290_not n42500_not ; n42501
g42246 and b[17] n42279_not ; n42502
g42247 and n42277_not n42502 ; n42503
g42248 and n42281_not n42503_not ; n42504
g42249 and n42501_not n42504 ; n42505
g42250 and n42281_not n42505_not ; n42506
g42251 and b[18] n42270_not ; n42507
g42252 and n42268_not n42507 ; n42508
g42253 and n42272_not n42508_not ; n42509
g42254 and n42506_not n42509 ; n42510
g42255 and n42272_not n42510_not ; n42511
g42256 and b[19] n42261_not ; n42512
g42257 and n42259_not n42512 ; n42513
g42258 and n42263_not n42513_not ; n42514
g42259 and n42511_not n42514 ; n42515
g42260 and n42263_not n42515_not ; n42516
g42261 and b[20] n42252_not ; n42517
g42262 and n42250_not n42517 ; n42518
g42263 and n42254_not n42518_not ; n42519
g42264 and n42516_not n42519 ; n42520
g42265 and n42254_not n42520_not ; n42521
g42266 and b[21] n42243_not ; n42522
g42267 and n42241_not n42522 ; n42523
g42268 and n42245_not n42523_not ; n42524
g42269 and n42521_not n42524 ; n42525
g42270 and n42245_not n42525_not ; n42526
g42271 and b[22] n42234_not ; n42527
g42272 and n42232_not n42527 ; n42528
g42273 and n42236_not n42528_not ; n42529
g42274 and n42526_not n42529 ; n42530
g42275 and n42236_not n42530_not ; n42531
g42276 and b[23] n42225_not ; n42532
g42277 and n42223_not n42532 ; n42533
g42278 and n42227_not n42533_not ; n42534
g42279 and n42531_not n42534 ; n42535
g42280 and n42227_not n42535_not ; n42536
g42281 and b[24] n42216_not ; n42537
g42282 and n42214_not n42537 ; n42538
g42283 and n42218_not n42538_not ; n42539
g42284 and n42536_not n42539 ; n42540
g42285 and n42218_not n42540_not ; n42541
g42286 and b[25] n42207_not ; n42542
g42287 and n42205_not n42542 ; n42543
g42288 and n42209_not n42543_not ; n42544
g42289 and n42541_not n42544 ; n42545
g42290 and n42209_not n42545_not ; n42546
g42291 and b[26] n42198_not ; n42547
g42292 and n42196_not n42547 ; n42548
g42293 and n42200_not n42548_not ; n42549
g42294 and n42546_not n42549 ; n42550
g42295 and n42200_not n42550_not ; n42551
g42296 and b[27] n42189_not ; n42552
g42297 and n42187_not n42552 ; n42553
g42298 and n42191_not n42553_not ; n42554
g42299 and n42551_not n42554 ; n42555
g42300 and n42191_not n42555_not ; n42556
g42301 and b[28] n42180_not ; n42557
g42302 and n42178_not n42557 ; n42558
g42303 and n42182_not n42558_not ; n42559
g42304 and n42556_not n42559 ; n42560
g42305 and n42182_not n42560_not ; n42561
g42306 and b[29] n42171_not ; n42562
g42307 and n42169_not n42562 ; n42563
g42308 and n42173_not n42563_not ; n42564
g42309 and n42561_not n42564 ; n42565
g42310 and n42173_not n42565_not ; n42566
g42311 and b[30] n42162_not ; n42567
g42312 and n42160_not n42567 ; n42568
g42313 and n42164_not n42568_not ; n42569
g42314 and n42566_not n42569 ; n42570
g42315 and n42164_not n42570_not ; n42571
g42316 and b[31] n42153_not ; n42572
g42317 and n42151_not n42572 ; n42573
g42318 and n42155_not n42573_not ; n42574
g42319 and n42571_not n42574 ; n42575
g42320 and n42155_not n42575_not ; n42576
g42321 and b[32] n42144_not ; n42577
g42322 and n42142_not n42577 ; n42578
g42323 and n42146_not n42578_not ; n42579
g42324 and n42576_not n42579 ; n42580
g42325 and n42146_not n42580_not ; n42581
g42326 and b[33] n42135_not ; n42582
g42327 and n42133_not n42582 ; n42583
g42328 and n42137_not n42583_not ; n42584
g42329 and n42581_not n42584 ; n42585
g42330 and n42137_not n42585_not ; n42586
g42331 and b[34] n42126_not ; n42587
g42332 and n42124_not n42587 ; n42588
g42333 and n42128_not n42588_not ; n42589
g42334 and n42586_not n42589 ; n42590
g42335 and n42128_not n42590_not ; n42591
g42336 and b[35] n42117_not ; n42592
g42337 and n42115_not n42592 ; n42593
g42338 and n42119_not n42593_not ; n42594
g42339 and n42591_not n42594 ; n42595
g42340 and n42119_not n42595_not ; n42596
g42341 and b[36] n42108_not ; n42597
g42342 and n42106_not n42597 ; n42598
g42343 and n42110_not n42598_not ; n42599
g42344 and n42596_not n42599 ; n42600
g42345 and n42110_not n42600_not ; n42601
g42346 and b[37] n42099_not ; n42602
g42347 and n42097_not n42602 ; n42603
g42348 and n42101_not n42603_not ; n42604
g42349 and n42601_not n42604 ; n42605
g42350 and n42101_not n42605_not ; n42606
g42351 and b[38] n42090_not ; n42607
g42352 and n42088_not n42607 ; n42608
g42353 and n42092_not n42608_not ; n42609
g42354 and n42606_not n42609 ; n42610
g42355 and n42092_not n42610_not ; n42611
g42356 and b[39] n42081_not ; n42612
g42357 and n42079_not n42612 ; n42613
g42358 and n42083_not n42613_not ; n42614
g42359 and n42611_not n42614 ; n42615
g42360 and n42083_not n42615_not ; n42616
g42361 and b[40] n42072_not ; n42617
g42362 and n42070_not n42617 ; n42618
g42363 and n42074_not n42618_not ; n42619
g42364 and n42616_not n42619 ; n42620
g42365 and n42074_not n42620_not ; n42621
g42366 and b[41] n42063_not ; n42622
g42367 and n42061_not n42622 ; n42623
g42368 and n42065_not n42623_not ; n42624
g42369 and n42621_not n42624 ; n42625
g42370 and n42065_not n42625_not ; n42626
g42371 and b[42] n42054_not ; n42627
g42372 and n42052_not n42627 ; n42628
g42373 and n42056_not n42628_not ; n42629
g42374 and n42626_not n42629 ; n42630
g42375 and n42056_not n42630_not ; n42631
g42376 and b[43] n42045_not ; n42632
g42377 and n42043_not n42632 ; n42633
g42378 and n42047_not n42633_not ; n42634
g42379 and n42631_not n42634 ; n42635
g42380 and n42047_not n42635_not ; n42636
g42381 and n41448_not n42033_not ; n42637
g42382 and n42031_not n42637 ; n42638
g42383 and n42022_not n42638 ; n42639
g42384 and n42031_not n42033_not ; n42640
g42385 and n42023_not n42640_not ; n42641
g42386 and n42639_not n42641_not ; n42642
g42387 and n42038_not n42642_not ; n42643
g42388 and n42030_not n42037_not ; n42644
g42389 and n42036_not n42644 ; n42645
g42390 and n42643_not n42645_not ; n42646
g42391 and b[44]_not n42646_not ; n42647
g42392 and b[44] n42645_not ; n42648
g42393 and n42643_not n42648 ; n42649
g42394 and n14576 n42649_not ; n42650
g42395 and n42647_not n42650 ; n42651
g42396 and n42636_not n42651 ; n42652
g42397 and n13958 n42646_not ; n42653
g42398 and n42652_not n42653_not ; n42654
g42399 and n42056_not n42634 ; n42655
g42400 and n42630_not n42655 ; n42656
g42401 and n42631_not n42634_not ; n42657
g42402 and n42656_not n42657_not ; n42658
g42403 and n42654_not n42658_not ; n42659
g42404 and n42046_not n42653_not ; n42660
g42405 and n42652_not n42660 ; n42661
g42406 and n42659_not n42661_not ; n42662
g42407 and n42047_not n42649_not ; n42663
g42408 and n42647_not n42663 ; n42664
g42409 and n42635_not n42664 ; n42665
g42410 and n42647_not n42649_not ; n42666
g42411 and n42636_not n42666_not ; n42667
g42412 and n42665_not n42667_not ; n42668
g42413 and n42654_not n42668_not ; n42669
g42414 and n42646_not n42653_not ; n42670
g42415 and n42652_not n42670 ; n42671
g42416 and n42669_not n42671_not ; n42672
g42417 and b[45]_not n42672_not ; n42673
g42418 and b[44]_not n42662_not ; n42674
g42419 and n42065_not n42629 ; n42675
g42420 and n42625_not n42675 ; n42676
g42421 and n42626_not n42629_not ; n42677
g42422 and n42676_not n42677_not ; n42678
g42423 and n42654_not n42678_not ; n42679
g42424 and n42055_not n42653_not ; n42680
g42425 and n42652_not n42680 ; n42681
g42426 and n42679_not n42681_not ; n42682
g42427 and b[43]_not n42682_not ; n42683
g42428 and n42074_not n42624 ; n42684
g42429 and n42620_not n42684 ; n42685
g42430 and n42621_not n42624_not ; n42686
g42431 and n42685_not n42686_not ; n42687
g42432 and n42654_not n42687_not ; n42688
g42433 and n42064_not n42653_not ; n42689
g42434 and n42652_not n42689 ; n42690
g42435 and n42688_not n42690_not ; n42691
g42436 and b[42]_not n42691_not ; n42692
g42437 and n42083_not n42619 ; n42693
g42438 and n42615_not n42693 ; n42694
g42439 and n42616_not n42619_not ; n42695
g42440 and n42694_not n42695_not ; n42696
g42441 and n42654_not n42696_not ; n42697
g42442 and n42073_not n42653_not ; n42698
g42443 and n42652_not n42698 ; n42699
g42444 and n42697_not n42699_not ; n42700
g42445 and b[41]_not n42700_not ; n42701
g42446 and n42092_not n42614 ; n42702
g42447 and n42610_not n42702 ; n42703
g42448 and n42611_not n42614_not ; n42704
g42449 and n42703_not n42704_not ; n42705
g42450 and n42654_not n42705_not ; n42706
g42451 and n42082_not n42653_not ; n42707
g42452 and n42652_not n42707 ; n42708
g42453 and n42706_not n42708_not ; n42709
g42454 and b[40]_not n42709_not ; n42710
g42455 and n42101_not n42609 ; n42711
g42456 and n42605_not n42711 ; n42712
g42457 and n42606_not n42609_not ; n42713
g42458 and n42712_not n42713_not ; n42714
g42459 and n42654_not n42714_not ; n42715
g42460 and n42091_not n42653_not ; n42716
g42461 and n42652_not n42716 ; n42717
g42462 and n42715_not n42717_not ; n42718
g42463 and b[39]_not n42718_not ; n42719
g42464 and n42110_not n42604 ; n42720
g42465 and n42600_not n42720 ; n42721
g42466 and n42601_not n42604_not ; n42722
g42467 and n42721_not n42722_not ; n42723
g42468 and n42654_not n42723_not ; n42724
g42469 and n42100_not n42653_not ; n42725
g42470 and n42652_not n42725 ; n42726
g42471 and n42724_not n42726_not ; n42727
g42472 and b[38]_not n42727_not ; n42728
g42473 and n42119_not n42599 ; n42729
g42474 and n42595_not n42729 ; n42730
g42475 and n42596_not n42599_not ; n42731
g42476 and n42730_not n42731_not ; n42732
g42477 and n42654_not n42732_not ; n42733
g42478 and n42109_not n42653_not ; n42734
g42479 and n42652_not n42734 ; n42735
g42480 and n42733_not n42735_not ; n42736
g42481 and b[37]_not n42736_not ; n42737
g42482 and n42128_not n42594 ; n42738
g42483 and n42590_not n42738 ; n42739
g42484 and n42591_not n42594_not ; n42740
g42485 and n42739_not n42740_not ; n42741
g42486 and n42654_not n42741_not ; n42742
g42487 and n42118_not n42653_not ; n42743
g42488 and n42652_not n42743 ; n42744
g42489 and n42742_not n42744_not ; n42745
g42490 and b[36]_not n42745_not ; n42746
g42491 and n42137_not n42589 ; n42747
g42492 and n42585_not n42747 ; n42748
g42493 and n42586_not n42589_not ; n42749
g42494 and n42748_not n42749_not ; n42750
g42495 and n42654_not n42750_not ; n42751
g42496 and n42127_not n42653_not ; n42752
g42497 and n42652_not n42752 ; n42753
g42498 and n42751_not n42753_not ; n42754
g42499 and b[35]_not n42754_not ; n42755
g42500 and n42146_not n42584 ; n42756
g42501 and n42580_not n42756 ; n42757
g42502 and n42581_not n42584_not ; n42758
g42503 and n42757_not n42758_not ; n42759
g42504 and n42654_not n42759_not ; n42760
g42505 and n42136_not n42653_not ; n42761
g42506 and n42652_not n42761 ; n42762
g42507 and n42760_not n42762_not ; n42763
g42508 and b[34]_not n42763_not ; n42764
g42509 and n42155_not n42579 ; n42765
g42510 and n42575_not n42765 ; n42766
g42511 and n42576_not n42579_not ; n42767
g42512 and n42766_not n42767_not ; n42768
g42513 and n42654_not n42768_not ; n42769
g42514 and n42145_not n42653_not ; n42770
g42515 and n42652_not n42770 ; n42771
g42516 and n42769_not n42771_not ; n42772
g42517 and b[33]_not n42772_not ; n42773
g42518 and n42164_not n42574 ; n42774
g42519 and n42570_not n42774 ; n42775
g42520 and n42571_not n42574_not ; n42776
g42521 and n42775_not n42776_not ; n42777
g42522 and n42654_not n42777_not ; n42778
g42523 and n42154_not n42653_not ; n42779
g42524 and n42652_not n42779 ; n42780
g42525 and n42778_not n42780_not ; n42781
g42526 and b[32]_not n42781_not ; n42782
g42527 and n42173_not n42569 ; n42783
g42528 and n42565_not n42783 ; n42784
g42529 and n42566_not n42569_not ; n42785
g42530 and n42784_not n42785_not ; n42786
g42531 and n42654_not n42786_not ; n42787
g42532 and n42163_not n42653_not ; n42788
g42533 and n42652_not n42788 ; n42789
g42534 and n42787_not n42789_not ; n42790
g42535 and b[31]_not n42790_not ; n42791
g42536 and n42182_not n42564 ; n42792
g42537 and n42560_not n42792 ; n42793
g42538 and n42561_not n42564_not ; n42794
g42539 and n42793_not n42794_not ; n42795
g42540 and n42654_not n42795_not ; n42796
g42541 and n42172_not n42653_not ; n42797
g42542 and n42652_not n42797 ; n42798
g42543 and n42796_not n42798_not ; n42799
g42544 and b[30]_not n42799_not ; n42800
g42545 and n42191_not n42559 ; n42801
g42546 and n42555_not n42801 ; n42802
g42547 and n42556_not n42559_not ; n42803
g42548 and n42802_not n42803_not ; n42804
g42549 and n42654_not n42804_not ; n42805
g42550 and n42181_not n42653_not ; n42806
g42551 and n42652_not n42806 ; n42807
g42552 and n42805_not n42807_not ; n42808
g42553 and b[29]_not n42808_not ; n42809
g42554 and n42200_not n42554 ; n42810
g42555 and n42550_not n42810 ; n42811
g42556 and n42551_not n42554_not ; n42812
g42557 and n42811_not n42812_not ; n42813
g42558 and n42654_not n42813_not ; n42814
g42559 and n42190_not n42653_not ; n42815
g42560 and n42652_not n42815 ; n42816
g42561 and n42814_not n42816_not ; n42817
g42562 and b[28]_not n42817_not ; n42818
g42563 and n42209_not n42549 ; n42819
g42564 and n42545_not n42819 ; n42820
g42565 and n42546_not n42549_not ; n42821
g42566 and n42820_not n42821_not ; n42822
g42567 and n42654_not n42822_not ; n42823
g42568 and n42199_not n42653_not ; n42824
g42569 and n42652_not n42824 ; n42825
g42570 and n42823_not n42825_not ; n42826
g42571 and b[27]_not n42826_not ; n42827
g42572 and n42218_not n42544 ; n42828
g42573 and n42540_not n42828 ; n42829
g42574 and n42541_not n42544_not ; n42830
g42575 and n42829_not n42830_not ; n42831
g42576 and n42654_not n42831_not ; n42832
g42577 and n42208_not n42653_not ; n42833
g42578 and n42652_not n42833 ; n42834
g42579 and n42832_not n42834_not ; n42835
g42580 and b[26]_not n42835_not ; n42836
g42581 and n42227_not n42539 ; n42837
g42582 and n42535_not n42837 ; n42838
g42583 and n42536_not n42539_not ; n42839
g42584 and n42838_not n42839_not ; n42840
g42585 and n42654_not n42840_not ; n42841
g42586 and n42217_not n42653_not ; n42842
g42587 and n42652_not n42842 ; n42843
g42588 and n42841_not n42843_not ; n42844
g42589 and b[25]_not n42844_not ; n42845
g42590 and n42236_not n42534 ; n42846
g42591 and n42530_not n42846 ; n42847
g42592 and n42531_not n42534_not ; n42848
g42593 and n42847_not n42848_not ; n42849
g42594 and n42654_not n42849_not ; n42850
g42595 and n42226_not n42653_not ; n42851
g42596 and n42652_not n42851 ; n42852
g42597 and n42850_not n42852_not ; n42853
g42598 and b[24]_not n42853_not ; n42854
g42599 and n42245_not n42529 ; n42855
g42600 and n42525_not n42855 ; n42856
g42601 and n42526_not n42529_not ; n42857
g42602 and n42856_not n42857_not ; n42858
g42603 and n42654_not n42858_not ; n42859
g42604 and n42235_not n42653_not ; n42860
g42605 and n42652_not n42860 ; n42861
g42606 and n42859_not n42861_not ; n42862
g42607 and b[23]_not n42862_not ; n42863
g42608 and n42254_not n42524 ; n42864
g42609 and n42520_not n42864 ; n42865
g42610 and n42521_not n42524_not ; n42866
g42611 and n42865_not n42866_not ; n42867
g42612 and n42654_not n42867_not ; n42868
g42613 and n42244_not n42653_not ; n42869
g42614 and n42652_not n42869 ; n42870
g42615 and n42868_not n42870_not ; n42871
g42616 and b[22]_not n42871_not ; n42872
g42617 and n42263_not n42519 ; n42873
g42618 and n42515_not n42873 ; n42874
g42619 and n42516_not n42519_not ; n42875
g42620 and n42874_not n42875_not ; n42876
g42621 and n42654_not n42876_not ; n42877
g42622 and n42253_not n42653_not ; n42878
g42623 and n42652_not n42878 ; n42879
g42624 and n42877_not n42879_not ; n42880
g42625 and b[21]_not n42880_not ; n42881
g42626 and n42272_not n42514 ; n42882
g42627 and n42510_not n42882 ; n42883
g42628 and n42511_not n42514_not ; n42884
g42629 and n42883_not n42884_not ; n42885
g42630 and n42654_not n42885_not ; n42886
g42631 and n42262_not n42653_not ; n42887
g42632 and n42652_not n42887 ; n42888
g42633 and n42886_not n42888_not ; n42889
g42634 and b[20]_not n42889_not ; n42890
g42635 and n42281_not n42509 ; n42891
g42636 and n42505_not n42891 ; n42892
g42637 and n42506_not n42509_not ; n42893
g42638 and n42892_not n42893_not ; n42894
g42639 and n42654_not n42894_not ; n42895
g42640 and n42271_not n42653_not ; n42896
g42641 and n42652_not n42896 ; n42897
g42642 and n42895_not n42897_not ; n42898
g42643 and b[19]_not n42898_not ; n42899
g42644 and n42290_not n42504 ; n42900
g42645 and n42500_not n42900 ; n42901
g42646 and n42501_not n42504_not ; n42902
g42647 and n42901_not n42902_not ; n42903
g42648 and n42654_not n42903_not ; n42904
g42649 and n42280_not n42653_not ; n42905
g42650 and n42652_not n42905 ; n42906
g42651 and n42904_not n42906_not ; n42907
g42652 and b[18]_not n42907_not ; n42908
g42653 and n42299_not n42499 ; n42909
g42654 and n42495_not n42909 ; n42910
g42655 and n42496_not n42499_not ; n42911
g42656 and n42910_not n42911_not ; n42912
g42657 and n42654_not n42912_not ; n42913
g42658 and n42289_not n42653_not ; n42914
g42659 and n42652_not n42914 ; n42915
g42660 and n42913_not n42915_not ; n42916
g42661 and b[17]_not n42916_not ; n42917
g42662 and n42308_not n42494 ; n42918
g42663 and n42490_not n42918 ; n42919
g42664 and n42491_not n42494_not ; n42920
g42665 and n42919_not n42920_not ; n42921
g42666 and n42654_not n42921_not ; n42922
g42667 and n42298_not n42653_not ; n42923
g42668 and n42652_not n42923 ; n42924
g42669 and n42922_not n42924_not ; n42925
g42670 and b[16]_not n42925_not ; n42926
g42671 and n42317_not n42489 ; n42927
g42672 and n42485_not n42927 ; n42928
g42673 and n42486_not n42489_not ; n42929
g42674 and n42928_not n42929_not ; n42930
g42675 and n42654_not n42930_not ; n42931
g42676 and n42307_not n42653_not ; n42932
g42677 and n42652_not n42932 ; n42933
g42678 and n42931_not n42933_not ; n42934
g42679 and b[15]_not n42934_not ; n42935
g42680 and n42326_not n42484 ; n42936
g42681 and n42480_not n42936 ; n42937
g42682 and n42481_not n42484_not ; n42938
g42683 and n42937_not n42938_not ; n42939
g42684 and n42654_not n42939_not ; n42940
g42685 and n42316_not n42653_not ; n42941
g42686 and n42652_not n42941 ; n42942
g42687 and n42940_not n42942_not ; n42943
g42688 and b[14]_not n42943_not ; n42944
g42689 and n42335_not n42479 ; n42945
g42690 and n42475_not n42945 ; n42946
g42691 and n42476_not n42479_not ; n42947
g42692 and n42946_not n42947_not ; n42948
g42693 and n42654_not n42948_not ; n42949
g42694 and n42325_not n42653_not ; n42950
g42695 and n42652_not n42950 ; n42951
g42696 and n42949_not n42951_not ; n42952
g42697 and b[13]_not n42952_not ; n42953
g42698 and n42344_not n42474 ; n42954
g42699 and n42470_not n42954 ; n42955
g42700 and n42471_not n42474_not ; n42956
g42701 and n42955_not n42956_not ; n42957
g42702 and n42654_not n42957_not ; n42958
g42703 and n42334_not n42653_not ; n42959
g42704 and n42652_not n42959 ; n42960
g42705 and n42958_not n42960_not ; n42961
g42706 and b[12]_not n42961_not ; n42962
g42707 and n42353_not n42469 ; n42963
g42708 and n42465_not n42963 ; n42964
g42709 and n42466_not n42469_not ; n42965
g42710 and n42964_not n42965_not ; n42966
g42711 and n42654_not n42966_not ; n42967
g42712 and n42343_not n42653_not ; n42968
g42713 and n42652_not n42968 ; n42969
g42714 and n42967_not n42969_not ; n42970
g42715 and b[11]_not n42970_not ; n42971
g42716 and n42362_not n42464 ; n42972
g42717 and n42460_not n42972 ; n42973
g42718 and n42461_not n42464_not ; n42974
g42719 and n42973_not n42974_not ; n42975
g42720 and n42654_not n42975_not ; n42976
g42721 and n42352_not n42653_not ; n42977
g42722 and n42652_not n42977 ; n42978
g42723 and n42976_not n42978_not ; n42979
g42724 and b[10]_not n42979_not ; n42980
g42725 and n42371_not n42459 ; n42981
g42726 and n42455_not n42981 ; n42982
g42727 and n42456_not n42459_not ; n42983
g42728 and n42982_not n42983_not ; n42984
g42729 and n42654_not n42984_not ; n42985
g42730 and n42361_not n42653_not ; n42986
g42731 and n42652_not n42986 ; n42987
g42732 and n42985_not n42987_not ; n42988
g42733 and b[9]_not n42988_not ; n42989
g42734 and n42380_not n42454 ; n42990
g42735 and n42450_not n42990 ; n42991
g42736 and n42451_not n42454_not ; n42992
g42737 and n42991_not n42992_not ; n42993
g42738 and n42654_not n42993_not ; n42994
g42739 and n42370_not n42653_not ; n42995
g42740 and n42652_not n42995 ; n42996
g42741 and n42994_not n42996_not ; n42997
g42742 and b[8]_not n42997_not ; n42998
g42743 and n42389_not n42449 ; n42999
g42744 and n42445_not n42999 ; n43000
g42745 and n42446_not n42449_not ; n43001
g42746 and n43000_not n43001_not ; n43002
g42747 and n42654_not n43002_not ; n43003
g42748 and n42379_not n42653_not ; n43004
g42749 and n42652_not n43004 ; n43005
g42750 and n43003_not n43005_not ; n43006
g42751 and b[7]_not n43006_not ; n43007
g42752 and n42398_not n42444 ; n43008
g42753 and n42440_not n43008 ; n43009
g42754 and n42441_not n42444_not ; n43010
g42755 and n43009_not n43010_not ; n43011
g42756 and n42654_not n43011_not ; n43012
g42757 and n42388_not n42653_not ; n43013
g42758 and n42652_not n43013 ; n43014
g42759 and n43012_not n43014_not ; n43015
g42760 and b[6]_not n43015_not ; n43016
g42761 and n42407_not n42439 ; n43017
g42762 and n42435_not n43017 ; n43018
g42763 and n42436_not n42439_not ; n43019
g42764 and n43018_not n43019_not ; n43020
g42765 and n42654_not n43020_not ; n43021
g42766 and n42397_not n42653_not ; n43022
g42767 and n42652_not n43022 ; n43023
g42768 and n43021_not n43023_not ; n43024
g42769 and b[5]_not n43024_not ; n43025
g42770 and n42415_not n42434 ; n43026
g42771 and n42430_not n43026 ; n43027
g42772 and n42431_not n42434_not ; n43028
g42773 and n43027_not n43028_not ; n43029
g42774 and n42654_not n43029_not ; n43030
g42775 and n42406_not n42653_not ; n43031
g42776 and n42652_not n43031 ; n43032
g42777 and n43030_not n43032_not ; n43033
g42778 and b[4]_not n43033_not ; n43034
g42779 and n42425_not n42429 ; n43035
g42780 and n42424_not n43035 ; n43036
g42781 and n42426_not n42429_not ; n43037
g42782 and n43036_not n43037_not ; n43038
g42783 and n42654_not n43038_not ; n43039
g42784 and n42414_not n42653_not ; n43040
g42785 and n42652_not n43040 ; n43041
g42786 and n43039_not n43041_not ; n43042
g42787 and b[3]_not n43042_not ; n43043
g42788 and n14349 n42422_not ; n43044
g42789 and n42420_not n43044 ; n43045
g42790 and n42424_not n43045_not ; n43046
g42791 and n42654_not n43046 ; n43047
g42792 and n42419_not n42653_not ; n43048
g42793 and n42652_not n43048 ; n43049
g42794 and n43047_not n43049_not ; n43050
g42795 and b[2]_not n43050_not ; n43051
g42796 and b[0] n42654_not ; n43052
g42797 and a[19] n43052_not ; n43053
g42798 and n14349 n42654_not ; n43054
g42799 and n43053_not n43054_not ; n43055
g42800 and b[1] n43055_not ; n43056
g42801 and b[1]_not n43054_not ; n43057
g42802 and n43053_not n43057 ; n43058
g42803 and n43056_not n43058_not ; n43059
g42804 and n14987_not n43059_not ; n43060
g42805 and b[1]_not n43055_not ; n43061
g42806 and n43060_not n43061_not ; n43062
g42807 and b[2] n43049_not ; n43063
g42808 and n43047_not n43063 ; n43064
g42809 and n43051_not n43064_not ; n43065
g42810 and n43062_not n43065 ; n43066
g42811 and n43051_not n43066_not ; n43067
g42812 and b[3] n43041_not ; n43068
g42813 and n43039_not n43068 ; n43069
g42814 and n43043_not n43069_not ; n43070
g42815 and n43067_not n43070 ; n43071
g42816 and n43043_not n43071_not ; n43072
g42817 and b[4] n43032_not ; n43073
g42818 and n43030_not n43073 ; n43074
g42819 and n43034_not n43074_not ; n43075
g42820 and n43072_not n43075 ; n43076
g42821 and n43034_not n43076_not ; n43077
g42822 and b[5] n43023_not ; n43078
g42823 and n43021_not n43078 ; n43079
g42824 and n43025_not n43079_not ; n43080
g42825 and n43077_not n43080 ; n43081
g42826 and n43025_not n43081_not ; n43082
g42827 and b[6] n43014_not ; n43083
g42828 and n43012_not n43083 ; n43084
g42829 and n43016_not n43084_not ; n43085
g42830 and n43082_not n43085 ; n43086
g42831 and n43016_not n43086_not ; n43087
g42832 and b[7] n43005_not ; n43088
g42833 and n43003_not n43088 ; n43089
g42834 and n43007_not n43089_not ; n43090
g42835 and n43087_not n43090 ; n43091
g42836 and n43007_not n43091_not ; n43092
g42837 and b[8] n42996_not ; n43093
g42838 and n42994_not n43093 ; n43094
g42839 and n42998_not n43094_not ; n43095
g42840 and n43092_not n43095 ; n43096
g42841 and n42998_not n43096_not ; n43097
g42842 and b[9] n42987_not ; n43098
g42843 and n42985_not n43098 ; n43099
g42844 and n42989_not n43099_not ; n43100
g42845 and n43097_not n43100 ; n43101
g42846 and n42989_not n43101_not ; n43102
g42847 and b[10] n42978_not ; n43103
g42848 and n42976_not n43103 ; n43104
g42849 and n42980_not n43104_not ; n43105
g42850 and n43102_not n43105 ; n43106
g42851 and n42980_not n43106_not ; n43107
g42852 and b[11] n42969_not ; n43108
g42853 and n42967_not n43108 ; n43109
g42854 and n42971_not n43109_not ; n43110
g42855 and n43107_not n43110 ; n43111
g42856 and n42971_not n43111_not ; n43112
g42857 and b[12] n42960_not ; n43113
g42858 and n42958_not n43113 ; n43114
g42859 and n42962_not n43114_not ; n43115
g42860 and n43112_not n43115 ; n43116
g42861 and n42962_not n43116_not ; n43117
g42862 and b[13] n42951_not ; n43118
g42863 and n42949_not n43118 ; n43119
g42864 and n42953_not n43119_not ; n43120
g42865 and n43117_not n43120 ; n43121
g42866 and n42953_not n43121_not ; n43122
g42867 and b[14] n42942_not ; n43123
g42868 and n42940_not n43123 ; n43124
g42869 and n42944_not n43124_not ; n43125
g42870 and n43122_not n43125 ; n43126
g42871 and n42944_not n43126_not ; n43127
g42872 and b[15] n42933_not ; n43128
g42873 and n42931_not n43128 ; n43129
g42874 and n42935_not n43129_not ; n43130
g42875 and n43127_not n43130 ; n43131
g42876 and n42935_not n43131_not ; n43132
g42877 and b[16] n42924_not ; n43133
g42878 and n42922_not n43133 ; n43134
g42879 and n42926_not n43134_not ; n43135
g42880 and n43132_not n43135 ; n43136
g42881 and n42926_not n43136_not ; n43137
g42882 and b[17] n42915_not ; n43138
g42883 and n42913_not n43138 ; n43139
g42884 and n42917_not n43139_not ; n43140
g42885 and n43137_not n43140 ; n43141
g42886 and n42917_not n43141_not ; n43142
g42887 and b[18] n42906_not ; n43143
g42888 and n42904_not n43143 ; n43144
g42889 and n42908_not n43144_not ; n43145
g42890 and n43142_not n43145 ; n43146
g42891 and n42908_not n43146_not ; n43147
g42892 and b[19] n42897_not ; n43148
g42893 and n42895_not n43148 ; n43149
g42894 and n42899_not n43149_not ; n43150
g42895 and n43147_not n43150 ; n43151
g42896 and n42899_not n43151_not ; n43152
g42897 and b[20] n42888_not ; n43153
g42898 and n42886_not n43153 ; n43154
g42899 and n42890_not n43154_not ; n43155
g42900 and n43152_not n43155 ; n43156
g42901 and n42890_not n43156_not ; n43157
g42902 and b[21] n42879_not ; n43158
g42903 and n42877_not n43158 ; n43159
g42904 and n42881_not n43159_not ; n43160
g42905 and n43157_not n43160 ; n43161
g42906 and n42881_not n43161_not ; n43162
g42907 and b[22] n42870_not ; n43163
g42908 and n42868_not n43163 ; n43164
g42909 and n42872_not n43164_not ; n43165
g42910 and n43162_not n43165 ; n43166
g42911 and n42872_not n43166_not ; n43167
g42912 and b[23] n42861_not ; n43168
g42913 and n42859_not n43168 ; n43169
g42914 and n42863_not n43169_not ; n43170
g42915 and n43167_not n43170 ; n43171
g42916 and n42863_not n43171_not ; n43172
g42917 and b[24] n42852_not ; n43173
g42918 and n42850_not n43173 ; n43174
g42919 and n42854_not n43174_not ; n43175
g42920 and n43172_not n43175 ; n43176
g42921 and n42854_not n43176_not ; n43177
g42922 and b[25] n42843_not ; n43178
g42923 and n42841_not n43178 ; n43179
g42924 and n42845_not n43179_not ; n43180
g42925 and n43177_not n43180 ; n43181
g42926 and n42845_not n43181_not ; n43182
g42927 and b[26] n42834_not ; n43183
g42928 and n42832_not n43183 ; n43184
g42929 and n42836_not n43184_not ; n43185
g42930 and n43182_not n43185 ; n43186
g42931 and n42836_not n43186_not ; n43187
g42932 and b[27] n42825_not ; n43188
g42933 and n42823_not n43188 ; n43189
g42934 and n42827_not n43189_not ; n43190
g42935 and n43187_not n43190 ; n43191
g42936 and n42827_not n43191_not ; n43192
g42937 and b[28] n42816_not ; n43193
g42938 and n42814_not n43193 ; n43194
g42939 and n42818_not n43194_not ; n43195
g42940 and n43192_not n43195 ; n43196
g42941 and n42818_not n43196_not ; n43197
g42942 and b[29] n42807_not ; n43198
g42943 and n42805_not n43198 ; n43199
g42944 and n42809_not n43199_not ; n43200
g42945 and n43197_not n43200 ; n43201
g42946 and n42809_not n43201_not ; n43202
g42947 and b[30] n42798_not ; n43203
g42948 and n42796_not n43203 ; n43204
g42949 and n42800_not n43204_not ; n43205
g42950 and n43202_not n43205 ; n43206
g42951 and n42800_not n43206_not ; n43207
g42952 and b[31] n42789_not ; n43208
g42953 and n42787_not n43208 ; n43209
g42954 and n42791_not n43209_not ; n43210
g42955 and n43207_not n43210 ; n43211
g42956 and n42791_not n43211_not ; n43212
g42957 and b[32] n42780_not ; n43213
g42958 and n42778_not n43213 ; n43214
g42959 and n42782_not n43214_not ; n43215
g42960 and n43212_not n43215 ; n43216
g42961 and n42782_not n43216_not ; n43217
g42962 and b[33] n42771_not ; n43218
g42963 and n42769_not n43218 ; n43219
g42964 and n42773_not n43219_not ; n43220
g42965 and n43217_not n43220 ; n43221
g42966 and n42773_not n43221_not ; n43222
g42967 and b[34] n42762_not ; n43223
g42968 and n42760_not n43223 ; n43224
g42969 and n42764_not n43224_not ; n43225
g42970 and n43222_not n43225 ; n43226
g42971 and n42764_not n43226_not ; n43227
g42972 and b[35] n42753_not ; n43228
g42973 and n42751_not n43228 ; n43229
g42974 and n42755_not n43229_not ; n43230
g42975 and n43227_not n43230 ; n43231
g42976 and n42755_not n43231_not ; n43232
g42977 and b[36] n42744_not ; n43233
g42978 and n42742_not n43233 ; n43234
g42979 and n42746_not n43234_not ; n43235
g42980 and n43232_not n43235 ; n43236
g42981 and n42746_not n43236_not ; n43237
g42982 and b[37] n42735_not ; n43238
g42983 and n42733_not n43238 ; n43239
g42984 and n42737_not n43239_not ; n43240
g42985 and n43237_not n43240 ; n43241
g42986 and n42737_not n43241_not ; n43242
g42987 and b[38] n42726_not ; n43243
g42988 and n42724_not n43243 ; n43244
g42989 and n42728_not n43244_not ; n43245
g42990 and n43242_not n43245 ; n43246
g42991 and n42728_not n43246_not ; n43247
g42992 and b[39] n42717_not ; n43248
g42993 and n42715_not n43248 ; n43249
g42994 and n42719_not n43249_not ; n43250
g42995 and n43247_not n43250 ; n43251
g42996 and n42719_not n43251_not ; n43252
g42997 and b[40] n42708_not ; n43253
g42998 and n42706_not n43253 ; n43254
g42999 and n42710_not n43254_not ; n43255
g43000 and n43252_not n43255 ; n43256
g43001 and n42710_not n43256_not ; n43257
g43002 and b[41] n42699_not ; n43258
g43003 and n42697_not n43258 ; n43259
g43004 and n42701_not n43259_not ; n43260
g43005 and n43257_not n43260 ; n43261
g43006 and n42701_not n43261_not ; n43262
g43007 and b[42] n42690_not ; n43263
g43008 and n42688_not n43263 ; n43264
g43009 and n42692_not n43264_not ; n43265
g43010 and n43262_not n43265 ; n43266
g43011 and n42692_not n43266_not ; n43267
g43012 and b[43] n42681_not ; n43268
g43013 and n42679_not n43268 ; n43269
g43014 and n42683_not n43269_not ; n43270
g43015 and n43267_not n43270 ; n43271
g43016 and n42683_not n43271_not ; n43272
g43017 and b[44] n42661_not ; n43273
g43018 and n42659_not n43273 ; n43274
g43019 and n42674_not n43274_not ; n43275
g43020 and n43272_not n43275 ; n43276
g43021 and n42674_not n43276_not ; n43277
g43022 and b[45] n42671_not ; n43278
g43023 and n42669_not n43278 ; n43279
g43024 and n42673_not n43279_not ; n43280
g43025 and n43277_not n43280 ; n43281
g43026 and n42673_not n43281_not ; n43282
g43027 and n15212 n43282_not ; n43283
g43028 and n42662_not n43283_not ; n43284
g43029 and n42683_not n43275 ; n43285
g43030 and n43271_not n43285 ; n43286
g43031 and n43272_not n43275_not ; n43287
g43032 and n43286_not n43287_not ; n43288
g43033 and n15212 n43288_not ; n43289
g43034 and n43282_not n43289 ; n43290
g43035 and n43284_not n43290_not ; n43291
g43036 and b[45]_not n43291_not ; n43292
g43037 and n42682_not n43283_not ; n43293
g43038 and n42692_not n43270 ; n43294
g43039 and n43266_not n43294 ; n43295
g43040 and n43267_not n43270_not ; n43296
g43041 and n43295_not n43296_not ; n43297
g43042 and n15212 n43297_not ; n43298
g43043 and n43282_not n43298 ; n43299
g43044 and n43293_not n43299_not ; n43300
g43045 and b[44]_not n43300_not ; n43301
g43046 and n42691_not n43283_not ; n43302
g43047 and n42701_not n43265 ; n43303
g43048 and n43261_not n43303 ; n43304
g43049 and n43262_not n43265_not ; n43305
g43050 and n43304_not n43305_not ; n43306
g43051 and n15212 n43306_not ; n43307
g43052 and n43282_not n43307 ; n43308
g43053 and n43302_not n43308_not ; n43309
g43054 and b[43]_not n43309_not ; n43310
g43055 and n42700_not n43283_not ; n43311
g43056 and n42710_not n43260 ; n43312
g43057 and n43256_not n43312 ; n43313
g43058 and n43257_not n43260_not ; n43314
g43059 and n43313_not n43314_not ; n43315
g43060 and n15212 n43315_not ; n43316
g43061 and n43282_not n43316 ; n43317
g43062 and n43311_not n43317_not ; n43318
g43063 and b[42]_not n43318_not ; n43319
g43064 and n42709_not n43283_not ; n43320
g43065 and n42719_not n43255 ; n43321
g43066 and n43251_not n43321 ; n43322
g43067 and n43252_not n43255_not ; n43323
g43068 and n43322_not n43323_not ; n43324
g43069 and n15212 n43324_not ; n43325
g43070 and n43282_not n43325 ; n43326
g43071 and n43320_not n43326_not ; n43327
g43072 and b[41]_not n43327_not ; n43328
g43073 and n42718_not n43283_not ; n43329
g43074 and n42728_not n43250 ; n43330
g43075 and n43246_not n43330 ; n43331
g43076 and n43247_not n43250_not ; n43332
g43077 and n43331_not n43332_not ; n43333
g43078 and n15212 n43333_not ; n43334
g43079 and n43282_not n43334 ; n43335
g43080 and n43329_not n43335_not ; n43336
g43081 and b[40]_not n43336_not ; n43337
g43082 and n42727_not n43283_not ; n43338
g43083 and n42737_not n43245 ; n43339
g43084 and n43241_not n43339 ; n43340
g43085 and n43242_not n43245_not ; n43341
g43086 and n43340_not n43341_not ; n43342
g43087 and n15212 n43342_not ; n43343
g43088 and n43282_not n43343 ; n43344
g43089 and n43338_not n43344_not ; n43345
g43090 and b[39]_not n43345_not ; n43346
g43091 and n42736_not n43283_not ; n43347
g43092 and n42746_not n43240 ; n43348
g43093 and n43236_not n43348 ; n43349
g43094 and n43237_not n43240_not ; n43350
g43095 and n43349_not n43350_not ; n43351
g43096 and n15212 n43351_not ; n43352
g43097 and n43282_not n43352 ; n43353
g43098 and n43347_not n43353_not ; n43354
g43099 and b[38]_not n43354_not ; n43355
g43100 and n42745_not n43283_not ; n43356
g43101 and n42755_not n43235 ; n43357
g43102 and n43231_not n43357 ; n43358
g43103 and n43232_not n43235_not ; n43359
g43104 and n43358_not n43359_not ; n43360
g43105 and n15212 n43360_not ; n43361
g43106 and n43282_not n43361 ; n43362
g43107 and n43356_not n43362_not ; n43363
g43108 and b[37]_not n43363_not ; n43364
g43109 and n42754_not n43283_not ; n43365
g43110 and n42764_not n43230 ; n43366
g43111 and n43226_not n43366 ; n43367
g43112 and n43227_not n43230_not ; n43368
g43113 and n43367_not n43368_not ; n43369
g43114 and n15212 n43369_not ; n43370
g43115 and n43282_not n43370 ; n43371
g43116 and n43365_not n43371_not ; n43372
g43117 and b[36]_not n43372_not ; n43373
g43118 and n42763_not n43283_not ; n43374
g43119 and n42773_not n43225 ; n43375
g43120 and n43221_not n43375 ; n43376
g43121 and n43222_not n43225_not ; n43377
g43122 and n43376_not n43377_not ; n43378
g43123 and n15212 n43378_not ; n43379
g43124 and n43282_not n43379 ; n43380
g43125 and n43374_not n43380_not ; n43381
g43126 and b[35]_not n43381_not ; n43382
g43127 and n42772_not n43283_not ; n43383
g43128 and n42782_not n43220 ; n43384
g43129 and n43216_not n43384 ; n43385
g43130 and n43217_not n43220_not ; n43386
g43131 and n43385_not n43386_not ; n43387
g43132 and n15212 n43387_not ; n43388
g43133 and n43282_not n43388 ; n43389
g43134 and n43383_not n43389_not ; n43390
g43135 and b[34]_not n43390_not ; n43391
g43136 and n42781_not n43283_not ; n43392
g43137 and n42791_not n43215 ; n43393
g43138 and n43211_not n43393 ; n43394
g43139 and n43212_not n43215_not ; n43395
g43140 and n43394_not n43395_not ; n43396
g43141 and n15212 n43396_not ; n43397
g43142 and n43282_not n43397 ; n43398
g43143 and n43392_not n43398_not ; n43399
g43144 and b[33]_not n43399_not ; n43400
g43145 and n42790_not n43283_not ; n43401
g43146 and n42800_not n43210 ; n43402
g43147 and n43206_not n43402 ; n43403
g43148 and n43207_not n43210_not ; n43404
g43149 and n43403_not n43404_not ; n43405
g43150 and n15212 n43405_not ; n43406
g43151 and n43282_not n43406 ; n43407
g43152 and n43401_not n43407_not ; n43408
g43153 and b[32]_not n43408_not ; n43409
g43154 and n42799_not n43283_not ; n43410
g43155 and n42809_not n43205 ; n43411
g43156 and n43201_not n43411 ; n43412
g43157 and n43202_not n43205_not ; n43413
g43158 and n43412_not n43413_not ; n43414
g43159 and n15212 n43414_not ; n43415
g43160 and n43282_not n43415 ; n43416
g43161 and n43410_not n43416_not ; n43417
g43162 and b[31]_not n43417_not ; n43418
g43163 and n42808_not n43283_not ; n43419
g43164 and n42818_not n43200 ; n43420
g43165 and n43196_not n43420 ; n43421
g43166 and n43197_not n43200_not ; n43422
g43167 and n43421_not n43422_not ; n43423
g43168 and n15212 n43423_not ; n43424
g43169 and n43282_not n43424 ; n43425
g43170 and n43419_not n43425_not ; n43426
g43171 and b[30]_not n43426_not ; n43427
g43172 and n42817_not n43283_not ; n43428
g43173 and n42827_not n43195 ; n43429
g43174 and n43191_not n43429 ; n43430
g43175 and n43192_not n43195_not ; n43431
g43176 and n43430_not n43431_not ; n43432
g43177 and n15212 n43432_not ; n43433
g43178 and n43282_not n43433 ; n43434
g43179 and n43428_not n43434_not ; n43435
g43180 and b[29]_not n43435_not ; n43436
g43181 and n42826_not n43283_not ; n43437
g43182 and n42836_not n43190 ; n43438
g43183 and n43186_not n43438 ; n43439
g43184 and n43187_not n43190_not ; n43440
g43185 and n43439_not n43440_not ; n43441
g43186 and n15212 n43441_not ; n43442
g43187 and n43282_not n43442 ; n43443
g43188 and n43437_not n43443_not ; n43444
g43189 and b[28]_not n43444_not ; n43445
g43190 and n42835_not n43283_not ; n43446
g43191 and n42845_not n43185 ; n43447
g43192 and n43181_not n43447 ; n43448
g43193 and n43182_not n43185_not ; n43449
g43194 and n43448_not n43449_not ; n43450
g43195 and n15212 n43450_not ; n43451
g43196 and n43282_not n43451 ; n43452
g43197 and n43446_not n43452_not ; n43453
g43198 and b[27]_not n43453_not ; n43454
g43199 and n42844_not n43283_not ; n43455
g43200 and n42854_not n43180 ; n43456
g43201 and n43176_not n43456 ; n43457
g43202 and n43177_not n43180_not ; n43458
g43203 and n43457_not n43458_not ; n43459
g43204 and n15212 n43459_not ; n43460
g43205 and n43282_not n43460 ; n43461
g43206 and n43455_not n43461_not ; n43462
g43207 and b[26]_not n43462_not ; n43463
g43208 and n42853_not n43283_not ; n43464
g43209 and n42863_not n43175 ; n43465
g43210 and n43171_not n43465 ; n43466
g43211 and n43172_not n43175_not ; n43467
g43212 and n43466_not n43467_not ; n43468
g43213 and n15212 n43468_not ; n43469
g43214 and n43282_not n43469 ; n43470
g43215 and n43464_not n43470_not ; n43471
g43216 and b[25]_not n43471_not ; n43472
g43217 and n42862_not n43283_not ; n43473
g43218 and n42872_not n43170 ; n43474
g43219 and n43166_not n43474 ; n43475
g43220 and n43167_not n43170_not ; n43476
g43221 and n43475_not n43476_not ; n43477
g43222 and n15212 n43477_not ; n43478
g43223 and n43282_not n43478 ; n43479
g43224 and n43473_not n43479_not ; n43480
g43225 and b[24]_not n43480_not ; n43481
g43226 and n42871_not n43283_not ; n43482
g43227 and n42881_not n43165 ; n43483
g43228 and n43161_not n43483 ; n43484
g43229 and n43162_not n43165_not ; n43485
g43230 and n43484_not n43485_not ; n43486
g43231 and n15212 n43486_not ; n43487
g43232 and n43282_not n43487 ; n43488
g43233 and n43482_not n43488_not ; n43489
g43234 and b[23]_not n43489_not ; n43490
g43235 and n42880_not n43283_not ; n43491
g43236 and n42890_not n43160 ; n43492
g43237 and n43156_not n43492 ; n43493
g43238 and n43157_not n43160_not ; n43494
g43239 and n43493_not n43494_not ; n43495
g43240 and n15212 n43495_not ; n43496
g43241 and n43282_not n43496 ; n43497
g43242 and n43491_not n43497_not ; n43498
g43243 and b[22]_not n43498_not ; n43499
g43244 and n42889_not n43283_not ; n43500
g43245 and n42899_not n43155 ; n43501
g43246 and n43151_not n43501 ; n43502
g43247 and n43152_not n43155_not ; n43503
g43248 and n43502_not n43503_not ; n43504
g43249 and n15212 n43504_not ; n43505
g43250 and n43282_not n43505 ; n43506
g43251 and n43500_not n43506_not ; n43507
g43252 and b[21]_not n43507_not ; n43508
g43253 and n42898_not n43283_not ; n43509
g43254 and n42908_not n43150 ; n43510
g43255 and n43146_not n43510 ; n43511
g43256 and n43147_not n43150_not ; n43512
g43257 and n43511_not n43512_not ; n43513
g43258 and n15212 n43513_not ; n43514
g43259 and n43282_not n43514 ; n43515
g43260 and n43509_not n43515_not ; n43516
g43261 and b[20]_not n43516_not ; n43517
g43262 and n42907_not n43283_not ; n43518
g43263 and n42917_not n43145 ; n43519
g43264 and n43141_not n43519 ; n43520
g43265 and n43142_not n43145_not ; n43521
g43266 and n43520_not n43521_not ; n43522
g43267 and n15212 n43522_not ; n43523
g43268 and n43282_not n43523 ; n43524
g43269 and n43518_not n43524_not ; n43525
g43270 and b[19]_not n43525_not ; n43526
g43271 and n42916_not n43283_not ; n43527
g43272 and n42926_not n43140 ; n43528
g43273 and n43136_not n43528 ; n43529
g43274 and n43137_not n43140_not ; n43530
g43275 and n43529_not n43530_not ; n43531
g43276 and n15212 n43531_not ; n43532
g43277 and n43282_not n43532 ; n43533
g43278 and n43527_not n43533_not ; n43534
g43279 and b[18]_not n43534_not ; n43535
g43280 and n42925_not n43283_not ; n43536
g43281 and n42935_not n43135 ; n43537
g43282 and n43131_not n43537 ; n43538
g43283 and n43132_not n43135_not ; n43539
g43284 and n43538_not n43539_not ; n43540
g43285 and n15212 n43540_not ; n43541
g43286 and n43282_not n43541 ; n43542
g43287 and n43536_not n43542_not ; n43543
g43288 and b[17]_not n43543_not ; n43544
g43289 and n42934_not n43283_not ; n43545
g43290 and n42944_not n43130 ; n43546
g43291 and n43126_not n43546 ; n43547
g43292 and n43127_not n43130_not ; n43548
g43293 and n43547_not n43548_not ; n43549
g43294 and n15212 n43549_not ; n43550
g43295 and n43282_not n43550 ; n43551
g43296 and n43545_not n43551_not ; n43552
g43297 and b[16]_not n43552_not ; n43553
g43298 and n42943_not n43283_not ; n43554
g43299 and n42953_not n43125 ; n43555
g43300 and n43121_not n43555 ; n43556
g43301 and n43122_not n43125_not ; n43557
g43302 and n43556_not n43557_not ; n43558
g43303 and n15212 n43558_not ; n43559
g43304 and n43282_not n43559 ; n43560
g43305 and n43554_not n43560_not ; n43561
g43306 and b[15]_not n43561_not ; n43562
g43307 and n42952_not n43283_not ; n43563
g43308 and n42962_not n43120 ; n43564
g43309 and n43116_not n43564 ; n43565
g43310 and n43117_not n43120_not ; n43566
g43311 and n43565_not n43566_not ; n43567
g43312 and n15212 n43567_not ; n43568
g43313 and n43282_not n43568 ; n43569
g43314 and n43563_not n43569_not ; n43570
g43315 and b[14]_not n43570_not ; n43571
g43316 and n42961_not n43283_not ; n43572
g43317 and n42971_not n43115 ; n43573
g43318 and n43111_not n43573 ; n43574
g43319 and n43112_not n43115_not ; n43575
g43320 and n43574_not n43575_not ; n43576
g43321 and n15212 n43576_not ; n43577
g43322 and n43282_not n43577 ; n43578
g43323 and n43572_not n43578_not ; n43579
g43324 and b[13]_not n43579_not ; n43580
g43325 and n42970_not n43283_not ; n43581
g43326 and n42980_not n43110 ; n43582
g43327 and n43106_not n43582 ; n43583
g43328 and n43107_not n43110_not ; n43584
g43329 and n43583_not n43584_not ; n43585
g43330 and n15212 n43585_not ; n43586
g43331 and n43282_not n43586 ; n43587
g43332 and n43581_not n43587_not ; n43588
g43333 and b[12]_not n43588_not ; n43589
g43334 and n42979_not n43283_not ; n43590
g43335 and n42989_not n43105 ; n43591
g43336 and n43101_not n43591 ; n43592
g43337 and n43102_not n43105_not ; n43593
g43338 and n43592_not n43593_not ; n43594
g43339 and n15212 n43594_not ; n43595
g43340 and n43282_not n43595 ; n43596
g43341 and n43590_not n43596_not ; n43597
g43342 and b[11]_not n43597_not ; n43598
g43343 and n42988_not n43283_not ; n43599
g43344 and n42998_not n43100 ; n43600
g43345 and n43096_not n43600 ; n43601
g43346 and n43097_not n43100_not ; n43602
g43347 and n43601_not n43602_not ; n43603
g43348 and n15212 n43603_not ; n43604
g43349 and n43282_not n43604 ; n43605
g43350 and n43599_not n43605_not ; n43606
g43351 and b[10]_not n43606_not ; n43607
g43352 and n42997_not n43283_not ; n43608
g43353 and n43007_not n43095 ; n43609
g43354 and n43091_not n43609 ; n43610
g43355 and n43092_not n43095_not ; n43611
g43356 and n43610_not n43611_not ; n43612
g43357 and n15212 n43612_not ; n43613
g43358 and n43282_not n43613 ; n43614
g43359 and n43608_not n43614_not ; n43615
g43360 and b[9]_not n43615_not ; n43616
g43361 and n43006_not n43283_not ; n43617
g43362 and n43016_not n43090 ; n43618
g43363 and n43086_not n43618 ; n43619
g43364 and n43087_not n43090_not ; n43620
g43365 and n43619_not n43620_not ; n43621
g43366 and n15212 n43621_not ; n43622
g43367 and n43282_not n43622 ; n43623
g43368 and n43617_not n43623_not ; n43624
g43369 and b[8]_not n43624_not ; n43625
g43370 and n43015_not n43283_not ; n43626
g43371 and n43025_not n43085 ; n43627
g43372 and n43081_not n43627 ; n43628
g43373 and n43082_not n43085_not ; n43629
g43374 and n43628_not n43629_not ; n43630
g43375 and n15212 n43630_not ; n43631
g43376 and n43282_not n43631 ; n43632
g43377 and n43626_not n43632_not ; n43633
g43378 and b[7]_not n43633_not ; n43634
g43379 and n43024_not n43283_not ; n43635
g43380 and n43034_not n43080 ; n43636
g43381 and n43076_not n43636 ; n43637
g43382 and n43077_not n43080_not ; n43638
g43383 and n43637_not n43638_not ; n43639
g43384 and n15212 n43639_not ; n43640
g43385 and n43282_not n43640 ; n43641
g43386 and n43635_not n43641_not ; n43642
g43387 and b[6]_not n43642_not ; n43643
g43388 and n43033_not n43283_not ; n43644
g43389 and n43043_not n43075 ; n43645
g43390 and n43071_not n43645 ; n43646
g43391 and n43072_not n43075_not ; n43647
g43392 and n43646_not n43647_not ; n43648
g43393 and n15212 n43648_not ; n43649
g43394 and n43282_not n43649 ; n43650
g43395 and n43644_not n43650_not ; n43651
g43396 and b[5]_not n43651_not ; n43652
g43397 and n43042_not n43283_not ; n43653
g43398 and n43051_not n43070 ; n43654
g43399 and n43066_not n43654 ; n43655
g43400 and n43067_not n43070_not ; n43656
g43401 and n43655_not n43656_not ; n43657
g43402 and n15212 n43657_not ; n43658
g43403 and n43282_not n43658 ; n43659
g43404 and n43653_not n43659_not ; n43660
g43405 and b[4]_not n43660_not ; n43661
g43406 and n43050_not n43283_not ; n43662
g43407 and n43061_not n43065 ; n43663
g43408 and n43060_not n43663 ; n43664
g43409 and n43062_not n43065_not ; n43665
g43410 and n43664_not n43665_not ; n43666
g43411 and n15212 n43666_not ; n43667
g43412 and n43282_not n43667 ; n43668
g43413 and n43662_not n43668_not ; n43669
g43414 and b[3]_not n43669_not ; n43670
g43415 and n43055_not n43283_not ; n43671
g43416 and n14987 n43058_not ; n43672
g43417 and n43056_not n43672 ; n43673
g43418 and n15212 n43673_not ; n43674
g43419 and n43060_not n43674 ; n43675
g43420 and n43282_not n43675 ; n43676
g43421 and n43671_not n43676_not ; n43677
g43422 and b[2]_not n43677_not ; n43678
g43423 and n15612 n43282_not ; n43679
g43424 and a[18] n43679_not ; n43680
g43425 and n15617 n43282_not ; n43681
g43426 and n43680_not n43681_not ; n43682
g43427 and b[1] n43682_not ; n43683
g43428 and b[1]_not n43681_not ; n43684
g43429 and n43680_not n43684 ; n43685
g43430 and n43683_not n43685_not ; n43686
g43431 and n15624_not n43686_not ; n43687
g43432 and b[1]_not n43682_not ; n43688
g43433 and n43687_not n43688_not ; n43689
g43434 and b[2] n43676_not ; n43690
g43435 and n43671_not n43690 ; n43691
g43436 and n43678_not n43691_not ; n43692
g43437 and n43689_not n43692 ; n43693
g43438 and n43678_not n43693_not ; n43694
g43439 and b[3] n43668_not ; n43695
g43440 and n43662_not n43695 ; n43696
g43441 and n43670_not n43696_not ; n43697
g43442 and n43694_not n43697 ; n43698
g43443 and n43670_not n43698_not ; n43699
g43444 and b[4] n43659_not ; n43700
g43445 and n43653_not n43700 ; n43701
g43446 and n43661_not n43701_not ; n43702
g43447 and n43699_not n43702 ; n43703
g43448 and n43661_not n43703_not ; n43704
g43449 and b[5] n43650_not ; n43705
g43450 and n43644_not n43705 ; n43706
g43451 and n43652_not n43706_not ; n43707
g43452 and n43704_not n43707 ; n43708
g43453 and n43652_not n43708_not ; n43709
g43454 and b[6] n43641_not ; n43710
g43455 and n43635_not n43710 ; n43711
g43456 and n43643_not n43711_not ; n43712
g43457 and n43709_not n43712 ; n43713
g43458 and n43643_not n43713_not ; n43714
g43459 and b[7] n43632_not ; n43715
g43460 and n43626_not n43715 ; n43716
g43461 and n43634_not n43716_not ; n43717
g43462 and n43714_not n43717 ; n43718
g43463 and n43634_not n43718_not ; n43719
g43464 and b[8] n43623_not ; n43720
g43465 and n43617_not n43720 ; n43721
g43466 and n43625_not n43721_not ; n43722
g43467 and n43719_not n43722 ; n43723
g43468 and n43625_not n43723_not ; n43724
g43469 and b[9] n43614_not ; n43725
g43470 and n43608_not n43725 ; n43726
g43471 and n43616_not n43726_not ; n43727
g43472 and n43724_not n43727 ; n43728
g43473 and n43616_not n43728_not ; n43729
g43474 and b[10] n43605_not ; n43730
g43475 and n43599_not n43730 ; n43731
g43476 and n43607_not n43731_not ; n43732
g43477 and n43729_not n43732 ; n43733
g43478 and n43607_not n43733_not ; n43734
g43479 and b[11] n43596_not ; n43735
g43480 and n43590_not n43735 ; n43736
g43481 and n43598_not n43736_not ; n43737
g43482 and n43734_not n43737 ; n43738
g43483 and n43598_not n43738_not ; n43739
g43484 and b[12] n43587_not ; n43740
g43485 and n43581_not n43740 ; n43741
g43486 and n43589_not n43741_not ; n43742
g43487 and n43739_not n43742 ; n43743
g43488 and n43589_not n43743_not ; n43744
g43489 and b[13] n43578_not ; n43745
g43490 and n43572_not n43745 ; n43746
g43491 and n43580_not n43746_not ; n43747
g43492 and n43744_not n43747 ; n43748
g43493 and n43580_not n43748_not ; n43749
g43494 and b[14] n43569_not ; n43750
g43495 and n43563_not n43750 ; n43751
g43496 and n43571_not n43751_not ; n43752
g43497 and n43749_not n43752 ; n43753
g43498 and n43571_not n43753_not ; n43754
g43499 and b[15] n43560_not ; n43755
g43500 and n43554_not n43755 ; n43756
g43501 and n43562_not n43756_not ; n43757
g43502 and n43754_not n43757 ; n43758
g43503 and n43562_not n43758_not ; n43759
g43504 and b[16] n43551_not ; n43760
g43505 and n43545_not n43760 ; n43761
g43506 and n43553_not n43761_not ; n43762
g43507 and n43759_not n43762 ; n43763
g43508 and n43553_not n43763_not ; n43764
g43509 and b[17] n43542_not ; n43765
g43510 and n43536_not n43765 ; n43766
g43511 and n43544_not n43766_not ; n43767
g43512 and n43764_not n43767 ; n43768
g43513 and n43544_not n43768_not ; n43769
g43514 and b[18] n43533_not ; n43770
g43515 and n43527_not n43770 ; n43771
g43516 and n43535_not n43771_not ; n43772
g43517 and n43769_not n43772 ; n43773
g43518 and n43535_not n43773_not ; n43774
g43519 and b[19] n43524_not ; n43775
g43520 and n43518_not n43775 ; n43776
g43521 and n43526_not n43776_not ; n43777
g43522 and n43774_not n43777 ; n43778
g43523 and n43526_not n43778_not ; n43779
g43524 and b[20] n43515_not ; n43780
g43525 and n43509_not n43780 ; n43781
g43526 and n43517_not n43781_not ; n43782
g43527 and n43779_not n43782 ; n43783
g43528 and n43517_not n43783_not ; n43784
g43529 and b[21] n43506_not ; n43785
g43530 and n43500_not n43785 ; n43786
g43531 and n43508_not n43786_not ; n43787
g43532 and n43784_not n43787 ; n43788
g43533 and n43508_not n43788_not ; n43789
g43534 and b[22] n43497_not ; n43790
g43535 and n43491_not n43790 ; n43791
g43536 and n43499_not n43791_not ; n43792
g43537 and n43789_not n43792 ; n43793
g43538 and n43499_not n43793_not ; n43794
g43539 and b[23] n43488_not ; n43795
g43540 and n43482_not n43795 ; n43796
g43541 and n43490_not n43796_not ; n43797
g43542 and n43794_not n43797 ; n43798
g43543 and n43490_not n43798_not ; n43799
g43544 and b[24] n43479_not ; n43800
g43545 and n43473_not n43800 ; n43801
g43546 and n43481_not n43801_not ; n43802
g43547 and n43799_not n43802 ; n43803
g43548 and n43481_not n43803_not ; n43804
g43549 and b[25] n43470_not ; n43805
g43550 and n43464_not n43805 ; n43806
g43551 and n43472_not n43806_not ; n43807
g43552 and n43804_not n43807 ; n43808
g43553 and n43472_not n43808_not ; n43809
g43554 and b[26] n43461_not ; n43810
g43555 and n43455_not n43810 ; n43811
g43556 and n43463_not n43811_not ; n43812
g43557 and n43809_not n43812 ; n43813
g43558 and n43463_not n43813_not ; n43814
g43559 and b[27] n43452_not ; n43815
g43560 and n43446_not n43815 ; n43816
g43561 and n43454_not n43816_not ; n43817
g43562 and n43814_not n43817 ; n43818
g43563 and n43454_not n43818_not ; n43819
g43564 and b[28] n43443_not ; n43820
g43565 and n43437_not n43820 ; n43821
g43566 and n43445_not n43821_not ; n43822
g43567 and n43819_not n43822 ; n43823
g43568 and n43445_not n43823_not ; n43824
g43569 and b[29] n43434_not ; n43825
g43570 and n43428_not n43825 ; n43826
g43571 and n43436_not n43826_not ; n43827
g43572 and n43824_not n43827 ; n43828
g43573 and n43436_not n43828_not ; n43829
g43574 and b[30] n43425_not ; n43830
g43575 and n43419_not n43830 ; n43831
g43576 and n43427_not n43831_not ; n43832
g43577 and n43829_not n43832 ; n43833
g43578 and n43427_not n43833_not ; n43834
g43579 and b[31] n43416_not ; n43835
g43580 and n43410_not n43835 ; n43836
g43581 and n43418_not n43836_not ; n43837
g43582 and n43834_not n43837 ; n43838
g43583 and n43418_not n43838_not ; n43839
g43584 and b[32] n43407_not ; n43840
g43585 and n43401_not n43840 ; n43841
g43586 and n43409_not n43841_not ; n43842
g43587 and n43839_not n43842 ; n43843
g43588 and n43409_not n43843_not ; n43844
g43589 and b[33] n43398_not ; n43845
g43590 and n43392_not n43845 ; n43846
g43591 and n43400_not n43846_not ; n43847
g43592 and n43844_not n43847 ; n43848
g43593 and n43400_not n43848_not ; n43849
g43594 and b[34] n43389_not ; n43850
g43595 and n43383_not n43850 ; n43851
g43596 and n43391_not n43851_not ; n43852
g43597 and n43849_not n43852 ; n43853
g43598 and n43391_not n43853_not ; n43854
g43599 and b[35] n43380_not ; n43855
g43600 and n43374_not n43855 ; n43856
g43601 and n43382_not n43856_not ; n43857
g43602 and n43854_not n43857 ; n43858
g43603 and n43382_not n43858_not ; n43859
g43604 and b[36] n43371_not ; n43860
g43605 and n43365_not n43860 ; n43861
g43606 and n43373_not n43861_not ; n43862
g43607 and n43859_not n43862 ; n43863
g43608 and n43373_not n43863_not ; n43864
g43609 and b[37] n43362_not ; n43865
g43610 and n43356_not n43865 ; n43866
g43611 and n43364_not n43866_not ; n43867
g43612 and n43864_not n43867 ; n43868
g43613 and n43364_not n43868_not ; n43869
g43614 and b[38] n43353_not ; n43870
g43615 and n43347_not n43870 ; n43871
g43616 and n43355_not n43871_not ; n43872
g43617 and n43869_not n43872 ; n43873
g43618 and n43355_not n43873_not ; n43874
g43619 and b[39] n43344_not ; n43875
g43620 and n43338_not n43875 ; n43876
g43621 and n43346_not n43876_not ; n43877
g43622 and n43874_not n43877 ; n43878
g43623 and n43346_not n43878_not ; n43879
g43624 and b[40] n43335_not ; n43880
g43625 and n43329_not n43880 ; n43881
g43626 and n43337_not n43881_not ; n43882
g43627 and n43879_not n43882 ; n43883
g43628 and n43337_not n43883_not ; n43884
g43629 and b[41] n43326_not ; n43885
g43630 and n43320_not n43885 ; n43886
g43631 and n43328_not n43886_not ; n43887
g43632 and n43884_not n43887 ; n43888
g43633 and n43328_not n43888_not ; n43889
g43634 and b[42] n43317_not ; n43890
g43635 and n43311_not n43890 ; n43891
g43636 and n43319_not n43891_not ; n43892
g43637 and n43889_not n43892 ; n43893
g43638 and n43319_not n43893_not ; n43894
g43639 and b[43] n43308_not ; n43895
g43640 and n43302_not n43895 ; n43896
g43641 and n43310_not n43896_not ; n43897
g43642 and n43894_not n43897 ; n43898
g43643 and n43310_not n43898_not ; n43899
g43644 and b[44] n43299_not ; n43900
g43645 and n43293_not n43900 ; n43901
g43646 and n43301_not n43901_not ; n43902
g43647 and n43899_not n43902 ; n43903
g43648 and n43301_not n43903_not ; n43904
g43649 and b[45] n43290_not ; n43905
g43650 and n43284_not n43905 ; n43906
g43651 and n43292_not n43906_not ; n43907
g43652 and n43904_not n43907 ; n43908
g43653 and n43292_not n43908_not ; n43909
g43654 and n42672_not n43283_not ; n43910
g43655 and n42674_not n43280 ; n43911
g43656 and n43276_not n43911 ; n43912
g43657 and n43277_not n43280_not ; n43913
g43658 and n43912_not n43913_not ; n43914
g43659 and n43283 n43914_not ; n43915
g43660 and n43910_not n43915_not ; n43916
g43661 and b[46]_not n43916_not ; n43917
g43662 and b[46] n43910_not ; n43918
g43663 and n43915_not n43918 ; n43919
g43664 and n15859 n43919_not ; n43920
g43665 and n43917_not n43920 ; n43921
g43666 and n43909_not n43921 ; n43922
g43667 and n15212 n43916_not ; n43923
g43668 and n43922_not n43923_not ; n43924
g43669 and n43301_not n43907 ; n43925
g43670 and n43903_not n43925 ; n43926
g43671 and n43904_not n43907_not ; n43927
g43672 and n43926_not n43927_not ; n43928
g43673 and n43924_not n43928_not ; n43929
g43674 and n43291_not n43923_not ; n43930
g43675 and n43922_not n43930 ; n43931
g43676 and n43929_not n43931_not ; n43932
g43677 and b[46]_not n43932_not ; n43933
g43678 and n43310_not n43902 ; n43934
g43679 and n43898_not n43934 ; n43935
g43680 and n43899_not n43902_not ; n43936
g43681 and n43935_not n43936_not ; n43937
g43682 and n43924_not n43937_not ; n43938
g43683 and n43300_not n43923_not ; n43939
g43684 and n43922_not n43939 ; n43940
g43685 and n43938_not n43940_not ; n43941
g43686 and b[45]_not n43941_not ; n43942
g43687 and n43319_not n43897 ; n43943
g43688 and n43893_not n43943 ; n43944
g43689 and n43894_not n43897_not ; n43945
g43690 and n43944_not n43945_not ; n43946
g43691 and n43924_not n43946_not ; n43947
g43692 and n43309_not n43923_not ; n43948
g43693 and n43922_not n43948 ; n43949
g43694 and n43947_not n43949_not ; n43950
g43695 and b[44]_not n43950_not ; n43951
g43696 and n43328_not n43892 ; n43952
g43697 and n43888_not n43952 ; n43953
g43698 and n43889_not n43892_not ; n43954
g43699 and n43953_not n43954_not ; n43955
g43700 and n43924_not n43955_not ; n43956
g43701 and n43318_not n43923_not ; n43957
g43702 and n43922_not n43957 ; n43958
g43703 and n43956_not n43958_not ; n43959
g43704 and b[43]_not n43959_not ; n43960
g43705 and n43337_not n43887 ; n43961
g43706 and n43883_not n43961 ; n43962
g43707 and n43884_not n43887_not ; n43963
g43708 and n43962_not n43963_not ; n43964
g43709 and n43924_not n43964_not ; n43965
g43710 and n43327_not n43923_not ; n43966
g43711 and n43922_not n43966 ; n43967
g43712 and n43965_not n43967_not ; n43968
g43713 and b[42]_not n43968_not ; n43969
g43714 and n43346_not n43882 ; n43970
g43715 and n43878_not n43970 ; n43971
g43716 and n43879_not n43882_not ; n43972
g43717 and n43971_not n43972_not ; n43973
g43718 and n43924_not n43973_not ; n43974
g43719 and n43336_not n43923_not ; n43975
g43720 and n43922_not n43975 ; n43976
g43721 and n43974_not n43976_not ; n43977
g43722 and b[41]_not n43977_not ; n43978
g43723 and n43355_not n43877 ; n43979
g43724 and n43873_not n43979 ; n43980
g43725 and n43874_not n43877_not ; n43981
g43726 and n43980_not n43981_not ; n43982
g43727 and n43924_not n43982_not ; n43983
g43728 and n43345_not n43923_not ; n43984
g43729 and n43922_not n43984 ; n43985
g43730 and n43983_not n43985_not ; n43986
g43731 and b[40]_not n43986_not ; n43987
g43732 and n43364_not n43872 ; n43988
g43733 and n43868_not n43988 ; n43989
g43734 and n43869_not n43872_not ; n43990
g43735 and n43989_not n43990_not ; n43991
g43736 and n43924_not n43991_not ; n43992
g43737 and n43354_not n43923_not ; n43993
g43738 and n43922_not n43993 ; n43994
g43739 and n43992_not n43994_not ; n43995
g43740 and b[39]_not n43995_not ; n43996
g43741 and n43373_not n43867 ; n43997
g43742 and n43863_not n43997 ; n43998
g43743 and n43864_not n43867_not ; n43999
g43744 and n43998_not n43999_not ; n44000
g43745 and n43924_not n44000_not ; n44001
g43746 and n43363_not n43923_not ; n44002
g43747 and n43922_not n44002 ; n44003
g43748 and n44001_not n44003_not ; n44004
g43749 and b[38]_not n44004_not ; n44005
g43750 and n43382_not n43862 ; n44006
g43751 and n43858_not n44006 ; n44007
g43752 and n43859_not n43862_not ; n44008
g43753 and n44007_not n44008_not ; n44009
g43754 and n43924_not n44009_not ; n44010
g43755 and n43372_not n43923_not ; n44011
g43756 and n43922_not n44011 ; n44012
g43757 and n44010_not n44012_not ; n44013
g43758 and b[37]_not n44013_not ; n44014
g43759 and n43391_not n43857 ; n44015
g43760 and n43853_not n44015 ; n44016
g43761 and n43854_not n43857_not ; n44017
g43762 and n44016_not n44017_not ; n44018
g43763 and n43924_not n44018_not ; n44019
g43764 and n43381_not n43923_not ; n44020
g43765 and n43922_not n44020 ; n44021
g43766 and n44019_not n44021_not ; n44022
g43767 and b[36]_not n44022_not ; n44023
g43768 and n43400_not n43852 ; n44024
g43769 and n43848_not n44024 ; n44025
g43770 and n43849_not n43852_not ; n44026
g43771 and n44025_not n44026_not ; n44027
g43772 and n43924_not n44027_not ; n44028
g43773 and n43390_not n43923_not ; n44029
g43774 and n43922_not n44029 ; n44030
g43775 and n44028_not n44030_not ; n44031
g43776 and b[35]_not n44031_not ; n44032
g43777 and n43409_not n43847 ; n44033
g43778 and n43843_not n44033 ; n44034
g43779 and n43844_not n43847_not ; n44035
g43780 and n44034_not n44035_not ; n44036
g43781 and n43924_not n44036_not ; n44037
g43782 and n43399_not n43923_not ; n44038
g43783 and n43922_not n44038 ; n44039
g43784 and n44037_not n44039_not ; n44040
g43785 and b[34]_not n44040_not ; n44041
g43786 and n43418_not n43842 ; n44042
g43787 and n43838_not n44042 ; n44043
g43788 and n43839_not n43842_not ; n44044
g43789 and n44043_not n44044_not ; n44045
g43790 and n43924_not n44045_not ; n44046
g43791 and n43408_not n43923_not ; n44047
g43792 and n43922_not n44047 ; n44048
g43793 and n44046_not n44048_not ; n44049
g43794 and b[33]_not n44049_not ; n44050
g43795 and n43427_not n43837 ; n44051
g43796 and n43833_not n44051 ; n44052
g43797 and n43834_not n43837_not ; n44053
g43798 and n44052_not n44053_not ; n44054
g43799 and n43924_not n44054_not ; n44055
g43800 and n43417_not n43923_not ; n44056
g43801 and n43922_not n44056 ; n44057
g43802 and n44055_not n44057_not ; n44058
g43803 and b[32]_not n44058_not ; n44059
g43804 and n43436_not n43832 ; n44060
g43805 and n43828_not n44060 ; n44061
g43806 and n43829_not n43832_not ; n44062
g43807 and n44061_not n44062_not ; n44063
g43808 and n43924_not n44063_not ; n44064
g43809 and n43426_not n43923_not ; n44065
g43810 and n43922_not n44065 ; n44066
g43811 and n44064_not n44066_not ; n44067
g43812 and b[31]_not n44067_not ; n44068
g43813 and n43445_not n43827 ; n44069
g43814 and n43823_not n44069 ; n44070
g43815 and n43824_not n43827_not ; n44071
g43816 and n44070_not n44071_not ; n44072
g43817 and n43924_not n44072_not ; n44073
g43818 and n43435_not n43923_not ; n44074
g43819 and n43922_not n44074 ; n44075
g43820 and n44073_not n44075_not ; n44076
g43821 and b[30]_not n44076_not ; n44077
g43822 and n43454_not n43822 ; n44078
g43823 and n43818_not n44078 ; n44079
g43824 and n43819_not n43822_not ; n44080
g43825 and n44079_not n44080_not ; n44081
g43826 and n43924_not n44081_not ; n44082
g43827 and n43444_not n43923_not ; n44083
g43828 and n43922_not n44083 ; n44084
g43829 and n44082_not n44084_not ; n44085
g43830 and b[29]_not n44085_not ; n44086
g43831 and n43463_not n43817 ; n44087
g43832 and n43813_not n44087 ; n44088
g43833 and n43814_not n43817_not ; n44089
g43834 and n44088_not n44089_not ; n44090
g43835 and n43924_not n44090_not ; n44091
g43836 and n43453_not n43923_not ; n44092
g43837 and n43922_not n44092 ; n44093
g43838 and n44091_not n44093_not ; n44094
g43839 and b[28]_not n44094_not ; n44095
g43840 and n43472_not n43812 ; n44096
g43841 and n43808_not n44096 ; n44097
g43842 and n43809_not n43812_not ; n44098
g43843 and n44097_not n44098_not ; n44099
g43844 and n43924_not n44099_not ; n44100
g43845 and n43462_not n43923_not ; n44101
g43846 and n43922_not n44101 ; n44102
g43847 and n44100_not n44102_not ; n44103
g43848 and b[27]_not n44103_not ; n44104
g43849 and n43481_not n43807 ; n44105
g43850 and n43803_not n44105 ; n44106
g43851 and n43804_not n43807_not ; n44107
g43852 and n44106_not n44107_not ; n44108
g43853 and n43924_not n44108_not ; n44109
g43854 and n43471_not n43923_not ; n44110
g43855 and n43922_not n44110 ; n44111
g43856 and n44109_not n44111_not ; n44112
g43857 and b[26]_not n44112_not ; n44113
g43858 and n43490_not n43802 ; n44114
g43859 and n43798_not n44114 ; n44115
g43860 and n43799_not n43802_not ; n44116
g43861 and n44115_not n44116_not ; n44117
g43862 and n43924_not n44117_not ; n44118
g43863 and n43480_not n43923_not ; n44119
g43864 and n43922_not n44119 ; n44120
g43865 and n44118_not n44120_not ; n44121
g43866 and b[25]_not n44121_not ; n44122
g43867 and n43499_not n43797 ; n44123
g43868 and n43793_not n44123 ; n44124
g43869 and n43794_not n43797_not ; n44125
g43870 and n44124_not n44125_not ; n44126
g43871 and n43924_not n44126_not ; n44127
g43872 and n43489_not n43923_not ; n44128
g43873 and n43922_not n44128 ; n44129
g43874 and n44127_not n44129_not ; n44130
g43875 and b[24]_not n44130_not ; n44131
g43876 and n43508_not n43792 ; n44132
g43877 and n43788_not n44132 ; n44133
g43878 and n43789_not n43792_not ; n44134
g43879 and n44133_not n44134_not ; n44135
g43880 and n43924_not n44135_not ; n44136
g43881 and n43498_not n43923_not ; n44137
g43882 and n43922_not n44137 ; n44138
g43883 and n44136_not n44138_not ; n44139
g43884 and b[23]_not n44139_not ; n44140
g43885 and n43517_not n43787 ; n44141
g43886 and n43783_not n44141 ; n44142
g43887 and n43784_not n43787_not ; n44143
g43888 and n44142_not n44143_not ; n44144
g43889 and n43924_not n44144_not ; n44145
g43890 and n43507_not n43923_not ; n44146
g43891 and n43922_not n44146 ; n44147
g43892 and n44145_not n44147_not ; n44148
g43893 and b[22]_not n44148_not ; n44149
g43894 and n43526_not n43782 ; n44150
g43895 and n43778_not n44150 ; n44151
g43896 and n43779_not n43782_not ; n44152
g43897 and n44151_not n44152_not ; n44153
g43898 and n43924_not n44153_not ; n44154
g43899 and n43516_not n43923_not ; n44155
g43900 and n43922_not n44155 ; n44156
g43901 and n44154_not n44156_not ; n44157
g43902 and b[21]_not n44157_not ; n44158
g43903 and n43535_not n43777 ; n44159
g43904 and n43773_not n44159 ; n44160
g43905 and n43774_not n43777_not ; n44161
g43906 and n44160_not n44161_not ; n44162
g43907 and n43924_not n44162_not ; n44163
g43908 and n43525_not n43923_not ; n44164
g43909 and n43922_not n44164 ; n44165
g43910 and n44163_not n44165_not ; n44166
g43911 and b[20]_not n44166_not ; n44167
g43912 and n43544_not n43772 ; n44168
g43913 and n43768_not n44168 ; n44169
g43914 and n43769_not n43772_not ; n44170
g43915 and n44169_not n44170_not ; n44171
g43916 and n43924_not n44171_not ; n44172
g43917 and n43534_not n43923_not ; n44173
g43918 and n43922_not n44173 ; n44174
g43919 and n44172_not n44174_not ; n44175
g43920 and b[19]_not n44175_not ; n44176
g43921 and n43553_not n43767 ; n44177
g43922 and n43763_not n44177 ; n44178
g43923 and n43764_not n43767_not ; n44179
g43924 and n44178_not n44179_not ; n44180
g43925 and n43924_not n44180_not ; n44181
g43926 and n43543_not n43923_not ; n44182
g43927 and n43922_not n44182 ; n44183
g43928 and n44181_not n44183_not ; n44184
g43929 and b[18]_not n44184_not ; n44185
g43930 and n43562_not n43762 ; n44186
g43931 and n43758_not n44186 ; n44187
g43932 and n43759_not n43762_not ; n44188
g43933 and n44187_not n44188_not ; n44189
g43934 and n43924_not n44189_not ; n44190
g43935 and n43552_not n43923_not ; n44191
g43936 and n43922_not n44191 ; n44192
g43937 and n44190_not n44192_not ; n44193
g43938 and b[17]_not n44193_not ; n44194
g43939 and n43571_not n43757 ; n44195
g43940 and n43753_not n44195 ; n44196
g43941 and n43754_not n43757_not ; n44197
g43942 and n44196_not n44197_not ; n44198
g43943 and n43924_not n44198_not ; n44199
g43944 and n43561_not n43923_not ; n44200
g43945 and n43922_not n44200 ; n44201
g43946 and n44199_not n44201_not ; n44202
g43947 and b[16]_not n44202_not ; n44203
g43948 and n43580_not n43752 ; n44204
g43949 and n43748_not n44204 ; n44205
g43950 and n43749_not n43752_not ; n44206
g43951 and n44205_not n44206_not ; n44207
g43952 and n43924_not n44207_not ; n44208
g43953 and n43570_not n43923_not ; n44209
g43954 and n43922_not n44209 ; n44210
g43955 and n44208_not n44210_not ; n44211
g43956 and b[15]_not n44211_not ; n44212
g43957 and n43589_not n43747 ; n44213
g43958 and n43743_not n44213 ; n44214
g43959 and n43744_not n43747_not ; n44215
g43960 and n44214_not n44215_not ; n44216
g43961 and n43924_not n44216_not ; n44217
g43962 and n43579_not n43923_not ; n44218
g43963 and n43922_not n44218 ; n44219
g43964 and n44217_not n44219_not ; n44220
g43965 and b[14]_not n44220_not ; n44221
g43966 and n43598_not n43742 ; n44222
g43967 and n43738_not n44222 ; n44223
g43968 and n43739_not n43742_not ; n44224
g43969 and n44223_not n44224_not ; n44225
g43970 and n43924_not n44225_not ; n44226
g43971 and n43588_not n43923_not ; n44227
g43972 and n43922_not n44227 ; n44228
g43973 and n44226_not n44228_not ; n44229
g43974 and b[13]_not n44229_not ; n44230
g43975 and n43607_not n43737 ; n44231
g43976 and n43733_not n44231 ; n44232
g43977 and n43734_not n43737_not ; n44233
g43978 and n44232_not n44233_not ; n44234
g43979 and n43924_not n44234_not ; n44235
g43980 and n43597_not n43923_not ; n44236
g43981 and n43922_not n44236 ; n44237
g43982 and n44235_not n44237_not ; n44238
g43983 and b[12]_not n44238_not ; n44239
g43984 and n43616_not n43732 ; n44240
g43985 and n43728_not n44240 ; n44241
g43986 and n43729_not n43732_not ; n44242
g43987 and n44241_not n44242_not ; n44243
g43988 and n43924_not n44243_not ; n44244
g43989 and n43606_not n43923_not ; n44245
g43990 and n43922_not n44245 ; n44246
g43991 and n44244_not n44246_not ; n44247
g43992 and b[11]_not n44247_not ; n44248
g43993 and n43625_not n43727 ; n44249
g43994 and n43723_not n44249 ; n44250
g43995 and n43724_not n43727_not ; n44251
g43996 and n44250_not n44251_not ; n44252
g43997 and n43924_not n44252_not ; n44253
g43998 and n43615_not n43923_not ; n44254
g43999 and n43922_not n44254 ; n44255
g44000 and n44253_not n44255_not ; n44256
g44001 and b[10]_not n44256_not ; n44257
g44002 and n43634_not n43722 ; n44258
g44003 and n43718_not n44258 ; n44259
g44004 and n43719_not n43722_not ; n44260
g44005 and n44259_not n44260_not ; n44261
g44006 and n43924_not n44261_not ; n44262
g44007 and n43624_not n43923_not ; n44263
g44008 and n43922_not n44263 ; n44264
g44009 and n44262_not n44264_not ; n44265
g44010 and b[9]_not n44265_not ; n44266
g44011 and n43643_not n43717 ; n44267
g44012 and n43713_not n44267 ; n44268
g44013 and n43714_not n43717_not ; n44269
g44014 and n44268_not n44269_not ; n44270
g44015 and n43924_not n44270_not ; n44271
g44016 and n43633_not n43923_not ; n44272
g44017 and n43922_not n44272 ; n44273
g44018 and n44271_not n44273_not ; n44274
g44019 and b[8]_not n44274_not ; n44275
g44020 and n43652_not n43712 ; n44276
g44021 and n43708_not n44276 ; n44277
g44022 and n43709_not n43712_not ; n44278
g44023 and n44277_not n44278_not ; n44279
g44024 and n43924_not n44279_not ; n44280
g44025 and n43642_not n43923_not ; n44281
g44026 and n43922_not n44281 ; n44282
g44027 and n44280_not n44282_not ; n44283
g44028 and b[7]_not n44283_not ; n44284
g44029 and n43661_not n43707 ; n44285
g44030 and n43703_not n44285 ; n44286
g44031 and n43704_not n43707_not ; n44287
g44032 and n44286_not n44287_not ; n44288
g44033 and n43924_not n44288_not ; n44289
g44034 and n43651_not n43923_not ; n44290
g44035 and n43922_not n44290 ; n44291
g44036 and n44289_not n44291_not ; n44292
g44037 and b[6]_not n44292_not ; n44293
g44038 and n43670_not n43702 ; n44294
g44039 and n43698_not n44294 ; n44295
g44040 and n43699_not n43702_not ; n44296
g44041 and n44295_not n44296_not ; n44297
g44042 and n43924_not n44297_not ; n44298
g44043 and n43660_not n43923_not ; n44299
g44044 and n43922_not n44299 ; n44300
g44045 and n44298_not n44300_not ; n44301
g44046 and b[5]_not n44301_not ; n44302
g44047 and n43678_not n43697 ; n44303
g44048 and n43693_not n44303 ; n44304
g44049 and n43694_not n43697_not ; n44305
g44050 and n44304_not n44305_not ; n44306
g44051 and n43924_not n44306_not ; n44307
g44052 and n43669_not n43923_not ; n44308
g44053 and n43922_not n44308 ; n44309
g44054 and n44307_not n44309_not ; n44310
g44055 and b[4]_not n44310_not ; n44311
g44056 and n43688_not n43692 ; n44312
g44057 and n43687_not n44312 ; n44313
g44058 and n43689_not n43692_not ; n44314
g44059 and n44313_not n44314_not ; n44315
g44060 and n43924_not n44315_not ; n44316
g44061 and n43677_not n43923_not ; n44317
g44062 and n43922_not n44317 ; n44318
g44063 and n44316_not n44318_not ; n44319
g44064 and b[3]_not n44319_not ; n44320
g44065 and n15624 n43685_not ; n44321
g44066 and n43683_not n44321 ; n44322
g44067 and n43687_not n44322_not ; n44323
g44068 and n43924_not n44323 ; n44324
g44069 and n43682_not n43923_not ; n44325
g44070 and n43922_not n44325 ; n44326
g44071 and n44324_not n44326_not ; n44327
g44072 and b[2]_not n44327_not ; n44328
g44073 and b[0] n43924_not ; n44329
g44074 and a[17] n44329_not ; n44330
g44075 and n15624 n43924_not ; n44331
g44076 and n44330_not n44331_not ; n44332
g44077 and b[1] n44332_not ; n44333
g44078 and b[1]_not n44331_not ; n44334
g44079 and n44330_not n44334 ; n44335
g44080 and n44333_not n44335_not ; n44336
g44081 and n16277_not n44336_not ; n44337
g44082 and b[1]_not n44332_not ; n44338
g44083 and n44337_not n44338_not ; n44339
g44084 and b[2] n44326_not ; n44340
g44085 and n44324_not n44340 ; n44341
g44086 and n44328_not n44341_not ; n44342
g44087 and n44339_not n44342 ; n44343
g44088 and n44328_not n44343_not ; n44344
g44089 and b[3] n44318_not ; n44345
g44090 and n44316_not n44345 ; n44346
g44091 and n44320_not n44346_not ; n44347
g44092 and n44344_not n44347 ; n44348
g44093 and n44320_not n44348_not ; n44349
g44094 and b[4] n44309_not ; n44350
g44095 and n44307_not n44350 ; n44351
g44096 and n44311_not n44351_not ; n44352
g44097 and n44349_not n44352 ; n44353
g44098 and n44311_not n44353_not ; n44354
g44099 and b[5] n44300_not ; n44355
g44100 and n44298_not n44355 ; n44356
g44101 and n44302_not n44356_not ; n44357
g44102 and n44354_not n44357 ; n44358
g44103 and n44302_not n44358_not ; n44359
g44104 and b[6] n44291_not ; n44360
g44105 and n44289_not n44360 ; n44361
g44106 and n44293_not n44361_not ; n44362
g44107 and n44359_not n44362 ; n44363
g44108 and n44293_not n44363_not ; n44364
g44109 and b[7] n44282_not ; n44365
g44110 and n44280_not n44365 ; n44366
g44111 and n44284_not n44366_not ; n44367
g44112 and n44364_not n44367 ; n44368
g44113 and n44284_not n44368_not ; n44369
g44114 and b[8] n44273_not ; n44370
g44115 and n44271_not n44370 ; n44371
g44116 and n44275_not n44371_not ; n44372
g44117 and n44369_not n44372 ; n44373
g44118 and n44275_not n44373_not ; n44374
g44119 and b[9] n44264_not ; n44375
g44120 and n44262_not n44375 ; n44376
g44121 and n44266_not n44376_not ; n44377
g44122 and n44374_not n44377 ; n44378
g44123 and n44266_not n44378_not ; n44379
g44124 and b[10] n44255_not ; n44380
g44125 and n44253_not n44380 ; n44381
g44126 and n44257_not n44381_not ; n44382
g44127 and n44379_not n44382 ; n44383
g44128 and n44257_not n44383_not ; n44384
g44129 and b[11] n44246_not ; n44385
g44130 and n44244_not n44385 ; n44386
g44131 and n44248_not n44386_not ; n44387
g44132 and n44384_not n44387 ; n44388
g44133 and n44248_not n44388_not ; n44389
g44134 and b[12] n44237_not ; n44390
g44135 and n44235_not n44390 ; n44391
g44136 and n44239_not n44391_not ; n44392
g44137 and n44389_not n44392 ; n44393
g44138 and n44239_not n44393_not ; n44394
g44139 and b[13] n44228_not ; n44395
g44140 and n44226_not n44395 ; n44396
g44141 and n44230_not n44396_not ; n44397
g44142 and n44394_not n44397 ; n44398
g44143 and n44230_not n44398_not ; n44399
g44144 and b[14] n44219_not ; n44400
g44145 and n44217_not n44400 ; n44401
g44146 and n44221_not n44401_not ; n44402
g44147 and n44399_not n44402 ; n44403
g44148 and n44221_not n44403_not ; n44404
g44149 and b[15] n44210_not ; n44405
g44150 and n44208_not n44405 ; n44406
g44151 and n44212_not n44406_not ; n44407
g44152 and n44404_not n44407 ; n44408
g44153 and n44212_not n44408_not ; n44409
g44154 and b[16] n44201_not ; n44410
g44155 and n44199_not n44410 ; n44411
g44156 and n44203_not n44411_not ; n44412
g44157 and n44409_not n44412 ; n44413
g44158 and n44203_not n44413_not ; n44414
g44159 and b[17] n44192_not ; n44415
g44160 and n44190_not n44415 ; n44416
g44161 and n44194_not n44416_not ; n44417
g44162 and n44414_not n44417 ; n44418
g44163 and n44194_not n44418_not ; n44419
g44164 and b[18] n44183_not ; n44420
g44165 and n44181_not n44420 ; n44421
g44166 and n44185_not n44421_not ; n44422
g44167 and n44419_not n44422 ; n44423
g44168 and n44185_not n44423_not ; n44424
g44169 and b[19] n44174_not ; n44425
g44170 and n44172_not n44425 ; n44426
g44171 and n44176_not n44426_not ; n44427
g44172 and n44424_not n44427 ; n44428
g44173 and n44176_not n44428_not ; n44429
g44174 and b[20] n44165_not ; n44430
g44175 and n44163_not n44430 ; n44431
g44176 and n44167_not n44431_not ; n44432
g44177 and n44429_not n44432 ; n44433
g44178 and n44167_not n44433_not ; n44434
g44179 and b[21] n44156_not ; n44435
g44180 and n44154_not n44435 ; n44436
g44181 and n44158_not n44436_not ; n44437
g44182 and n44434_not n44437 ; n44438
g44183 and n44158_not n44438_not ; n44439
g44184 and b[22] n44147_not ; n44440
g44185 and n44145_not n44440 ; n44441
g44186 and n44149_not n44441_not ; n44442
g44187 and n44439_not n44442 ; n44443
g44188 and n44149_not n44443_not ; n44444
g44189 and b[23] n44138_not ; n44445
g44190 and n44136_not n44445 ; n44446
g44191 and n44140_not n44446_not ; n44447
g44192 and n44444_not n44447 ; n44448
g44193 and n44140_not n44448_not ; n44449
g44194 and b[24] n44129_not ; n44450
g44195 and n44127_not n44450 ; n44451
g44196 and n44131_not n44451_not ; n44452
g44197 and n44449_not n44452 ; n44453
g44198 and n44131_not n44453_not ; n44454
g44199 and b[25] n44120_not ; n44455
g44200 and n44118_not n44455 ; n44456
g44201 and n44122_not n44456_not ; n44457
g44202 and n44454_not n44457 ; n44458
g44203 and n44122_not n44458_not ; n44459
g44204 and b[26] n44111_not ; n44460
g44205 and n44109_not n44460 ; n44461
g44206 and n44113_not n44461_not ; n44462
g44207 and n44459_not n44462 ; n44463
g44208 and n44113_not n44463_not ; n44464
g44209 and b[27] n44102_not ; n44465
g44210 and n44100_not n44465 ; n44466
g44211 and n44104_not n44466_not ; n44467
g44212 and n44464_not n44467 ; n44468
g44213 and n44104_not n44468_not ; n44469
g44214 and b[28] n44093_not ; n44470
g44215 and n44091_not n44470 ; n44471
g44216 and n44095_not n44471_not ; n44472
g44217 and n44469_not n44472 ; n44473
g44218 and n44095_not n44473_not ; n44474
g44219 and b[29] n44084_not ; n44475
g44220 and n44082_not n44475 ; n44476
g44221 and n44086_not n44476_not ; n44477
g44222 and n44474_not n44477 ; n44478
g44223 and n44086_not n44478_not ; n44479
g44224 and b[30] n44075_not ; n44480
g44225 and n44073_not n44480 ; n44481
g44226 and n44077_not n44481_not ; n44482
g44227 and n44479_not n44482 ; n44483
g44228 and n44077_not n44483_not ; n44484
g44229 and b[31] n44066_not ; n44485
g44230 and n44064_not n44485 ; n44486
g44231 and n44068_not n44486_not ; n44487
g44232 and n44484_not n44487 ; n44488
g44233 and n44068_not n44488_not ; n44489
g44234 and b[32] n44057_not ; n44490
g44235 and n44055_not n44490 ; n44491
g44236 and n44059_not n44491_not ; n44492
g44237 and n44489_not n44492 ; n44493
g44238 and n44059_not n44493_not ; n44494
g44239 and b[33] n44048_not ; n44495
g44240 and n44046_not n44495 ; n44496
g44241 and n44050_not n44496_not ; n44497
g44242 and n44494_not n44497 ; n44498
g44243 and n44050_not n44498_not ; n44499
g44244 and b[34] n44039_not ; n44500
g44245 and n44037_not n44500 ; n44501
g44246 and n44041_not n44501_not ; n44502
g44247 and n44499_not n44502 ; n44503
g44248 and n44041_not n44503_not ; n44504
g44249 and b[35] n44030_not ; n44505
g44250 and n44028_not n44505 ; n44506
g44251 and n44032_not n44506_not ; n44507
g44252 and n44504_not n44507 ; n44508
g44253 and n44032_not n44508_not ; n44509
g44254 and b[36] n44021_not ; n44510
g44255 and n44019_not n44510 ; n44511
g44256 and n44023_not n44511_not ; n44512
g44257 and n44509_not n44512 ; n44513
g44258 and n44023_not n44513_not ; n44514
g44259 and b[37] n44012_not ; n44515
g44260 and n44010_not n44515 ; n44516
g44261 and n44014_not n44516_not ; n44517
g44262 and n44514_not n44517 ; n44518
g44263 and n44014_not n44518_not ; n44519
g44264 and b[38] n44003_not ; n44520
g44265 and n44001_not n44520 ; n44521
g44266 and n44005_not n44521_not ; n44522
g44267 and n44519_not n44522 ; n44523
g44268 and n44005_not n44523_not ; n44524
g44269 and b[39] n43994_not ; n44525
g44270 and n43992_not n44525 ; n44526
g44271 and n43996_not n44526_not ; n44527
g44272 and n44524_not n44527 ; n44528
g44273 and n43996_not n44528_not ; n44529
g44274 and b[40] n43985_not ; n44530
g44275 and n43983_not n44530 ; n44531
g44276 and n43987_not n44531_not ; n44532
g44277 and n44529_not n44532 ; n44533
g44278 and n43987_not n44533_not ; n44534
g44279 and b[41] n43976_not ; n44535
g44280 and n43974_not n44535 ; n44536
g44281 and n43978_not n44536_not ; n44537
g44282 and n44534_not n44537 ; n44538
g44283 and n43978_not n44538_not ; n44539
g44284 and b[42] n43967_not ; n44540
g44285 and n43965_not n44540 ; n44541
g44286 and n43969_not n44541_not ; n44542
g44287 and n44539_not n44542 ; n44543
g44288 and n43969_not n44543_not ; n44544
g44289 and b[43] n43958_not ; n44545
g44290 and n43956_not n44545 ; n44546
g44291 and n43960_not n44546_not ; n44547
g44292 and n44544_not n44547 ; n44548
g44293 and n43960_not n44548_not ; n44549
g44294 and b[44] n43949_not ; n44550
g44295 and n43947_not n44550 ; n44551
g44296 and n43951_not n44551_not ; n44552
g44297 and n44549_not n44552 ; n44553
g44298 and n43951_not n44553_not ; n44554
g44299 and b[45] n43940_not ; n44555
g44300 and n43938_not n44555 ; n44556
g44301 and n43942_not n44556_not ; n44557
g44302 and n44554_not n44557 ; n44558
g44303 and n43942_not n44558_not ; n44559
g44304 and b[46] n43931_not ; n44560
g44305 and n43929_not n44560 ; n44561
g44306 and n43933_not n44561_not ; n44562
g44307 and n44559_not n44562 ; n44563
g44308 and n43933_not n44563_not ; n44564
g44309 and n43292_not n43919_not ; n44565
g44310 and n43917_not n44565 ; n44566
g44311 and n43908_not n44566 ; n44567
g44312 and n43917_not n43919_not ; n44568
g44313 and n43909_not n44568_not ; n44569
g44314 and n44567_not n44569_not ; n44570
g44315 and n43924_not n44570_not ; n44571
g44316 and n43916_not n43923_not ; n44572
g44317 and n43922_not n44572 ; n44573
g44318 and n44571_not n44573_not ; n44574
g44319 and b[47]_not n44574_not ; n44575
g44320 and b[47] n44573_not ; n44576
g44321 and n44571_not n44576 ; n44577
g44322 and n338 n44577_not ; n44578
g44323 and n44575_not n44578 ; n44579
g44324 and n44564_not n44579 ; n44580
g44325 and n15859 n44574_not ; n44581
g44326 and n44580_not n44581_not ; n44582
g44327 and n43942_not n44562 ; n44583
g44328 and n44558_not n44583 ; n44584
g44329 and n44559_not n44562_not ; n44585
g44330 and n44584_not n44585_not ; n44586
g44331 and n44582_not n44586_not ; n44587
g44332 and n43932_not n44581_not ; n44588
g44333 and n44580_not n44588 ; n44589
g44334 and n44587_not n44589_not ; n44590
g44335 and n43933_not n44577_not ; n44591
g44336 and n44575_not n44591 ; n44592
g44337 and n44563_not n44592 ; n44593
g44338 and n44575_not n44577_not ; n44594
g44339 and n44564_not n44594_not ; n44595
g44340 and n44593_not n44595_not ; n44596
g44341 and n44582_not n44596_not ; n44597
g44342 and n44574_not n44581_not ; n44598
g44343 and n44580_not n44598 ; n44599
g44344 and n44597_not n44599_not ; n44600
g44345 and b[48]_not n44600_not ; n44601
g44346 and b[47]_not n44590_not ; n44602
g44347 and n43951_not n44557 ; n44603
g44348 and n44553_not n44603 ; n44604
g44349 and n44554_not n44557_not ; n44605
g44350 and n44604_not n44605_not ; n44606
g44351 and n44582_not n44606_not ; n44607
g44352 and n43941_not n44581_not ; n44608
g44353 and n44580_not n44608 ; n44609
g44354 and n44607_not n44609_not ; n44610
g44355 and b[46]_not n44610_not ; n44611
g44356 and n43960_not n44552 ; n44612
g44357 and n44548_not n44612 ; n44613
g44358 and n44549_not n44552_not ; n44614
g44359 and n44613_not n44614_not ; n44615
g44360 and n44582_not n44615_not ; n44616
g44361 and n43950_not n44581_not ; n44617
g44362 and n44580_not n44617 ; n44618
g44363 and n44616_not n44618_not ; n44619
g44364 and b[45]_not n44619_not ; n44620
g44365 and n43969_not n44547 ; n44621
g44366 and n44543_not n44621 ; n44622
g44367 and n44544_not n44547_not ; n44623
g44368 and n44622_not n44623_not ; n44624
g44369 and n44582_not n44624_not ; n44625
g44370 and n43959_not n44581_not ; n44626
g44371 and n44580_not n44626 ; n44627
g44372 and n44625_not n44627_not ; n44628
g44373 and b[44]_not n44628_not ; n44629
g44374 and n43978_not n44542 ; n44630
g44375 and n44538_not n44630 ; n44631
g44376 and n44539_not n44542_not ; n44632
g44377 and n44631_not n44632_not ; n44633
g44378 and n44582_not n44633_not ; n44634
g44379 and n43968_not n44581_not ; n44635
g44380 and n44580_not n44635 ; n44636
g44381 and n44634_not n44636_not ; n44637
g44382 and b[43]_not n44637_not ; n44638
g44383 and n43987_not n44537 ; n44639
g44384 and n44533_not n44639 ; n44640
g44385 and n44534_not n44537_not ; n44641
g44386 and n44640_not n44641_not ; n44642
g44387 and n44582_not n44642_not ; n44643
g44388 and n43977_not n44581_not ; n44644
g44389 and n44580_not n44644 ; n44645
g44390 and n44643_not n44645_not ; n44646
g44391 and b[42]_not n44646_not ; n44647
g44392 and n43996_not n44532 ; n44648
g44393 and n44528_not n44648 ; n44649
g44394 and n44529_not n44532_not ; n44650
g44395 and n44649_not n44650_not ; n44651
g44396 and n44582_not n44651_not ; n44652
g44397 and n43986_not n44581_not ; n44653
g44398 and n44580_not n44653 ; n44654
g44399 and n44652_not n44654_not ; n44655
g44400 and b[41]_not n44655_not ; n44656
g44401 and n44005_not n44527 ; n44657
g44402 and n44523_not n44657 ; n44658
g44403 and n44524_not n44527_not ; n44659
g44404 and n44658_not n44659_not ; n44660
g44405 and n44582_not n44660_not ; n44661
g44406 and n43995_not n44581_not ; n44662
g44407 and n44580_not n44662 ; n44663
g44408 and n44661_not n44663_not ; n44664
g44409 and b[40]_not n44664_not ; n44665
g44410 and n44014_not n44522 ; n44666
g44411 and n44518_not n44666 ; n44667
g44412 and n44519_not n44522_not ; n44668
g44413 and n44667_not n44668_not ; n44669
g44414 and n44582_not n44669_not ; n44670
g44415 and n44004_not n44581_not ; n44671
g44416 and n44580_not n44671 ; n44672
g44417 and n44670_not n44672_not ; n44673
g44418 and b[39]_not n44673_not ; n44674
g44419 and n44023_not n44517 ; n44675
g44420 and n44513_not n44675 ; n44676
g44421 and n44514_not n44517_not ; n44677
g44422 and n44676_not n44677_not ; n44678
g44423 and n44582_not n44678_not ; n44679
g44424 and n44013_not n44581_not ; n44680
g44425 and n44580_not n44680 ; n44681
g44426 and n44679_not n44681_not ; n44682
g44427 and b[38]_not n44682_not ; n44683
g44428 and n44032_not n44512 ; n44684
g44429 and n44508_not n44684 ; n44685
g44430 and n44509_not n44512_not ; n44686
g44431 and n44685_not n44686_not ; n44687
g44432 and n44582_not n44687_not ; n44688
g44433 and n44022_not n44581_not ; n44689
g44434 and n44580_not n44689 ; n44690
g44435 and n44688_not n44690_not ; n44691
g44436 and b[37]_not n44691_not ; n44692
g44437 and n44041_not n44507 ; n44693
g44438 and n44503_not n44693 ; n44694
g44439 and n44504_not n44507_not ; n44695
g44440 and n44694_not n44695_not ; n44696
g44441 and n44582_not n44696_not ; n44697
g44442 and n44031_not n44581_not ; n44698
g44443 and n44580_not n44698 ; n44699
g44444 and n44697_not n44699_not ; n44700
g44445 and b[36]_not n44700_not ; n44701
g44446 and n44050_not n44502 ; n44702
g44447 and n44498_not n44702 ; n44703
g44448 and n44499_not n44502_not ; n44704
g44449 and n44703_not n44704_not ; n44705
g44450 and n44582_not n44705_not ; n44706
g44451 and n44040_not n44581_not ; n44707
g44452 and n44580_not n44707 ; n44708
g44453 and n44706_not n44708_not ; n44709
g44454 and b[35]_not n44709_not ; n44710
g44455 and n44059_not n44497 ; n44711
g44456 and n44493_not n44711 ; n44712
g44457 and n44494_not n44497_not ; n44713
g44458 and n44712_not n44713_not ; n44714
g44459 and n44582_not n44714_not ; n44715
g44460 and n44049_not n44581_not ; n44716
g44461 and n44580_not n44716 ; n44717
g44462 and n44715_not n44717_not ; n44718
g44463 and b[34]_not n44718_not ; n44719
g44464 and n44068_not n44492 ; n44720
g44465 and n44488_not n44720 ; n44721
g44466 and n44489_not n44492_not ; n44722
g44467 and n44721_not n44722_not ; n44723
g44468 and n44582_not n44723_not ; n44724
g44469 and n44058_not n44581_not ; n44725
g44470 and n44580_not n44725 ; n44726
g44471 and n44724_not n44726_not ; n44727
g44472 and b[33]_not n44727_not ; n44728
g44473 and n44077_not n44487 ; n44729
g44474 and n44483_not n44729 ; n44730
g44475 and n44484_not n44487_not ; n44731
g44476 and n44730_not n44731_not ; n44732
g44477 and n44582_not n44732_not ; n44733
g44478 and n44067_not n44581_not ; n44734
g44479 and n44580_not n44734 ; n44735
g44480 and n44733_not n44735_not ; n44736
g44481 and b[32]_not n44736_not ; n44737
g44482 and n44086_not n44482 ; n44738
g44483 and n44478_not n44738 ; n44739
g44484 and n44479_not n44482_not ; n44740
g44485 and n44739_not n44740_not ; n44741
g44486 and n44582_not n44741_not ; n44742
g44487 and n44076_not n44581_not ; n44743
g44488 and n44580_not n44743 ; n44744
g44489 and n44742_not n44744_not ; n44745
g44490 and b[31]_not n44745_not ; n44746
g44491 and n44095_not n44477 ; n44747
g44492 and n44473_not n44747 ; n44748
g44493 and n44474_not n44477_not ; n44749
g44494 and n44748_not n44749_not ; n44750
g44495 and n44582_not n44750_not ; n44751
g44496 and n44085_not n44581_not ; n44752
g44497 and n44580_not n44752 ; n44753
g44498 and n44751_not n44753_not ; n44754
g44499 and b[30]_not n44754_not ; n44755
g44500 and n44104_not n44472 ; n44756
g44501 and n44468_not n44756 ; n44757
g44502 and n44469_not n44472_not ; n44758
g44503 and n44757_not n44758_not ; n44759
g44504 and n44582_not n44759_not ; n44760
g44505 and n44094_not n44581_not ; n44761
g44506 and n44580_not n44761 ; n44762
g44507 and n44760_not n44762_not ; n44763
g44508 and b[29]_not n44763_not ; n44764
g44509 and n44113_not n44467 ; n44765
g44510 and n44463_not n44765 ; n44766
g44511 and n44464_not n44467_not ; n44767
g44512 and n44766_not n44767_not ; n44768
g44513 and n44582_not n44768_not ; n44769
g44514 and n44103_not n44581_not ; n44770
g44515 and n44580_not n44770 ; n44771
g44516 and n44769_not n44771_not ; n44772
g44517 and b[28]_not n44772_not ; n44773
g44518 and n44122_not n44462 ; n44774
g44519 and n44458_not n44774 ; n44775
g44520 and n44459_not n44462_not ; n44776
g44521 and n44775_not n44776_not ; n44777
g44522 and n44582_not n44777_not ; n44778
g44523 and n44112_not n44581_not ; n44779
g44524 and n44580_not n44779 ; n44780
g44525 and n44778_not n44780_not ; n44781
g44526 and b[27]_not n44781_not ; n44782
g44527 and n44131_not n44457 ; n44783
g44528 and n44453_not n44783 ; n44784
g44529 and n44454_not n44457_not ; n44785
g44530 and n44784_not n44785_not ; n44786
g44531 and n44582_not n44786_not ; n44787
g44532 and n44121_not n44581_not ; n44788
g44533 and n44580_not n44788 ; n44789
g44534 and n44787_not n44789_not ; n44790
g44535 and b[26]_not n44790_not ; n44791
g44536 and n44140_not n44452 ; n44792
g44537 and n44448_not n44792 ; n44793
g44538 and n44449_not n44452_not ; n44794
g44539 and n44793_not n44794_not ; n44795
g44540 and n44582_not n44795_not ; n44796
g44541 and n44130_not n44581_not ; n44797
g44542 and n44580_not n44797 ; n44798
g44543 and n44796_not n44798_not ; n44799
g44544 and b[25]_not n44799_not ; n44800
g44545 and n44149_not n44447 ; n44801
g44546 and n44443_not n44801 ; n44802
g44547 and n44444_not n44447_not ; n44803
g44548 and n44802_not n44803_not ; n44804
g44549 and n44582_not n44804_not ; n44805
g44550 and n44139_not n44581_not ; n44806
g44551 and n44580_not n44806 ; n44807
g44552 and n44805_not n44807_not ; n44808
g44553 and b[24]_not n44808_not ; n44809
g44554 and n44158_not n44442 ; n44810
g44555 and n44438_not n44810 ; n44811
g44556 and n44439_not n44442_not ; n44812
g44557 and n44811_not n44812_not ; n44813
g44558 and n44582_not n44813_not ; n44814
g44559 and n44148_not n44581_not ; n44815
g44560 and n44580_not n44815 ; n44816
g44561 and n44814_not n44816_not ; n44817
g44562 and b[23]_not n44817_not ; n44818
g44563 and n44167_not n44437 ; n44819
g44564 and n44433_not n44819 ; n44820
g44565 and n44434_not n44437_not ; n44821
g44566 and n44820_not n44821_not ; n44822
g44567 and n44582_not n44822_not ; n44823
g44568 and n44157_not n44581_not ; n44824
g44569 and n44580_not n44824 ; n44825
g44570 and n44823_not n44825_not ; n44826
g44571 and b[22]_not n44826_not ; n44827
g44572 and n44176_not n44432 ; n44828
g44573 and n44428_not n44828 ; n44829
g44574 and n44429_not n44432_not ; n44830
g44575 and n44829_not n44830_not ; n44831
g44576 and n44582_not n44831_not ; n44832
g44577 and n44166_not n44581_not ; n44833
g44578 and n44580_not n44833 ; n44834
g44579 and n44832_not n44834_not ; n44835
g44580 and b[21]_not n44835_not ; n44836
g44581 and n44185_not n44427 ; n44837
g44582 and n44423_not n44837 ; n44838
g44583 and n44424_not n44427_not ; n44839
g44584 and n44838_not n44839_not ; n44840
g44585 and n44582_not n44840_not ; n44841
g44586 and n44175_not n44581_not ; n44842
g44587 and n44580_not n44842 ; n44843
g44588 and n44841_not n44843_not ; n44844
g44589 and b[20]_not n44844_not ; n44845
g44590 and n44194_not n44422 ; n44846
g44591 and n44418_not n44846 ; n44847
g44592 and n44419_not n44422_not ; n44848
g44593 and n44847_not n44848_not ; n44849
g44594 and n44582_not n44849_not ; n44850
g44595 and n44184_not n44581_not ; n44851
g44596 and n44580_not n44851 ; n44852
g44597 and n44850_not n44852_not ; n44853
g44598 and b[19]_not n44853_not ; n44854
g44599 and n44203_not n44417 ; n44855
g44600 and n44413_not n44855 ; n44856
g44601 and n44414_not n44417_not ; n44857
g44602 and n44856_not n44857_not ; n44858
g44603 and n44582_not n44858_not ; n44859
g44604 and n44193_not n44581_not ; n44860
g44605 and n44580_not n44860 ; n44861
g44606 and n44859_not n44861_not ; n44862
g44607 and b[18]_not n44862_not ; n44863
g44608 and n44212_not n44412 ; n44864
g44609 and n44408_not n44864 ; n44865
g44610 and n44409_not n44412_not ; n44866
g44611 and n44865_not n44866_not ; n44867
g44612 and n44582_not n44867_not ; n44868
g44613 and n44202_not n44581_not ; n44869
g44614 and n44580_not n44869 ; n44870
g44615 and n44868_not n44870_not ; n44871
g44616 and b[17]_not n44871_not ; n44872
g44617 and n44221_not n44407 ; n44873
g44618 and n44403_not n44873 ; n44874
g44619 and n44404_not n44407_not ; n44875
g44620 and n44874_not n44875_not ; n44876
g44621 and n44582_not n44876_not ; n44877
g44622 and n44211_not n44581_not ; n44878
g44623 and n44580_not n44878 ; n44879
g44624 and n44877_not n44879_not ; n44880
g44625 and b[16]_not n44880_not ; n44881
g44626 and n44230_not n44402 ; n44882
g44627 and n44398_not n44882 ; n44883
g44628 and n44399_not n44402_not ; n44884
g44629 and n44883_not n44884_not ; n44885
g44630 and n44582_not n44885_not ; n44886
g44631 and n44220_not n44581_not ; n44887
g44632 and n44580_not n44887 ; n44888
g44633 and n44886_not n44888_not ; n44889
g44634 and b[15]_not n44889_not ; n44890
g44635 and n44239_not n44397 ; n44891
g44636 and n44393_not n44891 ; n44892
g44637 and n44394_not n44397_not ; n44893
g44638 and n44892_not n44893_not ; n44894
g44639 and n44582_not n44894_not ; n44895
g44640 and n44229_not n44581_not ; n44896
g44641 and n44580_not n44896 ; n44897
g44642 and n44895_not n44897_not ; n44898
g44643 and b[14]_not n44898_not ; n44899
g44644 and n44248_not n44392 ; n44900
g44645 and n44388_not n44900 ; n44901
g44646 and n44389_not n44392_not ; n44902
g44647 and n44901_not n44902_not ; n44903
g44648 and n44582_not n44903_not ; n44904
g44649 and n44238_not n44581_not ; n44905
g44650 and n44580_not n44905 ; n44906
g44651 and n44904_not n44906_not ; n44907
g44652 and b[13]_not n44907_not ; n44908
g44653 and n44257_not n44387 ; n44909
g44654 and n44383_not n44909 ; n44910
g44655 and n44384_not n44387_not ; n44911
g44656 and n44910_not n44911_not ; n44912
g44657 and n44582_not n44912_not ; n44913
g44658 and n44247_not n44581_not ; n44914
g44659 and n44580_not n44914 ; n44915
g44660 and n44913_not n44915_not ; n44916
g44661 and b[12]_not n44916_not ; n44917
g44662 and n44266_not n44382 ; n44918
g44663 and n44378_not n44918 ; n44919
g44664 and n44379_not n44382_not ; n44920
g44665 and n44919_not n44920_not ; n44921
g44666 and n44582_not n44921_not ; n44922
g44667 and n44256_not n44581_not ; n44923
g44668 and n44580_not n44923 ; n44924
g44669 and n44922_not n44924_not ; n44925
g44670 and b[11]_not n44925_not ; n44926
g44671 and n44275_not n44377 ; n44927
g44672 and n44373_not n44927 ; n44928
g44673 and n44374_not n44377_not ; n44929
g44674 and n44928_not n44929_not ; n44930
g44675 and n44582_not n44930_not ; n44931
g44676 and n44265_not n44581_not ; n44932
g44677 and n44580_not n44932 ; n44933
g44678 and n44931_not n44933_not ; n44934
g44679 and b[10]_not n44934_not ; n44935
g44680 and n44284_not n44372 ; n44936
g44681 and n44368_not n44936 ; n44937
g44682 and n44369_not n44372_not ; n44938
g44683 and n44937_not n44938_not ; n44939
g44684 and n44582_not n44939_not ; n44940
g44685 and n44274_not n44581_not ; n44941
g44686 and n44580_not n44941 ; n44942
g44687 and n44940_not n44942_not ; n44943
g44688 and b[9]_not n44943_not ; n44944
g44689 and n44293_not n44367 ; n44945
g44690 and n44363_not n44945 ; n44946
g44691 and n44364_not n44367_not ; n44947
g44692 and n44946_not n44947_not ; n44948
g44693 and n44582_not n44948_not ; n44949
g44694 and n44283_not n44581_not ; n44950
g44695 and n44580_not n44950 ; n44951
g44696 and n44949_not n44951_not ; n44952
g44697 and b[8]_not n44952_not ; n44953
g44698 and n44302_not n44362 ; n44954
g44699 and n44358_not n44954 ; n44955
g44700 and n44359_not n44362_not ; n44956
g44701 and n44955_not n44956_not ; n44957
g44702 and n44582_not n44957_not ; n44958
g44703 and n44292_not n44581_not ; n44959
g44704 and n44580_not n44959 ; n44960
g44705 and n44958_not n44960_not ; n44961
g44706 and b[7]_not n44961_not ; n44962
g44707 and n44311_not n44357 ; n44963
g44708 and n44353_not n44963 ; n44964
g44709 and n44354_not n44357_not ; n44965
g44710 and n44964_not n44965_not ; n44966
g44711 and n44582_not n44966_not ; n44967
g44712 and n44301_not n44581_not ; n44968
g44713 and n44580_not n44968 ; n44969
g44714 and n44967_not n44969_not ; n44970
g44715 and b[6]_not n44970_not ; n44971
g44716 and n44320_not n44352 ; n44972
g44717 and n44348_not n44972 ; n44973
g44718 and n44349_not n44352_not ; n44974
g44719 and n44973_not n44974_not ; n44975
g44720 and n44582_not n44975_not ; n44976
g44721 and n44310_not n44581_not ; n44977
g44722 and n44580_not n44977 ; n44978
g44723 and n44976_not n44978_not ; n44979
g44724 and b[5]_not n44979_not ; n44980
g44725 and n44328_not n44347 ; n44981
g44726 and n44343_not n44981 ; n44982
g44727 and n44344_not n44347_not ; n44983
g44728 and n44982_not n44983_not ; n44984
g44729 and n44582_not n44984_not ; n44985
g44730 and n44319_not n44581_not ; n44986
g44731 and n44580_not n44986 ; n44987
g44732 and n44985_not n44987_not ; n44988
g44733 and b[4]_not n44988_not ; n44989
g44734 and n44338_not n44342 ; n44990
g44735 and n44337_not n44990 ; n44991
g44736 and n44339_not n44342_not ; n44992
g44737 and n44991_not n44992_not ; n44993
g44738 and n44582_not n44993_not ; n44994
g44739 and n44327_not n44581_not ; n44995
g44740 and n44580_not n44995 ; n44996
g44741 and n44994_not n44996_not ; n44997
g44742 and b[3]_not n44997_not ; n44998
g44743 and n16277 n44335_not ; n44999
g44744 and n44333_not n44999 ; n45000
g44745 and n44337_not n45000_not ; n45001
g44746 and n44582_not n45001 ; n45002
g44747 and n44332_not n44581_not ; n45003
g44748 and n44580_not n45003 ; n45004
g44749 and n45002_not n45004_not ; n45005
g44750 and b[2]_not n45005_not ; n45006
g44751 and b[0] n44582_not ; n45007
g44752 and a[16] n45007_not ; n45008
g44753 and n16277 n44582_not ; n45009
g44754 and n45008_not n45009_not ; n45010
g44755 and b[1] n45010_not ; n45011
g44756 and b[1]_not n45009_not ; n45012
g44757 and n45008_not n45012 ; n45013
g44758 and n45011_not n45013_not ; n45014
g44759 and n16956_not n45014_not ; n45015
g44760 and b[1]_not n45010_not ; n45016
g44761 and n45015_not n45016_not ; n45017
g44762 and b[2] n45004_not ; n45018
g44763 and n45002_not n45018 ; n45019
g44764 and n45006_not n45019_not ; n45020
g44765 and n45017_not n45020 ; n45021
g44766 and n45006_not n45021_not ; n45022
g44767 and b[3] n44996_not ; n45023
g44768 and n44994_not n45023 ; n45024
g44769 and n44998_not n45024_not ; n45025
g44770 and n45022_not n45025 ; n45026
g44771 and n44998_not n45026_not ; n45027
g44772 and b[4] n44987_not ; n45028
g44773 and n44985_not n45028 ; n45029
g44774 and n44989_not n45029_not ; n45030
g44775 and n45027_not n45030 ; n45031
g44776 and n44989_not n45031_not ; n45032
g44777 and b[5] n44978_not ; n45033
g44778 and n44976_not n45033 ; n45034
g44779 and n44980_not n45034_not ; n45035
g44780 and n45032_not n45035 ; n45036
g44781 and n44980_not n45036_not ; n45037
g44782 and b[6] n44969_not ; n45038
g44783 and n44967_not n45038 ; n45039
g44784 and n44971_not n45039_not ; n45040
g44785 and n45037_not n45040 ; n45041
g44786 and n44971_not n45041_not ; n45042
g44787 and b[7] n44960_not ; n45043
g44788 and n44958_not n45043 ; n45044
g44789 and n44962_not n45044_not ; n45045
g44790 and n45042_not n45045 ; n45046
g44791 and n44962_not n45046_not ; n45047
g44792 and b[8] n44951_not ; n45048
g44793 and n44949_not n45048 ; n45049
g44794 and n44953_not n45049_not ; n45050
g44795 and n45047_not n45050 ; n45051
g44796 and n44953_not n45051_not ; n45052
g44797 and b[9] n44942_not ; n45053
g44798 and n44940_not n45053 ; n45054
g44799 and n44944_not n45054_not ; n45055
g44800 and n45052_not n45055 ; n45056
g44801 and n44944_not n45056_not ; n45057
g44802 and b[10] n44933_not ; n45058
g44803 and n44931_not n45058 ; n45059
g44804 and n44935_not n45059_not ; n45060
g44805 and n45057_not n45060 ; n45061
g44806 and n44935_not n45061_not ; n45062
g44807 and b[11] n44924_not ; n45063
g44808 and n44922_not n45063 ; n45064
g44809 and n44926_not n45064_not ; n45065
g44810 and n45062_not n45065 ; n45066
g44811 and n44926_not n45066_not ; n45067
g44812 and b[12] n44915_not ; n45068
g44813 and n44913_not n45068 ; n45069
g44814 and n44917_not n45069_not ; n45070
g44815 and n45067_not n45070 ; n45071
g44816 and n44917_not n45071_not ; n45072
g44817 and b[13] n44906_not ; n45073
g44818 and n44904_not n45073 ; n45074
g44819 and n44908_not n45074_not ; n45075
g44820 and n45072_not n45075 ; n45076
g44821 and n44908_not n45076_not ; n45077
g44822 and b[14] n44897_not ; n45078
g44823 and n44895_not n45078 ; n45079
g44824 and n44899_not n45079_not ; n45080
g44825 and n45077_not n45080 ; n45081
g44826 and n44899_not n45081_not ; n45082
g44827 and b[15] n44888_not ; n45083
g44828 and n44886_not n45083 ; n45084
g44829 and n44890_not n45084_not ; n45085
g44830 and n45082_not n45085 ; n45086
g44831 and n44890_not n45086_not ; n45087
g44832 and b[16] n44879_not ; n45088
g44833 and n44877_not n45088 ; n45089
g44834 and n44881_not n45089_not ; n45090
g44835 and n45087_not n45090 ; n45091
g44836 and n44881_not n45091_not ; n45092
g44837 and b[17] n44870_not ; n45093
g44838 and n44868_not n45093 ; n45094
g44839 and n44872_not n45094_not ; n45095
g44840 and n45092_not n45095 ; n45096
g44841 and n44872_not n45096_not ; n45097
g44842 and b[18] n44861_not ; n45098
g44843 and n44859_not n45098 ; n45099
g44844 and n44863_not n45099_not ; n45100
g44845 and n45097_not n45100 ; n45101
g44846 and n44863_not n45101_not ; n45102
g44847 and b[19] n44852_not ; n45103
g44848 and n44850_not n45103 ; n45104
g44849 and n44854_not n45104_not ; n45105
g44850 and n45102_not n45105 ; n45106
g44851 and n44854_not n45106_not ; n45107
g44852 and b[20] n44843_not ; n45108
g44853 and n44841_not n45108 ; n45109
g44854 and n44845_not n45109_not ; n45110
g44855 and n45107_not n45110 ; n45111
g44856 and n44845_not n45111_not ; n45112
g44857 and b[21] n44834_not ; n45113
g44858 and n44832_not n45113 ; n45114
g44859 and n44836_not n45114_not ; n45115
g44860 and n45112_not n45115 ; n45116
g44861 and n44836_not n45116_not ; n45117
g44862 and b[22] n44825_not ; n45118
g44863 and n44823_not n45118 ; n45119
g44864 and n44827_not n45119_not ; n45120
g44865 and n45117_not n45120 ; n45121
g44866 and n44827_not n45121_not ; n45122
g44867 and b[23] n44816_not ; n45123
g44868 and n44814_not n45123 ; n45124
g44869 and n44818_not n45124_not ; n45125
g44870 and n45122_not n45125 ; n45126
g44871 and n44818_not n45126_not ; n45127
g44872 and b[24] n44807_not ; n45128
g44873 and n44805_not n45128 ; n45129
g44874 and n44809_not n45129_not ; n45130
g44875 and n45127_not n45130 ; n45131
g44876 and n44809_not n45131_not ; n45132
g44877 and b[25] n44798_not ; n45133
g44878 and n44796_not n45133 ; n45134
g44879 and n44800_not n45134_not ; n45135
g44880 and n45132_not n45135 ; n45136
g44881 and n44800_not n45136_not ; n45137
g44882 and b[26] n44789_not ; n45138
g44883 and n44787_not n45138 ; n45139
g44884 and n44791_not n45139_not ; n45140
g44885 and n45137_not n45140 ; n45141
g44886 and n44791_not n45141_not ; n45142
g44887 and b[27] n44780_not ; n45143
g44888 and n44778_not n45143 ; n45144
g44889 and n44782_not n45144_not ; n45145
g44890 and n45142_not n45145 ; n45146
g44891 and n44782_not n45146_not ; n45147
g44892 and b[28] n44771_not ; n45148
g44893 and n44769_not n45148 ; n45149
g44894 and n44773_not n45149_not ; n45150
g44895 and n45147_not n45150 ; n45151
g44896 and n44773_not n45151_not ; n45152
g44897 and b[29] n44762_not ; n45153
g44898 and n44760_not n45153 ; n45154
g44899 and n44764_not n45154_not ; n45155
g44900 and n45152_not n45155 ; n45156
g44901 and n44764_not n45156_not ; n45157
g44902 and b[30] n44753_not ; n45158
g44903 and n44751_not n45158 ; n45159
g44904 and n44755_not n45159_not ; n45160
g44905 and n45157_not n45160 ; n45161
g44906 and n44755_not n45161_not ; n45162
g44907 and b[31] n44744_not ; n45163
g44908 and n44742_not n45163 ; n45164
g44909 and n44746_not n45164_not ; n45165
g44910 and n45162_not n45165 ; n45166
g44911 and n44746_not n45166_not ; n45167
g44912 and b[32] n44735_not ; n45168
g44913 and n44733_not n45168 ; n45169
g44914 and n44737_not n45169_not ; n45170
g44915 and n45167_not n45170 ; n45171
g44916 and n44737_not n45171_not ; n45172
g44917 and b[33] n44726_not ; n45173
g44918 and n44724_not n45173 ; n45174
g44919 and n44728_not n45174_not ; n45175
g44920 and n45172_not n45175 ; n45176
g44921 and n44728_not n45176_not ; n45177
g44922 and b[34] n44717_not ; n45178
g44923 and n44715_not n45178 ; n45179
g44924 and n44719_not n45179_not ; n45180
g44925 and n45177_not n45180 ; n45181
g44926 and n44719_not n45181_not ; n45182
g44927 and b[35] n44708_not ; n45183
g44928 and n44706_not n45183 ; n45184
g44929 and n44710_not n45184_not ; n45185
g44930 and n45182_not n45185 ; n45186
g44931 and n44710_not n45186_not ; n45187
g44932 and b[36] n44699_not ; n45188
g44933 and n44697_not n45188 ; n45189
g44934 and n44701_not n45189_not ; n45190
g44935 and n45187_not n45190 ; n45191
g44936 and n44701_not n45191_not ; n45192
g44937 and b[37] n44690_not ; n45193
g44938 and n44688_not n45193 ; n45194
g44939 and n44692_not n45194_not ; n45195
g44940 and n45192_not n45195 ; n45196
g44941 and n44692_not n45196_not ; n45197
g44942 and b[38] n44681_not ; n45198
g44943 and n44679_not n45198 ; n45199
g44944 and n44683_not n45199_not ; n45200
g44945 and n45197_not n45200 ; n45201
g44946 and n44683_not n45201_not ; n45202
g44947 and b[39] n44672_not ; n45203
g44948 and n44670_not n45203 ; n45204
g44949 and n44674_not n45204_not ; n45205
g44950 and n45202_not n45205 ; n45206
g44951 and n44674_not n45206_not ; n45207
g44952 and b[40] n44663_not ; n45208
g44953 and n44661_not n45208 ; n45209
g44954 and n44665_not n45209_not ; n45210
g44955 and n45207_not n45210 ; n45211
g44956 and n44665_not n45211_not ; n45212
g44957 and b[41] n44654_not ; n45213
g44958 and n44652_not n45213 ; n45214
g44959 and n44656_not n45214_not ; n45215
g44960 and n45212_not n45215 ; n45216
g44961 and n44656_not n45216_not ; n45217
g44962 and b[42] n44645_not ; n45218
g44963 and n44643_not n45218 ; n45219
g44964 and n44647_not n45219_not ; n45220
g44965 and n45217_not n45220 ; n45221
g44966 and n44647_not n45221_not ; n45222
g44967 and b[43] n44636_not ; n45223
g44968 and n44634_not n45223 ; n45224
g44969 and n44638_not n45224_not ; n45225
g44970 and n45222_not n45225 ; n45226
g44971 and n44638_not n45226_not ; n45227
g44972 and b[44] n44627_not ; n45228
g44973 and n44625_not n45228 ; n45229
g44974 and n44629_not n45229_not ; n45230
g44975 and n45227_not n45230 ; n45231
g44976 and n44629_not n45231_not ; n45232
g44977 and b[45] n44618_not ; n45233
g44978 and n44616_not n45233 ; n45234
g44979 and n44620_not n45234_not ; n45235
g44980 and n45232_not n45235 ; n45236
g44981 and n44620_not n45236_not ; n45237
g44982 and b[46] n44609_not ; n45238
g44983 and n44607_not n45238 ; n45239
g44984 and n44611_not n45239_not ; n45240
g44985 and n45237_not n45240 ; n45241
g44986 and n44611_not n45241_not ; n45242
g44987 and b[47] n44589_not ; n45243
g44988 and n44587_not n45243 ; n45244
g44989 and n44602_not n45244_not ; n45245
g44990 and n45242_not n45245 ; n45246
g44991 and n44602_not n45246_not ; n45247
g44992 and b[48] n44599_not ; n45248
g44993 and n44597_not n45248 ; n45249
g44994 and n44601_not n45249_not ; n45250
g44995 and n45247_not n45250 ; n45251
g44996 and n44601_not n45251_not ; n45252
g44997 and n408 n45252_not ; n45253
g44998 and n44590_not n45253_not ; n45254
g44999 and n44611_not n45245 ; n45255
g45000 and n45241_not n45255 ; n45256
g45001 and n45242_not n45245_not ; n45257
g45002 and n45256_not n45257_not ; n45258
g45003 and n408 n45258_not ; n45259
g45004 and n45252_not n45259 ; n45260
g45005 and n45254_not n45260_not ; n45261
g45006 and b[48]_not n45261_not ; n45262
g45007 and n44610_not n45253_not ; n45263
g45008 and n44620_not n45240 ; n45264
g45009 and n45236_not n45264 ; n45265
g45010 and n45237_not n45240_not ; n45266
g45011 and n45265_not n45266_not ; n45267
g45012 and n408 n45267_not ; n45268
g45013 and n45252_not n45268 ; n45269
g45014 and n45263_not n45269_not ; n45270
g45015 and b[47]_not n45270_not ; n45271
g45016 and n44619_not n45253_not ; n45272
g45017 and n44629_not n45235 ; n45273
g45018 and n45231_not n45273 ; n45274
g45019 and n45232_not n45235_not ; n45275
g45020 and n45274_not n45275_not ; n45276
g45021 and n408 n45276_not ; n45277
g45022 and n45252_not n45277 ; n45278
g45023 and n45272_not n45278_not ; n45279
g45024 and b[46]_not n45279_not ; n45280
g45025 and n44628_not n45253_not ; n45281
g45026 and n44638_not n45230 ; n45282
g45027 and n45226_not n45282 ; n45283
g45028 and n45227_not n45230_not ; n45284
g45029 and n45283_not n45284_not ; n45285
g45030 and n408 n45285_not ; n45286
g45031 and n45252_not n45286 ; n45287
g45032 and n45281_not n45287_not ; n45288
g45033 and b[45]_not n45288_not ; n45289
g45034 and n44637_not n45253_not ; n45290
g45035 and n44647_not n45225 ; n45291
g45036 and n45221_not n45291 ; n45292
g45037 and n45222_not n45225_not ; n45293
g45038 and n45292_not n45293_not ; n45294
g45039 and n408 n45294_not ; n45295
g45040 and n45252_not n45295 ; n45296
g45041 and n45290_not n45296_not ; n45297
g45042 and b[44]_not n45297_not ; n45298
g45043 and n44646_not n45253_not ; n45299
g45044 and n44656_not n45220 ; n45300
g45045 and n45216_not n45300 ; n45301
g45046 and n45217_not n45220_not ; n45302
g45047 and n45301_not n45302_not ; n45303
g45048 and n408 n45303_not ; n45304
g45049 and n45252_not n45304 ; n45305
g45050 and n45299_not n45305_not ; n45306
g45051 and b[43]_not n45306_not ; n45307
g45052 and n44655_not n45253_not ; n45308
g45053 and n44665_not n45215 ; n45309
g45054 and n45211_not n45309 ; n45310
g45055 and n45212_not n45215_not ; n45311
g45056 and n45310_not n45311_not ; n45312
g45057 and n408 n45312_not ; n45313
g45058 and n45252_not n45313 ; n45314
g45059 and n45308_not n45314_not ; n45315
g45060 and b[42]_not n45315_not ; n45316
g45061 and n44664_not n45253_not ; n45317
g45062 and n44674_not n45210 ; n45318
g45063 and n45206_not n45318 ; n45319
g45064 and n45207_not n45210_not ; n45320
g45065 and n45319_not n45320_not ; n45321
g45066 and n408 n45321_not ; n45322
g45067 and n45252_not n45322 ; n45323
g45068 and n45317_not n45323_not ; n45324
g45069 and b[41]_not n45324_not ; n45325
g45070 and n44673_not n45253_not ; n45326
g45071 and n44683_not n45205 ; n45327
g45072 and n45201_not n45327 ; n45328
g45073 and n45202_not n45205_not ; n45329
g45074 and n45328_not n45329_not ; n45330
g45075 and n408 n45330_not ; n45331
g45076 and n45252_not n45331 ; n45332
g45077 and n45326_not n45332_not ; n45333
g45078 and b[40]_not n45333_not ; n45334
g45079 and n44682_not n45253_not ; n45335
g45080 and n44692_not n45200 ; n45336
g45081 and n45196_not n45336 ; n45337
g45082 and n45197_not n45200_not ; n45338
g45083 and n45337_not n45338_not ; n45339
g45084 and n408 n45339_not ; n45340
g45085 and n45252_not n45340 ; n45341
g45086 and n45335_not n45341_not ; n45342
g45087 and b[39]_not n45342_not ; n45343
g45088 and n44691_not n45253_not ; n45344
g45089 and n44701_not n45195 ; n45345
g45090 and n45191_not n45345 ; n45346
g45091 and n45192_not n45195_not ; n45347
g45092 and n45346_not n45347_not ; n45348
g45093 and n408 n45348_not ; n45349
g45094 and n45252_not n45349 ; n45350
g45095 and n45344_not n45350_not ; n45351
g45096 and b[38]_not n45351_not ; n45352
g45097 and n44700_not n45253_not ; n45353
g45098 and n44710_not n45190 ; n45354
g45099 and n45186_not n45354 ; n45355
g45100 and n45187_not n45190_not ; n45356
g45101 and n45355_not n45356_not ; n45357
g45102 and n408 n45357_not ; n45358
g45103 and n45252_not n45358 ; n45359
g45104 and n45353_not n45359_not ; n45360
g45105 and b[37]_not n45360_not ; n45361
g45106 and n44709_not n45253_not ; n45362
g45107 and n44719_not n45185 ; n45363
g45108 and n45181_not n45363 ; n45364
g45109 and n45182_not n45185_not ; n45365
g45110 and n45364_not n45365_not ; n45366
g45111 and n408 n45366_not ; n45367
g45112 and n45252_not n45367 ; n45368
g45113 and n45362_not n45368_not ; n45369
g45114 and b[36]_not n45369_not ; n45370
g45115 and n44718_not n45253_not ; n45371
g45116 and n44728_not n45180 ; n45372
g45117 and n45176_not n45372 ; n45373
g45118 and n45177_not n45180_not ; n45374
g45119 and n45373_not n45374_not ; n45375
g45120 and n408 n45375_not ; n45376
g45121 and n45252_not n45376 ; n45377
g45122 and n45371_not n45377_not ; n45378
g45123 and b[35]_not n45378_not ; n45379
g45124 and n44727_not n45253_not ; n45380
g45125 and n44737_not n45175 ; n45381
g45126 and n45171_not n45381 ; n45382
g45127 and n45172_not n45175_not ; n45383
g45128 and n45382_not n45383_not ; n45384
g45129 and n408 n45384_not ; n45385
g45130 and n45252_not n45385 ; n45386
g45131 and n45380_not n45386_not ; n45387
g45132 and b[34]_not n45387_not ; n45388
g45133 and n44736_not n45253_not ; n45389
g45134 and n44746_not n45170 ; n45390
g45135 and n45166_not n45390 ; n45391
g45136 and n45167_not n45170_not ; n45392
g45137 and n45391_not n45392_not ; n45393
g45138 and n408 n45393_not ; n45394
g45139 and n45252_not n45394 ; n45395
g45140 and n45389_not n45395_not ; n45396
g45141 and b[33]_not n45396_not ; n45397
g45142 and n44745_not n45253_not ; n45398
g45143 and n44755_not n45165 ; n45399
g45144 and n45161_not n45399 ; n45400
g45145 and n45162_not n45165_not ; n45401
g45146 and n45400_not n45401_not ; n45402
g45147 and n408 n45402_not ; n45403
g45148 and n45252_not n45403 ; n45404
g45149 and n45398_not n45404_not ; n45405
g45150 and b[32]_not n45405_not ; n45406
g45151 and n44754_not n45253_not ; n45407
g45152 and n44764_not n45160 ; n45408
g45153 and n45156_not n45408 ; n45409
g45154 and n45157_not n45160_not ; n45410
g45155 and n45409_not n45410_not ; n45411
g45156 and n408 n45411_not ; n45412
g45157 and n45252_not n45412 ; n45413
g45158 and n45407_not n45413_not ; n45414
g45159 and b[31]_not n45414_not ; n45415
g45160 and n44763_not n45253_not ; n45416
g45161 and n44773_not n45155 ; n45417
g45162 and n45151_not n45417 ; n45418
g45163 and n45152_not n45155_not ; n45419
g45164 and n45418_not n45419_not ; n45420
g45165 and n408 n45420_not ; n45421
g45166 and n45252_not n45421 ; n45422
g45167 and n45416_not n45422_not ; n45423
g45168 and b[30]_not n45423_not ; n45424
g45169 and n44772_not n45253_not ; n45425
g45170 and n44782_not n45150 ; n45426
g45171 and n45146_not n45426 ; n45427
g45172 and n45147_not n45150_not ; n45428
g45173 and n45427_not n45428_not ; n45429
g45174 and n408 n45429_not ; n45430
g45175 and n45252_not n45430 ; n45431
g45176 and n45425_not n45431_not ; n45432
g45177 and b[29]_not n45432_not ; n45433
g45178 and n44781_not n45253_not ; n45434
g45179 and n44791_not n45145 ; n45435
g45180 and n45141_not n45435 ; n45436
g45181 and n45142_not n45145_not ; n45437
g45182 and n45436_not n45437_not ; n45438
g45183 and n408 n45438_not ; n45439
g45184 and n45252_not n45439 ; n45440
g45185 and n45434_not n45440_not ; n45441
g45186 and b[28]_not n45441_not ; n45442
g45187 and n44790_not n45253_not ; n45443
g45188 and n44800_not n45140 ; n45444
g45189 and n45136_not n45444 ; n45445
g45190 and n45137_not n45140_not ; n45446
g45191 and n45445_not n45446_not ; n45447
g45192 and n408 n45447_not ; n45448
g45193 and n45252_not n45448 ; n45449
g45194 and n45443_not n45449_not ; n45450
g45195 and b[27]_not n45450_not ; n45451
g45196 and n44799_not n45253_not ; n45452
g45197 and n44809_not n45135 ; n45453
g45198 and n45131_not n45453 ; n45454
g45199 and n45132_not n45135_not ; n45455
g45200 and n45454_not n45455_not ; n45456
g45201 and n408 n45456_not ; n45457
g45202 and n45252_not n45457 ; n45458
g45203 and n45452_not n45458_not ; n45459
g45204 and b[26]_not n45459_not ; n45460
g45205 and n44808_not n45253_not ; n45461
g45206 and n44818_not n45130 ; n45462
g45207 and n45126_not n45462 ; n45463
g45208 and n45127_not n45130_not ; n45464
g45209 and n45463_not n45464_not ; n45465
g45210 and n408 n45465_not ; n45466
g45211 and n45252_not n45466 ; n45467
g45212 and n45461_not n45467_not ; n45468
g45213 and b[25]_not n45468_not ; n45469
g45214 and n44817_not n45253_not ; n45470
g45215 and n44827_not n45125 ; n45471
g45216 and n45121_not n45471 ; n45472
g45217 and n45122_not n45125_not ; n45473
g45218 and n45472_not n45473_not ; n45474
g45219 and n408 n45474_not ; n45475
g45220 and n45252_not n45475 ; n45476
g45221 and n45470_not n45476_not ; n45477
g45222 and b[24]_not n45477_not ; n45478
g45223 and n44826_not n45253_not ; n45479
g45224 and n44836_not n45120 ; n45480
g45225 and n45116_not n45480 ; n45481
g45226 and n45117_not n45120_not ; n45482
g45227 and n45481_not n45482_not ; n45483
g45228 and n408 n45483_not ; n45484
g45229 and n45252_not n45484 ; n45485
g45230 and n45479_not n45485_not ; n45486
g45231 and b[23]_not n45486_not ; n45487
g45232 and n44835_not n45253_not ; n45488
g45233 and n44845_not n45115 ; n45489
g45234 and n45111_not n45489 ; n45490
g45235 and n45112_not n45115_not ; n45491
g45236 and n45490_not n45491_not ; n45492
g45237 and n408 n45492_not ; n45493
g45238 and n45252_not n45493 ; n45494
g45239 and n45488_not n45494_not ; n45495
g45240 and b[22]_not n45495_not ; n45496
g45241 and n44844_not n45253_not ; n45497
g45242 and n44854_not n45110 ; n45498
g45243 and n45106_not n45498 ; n45499
g45244 and n45107_not n45110_not ; n45500
g45245 and n45499_not n45500_not ; n45501
g45246 and n408 n45501_not ; n45502
g45247 and n45252_not n45502 ; n45503
g45248 and n45497_not n45503_not ; n45504
g45249 and b[21]_not n45504_not ; n45505
g45250 and n44853_not n45253_not ; n45506
g45251 and n44863_not n45105 ; n45507
g45252 and n45101_not n45507 ; n45508
g45253 and n45102_not n45105_not ; n45509
g45254 and n45508_not n45509_not ; n45510
g45255 and n408 n45510_not ; n45511
g45256 and n45252_not n45511 ; n45512
g45257 and n45506_not n45512_not ; n45513
g45258 and b[20]_not n45513_not ; n45514
g45259 and n44862_not n45253_not ; n45515
g45260 and n44872_not n45100 ; n45516
g45261 and n45096_not n45516 ; n45517
g45262 and n45097_not n45100_not ; n45518
g45263 and n45517_not n45518_not ; n45519
g45264 and n408 n45519_not ; n45520
g45265 and n45252_not n45520 ; n45521
g45266 and n45515_not n45521_not ; n45522
g45267 and b[19]_not n45522_not ; n45523
g45268 and n44871_not n45253_not ; n45524
g45269 and n44881_not n45095 ; n45525
g45270 and n45091_not n45525 ; n45526
g45271 and n45092_not n45095_not ; n45527
g45272 and n45526_not n45527_not ; n45528
g45273 and n408 n45528_not ; n45529
g45274 and n45252_not n45529 ; n45530
g45275 and n45524_not n45530_not ; n45531
g45276 and b[18]_not n45531_not ; n45532
g45277 and n44880_not n45253_not ; n45533
g45278 and n44890_not n45090 ; n45534
g45279 and n45086_not n45534 ; n45535
g45280 and n45087_not n45090_not ; n45536
g45281 and n45535_not n45536_not ; n45537
g45282 and n408 n45537_not ; n45538
g45283 and n45252_not n45538 ; n45539
g45284 and n45533_not n45539_not ; n45540
g45285 and b[17]_not n45540_not ; n45541
g45286 and n44889_not n45253_not ; n45542
g45287 and n44899_not n45085 ; n45543
g45288 and n45081_not n45543 ; n45544
g45289 and n45082_not n45085_not ; n45545
g45290 and n45544_not n45545_not ; n45546
g45291 and n408 n45546_not ; n45547
g45292 and n45252_not n45547 ; n45548
g45293 and n45542_not n45548_not ; n45549
g45294 and b[16]_not n45549_not ; n45550
g45295 and n44898_not n45253_not ; n45551
g45296 and n44908_not n45080 ; n45552
g45297 and n45076_not n45552 ; n45553
g45298 and n45077_not n45080_not ; n45554
g45299 and n45553_not n45554_not ; n45555
g45300 and n408 n45555_not ; n45556
g45301 and n45252_not n45556 ; n45557
g45302 and n45551_not n45557_not ; n45558
g45303 and b[15]_not n45558_not ; n45559
g45304 and n44907_not n45253_not ; n45560
g45305 and n44917_not n45075 ; n45561
g45306 and n45071_not n45561 ; n45562
g45307 and n45072_not n45075_not ; n45563
g45308 and n45562_not n45563_not ; n45564
g45309 and n408 n45564_not ; n45565
g45310 and n45252_not n45565 ; n45566
g45311 and n45560_not n45566_not ; n45567
g45312 and b[14]_not n45567_not ; n45568
g45313 and n44916_not n45253_not ; n45569
g45314 and n44926_not n45070 ; n45570
g45315 and n45066_not n45570 ; n45571
g45316 and n45067_not n45070_not ; n45572
g45317 and n45571_not n45572_not ; n45573
g45318 and n408 n45573_not ; n45574
g45319 and n45252_not n45574 ; n45575
g45320 and n45569_not n45575_not ; n45576
g45321 and b[13]_not n45576_not ; n45577
g45322 and n44925_not n45253_not ; n45578
g45323 and n44935_not n45065 ; n45579
g45324 and n45061_not n45579 ; n45580
g45325 and n45062_not n45065_not ; n45581
g45326 and n45580_not n45581_not ; n45582
g45327 and n408 n45582_not ; n45583
g45328 and n45252_not n45583 ; n45584
g45329 and n45578_not n45584_not ; n45585
g45330 and b[12]_not n45585_not ; n45586
g45331 and n44934_not n45253_not ; n45587
g45332 and n44944_not n45060 ; n45588
g45333 and n45056_not n45588 ; n45589
g45334 and n45057_not n45060_not ; n45590
g45335 and n45589_not n45590_not ; n45591
g45336 and n408 n45591_not ; n45592
g45337 and n45252_not n45592 ; n45593
g45338 and n45587_not n45593_not ; n45594
g45339 and b[11]_not n45594_not ; n45595
g45340 and n44943_not n45253_not ; n45596
g45341 and n44953_not n45055 ; n45597
g45342 and n45051_not n45597 ; n45598
g45343 and n45052_not n45055_not ; n45599
g45344 and n45598_not n45599_not ; n45600
g45345 and n408 n45600_not ; n45601
g45346 and n45252_not n45601 ; n45602
g45347 and n45596_not n45602_not ; n45603
g45348 and b[10]_not n45603_not ; n45604
g45349 and n44952_not n45253_not ; n45605
g45350 and n44962_not n45050 ; n45606
g45351 and n45046_not n45606 ; n45607
g45352 and n45047_not n45050_not ; n45608
g45353 and n45607_not n45608_not ; n45609
g45354 and n408 n45609_not ; n45610
g45355 and n45252_not n45610 ; n45611
g45356 and n45605_not n45611_not ; n45612
g45357 and b[9]_not n45612_not ; n45613
g45358 and n44961_not n45253_not ; n45614
g45359 and n44971_not n45045 ; n45615
g45360 and n45041_not n45615 ; n45616
g45361 and n45042_not n45045_not ; n45617
g45362 and n45616_not n45617_not ; n45618
g45363 and n408 n45618_not ; n45619
g45364 and n45252_not n45619 ; n45620
g45365 and n45614_not n45620_not ; n45621
g45366 and b[8]_not n45621_not ; n45622
g45367 and n44970_not n45253_not ; n45623
g45368 and n44980_not n45040 ; n45624
g45369 and n45036_not n45624 ; n45625
g45370 and n45037_not n45040_not ; n45626
g45371 and n45625_not n45626_not ; n45627
g45372 and n408 n45627_not ; n45628
g45373 and n45252_not n45628 ; n45629
g45374 and n45623_not n45629_not ; n45630
g45375 and b[7]_not n45630_not ; n45631
g45376 and n44979_not n45253_not ; n45632
g45377 and n44989_not n45035 ; n45633
g45378 and n45031_not n45633 ; n45634
g45379 and n45032_not n45035_not ; n45635
g45380 and n45634_not n45635_not ; n45636
g45381 and n408 n45636_not ; n45637
g45382 and n45252_not n45637 ; n45638
g45383 and n45632_not n45638_not ; n45639
g45384 and b[6]_not n45639_not ; n45640
g45385 and n44988_not n45253_not ; n45641
g45386 and n44998_not n45030 ; n45642
g45387 and n45026_not n45642 ; n45643
g45388 and n45027_not n45030_not ; n45644
g45389 and n45643_not n45644_not ; n45645
g45390 and n408 n45645_not ; n45646
g45391 and n45252_not n45646 ; n45647
g45392 and n45641_not n45647_not ; n45648
g45393 and b[5]_not n45648_not ; n45649
g45394 and n44997_not n45253_not ; n45650
g45395 and n45006_not n45025 ; n45651
g45396 and n45021_not n45651 ; n45652
g45397 and n45022_not n45025_not ; n45653
g45398 and n45652_not n45653_not ; n45654
g45399 and n408 n45654_not ; n45655
g45400 and n45252_not n45655 ; n45656
g45401 and n45650_not n45656_not ; n45657
g45402 and b[4]_not n45657_not ; n45658
g45403 and n45005_not n45253_not ; n45659
g45404 and n45016_not n45020 ; n45660
g45405 and n45015_not n45660 ; n45661
g45406 and n45017_not n45020_not ; n45662
g45407 and n45661_not n45662_not ; n45663
g45408 and n408 n45663_not ; n45664
g45409 and n45252_not n45664 ; n45665
g45410 and n45659_not n45665_not ; n45666
g45411 and b[3]_not n45666_not ; n45667
g45412 and n45010_not n45253_not ; n45668
g45413 and n16956 n45013_not ; n45669
g45414 and n45011_not n45669 ; n45670
g45415 and n408 n45670_not ; n45671
g45416 and n45015_not n45671 ; n45672
g45417 and n45252_not n45672 ; n45673
g45418 and n45668_not n45673_not ; n45674
g45419 and b[2]_not n45674_not ; n45675
g45420 and n17621 n45252_not ; n45676
g45421 and a[15] n45676_not ; n45677
g45422 and n17625 n45252_not ; n45678
g45423 and n45677_not n45678_not ; n45679
g45424 and b[1] n45679_not ; n45680
g45425 and b[1]_not n45678_not ; n45681
g45426 and n45677_not n45681 ; n45682
g45427 and n45680_not n45682_not ; n45683
g45428 and n17632_not n45683_not ; n45684
g45429 and b[1]_not n45679_not ; n45685
g45430 and n45684_not n45685_not ; n45686
g45431 and b[2] n45673_not ; n45687
g45432 and n45668_not n45687 ; n45688
g45433 and n45675_not n45688_not ; n45689
g45434 and n45686_not n45689 ; n45690
g45435 and n45675_not n45690_not ; n45691
g45436 and b[3] n45665_not ; n45692
g45437 and n45659_not n45692 ; n45693
g45438 and n45667_not n45693_not ; n45694
g45439 and n45691_not n45694 ; n45695
g45440 and n45667_not n45695_not ; n45696
g45441 and b[4] n45656_not ; n45697
g45442 and n45650_not n45697 ; n45698
g45443 and n45658_not n45698_not ; n45699
g45444 and n45696_not n45699 ; n45700
g45445 and n45658_not n45700_not ; n45701
g45446 and b[5] n45647_not ; n45702
g45447 and n45641_not n45702 ; n45703
g45448 and n45649_not n45703_not ; n45704
g45449 and n45701_not n45704 ; n45705
g45450 and n45649_not n45705_not ; n45706
g45451 and b[6] n45638_not ; n45707
g45452 and n45632_not n45707 ; n45708
g45453 and n45640_not n45708_not ; n45709
g45454 and n45706_not n45709 ; n45710
g45455 and n45640_not n45710_not ; n45711
g45456 and b[7] n45629_not ; n45712
g45457 and n45623_not n45712 ; n45713
g45458 and n45631_not n45713_not ; n45714
g45459 and n45711_not n45714 ; n45715
g45460 and n45631_not n45715_not ; n45716
g45461 and b[8] n45620_not ; n45717
g45462 and n45614_not n45717 ; n45718
g45463 and n45622_not n45718_not ; n45719
g45464 and n45716_not n45719 ; n45720
g45465 and n45622_not n45720_not ; n45721
g45466 and b[9] n45611_not ; n45722
g45467 and n45605_not n45722 ; n45723
g45468 and n45613_not n45723_not ; n45724
g45469 and n45721_not n45724 ; n45725
g45470 and n45613_not n45725_not ; n45726
g45471 and b[10] n45602_not ; n45727
g45472 and n45596_not n45727 ; n45728
g45473 and n45604_not n45728_not ; n45729
g45474 and n45726_not n45729 ; n45730
g45475 and n45604_not n45730_not ; n45731
g45476 and b[11] n45593_not ; n45732
g45477 and n45587_not n45732 ; n45733
g45478 and n45595_not n45733_not ; n45734
g45479 and n45731_not n45734 ; n45735
g45480 and n45595_not n45735_not ; n45736
g45481 and b[12] n45584_not ; n45737
g45482 and n45578_not n45737 ; n45738
g45483 and n45586_not n45738_not ; n45739
g45484 and n45736_not n45739 ; n45740
g45485 and n45586_not n45740_not ; n45741
g45486 and b[13] n45575_not ; n45742
g45487 and n45569_not n45742 ; n45743
g45488 and n45577_not n45743_not ; n45744
g45489 and n45741_not n45744 ; n45745
g45490 and n45577_not n45745_not ; n45746
g45491 and b[14] n45566_not ; n45747
g45492 and n45560_not n45747 ; n45748
g45493 and n45568_not n45748_not ; n45749
g45494 and n45746_not n45749 ; n45750
g45495 and n45568_not n45750_not ; n45751
g45496 and b[15] n45557_not ; n45752
g45497 and n45551_not n45752 ; n45753
g45498 and n45559_not n45753_not ; n45754
g45499 and n45751_not n45754 ; n45755
g45500 and n45559_not n45755_not ; n45756
g45501 and b[16] n45548_not ; n45757
g45502 and n45542_not n45757 ; n45758
g45503 and n45550_not n45758_not ; n45759
g45504 and n45756_not n45759 ; n45760
g45505 and n45550_not n45760_not ; n45761
g45506 and b[17] n45539_not ; n45762
g45507 and n45533_not n45762 ; n45763
g45508 and n45541_not n45763_not ; n45764
g45509 and n45761_not n45764 ; n45765
g45510 and n45541_not n45765_not ; n45766
g45511 and b[18] n45530_not ; n45767
g45512 and n45524_not n45767 ; n45768
g45513 and n45532_not n45768_not ; n45769
g45514 and n45766_not n45769 ; n45770
g45515 and n45532_not n45770_not ; n45771
g45516 and b[19] n45521_not ; n45772
g45517 and n45515_not n45772 ; n45773
g45518 and n45523_not n45773_not ; n45774
g45519 and n45771_not n45774 ; n45775
g45520 and n45523_not n45775_not ; n45776
g45521 and b[20] n45512_not ; n45777
g45522 and n45506_not n45777 ; n45778
g45523 and n45514_not n45778_not ; n45779
g45524 and n45776_not n45779 ; n45780
g45525 and n45514_not n45780_not ; n45781
g45526 and b[21] n45503_not ; n45782
g45527 and n45497_not n45782 ; n45783
g45528 and n45505_not n45783_not ; n45784
g45529 and n45781_not n45784 ; n45785
g45530 and n45505_not n45785_not ; n45786
g45531 and b[22] n45494_not ; n45787
g45532 and n45488_not n45787 ; n45788
g45533 and n45496_not n45788_not ; n45789
g45534 and n45786_not n45789 ; n45790
g45535 and n45496_not n45790_not ; n45791
g45536 and b[23] n45485_not ; n45792
g45537 and n45479_not n45792 ; n45793
g45538 and n45487_not n45793_not ; n45794
g45539 and n45791_not n45794 ; n45795
g45540 and n45487_not n45795_not ; n45796
g45541 and b[24] n45476_not ; n45797
g45542 and n45470_not n45797 ; n45798
g45543 and n45478_not n45798_not ; n45799
g45544 and n45796_not n45799 ; n45800
g45545 and n45478_not n45800_not ; n45801
g45546 and b[25] n45467_not ; n45802
g45547 and n45461_not n45802 ; n45803
g45548 and n45469_not n45803_not ; n45804
g45549 and n45801_not n45804 ; n45805
g45550 and n45469_not n45805_not ; n45806
g45551 and b[26] n45458_not ; n45807
g45552 and n45452_not n45807 ; n45808
g45553 and n45460_not n45808_not ; n45809
g45554 and n45806_not n45809 ; n45810
g45555 and n45460_not n45810_not ; n45811
g45556 and b[27] n45449_not ; n45812
g45557 and n45443_not n45812 ; n45813
g45558 and n45451_not n45813_not ; n45814
g45559 and n45811_not n45814 ; n45815
g45560 and n45451_not n45815_not ; n45816
g45561 and b[28] n45440_not ; n45817
g45562 and n45434_not n45817 ; n45818
g45563 and n45442_not n45818_not ; n45819
g45564 and n45816_not n45819 ; n45820
g45565 and n45442_not n45820_not ; n45821
g45566 and b[29] n45431_not ; n45822
g45567 and n45425_not n45822 ; n45823
g45568 and n45433_not n45823_not ; n45824
g45569 and n45821_not n45824 ; n45825
g45570 and n45433_not n45825_not ; n45826
g45571 and b[30] n45422_not ; n45827
g45572 and n45416_not n45827 ; n45828
g45573 and n45424_not n45828_not ; n45829
g45574 and n45826_not n45829 ; n45830
g45575 and n45424_not n45830_not ; n45831
g45576 and b[31] n45413_not ; n45832
g45577 and n45407_not n45832 ; n45833
g45578 and n45415_not n45833_not ; n45834
g45579 and n45831_not n45834 ; n45835
g45580 and n45415_not n45835_not ; n45836
g45581 and b[32] n45404_not ; n45837
g45582 and n45398_not n45837 ; n45838
g45583 and n45406_not n45838_not ; n45839
g45584 and n45836_not n45839 ; n45840
g45585 and n45406_not n45840_not ; n45841
g45586 and b[33] n45395_not ; n45842
g45587 and n45389_not n45842 ; n45843
g45588 and n45397_not n45843_not ; n45844
g45589 and n45841_not n45844 ; n45845
g45590 and n45397_not n45845_not ; n45846
g45591 and b[34] n45386_not ; n45847
g45592 and n45380_not n45847 ; n45848
g45593 and n45388_not n45848_not ; n45849
g45594 and n45846_not n45849 ; n45850
g45595 and n45388_not n45850_not ; n45851
g45596 and b[35] n45377_not ; n45852
g45597 and n45371_not n45852 ; n45853
g45598 and n45379_not n45853_not ; n45854
g45599 and n45851_not n45854 ; n45855
g45600 and n45379_not n45855_not ; n45856
g45601 and b[36] n45368_not ; n45857
g45602 and n45362_not n45857 ; n45858
g45603 and n45370_not n45858_not ; n45859
g45604 and n45856_not n45859 ; n45860
g45605 and n45370_not n45860_not ; n45861
g45606 and b[37] n45359_not ; n45862
g45607 and n45353_not n45862 ; n45863
g45608 and n45361_not n45863_not ; n45864
g45609 and n45861_not n45864 ; n45865
g45610 and n45361_not n45865_not ; n45866
g45611 and b[38] n45350_not ; n45867
g45612 and n45344_not n45867 ; n45868
g45613 and n45352_not n45868_not ; n45869
g45614 and n45866_not n45869 ; n45870
g45615 and n45352_not n45870_not ; n45871
g45616 and b[39] n45341_not ; n45872
g45617 and n45335_not n45872 ; n45873
g45618 and n45343_not n45873_not ; n45874
g45619 and n45871_not n45874 ; n45875
g45620 and n45343_not n45875_not ; n45876
g45621 and b[40] n45332_not ; n45877
g45622 and n45326_not n45877 ; n45878
g45623 and n45334_not n45878_not ; n45879
g45624 and n45876_not n45879 ; n45880
g45625 and n45334_not n45880_not ; n45881
g45626 and b[41] n45323_not ; n45882
g45627 and n45317_not n45882 ; n45883
g45628 and n45325_not n45883_not ; n45884
g45629 and n45881_not n45884 ; n45885
g45630 and n45325_not n45885_not ; n45886
g45631 and b[42] n45314_not ; n45887
g45632 and n45308_not n45887 ; n45888
g45633 and n45316_not n45888_not ; n45889
g45634 and n45886_not n45889 ; n45890
g45635 and n45316_not n45890_not ; n45891
g45636 and b[43] n45305_not ; n45892
g45637 and n45299_not n45892 ; n45893
g45638 and n45307_not n45893_not ; n45894
g45639 and n45891_not n45894 ; n45895
g45640 and n45307_not n45895_not ; n45896
g45641 and b[44] n45296_not ; n45897
g45642 and n45290_not n45897 ; n45898
g45643 and n45298_not n45898_not ; n45899
g45644 and n45896_not n45899 ; n45900
g45645 and n45298_not n45900_not ; n45901
g45646 and b[45] n45287_not ; n45902
g45647 and n45281_not n45902 ; n45903
g45648 and n45289_not n45903_not ; n45904
g45649 and n45901_not n45904 ; n45905
g45650 and n45289_not n45905_not ; n45906
g45651 and b[46] n45278_not ; n45907
g45652 and n45272_not n45907 ; n45908
g45653 and n45280_not n45908_not ; n45909
g45654 and n45906_not n45909 ; n45910
g45655 and n45280_not n45910_not ; n45911
g45656 and b[47] n45269_not ; n45912
g45657 and n45263_not n45912 ; n45913
g45658 and n45271_not n45913_not ; n45914
g45659 and n45911_not n45914 ; n45915
g45660 and n45271_not n45915_not ; n45916
g45661 and b[48] n45260_not ; n45917
g45662 and n45254_not n45917 ; n45918
g45663 and n45262_not n45918_not ; n45919
g45664 and n45916_not n45919 ; n45920
g45665 and n45262_not n45920_not ; n45921
g45666 and n44600_not n45253_not ; n45922
g45667 and n44602_not n45250 ; n45923
g45668 and n45246_not n45923 ; n45924
g45669 and n45247_not n45250_not ; n45925
g45670 and n45924_not n45925_not ; n45926
g45671 and n45253 n45926_not ; n45927
g45672 and n45922_not n45927_not ; n45928
g45673 and b[49]_not n45928_not ; n45929
g45674 and b[49] n45922_not ; n45930
g45675 and n45927_not n45930 ; n45931
g45676 and n17882 n45931_not ; n45932
g45677 and n45929_not n45932 ; n45933
g45678 and n45921_not n45933 ; n45934
g45679 and n408 n45928_not ; n45935
g45680 and n45934_not n45935_not ; n45936
g45681 and n45271_not n45919 ; n45937
g45682 and n45915_not n45937 ; n45938
g45683 and n45916_not n45919_not ; n45939
g45684 and n45938_not n45939_not ; n45940
g45685 and n45936_not n45940_not ; n45941
g45686 and n45261_not n45935_not ; n45942
g45687 and n45934_not n45942 ; n45943
g45688 and n45941_not n45943_not ; n45944
g45689 and b[49]_not n45944_not ; n45945
g45690 and n45280_not n45914 ; n45946
g45691 and n45910_not n45946 ; n45947
g45692 and n45911_not n45914_not ; n45948
g45693 and n45947_not n45948_not ; n45949
g45694 and n45936_not n45949_not ; n45950
g45695 and n45270_not n45935_not ; n45951
g45696 and n45934_not n45951 ; n45952
g45697 and n45950_not n45952_not ; n45953
g45698 and b[48]_not n45953_not ; n45954
g45699 and n45289_not n45909 ; n45955
g45700 and n45905_not n45955 ; n45956
g45701 and n45906_not n45909_not ; n45957
g45702 and n45956_not n45957_not ; n45958
g45703 and n45936_not n45958_not ; n45959
g45704 and n45279_not n45935_not ; n45960
g45705 and n45934_not n45960 ; n45961
g45706 and n45959_not n45961_not ; n45962
g45707 and b[47]_not n45962_not ; n45963
g45708 and n45298_not n45904 ; n45964
g45709 and n45900_not n45964 ; n45965
g45710 and n45901_not n45904_not ; n45966
g45711 and n45965_not n45966_not ; n45967
g45712 and n45936_not n45967_not ; n45968
g45713 and n45288_not n45935_not ; n45969
g45714 and n45934_not n45969 ; n45970
g45715 and n45968_not n45970_not ; n45971
g45716 and b[46]_not n45971_not ; n45972
g45717 and n45307_not n45899 ; n45973
g45718 and n45895_not n45973 ; n45974
g45719 and n45896_not n45899_not ; n45975
g45720 and n45974_not n45975_not ; n45976
g45721 and n45936_not n45976_not ; n45977
g45722 and n45297_not n45935_not ; n45978
g45723 and n45934_not n45978 ; n45979
g45724 and n45977_not n45979_not ; n45980
g45725 and b[45]_not n45980_not ; n45981
g45726 and n45316_not n45894 ; n45982
g45727 and n45890_not n45982 ; n45983
g45728 and n45891_not n45894_not ; n45984
g45729 and n45983_not n45984_not ; n45985
g45730 and n45936_not n45985_not ; n45986
g45731 and n45306_not n45935_not ; n45987
g45732 and n45934_not n45987 ; n45988
g45733 and n45986_not n45988_not ; n45989
g45734 and b[44]_not n45989_not ; n45990
g45735 and n45325_not n45889 ; n45991
g45736 and n45885_not n45991 ; n45992
g45737 and n45886_not n45889_not ; n45993
g45738 and n45992_not n45993_not ; n45994
g45739 and n45936_not n45994_not ; n45995
g45740 and n45315_not n45935_not ; n45996
g45741 and n45934_not n45996 ; n45997
g45742 and n45995_not n45997_not ; n45998
g45743 and b[43]_not n45998_not ; n45999
g45744 and n45334_not n45884 ; n46000
g45745 and n45880_not n46000 ; n46001
g45746 and n45881_not n45884_not ; n46002
g45747 and n46001_not n46002_not ; n46003
g45748 and n45936_not n46003_not ; n46004
g45749 and n45324_not n45935_not ; n46005
g45750 and n45934_not n46005 ; n46006
g45751 and n46004_not n46006_not ; n46007
g45752 and b[42]_not n46007_not ; n46008
g45753 and n45343_not n45879 ; n46009
g45754 and n45875_not n46009 ; n46010
g45755 and n45876_not n45879_not ; n46011
g45756 and n46010_not n46011_not ; n46012
g45757 and n45936_not n46012_not ; n46013
g45758 and n45333_not n45935_not ; n46014
g45759 and n45934_not n46014 ; n46015
g45760 and n46013_not n46015_not ; n46016
g45761 and b[41]_not n46016_not ; n46017
g45762 and n45352_not n45874 ; n46018
g45763 and n45870_not n46018 ; n46019
g45764 and n45871_not n45874_not ; n46020
g45765 and n46019_not n46020_not ; n46021
g45766 and n45936_not n46021_not ; n46022
g45767 and n45342_not n45935_not ; n46023
g45768 and n45934_not n46023 ; n46024
g45769 and n46022_not n46024_not ; n46025
g45770 and b[40]_not n46025_not ; n46026
g45771 and n45361_not n45869 ; n46027
g45772 and n45865_not n46027 ; n46028
g45773 and n45866_not n45869_not ; n46029
g45774 and n46028_not n46029_not ; n46030
g45775 and n45936_not n46030_not ; n46031
g45776 and n45351_not n45935_not ; n46032
g45777 and n45934_not n46032 ; n46033
g45778 and n46031_not n46033_not ; n46034
g45779 and b[39]_not n46034_not ; n46035
g45780 and n45370_not n45864 ; n46036
g45781 and n45860_not n46036 ; n46037
g45782 and n45861_not n45864_not ; n46038
g45783 and n46037_not n46038_not ; n46039
g45784 and n45936_not n46039_not ; n46040
g45785 and n45360_not n45935_not ; n46041
g45786 and n45934_not n46041 ; n46042
g45787 and n46040_not n46042_not ; n46043
g45788 and b[38]_not n46043_not ; n46044
g45789 and n45379_not n45859 ; n46045
g45790 and n45855_not n46045 ; n46046
g45791 and n45856_not n45859_not ; n46047
g45792 and n46046_not n46047_not ; n46048
g45793 and n45936_not n46048_not ; n46049
g45794 and n45369_not n45935_not ; n46050
g45795 and n45934_not n46050 ; n46051
g45796 and n46049_not n46051_not ; n46052
g45797 and b[37]_not n46052_not ; n46053
g45798 and n45388_not n45854 ; n46054
g45799 and n45850_not n46054 ; n46055
g45800 and n45851_not n45854_not ; n46056
g45801 and n46055_not n46056_not ; n46057
g45802 and n45936_not n46057_not ; n46058
g45803 and n45378_not n45935_not ; n46059
g45804 and n45934_not n46059 ; n46060
g45805 and n46058_not n46060_not ; n46061
g45806 and b[36]_not n46061_not ; n46062
g45807 and n45397_not n45849 ; n46063
g45808 and n45845_not n46063 ; n46064
g45809 and n45846_not n45849_not ; n46065
g45810 and n46064_not n46065_not ; n46066
g45811 and n45936_not n46066_not ; n46067
g45812 and n45387_not n45935_not ; n46068
g45813 and n45934_not n46068 ; n46069
g45814 and n46067_not n46069_not ; n46070
g45815 and b[35]_not n46070_not ; n46071
g45816 and n45406_not n45844 ; n46072
g45817 and n45840_not n46072 ; n46073
g45818 and n45841_not n45844_not ; n46074
g45819 and n46073_not n46074_not ; n46075
g45820 and n45936_not n46075_not ; n46076
g45821 and n45396_not n45935_not ; n46077
g45822 and n45934_not n46077 ; n46078
g45823 and n46076_not n46078_not ; n46079
g45824 and b[34]_not n46079_not ; n46080
g45825 and n45415_not n45839 ; n46081
g45826 and n45835_not n46081 ; n46082
g45827 and n45836_not n45839_not ; n46083
g45828 and n46082_not n46083_not ; n46084
g45829 and n45936_not n46084_not ; n46085
g45830 and n45405_not n45935_not ; n46086
g45831 and n45934_not n46086 ; n46087
g45832 and n46085_not n46087_not ; n46088
g45833 and b[33]_not n46088_not ; n46089
g45834 and n45424_not n45834 ; n46090
g45835 and n45830_not n46090 ; n46091
g45836 and n45831_not n45834_not ; n46092
g45837 and n46091_not n46092_not ; n46093
g45838 and n45936_not n46093_not ; n46094
g45839 and n45414_not n45935_not ; n46095
g45840 and n45934_not n46095 ; n46096
g45841 and n46094_not n46096_not ; n46097
g45842 and b[32]_not n46097_not ; n46098
g45843 and n45433_not n45829 ; n46099
g45844 and n45825_not n46099 ; n46100
g45845 and n45826_not n45829_not ; n46101
g45846 and n46100_not n46101_not ; n46102
g45847 and n45936_not n46102_not ; n46103
g45848 and n45423_not n45935_not ; n46104
g45849 and n45934_not n46104 ; n46105
g45850 and n46103_not n46105_not ; n46106
g45851 and b[31]_not n46106_not ; n46107
g45852 and n45442_not n45824 ; n46108
g45853 and n45820_not n46108 ; n46109
g45854 and n45821_not n45824_not ; n46110
g45855 and n46109_not n46110_not ; n46111
g45856 and n45936_not n46111_not ; n46112
g45857 and n45432_not n45935_not ; n46113
g45858 and n45934_not n46113 ; n46114
g45859 and n46112_not n46114_not ; n46115
g45860 and b[30]_not n46115_not ; n46116
g45861 and n45451_not n45819 ; n46117
g45862 and n45815_not n46117 ; n46118
g45863 and n45816_not n45819_not ; n46119
g45864 and n46118_not n46119_not ; n46120
g45865 and n45936_not n46120_not ; n46121
g45866 and n45441_not n45935_not ; n46122
g45867 and n45934_not n46122 ; n46123
g45868 and n46121_not n46123_not ; n46124
g45869 and b[29]_not n46124_not ; n46125
g45870 and n45460_not n45814 ; n46126
g45871 and n45810_not n46126 ; n46127
g45872 and n45811_not n45814_not ; n46128
g45873 and n46127_not n46128_not ; n46129
g45874 and n45936_not n46129_not ; n46130
g45875 and n45450_not n45935_not ; n46131
g45876 and n45934_not n46131 ; n46132
g45877 and n46130_not n46132_not ; n46133
g45878 and b[28]_not n46133_not ; n46134
g45879 and n45469_not n45809 ; n46135
g45880 and n45805_not n46135 ; n46136
g45881 and n45806_not n45809_not ; n46137
g45882 and n46136_not n46137_not ; n46138
g45883 and n45936_not n46138_not ; n46139
g45884 and n45459_not n45935_not ; n46140
g45885 and n45934_not n46140 ; n46141
g45886 and n46139_not n46141_not ; n46142
g45887 and b[27]_not n46142_not ; n46143
g45888 and n45478_not n45804 ; n46144
g45889 and n45800_not n46144 ; n46145
g45890 and n45801_not n45804_not ; n46146
g45891 and n46145_not n46146_not ; n46147
g45892 and n45936_not n46147_not ; n46148
g45893 and n45468_not n45935_not ; n46149
g45894 and n45934_not n46149 ; n46150
g45895 and n46148_not n46150_not ; n46151
g45896 and b[26]_not n46151_not ; n46152
g45897 and n45487_not n45799 ; n46153
g45898 and n45795_not n46153 ; n46154
g45899 and n45796_not n45799_not ; n46155
g45900 and n46154_not n46155_not ; n46156
g45901 and n45936_not n46156_not ; n46157
g45902 and n45477_not n45935_not ; n46158
g45903 and n45934_not n46158 ; n46159
g45904 and n46157_not n46159_not ; n46160
g45905 and b[25]_not n46160_not ; n46161
g45906 and n45496_not n45794 ; n46162
g45907 and n45790_not n46162 ; n46163
g45908 and n45791_not n45794_not ; n46164
g45909 and n46163_not n46164_not ; n46165
g45910 and n45936_not n46165_not ; n46166
g45911 and n45486_not n45935_not ; n46167
g45912 and n45934_not n46167 ; n46168
g45913 and n46166_not n46168_not ; n46169
g45914 and b[24]_not n46169_not ; n46170
g45915 and n45505_not n45789 ; n46171
g45916 and n45785_not n46171 ; n46172
g45917 and n45786_not n45789_not ; n46173
g45918 and n46172_not n46173_not ; n46174
g45919 and n45936_not n46174_not ; n46175
g45920 and n45495_not n45935_not ; n46176
g45921 and n45934_not n46176 ; n46177
g45922 and n46175_not n46177_not ; n46178
g45923 and b[23]_not n46178_not ; n46179
g45924 and n45514_not n45784 ; n46180
g45925 and n45780_not n46180 ; n46181
g45926 and n45781_not n45784_not ; n46182
g45927 and n46181_not n46182_not ; n46183
g45928 and n45936_not n46183_not ; n46184
g45929 and n45504_not n45935_not ; n46185
g45930 and n45934_not n46185 ; n46186
g45931 and n46184_not n46186_not ; n46187
g45932 and b[22]_not n46187_not ; n46188
g45933 and n45523_not n45779 ; n46189
g45934 and n45775_not n46189 ; n46190
g45935 and n45776_not n45779_not ; n46191
g45936 and n46190_not n46191_not ; n46192
g45937 and n45936_not n46192_not ; n46193
g45938 and n45513_not n45935_not ; n46194
g45939 and n45934_not n46194 ; n46195
g45940 and n46193_not n46195_not ; n46196
g45941 and b[21]_not n46196_not ; n46197
g45942 and n45532_not n45774 ; n46198
g45943 and n45770_not n46198 ; n46199
g45944 and n45771_not n45774_not ; n46200
g45945 and n46199_not n46200_not ; n46201
g45946 and n45936_not n46201_not ; n46202
g45947 and n45522_not n45935_not ; n46203
g45948 and n45934_not n46203 ; n46204
g45949 and n46202_not n46204_not ; n46205
g45950 and b[20]_not n46205_not ; n46206
g45951 and n45541_not n45769 ; n46207
g45952 and n45765_not n46207 ; n46208
g45953 and n45766_not n45769_not ; n46209
g45954 and n46208_not n46209_not ; n46210
g45955 and n45936_not n46210_not ; n46211
g45956 and n45531_not n45935_not ; n46212
g45957 and n45934_not n46212 ; n46213
g45958 and n46211_not n46213_not ; n46214
g45959 and b[19]_not n46214_not ; n46215
g45960 and n45550_not n45764 ; n46216
g45961 and n45760_not n46216 ; n46217
g45962 and n45761_not n45764_not ; n46218
g45963 and n46217_not n46218_not ; n46219
g45964 and n45936_not n46219_not ; n46220
g45965 and n45540_not n45935_not ; n46221
g45966 and n45934_not n46221 ; n46222
g45967 and n46220_not n46222_not ; n46223
g45968 and b[18]_not n46223_not ; n46224
g45969 and n45559_not n45759 ; n46225
g45970 and n45755_not n46225 ; n46226
g45971 and n45756_not n45759_not ; n46227
g45972 and n46226_not n46227_not ; n46228
g45973 and n45936_not n46228_not ; n46229
g45974 and n45549_not n45935_not ; n46230
g45975 and n45934_not n46230 ; n46231
g45976 and n46229_not n46231_not ; n46232
g45977 and b[17]_not n46232_not ; n46233
g45978 and n45568_not n45754 ; n46234
g45979 and n45750_not n46234 ; n46235
g45980 and n45751_not n45754_not ; n46236
g45981 and n46235_not n46236_not ; n46237
g45982 and n45936_not n46237_not ; n46238
g45983 and n45558_not n45935_not ; n46239
g45984 and n45934_not n46239 ; n46240
g45985 and n46238_not n46240_not ; n46241
g45986 and b[16]_not n46241_not ; n46242
g45987 and n45577_not n45749 ; n46243
g45988 and n45745_not n46243 ; n46244
g45989 and n45746_not n45749_not ; n46245
g45990 and n46244_not n46245_not ; n46246
g45991 and n45936_not n46246_not ; n46247
g45992 and n45567_not n45935_not ; n46248
g45993 and n45934_not n46248 ; n46249
g45994 and n46247_not n46249_not ; n46250
g45995 and b[15]_not n46250_not ; n46251
g45996 and n45586_not n45744 ; n46252
g45997 and n45740_not n46252 ; n46253
g45998 and n45741_not n45744_not ; n46254
g45999 and n46253_not n46254_not ; n46255
g46000 and n45936_not n46255_not ; n46256
g46001 and n45576_not n45935_not ; n46257
g46002 and n45934_not n46257 ; n46258
g46003 and n46256_not n46258_not ; n46259
g46004 and b[14]_not n46259_not ; n46260
g46005 and n45595_not n45739 ; n46261
g46006 and n45735_not n46261 ; n46262
g46007 and n45736_not n45739_not ; n46263
g46008 and n46262_not n46263_not ; n46264
g46009 and n45936_not n46264_not ; n46265
g46010 and n45585_not n45935_not ; n46266
g46011 and n45934_not n46266 ; n46267
g46012 and n46265_not n46267_not ; n46268
g46013 and b[13]_not n46268_not ; n46269
g46014 and n45604_not n45734 ; n46270
g46015 and n45730_not n46270 ; n46271
g46016 and n45731_not n45734_not ; n46272
g46017 and n46271_not n46272_not ; n46273
g46018 and n45936_not n46273_not ; n46274
g46019 and n45594_not n45935_not ; n46275
g46020 and n45934_not n46275 ; n46276
g46021 and n46274_not n46276_not ; n46277
g46022 and b[12]_not n46277_not ; n46278
g46023 and n45613_not n45729 ; n46279
g46024 and n45725_not n46279 ; n46280
g46025 and n45726_not n45729_not ; n46281
g46026 and n46280_not n46281_not ; n46282
g46027 and n45936_not n46282_not ; n46283
g46028 and n45603_not n45935_not ; n46284
g46029 and n45934_not n46284 ; n46285
g46030 and n46283_not n46285_not ; n46286
g46031 and b[11]_not n46286_not ; n46287
g46032 and n45622_not n45724 ; n46288
g46033 and n45720_not n46288 ; n46289
g46034 and n45721_not n45724_not ; n46290
g46035 and n46289_not n46290_not ; n46291
g46036 and n45936_not n46291_not ; n46292
g46037 and n45612_not n45935_not ; n46293
g46038 and n45934_not n46293 ; n46294
g46039 and n46292_not n46294_not ; n46295
g46040 and b[10]_not n46295_not ; n46296
g46041 and n45631_not n45719 ; n46297
g46042 and n45715_not n46297 ; n46298
g46043 and n45716_not n45719_not ; n46299
g46044 and n46298_not n46299_not ; n46300
g46045 and n45936_not n46300_not ; n46301
g46046 and n45621_not n45935_not ; n46302
g46047 and n45934_not n46302 ; n46303
g46048 and n46301_not n46303_not ; n46304
g46049 and b[9]_not n46304_not ; n46305
g46050 and n45640_not n45714 ; n46306
g46051 and n45710_not n46306 ; n46307
g46052 and n45711_not n45714_not ; n46308
g46053 and n46307_not n46308_not ; n46309
g46054 and n45936_not n46309_not ; n46310
g46055 and n45630_not n45935_not ; n46311
g46056 and n45934_not n46311 ; n46312
g46057 and n46310_not n46312_not ; n46313
g46058 and b[8]_not n46313_not ; n46314
g46059 and n45649_not n45709 ; n46315
g46060 and n45705_not n46315 ; n46316
g46061 and n45706_not n45709_not ; n46317
g46062 and n46316_not n46317_not ; n46318
g46063 and n45936_not n46318_not ; n46319
g46064 and n45639_not n45935_not ; n46320
g46065 and n45934_not n46320 ; n46321
g46066 and n46319_not n46321_not ; n46322
g46067 and b[7]_not n46322_not ; n46323
g46068 and n45658_not n45704 ; n46324
g46069 and n45700_not n46324 ; n46325
g46070 and n45701_not n45704_not ; n46326
g46071 and n46325_not n46326_not ; n46327
g46072 and n45936_not n46327_not ; n46328
g46073 and n45648_not n45935_not ; n46329
g46074 and n45934_not n46329 ; n46330
g46075 and n46328_not n46330_not ; n46331
g46076 and b[6]_not n46331_not ; n46332
g46077 and n45667_not n45699 ; n46333
g46078 and n45695_not n46333 ; n46334
g46079 and n45696_not n45699_not ; n46335
g46080 and n46334_not n46335_not ; n46336
g46081 and n45936_not n46336_not ; n46337
g46082 and n45657_not n45935_not ; n46338
g46083 and n45934_not n46338 ; n46339
g46084 and n46337_not n46339_not ; n46340
g46085 and b[5]_not n46340_not ; n46341
g46086 and n45675_not n45694 ; n46342
g46087 and n45690_not n46342 ; n46343
g46088 and n45691_not n45694_not ; n46344
g46089 and n46343_not n46344_not ; n46345
g46090 and n45936_not n46345_not ; n46346
g46091 and n45666_not n45935_not ; n46347
g46092 and n45934_not n46347 ; n46348
g46093 and n46346_not n46348_not ; n46349
g46094 and b[4]_not n46349_not ; n46350
g46095 and n45685_not n45689 ; n46351
g46096 and n45684_not n46351 ; n46352
g46097 and n45686_not n45689_not ; n46353
g46098 and n46352_not n46353_not ; n46354
g46099 and n45936_not n46354_not ; n46355
g46100 and n45674_not n45935_not ; n46356
g46101 and n45934_not n46356 ; n46357
g46102 and n46355_not n46357_not ; n46358
g46103 and b[3]_not n46358_not ; n46359
g46104 and n17632 n45682_not ; n46360
g46105 and n45680_not n46360 ; n46361
g46106 and n45684_not n46361_not ; n46362
g46107 and n45936_not n46362 ; n46363
g46108 and n45679_not n45935_not ; n46364
g46109 and n45934_not n46364 ; n46365
g46110 and n46363_not n46365_not ; n46366
g46111 and b[2]_not n46366_not ; n46367
g46112 and b[0] n45936_not ; n46368
g46113 and a[14] n46368_not ; n46369
g46114 and n17632 n45936_not ; n46370
g46115 and n46369_not n46370_not ; n46371
g46116 and b[1] n46371_not ; n46372
g46117 and b[1]_not n46370_not ; n46373
g46118 and n46369_not n46373 ; n46374
g46119 and n46372_not n46374_not ; n46375
g46120 and n18327_not n46375_not ; n46376
g46121 and b[1]_not n46371_not ; n46377
g46122 and n46376_not n46377_not ; n46378
g46123 and b[2] n46365_not ; n46379
g46124 and n46363_not n46379 ; n46380
g46125 and n46367_not n46380_not ; n46381
g46126 and n46378_not n46381 ; n46382
g46127 and n46367_not n46382_not ; n46383
g46128 and b[3] n46357_not ; n46384
g46129 and n46355_not n46384 ; n46385
g46130 and n46359_not n46385_not ; n46386
g46131 and n46383_not n46386 ; n46387
g46132 and n46359_not n46387_not ; n46388
g46133 and b[4] n46348_not ; n46389
g46134 and n46346_not n46389 ; n46390
g46135 and n46350_not n46390_not ; n46391
g46136 and n46388_not n46391 ; n46392
g46137 and n46350_not n46392_not ; n46393
g46138 and b[5] n46339_not ; n46394
g46139 and n46337_not n46394 ; n46395
g46140 and n46341_not n46395_not ; n46396
g46141 and n46393_not n46396 ; n46397
g46142 and n46341_not n46397_not ; n46398
g46143 and b[6] n46330_not ; n46399
g46144 and n46328_not n46399 ; n46400
g46145 and n46332_not n46400_not ; n46401
g46146 and n46398_not n46401 ; n46402
g46147 and n46332_not n46402_not ; n46403
g46148 and b[7] n46321_not ; n46404
g46149 and n46319_not n46404 ; n46405
g46150 and n46323_not n46405_not ; n46406
g46151 and n46403_not n46406 ; n46407
g46152 and n46323_not n46407_not ; n46408
g46153 and b[8] n46312_not ; n46409
g46154 and n46310_not n46409 ; n46410
g46155 and n46314_not n46410_not ; n46411
g46156 and n46408_not n46411 ; n46412
g46157 and n46314_not n46412_not ; n46413
g46158 and b[9] n46303_not ; n46414
g46159 and n46301_not n46414 ; n46415
g46160 and n46305_not n46415_not ; n46416
g46161 and n46413_not n46416 ; n46417
g46162 and n46305_not n46417_not ; n46418
g46163 and b[10] n46294_not ; n46419
g46164 and n46292_not n46419 ; n46420
g46165 and n46296_not n46420_not ; n46421
g46166 and n46418_not n46421 ; n46422
g46167 and n46296_not n46422_not ; n46423
g46168 and b[11] n46285_not ; n46424
g46169 and n46283_not n46424 ; n46425
g46170 and n46287_not n46425_not ; n46426
g46171 and n46423_not n46426 ; n46427
g46172 and n46287_not n46427_not ; n46428
g46173 and b[12] n46276_not ; n46429
g46174 and n46274_not n46429 ; n46430
g46175 and n46278_not n46430_not ; n46431
g46176 and n46428_not n46431 ; n46432
g46177 and n46278_not n46432_not ; n46433
g46178 and b[13] n46267_not ; n46434
g46179 and n46265_not n46434 ; n46435
g46180 and n46269_not n46435_not ; n46436
g46181 and n46433_not n46436 ; n46437
g46182 and n46269_not n46437_not ; n46438
g46183 and b[14] n46258_not ; n46439
g46184 and n46256_not n46439 ; n46440
g46185 and n46260_not n46440_not ; n46441
g46186 and n46438_not n46441 ; n46442
g46187 and n46260_not n46442_not ; n46443
g46188 and b[15] n46249_not ; n46444
g46189 and n46247_not n46444 ; n46445
g46190 and n46251_not n46445_not ; n46446
g46191 and n46443_not n46446 ; n46447
g46192 and n46251_not n46447_not ; n46448
g46193 and b[16] n46240_not ; n46449
g46194 and n46238_not n46449 ; n46450
g46195 and n46242_not n46450_not ; n46451
g46196 and n46448_not n46451 ; n46452
g46197 and n46242_not n46452_not ; n46453
g46198 and b[17] n46231_not ; n46454
g46199 and n46229_not n46454 ; n46455
g46200 and n46233_not n46455_not ; n46456
g46201 and n46453_not n46456 ; n46457
g46202 and n46233_not n46457_not ; n46458
g46203 and b[18] n46222_not ; n46459
g46204 and n46220_not n46459 ; n46460
g46205 and n46224_not n46460_not ; n46461
g46206 and n46458_not n46461 ; n46462
g46207 and n46224_not n46462_not ; n46463
g46208 and b[19] n46213_not ; n46464
g46209 and n46211_not n46464 ; n46465
g46210 and n46215_not n46465_not ; n46466
g46211 and n46463_not n46466 ; n46467
g46212 and n46215_not n46467_not ; n46468
g46213 and b[20] n46204_not ; n46469
g46214 and n46202_not n46469 ; n46470
g46215 and n46206_not n46470_not ; n46471
g46216 and n46468_not n46471 ; n46472
g46217 and n46206_not n46472_not ; n46473
g46218 and b[21] n46195_not ; n46474
g46219 and n46193_not n46474 ; n46475
g46220 and n46197_not n46475_not ; n46476
g46221 and n46473_not n46476 ; n46477
g46222 and n46197_not n46477_not ; n46478
g46223 and b[22] n46186_not ; n46479
g46224 and n46184_not n46479 ; n46480
g46225 and n46188_not n46480_not ; n46481
g46226 and n46478_not n46481 ; n46482
g46227 and n46188_not n46482_not ; n46483
g46228 and b[23] n46177_not ; n46484
g46229 and n46175_not n46484 ; n46485
g46230 and n46179_not n46485_not ; n46486
g46231 and n46483_not n46486 ; n46487
g46232 and n46179_not n46487_not ; n46488
g46233 and b[24] n46168_not ; n46489
g46234 and n46166_not n46489 ; n46490
g46235 and n46170_not n46490_not ; n46491
g46236 and n46488_not n46491 ; n46492
g46237 and n46170_not n46492_not ; n46493
g46238 and b[25] n46159_not ; n46494
g46239 and n46157_not n46494 ; n46495
g46240 and n46161_not n46495_not ; n46496
g46241 and n46493_not n46496 ; n46497
g46242 and n46161_not n46497_not ; n46498
g46243 and b[26] n46150_not ; n46499
g46244 and n46148_not n46499 ; n46500
g46245 and n46152_not n46500_not ; n46501
g46246 and n46498_not n46501 ; n46502
g46247 and n46152_not n46502_not ; n46503
g46248 and b[27] n46141_not ; n46504
g46249 and n46139_not n46504 ; n46505
g46250 and n46143_not n46505_not ; n46506
g46251 and n46503_not n46506 ; n46507
g46252 and n46143_not n46507_not ; n46508
g46253 and b[28] n46132_not ; n46509
g46254 and n46130_not n46509 ; n46510
g46255 and n46134_not n46510_not ; n46511
g46256 and n46508_not n46511 ; n46512
g46257 and n46134_not n46512_not ; n46513
g46258 and b[29] n46123_not ; n46514
g46259 and n46121_not n46514 ; n46515
g46260 and n46125_not n46515_not ; n46516
g46261 and n46513_not n46516 ; n46517
g46262 and n46125_not n46517_not ; n46518
g46263 and b[30] n46114_not ; n46519
g46264 and n46112_not n46519 ; n46520
g46265 and n46116_not n46520_not ; n46521
g46266 and n46518_not n46521 ; n46522
g46267 and n46116_not n46522_not ; n46523
g46268 and b[31] n46105_not ; n46524
g46269 and n46103_not n46524 ; n46525
g46270 and n46107_not n46525_not ; n46526
g46271 and n46523_not n46526 ; n46527
g46272 and n46107_not n46527_not ; n46528
g46273 and b[32] n46096_not ; n46529
g46274 and n46094_not n46529 ; n46530
g46275 and n46098_not n46530_not ; n46531
g46276 and n46528_not n46531 ; n46532
g46277 and n46098_not n46532_not ; n46533
g46278 and b[33] n46087_not ; n46534
g46279 and n46085_not n46534 ; n46535
g46280 and n46089_not n46535_not ; n46536
g46281 and n46533_not n46536 ; n46537
g46282 and n46089_not n46537_not ; n46538
g46283 and b[34] n46078_not ; n46539
g46284 and n46076_not n46539 ; n46540
g46285 and n46080_not n46540_not ; n46541
g46286 and n46538_not n46541 ; n46542
g46287 and n46080_not n46542_not ; n46543
g46288 and b[35] n46069_not ; n46544
g46289 and n46067_not n46544 ; n46545
g46290 and n46071_not n46545_not ; n46546
g46291 and n46543_not n46546 ; n46547
g46292 and n46071_not n46547_not ; n46548
g46293 and b[36] n46060_not ; n46549
g46294 and n46058_not n46549 ; n46550
g46295 and n46062_not n46550_not ; n46551
g46296 and n46548_not n46551 ; n46552
g46297 and n46062_not n46552_not ; n46553
g46298 and b[37] n46051_not ; n46554
g46299 and n46049_not n46554 ; n46555
g46300 and n46053_not n46555_not ; n46556
g46301 and n46553_not n46556 ; n46557
g46302 and n46053_not n46557_not ; n46558
g46303 and b[38] n46042_not ; n46559
g46304 and n46040_not n46559 ; n46560
g46305 and n46044_not n46560_not ; n46561
g46306 and n46558_not n46561 ; n46562
g46307 and n46044_not n46562_not ; n46563
g46308 and b[39] n46033_not ; n46564
g46309 and n46031_not n46564 ; n46565
g46310 and n46035_not n46565_not ; n46566
g46311 and n46563_not n46566 ; n46567
g46312 and n46035_not n46567_not ; n46568
g46313 and b[40] n46024_not ; n46569
g46314 and n46022_not n46569 ; n46570
g46315 and n46026_not n46570_not ; n46571
g46316 and n46568_not n46571 ; n46572
g46317 and n46026_not n46572_not ; n46573
g46318 and b[41] n46015_not ; n46574
g46319 and n46013_not n46574 ; n46575
g46320 and n46017_not n46575_not ; n46576
g46321 and n46573_not n46576 ; n46577
g46322 and n46017_not n46577_not ; n46578
g46323 and b[42] n46006_not ; n46579
g46324 and n46004_not n46579 ; n46580
g46325 and n46008_not n46580_not ; n46581
g46326 and n46578_not n46581 ; n46582
g46327 and n46008_not n46582_not ; n46583
g46328 and b[43] n45997_not ; n46584
g46329 and n45995_not n46584 ; n46585
g46330 and n45999_not n46585_not ; n46586
g46331 and n46583_not n46586 ; n46587
g46332 and n45999_not n46587_not ; n46588
g46333 and b[44] n45988_not ; n46589
g46334 and n45986_not n46589 ; n46590
g46335 and n45990_not n46590_not ; n46591
g46336 and n46588_not n46591 ; n46592
g46337 and n45990_not n46592_not ; n46593
g46338 and b[45] n45979_not ; n46594
g46339 and n45977_not n46594 ; n46595
g46340 and n45981_not n46595_not ; n46596
g46341 and n46593_not n46596 ; n46597
g46342 and n45981_not n46597_not ; n46598
g46343 and b[46] n45970_not ; n46599
g46344 and n45968_not n46599 ; n46600
g46345 and n45972_not n46600_not ; n46601
g46346 and n46598_not n46601 ; n46602
g46347 and n45972_not n46602_not ; n46603
g46348 and b[47] n45961_not ; n46604
g46349 and n45959_not n46604 ; n46605
g46350 and n45963_not n46605_not ; n46606
g46351 and n46603_not n46606 ; n46607
g46352 and n45963_not n46607_not ; n46608
g46353 and b[48] n45952_not ; n46609
g46354 and n45950_not n46609 ; n46610
g46355 and n45954_not n46610_not ; n46611
g46356 and n46608_not n46611 ; n46612
g46357 and n45954_not n46612_not ; n46613
g46358 and b[49] n45943_not ; n46614
g46359 and n45941_not n46614 ; n46615
g46360 and n45945_not n46615_not ; n46616
g46361 and n46613_not n46616 ; n46617
g46362 and n45945_not n46617_not ; n46618
g46363 and n45262_not n45931_not ; n46619
g46364 and n45929_not n46619 ; n46620
g46365 and n45920_not n46620 ; n46621
g46366 and n45929_not n45931_not ; n46622
g46367 and n45921_not n46622_not ; n46623
g46368 and n46621_not n46623_not ; n46624
g46369 and n45936_not n46624_not ; n46625
g46370 and n45928_not n45935_not ; n46626
g46371 and n45934_not n46626 ; n46627
g46372 and n46625_not n46627_not ; n46628
g46373 and b[50]_not n46628_not ; n46629
g46374 and b[50] n46627_not ; n46630
g46375 and n46625_not n46630 ; n46631
g46376 and n18585 n46631_not ; n46632
g46377 and n46629_not n46632 ; n46633
g46378 and n46618_not n46633 ; n46634
g46379 and n17882 n46628_not ; n46635
g46380 and n46634_not n46635_not ; n46636
g46381 and n45954_not n46616 ; n46637
g46382 and n46612_not n46637 ; n46638
g46383 and n46613_not n46616_not ; n46639
g46384 and n46638_not n46639_not ; n46640
g46385 and n46636_not n46640_not ; n46641
g46386 and n45944_not n46635_not ; n46642
g46387 and n46634_not n46642 ; n46643
g46388 and n46641_not n46643_not ; n46644
g46389 and n45945_not n46631_not ; n46645
g46390 and n46629_not n46645 ; n46646
g46391 and n46617_not n46646 ; n46647
g46392 and n46629_not n46631_not ; n46648
g46393 and n46618_not n46648_not ; n46649
g46394 and n46647_not n46649_not ; n46650
g46395 and n46636_not n46650_not ; n46651
g46396 and n46628_not n46635_not ; n46652
g46397 and n46634_not n46652 ; n46653
g46398 and n46651_not n46653_not ; n46654
g46399 and b[51]_not n46654_not ; n46655
g46400 and b[50]_not n46644_not ; n46656
g46401 and n45963_not n46611 ; n46657
g46402 and n46607_not n46657 ; n46658
g46403 and n46608_not n46611_not ; n46659
g46404 and n46658_not n46659_not ; n46660
g46405 and n46636_not n46660_not ; n46661
g46406 and n45953_not n46635_not ; n46662
g46407 and n46634_not n46662 ; n46663
g46408 and n46661_not n46663_not ; n46664
g46409 and b[49]_not n46664_not ; n46665
g46410 and n45972_not n46606 ; n46666
g46411 and n46602_not n46666 ; n46667
g46412 and n46603_not n46606_not ; n46668
g46413 and n46667_not n46668_not ; n46669
g46414 and n46636_not n46669_not ; n46670
g46415 and n45962_not n46635_not ; n46671
g46416 and n46634_not n46671 ; n46672
g46417 and n46670_not n46672_not ; n46673
g46418 and b[48]_not n46673_not ; n46674
g46419 and n45981_not n46601 ; n46675
g46420 and n46597_not n46675 ; n46676
g46421 and n46598_not n46601_not ; n46677
g46422 and n46676_not n46677_not ; n46678
g46423 and n46636_not n46678_not ; n46679
g46424 and n45971_not n46635_not ; n46680
g46425 and n46634_not n46680 ; n46681
g46426 and n46679_not n46681_not ; n46682
g46427 and b[47]_not n46682_not ; n46683
g46428 and n45990_not n46596 ; n46684
g46429 and n46592_not n46684 ; n46685
g46430 and n46593_not n46596_not ; n46686
g46431 and n46685_not n46686_not ; n46687
g46432 and n46636_not n46687_not ; n46688
g46433 and n45980_not n46635_not ; n46689
g46434 and n46634_not n46689 ; n46690
g46435 and n46688_not n46690_not ; n46691
g46436 and b[46]_not n46691_not ; n46692
g46437 and n45999_not n46591 ; n46693
g46438 and n46587_not n46693 ; n46694
g46439 and n46588_not n46591_not ; n46695
g46440 and n46694_not n46695_not ; n46696
g46441 and n46636_not n46696_not ; n46697
g46442 and n45989_not n46635_not ; n46698
g46443 and n46634_not n46698 ; n46699
g46444 and n46697_not n46699_not ; n46700
g46445 and b[45]_not n46700_not ; n46701
g46446 and n46008_not n46586 ; n46702
g46447 and n46582_not n46702 ; n46703
g46448 and n46583_not n46586_not ; n46704
g46449 and n46703_not n46704_not ; n46705
g46450 and n46636_not n46705_not ; n46706
g46451 and n45998_not n46635_not ; n46707
g46452 and n46634_not n46707 ; n46708
g46453 and n46706_not n46708_not ; n46709
g46454 and b[44]_not n46709_not ; n46710
g46455 and n46017_not n46581 ; n46711
g46456 and n46577_not n46711 ; n46712
g46457 and n46578_not n46581_not ; n46713
g46458 and n46712_not n46713_not ; n46714
g46459 and n46636_not n46714_not ; n46715
g46460 and n46007_not n46635_not ; n46716
g46461 and n46634_not n46716 ; n46717
g46462 and n46715_not n46717_not ; n46718
g46463 and b[43]_not n46718_not ; n46719
g46464 and n46026_not n46576 ; n46720
g46465 and n46572_not n46720 ; n46721
g46466 and n46573_not n46576_not ; n46722
g46467 and n46721_not n46722_not ; n46723
g46468 and n46636_not n46723_not ; n46724
g46469 and n46016_not n46635_not ; n46725
g46470 and n46634_not n46725 ; n46726
g46471 and n46724_not n46726_not ; n46727
g46472 and b[42]_not n46727_not ; n46728
g46473 and n46035_not n46571 ; n46729
g46474 and n46567_not n46729 ; n46730
g46475 and n46568_not n46571_not ; n46731
g46476 and n46730_not n46731_not ; n46732
g46477 and n46636_not n46732_not ; n46733
g46478 and n46025_not n46635_not ; n46734
g46479 and n46634_not n46734 ; n46735
g46480 and n46733_not n46735_not ; n46736
g46481 and b[41]_not n46736_not ; n46737
g46482 and n46044_not n46566 ; n46738
g46483 and n46562_not n46738 ; n46739
g46484 and n46563_not n46566_not ; n46740
g46485 and n46739_not n46740_not ; n46741
g46486 and n46636_not n46741_not ; n46742
g46487 and n46034_not n46635_not ; n46743
g46488 and n46634_not n46743 ; n46744
g46489 and n46742_not n46744_not ; n46745
g46490 and b[40]_not n46745_not ; n46746
g46491 and n46053_not n46561 ; n46747
g46492 and n46557_not n46747 ; n46748
g46493 and n46558_not n46561_not ; n46749
g46494 and n46748_not n46749_not ; n46750
g46495 and n46636_not n46750_not ; n46751
g46496 and n46043_not n46635_not ; n46752
g46497 and n46634_not n46752 ; n46753
g46498 and n46751_not n46753_not ; n46754
g46499 and b[39]_not n46754_not ; n46755
g46500 and n46062_not n46556 ; n46756
g46501 and n46552_not n46756 ; n46757
g46502 and n46553_not n46556_not ; n46758
g46503 and n46757_not n46758_not ; n46759
g46504 and n46636_not n46759_not ; n46760
g46505 and n46052_not n46635_not ; n46761
g46506 and n46634_not n46761 ; n46762
g46507 and n46760_not n46762_not ; n46763
g46508 and b[38]_not n46763_not ; n46764
g46509 and n46071_not n46551 ; n46765
g46510 and n46547_not n46765 ; n46766
g46511 and n46548_not n46551_not ; n46767
g46512 and n46766_not n46767_not ; n46768
g46513 and n46636_not n46768_not ; n46769
g46514 and n46061_not n46635_not ; n46770
g46515 and n46634_not n46770 ; n46771
g46516 and n46769_not n46771_not ; n46772
g46517 and b[37]_not n46772_not ; n46773
g46518 and n46080_not n46546 ; n46774
g46519 and n46542_not n46774 ; n46775
g46520 and n46543_not n46546_not ; n46776
g46521 and n46775_not n46776_not ; n46777
g46522 and n46636_not n46777_not ; n46778
g46523 and n46070_not n46635_not ; n46779
g46524 and n46634_not n46779 ; n46780
g46525 and n46778_not n46780_not ; n46781
g46526 and b[36]_not n46781_not ; n46782
g46527 and n46089_not n46541 ; n46783
g46528 and n46537_not n46783 ; n46784
g46529 and n46538_not n46541_not ; n46785
g46530 and n46784_not n46785_not ; n46786
g46531 and n46636_not n46786_not ; n46787
g46532 and n46079_not n46635_not ; n46788
g46533 and n46634_not n46788 ; n46789
g46534 and n46787_not n46789_not ; n46790
g46535 and b[35]_not n46790_not ; n46791
g46536 and n46098_not n46536 ; n46792
g46537 and n46532_not n46792 ; n46793
g46538 and n46533_not n46536_not ; n46794
g46539 and n46793_not n46794_not ; n46795
g46540 and n46636_not n46795_not ; n46796
g46541 and n46088_not n46635_not ; n46797
g46542 and n46634_not n46797 ; n46798
g46543 and n46796_not n46798_not ; n46799
g46544 and b[34]_not n46799_not ; n46800
g46545 and n46107_not n46531 ; n46801
g46546 and n46527_not n46801 ; n46802
g46547 and n46528_not n46531_not ; n46803
g46548 and n46802_not n46803_not ; n46804
g46549 and n46636_not n46804_not ; n46805
g46550 and n46097_not n46635_not ; n46806
g46551 and n46634_not n46806 ; n46807
g46552 and n46805_not n46807_not ; n46808
g46553 and b[33]_not n46808_not ; n46809
g46554 and n46116_not n46526 ; n46810
g46555 and n46522_not n46810 ; n46811
g46556 and n46523_not n46526_not ; n46812
g46557 and n46811_not n46812_not ; n46813
g46558 and n46636_not n46813_not ; n46814
g46559 and n46106_not n46635_not ; n46815
g46560 and n46634_not n46815 ; n46816
g46561 and n46814_not n46816_not ; n46817
g46562 and b[32]_not n46817_not ; n46818
g46563 and n46125_not n46521 ; n46819
g46564 and n46517_not n46819 ; n46820
g46565 and n46518_not n46521_not ; n46821
g46566 and n46820_not n46821_not ; n46822
g46567 and n46636_not n46822_not ; n46823
g46568 and n46115_not n46635_not ; n46824
g46569 and n46634_not n46824 ; n46825
g46570 and n46823_not n46825_not ; n46826
g46571 and b[31]_not n46826_not ; n46827
g46572 and n46134_not n46516 ; n46828
g46573 and n46512_not n46828 ; n46829
g46574 and n46513_not n46516_not ; n46830
g46575 and n46829_not n46830_not ; n46831
g46576 and n46636_not n46831_not ; n46832
g46577 and n46124_not n46635_not ; n46833
g46578 and n46634_not n46833 ; n46834
g46579 and n46832_not n46834_not ; n46835
g46580 and b[30]_not n46835_not ; n46836
g46581 and n46143_not n46511 ; n46837
g46582 and n46507_not n46837 ; n46838
g46583 and n46508_not n46511_not ; n46839
g46584 and n46838_not n46839_not ; n46840
g46585 and n46636_not n46840_not ; n46841
g46586 and n46133_not n46635_not ; n46842
g46587 and n46634_not n46842 ; n46843
g46588 and n46841_not n46843_not ; n46844
g46589 and b[29]_not n46844_not ; n46845
g46590 and n46152_not n46506 ; n46846
g46591 and n46502_not n46846 ; n46847
g46592 and n46503_not n46506_not ; n46848
g46593 and n46847_not n46848_not ; n46849
g46594 and n46636_not n46849_not ; n46850
g46595 and n46142_not n46635_not ; n46851
g46596 and n46634_not n46851 ; n46852
g46597 and n46850_not n46852_not ; n46853
g46598 and b[28]_not n46853_not ; n46854
g46599 and n46161_not n46501 ; n46855
g46600 and n46497_not n46855 ; n46856
g46601 and n46498_not n46501_not ; n46857
g46602 and n46856_not n46857_not ; n46858
g46603 and n46636_not n46858_not ; n46859
g46604 and n46151_not n46635_not ; n46860
g46605 and n46634_not n46860 ; n46861
g46606 and n46859_not n46861_not ; n46862
g46607 and b[27]_not n46862_not ; n46863
g46608 and n46170_not n46496 ; n46864
g46609 and n46492_not n46864 ; n46865
g46610 and n46493_not n46496_not ; n46866
g46611 and n46865_not n46866_not ; n46867
g46612 and n46636_not n46867_not ; n46868
g46613 and n46160_not n46635_not ; n46869
g46614 and n46634_not n46869 ; n46870
g46615 and n46868_not n46870_not ; n46871
g46616 and b[26]_not n46871_not ; n46872
g46617 and n46179_not n46491 ; n46873
g46618 and n46487_not n46873 ; n46874
g46619 and n46488_not n46491_not ; n46875
g46620 and n46874_not n46875_not ; n46876
g46621 and n46636_not n46876_not ; n46877
g46622 and n46169_not n46635_not ; n46878
g46623 and n46634_not n46878 ; n46879
g46624 and n46877_not n46879_not ; n46880
g46625 and b[25]_not n46880_not ; n46881
g46626 and n46188_not n46486 ; n46882
g46627 and n46482_not n46882 ; n46883
g46628 and n46483_not n46486_not ; n46884
g46629 and n46883_not n46884_not ; n46885
g46630 and n46636_not n46885_not ; n46886
g46631 and n46178_not n46635_not ; n46887
g46632 and n46634_not n46887 ; n46888
g46633 and n46886_not n46888_not ; n46889
g46634 and b[24]_not n46889_not ; n46890
g46635 and n46197_not n46481 ; n46891
g46636 and n46477_not n46891 ; n46892
g46637 and n46478_not n46481_not ; n46893
g46638 and n46892_not n46893_not ; n46894
g46639 and n46636_not n46894_not ; n46895
g46640 and n46187_not n46635_not ; n46896
g46641 and n46634_not n46896 ; n46897
g46642 and n46895_not n46897_not ; n46898
g46643 and b[23]_not n46898_not ; n46899
g46644 and n46206_not n46476 ; n46900
g46645 and n46472_not n46900 ; n46901
g46646 and n46473_not n46476_not ; n46902
g46647 and n46901_not n46902_not ; n46903
g46648 and n46636_not n46903_not ; n46904
g46649 and n46196_not n46635_not ; n46905
g46650 and n46634_not n46905 ; n46906
g46651 and n46904_not n46906_not ; n46907
g46652 and b[22]_not n46907_not ; n46908
g46653 and n46215_not n46471 ; n46909
g46654 and n46467_not n46909 ; n46910
g46655 and n46468_not n46471_not ; n46911
g46656 and n46910_not n46911_not ; n46912
g46657 and n46636_not n46912_not ; n46913
g46658 and n46205_not n46635_not ; n46914
g46659 and n46634_not n46914 ; n46915
g46660 and n46913_not n46915_not ; n46916
g46661 and b[21]_not n46916_not ; n46917
g46662 and n46224_not n46466 ; n46918
g46663 and n46462_not n46918 ; n46919
g46664 and n46463_not n46466_not ; n46920
g46665 and n46919_not n46920_not ; n46921
g46666 and n46636_not n46921_not ; n46922
g46667 and n46214_not n46635_not ; n46923
g46668 and n46634_not n46923 ; n46924
g46669 and n46922_not n46924_not ; n46925
g46670 and b[20]_not n46925_not ; n46926
g46671 and n46233_not n46461 ; n46927
g46672 and n46457_not n46927 ; n46928
g46673 and n46458_not n46461_not ; n46929
g46674 and n46928_not n46929_not ; n46930
g46675 and n46636_not n46930_not ; n46931
g46676 and n46223_not n46635_not ; n46932
g46677 and n46634_not n46932 ; n46933
g46678 and n46931_not n46933_not ; n46934
g46679 and b[19]_not n46934_not ; n46935
g46680 and n46242_not n46456 ; n46936
g46681 and n46452_not n46936 ; n46937
g46682 and n46453_not n46456_not ; n46938
g46683 and n46937_not n46938_not ; n46939
g46684 and n46636_not n46939_not ; n46940
g46685 and n46232_not n46635_not ; n46941
g46686 and n46634_not n46941 ; n46942
g46687 and n46940_not n46942_not ; n46943
g46688 and b[18]_not n46943_not ; n46944
g46689 and n46251_not n46451 ; n46945
g46690 and n46447_not n46945 ; n46946
g46691 and n46448_not n46451_not ; n46947
g46692 and n46946_not n46947_not ; n46948
g46693 and n46636_not n46948_not ; n46949
g46694 and n46241_not n46635_not ; n46950
g46695 and n46634_not n46950 ; n46951
g46696 and n46949_not n46951_not ; n46952
g46697 and b[17]_not n46952_not ; n46953
g46698 and n46260_not n46446 ; n46954
g46699 and n46442_not n46954 ; n46955
g46700 and n46443_not n46446_not ; n46956
g46701 and n46955_not n46956_not ; n46957
g46702 and n46636_not n46957_not ; n46958
g46703 and n46250_not n46635_not ; n46959
g46704 and n46634_not n46959 ; n46960
g46705 and n46958_not n46960_not ; n46961
g46706 and b[16]_not n46961_not ; n46962
g46707 and n46269_not n46441 ; n46963
g46708 and n46437_not n46963 ; n46964
g46709 and n46438_not n46441_not ; n46965
g46710 and n46964_not n46965_not ; n46966
g46711 and n46636_not n46966_not ; n46967
g46712 and n46259_not n46635_not ; n46968
g46713 and n46634_not n46968 ; n46969
g46714 and n46967_not n46969_not ; n46970
g46715 and b[15]_not n46970_not ; n46971
g46716 and n46278_not n46436 ; n46972
g46717 and n46432_not n46972 ; n46973
g46718 and n46433_not n46436_not ; n46974
g46719 and n46973_not n46974_not ; n46975
g46720 and n46636_not n46975_not ; n46976
g46721 and n46268_not n46635_not ; n46977
g46722 and n46634_not n46977 ; n46978
g46723 and n46976_not n46978_not ; n46979
g46724 and b[14]_not n46979_not ; n46980
g46725 and n46287_not n46431 ; n46981
g46726 and n46427_not n46981 ; n46982
g46727 and n46428_not n46431_not ; n46983
g46728 and n46982_not n46983_not ; n46984
g46729 and n46636_not n46984_not ; n46985
g46730 and n46277_not n46635_not ; n46986
g46731 and n46634_not n46986 ; n46987
g46732 and n46985_not n46987_not ; n46988
g46733 and b[13]_not n46988_not ; n46989
g46734 and n46296_not n46426 ; n46990
g46735 and n46422_not n46990 ; n46991
g46736 and n46423_not n46426_not ; n46992
g46737 and n46991_not n46992_not ; n46993
g46738 and n46636_not n46993_not ; n46994
g46739 and n46286_not n46635_not ; n46995
g46740 and n46634_not n46995 ; n46996
g46741 and n46994_not n46996_not ; n46997
g46742 and b[12]_not n46997_not ; n46998
g46743 and n46305_not n46421 ; n46999
g46744 and n46417_not n46999 ; n47000
g46745 and n46418_not n46421_not ; n47001
g46746 and n47000_not n47001_not ; n47002
g46747 and n46636_not n47002_not ; n47003
g46748 and n46295_not n46635_not ; n47004
g46749 and n46634_not n47004 ; n47005
g46750 and n47003_not n47005_not ; n47006
g46751 and b[11]_not n47006_not ; n47007
g46752 and n46314_not n46416 ; n47008
g46753 and n46412_not n47008 ; n47009
g46754 and n46413_not n46416_not ; n47010
g46755 and n47009_not n47010_not ; n47011
g46756 and n46636_not n47011_not ; n47012
g46757 and n46304_not n46635_not ; n47013
g46758 and n46634_not n47013 ; n47014
g46759 and n47012_not n47014_not ; n47015
g46760 and b[10]_not n47015_not ; n47016
g46761 and n46323_not n46411 ; n47017
g46762 and n46407_not n47017 ; n47018
g46763 and n46408_not n46411_not ; n47019
g46764 and n47018_not n47019_not ; n47020
g46765 and n46636_not n47020_not ; n47021
g46766 and n46313_not n46635_not ; n47022
g46767 and n46634_not n47022 ; n47023
g46768 and n47021_not n47023_not ; n47024
g46769 and b[9]_not n47024_not ; n47025
g46770 and n46332_not n46406 ; n47026
g46771 and n46402_not n47026 ; n47027
g46772 and n46403_not n46406_not ; n47028
g46773 and n47027_not n47028_not ; n47029
g46774 and n46636_not n47029_not ; n47030
g46775 and n46322_not n46635_not ; n47031
g46776 and n46634_not n47031 ; n47032
g46777 and n47030_not n47032_not ; n47033
g46778 and b[8]_not n47033_not ; n47034
g46779 and n46341_not n46401 ; n47035
g46780 and n46397_not n47035 ; n47036
g46781 and n46398_not n46401_not ; n47037
g46782 and n47036_not n47037_not ; n47038
g46783 and n46636_not n47038_not ; n47039
g46784 and n46331_not n46635_not ; n47040
g46785 and n46634_not n47040 ; n47041
g46786 and n47039_not n47041_not ; n47042
g46787 and b[7]_not n47042_not ; n47043
g46788 and n46350_not n46396 ; n47044
g46789 and n46392_not n47044 ; n47045
g46790 and n46393_not n46396_not ; n47046
g46791 and n47045_not n47046_not ; n47047
g46792 and n46636_not n47047_not ; n47048
g46793 and n46340_not n46635_not ; n47049
g46794 and n46634_not n47049 ; n47050
g46795 and n47048_not n47050_not ; n47051
g46796 and b[6]_not n47051_not ; n47052
g46797 and n46359_not n46391 ; n47053
g46798 and n46387_not n47053 ; n47054
g46799 and n46388_not n46391_not ; n47055
g46800 and n47054_not n47055_not ; n47056
g46801 and n46636_not n47056_not ; n47057
g46802 and n46349_not n46635_not ; n47058
g46803 and n46634_not n47058 ; n47059
g46804 and n47057_not n47059_not ; n47060
g46805 and b[5]_not n47060_not ; n47061
g46806 and n46367_not n46386 ; n47062
g46807 and n46382_not n47062 ; n47063
g46808 and n46383_not n46386_not ; n47064
g46809 and n47063_not n47064_not ; n47065
g46810 and n46636_not n47065_not ; n47066
g46811 and n46358_not n46635_not ; n47067
g46812 and n46634_not n47067 ; n47068
g46813 and n47066_not n47068_not ; n47069
g46814 and b[4]_not n47069_not ; n47070
g46815 and n46377_not n46381 ; n47071
g46816 and n46376_not n47071 ; n47072
g46817 and n46378_not n46381_not ; n47073
g46818 and n47072_not n47073_not ; n47074
g46819 and n46636_not n47074_not ; n47075
g46820 and n46366_not n46635_not ; n47076
g46821 and n46634_not n47076 ; n47077
g46822 and n47075_not n47077_not ; n47078
g46823 and b[3]_not n47078_not ; n47079
g46824 and n18327 n46374_not ; n47080
g46825 and n46372_not n47080 ; n47081
g46826 and n46376_not n47081_not ; n47082
g46827 and n46636_not n47082 ; n47083
g46828 and n46371_not n46635_not ; n47084
g46829 and n46634_not n47084 ; n47085
g46830 and n47083_not n47085_not ; n47086
g46831 and b[2]_not n47086_not ; n47087
g46832 and b[0] n46636_not ; n47088
g46833 and a[13] n47088_not ; n47089
g46834 and n18327 n46636_not ; n47090
g46835 and n47089_not n47090_not ; n47091
g46836 and b[1] n47091_not ; n47092
g46837 and b[1]_not n47090_not ; n47093
g46838 and n47089_not n47093 ; n47094
g46839 and n47092_not n47094_not ; n47095
g46840 and n19050_not n47095_not ; n47096
g46841 and b[1]_not n47091_not ; n47097
g46842 and n47096_not n47097_not ; n47098
g46843 and b[2] n47085_not ; n47099
g46844 and n47083_not n47099 ; n47100
g46845 and n47087_not n47100_not ; n47101
g46846 and n47098_not n47101 ; n47102
g46847 and n47087_not n47102_not ; n47103
g46848 and b[3] n47077_not ; n47104
g46849 and n47075_not n47104 ; n47105
g46850 and n47079_not n47105_not ; n47106
g46851 and n47103_not n47106 ; n47107
g46852 and n47079_not n47107_not ; n47108
g46853 and b[4] n47068_not ; n47109
g46854 and n47066_not n47109 ; n47110
g46855 and n47070_not n47110_not ; n47111
g46856 and n47108_not n47111 ; n47112
g46857 and n47070_not n47112_not ; n47113
g46858 and b[5] n47059_not ; n47114
g46859 and n47057_not n47114 ; n47115
g46860 and n47061_not n47115_not ; n47116
g46861 and n47113_not n47116 ; n47117
g46862 and n47061_not n47117_not ; n47118
g46863 and b[6] n47050_not ; n47119
g46864 and n47048_not n47119 ; n47120
g46865 and n47052_not n47120_not ; n47121
g46866 and n47118_not n47121 ; n47122
g46867 and n47052_not n47122_not ; n47123
g46868 and b[7] n47041_not ; n47124
g46869 and n47039_not n47124 ; n47125
g46870 and n47043_not n47125_not ; n47126
g46871 and n47123_not n47126 ; n47127
g46872 and n47043_not n47127_not ; n47128
g46873 and b[8] n47032_not ; n47129
g46874 and n47030_not n47129 ; n47130
g46875 and n47034_not n47130_not ; n47131
g46876 and n47128_not n47131 ; n47132
g46877 and n47034_not n47132_not ; n47133
g46878 and b[9] n47023_not ; n47134
g46879 and n47021_not n47134 ; n47135
g46880 and n47025_not n47135_not ; n47136
g46881 and n47133_not n47136 ; n47137
g46882 and n47025_not n47137_not ; n47138
g46883 and b[10] n47014_not ; n47139
g46884 and n47012_not n47139 ; n47140
g46885 and n47016_not n47140_not ; n47141
g46886 and n47138_not n47141 ; n47142
g46887 and n47016_not n47142_not ; n47143
g46888 and b[11] n47005_not ; n47144
g46889 and n47003_not n47144 ; n47145
g46890 and n47007_not n47145_not ; n47146
g46891 and n47143_not n47146 ; n47147
g46892 and n47007_not n47147_not ; n47148
g46893 and b[12] n46996_not ; n47149
g46894 and n46994_not n47149 ; n47150
g46895 and n46998_not n47150_not ; n47151
g46896 and n47148_not n47151 ; n47152
g46897 and n46998_not n47152_not ; n47153
g46898 and b[13] n46987_not ; n47154
g46899 and n46985_not n47154 ; n47155
g46900 and n46989_not n47155_not ; n47156
g46901 and n47153_not n47156 ; n47157
g46902 and n46989_not n47157_not ; n47158
g46903 and b[14] n46978_not ; n47159
g46904 and n46976_not n47159 ; n47160
g46905 and n46980_not n47160_not ; n47161
g46906 and n47158_not n47161 ; n47162
g46907 and n46980_not n47162_not ; n47163
g46908 and b[15] n46969_not ; n47164
g46909 and n46967_not n47164 ; n47165
g46910 and n46971_not n47165_not ; n47166
g46911 and n47163_not n47166 ; n47167
g46912 and n46971_not n47167_not ; n47168
g46913 and b[16] n46960_not ; n47169
g46914 and n46958_not n47169 ; n47170
g46915 and n46962_not n47170_not ; n47171
g46916 and n47168_not n47171 ; n47172
g46917 and n46962_not n47172_not ; n47173
g46918 and b[17] n46951_not ; n47174
g46919 and n46949_not n47174 ; n47175
g46920 and n46953_not n47175_not ; n47176
g46921 and n47173_not n47176 ; n47177
g46922 and n46953_not n47177_not ; n47178
g46923 and b[18] n46942_not ; n47179
g46924 and n46940_not n47179 ; n47180
g46925 and n46944_not n47180_not ; n47181
g46926 and n47178_not n47181 ; n47182
g46927 and n46944_not n47182_not ; n47183
g46928 and b[19] n46933_not ; n47184
g46929 and n46931_not n47184 ; n47185
g46930 and n46935_not n47185_not ; n47186
g46931 and n47183_not n47186 ; n47187
g46932 and n46935_not n47187_not ; n47188
g46933 and b[20] n46924_not ; n47189
g46934 and n46922_not n47189 ; n47190
g46935 and n46926_not n47190_not ; n47191
g46936 and n47188_not n47191 ; n47192
g46937 and n46926_not n47192_not ; n47193
g46938 and b[21] n46915_not ; n47194
g46939 and n46913_not n47194 ; n47195
g46940 and n46917_not n47195_not ; n47196
g46941 and n47193_not n47196 ; n47197
g46942 and n46917_not n47197_not ; n47198
g46943 and b[22] n46906_not ; n47199
g46944 and n46904_not n47199 ; n47200
g46945 and n46908_not n47200_not ; n47201
g46946 and n47198_not n47201 ; n47202
g46947 and n46908_not n47202_not ; n47203
g46948 and b[23] n46897_not ; n47204
g46949 and n46895_not n47204 ; n47205
g46950 and n46899_not n47205_not ; n47206
g46951 and n47203_not n47206 ; n47207
g46952 and n46899_not n47207_not ; n47208
g46953 and b[24] n46888_not ; n47209
g46954 and n46886_not n47209 ; n47210
g46955 and n46890_not n47210_not ; n47211
g46956 and n47208_not n47211 ; n47212
g46957 and n46890_not n47212_not ; n47213
g46958 and b[25] n46879_not ; n47214
g46959 and n46877_not n47214 ; n47215
g46960 and n46881_not n47215_not ; n47216
g46961 and n47213_not n47216 ; n47217
g46962 and n46881_not n47217_not ; n47218
g46963 and b[26] n46870_not ; n47219
g46964 and n46868_not n47219 ; n47220
g46965 and n46872_not n47220_not ; n47221
g46966 and n47218_not n47221 ; n47222
g46967 and n46872_not n47222_not ; n47223
g46968 and b[27] n46861_not ; n47224
g46969 and n46859_not n47224 ; n47225
g46970 and n46863_not n47225_not ; n47226
g46971 and n47223_not n47226 ; n47227
g46972 and n46863_not n47227_not ; n47228
g46973 and b[28] n46852_not ; n47229
g46974 and n46850_not n47229 ; n47230
g46975 and n46854_not n47230_not ; n47231
g46976 and n47228_not n47231 ; n47232
g46977 and n46854_not n47232_not ; n47233
g46978 and b[29] n46843_not ; n47234
g46979 and n46841_not n47234 ; n47235
g46980 and n46845_not n47235_not ; n47236
g46981 and n47233_not n47236 ; n47237
g46982 and n46845_not n47237_not ; n47238
g46983 and b[30] n46834_not ; n47239
g46984 and n46832_not n47239 ; n47240
g46985 and n46836_not n47240_not ; n47241
g46986 and n47238_not n47241 ; n47242
g46987 and n46836_not n47242_not ; n47243
g46988 and b[31] n46825_not ; n47244
g46989 and n46823_not n47244 ; n47245
g46990 and n46827_not n47245_not ; n47246
g46991 and n47243_not n47246 ; n47247
g46992 and n46827_not n47247_not ; n47248
g46993 and b[32] n46816_not ; n47249
g46994 and n46814_not n47249 ; n47250
g46995 and n46818_not n47250_not ; n47251
g46996 and n47248_not n47251 ; n47252
g46997 and n46818_not n47252_not ; n47253
g46998 and b[33] n46807_not ; n47254
g46999 and n46805_not n47254 ; n47255
g47000 and n46809_not n47255_not ; n47256
g47001 and n47253_not n47256 ; n47257
g47002 and n46809_not n47257_not ; n47258
g47003 and b[34] n46798_not ; n47259
g47004 and n46796_not n47259 ; n47260
g47005 and n46800_not n47260_not ; n47261
g47006 and n47258_not n47261 ; n47262
g47007 and n46800_not n47262_not ; n47263
g47008 and b[35] n46789_not ; n47264
g47009 and n46787_not n47264 ; n47265
g47010 and n46791_not n47265_not ; n47266
g47011 and n47263_not n47266 ; n47267
g47012 and n46791_not n47267_not ; n47268
g47013 and b[36] n46780_not ; n47269
g47014 and n46778_not n47269 ; n47270
g47015 and n46782_not n47270_not ; n47271
g47016 and n47268_not n47271 ; n47272
g47017 and n46782_not n47272_not ; n47273
g47018 and b[37] n46771_not ; n47274
g47019 and n46769_not n47274 ; n47275
g47020 and n46773_not n47275_not ; n47276
g47021 and n47273_not n47276 ; n47277
g47022 and n46773_not n47277_not ; n47278
g47023 and b[38] n46762_not ; n47279
g47024 and n46760_not n47279 ; n47280
g47025 and n46764_not n47280_not ; n47281
g47026 and n47278_not n47281 ; n47282
g47027 and n46764_not n47282_not ; n47283
g47028 and b[39] n46753_not ; n47284
g47029 and n46751_not n47284 ; n47285
g47030 and n46755_not n47285_not ; n47286
g47031 and n47283_not n47286 ; n47287
g47032 and n46755_not n47287_not ; n47288
g47033 and b[40] n46744_not ; n47289
g47034 and n46742_not n47289 ; n47290
g47035 and n46746_not n47290_not ; n47291
g47036 and n47288_not n47291 ; n47292
g47037 and n46746_not n47292_not ; n47293
g47038 and b[41] n46735_not ; n47294
g47039 and n46733_not n47294 ; n47295
g47040 and n46737_not n47295_not ; n47296
g47041 and n47293_not n47296 ; n47297
g47042 and n46737_not n47297_not ; n47298
g47043 and b[42] n46726_not ; n47299
g47044 and n46724_not n47299 ; n47300
g47045 and n46728_not n47300_not ; n47301
g47046 and n47298_not n47301 ; n47302
g47047 and n46728_not n47302_not ; n47303
g47048 and b[43] n46717_not ; n47304
g47049 and n46715_not n47304 ; n47305
g47050 and n46719_not n47305_not ; n47306
g47051 and n47303_not n47306 ; n47307
g47052 and n46719_not n47307_not ; n47308
g47053 and b[44] n46708_not ; n47309
g47054 and n46706_not n47309 ; n47310
g47055 and n46710_not n47310_not ; n47311
g47056 and n47308_not n47311 ; n47312
g47057 and n46710_not n47312_not ; n47313
g47058 and b[45] n46699_not ; n47314
g47059 and n46697_not n47314 ; n47315
g47060 and n46701_not n47315_not ; n47316
g47061 and n47313_not n47316 ; n47317
g47062 and n46701_not n47317_not ; n47318
g47063 and b[46] n46690_not ; n47319
g47064 and n46688_not n47319 ; n47320
g47065 and n46692_not n47320_not ; n47321
g47066 and n47318_not n47321 ; n47322
g47067 and n46692_not n47322_not ; n47323
g47068 and b[47] n46681_not ; n47324
g47069 and n46679_not n47324 ; n47325
g47070 and n46683_not n47325_not ; n47326
g47071 and n47323_not n47326 ; n47327
g47072 and n46683_not n47327_not ; n47328
g47073 and b[48] n46672_not ; n47329
g47074 and n46670_not n47329 ; n47330
g47075 and n46674_not n47330_not ; n47331
g47076 and n47328_not n47331 ; n47332
g47077 and n46674_not n47332_not ; n47333
g47078 and b[49] n46663_not ; n47334
g47079 and n46661_not n47334 ; n47335
g47080 and n46665_not n47335_not ; n47336
g47081 and n47333_not n47336 ; n47337
g47082 and n46665_not n47337_not ; n47338
g47083 and b[50] n46643_not ; n47339
g47084 and n46641_not n47339 ; n47340
g47085 and n46656_not n47340_not ; n47341
g47086 and n47338_not n47341 ; n47342
g47087 and n46656_not n47342_not ; n47343
g47088 and b[51] n46653_not ; n47344
g47089 and n46651_not n47344 ; n47345
g47090 and n46655_not n47345_not ; n47346
g47091 and n47343_not n47346 ; n47347
g47092 and n46655_not n47347_not ; n47348
g47093 and n288 n47348_not ; n47349
g47094 and n46644_not n47349_not ; n47350
g47095 and n46665_not n47341 ; n47351
g47096 and n47337_not n47351 ; n47352
g47097 and n47338_not n47341_not ; n47353
g47098 and n47352_not n47353_not ; n47354
g47099 and n288 n47354_not ; n47355
g47100 and n47348_not n47355 ; n47356
g47101 and n47350_not n47356_not ; n47357
g47102 and b[51]_not n47357_not ; n47358
g47103 and n46664_not n47349_not ; n47359
g47104 and n46674_not n47336 ; n47360
g47105 and n47332_not n47360 ; n47361
g47106 and n47333_not n47336_not ; n47362
g47107 and n47361_not n47362_not ; n47363
g47108 and n288 n47363_not ; n47364
g47109 and n47348_not n47364 ; n47365
g47110 and n47359_not n47365_not ; n47366
g47111 and b[50]_not n47366_not ; n47367
g47112 and n46673_not n47349_not ; n47368
g47113 and n46683_not n47331 ; n47369
g47114 and n47327_not n47369 ; n47370
g47115 and n47328_not n47331_not ; n47371
g47116 and n47370_not n47371_not ; n47372
g47117 and n288 n47372_not ; n47373
g47118 and n47348_not n47373 ; n47374
g47119 and n47368_not n47374_not ; n47375
g47120 and b[49]_not n47375_not ; n47376
g47121 and n46682_not n47349_not ; n47377
g47122 and n46692_not n47326 ; n47378
g47123 and n47322_not n47378 ; n47379
g47124 and n47323_not n47326_not ; n47380
g47125 and n47379_not n47380_not ; n47381
g47126 and n288 n47381_not ; n47382
g47127 and n47348_not n47382 ; n47383
g47128 and n47377_not n47383_not ; n47384
g47129 and b[48]_not n47384_not ; n47385
g47130 and n46691_not n47349_not ; n47386
g47131 and n46701_not n47321 ; n47387
g47132 and n47317_not n47387 ; n47388
g47133 and n47318_not n47321_not ; n47389
g47134 and n47388_not n47389_not ; n47390
g47135 and n288 n47390_not ; n47391
g47136 and n47348_not n47391 ; n47392
g47137 and n47386_not n47392_not ; n47393
g47138 and b[47]_not n47393_not ; n47394
g47139 and n46700_not n47349_not ; n47395
g47140 and n46710_not n47316 ; n47396
g47141 and n47312_not n47396 ; n47397
g47142 and n47313_not n47316_not ; n47398
g47143 and n47397_not n47398_not ; n47399
g47144 and n288 n47399_not ; n47400
g47145 and n47348_not n47400 ; n47401
g47146 and n47395_not n47401_not ; n47402
g47147 and b[46]_not n47402_not ; n47403
g47148 and n46709_not n47349_not ; n47404
g47149 and n46719_not n47311 ; n47405
g47150 and n47307_not n47405 ; n47406
g47151 and n47308_not n47311_not ; n47407
g47152 and n47406_not n47407_not ; n47408
g47153 and n288 n47408_not ; n47409
g47154 and n47348_not n47409 ; n47410
g47155 and n47404_not n47410_not ; n47411
g47156 and b[45]_not n47411_not ; n47412
g47157 and n46718_not n47349_not ; n47413
g47158 and n46728_not n47306 ; n47414
g47159 and n47302_not n47414 ; n47415
g47160 and n47303_not n47306_not ; n47416
g47161 and n47415_not n47416_not ; n47417
g47162 and n288 n47417_not ; n47418
g47163 and n47348_not n47418 ; n47419
g47164 and n47413_not n47419_not ; n47420
g47165 and b[44]_not n47420_not ; n47421
g47166 and n46727_not n47349_not ; n47422
g47167 and n46737_not n47301 ; n47423
g47168 and n47297_not n47423 ; n47424
g47169 and n47298_not n47301_not ; n47425
g47170 and n47424_not n47425_not ; n47426
g47171 and n288 n47426_not ; n47427
g47172 and n47348_not n47427 ; n47428
g47173 and n47422_not n47428_not ; n47429
g47174 and b[43]_not n47429_not ; n47430
g47175 and n46736_not n47349_not ; n47431
g47176 and n46746_not n47296 ; n47432
g47177 and n47292_not n47432 ; n47433
g47178 and n47293_not n47296_not ; n47434
g47179 and n47433_not n47434_not ; n47435
g47180 and n288 n47435_not ; n47436
g47181 and n47348_not n47436 ; n47437
g47182 and n47431_not n47437_not ; n47438
g47183 and b[42]_not n47438_not ; n47439
g47184 and n46745_not n47349_not ; n47440
g47185 and n46755_not n47291 ; n47441
g47186 and n47287_not n47441 ; n47442
g47187 and n47288_not n47291_not ; n47443
g47188 and n47442_not n47443_not ; n47444
g47189 and n288 n47444_not ; n47445
g47190 and n47348_not n47445 ; n47446
g47191 and n47440_not n47446_not ; n47447
g47192 and b[41]_not n47447_not ; n47448
g47193 and n46754_not n47349_not ; n47449
g47194 and n46764_not n47286 ; n47450
g47195 and n47282_not n47450 ; n47451
g47196 and n47283_not n47286_not ; n47452
g47197 and n47451_not n47452_not ; n47453
g47198 and n288 n47453_not ; n47454
g47199 and n47348_not n47454 ; n47455
g47200 and n47449_not n47455_not ; n47456
g47201 and b[40]_not n47456_not ; n47457
g47202 and n46763_not n47349_not ; n47458
g47203 and n46773_not n47281 ; n47459
g47204 and n47277_not n47459 ; n47460
g47205 and n47278_not n47281_not ; n47461
g47206 and n47460_not n47461_not ; n47462
g47207 and n288 n47462_not ; n47463
g47208 and n47348_not n47463 ; n47464
g47209 and n47458_not n47464_not ; n47465
g47210 and b[39]_not n47465_not ; n47466
g47211 and n46772_not n47349_not ; n47467
g47212 and n46782_not n47276 ; n47468
g47213 and n47272_not n47468 ; n47469
g47214 and n47273_not n47276_not ; n47470
g47215 and n47469_not n47470_not ; n47471
g47216 and n288 n47471_not ; n47472
g47217 and n47348_not n47472 ; n47473
g47218 and n47467_not n47473_not ; n47474
g47219 and b[38]_not n47474_not ; n47475
g47220 and n46781_not n47349_not ; n47476
g47221 and n46791_not n47271 ; n47477
g47222 and n47267_not n47477 ; n47478
g47223 and n47268_not n47271_not ; n47479
g47224 and n47478_not n47479_not ; n47480
g47225 and n288 n47480_not ; n47481
g47226 and n47348_not n47481 ; n47482
g47227 and n47476_not n47482_not ; n47483
g47228 and b[37]_not n47483_not ; n47484
g47229 and n46790_not n47349_not ; n47485
g47230 and n46800_not n47266 ; n47486
g47231 and n47262_not n47486 ; n47487
g47232 and n47263_not n47266_not ; n47488
g47233 and n47487_not n47488_not ; n47489
g47234 and n288 n47489_not ; n47490
g47235 and n47348_not n47490 ; n47491
g47236 and n47485_not n47491_not ; n47492
g47237 and b[36]_not n47492_not ; n47493
g47238 and n46799_not n47349_not ; n47494
g47239 and n46809_not n47261 ; n47495
g47240 and n47257_not n47495 ; n47496
g47241 and n47258_not n47261_not ; n47497
g47242 and n47496_not n47497_not ; n47498
g47243 and n288 n47498_not ; n47499
g47244 and n47348_not n47499 ; n47500
g47245 and n47494_not n47500_not ; n47501
g47246 and b[35]_not n47501_not ; n47502
g47247 and n46808_not n47349_not ; n47503
g47248 and n46818_not n47256 ; n47504
g47249 and n47252_not n47504 ; n47505
g47250 and n47253_not n47256_not ; n47506
g47251 and n47505_not n47506_not ; n47507
g47252 and n288 n47507_not ; n47508
g47253 and n47348_not n47508 ; n47509
g47254 and n47503_not n47509_not ; n47510
g47255 and b[34]_not n47510_not ; n47511
g47256 and n46817_not n47349_not ; n47512
g47257 and n46827_not n47251 ; n47513
g47258 and n47247_not n47513 ; n47514
g47259 and n47248_not n47251_not ; n47515
g47260 and n47514_not n47515_not ; n47516
g47261 and n288 n47516_not ; n47517
g47262 and n47348_not n47517 ; n47518
g47263 and n47512_not n47518_not ; n47519
g47264 and b[33]_not n47519_not ; n47520
g47265 and n46826_not n47349_not ; n47521
g47266 and n46836_not n47246 ; n47522
g47267 and n47242_not n47522 ; n47523
g47268 and n47243_not n47246_not ; n47524
g47269 and n47523_not n47524_not ; n47525
g47270 and n288 n47525_not ; n47526
g47271 and n47348_not n47526 ; n47527
g47272 and n47521_not n47527_not ; n47528
g47273 and b[32]_not n47528_not ; n47529
g47274 and n46835_not n47349_not ; n47530
g47275 and n46845_not n47241 ; n47531
g47276 and n47237_not n47531 ; n47532
g47277 and n47238_not n47241_not ; n47533
g47278 and n47532_not n47533_not ; n47534
g47279 and n288 n47534_not ; n47535
g47280 and n47348_not n47535 ; n47536
g47281 and n47530_not n47536_not ; n47537
g47282 and b[31]_not n47537_not ; n47538
g47283 and n46844_not n47349_not ; n47539
g47284 and n46854_not n47236 ; n47540
g47285 and n47232_not n47540 ; n47541
g47286 and n47233_not n47236_not ; n47542
g47287 and n47541_not n47542_not ; n47543
g47288 and n288 n47543_not ; n47544
g47289 and n47348_not n47544 ; n47545
g47290 and n47539_not n47545_not ; n47546
g47291 and b[30]_not n47546_not ; n47547
g47292 and n46853_not n47349_not ; n47548
g47293 and n46863_not n47231 ; n47549
g47294 and n47227_not n47549 ; n47550
g47295 and n47228_not n47231_not ; n47551
g47296 and n47550_not n47551_not ; n47552
g47297 and n288 n47552_not ; n47553
g47298 and n47348_not n47553 ; n47554
g47299 and n47548_not n47554_not ; n47555
g47300 and b[29]_not n47555_not ; n47556
g47301 and n46862_not n47349_not ; n47557
g47302 and n46872_not n47226 ; n47558
g47303 and n47222_not n47558 ; n47559
g47304 and n47223_not n47226_not ; n47560
g47305 and n47559_not n47560_not ; n47561
g47306 and n288 n47561_not ; n47562
g47307 and n47348_not n47562 ; n47563
g47308 and n47557_not n47563_not ; n47564
g47309 and b[28]_not n47564_not ; n47565
g47310 and n46871_not n47349_not ; n47566
g47311 and n46881_not n47221 ; n47567
g47312 and n47217_not n47567 ; n47568
g47313 and n47218_not n47221_not ; n47569
g47314 and n47568_not n47569_not ; n47570
g47315 and n288 n47570_not ; n47571
g47316 and n47348_not n47571 ; n47572
g47317 and n47566_not n47572_not ; n47573
g47318 and b[27]_not n47573_not ; n47574
g47319 and n46880_not n47349_not ; n47575
g47320 and n46890_not n47216 ; n47576
g47321 and n47212_not n47576 ; n47577
g47322 and n47213_not n47216_not ; n47578
g47323 and n47577_not n47578_not ; n47579
g47324 and n288 n47579_not ; n47580
g47325 and n47348_not n47580 ; n47581
g47326 and n47575_not n47581_not ; n47582
g47327 and b[26]_not n47582_not ; n47583
g47328 and n46889_not n47349_not ; n47584
g47329 and n46899_not n47211 ; n47585
g47330 and n47207_not n47585 ; n47586
g47331 and n47208_not n47211_not ; n47587
g47332 and n47586_not n47587_not ; n47588
g47333 and n288 n47588_not ; n47589
g47334 and n47348_not n47589 ; n47590
g47335 and n47584_not n47590_not ; n47591
g47336 and b[25]_not n47591_not ; n47592
g47337 and n46898_not n47349_not ; n47593
g47338 and n46908_not n47206 ; n47594
g47339 and n47202_not n47594 ; n47595
g47340 and n47203_not n47206_not ; n47596
g47341 and n47595_not n47596_not ; n47597
g47342 and n288 n47597_not ; n47598
g47343 and n47348_not n47598 ; n47599
g47344 and n47593_not n47599_not ; n47600
g47345 and b[24]_not n47600_not ; n47601
g47346 and n46907_not n47349_not ; n47602
g47347 and n46917_not n47201 ; n47603
g47348 and n47197_not n47603 ; n47604
g47349 and n47198_not n47201_not ; n47605
g47350 and n47604_not n47605_not ; n47606
g47351 and n288 n47606_not ; n47607
g47352 and n47348_not n47607 ; n47608
g47353 and n47602_not n47608_not ; n47609
g47354 and b[23]_not n47609_not ; n47610
g47355 and n46916_not n47349_not ; n47611
g47356 and n46926_not n47196 ; n47612
g47357 and n47192_not n47612 ; n47613
g47358 and n47193_not n47196_not ; n47614
g47359 and n47613_not n47614_not ; n47615
g47360 and n288 n47615_not ; n47616
g47361 and n47348_not n47616 ; n47617
g47362 and n47611_not n47617_not ; n47618
g47363 and b[22]_not n47618_not ; n47619
g47364 and n46925_not n47349_not ; n47620
g47365 and n46935_not n47191 ; n47621
g47366 and n47187_not n47621 ; n47622
g47367 and n47188_not n47191_not ; n47623
g47368 and n47622_not n47623_not ; n47624
g47369 and n288 n47624_not ; n47625
g47370 and n47348_not n47625 ; n47626
g47371 and n47620_not n47626_not ; n47627
g47372 and b[21]_not n47627_not ; n47628
g47373 and n46934_not n47349_not ; n47629
g47374 and n46944_not n47186 ; n47630
g47375 and n47182_not n47630 ; n47631
g47376 and n47183_not n47186_not ; n47632
g47377 and n47631_not n47632_not ; n47633
g47378 and n288 n47633_not ; n47634
g47379 and n47348_not n47634 ; n47635
g47380 and n47629_not n47635_not ; n47636
g47381 and b[20]_not n47636_not ; n47637
g47382 and n46943_not n47349_not ; n47638
g47383 and n46953_not n47181 ; n47639
g47384 and n47177_not n47639 ; n47640
g47385 and n47178_not n47181_not ; n47641
g47386 and n47640_not n47641_not ; n47642
g47387 and n288 n47642_not ; n47643
g47388 and n47348_not n47643 ; n47644
g47389 and n47638_not n47644_not ; n47645
g47390 and b[19]_not n47645_not ; n47646
g47391 and n46952_not n47349_not ; n47647
g47392 and n46962_not n47176 ; n47648
g47393 and n47172_not n47648 ; n47649
g47394 and n47173_not n47176_not ; n47650
g47395 and n47649_not n47650_not ; n47651
g47396 and n288 n47651_not ; n47652
g47397 and n47348_not n47652 ; n47653
g47398 and n47647_not n47653_not ; n47654
g47399 and b[18]_not n47654_not ; n47655
g47400 and n46961_not n47349_not ; n47656
g47401 and n46971_not n47171 ; n47657
g47402 and n47167_not n47657 ; n47658
g47403 and n47168_not n47171_not ; n47659
g47404 and n47658_not n47659_not ; n47660
g47405 and n288 n47660_not ; n47661
g47406 and n47348_not n47661 ; n47662
g47407 and n47656_not n47662_not ; n47663
g47408 and b[17]_not n47663_not ; n47664
g47409 and n46970_not n47349_not ; n47665
g47410 and n46980_not n47166 ; n47666
g47411 and n47162_not n47666 ; n47667
g47412 and n47163_not n47166_not ; n47668
g47413 and n47667_not n47668_not ; n47669
g47414 and n288 n47669_not ; n47670
g47415 and n47348_not n47670 ; n47671
g47416 and n47665_not n47671_not ; n47672
g47417 and b[16]_not n47672_not ; n47673
g47418 and n46979_not n47349_not ; n47674
g47419 and n46989_not n47161 ; n47675
g47420 and n47157_not n47675 ; n47676
g47421 and n47158_not n47161_not ; n47677
g47422 and n47676_not n47677_not ; n47678
g47423 and n288 n47678_not ; n47679
g47424 and n47348_not n47679 ; n47680
g47425 and n47674_not n47680_not ; n47681
g47426 and b[15]_not n47681_not ; n47682
g47427 and n46988_not n47349_not ; n47683
g47428 and n46998_not n47156 ; n47684
g47429 and n47152_not n47684 ; n47685
g47430 and n47153_not n47156_not ; n47686
g47431 and n47685_not n47686_not ; n47687
g47432 and n288 n47687_not ; n47688
g47433 and n47348_not n47688 ; n47689
g47434 and n47683_not n47689_not ; n47690
g47435 and b[14]_not n47690_not ; n47691
g47436 and n46997_not n47349_not ; n47692
g47437 and n47007_not n47151 ; n47693
g47438 and n47147_not n47693 ; n47694
g47439 and n47148_not n47151_not ; n47695
g47440 and n47694_not n47695_not ; n47696
g47441 and n288 n47696_not ; n47697
g47442 and n47348_not n47697 ; n47698
g47443 and n47692_not n47698_not ; n47699
g47444 and b[13]_not n47699_not ; n47700
g47445 and n47006_not n47349_not ; n47701
g47446 and n47016_not n47146 ; n47702
g47447 and n47142_not n47702 ; n47703
g47448 and n47143_not n47146_not ; n47704
g47449 and n47703_not n47704_not ; n47705
g47450 and n288 n47705_not ; n47706
g47451 and n47348_not n47706 ; n47707
g47452 and n47701_not n47707_not ; n47708
g47453 and b[12]_not n47708_not ; n47709
g47454 and n47015_not n47349_not ; n47710
g47455 and n47025_not n47141 ; n47711
g47456 and n47137_not n47711 ; n47712
g47457 and n47138_not n47141_not ; n47713
g47458 and n47712_not n47713_not ; n47714
g47459 and n288 n47714_not ; n47715
g47460 and n47348_not n47715 ; n47716
g47461 and n47710_not n47716_not ; n47717
g47462 and b[11]_not n47717_not ; n47718
g47463 and n47024_not n47349_not ; n47719
g47464 and n47034_not n47136 ; n47720
g47465 and n47132_not n47720 ; n47721
g47466 and n47133_not n47136_not ; n47722
g47467 and n47721_not n47722_not ; n47723
g47468 and n288 n47723_not ; n47724
g47469 and n47348_not n47724 ; n47725
g47470 and n47719_not n47725_not ; n47726
g47471 and b[10]_not n47726_not ; n47727
g47472 and n47033_not n47349_not ; n47728
g47473 and n47043_not n47131 ; n47729
g47474 and n47127_not n47729 ; n47730
g47475 and n47128_not n47131_not ; n47731
g47476 and n47730_not n47731_not ; n47732
g47477 and n288 n47732_not ; n47733
g47478 and n47348_not n47733 ; n47734
g47479 and n47728_not n47734_not ; n47735
g47480 and b[9]_not n47735_not ; n47736
g47481 and n47042_not n47349_not ; n47737
g47482 and n47052_not n47126 ; n47738
g47483 and n47122_not n47738 ; n47739
g47484 and n47123_not n47126_not ; n47740
g47485 and n47739_not n47740_not ; n47741
g47486 and n288 n47741_not ; n47742
g47487 and n47348_not n47742 ; n47743
g47488 and n47737_not n47743_not ; n47744
g47489 and b[8]_not n47744_not ; n47745
g47490 and n47051_not n47349_not ; n47746
g47491 and n47061_not n47121 ; n47747
g47492 and n47117_not n47747 ; n47748
g47493 and n47118_not n47121_not ; n47749
g47494 and n47748_not n47749_not ; n47750
g47495 and n288 n47750_not ; n47751
g47496 and n47348_not n47751 ; n47752
g47497 and n47746_not n47752_not ; n47753
g47498 and b[7]_not n47753_not ; n47754
g47499 and n47060_not n47349_not ; n47755
g47500 and n47070_not n47116 ; n47756
g47501 and n47112_not n47756 ; n47757
g47502 and n47113_not n47116_not ; n47758
g47503 and n47757_not n47758_not ; n47759
g47504 and n288 n47759_not ; n47760
g47505 and n47348_not n47760 ; n47761
g47506 and n47755_not n47761_not ; n47762
g47507 and b[6]_not n47762_not ; n47763
g47508 and n47069_not n47349_not ; n47764
g47509 and n47079_not n47111 ; n47765
g47510 and n47107_not n47765 ; n47766
g47511 and n47108_not n47111_not ; n47767
g47512 and n47766_not n47767_not ; n47768
g47513 and n288 n47768_not ; n47769
g47514 and n47348_not n47769 ; n47770
g47515 and n47764_not n47770_not ; n47771
g47516 and b[5]_not n47771_not ; n47772
g47517 and n47078_not n47349_not ; n47773
g47518 and n47087_not n47106 ; n47774
g47519 and n47102_not n47774 ; n47775
g47520 and n47103_not n47106_not ; n47776
g47521 and n47775_not n47776_not ; n47777
g47522 and n288 n47777_not ; n47778
g47523 and n47348_not n47778 ; n47779
g47524 and n47773_not n47779_not ; n47780
g47525 and b[4]_not n47780_not ; n47781
g47526 and n47086_not n47349_not ; n47782
g47527 and n47097_not n47101 ; n47783
g47528 and n47096_not n47783 ; n47784
g47529 and n47098_not n47101_not ; n47785
g47530 and n47784_not n47785_not ; n47786
g47531 and n288 n47786_not ; n47787
g47532 and n47348_not n47787 ; n47788
g47533 and n47782_not n47788_not ; n47789
g47534 and b[3]_not n47789_not ; n47790
g47535 and n47091_not n47349_not ; n47791
g47536 and n19050 n47094_not ; n47792
g47537 and n47092_not n47792 ; n47793
g47538 and n288 n47793_not ; n47794
g47539 and n47096_not n47794 ; n47795
g47540 and n47348_not n47795 ; n47796
g47541 and n47791_not n47796_not ; n47797
g47542 and b[2]_not n47797_not ; n47798
g47543 and n19756 n47348_not ; n47799
g47544 and a[12] n47799_not ; n47800
g47545 and n19760 n47348_not ; n47801
g47546 and n47800_not n47801_not ; n47802
g47547 and b[1] n47802_not ; n47803
g47548 and b[1]_not n47801_not ; n47804
g47549 and n47800_not n47804 ; n47805
g47550 and n47803_not n47805_not ; n47806
g47551 and n19767_not n47806_not ; n47807
g47552 and b[1]_not n47802_not ; n47808
g47553 and n47807_not n47808_not ; n47809
g47554 and b[2] n47796_not ; n47810
g47555 and n47791_not n47810 ; n47811
g47556 and n47798_not n47811_not ; n47812
g47557 and n47809_not n47812 ; n47813
g47558 and n47798_not n47813_not ; n47814
g47559 and b[3] n47788_not ; n47815
g47560 and n47782_not n47815 ; n47816
g47561 and n47790_not n47816_not ; n47817
g47562 and n47814_not n47817 ; n47818
g47563 and n47790_not n47818_not ; n47819
g47564 and b[4] n47779_not ; n47820
g47565 and n47773_not n47820 ; n47821
g47566 and n47781_not n47821_not ; n47822
g47567 and n47819_not n47822 ; n47823
g47568 and n47781_not n47823_not ; n47824
g47569 and b[5] n47770_not ; n47825
g47570 and n47764_not n47825 ; n47826
g47571 and n47772_not n47826_not ; n47827
g47572 and n47824_not n47827 ; n47828
g47573 and n47772_not n47828_not ; n47829
g47574 and b[6] n47761_not ; n47830
g47575 and n47755_not n47830 ; n47831
g47576 and n47763_not n47831_not ; n47832
g47577 and n47829_not n47832 ; n47833
g47578 and n47763_not n47833_not ; n47834
g47579 and b[7] n47752_not ; n47835
g47580 and n47746_not n47835 ; n47836
g47581 and n47754_not n47836_not ; n47837
g47582 and n47834_not n47837 ; n47838
g47583 and n47754_not n47838_not ; n47839
g47584 and b[8] n47743_not ; n47840
g47585 and n47737_not n47840 ; n47841
g47586 and n47745_not n47841_not ; n47842
g47587 and n47839_not n47842 ; n47843
g47588 and n47745_not n47843_not ; n47844
g47589 and b[9] n47734_not ; n47845
g47590 and n47728_not n47845 ; n47846
g47591 and n47736_not n47846_not ; n47847
g47592 and n47844_not n47847 ; n47848
g47593 and n47736_not n47848_not ; n47849
g47594 and b[10] n47725_not ; n47850
g47595 and n47719_not n47850 ; n47851
g47596 and n47727_not n47851_not ; n47852
g47597 and n47849_not n47852 ; n47853
g47598 and n47727_not n47853_not ; n47854
g47599 and b[11] n47716_not ; n47855
g47600 and n47710_not n47855 ; n47856
g47601 and n47718_not n47856_not ; n47857
g47602 and n47854_not n47857 ; n47858
g47603 and n47718_not n47858_not ; n47859
g47604 and b[12] n47707_not ; n47860
g47605 and n47701_not n47860 ; n47861
g47606 and n47709_not n47861_not ; n47862
g47607 and n47859_not n47862 ; n47863
g47608 and n47709_not n47863_not ; n47864
g47609 and b[13] n47698_not ; n47865
g47610 and n47692_not n47865 ; n47866
g47611 and n47700_not n47866_not ; n47867
g47612 and n47864_not n47867 ; n47868
g47613 and n47700_not n47868_not ; n47869
g47614 and b[14] n47689_not ; n47870
g47615 and n47683_not n47870 ; n47871
g47616 and n47691_not n47871_not ; n47872
g47617 and n47869_not n47872 ; n47873
g47618 and n47691_not n47873_not ; n47874
g47619 and b[15] n47680_not ; n47875
g47620 and n47674_not n47875 ; n47876
g47621 and n47682_not n47876_not ; n47877
g47622 and n47874_not n47877 ; n47878
g47623 and n47682_not n47878_not ; n47879
g47624 and b[16] n47671_not ; n47880
g47625 and n47665_not n47880 ; n47881
g47626 and n47673_not n47881_not ; n47882
g47627 and n47879_not n47882 ; n47883
g47628 and n47673_not n47883_not ; n47884
g47629 and b[17] n47662_not ; n47885
g47630 and n47656_not n47885 ; n47886
g47631 and n47664_not n47886_not ; n47887
g47632 and n47884_not n47887 ; n47888
g47633 and n47664_not n47888_not ; n47889
g47634 and b[18] n47653_not ; n47890
g47635 and n47647_not n47890 ; n47891
g47636 and n47655_not n47891_not ; n47892
g47637 and n47889_not n47892 ; n47893
g47638 and n47655_not n47893_not ; n47894
g47639 and b[19] n47644_not ; n47895
g47640 and n47638_not n47895 ; n47896
g47641 and n47646_not n47896_not ; n47897
g47642 and n47894_not n47897 ; n47898
g47643 and n47646_not n47898_not ; n47899
g47644 and b[20] n47635_not ; n47900
g47645 and n47629_not n47900 ; n47901
g47646 and n47637_not n47901_not ; n47902
g47647 and n47899_not n47902 ; n47903
g47648 and n47637_not n47903_not ; n47904
g47649 and b[21] n47626_not ; n47905
g47650 and n47620_not n47905 ; n47906
g47651 and n47628_not n47906_not ; n47907
g47652 and n47904_not n47907 ; n47908
g47653 and n47628_not n47908_not ; n47909
g47654 and b[22] n47617_not ; n47910
g47655 and n47611_not n47910 ; n47911
g47656 and n47619_not n47911_not ; n47912
g47657 and n47909_not n47912 ; n47913
g47658 and n47619_not n47913_not ; n47914
g47659 and b[23] n47608_not ; n47915
g47660 and n47602_not n47915 ; n47916
g47661 and n47610_not n47916_not ; n47917
g47662 and n47914_not n47917 ; n47918
g47663 and n47610_not n47918_not ; n47919
g47664 and b[24] n47599_not ; n47920
g47665 and n47593_not n47920 ; n47921
g47666 and n47601_not n47921_not ; n47922
g47667 and n47919_not n47922 ; n47923
g47668 and n47601_not n47923_not ; n47924
g47669 and b[25] n47590_not ; n47925
g47670 and n47584_not n47925 ; n47926
g47671 and n47592_not n47926_not ; n47927
g47672 and n47924_not n47927 ; n47928
g47673 and n47592_not n47928_not ; n47929
g47674 and b[26] n47581_not ; n47930
g47675 and n47575_not n47930 ; n47931
g47676 and n47583_not n47931_not ; n47932
g47677 and n47929_not n47932 ; n47933
g47678 and n47583_not n47933_not ; n47934
g47679 and b[27] n47572_not ; n47935
g47680 and n47566_not n47935 ; n47936
g47681 and n47574_not n47936_not ; n47937
g47682 and n47934_not n47937 ; n47938
g47683 and n47574_not n47938_not ; n47939
g47684 and b[28] n47563_not ; n47940
g47685 and n47557_not n47940 ; n47941
g47686 and n47565_not n47941_not ; n47942
g47687 and n47939_not n47942 ; n47943
g47688 and n47565_not n47943_not ; n47944
g47689 and b[29] n47554_not ; n47945
g47690 and n47548_not n47945 ; n47946
g47691 and n47556_not n47946_not ; n47947
g47692 and n47944_not n47947 ; n47948
g47693 and n47556_not n47948_not ; n47949
g47694 and b[30] n47545_not ; n47950
g47695 and n47539_not n47950 ; n47951
g47696 and n47547_not n47951_not ; n47952
g47697 and n47949_not n47952 ; n47953
g47698 and n47547_not n47953_not ; n47954
g47699 and b[31] n47536_not ; n47955
g47700 and n47530_not n47955 ; n47956
g47701 and n47538_not n47956_not ; n47957
g47702 and n47954_not n47957 ; n47958
g47703 and n47538_not n47958_not ; n47959
g47704 and b[32] n47527_not ; n47960
g47705 and n47521_not n47960 ; n47961
g47706 and n47529_not n47961_not ; n47962
g47707 and n47959_not n47962 ; n47963
g47708 and n47529_not n47963_not ; n47964
g47709 and b[33] n47518_not ; n47965
g47710 and n47512_not n47965 ; n47966
g47711 and n47520_not n47966_not ; n47967
g47712 and n47964_not n47967 ; n47968
g47713 and n47520_not n47968_not ; n47969
g47714 and b[34] n47509_not ; n47970
g47715 and n47503_not n47970 ; n47971
g47716 and n47511_not n47971_not ; n47972
g47717 and n47969_not n47972 ; n47973
g47718 and n47511_not n47973_not ; n47974
g47719 and b[35] n47500_not ; n47975
g47720 and n47494_not n47975 ; n47976
g47721 and n47502_not n47976_not ; n47977
g47722 and n47974_not n47977 ; n47978
g47723 and n47502_not n47978_not ; n47979
g47724 and b[36] n47491_not ; n47980
g47725 and n47485_not n47980 ; n47981
g47726 and n47493_not n47981_not ; n47982
g47727 and n47979_not n47982 ; n47983
g47728 and n47493_not n47983_not ; n47984
g47729 and b[37] n47482_not ; n47985
g47730 and n47476_not n47985 ; n47986
g47731 and n47484_not n47986_not ; n47987
g47732 and n47984_not n47987 ; n47988
g47733 and n47484_not n47988_not ; n47989
g47734 and b[38] n47473_not ; n47990
g47735 and n47467_not n47990 ; n47991
g47736 and n47475_not n47991_not ; n47992
g47737 and n47989_not n47992 ; n47993
g47738 and n47475_not n47993_not ; n47994
g47739 and b[39] n47464_not ; n47995
g47740 and n47458_not n47995 ; n47996
g47741 and n47466_not n47996_not ; n47997
g47742 and n47994_not n47997 ; n47998
g47743 and n47466_not n47998_not ; n47999
g47744 and b[40] n47455_not ; n48000
g47745 and n47449_not n48000 ; n48001
g47746 and n47457_not n48001_not ; n48002
g47747 and n47999_not n48002 ; n48003
g47748 and n47457_not n48003_not ; n48004
g47749 and b[41] n47446_not ; n48005
g47750 and n47440_not n48005 ; n48006
g47751 and n47448_not n48006_not ; n48007
g47752 and n48004_not n48007 ; n48008
g47753 and n47448_not n48008_not ; n48009
g47754 and b[42] n47437_not ; n48010
g47755 and n47431_not n48010 ; n48011
g47756 and n47439_not n48011_not ; n48012
g47757 and n48009_not n48012 ; n48013
g47758 and n47439_not n48013_not ; n48014
g47759 and b[43] n47428_not ; n48015
g47760 and n47422_not n48015 ; n48016
g47761 and n47430_not n48016_not ; n48017
g47762 and n48014_not n48017 ; n48018
g47763 and n47430_not n48018_not ; n48019
g47764 and b[44] n47419_not ; n48020
g47765 and n47413_not n48020 ; n48021
g47766 and n47421_not n48021_not ; n48022
g47767 and n48019_not n48022 ; n48023
g47768 and n47421_not n48023_not ; n48024
g47769 and b[45] n47410_not ; n48025
g47770 and n47404_not n48025 ; n48026
g47771 and n47412_not n48026_not ; n48027
g47772 and n48024_not n48027 ; n48028
g47773 and n47412_not n48028_not ; n48029
g47774 and b[46] n47401_not ; n48030
g47775 and n47395_not n48030 ; n48031
g47776 and n47403_not n48031_not ; n48032
g47777 and n48029_not n48032 ; n48033
g47778 and n47403_not n48033_not ; n48034
g47779 and b[47] n47392_not ; n48035
g47780 and n47386_not n48035 ; n48036
g47781 and n47394_not n48036_not ; n48037
g47782 and n48034_not n48037 ; n48038
g47783 and n47394_not n48038_not ; n48039
g47784 and b[48] n47383_not ; n48040
g47785 and n47377_not n48040 ; n48041
g47786 and n47385_not n48041_not ; n48042
g47787 and n48039_not n48042 ; n48043
g47788 and n47385_not n48043_not ; n48044
g47789 and b[49] n47374_not ; n48045
g47790 and n47368_not n48045 ; n48046
g47791 and n47376_not n48046_not ; n48047
g47792 and n48044_not n48047 ; n48048
g47793 and n47376_not n48048_not ; n48049
g47794 and b[50] n47365_not ; n48050
g47795 and n47359_not n48050 ; n48051
g47796 and n47367_not n48051_not ; n48052
g47797 and n48049_not n48052 ; n48053
g47798 and n47367_not n48053_not ; n48054
g47799 and b[51] n47356_not ; n48055
g47800 and n47350_not n48055 ; n48056
g47801 and n47358_not n48056_not ; n48057
g47802 and n48054_not n48057 ; n48058
g47803 and n47358_not n48058_not ; n48059
g47804 and n46654_not n47349_not ; n48060
g47805 and n46656_not n47346 ; n48061
g47806 and n47342_not n48061 ; n48062
g47807 and n47343_not n47346_not ; n48063
g47808 and n48062_not n48063_not ; n48064
g47809 and n47349 n48064_not ; n48065
g47810 and n48060_not n48065_not ; n48066
g47811 and b[52]_not n48066_not ; n48067
g47812 and b[52] n48060_not ; n48068
g47813 and n48065_not n48068 ; n48069
g47814 and n595 n48069_not ; n48070
g47815 and n48067_not n48070 ; n48071
g47816 and n48059_not n48071 ; n48072
g47817 and n288 n48066_not ; n48073
g47818 and n48072_not n48073_not ; n48074
g47819 and n47367_not n48057 ; n48075
g47820 and n48053_not n48075 ; n48076
g47821 and n48054_not n48057_not ; n48077
g47822 and n48076_not n48077_not ; n48078
g47823 and n48074_not n48078_not ; n48079
g47824 and n47357_not n48073_not ; n48080
g47825 and n48072_not n48080 ; n48081
g47826 and n48079_not n48081_not ; n48082
g47827 and b[52]_not n48082_not ; n48083
g47828 and n47376_not n48052 ; n48084
g47829 and n48048_not n48084 ; n48085
g47830 and n48049_not n48052_not ; n48086
g47831 and n48085_not n48086_not ; n48087
g47832 and n48074_not n48087_not ; n48088
g47833 and n47366_not n48073_not ; n48089
g47834 and n48072_not n48089 ; n48090
g47835 and n48088_not n48090_not ; n48091
g47836 and b[51]_not n48091_not ; n48092
g47837 and n47385_not n48047 ; n48093
g47838 and n48043_not n48093 ; n48094
g47839 and n48044_not n48047_not ; n48095
g47840 and n48094_not n48095_not ; n48096
g47841 and n48074_not n48096_not ; n48097
g47842 and n47375_not n48073_not ; n48098
g47843 and n48072_not n48098 ; n48099
g47844 and n48097_not n48099_not ; n48100
g47845 and b[50]_not n48100_not ; n48101
g47846 and n47394_not n48042 ; n48102
g47847 and n48038_not n48102 ; n48103
g47848 and n48039_not n48042_not ; n48104
g47849 and n48103_not n48104_not ; n48105
g47850 and n48074_not n48105_not ; n48106
g47851 and n47384_not n48073_not ; n48107
g47852 and n48072_not n48107 ; n48108
g47853 and n48106_not n48108_not ; n48109
g47854 and b[49]_not n48109_not ; n48110
g47855 and n47403_not n48037 ; n48111
g47856 and n48033_not n48111 ; n48112
g47857 and n48034_not n48037_not ; n48113
g47858 and n48112_not n48113_not ; n48114
g47859 and n48074_not n48114_not ; n48115
g47860 and n47393_not n48073_not ; n48116
g47861 and n48072_not n48116 ; n48117
g47862 and n48115_not n48117_not ; n48118
g47863 and b[48]_not n48118_not ; n48119
g47864 and n47412_not n48032 ; n48120
g47865 and n48028_not n48120 ; n48121
g47866 and n48029_not n48032_not ; n48122
g47867 and n48121_not n48122_not ; n48123
g47868 and n48074_not n48123_not ; n48124
g47869 and n47402_not n48073_not ; n48125
g47870 and n48072_not n48125 ; n48126
g47871 and n48124_not n48126_not ; n48127
g47872 and b[47]_not n48127_not ; n48128
g47873 and n47421_not n48027 ; n48129
g47874 and n48023_not n48129 ; n48130
g47875 and n48024_not n48027_not ; n48131
g47876 and n48130_not n48131_not ; n48132
g47877 and n48074_not n48132_not ; n48133
g47878 and n47411_not n48073_not ; n48134
g47879 and n48072_not n48134 ; n48135
g47880 and n48133_not n48135_not ; n48136
g47881 and b[46]_not n48136_not ; n48137
g47882 and n47430_not n48022 ; n48138
g47883 and n48018_not n48138 ; n48139
g47884 and n48019_not n48022_not ; n48140
g47885 and n48139_not n48140_not ; n48141
g47886 and n48074_not n48141_not ; n48142
g47887 and n47420_not n48073_not ; n48143
g47888 and n48072_not n48143 ; n48144
g47889 and n48142_not n48144_not ; n48145
g47890 and b[45]_not n48145_not ; n48146
g47891 and n47439_not n48017 ; n48147
g47892 and n48013_not n48147 ; n48148
g47893 and n48014_not n48017_not ; n48149
g47894 and n48148_not n48149_not ; n48150
g47895 and n48074_not n48150_not ; n48151
g47896 and n47429_not n48073_not ; n48152
g47897 and n48072_not n48152 ; n48153
g47898 and n48151_not n48153_not ; n48154
g47899 and b[44]_not n48154_not ; n48155
g47900 and n47448_not n48012 ; n48156
g47901 and n48008_not n48156 ; n48157
g47902 and n48009_not n48012_not ; n48158
g47903 and n48157_not n48158_not ; n48159
g47904 and n48074_not n48159_not ; n48160
g47905 and n47438_not n48073_not ; n48161
g47906 and n48072_not n48161 ; n48162
g47907 and n48160_not n48162_not ; n48163
g47908 and b[43]_not n48163_not ; n48164
g47909 and n47457_not n48007 ; n48165
g47910 and n48003_not n48165 ; n48166
g47911 and n48004_not n48007_not ; n48167
g47912 and n48166_not n48167_not ; n48168
g47913 and n48074_not n48168_not ; n48169
g47914 and n47447_not n48073_not ; n48170
g47915 and n48072_not n48170 ; n48171
g47916 and n48169_not n48171_not ; n48172
g47917 and b[42]_not n48172_not ; n48173
g47918 and n47466_not n48002 ; n48174
g47919 and n47998_not n48174 ; n48175
g47920 and n47999_not n48002_not ; n48176
g47921 and n48175_not n48176_not ; n48177
g47922 and n48074_not n48177_not ; n48178
g47923 and n47456_not n48073_not ; n48179
g47924 and n48072_not n48179 ; n48180
g47925 and n48178_not n48180_not ; n48181
g47926 and b[41]_not n48181_not ; n48182
g47927 and n47475_not n47997 ; n48183
g47928 and n47993_not n48183 ; n48184
g47929 and n47994_not n47997_not ; n48185
g47930 and n48184_not n48185_not ; n48186
g47931 and n48074_not n48186_not ; n48187
g47932 and n47465_not n48073_not ; n48188
g47933 and n48072_not n48188 ; n48189
g47934 and n48187_not n48189_not ; n48190
g47935 and b[40]_not n48190_not ; n48191
g47936 and n47484_not n47992 ; n48192
g47937 and n47988_not n48192 ; n48193
g47938 and n47989_not n47992_not ; n48194
g47939 and n48193_not n48194_not ; n48195
g47940 and n48074_not n48195_not ; n48196
g47941 and n47474_not n48073_not ; n48197
g47942 and n48072_not n48197 ; n48198
g47943 and n48196_not n48198_not ; n48199
g47944 and b[39]_not n48199_not ; n48200
g47945 and n47493_not n47987 ; n48201
g47946 and n47983_not n48201 ; n48202
g47947 and n47984_not n47987_not ; n48203
g47948 and n48202_not n48203_not ; n48204
g47949 and n48074_not n48204_not ; n48205
g47950 and n47483_not n48073_not ; n48206
g47951 and n48072_not n48206 ; n48207
g47952 and n48205_not n48207_not ; n48208
g47953 and b[38]_not n48208_not ; n48209
g47954 and n47502_not n47982 ; n48210
g47955 and n47978_not n48210 ; n48211
g47956 and n47979_not n47982_not ; n48212
g47957 and n48211_not n48212_not ; n48213
g47958 and n48074_not n48213_not ; n48214
g47959 and n47492_not n48073_not ; n48215
g47960 and n48072_not n48215 ; n48216
g47961 and n48214_not n48216_not ; n48217
g47962 and b[37]_not n48217_not ; n48218
g47963 and n47511_not n47977 ; n48219
g47964 and n47973_not n48219 ; n48220
g47965 and n47974_not n47977_not ; n48221
g47966 and n48220_not n48221_not ; n48222
g47967 and n48074_not n48222_not ; n48223
g47968 and n47501_not n48073_not ; n48224
g47969 and n48072_not n48224 ; n48225
g47970 and n48223_not n48225_not ; n48226
g47971 and b[36]_not n48226_not ; n48227
g47972 and n47520_not n47972 ; n48228
g47973 and n47968_not n48228 ; n48229
g47974 and n47969_not n47972_not ; n48230
g47975 and n48229_not n48230_not ; n48231
g47976 and n48074_not n48231_not ; n48232
g47977 and n47510_not n48073_not ; n48233
g47978 and n48072_not n48233 ; n48234
g47979 and n48232_not n48234_not ; n48235
g47980 and b[35]_not n48235_not ; n48236
g47981 and n47529_not n47967 ; n48237
g47982 and n47963_not n48237 ; n48238
g47983 and n47964_not n47967_not ; n48239
g47984 and n48238_not n48239_not ; n48240
g47985 and n48074_not n48240_not ; n48241
g47986 and n47519_not n48073_not ; n48242
g47987 and n48072_not n48242 ; n48243
g47988 and n48241_not n48243_not ; n48244
g47989 and b[34]_not n48244_not ; n48245
g47990 and n47538_not n47962 ; n48246
g47991 and n47958_not n48246 ; n48247
g47992 and n47959_not n47962_not ; n48248
g47993 and n48247_not n48248_not ; n48249
g47994 and n48074_not n48249_not ; n48250
g47995 and n47528_not n48073_not ; n48251
g47996 and n48072_not n48251 ; n48252
g47997 and n48250_not n48252_not ; n48253
g47998 and b[33]_not n48253_not ; n48254
g47999 and n47547_not n47957 ; n48255
g48000 and n47953_not n48255 ; n48256
g48001 and n47954_not n47957_not ; n48257
g48002 and n48256_not n48257_not ; n48258
g48003 and n48074_not n48258_not ; n48259
g48004 and n47537_not n48073_not ; n48260
g48005 and n48072_not n48260 ; n48261
g48006 and n48259_not n48261_not ; n48262
g48007 and b[32]_not n48262_not ; n48263
g48008 and n47556_not n47952 ; n48264
g48009 and n47948_not n48264 ; n48265
g48010 and n47949_not n47952_not ; n48266
g48011 and n48265_not n48266_not ; n48267
g48012 and n48074_not n48267_not ; n48268
g48013 and n47546_not n48073_not ; n48269
g48014 and n48072_not n48269 ; n48270
g48015 and n48268_not n48270_not ; n48271
g48016 and b[31]_not n48271_not ; n48272
g48017 and n47565_not n47947 ; n48273
g48018 and n47943_not n48273 ; n48274
g48019 and n47944_not n47947_not ; n48275
g48020 and n48274_not n48275_not ; n48276
g48021 and n48074_not n48276_not ; n48277
g48022 and n47555_not n48073_not ; n48278
g48023 and n48072_not n48278 ; n48279
g48024 and n48277_not n48279_not ; n48280
g48025 and b[30]_not n48280_not ; n48281
g48026 and n47574_not n47942 ; n48282
g48027 and n47938_not n48282 ; n48283
g48028 and n47939_not n47942_not ; n48284
g48029 and n48283_not n48284_not ; n48285
g48030 and n48074_not n48285_not ; n48286
g48031 and n47564_not n48073_not ; n48287
g48032 and n48072_not n48287 ; n48288
g48033 and n48286_not n48288_not ; n48289
g48034 and b[29]_not n48289_not ; n48290
g48035 and n47583_not n47937 ; n48291
g48036 and n47933_not n48291 ; n48292
g48037 and n47934_not n47937_not ; n48293
g48038 and n48292_not n48293_not ; n48294
g48039 and n48074_not n48294_not ; n48295
g48040 and n47573_not n48073_not ; n48296
g48041 and n48072_not n48296 ; n48297
g48042 and n48295_not n48297_not ; n48298
g48043 and b[28]_not n48298_not ; n48299
g48044 and n47592_not n47932 ; n48300
g48045 and n47928_not n48300 ; n48301
g48046 and n47929_not n47932_not ; n48302
g48047 and n48301_not n48302_not ; n48303
g48048 and n48074_not n48303_not ; n48304
g48049 and n47582_not n48073_not ; n48305
g48050 and n48072_not n48305 ; n48306
g48051 and n48304_not n48306_not ; n48307
g48052 and b[27]_not n48307_not ; n48308
g48053 and n47601_not n47927 ; n48309
g48054 and n47923_not n48309 ; n48310
g48055 and n47924_not n47927_not ; n48311
g48056 and n48310_not n48311_not ; n48312
g48057 and n48074_not n48312_not ; n48313
g48058 and n47591_not n48073_not ; n48314
g48059 and n48072_not n48314 ; n48315
g48060 and n48313_not n48315_not ; n48316
g48061 and b[26]_not n48316_not ; n48317
g48062 and n47610_not n47922 ; n48318
g48063 and n47918_not n48318 ; n48319
g48064 and n47919_not n47922_not ; n48320
g48065 and n48319_not n48320_not ; n48321
g48066 and n48074_not n48321_not ; n48322
g48067 and n47600_not n48073_not ; n48323
g48068 and n48072_not n48323 ; n48324
g48069 and n48322_not n48324_not ; n48325
g48070 and b[25]_not n48325_not ; n48326
g48071 and n47619_not n47917 ; n48327
g48072 and n47913_not n48327 ; n48328
g48073 and n47914_not n47917_not ; n48329
g48074 and n48328_not n48329_not ; n48330
g48075 and n48074_not n48330_not ; n48331
g48076 and n47609_not n48073_not ; n48332
g48077 and n48072_not n48332 ; n48333
g48078 and n48331_not n48333_not ; n48334
g48079 and b[24]_not n48334_not ; n48335
g48080 and n47628_not n47912 ; n48336
g48081 and n47908_not n48336 ; n48337
g48082 and n47909_not n47912_not ; n48338
g48083 and n48337_not n48338_not ; n48339
g48084 and n48074_not n48339_not ; n48340
g48085 and n47618_not n48073_not ; n48341
g48086 and n48072_not n48341 ; n48342
g48087 and n48340_not n48342_not ; n48343
g48088 and b[23]_not n48343_not ; n48344
g48089 and n47637_not n47907 ; n48345
g48090 and n47903_not n48345 ; n48346
g48091 and n47904_not n47907_not ; n48347
g48092 and n48346_not n48347_not ; n48348
g48093 and n48074_not n48348_not ; n48349
g48094 and n47627_not n48073_not ; n48350
g48095 and n48072_not n48350 ; n48351
g48096 and n48349_not n48351_not ; n48352
g48097 and b[22]_not n48352_not ; n48353
g48098 and n47646_not n47902 ; n48354
g48099 and n47898_not n48354 ; n48355
g48100 and n47899_not n47902_not ; n48356
g48101 and n48355_not n48356_not ; n48357
g48102 and n48074_not n48357_not ; n48358
g48103 and n47636_not n48073_not ; n48359
g48104 and n48072_not n48359 ; n48360
g48105 and n48358_not n48360_not ; n48361
g48106 and b[21]_not n48361_not ; n48362
g48107 and n47655_not n47897 ; n48363
g48108 and n47893_not n48363 ; n48364
g48109 and n47894_not n47897_not ; n48365
g48110 and n48364_not n48365_not ; n48366
g48111 and n48074_not n48366_not ; n48367
g48112 and n47645_not n48073_not ; n48368
g48113 and n48072_not n48368 ; n48369
g48114 and n48367_not n48369_not ; n48370
g48115 and b[20]_not n48370_not ; n48371
g48116 and n47664_not n47892 ; n48372
g48117 and n47888_not n48372 ; n48373
g48118 and n47889_not n47892_not ; n48374
g48119 and n48373_not n48374_not ; n48375
g48120 and n48074_not n48375_not ; n48376
g48121 and n47654_not n48073_not ; n48377
g48122 and n48072_not n48377 ; n48378
g48123 and n48376_not n48378_not ; n48379
g48124 and b[19]_not n48379_not ; n48380
g48125 and n47673_not n47887 ; n48381
g48126 and n47883_not n48381 ; n48382
g48127 and n47884_not n47887_not ; n48383
g48128 and n48382_not n48383_not ; n48384
g48129 and n48074_not n48384_not ; n48385
g48130 and n47663_not n48073_not ; n48386
g48131 and n48072_not n48386 ; n48387
g48132 and n48385_not n48387_not ; n48388
g48133 and b[18]_not n48388_not ; n48389
g48134 and n47682_not n47882 ; n48390
g48135 and n47878_not n48390 ; n48391
g48136 and n47879_not n47882_not ; n48392
g48137 and n48391_not n48392_not ; n48393
g48138 and n48074_not n48393_not ; n48394
g48139 and n47672_not n48073_not ; n48395
g48140 and n48072_not n48395 ; n48396
g48141 and n48394_not n48396_not ; n48397
g48142 and b[17]_not n48397_not ; n48398
g48143 and n47691_not n47877 ; n48399
g48144 and n47873_not n48399 ; n48400
g48145 and n47874_not n47877_not ; n48401
g48146 and n48400_not n48401_not ; n48402
g48147 and n48074_not n48402_not ; n48403
g48148 and n47681_not n48073_not ; n48404
g48149 and n48072_not n48404 ; n48405
g48150 and n48403_not n48405_not ; n48406
g48151 and b[16]_not n48406_not ; n48407
g48152 and n47700_not n47872 ; n48408
g48153 and n47868_not n48408 ; n48409
g48154 and n47869_not n47872_not ; n48410
g48155 and n48409_not n48410_not ; n48411
g48156 and n48074_not n48411_not ; n48412
g48157 and n47690_not n48073_not ; n48413
g48158 and n48072_not n48413 ; n48414
g48159 and n48412_not n48414_not ; n48415
g48160 and b[15]_not n48415_not ; n48416
g48161 and n47709_not n47867 ; n48417
g48162 and n47863_not n48417 ; n48418
g48163 and n47864_not n47867_not ; n48419
g48164 and n48418_not n48419_not ; n48420
g48165 and n48074_not n48420_not ; n48421
g48166 and n47699_not n48073_not ; n48422
g48167 and n48072_not n48422 ; n48423
g48168 and n48421_not n48423_not ; n48424
g48169 and b[14]_not n48424_not ; n48425
g48170 and n47718_not n47862 ; n48426
g48171 and n47858_not n48426 ; n48427
g48172 and n47859_not n47862_not ; n48428
g48173 and n48427_not n48428_not ; n48429
g48174 and n48074_not n48429_not ; n48430
g48175 and n47708_not n48073_not ; n48431
g48176 and n48072_not n48431 ; n48432
g48177 and n48430_not n48432_not ; n48433
g48178 and b[13]_not n48433_not ; n48434
g48179 and n47727_not n47857 ; n48435
g48180 and n47853_not n48435 ; n48436
g48181 and n47854_not n47857_not ; n48437
g48182 and n48436_not n48437_not ; n48438
g48183 and n48074_not n48438_not ; n48439
g48184 and n47717_not n48073_not ; n48440
g48185 and n48072_not n48440 ; n48441
g48186 and n48439_not n48441_not ; n48442
g48187 and b[12]_not n48442_not ; n48443
g48188 and n47736_not n47852 ; n48444
g48189 and n47848_not n48444 ; n48445
g48190 and n47849_not n47852_not ; n48446
g48191 and n48445_not n48446_not ; n48447
g48192 and n48074_not n48447_not ; n48448
g48193 and n47726_not n48073_not ; n48449
g48194 and n48072_not n48449 ; n48450
g48195 and n48448_not n48450_not ; n48451
g48196 and b[11]_not n48451_not ; n48452
g48197 and n47745_not n47847 ; n48453
g48198 and n47843_not n48453 ; n48454
g48199 and n47844_not n47847_not ; n48455
g48200 and n48454_not n48455_not ; n48456
g48201 and n48074_not n48456_not ; n48457
g48202 and n47735_not n48073_not ; n48458
g48203 and n48072_not n48458 ; n48459
g48204 and n48457_not n48459_not ; n48460
g48205 and b[10]_not n48460_not ; n48461
g48206 and n47754_not n47842 ; n48462
g48207 and n47838_not n48462 ; n48463
g48208 and n47839_not n47842_not ; n48464
g48209 and n48463_not n48464_not ; n48465
g48210 and n48074_not n48465_not ; n48466
g48211 and n47744_not n48073_not ; n48467
g48212 and n48072_not n48467 ; n48468
g48213 and n48466_not n48468_not ; n48469
g48214 and b[9]_not n48469_not ; n48470
g48215 and n47763_not n47837 ; n48471
g48216 and n47833_not n48471 ; n48472
g48217 and n47834_not n47837_not ; n48473
g48218 and n48472_not n48473_not ; n48474
g48219 and n48074_not n48474_not ; n48475
g48220 and n47753_not n48073_not ; n48476
g48221 and n48072_not n48476 ; n48477
g48222 and n48475_not n48477_not ; n48478
g48223 and b[8]_not n48478_not ; n48479
g48224 and n47772_not n47832 ; n48480
g48225 and n47828_not n48480 ; n48481
g48226 and n47829_not n47832_not ; n48482
g48227 and n48481_not n48482_not ; n48483
g48228 and n48074_not n48483_not ; n48484
g48229 and n47762_not n48073_not ; n48485
g48230 and n48072_not n48485 ; n48486
g48231 and n48484_not n48486_not ; n48487
g48232 and b[7]_not n48487_not ; n48488
g48233 and n47781_not n47827 ; n48489
g48234 and n47823_not n48489 ; n48490
g48235 and n47824_not n47827_not ; n48491
g48236 and n48490_not n48491_not ; n48492
g48237 and n48074_not n48492_not ; n48493
g48238 and n47771_not n48073_not ; n48494
g48239 and n48072_not n48494 ; n48495
g48240 and n48493_not n48495_not ; n48496
g48241 and b[6]_not n48496_not ; n48497
g48242 and n47790_not n47822 ; n48498
g48243 and n47818_not n48498 ; n48499
g48244 and n47819_not n47822_not ; n48500
g48245 and n48499_not n48500_not ; n48501
g48246 and n48074_not n48501_not ; n48502
g48247 and n47780_not n48073_not ; n48503
g48248 and n48072_not n48503 ; n48504
g48249 and n48502_not n48504_not ; n48505
g48250 and b[5]_not n48505_not ; n48506
g48251 and n47798_not n47817 ; n48507
g48252 and n47813_not n48507 ; n48508
g48253 and n47814_not n47817_not ; n48509
g48254 and n48508_not n48509_not ; n48510
g48255 and n48074_not n48510_not ; n48511
g48256 and n47789_not n48073_not ; n48512
g48257 and n48072_not n48512 ; n48513
g48258 and n48511_not n48513_not ; n48514
g48259 and b[4]_not n48514_not ; n48515
g48260 and n47808_not n47812 ; n48516
g48261 and n47807_not n48516 ; n48517
g48262 and n47809_not n47812_not ; n48518
g48263 and n48517_not n48518_not ; n48519
g48264 and n48074_not n48519_not ; n48520
g48265 and n47797_not n48073_not ; n48521
g48266 and n48072_not n48521 ; n48522
g48267 and n48520_not n48522_not ; n48523
g48268 and b[3]_not n48523_not ; n48524
g48269 and n19767 n47805_not ; n48525
g48270 and n47803_not n48525 ; n48526
g48271 and n47807_not n48526_not ; n48527
g48272 and n48074_not n48527 ; n48528
g48273 and n47802_not n48073_not ; n48529
g48274 and n48072_not n48529 ; n48530
g48275 and n48528_not n48530_not ; n48531
g48276 and b[2]_not n48531_not ; n48532
g48277 and b[0] n48074_not ; n48533
g48278 and a[11] n48533_not ; n48534
g48279 and n19767 n48074_not ; n48535
g48280 and n48534_not n48535_not ; n48536
g48281 and b[1] n48536_not ; n48537
g48282 and b[1]_not n48535_not ; n48538
g48283 and n48534_not n48538 ; n48539
g48284 and n48537_not n48539_not ; n48540
g48285 and n20502_not n48540_not ; n48541
g48286 and b[1]_not n48536_not ; n48542
g48287 and n48541_not n48542_not ; n48543
g48288 and b[2] n48530_not ; n48544
g48289 and n48528_not n48544 ; n48545
g48290 and n48532_not n48545_not ; n48546
g48291 and n48543_not n48546 ; n48547
g48292 and n48532_not n48547_not ; n48548
g48293 and b[3] n48522_not ; n48549
g48294 and n48520_not n48549 ; n48550
g48295 and n48524_not n48550_not ; n48551
g48296 and n48548_not n48551 ; n48552
g48297 and n48524_not n48552_not ; n48553
g48298 and b[4] n48513_not ; n48554
g48299 and n48511_not n48554 ; n48555
g48300 and n48515_not n48555_not ; n48556
g48301 and n48553_not n48556 ; n48557
g48302 and n48515_not n48557_not ; n48558
g48303 and b[5] n48504_not ; n48559
g48304 and n48502_not n48559 ; n48560
g48305 and n48506_not n48560_not ; n48561
g48306 and n48558_not n48561 ; n48562
g48307 and n48506_not n48562_not ; n48563
g48308 and b[6] n48495_not ; n48564
g48309 and n48493_not n48564 ; n48565
g48310 and n48497_not n48565_not ; n48566
g48311 and n48563_not n48566 ; n48567
g48312 and n48497_not n48567_not ; n48568
g48313 and b[7] n48486_not ; n48569
g48314 and n48484_not n48569 ; n48570
g48315 and n48488_not n48570_not ; n48571
g48316 and n48568_not n48571 ; n48572
g48317 and n48488_not n48572_not ; n48573
g48318 and b[8] n48477_not ; n48574
g48319 and n48475_not n48574 ; n48575
g48320 and n48479_not n48575_not ; n48576
g48321 and n48573_not n48576 ; n48577
g48322 and n48479_not n48577_not ; n48578
g48323 and b[9] n48468_not ; n48579
g48324 and n48466_not n48579 ; n48580
g48325 and n48470_not n48580_not ; n48581
g48326 and n48578_not n48581 ; n48582
g48327 and n48470_not n48582_not ; n48583
g48328 and b[10] n48459_not ; n48584
g48329 and n48457_not n48584 ; n48585
g48330 and n48461_not n48585_not ; n48586
g48331 and n48583_not n48586 ; n48587
g48332 and n48461_not n48587_not ; n48588
g48333 and b[11] n48450_not ; n48589
g48334 and n48448_not n48589 ; n48590
g48335 and n48452_not n48590_not ; n48591
g48336 and n48588_not n48591 ; n48592
g48337 and n48452_not n48592_not ; n48593
g48338 and b[12] n48441_not ; n48594
g48339 and n48439_not n48594 ; n48595
g48340 and n48443_not n48595_not ; n48596
g48341 and n48593_not n48596 ; n48597
g48342 and n48443_not n48597_not ; n48598
g48343 and b[13] n48432_not ; n48599
g48344 and n48430_not n48599 ; n48600
g48345 and n48434_not n48600_not ; n48601
g48346 and n48598_not n48601 ; n48602
g48347 and n48434_not n48602_not ; n48603
g48348 and b[14] n48423_not ; n48604
g48349 and n48421_not n48604 ; n48605
g48350 and n48425_not n48605_not ; n48606
g48351 and n48603_not n48606 ; n48607
g48352 and n48425_not n48607_not ; n48608
g48353 and b[15] n48414_not ; n48609
g48354 and n48412_not n48609 ; n48610
g48355 and n48416_not n48610_not ; n48611
g48356 and n48608_not n48611 ; n48612
g48357 and n48416_not n48612_not ; n48613
g48358 and b[16] n48405_not ; n48614
g48359 and n48403_not n48614 ; n48615
g48360 and n48407_not n48615_not ; n48616
g48361 and n48613_not n48616 ; n48617
g48362 and n48407_not n48617_not ; n48618
g48363 and b[17] n48396_not ; n48619
g48364 and n48394_not n48619 ; n48620
g48365 and n48398_not n48620_not ; n48621
g48366 and n48618_not n48621 ; n48622
g48367 and n48398_not n48622_not ; n48623
g48368 and b[18] n48387_not ; n48624
g48369 and n48385_not n48624 ; n48625
g48370 and n48389_not n48625_not ; n48626
g48371 and n48623_not n48626 ; n48627
g48372 and n48389_not n48627_not ; n48628
g48373 and b[19] n48378_not ; n48629
g48374 and n48376_not n48629 ; n48630
g48375 and n48380_not n48630_not ; n48631
g48376 and n48628_not n48631 ; n48632
g48377 and n48380_not n48632_not ; n48633
g48378 and b[20] n48369_not ; n48634
g48379 and n48367_not n48634 ; n48635
g48380 and n48371_not n48635_not ; n48636
g48381 and n48633_not n48636 ; n48637
g48382 and n48371_not n48637_not ; n48638
g48383 and b[21] n48360_not ; n48639
g48384 and n48358_not n48639 ; n48640
g48385 and n48362_not n48640_not ; n48641
g48386 and n48638_not n48641 ; n48642
g48387 and n48362_not n48642_not ; n48643
g48388 and b[22] n48351_not ; n48644
g48389 and n48349_not n48644 ; n48645
g48390 and n48353_not n48645_not ; n48646
g48391 and n48643_not n48646 ; n48647
g48392 and n48353_not n48647_not ; n48648
g48393 and b[23] n48342_not ; n48649
g48394 and n48340_not n48649 ; n48650
g48395 and n48344_not n48650_not ; n48651
g48396 and n48648_not n48651 ; n48652
g48397 and n48344_not n48652_not ; n48653
g48398 and b[24] n48333_not ; n48654
g48399 and n48331_not n48654 ; n48655
g48400 and n48335_not n48655_not ; n48656
g48401 and n48653_not n48656 ; n48657
g48402 and n48335_not n48657_not ; n48658
g48403 and b[25] n48324_not ; n48659
g48404 and n48322_not n48659 ; n48660
g48405 and n48326_not n48660_not ; n48661
g48406 and n48658_not n48661 ; n48662
g48407 and n48326_not n48662_not ; n48663
g48408 and b[26] n48315_not ; n48664
g48409 and n48313_not n48664 ; n48665
g48410 and n48317_not n48665_not ; n48666
g48411 and n48663_not n48666 ; n48667
g48412 and n48317_not n48667_not ; n48668
g48413 and b[27] n48306_not ; n48669
g48414 and n48304_not n48669 ; n48670
g48415 and n48308_not n48670_not ; n48671
g48416 and n48668_not n48671 ; n48672
g48417 and n48308_not n48672_not ; n48673
g48418 and b[28] n48297_not ; n48674
g48419 and n48295_not n48674 ; n48675
g48420 and n48299_not n48675_not ; n48676
g48421 and n48673_not n48676 ; n48677
g48422 and n48299_not n48677_not ; n48678
g48423 and b[29] n48288_not ; n48679
g48424 and n48286_not n48679 ; n48680
g48425 and n48290_not n48680_not ; n48681
g48426 and n48678_not n48681 ; n48682
g48427 and n48290_not n48682_not ; n48683
g48428 and b[30] n48279_not ; n48684
g48429 and n48277_not n48684 ; n48685
g48430 and n48281_not n48685_not ; n48686
g48431 and n48683_not n48686 ; n48687
g48432 and n48281_not n48687_not ; n48688
g48433 and b[31] n48270_not ; n48689
g48434 and n48268_not n48689 ; n48690
g48435 and n48272_not n48690_not ; n48691
g48436 and n48688_not n48691 ; n48692
g48437 and n48272_not n48692_not ; n48693
g48438 and b[32] n48261_not ; n48694
g48439 and n48259_not n48694 ; n48695
g48440 and n48263_not n48695_not ; n48696
g48441 and n48693_not n48696 ; n48697
g48442 and n48263_not n48697_not ; n48698
g48443 and b[33] n48252_not ; n48699
g48444 and n48250_not n48699 ; n48700
g48445 and n48254_not n48700_not ; n48701
g48446 and n48698_not n48701 ; n48702
g48447 and n48254_not n48702_not ; n48703
g48448 and b[34] n48243_not ; n48704
g48449 and n48241_not n48704 ; n48705
g48450 and n48245_not n48705_not ; n48706
g48451 and n48703_not n48706 ; n48707
g48452 and n48245_not n48707_not ; n48708
g48453 and b[35] n48234_not ; n48709
g48454 and n48232_not n48709 ; n48710
g48455 and n48236_not n48710_not ; n48711
g48456 and n48708_not n48711 ; n48712
g48457 and n48236_not n48712_not ; n48713
g48458 and b[36] n48225_not ; n48714
g48459 and n48223_not n48714 ; n48715
g48460 and n48227_not n48715_not ; n48716
g48461 and n48713_not n48716 ; n48717
g48462 and n48227_not n48717_not ; n48718
g48463 and b[37] n48216_not ; n48719
g48464 and n48214_not n48719 ; n48720
g48465 and n48218_not n48720_not ; n48721
g48466 and n48718_not n48721 ; n48722
g48467 and n48218_not n48722_not ; n48723
g48468 and b[38] n48207_not ; n48724
g48469 and n48205_not n48724 ; n48725
g48470 and n48209_not n48725_not ; n48726
g48471 and n48723_not n48726 ; n48727
g48472 and n48209_not n48727_not ; n48728
g48473 and b[39] n48198_not ; n48729
g48474 and n48196_not n48729 ; n48730
g48475 and n48200_not n48730_not ; n48731
g48476 and n48728_not n48731 ; n48732
g48477 and n48200_not n48732_not ; n48733
g48478 and b[40] n48189_not ; n48734
g48479 and n48187_not n48734 ; n48735
g48480 and n48191_not n48735_not ; n48736
g48481 and n48733_not n48736 ; n48737
g48482 and n48191_not n48737_not ; n48738
g48483 and b[41] n48180_not ; n48739
g48484 and n48178_not n48739 ; n48740
g48485 and n48182_not n48740_not ; n48741
g48486 and n48738_not n48741 ; n48742
g48487 and n48182_not n48742_not ; n48743
g48488 and b[42] n48171_not ; n48744
g48489 and n48169_not n48744 ; n48745
g48490 and n48173_not n48745_not ; n48746
g48491 and n48743_not n48746 ; n48747
g48492 and n48173_not n48747_not ; n48748
g48493 and b[43] n48162_not ; n48749
g48494 and n48160_not n48749 ; n48750
g48495 and n48164_not n48750_not ; n48751
g48496 and n48748_not n48751 ; n48752
g48497 and n48164_not n48752_not ; n48753
g48498 and b[44] n48153_not ; n48754
g48499 and n48151_not n48754 ; n48755
g48500 and n48155_not n48755_not ; n48756
g48501 and n48753_not n48756 ; n48757
g48502 and n48155_not n48757_not ; n48758
g48503 and b[45] n48144_not ; n48759
g48504 and n48142_not n48759 ; n48760
g48505 and n48146_not n48760_not ; n48761
g48506 and n48758_not n48761 ; n48762
g48507 and n48146_not n48762_not ; n48763
g48508 and b[46] n48135_not ; n48764
g48509 and n48133_not n48764 ; n48765
g48510 and n48137_not n48765_not ; n48766
g48511 and n48763_not n48766 ; n48767
g48512 and n48137_not n48767_not ; n48768
g48513 and b[47] n48126_not ; n48769
g48514 and n48124_not n48769 ; n48770
g48515 and n48128_not n48770_not ; n48771
g48516 and n48768_not n48771 ; n48772
g48517 and n48128_not n48772_not ; n48773
g48518 and b[48] n48117_not ; n48774
g48519 and n48115_not n48774 ; n48775
g48520 and n48119_not n48775_not ; n48776
g48521 and n48773_not n48776 ; n48777
g48522 and n48119_not n48777_not ; n48778
g48523 and b[49] n48108_not ; n48779
g48524 and n48106_not n48779 ; n48780
g48525 and n48110_not n48780_not ; n48781
g48526 and n48778_not n48781 ; n48782
g48527 and n48110_not n48782_not ; n48783
g48528 and b[50] n48099_not ; n48784
g48529 and n48097_not n48784 ; n48785
g48530 and n48101_not n48785_not ; n48786
g48531 and n48783_not n48786 ; n48787
g48532 and n48101_not n48787_not ; n48788
g48533 and b[51] n48090_not ; n48789
g48534 and n48088_not n48789 ; n48790
g48535 and n48092_not n48790_not ; n48791
g48536 and n48788_not n48791 ; n48792
g48537 and n48092_not n48792_not ; n48793
g48538 and b[52] n48081_not ; n48794
g48539 and n48079_not n48794 ; n48795
g48540 and n48083_not n48795_not ; n48796
g48541 and n48793_not n48796 ; n48797
g48542 and n48083_not n48797_not ; n48798
g48543 and n47358_not n48069_not ; n48799
g48544 and n48067_not n48799 ; n48800
g48545 and n48058_not n48800 ; n48801
g48546 and n48067_not n48069_not ; n48802
g48547 and n48059_not n48802_not ; n48803
g48548 and n48801_not n48803_not ; n48804
g48549 and n48074_not n48804_not ; n48805
g48550 and n48066_not n48073_not ; n48806
g48551 and n48072_not n48806 ; n48807
g48552 and n48805_not n48807_not ; n48808
g48553 and b[53]_not n48808_not ; n48809
g48554 and b[53] n48807_not ; n48810
g48555 and n48805_not n48810 ; n48811
g48556 and n20775 n48811_not ; n48812
g48557 and n48809_not n48812 ; n48813
g48558 and n48798_not n48813 ; n48814
g48559 and n595 n48808_not ; n48815
g48560 and n48814_not n48815_not ; n48816
g48561 and n48092_not n48796 ; n48817
g48562 and n48792_not n48817 ; n48818
g48563 and n48793_not n48796_not ; n48819
g48564 and n48818_not n48819_not ; n48820
g48565 and n48816_not n48820_not ; n48821
g48566 and n48082_not n48815_not ; n48822
g48567 and n48814_not n48822 ; n48823
g48568 and n48821_not n48823_not ; n48824
g48569 and n48083_not n48811_not ; n48825
g48570 and n48809_not n48825 ; n48826
g48571 and n48797_not n48826 ; n48827
g48572 and n48809_not n48811_not ; n48828
g48573 and n48798_not n48828_not ; n48829
g48574 and n48827_not n48829_not ; n48830
g48575 and n48816_not n48830_not ; n48831
g48576 and n48808_not n48815_not ; n48832
g48577 and n48814_not n48832 ; n48833
g48578 and n48831_not n48833_not ; n48834
g48579 and b[54]_not n48834_not ; n48835
g48580 and b[53]_not n48824_not ; n48836
g48581 and n48101_not n48791 ; n48837
g48582 and n48787_not n48837 ; n48838
g48583 and n48788_not n48791_not ; n48839
g48584 and n48838_not n48839_not ; n48840
g48585 and n48816_not n48840_not ; n48841
g48586 and n48091_not n48815_not ; n48842
g48587 and n48814_not n48842 ; n48843
g48588 and n48841_not n48843_not ; n48844
g48589 and b[52]_not n48844_not ; n48845
g48590 and n48110_not n48786 ; n48846
g48591 and n48782_not n48846 ; n48847
g48592 and n48783_not n48786_not ; n48848
g48593 and n48847_not n48848_not ; n48849
g48594 and n48816_not n48849_not ; n48850
g48595 and n48100_not n48815_not ; n48851
g48596 and n48814_not n48851 ; n48852
g48597 and n48850_not n48852_not ; n48853
g48598 and b[51]_not n48853_not ; n48854
g48599 and n48119_not n48781 ; n48855
g48600 and n48777_not n48855 ; n48856
g48601 and n48778_not n48781_not ; n48857
g48602 and n48856_not n48857_not ; n48858
g48603 and n48816_not n48858_not ; n48859
g48604 and n48109_not n48815_not ; n48860
g48605 and n48814_not n48860 ; n48861
g48606 and n48859_not n48861_not ; n48862
g48607 and b[50]_not n48862_not ; n48863
g48608 and n48128_not n48776 ; n48864
g48609 and n48772_not n48864 ; n48865
g48610 and n48773_not n48776_not ; n48866
g48611 and n48865_not n48866_not ; n48867
g48612 and n48816_not n48867_not ; n48868
g48613 and n48118_not n48815_not ; n48869
g48614 and n48814_not n48869 ; n48870
g48615 and n48868_not n48870_not ; n48871
g48616 and b[49]_not n48871_not ; n48872
g48617 and n48137_not n48771 ; n48873
g48618 and n48767_not n48873 ; n48874
g48619 and n48768_not n48771_not ; n48875
g48620 and n48874_not n48875_not ; n48876
g48621 and n48816_not n48876_not ; n48877
g48622 and n48127_not n48815_not ; n48878
g48623 and n48814_not n48878 ; n48879
g48624 and n48877_not n48879_not ; n48880
g48625 and b[48]_not n48880_not ; n48881
g48626 and n48146_not n48766 ; n48882
g48627 and n48762_not n48882 ; n48883
g48628 and n48763_not n48766_not ; n48884
g48629 and n48883_not n48884_not ; n48885
g48630 and n48816_not n48885_not ; n48886
g48631 and n48136_not n48815_not ; n48887
g48632 and n48814_not n48887 ; n48888
g48633 and n48886_not n48888_not ; n48889
g48634 and b[47]_not n48889_not ; n48890
g48635 and n48155_not n48761 ; n48891
g48636 and n48757_not n48891 ; n48892
g48637 and n48758_not n48761_not ; n48893
g48638 and n48892_not n48893_not ; n48894
g48639 and n48816_not n48894_not ; n48895
g48640 and n48145_not n48815_not ; n48896
g48641 and n48814_not n48896 ; n48897
g48642 and n48895_not n48897_not ; n48898
g48643 and b[46]_not n48898_not ; n48899
g48644 and n48164_not n48756 ; n48900
g48645 and n48752_not n48900 ; n48901
g48646 and n48753_not n48756_not ; n48902
g48647 and n48901_not n48902_not ; n48903
g48648 and n48816_not n48903_not ; n48904
g48649 and n48154_not n48815_not ; n48905
g48650 and n48814_not n48905 ; n48906
g48651 and n48904_not n48906_not ; n48907
g48652 and b[45]_not n48907_not ; n48908
g48653 and n48173_not n48751 ; n48909
g48654 and n48747_not n48909 ; n48910
g48655 and n48748_not n48751_not ; n48911
g48656 and n48910_not n48911_not ; n48912
g48657 and n48816_not n48912_not ; n48913
g48658 and n48163_not n48815_not ; n48914
g48659 and n48814_not n48914 ; n48915
g48660 and n48913_not n48915_not ; n48916
g48661 and b[44]_not n48916_not ; n48917
g48662 and n48182_not n48746 ; n48918
g48663 and n48742_not n48918 ; n48919
g48664 and n48743_not n48746_not ; n48920
g48665 and n48919_not n48920_not ; n48921
g48666 and n48816_not n48921_not ; n48922
g48667 and n48172_not n48815_not ; n48923
g48668 and n48814_not n48923 ; n48924
g48669 and n48922_not n48924_not ; n48925
g48670 and b[43]_not n48925_not ; n48926
g48671 and n48191_not n48741 ; n48927
g48672 and n48737_not n48927 ; n48928
g48673 and n48738_not n48741_not ; n48929
g48674 and n48928_not n48929_not ; n48930
g48675 and n48816_not n48930_not ; n48931
g48676 and n48181_not n48815_not ; n48932
g48677 and n48814_not n48932 ; n48933
g48678 and n48931_not n48933_not ; n48934
g48679 and b[42]_not n48934_not ; n48935
g48680 and n48200_not n48736 ; n48936
g48681 and n48732_not n48936 ; n48937
g48682 and n48733_not n48736_not ; n48938
g48683 and n48937_not n48938_not ; n48939
g48684 and n48816_not n48939_not ; n48940
g48685 and n48190_not n48815_not ; n48941
g48686 and n48814_not n48941 ; n48942
g48687 and n48940_not n48942_not ; n48943
g48688 and b[41]_not n48943_not ; n48944
g48689 and n48209_not n48731 ; n48945
g48690 and n48727_not n48945 ; n48946
g48691 and n48728_not n48731_not ; n48947
g48692 and n48946_not n48947_not ; n48948
g48693 and n48816_not n48948_not ; n48949
g48694 and n48199_not n48815_not ; n48950
g48695 and n48814_not n48950 ; n48951
g48696 and n48949_not n48951_not ; n48952
g48697 and b[40]_not n48952_not ; n48953
g48698 and n48218_not n48726 ; n48954
g48699 and n48722_not n48954 ; n48955
g48700 and n48723_not n48726_not ; n48956
g48701 and n48955_not n48956_not ; n48957
g48702 and n48816_not n48957_not ; n48958
g48703 and n48208_not n48815_not ; n48959
g48704 and n48814_not n48959 ; n48960
g48705 and n48958_not n48960_not ; n48961
g48706 and b[39]_not n48961_not ; n48962
g48707 and n48227_not n48721 ; n48963
g48708 and n48717_not n48963 ; n48964
g48709 and n48718_not n48721_not ; n48965
g48710 and n48964_not n48965_not ; n48966
g48711 and n48816_not n48966_not ; n48967
g48712 and n48217_not n48815_not ; n48968
g48713 and n48814_not n48968 ; n48969
g48714 and n48967_not n48969_not ; n48970
g48715 and b[38]_not n48970_not ; n48971
g48716 and n48236_not n48716 ; n48972
g48717 and n48712_not n48972 ; n48973
g48718 and n48713_not n48716_not ; n48974
g48719 and n48973_not n48974_not ; n48975
g48720 and n48816_not n48975_not ; n48976
g48721 and n48226_not n48815_not ; n48977
g48722 and n48814_not n48977 ; n48978
g48723 and n48976_not n48978_not ; n48979
g48724 and b[37]_not n48979_not ; n48980
g48725 and n48245_not n48711 ; n48981
g48726 and n48707_not n48981 ; n48982
g48727 and n48708_not n48711_not ; n48983
g48728 and n48982_not n48983_not ; n48984
g48729 and n48816_not n48984_not ; n48985
g48730 and n48235_not n48815_not ; n48986
g48731 and n48814_not n48986 ; n48987
g48732 and n48985_not n48987_not ; n48988
g48733 and b[36]_not n48988_not ; n48989
g48734 and n48254_not n48706 ; n48990
g48735 and n48702_not n48990 ; n48991
g48736 and n48703_not n48706_not ; n48992
g48737 and n48991_not n48992_not ; n48993
g48738 and n48816_not n48993_not ; n48994
g48739 and n48244_not n48815_not ; n48995
g48740 and n48814_not n48995 ; n48996
g48741 and n48994_not n48996_not ; n48997
g48742 and b[35]_not n48997_not ; n48998
g48743 and n48263_not n48701 ; n48999
g48744 and n48697_not n48999 ; n49000
g48745 and n48698_not n48701_not ; n49001
g48746 and n49000_not n49001_not ; n49002
g48747 and n48816_not n49002_not ; n49003
g48748 and n48253_not n48815_not ; n49004
g48749 and n48814_not n49004 ; n49005
g48750 and n49003_not n49005_not ; n49006
g48751 and b[34]_not n49006_not ; n49007
g48752 and n48272_not n48696 ; n49008
g48753 and n48692_not n49008 ; n49009
g48754 and n48693_not n48696_not ; n49010
g48755 and n49009_not n49010_not ; n49011
g48756 and n48816_not n49011_not ; n49012
g48757 and n48262_not n48815_not ; n49013
g48758 and n48814_not n49013 ; n49014
g48759 and n49012_not n49014_not ; n49015
g48760 and b[33]_not n49015_not ; n49016
g48761 and n48281_not n48691 ; n49017
g48762 and n48687_not n49017 ; n49018
g48763 and n48688_not n48691_not ; n49019
g48764 and n49018_not n49019_not ; n49020
g48765 and n48816_not n49020_not ; n49021
g48766 and n48271_not n48815_not ; n49022
g48767 and n48814_not n49022 ; n49023
g48768 and n49021_not n49023_not ; n49024
g48769 and b[32]_not n49024_not ; n49025
g48770 and n48290_not n48686 ; n49026
g48771 and n48682_not n49026 ; n49027
g48772 and n48683_not n48686_not ; n49028
g48773 and n49027_not n49028_not ; n49029
g48774 and n48816_not n49029_not ; n49030
g48775 and n48280_not n48815_not ; n49031
g48776 and n48814_not n49031 ; n49032
g48777 and n49030_not n49032_not ; n49033
g48778 and b[31]_not n49033_not ; n49034
g48779 and n48299_not n48681 ; n49035
g48780 and n48677_not n49035 ; n49036
g48781 and n48678_not n48681_not ; n49037
g48782 and n49036_not n49037_not ; n49038
g48783 and n48816_not n49038_not ; n49039
g48784 and n48289_not n48815_not ; n49040
g48785 and n48814_not n49040 ; n49041
g48786 and n49039_not n49041_not ; n49042
g48787 and b[30]_not n49042_not ; n49043
g48788 and n48308_not n48676 ; n49044
g48789 and n48672_not n49044 ; n49045
g48790 and n48673_not n48676_not ; n49046
g48791 and n49045_not n49046_not ; n49047
g48792 and n48816_not n49047_not ; n49048
g48793 and n48298_not n48815_not ; n49049
g48794 and n48814_not n49049 ; n49050
g48795 and n49048_not n49050_not ; n49051
g48796 and b[29]_not n49051_not ; n49052
g48797 and n48317_not n48671 ; n49053
g48798 and n48667_not n49053 ; n49054
g48799 and n48668_not n48671_not ; n49055
g48800 and n49054_not n49055_not ; n49056
g48801 and n48816_not n49056_not ; n49057
g48802 and n48307_not n48815_not ; n49058
g48803 and n48814_not n49058 ; n49059
g48804 and n49057_not n49059_not ; n49060
g48805 and b[28]_not n49060_not ; n49061
g48806 and n48326_not n48666 ; n49062
g48807 and n48662_not n49062 ; n49063
g48808 and n48663_not n48666_not ; n49064
g48809 and n49063_not n49064_not ; n49065
g48810 and n48816_not n49065_not ; n49066
g48811 and n48316_not n48815_not ; n49067
g48812 and n48814_not n49067 ; n49068
g48813 and n49066_not n49068_not ; n49069
g48814 and b[27]_not n49069_not ; n49070
g48815 and n48335_not n48661 ; n49071
g48816 and n48657_not n49071 ; n49072
g48817 and n48658_not n48661_not ; n49073
g48818 and n49072_not n49073_not ; n49074
g48819 and n48816_not n49074_not ; n49075
g48820 and n48325_not n48815_not ; n49076
g48821 and n48814_not n49076 ; n49077
g48822 and n49075_not n49077_not ; n49078
g48823 and b[26]_not n49078_not ; n49079
g48824 and n48344_not n48656 ; n49080
g48825 and n48652_not n49080 ; n49081
g48826 and n48653_not n48656_not ; n49082
g48827 and n49081_not n49082_not ; n49083
g48828 and n48816_not n49083_not ; n49084
g48829 and n48334_not n48815_not ; n49085
g48830 and n48814_not n49085 ; n49086
g48831 and n49084_not n49086_not ; n49087
g48832 and b[25]_not n49087_not ; n49088
g48833 and n48353_not n48651 ; n49089
g48834 and n48647_not n49089 ; n49090
g48835 and n48648_not n48651_not ; n49091
g48836 and n49090_not n49091_not ; n49092
g48837 and n48816_not n49092_not ; n49093
g48838 and n48343_not n48815_not ; n49094
g48839 and n48814_not n49094 ; n49095
g48840 and n49093_not n49095_not ; n49096
g48841 and b[24]_not n49096_not ; n49097
g48842 and n48362_not n48646 ; n49098
g48843 and n48642_not n49098 ; n49099
g48844 and n48643_not n48646_not ; n49100
g48845 and n49099_not n49100_not ; n49101
g48846 and n48816_not n49101_not ; n49102
g48847 and n48352_not n48815_not ; n49103
g48848 and n48814_not n49103 ; n49104
g48849 and n49102_not n49104_not ; n49105
g48850 and b[23]_not n49105_not ; n49106
g48851 and n48371_not n48641 ; n49107
g48852 and n48637_not n49107 ; n49108
g48853 and n48638_not n48641_not ; n49109
g48854 and n49108_not n49109_not ; n49110
g48855 and n48816_not n49110_not ; n49111
g48856 and n48361_not n48815_not ; n49112
g48857 and n48814_not n49112 ; n49113
g48858 and n49111_not n49113_not ; n49114
g48859 and b[22]_not n49114_not ; n49115
g48860 and n48380_not n48636 ; n49116
g48861 and n48632_not n49116 ; n49117
g48862 and n48633_not n48636_not ; n49118
g48863 and n49117_not n49118_not ; n49119
g48864 and n48816_not n49119_not ; n49120
g48865 and n48370_not n48815_not ; n49121
g48866 and n48814_not n49121 ; n49122
g48867 and n49120_not n49122_not ; n49123
g48868 and b[21]_not n49123_not ; n49124
g48869 and n48389_not n48631 ; n49125
g48870 and n48627_not n49125 ; n49126
g48871 and n48628_not n48631_not ; n49127
g48872 and n49126_not n49127_not ; n49128
g48873 and n48816_not n49128_not ; n49129
g48874 and n48379_not n48815_not ; n49130
g48875 and n48814_not n49130 ; n49131
g48876 and n49129_not n49131_not ; n49132
g48877 and b[20]_not n49132_not ; n49133
g48878 and n48398_not n48626 ; n49134
g48879 and n48622_not n49134 ; n49135
g48880 and n48623_not n48626_not ; n49136
g48881 and n49135_not n49136_not ; n49137
g48882 and n48816_not n49137_not ; n49138
g48883 and n48388_not n48815_not ; n49139
g48884 and n48814_not n49139 ; n49140
g48885 and n49138_not n49140_not ; n49141
g48886 and b[19]_not n49141_not ; n49142
g48887 and n48407_not n48621 ; n49143
g48888 and n48617_not n49143 ; n49144
g48889 and n48618_not n48621_not ; n49145
g48890 and n49144_not n49145_not ; n49146
g48891 and n48816_not n49146_not ; n49147
g48892 and n48397_not n48815_not ; n49148
g48893 and n48814_not n49148 ; n49149
g48894 and n49147_not n49149_not ; n49150
g48895 and b[18]_not n49150_not ; n49151
g48896 and n48416_not n48616 ; n49152
g48897 and n48612_not n49152 ; n49153
g48898 and n48613_not n48616_not ; n49154
g48899 and n49153_not n49154_not ; n49155
g48900 and n48816_not n49155_not ; n49156
g48901 and n48406_not n48815_not ; n49157
g48902 and n48814_not n49157 ; n49158
g48903 and n49156_not n49158_not ; n49159
g48904 and b[17]_not n49159_not ; n49160
g48905 and n48425_not n48611 ; n49161
g48906 and n48607_not n49161 ; n49162
g48907 and n48608_not n48611_not ; n49163
g48908 and n49162_not n49163_not ; n49164
g48909 and n48816_not n49164_not ; n49165
g48910 and n48415_not n48815_not ; n49166
g48911 and n48814_not n49166 ; n49167
g48912 and n49165_not n49167_not ; n49168
g48913 and b[16]_not n49168_not ; n49169
g48914 and n48434_not n48606 ; n49170
g48915 and n48602_not n49170 ; n49171
g48916 and n48603_not n48606_not ; n49172
g48917 and n49171_not n49172_not ; n49173
g48918 and n48816_not n49173_not ; n49174
g48919 and n48424_not n48815_not ; n49175
g48920 and n48814_not n49175 ; n49176
g48921 and n49174_not n49176_not ; n49177
g48922 and b[15]_not n49177_not ; n49178
g48923 and n48443_not n48601 ; n49179
g48924 and n48597_not n49179 ; n49180
g48925 and n48598_not n48601_not ; n49181
g48926 and n49180_not n49181_not ; n49182
g48927 and n48816_not n49182_not ; n49183
g48928 and n48433_not n48815_not ; n49184
g48929 and n48814_not n49184 ; n49185
g48930 and n49183_not n49185_not ; n49186
g48931 and b[14]_not n49186_not ; n49187
g48932 and n48452_not n48596 ; n49188
g48933 and n48592_not n49188 ; n49189
g48934 and n48593_not n48596_not ; n49190
g48935 and n49189_not n49190_not ; n49191
g48936 and n48816_not n49191_not ; n49192
g48937 and n48442_not n48815_not ; n49193
g48938 and n48814_not n49193 ; n49194
g48939 and n49192_not n49194_not ; n49195
g48940 and b[13]_not n49195_not ; n49196
g48941 and n48461_not n48591 ; n49197
g48942 and n48587_not n49197 ; n49198
g48943 and n48588_not n48591_not ; n49199
g48944 and n49198_not n49199_not ; n49200
g48945 and n48816_not n49200_not ; n49201
g48946 and n48451_not n48815_not ; n49202
g48947 and n48814_not n49202 ; n49203
g48948 and n49201_not n49203_not ; n49204
g48949 and b[12]_not n49204_not ; n49205
g48950 and n48470_not n48586 ; n49206
g48951 and n48582_not n49206 ; n49207
g48952 and n48583_not n48586_not ; n49208
g48953 and n49207_not n49208_not ; n49209
g48954 and n48816_not n49209_not ; n49210
g48955 and n48460_not n48815_not ; n49211
g48956 and n48814_not n49211 ; n49212
g48957 and n49210_not n49212_not ; n49213
g48958 and b[11]_not n49213_not ; n49214
g48959 and n48479_not n48581 ; n49215
g48960 and n48577_not n49215 ; n49216
g48961 and n48578_not n48581_not ; n49217
g48962 and n49216_not n49217_not ; n49218
g48963 and n48816_not n49218_not ; n49219
g48964 and n48469_not n48815_not ; n49220
g48965 and n48814_not n49220 ; n49221
g48966 and n49219_not n49221_not ; n49222
g48967 and b[10]_not n49222_not ; n49223
g48968 and n48488_not n48576 ; n49224
g48969 and n48572_not n49224 ; n49225
g48970 and n48573_not n48576_not ; n49226
g48971 and n49225_not n49226_not ; n49227
g48972 and n48816_not n49227_not ; n49228
g48973 and n48478_not n48815_not ; n49229
g48974 and n48814_not n49229 ; n49230
g48975 and n49228_not n49230_not ; n49231
g48976 and b[9]_not n49231_not ; n49232
g48977 and n48497_not n48571 ; n49233
g48978 and n48567_not n49233 ; n49234
g48979 and n48568_not n48571_not ; n49235
g48980 and n49234_not n49235_not ; n49236
g48981 and n48816_not n49236_not ; n49237
g48982 and n48487_not n48815_not ; n49238
g48983 and n48814_not n49238 ; n49239
g48984 and n49237_not n49239_not ; n49240
g48985 and b[8]_not n49240_not ; n49241
g48986 and n48506_not n48566 ; n49242
g48987 and n48562_not n49242 ; n49243
g48988 and n48563_not n48566_not ; n49244
g48989 and n49243_not n49244_not ; n49245
g48990 and n48816_not n49245_not ; n49246
g48991 and n48496_not n48815_not ; n49247
g48992 and n48814_not n49247 ; n49248
g48993 and n49246_not n49248_not ; n49249
g48994 and b[7]_not n49249_not ; n49250
g48995 and n48515_not n48561 ; n49251
g48996 and n48557_not n49251 ; n49252
g48997 and n48558_not n48561_not ; n49253
g48998 and n49252_not n49253_not ; n49254
g48999 and n48816_not n49254_not ; n49255
g49000 and n48505_not n48815_not ; n49256
g49001 and n48814_not n49256 ; n49257
g49002 and n49255_not n49257_not ; n49258
g49003 and b[6]_not n49258_not ; n49259
g49004 and n48524_not n48556 ; n49260
g49005 and n48552_not n49260 ; n49261
g49006 and n48553_not n48556_not ; n49262
g49007 and n49261_not n49262_not ; n49263
g49008 and n48816_not n49263_not ; n49264
g49009 and n48514_not n48815_not ; n49265
g49010 and n48814_not n49265 ; n49266
g49011 and n49264_not n49266_not ; n49267
g49012 and b[5]_not n49267_not ; n49268
g49013 and n48532_not n48551 ; n49269
g49014 and n48547_not n49269 ; n49270
g49015 and n48548_not n48551_not ; n49271
g49016 and n49270_not n49271_not ; n49272
g49017 and n48816_not n49272_not ; n49273
g49018 and n48523_not n48815_not ; n49274
g49019 and n48814_not n49274 ; n49275
g49020 and n49273_not n49275_not ; n49276
g49021 and b[4]_not n49276_not ; n49277
g49022 and n48542_not n48546 ; n49278
g49023 and n48541_not n49278 ; n49279
g49024 and n48543_not n48546_not ; n49280
g49025 and n49279_not n49280_not ; n49281
g49026 and n48816_not n49281_not ; n49282
g49027 and n48531_not n48815_not ; n49283
g49028 and n48814_not n49283 ; n49284
g49029 and n49282_not n49284_not ; n49285
g49030 and b[3]_not n49285_not ; n49286
g49031 and n20502 n48539_not ; n49287
g49032 and n48537_not n49287 ; n49288
g49033 and n48541_not n49288_not ; n49289
g49034 and n48816_not n49289 ; n49290
g49035 and n48536_not n48815_not ; n49291
g49036 and n48814_not n49291 ; n49292
g49037 and n49290_not n49292_not ; n49293
g49038 and b[2]_not n49293_not ; n49294
g49039 and b[0] n48816_not ; n49295
g49040 and a[10] n49295_not ; n49296
g49041 and n20502 n48816_not ; n49297
g49042 and n49296_not n49297_not ; n49298
g49043 and b[1] n49298_not ; n49299
g49044 and b[1]_not n49297_not ; n49300
g49045 and n49296_not n49300 ; n49301
g49046 and n49299_not n49301_not ; n49302
g49047 and n21267_not n49302_not ; n49303
g49048 and b[1]_not n49298_not ; n49304
g49049 and n49303_not n49304_not ; n49305
g49050 and b[2] n49292_not ; n49306
g49051 and n49290_not n49306 ; n49307
g49052 and n49294_not n49307_not ; n49308
g49053 and n49305_not n49308 ; n49309
g49054 and n49294_not n49309_not ; n49310
g49055 and b[3] n49284_not ; n49311
g49056 and n49282_not n49311 ; n49312
g49057 and n49286_not n49312_not ; n49313
g49058 and n49310_not n49313 ; n49314
g49059 and n49286_not n49314_not ; n49315
g49060 and b[4] n49275_not ; n49316
g49061 and n49273_not n49316 ; n49317
g49062 and n49277_not n49317_not ; n49318
g49063 and n49315_not n49318 ; n49319
g49064 and n49277_not n49319_not ; n49320
g49065 and b[5] n49266_not ; n49321
g49066 and n49264_not n49321 ; n49322
g49067 and n49268_not n49322_not ; n49323
g49068 and n49320_not n49323 ; n49324
g49069 and n49268_not n49324_not ; n49325
g49070 and b[6] n49257_not ; n49326
g49071 and n49255_not n49326 ; n49327
g49072 and n49259_not n49327_not ; n49328
g49073 and n49325_not n49328 ; n49329
g49074 and n49259_not n49329_not ; n49330
g49075 and b[7] n49248_not ; n49331
g49076 and n49246_not n49331 ; n49332
g49077 and n49250_not n49332_not ; n49333
g49078 and n49330_not n49333 ; n49334
g49079 and n49250_not n49334_not ; n49335
g49080 and b[8] n49239_not ; n49336
g49081 and n49237_not n49336 ; n49337
g49082 and n49241_not n49337_not ; n49338
g49083 and n49335_not n49338 ; n49339
g49084 and n49241_not n49339_not ; n49340
g49085 and b[9] n49230_not ; n49341
g49086 and n49228_not n49341 ; n49342
g49087 and n49232_not n49342_not ; n49343
g49088 and n49340_not n49343 ; n49344
g49089 and n49232_not n49344_not ; n49345
g49090 and b[10] n49221_not ; n49346
g49091 and n49219_not n49346 ; n49347
g49092 and n49223_not n49347_not ; n49348
g49093 and n49345_not n49348 ; n49349
g49094 and n49223_not n49349_not ; n49350
g49095 and b[11] n49212_not ; n49351
g49096 and n49210_not n49351 ; n49352
g49097 and n49214_not n49352_not ; n49353
g49098 and n49350_not n49353 ; n49354
g49099 and n49214_not n49354_not ; n49355
g49100 and b[12] n49203_not ; n49356
g49101 and n49201_not n49356 ; n49357
g49102 and n49205_not n49357_not ; n49358
g49103 and n49355_not n49358 ; n49359
g49104 and n49205_not n49359_not ; n49360
g49105 and b[13] n49194_not ; n49361
g49106 and n49192_not n49361 ; n49362
g49107 and n49196_not n49362_not ; n49363
g49108 and n49360_not n49363 ; n49364
g49109 and n49196_not n49364_not ; n49365
g49110 and b[14] n49185_not ; n49366
g49111 and n49183_not n49366 ; n49367
g49112 and n49187_not n49367_not ; n49368
g49113 and n49365_not n49368 ; n49369
g49114 and n49187_not n49369_not ; n49370
g49115 and b[15] n49176_not ; n49371
g49116 and n49174_not n49371 ; n49372
g49117 and n49178_not n49372_not ; n49373
g49118 and n49370_not n49373 ; n49374
g49119 and n49178_not n49374_not ; n49375
g49120 and b[16] n49167_not ; n49376
g49121 and n49165_not n49376 ; n49377
g49122 and n49169_not n49377_not ; n49378
g49123 and n49375_not n49378 ; n49379
g49124 and n49169_not n49379_not ; n49380
g49125 and b[17] n49158_not ; n49381
g49126 and n49156_not n49381 ; n49382
g49127 and n49160_not n49382_not ; n49383
g49128 and n49380_not n49383 ; n49384
g49129 and n49160_not n49384_not ; n49385
g49130 and b[18] n49149_not ; n49386
g49131 and n49147_not n49386 ; n49387
g49132 and n49151_not n49387_not ; n49388
g49133 and n49385_not n49388 ; n49389
g49134 and n49151_not n49389_not ; n49390
g49135 and b[19] n49140_not ; n49391
g49136 and n49138_not n49391 ; n49392
g49137 and n49142_not n49392_not ; n49393
g49138 and n49390_not n49393 ; n49394
g49139 and n49142_not n49394_not ; n49395
g49140 and b[20] n49131_not ; n49396
g49141 and n49129_not n49396 ; n49397
g49142 and n49133_not n49397_not ; n49398
g49143 and n49395_not n49398 ; n49399
g49144 and n49133_not n49399_not ; n49400
g49145 and b[21] n49122_not ; n49401
g49146 and n49120_not n49401 ; n49402
g49147 and n49124_not n49402_not ; n49403
g49148 and n49400_not n49403 ; n49404
g49149 and n49124_not n49404_not ; n49405
g49150 and b[22] n49113_not ; n49406
g49151 and n49111_not n49406 ; n49407
g49152 and n49115_not n49407_not ; n49408
g49153 and n49405_not n49408 ; n49409
g49154 and n49115_not n49409_not ; n49410
g49155 and b[23] n49104_not ; n49411
g49156 and n49102_not n49411 ; n49412
g49157 and n49106_not n49412_not ; n49413
g49158 and n49410_not n49413 ; n49414
g49159 and n49106_not n49414_not ; n49415
g49160 and b[24] n49095_not ; n49416
g49161 and n49093_not n49416 ; n49417
g49162 and n49097_not n49417_not ; n49418
g49163 and n49415_not n49418 ; n49419
g49164 and n49097_not n49419_not ; n49420
g49165 and b[25] n49086_not ; n49421
g49166 and n49084_not n49421 ; n49422
g49167 and n49088_not n49422_not ; n49423
g49168 and n49420_not n49423 ; n49424
g49169 and n49088_not n49424_not ; n49425
g49170 and b[26] n49077_not ; n49426
g49171 and n49075_not n49426 ; n49427
g49172 and n49079_not n49427_not ; n49428
g49173 and n49425_not n49428 ; n49429
g49174 and n49079_not n49429_not ; n49430
g49175 and b[27] n49068_not ; n49431
g49176 and n49066_not n49431 ; n49432
g49177 and n49070_not n49432_not ; n49433
g49178 and n49430_not n49433 ; n49434
g49179 and n49070_not n49434_not ; n49435
g49180 and b[28] n49059_not ; n49436
g49181 and n49057_not n49436 ; n49437
g49182 and n49061_not n49437_not ; n49438
g49183 and n49435_not n49438 ; n49439
g49184 and n49061_not n49439_not ; n49440
g49185 and b[29] n49050_not ; n49441
g49186 and n49048_not n49441 ; n49442
g49187 and n49052_not n49442_not ; n49443
g49188 and n49440_not n49443 ; n49444
g49189 and n49052_not n49444_not ; n49445
g49190 and b[30] n49041_not ; n49446
g49191 and n49039_not n49446 ; n49447
g49192 and n49043_not n49447_not ; n49448
g49193 and n49445_not n49448 ; n49449
g49194 and n49043_not n49449_not ; n49450
g49195 and b[31] n49032_not ; n49451
g49196 and n49030_not n49451 ; n49452
g49197 and n49034_not n49452_not ; n49453
g49198 and n49450_not n49453 ; n49454
g49199 and n49034_not n49454_not ; n49455
g49200 and b[32] n49023_not ; n49456
g49201 and n49021_not n49456 ; n49457
g49202 and n49025_not n49457_not ; n49458
g49203 and n49455_not n49458 ; n49459
g49204 and n49025_not n49459_not ; n49460
g49205 and b[33] n49014_not ; n49461
g49206 and n49012_not n49461 ; n49462
g49207 and n49016_not n49462_not ; n49463
g49208 and n49460_not n49463 ; n49464
g49209 and n49016_not n49464_not ; n49465
g49210 and b[34] n49005_not ; n49466
g49211 and n49003_not n49466 ; n49467
g49212 and n49007_not n49467_not ; n49468
g49213 and n49465_not n49468 ; n49469
g49214 and n49007_not n49469_not ; n49470
g49215 and b[35] n48996_not ; n49471
g49216 and n48994_not n49471 ; n49472
g49217 and n48998_not n49472_not ; n49473
g49218 and n49470_not n49473 ; n49474
g49219 and n48998_not n49474_not ; n49475
g49220 and b[36] n48987_not ; n49476
g49221 and n48985_not n49476 ; n49477
g49222 and n48989_not n49477_not ; n49478
g49223 and n49475_not n49478 ; n49479
g49224 and n48989_not n49479_not ; n49480
g49225 and b[37] n48978_not ; n49481
g49226 and n48976_not n49481 ; n49482
g49227 and n48980_not n49482_not ; n49483
g49228 and n49480_not n49483 ; n49484
g49229 and n48980_not n49484_not ; n49485
g49230 and b[38] n48969_not ; n49486
g49231 and n48967_not n49486 ; n49487
g49232 and n48971_not n49487_not ; n49488
g49233 and n49485_not n49488 ; n49489
g49234 and n48971_not n49489_not ; n49490
g49235 and b[39] n48960_not ; n49491
g49236 and n48958_not n49491 ; n49492
g49237 and n48962_not n49492_not ; n49493
g49238 and n49490_not n49493 ; n49494
g49239 and n48962_not n49494_not ; n49495
g49240 and b[40] n48951_not ; n49496
g49241 and n48949_not n49496 ; n49497
g49242 and n48953_not n49497_not ; n49498
g49243 and n49495_not n49498 ; n49499
g49244 and n48953_not n49499_not ; n49500
g49245 and b[41] n48942_not ; n49501
g49246 and n48940_not n49501 ; n49502
g49247 and n48944_not n49502_not ; n49503
g49248 and n49500_not n49503 ; n49504
g49249 and n48944_not n49504_not ; n49505
g49250 and b[42] n48933_not ; n49506
g49251 and n48931_not n49506 ; n49507
g49252 and n48935_not n49507_not ; n49508
g49253 and n49505_not n49508 ; n49509
g49254 and n48935_not n49509_not ; n49510
g49255 and b[43] n48924_not ; n49511
g49256 and n48922_not n49511 ; n49512
g49257 and n48926_not n49512_not ; n49513
g49258 and n49510_not n49513 ; n49514
g49259 and n48926_not n49514_not ; n49515
g49260 and b[44] n48915_not ; n49516
g49261 and n48913_not n49516 ; n49517
g49262 and n48917_not n49517_not ; n49518
g49263 and n49515_not n49518 ; n49519
g49264 and n48917_not n49519_not ; n49520
g49265 and b[45] n48906_not ; n49521
g49266 and n48904_not n49521 ; n49522
g49267 and n48908_not n49522_not ; n49523
g49268 and n49520_not n49523 ; n49524
g49269 and n48908_not n49524_not ; n49525
g49270 and b[46] n48897_not ; n49526
g49271 and n48895_not n49526 ; n49527
g49272 and n48899_not n49527_not ; n49528
g49273 and n49525_not n49528 ; n49529
g49274 and n48899_not n49529_not ; n49530
g49275 and b[47] n48888_not ; n49531
g49276 and n48886_not n49531 ; n49532
g49277 and n48890_not n49532_not ; n49533
g49278 and n49530_not n49533 ; n49534
g49279 and n48890_not n49534_not ; n49535
g49280 and b[48] n48879_not ; n49536
g49281 and n48877_not n49536 ; n49537
g49282 and n48881_not n49537_not ; n49538
g49283 and n49535_not n49538 ; n49539
g49284 and n48881_not n49539_not ; n49540
g49285 and b[49] n48870_not ; n49541
g49286 and n48868_not n49541 ; n49542
g49287 and n48872_not n49542_not ; n49543
g49288 and n49540_not n49543 ; n49544
g49289 and n48872_not n49544_not ; n49545
g49290 and b[50] n48861_not ; n49546
g49291 and n48859_not n49546 ; n49547
g49292 and n48863_not n49547_not ; n49548
g49293 and n49545_not n49548 ; n49549
g49294 and n48863_not n49549_not ; n49550
g49295 and b[51] n48852_not ; n49551
g49296 and n48850_not n49551 ; n49552
g49297 and n48854_not n49552_not ; n49553
g49298 and n49550_not n49553 ; n49554
g49299 and n48854_not n49554_not ; n49555
g49300 and b[52] n48843_not ; n49556
g49301 and n48841_not n49556 ; n49557
g49302 and n48845_not n49557_not ; n49558
g49303 and n49555_not n49558 ; n49559
g49304 and n48845_not n49559_not ; n49560
g49305 and b[53] n48823_not ; n49561
g49306 and n48821_not n49561 ; n49562
g49307 and n48836_not n49562_not ; n49563
g49308 and n49560_not n49563 ; n49564
g49309 and n48836_not n49564_not ; n49565
g49310 and b[54] n48833_not ; n49566
g49311 and n48831_not n49566 ; n49567
g49312 and n48835_not n49567_not ; n49568
g49313 and n49565_not n49568 ; n49569
g49314 and n48835_not n49569_not ; n49570
g49315 and n21537 n49570_not ; n49571
g49316 and n48824_not n49571_not ; n49572
g49317 and n48845_not n49563 ; n49573
g49318 and n49559_not n49573 ; n49574
g49319 and n49560_not n49563_not ; n49575
g49320 and n49574_not n49575_not ; n49576
g49321 and n21537 n49576_not ; n49577
g49322 and n49570_not n49577 ; n49578
g49323 and n49572_not n49578_not ; n49579
g49324 and b[54]_not n49579_not ; n49580
g49325 and n48844_not n49571_not ; n49581
g49326 and n48854_not n49558 ; n49582
g49327 and n49554_not n49582 ; n49583
g49328 and n49555_not n49558_not ; n49584
g49329 and n49583_not n49584_not ; n49585
g49330 and n21537 n49585_not ; n49586
g49331 and n49570_not n49586 ; n49587
g49332 and n49581_not n49587_not ; n49588
g49333 and b[53]_not n49588_not ; n49589
g49334 and n48853_not n49571_not ; n49590
g49335 and n48863_not n49553 ; n49591
g49336 and n49549_not n49591 ; n49592
g49337 and n49550_not n49553_not ; n49593
g49338 and n49592_not n49593_not ; n49594
g49339 and n21537 n49594_not ; n49595
g49340 and n49570_not n49595 ; n49596
g49341 and n49590_not n49596_not ; n49597
g49342 and b[52]_not n49597_not ; n49598
g49343 and n48862_not n49571_not ; n49599
g49344 and n48872_not n49548 ; n49600
g49345 and n49544_not n49600 ; n49601
g49346 and n49545_not n49548_not ; n49602
g49347 and n49601_not n49602_not ; n49603
g49348 and n21537 n49603_not ; n49604
g49349 and n49570_not n49604 ; n49605
g49350 and n49599_not n49605_not ; n49606
g49351 and b[51]_not n49606_not ; n49607
g49352 and n48871_not n49571_not ; n49608
g49353 and n48881_not n49543 ; n49609
g49354 and n49539_not n49609 ; n49610
g49355 and n49540_not n49543_not ; n49611
g49356 and n49610_not n49611_not ; n49612
g49357 and n21537 n49612_not ; n49613
g49358 and n49570_not n49613 ; n49614
g49359 and n49608_not n49614_not ; n49615
g49360 and b[50]_not n49615_not ; n49616
g49361 and n48880_not n49571_not ; n49617
g49362 and n48890_not n49538 ; n49618
g49363 and n49534_not n49618 ; n49619
g49364 and n49535_not n49538_not ; n49620
g49365 and n49619_not n49620_not ; n49621
g49366 and n21537 n49621_not ; n49622
g49367 and n49570_not n49622 ; n49623
g49368 and n49617_not n49623_not ; n49624
g49369 and b[49]_not n49624_not ; n49625
g49370 and n48889_not n49571_not ; n49626
g49371 and n48899_not n49533 ; n49627
g49372 and n49529_not n49627 ; n49628
g49373 and n49530_not n49533_not ; n49629
g49374 and n49628_not n49629_not ; n49630
g49375 and n21537 n49630_not ; n49631
g49376 and n49570_not n49631 ; n49632
g49377 and n49626_not n49632_not ; n49633
g49378 and b[48]_not n49633_not ; n49634
g49379 and n48898_not n49571_not ; n49635
g49380 and n48908_not n49528 ; n49636
g49381 and n49524_not n49636 ; n49637
g49382 and n49525_not n49528_not ; n49638
g49383 and n49637_not n49638_not ; n49639
g49384 and n21537 n49639_not ; n49640
g49385 and n49570_not n49640 ; n49641
g49386 and n49635_not n49641_not ; n49642
g49387 and b[47]_not n49642_not ; n49643
g49388 and n48907_not n49571_not ; n49644
g49389 and n48917_not n49523 ; n49645
g49390 and n49519_not n49645 ; n49646
g49391 and n49520_not n49523_not ; n49647
g49392 and n49646_not n49647_not ; n49648
g49393 and n21537 n49648_not ; n49649
g49394 and n49570_not n49649 ; n49650
g49395 and n49644_not n49650_not ; n49651
g49396 and b[46]_not n49651_not ; n49652
g49397 and n48916_not n49571_not ; n49653
g49398 and n48926_not n49518 ; n49654
g49399 and n49514_not n49654 ; n49655
g49400 and n49515_not n49518_not ; n49656
g49401 and n49655_not n49656_not ; n49657
g49402 and n21537 n49657_not ; n49658
g49403 and n49570_not n49658 ; n49659
g49404 and n49653_not n49659_not ; n49660
g49405 and b[45]_not n49660_not ; n49661
g49406 and n48925_not n49571_not ; n49662
g49407 and n48935_not n49513 ; n49663
g49408 and n49509_not n49663 ; n49664
g49409 and n49510_not n49513_not ; n49665
g49410 and n49664_not n49665_not ; n49666
g49411 and n21537 n49666_not ; n49667
g49412 and n49570_not n49667 ; n49668
g49413 and n49662_not n49668_not ; n49669
g49414 and b[44]_not n49669_not ; n49670
g49415 and n48934_not n49571_not ; n49671
g49416 and n48944_not n49508 ; n49672
g49417 and n49504_not n49672 ; n49673
g49418 and n49505_not n49508_not ; n49674
g49419 and n49673_not n49674_not ; n49675
g49420 and n21537 n49675_not ; n49676
g49421 and n49570_not n49676 ; n49677
g49422 and n49671_not n49677_not ; n49678
g49423 and b[43]_not n49678_not ; n49679
g49424 and n48943_not n49571_not ; n49680
g49425 and n48953_not n49503 ; n49681
g49426 and n49499_not n49681 ; n49682
g49427 and n49500_not n49503_not ; n49683
g49428 and n49682_not n49683_not ; n49684
g49429 and n21537 n49684_not ; n49685
g49430 and n49570_not n49685 ; n49686
g49431 and n49680_not n49686_not ; n49687
g49432 and b[42]_not n49687_not ; n49688
g49433 and n48952_not n49571_not ; n49689
g49434 and n48962_not n49498 ; n49690
g49435 and n49494_not n49690 ; n49691
g49436 and n49495_not n49498_not ; n49692
g49437 and n49691_not n49692_not ; n49693
g49438 and n21537 n49693_not ; n49694
g49439 and n49570_not n49694 ; n49695
g49440 and n49689_not n49695_not ; n49696
g49441 and b[41]_not n49696_not ; n49697
g49442 and n48961_not n49571_not ; n49698
g49443 and n48971_not n49493 ; n49699
g49444 and n49489_not n49699 ; n49700
g49445 and n49490_not n49493_not ; n49701
g49446 and n49700_not n49701_not ; n49702
g49447 and n21537 n49702_not ; n49703
g49448 and n49570_not n49703 ; n49704
g49449 and n49698_not n49704_not ; n49705
g49450 and b[40]_not n49705_not ; n49706
g49451 and n48970_not n49571_not ; n49707
g49452 and n48980_not n49488 ; n49708
g49453 and n49484_not n49708 ; n49709
g49454 and n49485_not n49488_not ; n49710
g49455 and n49709_not n49710_not ; n49711
g49456 and n21537 n49711_not ; n49712
g49457 and n49570_not n49712 ; n49713
g49458 and n49707_not n49713_not ; n49714
g49459 and b[39]_not n49714_not ; n49715
g49460 and n48979_not n49571_not ; n49716
g49461 and n48989_not n49483 ; n49717
g49462 and n49479_not n49717 ; n49718
g49463 and n49480_not n49483_not ; n49719
g49464 and n49718_not n49719_not ; n49720
g49465 and n21537 n49720_not ; n49721
g49466 and n49570_not n49721 ; n49722
g49467 and n49716_not n49722_not ; n49723
g49468 and b[38]_not n49723_not ; n49724
g49469 and n48988_not n49571_not ; n49725
g49470 and n48998_not n49478 ; n49726
g49471 and n49474_not n49726 ; n49727
g49472 and n49475_not n49478_not ; n49728
g49473 and n49727_not n49728_not ; n49729
g49474 and n21537 n49729_not ; n49730
g49475 and n49570_not n49730 ; n49731
g49476 and n49725_not n49731_not ; n49732
g49477 and b[37]_not n49732_not ; n49733
g49478 and n48997_not n49571_not ; n49734
g49479 and n49007_not n49473 ; n49735
g49480 and n49469_not n49735 ; n49736
g49481 and n49470_not n49473_not ; n49737
g49482 and n49736_not n49737_not ; n49738
g49483 and n21537 n49738_not ; n49739
g49484 and n49570_not n49739 ; n49740
g49485 and n49734_not n49740_not ; n49741
g49486 and b[36]_not n49741_not ; n49742
g49487 and n49006_not n49571_not ; n49743
g49488 and n49016_not n49468 ; n49744
g49489 and n49464_not n49744 ; n49745
g49490 and n49465_not n49468_not ; n49746
g49491 and n49745_not n49746_not ; n49747
g49492 and n21537 n49747_not ; n49748
g49493 and n49570_not n49748 ; n49749
g49494 and n49743_not n49749_not ; n49750
g49495 and b[35]_not n49750_not ; n49751
g49496 and n49015_not n49571_not ; n49752
g49497 and n49025_not n49463 ; n49753
g49498 and n49459_not n49753 ; n49754
g49499 and n49460_not n49463_not ; n49755
g49500 and n49754_not n49755_not ; n49756
g49501 and n21537 n49756_not ; n49757
g49502 and n49570_not n49757 ; n49758
g49503 and n49752_not n49758_not ; n49759
g49504 and b[34]_not n49759_not ; n49760
g49505 and n49024_not n49571_not ; n49761
g49506 and n49034_not n49458 ; n49762
g49507 and n49454_not n49762 ; n49763
g49508 and n49455_not n49458_not ; n49764
g49509 and n49763_not n49764_not ; n49765
g49510 and n21537 n49765_not ; n49766
g49511 and n49570_not n49766 ; n49767
g49512 and n49761_not n49767_not ; n49768
g49513 and b[33]_not n49768_not ; n49769
g49514 and n49033_not n49571_not ; n49770
g49515 and n49043_not n49453 ; n49771
g49516 and n49449_not n49771 ; n49772
g49517 and n49450_not n49453_not ; n49773
g49518 and n49772_not n49773_not ; n49774
g49519 and n21537 n49774_not ; n49775
g49520 and n49570_not n49775 ; n49776
g49521 and n49770_not n49776_not ; n49777
g49522 and b[32]_not n49777_not ; n49778
g49523 and n49042_not n49571_not ; n49779
g49524 and n49052_not n49448 ; n49780
g49525 and n49444_not n49780 ; n49781
g49526 and n49445_not n49448_not ; n49782
g49527 and n49781_not n49782_not ; n49783
g49528 and n21537 n49783_not ; n49784
g49529 and n49570_not n49784 ; n49785
g49530 and n49779_not n49785_not ; n49786
g49531 and b[31]_not n49786_not ; n49787
g49532 and n49051_not n49571_not ; n49788
g49533 and n49061_not n49443 ; n49789
g49534 and n49439_not n49789 ; n49790
g49535 and n49440_not n49443_not ; n49791
g49536 and n49790_not n49791_not ; n49792
g49537 and n21537 n49792_not ; n49793
g49538 and n49570_not n49793 ; n49794
g49539 and n49788_not n49794_not ; n49795
g49540 and b[30]_not n49795_not ; n49796
g49541 and n49060_not n49571_not ; n49797
g49542 and n49070_not n49438 ; n49798
g49543 and n49434_not n49798 ; n49799
g49544 and n49435_not n49438_not ; n49800
g49545 and n49799_not n49800_not ; n49801
g49546 and n21537 n49801_not ; n49802
g49547 and n49570_not n49802 ; n49803
g49548 and n49797_not n49803_not ; n49804
g49549 and b[29]_not n49804_not ; n49805
g49550 and n49069_not n49571_not ; n49806
g49551 and n49079_not n49433 ; n49807
g49552 and n49429_not n49807 ; n49808
g49553 and n49430_not n49433_not ; n49809
g49554 and n49808_not n49809_not ; n49810
g49555 and n21537 n49810_not ; n49811
g49556 and n49570_not n49811 ; n49812
g49557 and n49806_not n49812_not ; n49813
g49558 and b[28]_not n49813_not ; n49814
g49559 and n49078_not n49571_not ; n49815
g49560 and n49088_not n49428 ; n49816
g49561 and n49424_not n49816 ; n49817
g49562 and n49425_not n49428_not ; n49818
g49563 and n49817_not n49818_not ; n49819
g49564 and n21537 n49819_not ; n49820
g49565 and n49570_not n49820 ; n49821
g49566 and n49815_not n49821_not ; n49822
g49567 and b[27]_not n49822_not ; n49823
g49568 and n49087_not n49571_not ; n49824
g49569 and n49097_not n49423 ; n49825
g49570 and n49419_not n49825 ; n49826
g49571 and n49420_not n49423_not ; n49827
g49572 and n49826_not n49827_not ; n49828
g49573 and n21537 n49828_not ; n49829
g49574 and n49570_not n49829 ; n49830
g49575 and n49824_not n49830_not ; n49831
g49576 and b[26]_not n49831_not ; n49832
g49577 and n49096_not n49571_not ; n49833
g49578 and n49106_not n49418 ; n49834
g49579 and n49414_not n49834 ; n49835
g49580 and n49415_not n49418_not ; n49836
g49581 and n49835_not n49836_not ; n49837
g49582 and n21537 n49837_not ; n49838
g49583 and n49570_not n49838 ; n49839
g49584 and n49833_not n49839_not ; n49840
g49585 and b[25]_not n49840_not ; n49841
g49586 and n49105_not n49571_not ; n49842
g49587 and n49115_not n49413 ; n49843
g49588 and n49409_not n49843 ; n49844
g49589 and n49410_not n49413_not ; n49845
g49590 and n49844_not n49845_not ; n49846
g49591 and n21537 n49846_not ; n49847
g49592 and n49570_not n49847 ; n49848
g49593 and n49842_not n49848_not ; n49849
g49594 and b[24]_not n49849_not ; n49850
g49595 and n49114_not n49571_not ; n49851
g49596 and n49124_not n49408 ; n49852
g49597 and n49404_not n49852 ; n49853
g49598 and n49405_not n49408_not ; n49854
g49599 and n49853_not n49854_not ; n49855
g49600 and n21537 n49855_not ; n49856
g49601 and n49570_not n49856 ; n49857
g49602 and n49851_not n49857_not ; n49858
g49603 and b[23]_not n49858_not ; n49859
g49604 and n49123_not n49571_not ; n49860
g49605 and n49133_not n49403 ; n49861
g49606 and n49399_not n49861 ; n49862
g49607 and n49400_not n49403_not ; n49863
g49608 and n49862_not n49863_not ; n49864
g49609 and n21537 n49864_not ; n49865
g49610 and n49570_not n49865 ; n49866
g49611 and n49860_not n49866_not ; n49867
g49612 and b[22]_not n49867_not ; n49868
g49613 and n49132_not n49571_not ; n49869
g49614 and n49142_not n49398 ; n49870
g49615 and n49394_not n49870 ; n49871
g49616 and n49395_not n49398_not ; n49872
g49617 and n49871_not n49872_not ; n49873
g49618 and n21537 n49873_not ; n49874
g49619 and n49570_not n49874 ; n49875
g49620 and n49869_not n49875_not ; n49876
g49621 and b[21]_not n49876_not ; n49877
g49622 and n49141_not n49571_not ; n49878
g49623 and n49151_not n49393 ; n49879
g49624 and n49389_not n49879 ; n49880
g49625 and n49390_not n49393_not ; n49881
g49626 and n49880_not n49881_not ; n49882
g49627 and n21537 n49882_not ; n49883
g49628 and n49570_not n49883 ; n49884
g49629 and n49878_not n49884_not ; n49885
g49630 and b[20]_not n49885_not ; n49886
g49631 and n49150_not n49571_not ; n49887
g49632 and n49160_not n49388 ; n49888
g49633 and n49384_not n49888 ; n49889
g49634 and n49385_not n49388_not ; n49890
g49635 and n49889_not n49890_not ; n49891
g49636 and n21537 n49891_not ; n49892
g49637 and n49570_not n49892 ; n49893
g49638 and n49887_not n49893_not ; n49894
g49639 and b[19]_not n49894_not ; n49895
g49640 and n49159_not n49571_not ; n49896
g49641 and n49169_not n49383 ; n49897
g49642 and n49379_not n49897 ; n49898
g49643 and n49380_not n49383_not ; n49899
g49644 and n49898_not n49899_not ; n49900
g49645 and n21537 n49900_not ; n49901
g49646 and n49570_not n49901 ; n49902
g49647 and n49896_not n49902_not ; n49903
g49648 and b[18]_not n49903_not ; n49904
g49649 and n49168_not n49571_not ; n49905
g49650 and n49178_not n49378 ; n49906
g49651 and n49374_not n49906 ; n49907
g49652 and n49375_not n49378_not ; n49908
g49653 and n49907_not n49908_not ; n49909
g49654 and n21537 n49909_not ; n49910
g49655 and n49570_not n49910 ; n49911
g49656 and n49905_not n49911_not ; n49912
g49657 and b[17]_not n49912_not ; n49913
g49658 and n49177_not n49571_not ; n49914
g49659 and n49187_not n49373 ; n49915
g49660 and n49369_not n49915 ; n49916
g49661 and n49370_not n49373_not ; n49917
g49662 and n49916_not n49917_not ; n49918
g49663 and n21537 n49918_not ; n49919
g49664 and n49570_not n49919 ; n49920
g49665 and n49914_not n49920_not ; n49921
g49666 and b[16]_not n49921_not ; n49922
g49667 and n49186_not n49571_not ; n49923
g49668 and n49196_not n49368 ; n49924
g49669 and n49364_not n49924 ; n49925
g49670 and n49365_not n49368_not ; n49926
g49671 and n49925_not n49926_not ; n49927
g49672 and n21537 n49927_not ; n49928
g49673 and n49570_not n49928 ; n49929
g49674 and n49923_not n49929_not ; n49930
g49675 and b[15]_not n49930_not ; n49931
g49676 and n49195_not n49571_not ; n49932
g49677 and n49205_not n49363 ; n49933
g49678 and n49359_not n49933 ; n49934
g49679 and n49360_not n49363_not ; n49935
g49680 and n49934_not n49935_not ; n49936
g49681 and n21537 n49936_not ; n49937
g49682 and n49570_not n49937 ; n49938
g49683 and n49932_not n49938_not ; n49939
g49684 and b[14]_not n49939_not ; n49940
g49685 and n49204_not n49571_not ; n49941
g49686 and n49214_not n49358 ; n49942
g49687 and n49354_not n49942 ; n49943
g49688 and n49355_not n49358_not ; n49944
g49689 and n49943_not n49944_not ; n49945
g49690 and n21537 n49945_not ; n49946
g49691 and n49570_not n49946 ; n49947
g49692 and n49941_not n49947_not ; n49948
g49693 and b[13]_not n49948_not ; n49949
g49694 and n49213_not n49571_not ; n49950
g49695 and n49223_not n49353 ; n49951
g49696 and n49349_not n49951 ; n49952
g49697 and n49350_not n49353_not ; n49953
g49698 and n49952_not n49953_not ; n49954
g49699 and n21537 n49954_not ; n49955
g49700 and n49570_not n49955 ; n49956
g49701 and n49950_not n49956_not ; n49957
g49702 and b[12]_not n49957_not ; n49958
g49703 and n49222_not n49571_not ; n49959
g49704 and n49232_not n49348 ; n49960
g49705 and n49344_not n49960 ; n49961
g49706 and n49345_not n49348_not ; n49962
g49707 and n49961_not n49962_not ; n49963
g49708 and n21537 n49963_not ; n49964
g49709 and n49570_not n49964 ; n49965
g49710 and n49959_not n49965_not ; n49966
g49711 and b[11]_not n49966_not ; n49967
g49712 and n49231_not n49571_not ; n49968
g49713 and n49241_not n49343 ; n49969
g49714 and n49339_not n49969 ; n49970
g49715 and n49340_not n49343_not ; n49971
g49716 and n49970_not n49971_not ; n49972
g49717 and n21537 n49972_not ; n49973
g49718 and n49570_not n49973 ; n49974
g49719 and n49968_not n49974_not ; n49975
g49720 and b[10]_not n49975_not ; n49976
g49721 and n49240_not n49571_not ; n49977
g49722 and n49250_not n49338 ; n49978
g49723 and n49334_not n49978 ; n49979
g49724 and n49335_not n49338_not ; n49980
g49725 and n49979_not n49980_not ; n49981
g49726 and n21537 n49981_not ; n49982
g49727 and n49570_not n49982 ; n49983
g49728 and n49977_not n49983_not ; n49984
g49729 and b[9]_not n49984_not ; n49985
g49730 and n49249_not n49571_not ; n49986
g49731 and n49259_not n49333 ; n49987
g49732 and n49329_not n49987 ; n49988
g49733 and n49330_not n49333_not ; n49989
g49734 and n49988_not n49989_not ; n49990
g49735 and n21537 n49990_not ; n49991
g49736 and n49570_not n49991 ; n49992
g49737 and n49986_not n49992_not ; n49993
g49738 and b[8]_not n49993_not ; n49994
g49739 and n49258_not n49571_not ; n49995
g49740 and n49268_not n49328 ; n49996
g49741 and n49324_not n49996 ; n49997
g49742 and n49325_not n49328_not ; n49998
g49743 and n49997_not n49998_not ; n49999
g49744 and n21537 n49999_not ; n50000
g49745 and n49570_not n50000 ; n50001
g49746 and n49995_not n50001_not ; n50002
g49747 and b[7]_not n50002_not ; n50003
g49748 and n49267_not n49571_not ; n50004
g49749 and n49277_not n49323 ; n50005
g49750 and n49319_not n50005 ; n50006
g49751 and n49320_not n49323_not ; n50007
g49752 and n50006_not n50007_not ; n50008
g49753 and n21537 n50008_not ; n50009
g49754 and n49570_not n50009 ; n50010
g49755 and n50004_not n50010_not ; n50011
g49756 and b[6]_not n50011_not ; n50012
g49757 and n49276_not n49571_not ; n50013
g49758 and n49286_not n49318 ; n50014
g49759 and n49314_not n50014 ; n50015
g49760 and n49315_not n49318_not ; n50016
g49761 and n50015_not n50016_not ; n50017
g49762 and n21537 n50017_not ; n50018
g49763 and n49570_not n50018 ; n50019
g49764 and n50013_not n50019_not ; n50020
g49765 and b[5]_not n50020_not ; n50021
g49766 and n49285_not n49571_not ; n50022
g49767 and n49294_not n49313 ; n50023
g49768 and n49309_not n50023 ; n50024
g49769 and n49310_not n49313_not ; n50025
g49770 and n50024_not n50025_not ; n50026
g49771 and n21537 n50026_not ; n50027
g49772 and n49570_not n50027 ; n50028
g49773 and n50022_not n50028_not ; n50029
g49774 and b[4]_not n50029_not ; n50030
g49775 and n49293_not n49571_not ; n50031
g49776 and n49304_not n49308 ; n50032
g49777 and n49303_not n50032 ; n50033
g49778 and n49305_not n49308_not ; n50034
g49779 and n50033_not n50034_not ; n50035
g49780 and n21537 n50035_not ; n50036
g49781 and n49570_not n50036 ; n50037
g49782 and n50031_not n50037_not ; n50038
g49783 and b[3]_not n50038_not ; n50039
g49784 and n49298_not n49571_not ; n50040
g49785 and n21267 n49301_not ; n50041
g49786 and n49299_not n50041 ; n50042
g49787 and n21537 n50042_not ; n50043
g49788 and n49303_not n50043 ; n50044
g49789 and n49570_not n50044 ; n50045
g49790 and n50040_not n50045_not ; n50046
g49791 and b[2]_not n50046_not ; n50047
g49792 and n22017 n49570_not ; n50048
g49793 and a[9] n50048_not ; n50049
g49794 and n22022 n49570_not ; n50050
g49795 and n50049_not n50050_not ; n50051
g49796 and b[1] n50051_not ; n50052
g49797 and b[1]_not n50050_not ; n50053
g49798 and n50049_not n50053 ; n50054
g49799 and n50052_not n50054_not ; n50055
g49800 and n22029_not n50055_not ; n50056
g49801 and b[1]_not n50051_not ; n50057
g49802 and n50056_not n50057_not ; n50058
g49803 and b[2] n50045_not ; n50059
g49804 and n50040_not n50059 ; n50060
g49805 and n50047_not n50060_not ; n50061
g49806 and n50058_not n50061 ; n50062
g49807 and n50047_not n50062_not ; n50063
g49808 and b[3] n50037_not ; n50064
g49809 and n50031_not n50064 ; n50065
g49810 and n50039_not n50065_not ; n50066
g49811 and n50063_not n50066 ; n50067
g49812 and n50039_not n50067_not ; n50068
g49813 and b[4] n50028_not ; n50069
g49814 and n50022_not n50069 ; n50070
g49815 and n50030_not n50070_not ; n50071
g49816 and n50068_not n50071 ; n50072
g49817 and n50030_not n50072_not ; n50073
g49818 and b[5] n50019_not ; n50074
g49819 and n50013_not n50074 ; n50075
g49820 and n50021_not n50075_not ; n50076
g49821 and n50073_not n50076 ; n50077
g49822 and n50021_not n50077_not ; n50078
g49823 and b[6] n50010_not ; n50079
g49824 and n50004_not n50079 ; n50080
g49825 and n50012_not n50080_not ; n50081
g49826 and n50078_not n50081 ; n50082
g49827 and n50012_not n50082_not ; n50083
g49828 and b[7] n50001_not ; n50084
g49829 and n49995_not n50084 ; n50085
g49830 and n50003_not n50085_not ; n50086
g49831 and n50083_not n50086 ; n50087
g49832 and n50003_not n50087_not ; n50088
g49833 and b[8] n49992_not ; n50089
g49834 and n49986_not n50089 ; n50090
g49835 and n49994_not n50090_not ; n50091
g49836 and n50088_not n50091 ; n50092
g49837 and n49994_not n50092_not ; n50093
g49838 and b[9] n49983_not ; n50094
g49839 and n49977_not n50094 ; n50095
g49840 and n49985_not n50095_not ; n50096
g49841 and n50093_not n50096 ; n50097
g49842 and n49985_not n50097_not ; n50098
g49843 and b[10] n49974_not ; n50099
g49844 and n49968_not n50099 ; n50100
g49845 and n49976_not n50100_not ; n50101
g49846 and n50098_not n50101 ; n50102
g49847 and n49976_not n50102_not ; n50103
g49848 and b[11] n49965_not ; n50104
g49849 and n49959_not n50104 ; n50105
g49850 and n49967_not n50105_not ; n50106
g49851 and n50103_not n50106 ; n50107
g49852 and n49967_not n50107_not ; n50108
g49853 and b[12] n49956_not ; n50109
g49854 and n49950_not n50109 ; n50110
g49855 and n49958_not n50110_not ; n50111
g49856 and n50108_not n50111 ; n50112
g49857 and n49958_not n50112_not ; n50113
g49858 and b[13] n49947_not ; n50114
g49859 and n49941_not n50114 ; n50115
g49860 and n49949_not n50115_not ; n50116
g49861 and n50113_not n50116 ; n50117
g49862 and n49949_not n50117_not ; n50118
g49863 and b[14] n49938_not ; n50119
g49864 and n49932_not n50119 ; n50120
g49865 and n49940_not n50120_not ; n50121
g49866 and n50118_not n50121 ; n50122
g49867 and n49940_not n50122_not ; n50123
g49868 and b[15] n49929_not ; n50124
g49869 and n49923_not n50124 ; n50125
g49870 and n49931_not n50125_not ; n50126
g49871 and n50123_not n50126 ; n50127
g49872 and n49931_not n50127_not ; n50128
g49873 and b[16] n49920_not ; n50129
g49874 and n49914_not n50129 ; n50130
g49875 and n49922_not n50130_not ; n50131
g49876 and n50128_not n50131 ; n50132
g49877 and n49922_not n50132_not ; n50133
g49878 and b[17] n49911_not ; n50134
g49879 and n49905_not n50134 ; n50135
g49880 and n49913_not n50135_not ; n50136
g49881 and n50133_not n50136 ; n50137
g49882 and n49913_not n50137_not ; n50138
g49883 and b[18] n49902_not ; n50139
g49884 and n49896_not n50139 ; n50140
g49885 and n49904_not n50140_not ; n50141
g49886 and n50138_not n50141 ; n50142
g49887 and n49904_not n50142_not ; n50143
g49888 and b[19] n49893_not ; n50144
g49889 and n49887_not n50144 ; n50145
g49890 and n49895_not n50145_not ; n50146
g49891 and n50143_not n50146 ; n50147
g49892 and n49895_not n50147_not ; n50148
g49893 and b[20] n49884_not ; n50149
g49894 and n49878_not n50149 ; n50150
g49895 and n49886_not n50150_not ; n50151
g49896 and n50148_not n50151 ; n50152
g49897 and n49886_not n50152_not ; n50153
g49898 and b[21] n49875_not ; n50154
g49899 and n49869_not n50154 ; n50155
g49900 and n49877_not n50155_not ; n50156
g49901 and n50153_not n50156 ; n50157
g49902 and n49877_not n50157_not ; n50158
g49903 and b[22] n49866_not ; n50159
g49904 and n49860_not n50159 ; n50160
g49905 and n49868_not n50160_not ; n50161
g49906 and n50158_not n50161 ; n50162
g49907 and n49868_not n50162_not ; n50163
g49908 and b[23] n49857_not ; n50164
g49909 and n49851_not n50164 ; n50165
g49910 and n49859_not n50165_not ; n50166
g49911 and n50163_not n50166 ; n50167
g49912 and n49859_not n50167_not ; n50168
g49913 and b[24] n49848_not ; n50169
g49914 and n49842_not n50169 ; n50170
g49915 and n49850_not n50170_not ; n50171
g49916 and n50168_not n50171 ; n50172
g49917 and n49850_not n50172_not ; n50173
g49918 and b[25] n49839_not ; n50174
g49919 and n49833_not n50174 ; n50175
g49920 and n49841_not n50175_not ; n50176
g49921 and n50173_not n50176 ; n50177
g49922 and n49841_not n50177_not ; n50178
g49923 and b[26] n49830_not ; n50179
g49924 and n49824_not n50179 ; n50180
g49925 and n49832_not n50180_not ; n50181
g49926 and n50178_not n50181 ; n50182
g49927 and n49832_not n50182_not ; n50183
g49928 and b[27] n49821_not ; n50184
g49929 and n49815_not n50184 ; n50185
g49930 and n49823_not n50185_not ; n50186
g49931 and n50183_not n50186 ; n50187
g49932 and n49823_not n50187_not ; n50188
g49933 and b[28] n49812_not ; n50189
g49934 and n49806_not n50189 ; n50190
g49935 and n49814_not n50190_not ; n50191
g49936 and n50188_not n50191 ; n50192
g49937 and n49814_not n50192_not ; n50193
g49938 and b[29] n49803_not ; n50194
g49939 and n49797_not n50194 ; n50195
g49940 and n49805_not n50195_not ; n50196
g49941 and n50193_not n50196 ; n50197
g49942 and n49805_not n50197_not ; n50198
g49943 and b[30] n49794_not ; n50199
g49944 and n49788_not n50199 ; n50200
g49945 and n49796_not n50200_not ; n50201
g49946 and n50198_not n50201 ; n50202
g49947 and n49796_not n50202_not ; n50203
g49948 and b[31] n49785_not ; n50204
g49949 and n49779_not n50204 ; n50205
g49950 and n49787_not n50205_not ; n50206
g49951 and n50203_not n50206 ; n50207
g49952 and n49787_not n50207_not ; n50208
g49953 and b[32] n49776_not ; n50209
g49954 and n49770_not n50209 ; n50210
g49955 and n49778_not n50210_not ; n50211
g49956 and n50208_not n50211 ; n50212
g49957 and n49778_not n50212_not ; n50213
g49958 and b[33] n49767_not ; n50214
g49959 and n49761_not n50214 ; n50215
g49960 and n49769_not n50215_not ; n50216
g49961 and n50213_not n50216 ; n50217
g49962 and n49769_not n50217_not ; n50218
g49963 and b[34] n49758_not ; n50219
g49964 and n49752_not n50219 ; n50220
g49965 and n49760_not n50220_not ; n50221
g49966 and n50218_not n50221 ; n50222
g49967 and n49760_not n50222_not ; n50223
g49968 and b[35] n49749_not ; n50224
g49969 and n49743_not n50224 ; n50225
g49970 and n49751_not n50225_not ; n50226
g49971 and n50223_not n50226 ; n50227
g49972 and n49751_not n50227_not ; n50228
g49973 and b[36] n49740_not ; n50229
g49974 and n49734_not n50229 ; n50230
g49975 and n49742_not n50230_not ; n50231
g49976 and n50228_not n50231 ; n50232
g49977 and n49742_not n50232_not ; n50233
g49978 and b[37] n49731_not ; n50234
g49979 and n49725_not n50234 ; n50235
g49980 and n49733_not n50235_not ; n50236
g49981 and n50233_not n50236 ; n50237
g49982 and n49733_not n50237_not ; n50238
g49983 and b[38] n49722_not ; n50239
g49984 and n49716_not n50239 ; n50240
g49985 and n49724_not n50240_not ; n50241
g49986 and n50238_not n50241 ; n50242
g49987 and n49724_not n50242_not ; n50243
g49988 and b[39] n49713_not ; n50244
g49989 and n49707_not n50244 ; n50245
g49990 and n49715_not n50245_not ; n50246
g49991 and n50243_not n50246 ; n50247
g49992 and n49715_not n50247_not ; n50248
g49993 and b[40] n49704_not ; n50249
g49994 and n49698_not n50249 ; n50250
g49995 and n49706_not n50250_not ; n50251
g49996 and n50248_not n50251 ; n50252
g49997 and n49706_not n50252_not ; n50253
g49998 and b[41] n49695_not ; n50254
g49999 and n49689_not n50254 ; n50255
g50000 and n49697_not n50255_not ; n50256
g50001 and n50253_not n50256 ; n50257
g50002 and n49697_not n50257_not ; n50258
g50003 and b[42] n49686_not ; n50259
g50004 and n49680_not n50259 ; n50260
g50005 and n49688_not n50260_not ; n50261
g50006 and n50258_not n50261 ; n50262
g50007 and n49688_not n50262_not ; n50263
g50008 and b[43] n49677_not ; n50264
g50009 and n49671_not n50264 ; n50265
g50010 and n49679_not n50265_not ; n50266
g50011 and n50263_not n50266 ; n50267
g50012 and n49679_not n50267_not ; n50268
g50013 and b[44] n49668_not ; n50269
g50014 and n49662_not n50269 ; n50270
g50015 and n49670_not n50270_not ; n50271
g50016 and n50268_not n50271 ; n50272
g50017 and n49670_not n50272_not ; n50273
g50018 and b[45] n49659_not ; n50274
g50019 and n49653_not n50274 ; n50275
g50020 and n49661_not n50275_not ; n50276
g50021 and n50273_not n50276 ; n50277
g50022 and n49661_not n50277_not ; n50278
g50023 and b[46] n49650_not ; n50279
g50024 and n49644_not n50279 ; n50280
g50025 and n49652_not n50280_not ; n50281
g50026 and n50278_not n50281 ; n50282
g50027 and n49652_not n50282_not ; n50283
g50028 and b[47] n49641_not ; n50284
g50029 and n49635_not n50284 ; n50285
g50030 and n49643_not n50285_not ; n50286
g50031 and n50283_not n50286 ; n50287
g50032 and n49643_not n50287_not ; n50288
g50033 and b[48] n49632_not ; n50289
g50034 and n49626_not n50289 ; n50290
g50035 and n49634_not n50290_not ; n50291
g50036 and n50288_not n50291 ; n50292
g50037 and n49634_not n50292_not ; n50293
g50038 and b[49] n49623_not ; n50294
g50039 and n49617_not n50294 ; n50295
g50040 and n49625_not n50295_not ; n50296
g50041 and n50293_not n50296 ; n50297
g50042 and n49625_not n50297_not ; n50298
g50043 and b[50] n49614_not ; n50299
g50044 and n49608_not n50299 ; n50300
g50045 and n49616_not n50300_not ; n50301
g50046 and n50298_not n50301 ; n50302
g50047 and n49616_not n50302_not ; n50303
g50048 and b[51] n49605_not ; n50304
g50049 and n49599_not n50304 ; n50305
g50050 and n49607_not n50305_not ; n50306
g50051 and n50303_not n50306 ; n50307
g50052 and n49607_not n50307_not ; n50308
g50053 and b[52] n49596_not ; n50309
g50054 and n49590_not n50309 ; n50310
g50055 and n49598_not n50310_not ; n50311
g50056 and n50308_not n50311 ; n50312
g50057 and n49598_not n50312_not ; n50313
g50058 and b[53] n49587_not ; n50314
g50059 and n49581_not n50314 ; n50315
g50060 and n49589_not n50315_not ; n50316
g50061 and n50313_not n50316 ; n50317
g50062 and n49589_not n50317_not ; n50318
g50063 and b[54] n49578_not ; n50319
g50064 and n49572_not n50319 ; n50320
g50065 and n49580_not n50320_not ; n50321
g50066 and n50318_not n50321 ; n50322
g50067 and n49580_not n50322_not ; n50323
g50068 and n48834_not n49571_not ; n50324
g50069 and n48836_not n49568 ; n50325
g50070 and n49564_not n50325 ; n50326
g50071 and n49565_not n49568_not ; n50327
g50072 and n50326_not n50327_not ; n50328
g50073 and n49571 n50328_not ; n50329
g50074 and n50324_not n50329_not ; n50330
g50075 and b[55]_not n50330_not ; n50331
g50076 and b[55] n50324_not ; n50332
g50077 and n50329_not n50332 ; n50333
g50078 and n337 n50333_not ; n50334
g50079 and n50331_not n50334 ; n50335
g50080 and n50323_not n50335 ; n50336
g50081 and n21537 n50330_not ; n50337
g50082 and n50336_not n50337_not ; n50338
g50083 and n49589_not n50321 ; n50339
g50084 and n50317_not n50339 ; n50340
g50085 and n50318_not n50321_not ; n50341
g50086 and n50340_not n50341_not ; n50342
g50087 and n50338_not n50342_not ; n50343
g50088 and n49579_not n50337_not ; n50344
g50089 and n50336_not n50344 ; n50345
g50090 and n50343_not n50345_not ; n50346
g50091 and b[55]_not n50346_not ; n50347
g50092 and n49598_not n50316 ; n50348
g50093 and n50312_not n50348 ; n50349
g50094 and n50313_not n50316_not ; n50350
g50095 and n50349_not n50350_not ; n50351
g50096 and n50338_not n50351_not ; n50352
g50097 and n49588_not n50337_not ; n50353
g50098 and n50336_not n50353 ; n50354
g50099 and n50352_not n50354_not ; n50355
g50100 and b[54]_not n50355_not ; n50356
g50101 and n49607_not n50311 ; n50357
g50102 and n50307_not n50357 ; n50358
g50103 and n50308_not n50311_not ; n50359
g50104 and n50358_not n50359_not ; n50360
g50105 and n50338_not n50360_not ; n50361
g50106 and n49597_not n50337_not ; n50362
g50107 and n50336_not n50362 ; n50363
g50108 and n50361_not n50363_not ; n50364
g50109 and b[53]_not n50364_not ; n50365
g50110 and n49616_not n50306 ; n50366
g50111 and n50302_not n50366 ; n50367
g50112 and n50303_not n50306_not ; n50368
g50113 and n50367_not n50368_not ; n50369
g50114 and n50338_not n50369_not ; n50370
g50115 and n49606_not n50337_not ; n50371
g50116 and n50336_not n50371 ; n50372
g50117 and n50370_not n50372_not ; n50373
g50118 and b[52]_not n50373_not ; n50374
g50119 and n49625_not n50301 ; n50375
g50120 and n50297_not n50375 ; n50376
g50121 and n50298_not n50301_not ; n50377
g50122 and n50376_not n50377_not ; n50378
g50123 and n50338_not n50378_not ; n50379
g50124 and n49615_not n50337_not ; n50380
g50125 and n50336_not n50380 ; n50381
g50126 and n50379_not n50381_not ; n50382
g50127 and b[51]_not n50382_not ; n50383
g50128 and n49634_not n50296 ; n50384
g50129 and n50292_not n50384 ; n50385
g50130 and n50293_not n50296_not ; n50386
g50131 and n50385_not n50386_not ; n50387
g50132 and n50338_not n50387_not ; n50388
g50133 and n49624_not n50337_not ; n50389
g50134 and n50336_not n50389 ; n50390
g50135 and n50388_not n50390_not ; n50391
g50136 and b[50]_not n50391_not ; n50392
g50137 and n49643_not n50291 ; n50393
g50138 and n50287_not n50393 ; n50394
g50139 and n50288_not n50291_not ; n50395
g50140 and n50394_not n50395_not ; n50396
g50141 and n50338_not n50396_not ; n50397
g50142 and n49633_not n50337_not ; n50398
g50143 and n50336_not n50398 ; n50399
g50144 and n50397_not n50399_not ; n50400
g50145 and b[49]_not n50400_not ; n50401
g50146 and n49652_not n50286 ; n50402
g50147 and n50282_not n50402 ; n50403
g50148 and n50283_not n50286_not ; n50404
g50149 and n50403_not n50404_not ; n50405
g50150 and n50338_not n50405_not ; n50406
g50151 and n49642_not n50337_not ; n50407
g50152 and n50336_not n50407 ; n50408
g50153 and n50406_not n50408_not ; n50409
g50154 and b[48]_not n50409_not ; n50410
g50155 and n49661_not n50281 ; n50411
g50156 and n50277_not n50411 ; n50412
g50157 and n50278_not n50281_not ; n50413
g50158 and n50412_not n50413_not ; n50414
g50159 and n50338_not n50414_not ; n50415
g50160 and n49651_not n50337_not ; n50416
g50161 and n50336_not n50416 ; n50417
g50162 and n50415_not n50417_not ; n50418
g50163 and b[47]_not n50418_not ; n50419
g50164 and n49670_not n50276 ; n50420
g50165 and n50272_not n50420 ; n50421
g50166 and n50273_not n50276_not ; n50422
g50167 and n50421_not n50422_not ; n50423
g50168 and n50338_not n50423_not ; n50424
g50169 and n49660_not n50337_not ; n50425
g50170 and n50336_not n50425 ; n50426
g50171 and n50424_not n50426_not ; n50427
g50172 and b[46]_not n50427_not ; n50428
g50173 and n49679_not n50271 ; n50429
g50174 and n50267_not n50429 ; n50430
g50175 and n50268_not n50271_not ; n50431
g50176 and n50430_not n50431_not ; n50432
g50177 and n50338_not n50432_not ; n50433
g50178 and n49669_not n50337_not ; n50434
g50179 and n50336_not n50434 ; n50435
g50180 and n50433_not n50435_not ; n50436
g50181 and b[45]_not n50436_not ; n50437
g50182 and n49688_not n50266 ; n50438
g50183 and n50262_not n50438 ; n50439
g50184 and n50263_not n50266_not ; n50440
g50185 and n50439_not n50440_not ; n50441
g50186 and n50338_not n50441_not ; n50442
g50187 and n49678_not n50337_not ; n50443
g50188 and n50336_not n50443 ; n50444
g50189 and n50442_not n50444_not ; n50445
g50190 and b[44]_not n50445_not ; n50446
g50191 and n49697_not n50261 ; n50447
g50192 and n50257_not n50447 ; n50448
g50193 and n50258_not n50261_not ; n50449
g50194 and n50448_not n50449_not ; n50450
g50195 and n50338_not n50450_not ; n50451
g50196 and n49687_not n50337_not ; n50452
g50197 and n50336_not n50452 ; n50453
g50198 and n50451_not n50453_not ; n50454
g50199 and b[43]_not n50454_not ; n50455
g50200 and n49706_not n50256 ; n50456
g50201 and n50252_not n50456 ; n50457
g50202 and n50253_not n50256_not ; n50458
g50203 and n50457_not n50458_not ; n50459
g50204 and n50338_not n50459_not ; n50460
g50205 and n49696_not n50337_not ; n50461
g50206 and n50336_not n50461 ; n50462
g50207 and n50460_not n50462_not ; n50463
g50208 and b[42]_not n50463_not ; n50464
g50209 and n49715_not n50251 ; n50465
g50210 and n50247_not n50465 ; n50466
g50211 and n50248_not n50251_not ; n50467
g50212 and n50466_not n50467_not ; n50468
g50213 and n50338_not n50468_not ; n50469
g50214 and n49705_not n50337_not ; n50470
g50215 and n50336_not n50470 ; n50471
g50216 and n50469_not n50471_not ; n50472
g50217 and b[41]_not n50472_not ; n50473
g50218 and n49724_not n50246 ; n50474
g50219 and n50242_not n50474 ; n50475
g50220 and n50243_not n50246_not ; n50476
g50221 and n50475_not n50476_not ; n50477
g50222 and n50338_not n50477_not ; n50478
g50223 and n49714_not n50337_not ; n50479
g50224 and n50336_not n50479 ; n50480
g50225 and n50478_not n50480_not ; n50481
g50226 and b[40]_not n50481_not ; n50482
g50227 and n49733_not n50241 ; n50483
g50228 and n50237_not n50483 ; n50484
g50229 and n50238_not n50241_not ; n50485
g50230 and n50484_not n50485_not ; n50486
g50231 and n50338_not n50486_not ; n50487
g50232 and n49723_not n50337_not ; n50488
g50233 and n50336_not n50488 ; n50489
g50234 and n50487_not n50489_not ; n50490
g50235 and b[39]_not n50490_not ; n50491
g50236 and n49742_not n50236 ; n50492
g50237 and n50232_not n50492 ; n50493
g50238 and n50233_not n50236_not ; n50494
g50239 and n50493_not n50494_not ; n50495
g50240 and n50338_not n50495_not ; n50496
g50241 and n49732_not n50337_not ; n50497
g50242 and n50336_not n50497 ; n50498
g50243 and n50496_not n50498_not ; n50499
g50244 and b[38]_not n50499_not ; n50500
g50245 and n49751_not n50231 ; n50501
g50246 and n50227_not n50501 ; n50502
g50247 and n50228_not n50231_not ; n50503
g50248 and n50502_not n50503_not ; n50504
g50249 and n50338_not n50504_not ; n50505
g50250 and n49741_not n50337_not ; n50506
g50251 and n50336_not n50506 ; n50507
g50252 and n50505_not n50507_not ; n50508
g50253 and b[37]_not n50508_not ; n50509
g50254 and n49760_not n50226 ; n50510
g50255 and n50222_not n50510 ; n50511
g50256 and n50223_not n50226_not ; n50512
g50257 and n50511_not n50512_not ; n50513
g50258 and n50338_not n50513_not ; n50514
g50259 and n49750_not n50337_not ; n50515
g50260 and n50336_not n50515 ; n50516
g50261 and n50514_not n50516_not ; n50517
g50262 and b[36]_not n50517_not ; n50518
g50263 and n49769_not n50221 ; n50519
g50264 and n50217_not n50519 ; n50520
g50265 and n50218_not n50221_not ; n50521
g50266 and n50520_not n50521_not ; n50522
g50267 and n50338_not n50522_not ; n50523
g50268 and n49759_not n50337_not ; n50524
g50269 and n50336_not n50524 ; n50525
g50270 and n50523_not n50525_not ; n50526
g50271 and b[35]_not n50526_not ; n50527
g50272 and n49778_not n50216 ; n50528
g50273 and n50212_not n50528 ; n50529
g50274 and n50213_not n50216_not ; n50530
g50275 and n50529_not n50530_not ; n50531
g50276 and n50338_not n50531_not ; n50532
g50277 and n49768_not n50337_not ; n50533
g50278 and n50336_not n50533 ; n50534
g50279 and n50532_not n50534_not ; n50535
g50280 and b[34]_not n50535_not ; n50536
g50281 and n49787_not n50211 ; n50537
g50282 and n50207_not n50537 ; n50538
g50283 and n50208_not n50211_not ; n50539
g50284 and n50538_not n50539_not ; n50540
g50285 and n50338_not n50540_not ; n50541
g50286 and n49777_not n50337_not ; n50542
g50287 and n50336_not n50542 ; n50543
g50288 and n50541_not n50543_not ; n50544
g50289 and b[33]_not n50544_not ; n50545
g50290 and n49796_not n50206 ; n50546
g50291 and n50202_not n50546 ; n50547
g50292 and n50203_not n50206_not ; n50548
g50293 and n50547_not n50548_not ; n50549
g50294 and n50338_not n50549_not ; n50550
g50295 and n49786_not n50337_not ; n50551
g50296 and n50336_not n50551 ; n50552
g50297 and n50550_not n50552_not ; n50553
g50298 and b[32]_not n50553_not ; n50554
g50299 and n49805_not n50201 ; n50555
g50300 and n50197_not n50555 ; n50556
g50301 and n50198_not n50201_not ; n50557
g50302 and n50556_not n50557_not ; n50558
g50303 and n50338_not n50558_not ; n50559
g50304 and n49795_not n50337_not ; n50560
g50305 and n50336_not n50560 ; n50561
g50306 and n50559_not n50561_not ; n50562
g50307 and b[31]_not n50562_not ; n50563
g50308 and n49814_not n50196 ; n50564
g50309 and n50192_not n50564 ; n50565
g50310 and n50193_not n50196_not ; n50566
g50311 and n50565_not n50566_not ; n50567
g50312 and n50338_not n50567_not ; n50568
g50313 and n49804_not n50337_not ; n50569
g50314 and n50336_not n50569 ; n50570
g50315 and n50568_not n50570_not ; n50571
g50316 and b[30]_not n50571_not ; n50572
g50317 and n49823_not n50191 ; n50573
g50318 and n50187_not n50573 ; n50574
g50319 and n50188_not n50191_not ; n50575
g50320 and n50574_not n50575_not ; n50576
g50321 and n50338_not n50576_not ; n50577
g50322 and n49813_not n50337_not ; n50578
g50323 and n50336_not n50578 ; n50579
g50324 and n50577_not n50579_not ; n50580
g50325 and b[29]_not n50580_not ; n50581
g50326 and n49832_not n50186 ; n50582
g50327 and n50182_not n50582 ; n50583
g50328 and n50183_not n50186_not ; n50584
g50329 and n50583_not n50584_not ; n50585
g50330 and n50338_not n50585_not ; n50586
g50331 and n49822_not n50337_not ; n50587
g50332 and n50336_not n50587 ; n50588
g50333 and n50586_not n50588_not ; n50589
g50334 and b[28]_not n50589_not ; n50590
g50335 and n49841_not n50181 ; n50591
g50336 and n50177_not n50591 ; n50592
g50337 and n50178_not n50181_not ; n50593
g50338 and n50592_not n50593_not ; n50594
g50339 and n50338_not n50594_not ; n50595
g50340 and n49831_not n50337_not ; n50596
g50341 and n50336_not n50596 ; n50597
g50342 and n50595_not n50597_not ; n50598
g50343 and b[27]_not n50598_not ; n50599
g50344 and n49850_not n50176 ; n50600
g50345 and n50172_not n50600 ; n50601
g50346 and n50173_not n50176_not ; n50602
g50347 and n50601_not n50602_not ; n50603
g50348 and n50338_not n50603_not ; n50604
g50349 and n49840_not n50337_not ; n50605
g50350 and n50336_not n50605 ; n50606
g50351 and n50604_not n50606_not ; n50607
g50352 and b[26]_not n50607_not ; n50608
g50353 and n49859_not n50171 ; n50609
g50354 and n50167_not n50609 ; n50610
g50355 and n50168_not n50171_not ; n50611
g50356 and n50610_not n50611_not ; n50612
g50357 and n50338_not n50612_not ; n50613
g50358 and n49849_not n50337_not ; n50614
g50359 and n50336_not n50614 ; n50615
g50360 and n50613_not n50615_not ; n50616
g50361 and b[25]_not n50616_not ; n50617
g50362 and n49868_not n50166 ; n50618
g50363 and n50162_not n50618 ; n50619
g50364 and n50163_not n50166_not ; n50620
g50365 and n50619_not n50620_not ; n50621
g50366 and n50338_not n50621_not ; n50622
g50367 and n49858_not n50337_not ; n50623
g50368 and n50336_not n50623 ; n50624
g50369 and n50622_not n50624_not ; n50625
g50370 and b[24]_not n50625_not ; n50626
g50371 and n49877_not n50161 ; n50627
g50372 and n50157_not n50627 ; n50628
g50373 and n50158_not n50161_not ; n50629
g50374 and n50628_not n50629_not ; n50630
g50375 and n50338_not n50630_not ; n50631
g50376 and n49867_not n50337_not ; n50632
g50377 and n50336_not n50632 ; n50633
g50378 and n50631_not n50633_not ; n50634
g50379 and b[23]_not n50634_not ; n50635
g50380 and n49886_not n50156 ; n50636
g50381 and n50152_not n50636 ; n50637
g50382 and n50153_not n50156_not ; n50638
g50383 and n50637_not n50638_not ; n50639
g50384 and n50338_not n50639_not ; n50640
g50385 and n49876_not n50337_not ; n50641
g50386 and n50336_not n50641 ; n50642
g50387 and n50640_not n50642_not ; n50643
g50388 and b[22]_not n50643_not ; n50644
g50389 and n49895_not n50151 ; n50645
g50390 and n50147_not n50645 ; n50646
g50391 and n50148_not n50151_not ; n50647
g50392 and n50646_not n50647_not ; n50648
g50393 and n50338_not n50648_not ; n50649
g50394 and n49885_not n50337_not ; n50650
g50395 and n50336_not n50650 ; n50651
g50396 and n50649_not n50651_not ; n50652
g50397 and b[21]_not n50652_not ; n50653
g50398 and n49904_not n50146 ; n50654
g50399 and n50142_not n50654 ; n50655
g50400 and n50143_not n50146_not ; n50656
g50401 and n50655_not n50656_not ; n50657
g50402 and n50338_not n50657_not ; n50658
g50403 and n49894_not n50337_not ; n50659
g50404 and n50336_not n50659 ; n50660
g50405 and n50658_not n50660_not ; n50661
g50406 and b[20]_not n50661_not ; n50662
g50407 and n49913_not n50141 ; n50663
g50408 and n50137_not n50663 ; n50664
g50409 and n50138_not n50141_not ; n50665
g50410 and n50664_not n50665_not ; n50666
g50411 and n50338_not n50666_not ; n50667
g50412 and n49903_not n50337_not ; n50668
g50413 and n50336_not n50668 ; n50669
g50414 and n50667_not n50669_not ; n50670
g50415 and b[19]_not n50670_not ; n50671
g50416 and n49922_not n50136 ; n50672
g50417 and n50132_not n50672 ; n50673
g50418 and n50133_not n50136_not ; n50674
g50419 and n50673_not n50674_not ; n50675
g50420 and n50338_not n50675_not ; n50676
g50421 and n49912_not n50337_not ; n50677
g50422 and n50336_not n50677 ; n50678
g50423 and n50676_not n50678_not ; n50679
g50424 and b[18]_not n50679_not ; n50680
g50425 and n49931_not n50131 ; n50681
g50426 and n50127_not n50681 ; n50682
g50427 and n50128_not n50131_not ; n50683
g50428 and n50682_not n50683_not ; n50684
g50429 and n50338_not n50684_not ; n50685
g50430 and n49921_not n50337_not ; n50686
g50431 and n50336_not n50686 ; n50687
g50432 and n50685_not n50687_not ; n50688
g50433 and b[17]_not n50688_not ; n50689
g50434 and n49940_not n50126 ; n50690
g50435 and n50122_not n50690 ; n50691
g50436 and n50123_not n50126_not ; n50692
g50437 and n50691_not n50692_not ; n50693
g50438 and n50338_not n50693_not ; n50694
g50439 and n49930_not n50337_not ; n50695
g50440 and n50336_not n50695 ; n50696
g50441 and n50694_not n50696_not ; n50697
g50442 and b[16]_not n50697_not ; n50698
g50443 and n49949_not n50121 ; n50699
g50444 and n50117_not n50699 ; n50700
g50445 and n50118_not n50121_not ; n50701
g50446 and n50700_not n50701_not ; n50702
g50447 and n50338_not n50702_not ; n50703
g50448 and n49939_not n50337_not ; n50704
g50449 and n50336_not n50704 ; n50705
g50450 and n50703_not n50705_not ; n50706
g50451 and b[15]_not n50706_not ; n50707
g50452 and n49958_not n50116 ; n50708
g50453 and n50112_not n50708 ; n50709
g50454 and n50113_not n50116_not ; n50710
g50455 and n50709_not n50710_not ; n50711
g50456 and n50338_not n50711_not ; n50712
g50457 and n49948_not n50337_not ; n50713
g50458 and n50336_not n50713 ; n50714
g50459 and n50712_not n50714_not ; n50715
g50460 and b[14]_not n50715_not ; n50716
g50461 and n49967_not n50111 ; n50717
g50462 and n50107_not n50717 ; n50718
g50463 and n50108_not n50111_not ; n50719
g50464 and n50718_not n50719_not ; n50720
g50465 and n50338_not n50720_not ; n50721
g50466 and n49957_not n50337_not ; n50722
g50467 and n50336_not n50722 ; n50723
g50468 and n50721_not n50723_not ; n50724
g50469 and b[13]_not n50724_not ; n50725
g50470 and n49976_not n50106 ; n50726
g50471 and n50102_not n50726 ; n50727
g50472 and n50103_not n50106_not ; n50728
g50473 and n50727_not n50728_not ; n50729
g50474 and n50338_not n50729_not ; n50730
g50475 and n49966_not n50337_not ; n50731
g50476 and n50336_not n50731 ; n50732
g50477 and n50730_not n50732_not ; n50733
g50478 and b[12]_not n50733_not ; n50734
g50479 and n49985_not n50101 ; n50735
g50480 and n50097_not n50735 ; n50736
g50481 and n50098_not n50101_not ; n50737
g50482 and n50736_not n50737_not ; n50738
g50483 and n50338_not n50738_not ; n50739
g50484 and n49975_not n50337_not ; n50740
g50485 and n50336_not n50740 ; n50741
g50486 and n50739_not n50741_not ; n50742
g50487 and b[11]_not n50742_not ; n50743
g50488 and n49994_not n50096 ; n50744
g50489 and n50092_not n50744 ; n50745
g50490 and n50093_not n50096_not ; n50746
g50491 and n50745_not n50746_not ; n50747
g50492 and n50338_not n50747_not ; n50748
g50493 and n49984_not n50337_not ; n50749
g50494 and n50336_not n50749 ; n50750
g50495 and n50748_not n50750_not ; n50751
g50496 and b[10]_not n50751_not ; n50752
g50497 and n50003_not n50091 ; n50753
g50498 and n50087_not n50753 ; n50754
g50499 and n50088_not n50091_not ; n50755
g50500 and n50754_not n50755_not ; n50756
g50501 and n50338_not n50756_not ; n50757
g50502 and n49993_not n50337_not ; n50758
g50503 and n50336_not n50758 ; n50759
g50504 and n50757_not n50759_not ; n50760
g50505 and b[9]_not n50760_not ; n50761
g50506 and n50012_not n50086 ; n50762
g50507 and n50082_not n50762 ; n50763
g50508 and n50083_not n50086_not ; n50764
g50509 and n50763_not n50764_not ; n50765
g50510 and n50338_not n50765_not ; n50766
g50511 and n50002_not n50337_not ; n50767
g50512 and n50336_not n50767 ; n50768
g50513 and n50766_not n50768_not ; n50769
g50514 and b[8]_not n50769_not ; n50770
g50515 and n50021_not n50081 ; n50771
g50516 and n50077_not n50771 ; n50772
g50517 and n50078_not n50081_not ; n50773
g50518 and n50772_not n50773_not ; n50774
g50519 and n50338_not n50774_not ; n50775
g50520 and n50011_not n50337_not ; n50776
g50521 and n50336_not n50776 ; n50777
g50522 and n50775_not n50777_not ; n50778
g50523 and b[7]_not n50778_not ; n50779
g50524 and n50030_not n50076 ; n50780
g50525 and n50072_not n50780 ; n50781
g50526 and n50073_not n50076_not ; n50782
g50527 and n50781_not n50782_not ; n50783
g50528 and n50338_not n50783_not ; n50784
g50529 and n50020_not n50337_not ; n50785
g50530 and n50336_not n50785 ; n50786
g50531 and n50784_not n50786_not ; n50787
g50532 and b[6]_not n50787_not ; n50788
g50533 and n50039_not n50071 ; n50789
g50534 and n50067_not n50789 ; n50790
g50535 and n50068_not n50071_not ; n50791
g50536 and n50790_not n50791_not ; n50792
g50537 and n50338_not n50792_not ; n50793
g50538 and n50029_not n50337_not ; n50794
g50539 and n50336_not n50794 ; n50795
g50540 and n50793_not n50795_not ; n50796
g50541 and b[5]_not n50796_not ; n50797
g50542 and n50047_not n50066 ; n50798
g50543 and n50062_not n50798 ; n50799
g50544 and n50063_not n50066_not ; n50800
g50545 and n50799_not n50800_not ; n50801
g50546 and n50338_not n50801_not ; n50802
g50547 and n50038_not n50337_not ; n50803
g50548 and n50336_not n50803 ; n50804
g50549 and n50802_not n50804_not ; n50805
g50550 and b[4]_not n50805_not ; n50806
g50551 and n50057_not n50061 ; n50807
g50552 and n50056_not n50807 ; n50808
g50553 and n50058_not n50061_not ; n50809
g50554 and n50808_not n50809_not ; n50810
g50555 and n50338_not n50810_not ; n50811
g50556 and n50046_not n50337_not ; n50812
g50557 and n50336_not n50812 ; n50813
g50558 and n50811_not n50813_not ; n50814
g50559 and b[3]_not n50814_not ; n50815
g50560 and n22029 n50054_not ; n50816
g50561 and n50052_not n50816 ; n50817
g50562 and n50056_not n50817_not ; n50818
g50563 and n50338_not n50818 ; n50819
g50564 and n50051_not n50337_not ; n50820
g50565 and n50336_not n50820 ; n50821
g50566 and n50819_not n50821_not ; n50822
g50567 and b[2]_not n50822_not ; n50823
g50568 and b[0] n50338_not ; n50824
g50569 and a[8] n50824_not ; n50825
g50570 and n22029 n50338_not ; n50826
g50571 and n50825_not n50826_not ; n50827
g50572 and b[1] n50827_not ; n50828
g50573 and b[1]_not n50826_not ; n50829
g50574 and n50825_not n50829 ; n50830
g50575 and n50828_not n50830_not ; n50831
g50576 and n22806_not n50831_not ; n50832
g50577 and b[1]_not n50827_not ; n50833
g50578 and n50832_not n50833_not ; n50834
g50579 and b[2] n50821_not ; n50835
g50580 and n50819_not n50835 ; n50836
g50581 and n50823_not n50836_not ; n50837
g50582 and n50834_not n50837 ; n50838
g50583 and n50823_not n50838_not ; n50839
g50584 and b[3] n50813_not ; n50840
g50585 and n50811_not n50840 ; n50841
g50586 and n50815_not n50841_not ; n50842
g50587 and n50839_not n50842 ; n50843
g50588 and n50815_not n50843_not ; n50844
g50589 and b[4] n50804_not ; n50845
g50590 and n50802_not n50845 ; n50846
g50591 and n50806_not n50846_not ; n50847
g50592 and n50844_not n50847 ; n50848
g50593 and n50806_not n50848_not ; n50849
g50594 and b[5] n50795_not ; n50850
g50595 and n50793_not n50850 ; n50851
g50596 and n50797_not n50851_not ; n50852
g50597 and n50849_not n50852 ; n50853
g50598 and n50797_not n50853_not ; n50854
g50599 and b[6] n50786_not ; n50855
g50600 and n50784_not n50855 ; n50856
g50601 and n50788_not n50856_not ; n50857
g50602 and n50854_not n50857 ; n50858
g50603 and n50788_not n50858_not ; n50859
g50604 and b[7] n50777_not ; n50860
g50605 and n50775_not n50860 ; n50861
g50606 and n50779_not n50861_not ; n50862
g50607 and n50859_not n50862 ; n50863
g50608 and n50779_not n50863_not ; n50864
g50609 and b[8] n50768_not ; n50865
g50610 and n50766_not n50865 ; n50866
g50611 and n50770_not n50866_not ; n50867
g50612 and n50864_not n50867 ; n50868
g50613 and n50770_not n50868_not ; n50869
g50614 and b[9] n50759_not ; n50870
g50615 and n50757_not n50870 ; n50871
g50616 and n50761_not n50871_not ; n50872
g50617 and n50869_not n50872 ; n50873
g50618 and n50761_not n50873_not ; n50874
g50619 and b[10] n50750_not ; n50875
g50620 and n50748_not n50875 ; n50876
g50621 and n50752_not n50876_not ; n50877
g50622 and n50874_not n50877 ; n50878
g50623 and n50752_not n50878_not ; n50879
g50624 and b[11] n50741_not ; n50880
g50625 and n50739_not n50880 ; n50881
g50626 and n50743_not n50881_not ; n50882
g50627 and n50879_not n50882 ; n50883
g50628 and n50743_not n50883_not ; n50884
g50629 and b[12] n50732_not ; n50885
g50630 and n50730_not n50885 ; n50886
g50631 and n50734_not n50886_not ; n50887
g50632 and n50884_not n50887 ; n50888
g50633 and n50734_not n50888_not ; n50889
g50634 and b[13] n50723_not ; n50890
g50635 and n50721_not n50890 ; n50891
g50636 and n50725_not n50891_not ; n50892
g50637 and n50889_not n50892 ; n50893
g50638 and n50725_not n50893_not ; n50894
g50639 and b[14] n50714_not ; n50895
g50640 and n50712_not n50895 ; n50896
g50641 and n50716_not n50896_not ; n50897
g50642 and n50894_not n50897 ; n50898
g50643 and n50716_not n50898_not ; n50899
g50644 and b[15] n50705_not ; n50900
g50645 and n50703_not n50900 ; n50901
g50646 and n50707_not n50901_not ; n50902
g50647 and n50899_not n50902 ; n50903
g50648 and n50707_not n50903_not ; n50904
g50649 and b[16] n50696_not ; n50905
g50650 and n50694_not n50905 ; n50906
g50651 and n50698_not n50906_not ; n50907
g50652 and n50904_not n50907 ; n50908
g50653 and n50698_not n50908_not ; n50909
g50654 and b[17] n50687_not ; n50910
g50655 and n50685_not n50910 ; n50911
g50656 and n50689_not n50911_not ; n50912
g50657 and n50909_not n50912 ; n50913
g50658 and n50689_not n50913_not ; n50914
g50659 and b[18] n50678_not ; n50915
g50660 and n50676_not n50915 ; n50916
g50661 and n50680_not n50916_not ; n50917
g50662 and n50914_not n50917 ; n50918
g50663 and n50680_not n50918_not ; n50919
g50664 and b[19] n50669_not ; n50920
g50665 and n50667_not n50920 ; n50921
g50666 and n50671_not n50921_not ; n50922
g50667 and n50919_not n50922 ; n50923
g50668 and n50671_not n50923_not ; n50924
g50669 and b[20] n50660_not ; n50925
g50670 and n50658_not n50925 ; n50926
g50671 and n50662_not n50926_not ; n50927
g50672 and n50924_not n50927 ; n50928
g50673 and n50662_not n50928_not ; n50929
g50674 and b[21] n50651_not ; n50930
g50675 and n50649_not n50930 ; n50931
g50676 and n50653_not n50931_not ; n50932
g50677 and n50929_not n50932 ; n50933
g50678 and n50653_not n50933_not ; n50934
g50679 and b[22] n50642_not ; n50935
g50680 and n50640_not n50935 ; n50936
g50681 and n50644_not n50936_not ; n50937
g50682 and n50934_not n50937 ; n50938
g50683 and n50644_not n50938_not ; n50939
g50684 and b[23] n50633_not ; n50940
g50685 and n50631_not n50940 ; n50941
g50686 and n50635_not n50941_not ; n50942
g50687 and n50939_not n50942 ; n50943
g50688 and n50635_not n50943_not ; n50944
g50689 and b[24] n50624_not ; n50945
g50690 and n50622_not n50945 ; n50946
g50691 and n50626_not n50946_not ; n50947
g50692 and n50944_not n50947 ; n50948
g50693 and n50626_not n50948_not ; n50949
g50694 and b[25] n50615_not ; n50950
g50695 and n50613_not n50950 ; n50951
g50696 and n50617_not n50951_not ; n50952
g50697 and n50949_not n50952 ; n50953
g50698 and n50617_not n50953_not ; n50954
g50699 and b[26] n50606_not ; n50955
g50700 and n50604_not n50955 ; n50956
g50701 and n50608_not n50956_not ; n50957
g50702 and n50954_not n50957 ; n50958
g50703 and n50608_not n50958_not ; n50959
g50704 and b[27] n50597_not ; n50960
g50705 and n50595_not n50960 ; n50961
g50706 and n50599_not n50961_not ; n50962
g50707 and n50959_not n50962 ; n50963
g50708 and n50599_not n50963_not ; n50964
g50709 and b[28] n50588_not ; n50965
g50710 and n50586_not n50965 ; n50966
g50711 and n50590_not n50966_not ; n50967
g50712 and n50964_not n50967 ; n50968
g50713 and n50590_not n50968_not ; n50969
g50714 and b[29] n50579_not ; n50970
g50715 and n50577_not n50970 ; n50971
g50716 and n50581_not n50971_not ; n50972
g50717 and n50969_not n50972 ; n50973
g50718 and n50581_not n50973_not ; n50974
g50719 and b[30] n50570_not ; n50975
g50720 and n50568_not n50975 ; n50976
g50721 and n50572_not n50976_not ; n50977
g50722 and n50974_not n50977 ; n50978
g50723 and n50572_not n50978_not ; n50979
g50724 and b[31] n50561_not ; n50980
g50725 and n50559_not n50980 ; n50981
g50726 and n50563_not n50981_not ; n50982
g50727 and n50979_not n50982 ; n50983
g50728 and n50563_not n50983_not ; n50984
g50729 and b[32] n50552_not ; n50985
g50730 and n50550_not n50985 ; n50986
g50731 and n50554_not n50986_not ; n50987
g50732 and n50984_not n50987 ; n50988
g50733 and n50554_not n50988_not ; n50989
g50734 and b[33] n50543_not ; n50990
g50735 and n50541_not n50990 ; n50991
g50736 and n50545_not n50991_not ; n50992
g50737 and n50989_not n50992 ; n50993
g50738 and n50545_not n50993_not ; n50994
g50739 and b[34] n50534_not ; n50995
g50740 and n50532_not n50995 ; n50996
g50741 and n50536_not n50996_not ; n50997
g50742 and n50994_not n50997 ; n50998
g50743 and n50536_not n50998_not ; n50999
g50744 and b[35] n50525_not ; n51000
g50745 and n50523_not n51000 ; n51001
g50746 and n50527_not n51001_not ; n51002
g50747 and n50999_not n51002 ; n51003
g50748 and n50527_not n51003_not ; n51004
g50749 and b[36] n50516_not ; n51005
g50750 and n50514_not n51005 ; n51006
g50751 and n50518_not n51006_not ; n51007
g50752 and n51004_not n51007 ; n51008
g50753 and n50518_not n51008_not ; n51009
g50754 and b[37] n50507_not ; n51010
g50755 and n50505_not n51010 ; n51011
g50756 and n50509_not n51011_not ; n51012
g50757 and n51009_not n51012 ; n51013
g50758 and n50509_not n51013_not ; n51014
g50759 and b[38] n50498_not ; n51015
g50760 and n50496_not n51015 ; n51016
g50761 and n50500_not n51016_not ; n51017
g50762 and n51014_not n51017 ; n51018
g50763 and n50500_not n51018_not ; n51019
g50764 and b[39] n50489_not ; n51020
g50765 and n50487_not n51020 ; n51021
g50766 and n50491_not n51021_not ; n51022
g50767 and n51019_not n51022 ; n51023
g50768 and n50491_not n51023_not ; n51024
g50769 and b[40] n50480_not ; n51025
g50770 and n50478_not n51025 ; n51026
g50771 and n50482_not n51026_not ; n51027
g50772 and n51024_not n51027 ; n51028
g50773 and n50482_not n51028_not ; n51029
g50774 and b[41] n50471_not ; n51030
g50775 and n50469_not n51030 ; n51031
g50776 and n50473_not n51031_not ; n51032
g50777 and n51029_not n51032 ; n51033
g50778 and n50473_not n51033_not ; n51034
g50779 and b[42] n50462_not ; n51035
g50780 and n50460_not n51035 ; n51036
g50781 and n50464_not n51036_not ; n51037
g50782 and n51034_not n51037 ; n51038
g50783 and n50464_not n51038_not ; n51039
g50784 and b[43] n50453_not ; n51040
g50785 and n50451_not n51040 ; n51041
g50786 and n50455_not n51041_not ; n51042
g50787 and n51039_not n51042 ; n51043
g50788 and n50455_not n51043_not ; n51044
g50789 and b[44] n50444_not ; n51045
g50790 and n50442_not n51045 ; n51046
g50791 and n50446_not n51046_not ; n51047
g50792 and n51044_not n51047 ; n51048
g50793 and n50446_not n51048_not ; n51049
g50794 and b[45] n50435_not ; n51050
g50795 and n50433_not n51050 ; n51051
g50796 and n50437_not n51051_not ; n51052
g50797 and n51049_not n51052 ; n51053
g50798 and n50437_not n51053_not ; n51054
g50799 and b[46] n50426_not ; n51055
g50800 and n50424_not n51055 ; n51056
g50801 and n50428_not n51056_not ; n51057
g50802 and n51054_not n51057 ; n51058
g50803 and n50428_not n51058_not ; n51059
g50804 and b[47] n50417_not ; n51060
g50805 and n50415_not n51060 ; n51061
g50806 and n50419_not n51061_not ; n51062
g50807 and n51059_not n51062 ; n51063
g50808 and n50419_not n51063_not ; n51064
g50809 and b[48] n50408_not ; n51065
g50810 and n50406_not n51065 ; n51066
g50811 and n50410_not n51066_not ; n51067
g50812 and n51064_not n51067 ; n51068
g50813 and n50410_not n51068_not ; n51069
g50814 and b[49] n50399_not ; n51070
g50815 and n50397_not n51070 ; n51071
g50816 and n50401_not n51071_not ; n51072
g50817 and n51069_not n51072 ; n51073
g50818 and n50401_not n51073_not ; n51074
g50819 and b[50] n50390_not ; n51075
g50820 and n50388_not n51075 ; n51076
g50821 and n50392_not n51076_not ; n51077
g50822 and n51074_not n51077 ; n51078
g50823 and n50392_not n51078_not ; n51079
g50824 and b[51] n50381_not ; n51080
g50825 and n50379_not n51080 ; n51081
g50826 and n50383_not n51081_not ; n51082
g50827 and n51079_not n51082 ; n51083
g50828 and n50383_not n51083_not ; n51084
g50829 and b[52] n50372_not ; n51085
g50830 and n50370_not n51085 ; n51086
g50831 and n50374_not n51086_not ; n51087
g50832 and n51084_not n51087 ; n51088
g50833 and n50374_not n51088_not ; n51089
g50834 and b[53] n50363_not ; n51090
g50835 and n50361_not n51090 ; n51091
g50836 and n50365_not n51091_not ; n51092
g50837 and n51089_not n51092 ; n51093
g50838 and n50365_not n51093_not ; n51094
g50839 and b[54] n50354_not ; n51095
g50840 and n50352_not n51095 ; n51096
g50841 and n50356_not n51096_not ; n51097
g50842 and n51094_not n51097 ; n51098
g50843 and n50356_not n51098_not ; n51099
g50844 and b[55] n50345_not ; n51100
g50845 and n50343_not n51100 ; n51101
g50846 and n50347_not n51101_not ; n51102
g50847 and n51099_not n51102 ; n51103
g50848 and n50347_not n51103_not ; n51104
g50849 and n49580_not n50333_not ; n51105
g50850 and n50331_not n51105 ; n51106
g50851 and n50322_not n51106 ; n51107
g50852 and n50331_not n50333_not ; n51108
g50853 and n50323_not n51108_not ; n51109
g50854 and n51107_not n51109_not ; n51110
g50855 and n50338_not n51110_not ; n51111
g50856 and n50330_not n50337_not ; n51112
g50857 and n50336_not n51112 ; n51113
g50858 and n51111_not n51113_not ; n51114
g50859 and b[56]_not n51114_not ; n51115
g50860 and b[56] n51113_not ; n51116
g50861 and n51111_not n51116 ; n51117
g50862 and n407 n51117_not ; n51118
g50863 and n51115_not n51118 ; n51119
g50864 and n51104_not n51119 ; n51120
g50865 and n337 n51114_not ; n51121
g50866 and n51120_not n51121_not ; n51122
g50867 and n50356_not n51102 ; n51123
g50868 and n51098_not n51123 ; n51124
g50869 and n51099_not n51102_not ; n51125
g50870 and n51124_not n51125_not ; n51126
g50871 and n51122_not n51126_not ; n51127
g50872 and n50346_not n51121_not ; n51128
g50873 and n51120_not n51128 ; n51129
g50874 and n51127_not n51129_not ; n51130
g50875 and n50347_not n51117_not ; n51131
g50876 and n51115_not n51131 ; n51132
g50877 and n51103_not n51132 ; n51133
g50878 and n51115_not n51117_not ; n51134
g50879 and n51104_not n51134_not ; n51135
g50880 and n51133_not n51135_not ; n51136
g50881 and n51122_not n51136_not ; n51137
g50882 and n51114_not n51121_not ; n51138
g50883 and n51120_not n51138 ; n51139
g50884 and n51137_not n51139_not ; n51140
g50885 and b[57]_not n51140_not ; n51141
g50886 and b[56]_not n51130_not ; n51142
g50887 and n50365_not n51097 ; n51143
g50888 and n51093_not n51143 ; n51144
g50889 and n51094_not n51097_not ; n51145
g50890 and n51144_not n51145_not ; n51146
g50891 and n51122_not n51146_not ; n51147
g50892 and n50355_not n51121_not ; n51148
g50893 and n51120_not n51148 ; n51149
g50894 and n51147_not n51149_not ; n51150
g50895 and b[55]_not n51150_not ; n51151
g50896 and n50374_not n51092 ; n51152
g50897 and n51088_not n51152 ; n51153
g50898 and n51089_not n51092_not ; n51154
g50899 and n51153_not n51154_not ; n51155
g50900 and n51122_not n51155_not ; n51156
g50901 and n50364_not n51121_not ; n51157
g50902 and n51120_not n51157 ; n51158
g50903 and n51156_not n51158_not ; n51159
g50904 and b[54]_not n51159_not ; n51160
g50905 and n50383_not n51087 ; n51161
g50906 and n51083_not n51161 ; n51162
g50907 and n51084_not n51087_not ; n51163
g50908 and n51162_not n51163_not ; n51164
g50909 and n51122_not n51164_not ; n51165
g50910 and n50373_not n51121_not ; n51166
g50911 and n51120_not n51166 ; n51167
g50912 and n51165_not n51167_not ; n51168
g50913 and b[53]_not n51168_not ; n51169
g50914 and n50392_not n51082 ; n51170
g50915 and n51078_not n51170 ; n51171
g50916 and n51079_not n51082_not ; n51172
g50917 and n51171_not n51172_not ; n51173
g50918 and n51122_not n51173_not ; n51174
g50919 and n50382_not n51121_not ; n51175
g50920 and n51120_not n51175 ; n51176
g50921 and n51174_not n51176_not ; n51177
g50922 and b[52]_not n51177_not ; n51178
g50923 and n50401_not n51077 ; n51179
g50924 and n51073_not n51179 ; n51180
g50925 and n51074_not n51077_not ; n51181
g50926 and n51180_not n51181_not ; n51182
g50927 and n51122_not n51182_not ; n51183
g50928 and n50391_not n51121_not ; n51184
g50929 and n51120_not n51184 ; n51185
g50930 and n51183_not n51185_not ; n51186
g50931 and b[51]_not n51186_not ; n51187
g50932 and n50410_not n51072 ; n51188
g50933 and n51068_not n51188 ; n51189
g50934 and n51069_not n51072_not ; n51190
g50935 and n51189_not n51190_not ; n51191
g50936 and n51122_not n51191_not ; n51192
g50937 and n50400_not n51121_not ; n51193
g50938 and n51120_not n51193 ; n51194
g50939 and n51192_not n51194_not ; n51195
g50940 and b[50]_not n51195_not ; n51196
g50941 and n50419_not n51067 ; n51197
g50942 and n51063_not n51197 ; n51198
g50943 and n51064_not n51067_not ; n51199
g50944 and n51198_not n51199_not ; n51200
g50945 and n51122_not n51200_not ; n51201
g50946 and n50409_not n51121_not ; n51202
g50947 and n51120_not n51202 ; n51203
g50948 and n51201_not n51203_not ; n51204
g50949 and b[49]_not n51204_not ; n51205
g50950 and n50428_not n51062 ; n51206
g50951 and n51058_not n51206 ; n51207
g50952 and n51059_not n51062_not ; n51208
g50953 and n51207_not n51208_not ; n51209
g50954 and n51122_not n51209_not ; n51210
g50955 and n50418_not n51121_not ; n51211
g50956 and n51120_not n51211 ; n51212
g50957 and n51210_not n51212_not ; n51213
g50958 and b[48]_not n51213_not ; n51214
g50959 and n50437_not n51057 ; n51215
g50960 and n51053_not n51215 ; n51216
g50961 and n51054_not n51057_not ; n51217
g50962 and n51216_not n51217_not ; n51218
g50963 and n51122_not n51218_not ; n51219
g50964 and n50427_not n51121_not ; n51220
g50965 and n51120_not n51220 ; n51221
g50966 and n51219_not n51221_not ; n51222
g50967 and b[47]_not n51222_not ; n51223
g50968 and n50446_not n51052 ; n51224
g50969 and n51048_not n51224 ; n51225
g50970 and n51049_not n51052_not ; n51226
g50971 and n51225_not n51226_not ; n51227
g50972 and n51122_not n51227_not ; n51228
g50973 and n50436_not n51121_not ; n51229
g50974 and n51120_not n51229 ; n51230
g50975 and n51228_not n51230_not ; n51231
g50976 and b[46]_not n51231_not ; n51232
g50977 and n50455_not n51047 ; n51233
g50978 and n51043_not n51233 ; n51234
g50979 and n51044_not n51047_not ; n51235
g50980 and n51234_not n51235_not ; n51236
g50981 and n51122_not n51236_not ; n51237
g50982 and n50445_not n51121_not ; n51238
g50983 and n51120_not n51238 ; n51239
g50984 and n51237_not n51239_not ; n51240
g50985 and b[45]_not n51240_not ; n51241
g50986 and n50464_not n51042 ; n51242
g50987 and n51038_not n51242 ; n51243
g50988 and n51039_not n51042_not ; n51244
g50989 and n51243_not n51244_not ; n51245
g50990 and n51122_not n51245_not ; n51246
g50991 and n50454_not n51121_not ; n51247
g50992 and n51120_not n51247 ; n51248
g50993 and n51246_not n51248_not ; n51249
g50994 and b[44]_not n51249_not ; n51250
g50995 and n50473_not n51037 ; n51251
g50996 and n51033_not n51251 ; n51252
g50997 and n51034_not n51037_not ; n51253
g50998 and n51252_not n51253_not ; n51254
g50999 and n51122_not n51254_not ; n51255
g51000 and n50463_not n51121_not ; n51256
g51001 and n51120_not n51256 ; n51257
g51002 and n51255_not n51257_not ; n51258
g51003 and b[43]_not n51258_not ; n51259
g51004 and n50482_not n51032 ; n51260
g51005 and n51028_not n51260 ; n51261
g51006 and n51029_not n51032_not ; n51262
g51007 and n51261_not n51262_not ; n51263
g51008 and n51122_not n51263_not ; n51264
g51009 and n50472_not n51121_not ; n51265
g51010 and n51120_not n51265 ; n51266
g51011 and n51264_not n51266_not ; n51267
g51012 and b[42]_not n51267_not ; n51268
g51013 and n50491_not n51027 ; n51269
g51014 and n51023_not n51269 ; n51270
g51015 and n51024_not n51027_not ; n51271
g51016 and n51270_not n51271_not ; n51272
g51017 and n51122_not n51272_not ; n51273
g51018 and n50481_not n51121_not ; n51274
g51019 and n51120_not n51274 ; n51275
g51020 and n51273_not n51275_not ; n51276
g51021 and b[41]_not n51276_not ; n51277
g51022 and n50500_not n51022 ; n51278
g51023 and n51018_not n51278 ; n51279
g51024 and n51019_not n51022_not ; n51280
g51025 and n51279_not n51280_not ; n51281
g51026 and n51122_not n51281_not ; n51282
g51027 and n50490_not n51121_not ; n51283
g51028 and n51120_not n51283 ; n51284
g51029 and n51282_not n51284_not ; n51285
g51030 and b[40]_not n51285_not ; n51286
g51031 and n50509_not n51017 ; n51287
g51032 and n51013_not n51287 ; n51288
g51033 and n51014_not n51017_not ; n51289
g51034 and n51288_not n51289_not ; n51290
g51035 and n51122_not n51290_not ; n51291
g51036 and n50499_not n51121_not ; n51292
g51037 and n51120_not n51292 ; n51293
g51038 and n51291_not n51293_not ; n51294
g51039 and b[39]_not n51294_not ; n51295
g51040 and n50518_not n51012 ; n51296
g51041 and n51008_not n51296 ; n51297
g51042 and n51009_not n51012_not ; n51298
g51043 and n51297_not n51298_not ; n51299
g51044 and n51122_not n51299_not ; n51300
g51045 and n50508_not n51121_not ; n51301
g51046 and n51120_not n51301 ; n51302
g51047 and n51300_not n51302_not ; n51303
g51048 and b[38]_not n51303_not ; n51304
g51049 and n50527_not n51007 ; n51305
g51050 and n51003_not n51305 ; n51306
g51051 and n51004_not n51007_not ; n51307
g51052 and n51306_not n51307_not ; n51308
g51053 and n51122_not n51308_not ; n51309
g51054 and n50517_not n51121_not ; n51310
g51055 and n51120_not n51310 ; n51311
g51056 and n51309_not n51311_not ; n51312
g51057 and b[37]_not n51312_not ; n51313
g51058 and n50536_not n51002 ; n51314
g51059 and n50998_not n51314 ; n51315
g51060 and n50999_not n51002_not ; n51316
g51061 and n51315_not n51316_not ; n51317
g51062 and n51122_not n51317_not ; n51318
g51063 and n50526_not n51121_not ; n51319
g51064 and n51120_not n51319 ; n51320
g51065 and n51318_not n51320_not ; n51321
g51066 and b[36]_not n51321_not ; n51322
g51067 and n50545_not n50997 ; n51323
g51068 and n50993_not n51323 ; n51324
g51069 and n50994_not n50997_not ; n51325
g51070 and n51324_not n51325_not ; n51326
g51071 and n51122_not n51326_not ; n51327
g51072 and n50535_not n51121_not ; n51328
g51073 and n51120_not n51328 ; n51329
g51074 and n51327_not n51329_not ; n51330
g51075 and b[35]_not n51330_not ; n51331
g51076 and n50554_not n50992 ; n51332
g51077 and n50988_not n51332 ; n51333
g51078 and n50989_not n50992_not ; n51334
g51079 and n51333_not n51334_not ; n51335
g51080 and n51122_not n51335_not ; n51336
g51081 and n50544_not n51121_not ; n51337
g51082 and n51120_not n51337 ; n51338
g51083 and n51336_not n51338_not ; n51339
g51084 and b[34]_not n51339_not ; n51340
g51085 and n50563_not n50987 ; n51341
g51086 and n50983_not n51341 ; n51342
g51087 and n50984_not n50987_not ; n51343
g51088 and n51342_not n51343_not ; n51344
g51089 and n51122_not n51344_not ; n51345
g51090 and n50553_not n51121_not ; n51346
g51091 and n51120_not n51346 ; n51347
g51092 and n51345_not n51347_not ; n51348
g51093 and b[33]_not n51348_not ; n51349
g51094 and n50572_not n50982 ; n51350
g51095 and n50978_not n51350 ; n51351
g51096 and n50979_not n50982_not ; n51352
g51097 and n51351_not n51352_not ; n51353
g51098 and n51122_not n51353_not ; n51354
g51099 and n50562_not n51121_not ; n51355
g51100 and n51120_not n51355 ; n51356
g51101 and n51354_not n51356_not ; n51357
g51102 and b[32]_not n51357_not ; n51358
g51103 and n50581_not n50977 ; n51359
g51104 and n50973_not n51359 ; n51360
g51105 and n50974_not n50977_not ; n51361
g51106 and n51360_not n51361_not ; n51362
g51107 and n51122_not n51362_not ; n51363
g51108 and n50571_not n51121_not ; n51364
g51109 and n51120_not n51364 ; n51365
g51110 and n51363_not n51365_not ; n51366
g51111 and b[31]_not n51366_not ; n51367
g51112 and n50590_not n50972 ; n51368
g51113 and n50968_not n51368 ; n51369
g51114 and n50969_not n50972_not ; n51370
g51115 and n51369_not n51370_not ; n51371
g51116 and n51122_not n51371_not ; n51372
g51117 and n50580_not n51121_not ; n51373
g51118 and n51120_not n51373 ; n51374
g51119 and n51372_not n51374_not ; n51375
g51120 and b[30]_not n51375_not ; n51376
g51121 and n50599_not n50967 ; n51377
g51122 and n50963_not n51377 ; n51378
g51123 and n50964_not n50967_not ; n51379
g51124 and n51378_not n51379_not ; n51380
g51125 and n51122_not n51380_not ; n51381
g51126 and n50589_not n51121_not ; n51382
g51127 and n51120_not n51382 ; n51383
g51128 and n51381_not n51383_not ; n51384
g51129 and b[29]_not n51384_not ; n51385
g51130 and n50608_not n50962 ; n51386
g51131 and n50958_not n51386 ; n51387
g51132 and n50959_not n50962_not ; n51388
g51133 and n51387_not n51388_not ; n51389
g51134 and n51122_not n51389_not ; n51390
g51135 and n50598_not n51121_not ; n51391
g51136 and n51120_not n51391 ; n51392
g51137 and n51390_not n51392_not ; n51393
g51138 and b[28]_not n51393_not ; n51394
g51139 and n50617_not n50957 ; n51395
g51140 and n50953_not n51395 ; n51396
g51141 and n50954_not n50957_not ; n51397
g51142 and n51396_not n51397_not ; n51398
g51143 and n51122_not n51398_not ; n51399
g51144 and n50607_not n51121_not ; n51400
g51145 and n51120_not n51400 ; n51401
g51146 and n51399_not n51401_not ; n51402
g51147 and b[27]_not n51402_not ; n51403
g51148 and n50626_not n50952 ; n51404
g51149 and n50948_not n51404 ; n51405
g51150 and n50949_not n50952_not ; n51406
g51151 and n51405_not n51406_not ; n51407
g51152 and n51122_not n51407_not ; n51408
g51153 and n50616_not n51121_not ; n51409
g51154 and n51120_not n51409 ; n51410
g51155 and n51408_not n51410_not ; n51411
g51156 and b[26]_not n51411_not ; n51412
g51157 and n50635_not n50947 ; n51413
g51158 and n50943_not n51413 ; n51414
g51159 and n50944_not n50947_not ; n51415
g51160 and n51414_not n51415_not ; n51416
g51161 and n51122_not n51416_not ; n51417
g51162 and n50625_not n51121_not ; n51418
g51163 and n51120_not n51418 ; n51419
g51164 and n51417_not n51419_not ; n51420
g51165 and b[25]_not n51420_not ; n51421
g51166 and n50644_not n50942 ; n51422
g51167 and n50938_not n51422 ; n51423
g51168 and n50939_not n50942_not ; n51424
g51169 and n51423_not n51424_not ; n51425
g51170 and n51122_not n51425_not ; n51426
g51171 and n50634_not n51121_not ; n51427
g51172 and n51120_not n51427 ; n51428
g51173 and n51426_not n51428_not ; n51429
g51174 and b[24]_not n51429_not ; n51430
g51175 and n50653_not n50937 ; n51431
g51176 and n50933_not n51431 ; n51432
g51177 and n50934_not n50937_not ; n51433
g51178 and n51432_not n51433_not ; n51434
g51179 and n51122_not n51434_not ; n51435
g51180 and n50643_not n51121_not ; n51436
g51181 and n51120_not n51436 ; n51437
g51182 and n51435_not n51437_not ; n51438
g51183 and b[23]_not n51438_not ; n51439
g51184 and n50662_not n50932 ; n51440
g51185 and n50928_not n51440 ; n51441
g51186 and n50929_not n50932_not ; n51442
g51187 and n51441_not n51442_not ; n51443
g51188 and n51122_not n51443_not ; n51444
g51189 and n50652_not n51121_not ; n51445
g51190 and n51120_not n51445 ; n51446
g51191 and n51444_not n51446_not ; n51447
g51192 and b[22]_not n51447_not ; n51448
g51193 and n50671_not n50927 ; n51449
g51194 and n50923_not n51449 ; n51450
g51195 and n50924_not n50927_not ; n51451
g51196 and n51450_not n51451_not ; n51452
g51197 and n51122_not n51452_not ; n51453
g51198 and n50661_not n51121_not ; n51454
g51199 and n51120_not n51454 ; n51455
g51200 and n51453_not n51455_not ; n51456
g51201 and b[21]_not n51456_not ; n51457
g51202 and n50680_not n50922 ; n51458
g51203 and n50918_not n51458 ; n51459
g51204 and n50919_not n50922_not ; n51460
g51205 and n51459_not n51460_not ; n51461
g51206 and n51122_not n51461_not ; n51462
g51207 and n50670_not n51121_not ; n51463
g51208 and n51120_not n51463 ; n51464
g51209 and n51462_not n51464_not ; n51465
g51210 and b[20]_not n51465_not ; n51466
g51211 and n50689_not n50917 ; n51467
g51212 and n50913_not n51467 ; n51468
g51213 and n50914_not n50917_not ; n51469
g51214 and n51468_not n51469_not ; n51470
g51215 and n51122_not n51470_not ; n51471
g51216 and n50679_not n51121_not ; n51472
g51217 and n51120_not n51472 ; n51473
g51218 and n51471_not n51473_not ; n51474
g51219 and b[19]_not n51474_not ; n51475
g51220 and n50698_not n50912 ; n51476
g51221 and n50908_not n51476 ; n51477
g51222 and n50909_not n50912_not ; n51478
g51223 and n51477_not n51478_not ; n51479
g51224 and n51122_not n51479_not ; n51480
g51225 and n50688_not n51121_not ; n51481
g51226 and n51120_not n51481 ; n51482
g51227 and n51480_not n51482_not ; n51483
g51228 and b[18]_not n51483_not ; n51484
g51229 and n50707_not n50907 ; n51485
g51230 and n50903_not n51485 ; n51486
g51231 and n50904_not n50907_not ; n51487
g51232 and n51486_not n51487_not ; n51488
g51233 and n51122_not n51488_not ; n51489
g51234 and n50697_not n51121_not ; n51490
g51235 and n51120_not n51490 ; n51491
g51236 and n51489_not n51491_not ; n51492
g51237 and b[17]_not n51492_not ; n51493
g51238 and n50716_not n50902 ; n51494
g51239 and n50898_not n51494 ; n51495
g51240 and n50899_not n50902_not ; n51496
g51241 and n51495_not n51496_not ; n51497
g51242 and n51122_not n51497_not ; n51498
g51243 and n50706_not n51121_not ; n51499
g51244 and n51120_not n51499 ; n51500
g51245 and n51498_not n51500_not ; n51501
g51246 and b[16]_not n51501_not ; n51502
g51247 and n50725_not n50897 ; n51503
g51248 and n50893_not n51503 ; n51504
g51249 and n50894_not n50897_not ; n51505
g51250 and n51504_not n51505_not ; n51506
g51251 and n51122_not n51506_not ; n51507
g51252 and n50715_not n51121_not ; n51508
g51253 and n51120_not n51508 ; n51509
g51254 and n51507_not n51509_not ; n51510
g51255 and b[15]_not n51510_not ; n51511
g51256 and n50734_not n50892 ; n51512
g51257 and n50888_not n51512 ; n51513
g51258 and n50889_not n50892_not ; n51514
g51259 and n51513_not n51514_not ; n51515
g51260 and n51122_not n51515_not ; n51516
g51261 and n50724_not n51121_not ; n51517
g51262 and n51120_not n51517 ; n51518
g51263 and n51516_not n51518_not ; n51519
g51264 and b[14]_not n51519_not ; n51520
g51265 and n50743_not n50887 ; n51521
g51266 and n50883_not n51521 ; n51522
g51267 and n50884_not n50887_not ; n51523
g51268 and n51522_not n51523_not ; n51524
g51269 and n51122_not n51524_not ; n51525
g51270 and n50733_not n51121_not ; n51526
g51271 and n51120_not n51526 ; n51527
g51272 and n51525_not n51527_not ; n51528
g51273 and b[13]_not n51528_not ; n51529
g51274 and n50752_not n50882 ; n51530
g51275 and n50878_not n51530 ; n51531
g51276 and n50879_not n50882_not ; n51532
g51277 and n51531_not n51532_not ; n51533
g51278 and n51122_not n51533_not ; n51534
g51279 and n50742_not n51121_not ; n51535
g51280 and n51120_not n51535 ; n51536
g51281 and n51534_not n51536_not ; n51537
g51282 and b[12]_not n51537_not ; n51538
g51283 and n50761_not n50877 ; n51539
g51284 and n50873_not n51539 ; n51540
g51285 and n50874_not n50877_not ; n51541
g51286 and n51540_not n51541_not ; n51542
g51287 and n51122_not n51542_not ; n51543
g51288 and n50751_not n51121_not ; n51544
g51289 and n51120_not n51544 ; n51545
g51290 and n51543_not n51545_not ; n51546
g51291 and b[11]_not n51546_not ; n51547
g51292 and n50770_not n50872 ; n51548
g51293 and n50868_not n51548 ; n51549
g51294 and n50869_not n50872_not ; n51550
g51295 and n51549_not n51550_not ; n51551
g51296 and n51122_not n51551_not ; n51552
g51297 and n50760_not n51121_not ; n51553
g51298 and n51120_not n51553 ; n51554
g51299 and n51552_not n51554_not ; n51555
g51300 and b[10]_not n51555_not ; n51556
g51301 and n50779_not n50867 ; n51557
g51302 and n50863_not n51557 ; n51558
g51303 and n50864_not n50867_not ; n51559
g51304 and n51558_not n51559_not ; n51560
g51305 and n51122_not n51560_not ; n51561
g51306 and n50769_not n51121_not ; n51562
g51307 and n51120_not n51562 ; n51563
g51308 and n51561_not n51563_not ; n51564
g51309 and b[9]_not n51564_not ; n51565
g51310 and n50788_not n50862 ; n51566
g51311 and n50858_not n51566 ; n51567
g51312 and n50859_not n50862_not ; n51568
g51313 and n51567_not n51568_not ; n51569
g51314 and n51122_not n51569_not ; n51570
g51315 and n50778_not n51121_not ; n51571
g51316 and n51120_not n51571 ; n51572
g51317 and n51570_not n51572_not ; n51573
g51318 and b[8]_not n51573_not ; n51574
g51319 and n50797_not n50857 ; n51575
g51320 and n50853_not n51575 ; n51576
g51321 and n50854_not n50857_not ; n51577
g51322 and n51576_not n51577_not ; n51578
g51323 and n51122_not n51578_not ; n51579
g51324 and n50787_not n51121_not ; n51580
g51325 and n51120_not n51580 ; n51581
g51326 and n51579_not n51581_not ; n51582
g51327 and b[7]_not n51582_not ; n51583
g51328 and n50806_not n50852 ; n51584
g51329 and n50848_not n51584 ; n51585
g51330 and n50849_not n50852_not ; n51586
g51331 and n51585_not n51586_not ; n51587
g51332 and n51122_not n51587_not ; n51588
g51333 and n50796_not n51121_not ; n51589
g51334 and n51120_not n51589 ; n51590
g51335 and n51588_not n51590_not ; n51591
g51336 and b[6]_not n51591_not ; n51592
g51337 and n50815_not n50847 ; n51593
g51338 and n50843_not n51593 ; n51594
g51339 and n50844_not n50847_not ; n51595
g51340 and n51594_not n51595_not ; n51596
g51341 and n51122_not n51596_not ; n51597
g51342 and n50805_not n51121_not ; n51598
g51343 and n51120_not n51598 ; n51599
g51344 and n51597_not n51599_not ; n51600
g51345 and b[5]_not n51600_not ; n51601
g51346 and n50823_not n50842 ; n51602
g51347 and n50838_not n51602 ; n51603
g51348 and n50839_not n50842_not ; n51604
g51349 and n51603_not n51604_not ; n51605
g51350 and n51122_not n51605_not ; n51606
g51351 and n50814_not n51121_not ; n51607
g51352 and n51120_not n51607 ; n51608
g51353 and n51606_not n51608_not ; n51609
g51354 and b[4]_not n51609_not ; n51610
g51355 and n50833_not n50837 ; n51611
g51356 and n50832_not n51611 ; n51612
g51357 and n50834_not n50837_not ; n51613
g51358 and n51612_not n51613_not ; n51614
g51359 and n51122_not n51614_not ; n51615
g51360 and n50822_not n51121_not ; n51616
g51361 and n51120_not n51616 ; n51617
g51362 and n51615_not n51617_not ; n51618
g51363 and b[3]_not n51618_not ; n51619
g51364 and n22806 n50830_not ; n51620
g51365 and n50828_not n51620 ; n51621
g51366 and n50832_not n51621_not ; n51622
g51367 and n51122_not n51622 ; n51623
g51368 and n50827_not n51121_not ; n51624
g51369 and n51120_not n51624 ; n51625
g51370 and n51623_not n51625_not ; n51626
g51371 and b[2]_not n51626_not ; n51627
g51372 and b[0] n51122_not ; n51628
g51373 and a[7] n51628_not ; n51629
g51374 and n22806 n51122_not ; n51630
g51375 and n51629_not n51630_not ; n51631
g51376 and b[1] n51631_not ; n51632
g51377 and b[1]_not n51630_not ; n51633
g51378 and n51629_not n51633 ; n51634
g51379 and n51632_not n51634_not ; n51635
g51380 and n23611_not n51635_not ; n51636
g51381 and b[1]_not n51631_not ; n51637
g51382 and n51636_not n51637_not ; n51638
g51383 and b[2] n51625_not ; n51639
g51384 and n51623_not n51639 ; n51640
g51385 and n51627_not n51640_not ; n51641
g51386 and n51638_not n51641 ; n51642
g51387 and n51627_not n51642_not ; n51643
g51388 and b[3] n51617_not ; n51644
g51389 and n51615_not n51644 ; n51645
g51390 and n51619_not n51645_not ; n51646
g51391 and n51643_not n51646 ; n51647
g51392 and n51619_not n51647_not ; n51648
g51393 and b[4] n51608_not ; n51649
g51394 and n51606_not n51649 ; n51650
g51395 and n51610_not n51650_not ; n51651
g51396 and n51648_not n51651 ; n51652
g51397 and n51610_not n51652_not ; n51653
g51398 and b[5] n51599_not ; n51654
g51399 and n51597_not n51654 ; n51655
g51400 and n51601_not n51655_not ; n51656
g51401 and n51653_not n51656 ; n51657
g51402 and n51601_not n51657_not ; n51658
g51403 and b[6] n51590_not ; n51659
g51404 and n51588_not n51659 ; n51660
g51405 and n51592_not n51660_not ; n51661
g51406 and n51658_not n51661 ; n51662
g51407 and n51592_not n51662_not ; n51663
g51408 and b[7] n51581_not ; n51664
g51409 and n51579_not n51664 ; n51665
g51410 and n51583_not n51665_not ; n51666
g51411 and n51663_not n51666 ; n51667
g51412 and n51583_not n51667_not ; n51668
g51413 and b[8] n51572_not ; n51669
g51414 and n51570_not n51669 ; n51670
g51415 and n51574_not n51670_not ; n51671
g51416 and n51668_not n51671 ; n51672
g51417 and n51574_not n51672_not ; n51673
g51418 and b[9] n51563_not ; n51674
g51419 and n51561_not n51674 ; n51675
g51420 and n51565_not n51675_not ; n51676
g51421 and n51673_not n51676 ; n51677
g51422 and n51565_not n51677_not ; n51678
g51423 and b[10] n51554_not ; n51679
g51424 and n51552_not n51679 ; n51680
g51425 and n51556_not n51680_not ; n51681
g51426 and n51678_not n51681 ; n51682
g51427 and n51556_not n51682_not ; n51683
g51428 and b[11] n51545_not ; n51684
g51429 and n51543_not n51684 ; n51685
g51430 and n51547_not n51685_not ; n51686
g51431 and n51683_not n51686 ; n51687
g51432 and n51547_not n51687_not ; n51688
g51433 and b[12] n51536_not ; n51689
g51434 and n51534_not n51689 ; n51690
g51435 and n51538_not n51690_not ; n51691
g51436 and n51688_not n51691 ; n51692
g51437 and n51538_not n51692_not ; n51693
g51438 and b[13] n51527_not ; n51694
g51439 and n51525_not n51694 ; n51695
g51440 and n51529_not n51695_not ; n51696
g51441 and n51693_not n51696 ; n51697
g51442 and n51529_not n51697_not ; n51698
g51443 and b[14] n51518_not ; n51699
g51444 and n51516_not n51699 ; n51700
g51445 and n51520_not n51700_not ; n51701
g51446 and n51698_not n51701 ; n51702
g51447 and n51520_not n51702_not ; n51703
g51448 and b[15] n51509_not ; n51704
g51449 and n51507_not n51704 ; n51705
g51450 and n51511_not n51705_not ; n51706
g51451 and n51703_not n51706 ; n51707
g51452 and n51511_not n51707_not ; n51708
g51453 and b[16] n51500_not ; n51709
g51454 and n51498_not n51709 ; n51710
g51455 and n51502_not n51710_not ; n51711
g51456 and n51708_not n51711 ; n51712
g51457 and n51502_not n51712_not ; n51713
g51458 and b[17] n51491_not ; n51714
g51459 and n51489_not n51714 ; n51715
g51460 and n51493_not n51715_not ; n51716
g51461 and n51713_not n51716 ; n51717
g51462 and n51493_not n51717_not ; n51718
g51463 and b[18] n51482_not ; n51719
g51464 and n51480_not n51719 ; n51720
g51465 and n51484_not n51720_not ; n51721
g51466 and n51718_not n51721 ; n51722
g51467 and n51484_not n51722_not ; n51723
g51468 and b[19] n51473_not ; n51724
g51469 and n51471_not n51724 ; n51725
g51470 and n51475_not n51725_not ; n51726
g51471 and n51723_not n51726 ; n51727
g51472 and n51475_not n51727_not ; n51728
g51473 and b[20] n51464_not ; n51729
g51474 and n51462_not n51729 ; n51730
g51475 and n51466_not n51730_not ; n51731
g51476 and n51728_not n51731 ; n51732
g51477 and n51466_not n51732_not ; n51733
g51478 and b[21] n51455_not ; n51734
g51479 and n51453_not n51734 ; n51735
g51480 and n51457_not n51735_not ; n51736
g51481 and n51733_not n51736 ; n51737
g51482 and n51457_not n51737_not ; n51738
g51483 and b[22] n51446_not ; n51739
g51484 and n51444_not n51739 ; n51740
g51485 and n51448_not n51740_not ; n51741
g51486 and n51738_not n51741 ; n51742
g51487 and n51448_not n51742_not ; n51743
g51488 and b[23] n51437_not ; n51744
g51489 and n51435_not n51744 ; n51745
g51490 and n51439_not n51745_not ; n51746
g51491 and n51743_not n51746 ; n51747
g51492 and n51439_not n51747_not ; n51748
g51493 and b[24] n51428_not ; n51749
g51494 and n51426_not n51749 ; n51750
g51495 and n51430_not n51750_not ; n51751
g51496 and n51748_not n51751 ; n51752
g51497 and n51430_not n51752_not ; n51753
g51498 and b[25] n51419_not ; n51754
g51499 and n51417_not n51754 ; n51755
g51500 and n51421_not n51755_not ; n51756
g51501 and n51753_not n51756 ; n51757
g51502 and n51421_not n51757_not ; n51758
g51503 and b[26] n51410_not ; n51759
g51504 and n51408_not n51759 ; n51760
g51505 and n51412_not n51760_not ; n51761
g51506 and n51758_not n51761 ; n51762
g51507 and n51412_not n51762_not ; n51763
g51508 and b[27] n51401_not ; n51764
g51509 and n51399_not n51764 ; n51765
g51510 and n51403_not n51765_not ; n51766
g51511 and n51763_not n51766 ; n51767
g51512 and n51403_not n51767_not ; n51768
g51513 and b[28] n51392_not ; n51769
g51514 and n51390_not n51769 ; n51770
g51515 and n51394_not n51770_not ; n51771
g51516 and n51768_not n51771 ; n51772
g51517 and n51394_not n51772_not ; n51773
g51518 and b[29] n51383_not ; n51774
g51519 and n51381_not n51774 ; n51775
g51520 and n51385_not n51775_not ; n51776
g51521 and n51773_not n51776 ; n51777
g51522 and n51385_not n51777_not ; n51778
g51523 and b[30] n51374_not ; n51779
g51524 and n51372_not n51779 ; n51780
g51525 and n51376_not n51780_not ; n51781
g51526 and n51778_not n51781 ; n51782
g51527 and n51376_not n51782_not ; n51783
g51528 and b[31] n51365_not ; n51784
g51529 and n51363_not n51784 ; n51785
g51530 and n51367_not n51785_not ; n51786
g51531 and n51783_not n51786 ; n51787
g51532 and n51367_not n51787_not ; n51788
g51533 and b[32] n51356_not ; n51789
g51534 and n51354_not n51789 ; n51790
g51535 and n51358_not n51790_not ; n51791
g51536 and n51788_not n51791 ; n51792
g51537 and n51358_not n51792_not ; n51793
g51538 and b[33] n51347_not ; n51794
g51539 and n51345_not n51794 ; n51795
g51540 and n51349_not n51795_not ; n51796
g51541 and n51793_not n51796 ; n51797
g51542 and n51349_not n51797_not ; n51798
g51543 and b[34] n51338_not ; n51799
g51544 and n51336_not n51799 ; n51800
g51545 and n51340_not n51800_not ; n51801
g51546 and n51798_not n51801 ; n51802
g51547 and n51340_not n51802_not ; n51803
g51548 and b[35] n51329_not ; n51804
g51549 and n51327_not n51804 ; n51805
g51550 and n51331_not n51805_not ; n51806
g51551 and n51803_not n51806 ; n51807
g51552 and n51331_not n51807_not ; n51808
g51553 and b[36] n51320_not ; n51809
g51554 and n51318_not n51809 ; n51810
g51555 and n51322_not n51810_not ; n51811
g51556 and n51808_not n51811 ; n51812
g51557 and n51322_not n51812_not ; n51813
g51558 and b[37] n51311_not ; n51814
g51559 and n51309_not n51814 ; n51815
g51560 and n51313_not n51815_not ; n51816
g51561 and n51813_not n51816 ; n51817
g51562 and n51313_not n51817_not ; n51818
g51563 and b[38] n51302_not ; n51819
g51564 and n51300_not n51819 ; n51820
g51565 and n51304_not n51820_not ; n51821
g51566 and n51818_not n51821 ; n51822
g51567 and n51304_not n51822_not ; n51823
g51568 and b[39] n51293_not ; n51824
g51569 and n51291_not n51824 ; n51825
g51570 and n51295_not n51825_not ; n51826
g51571 and n51823_not n51826 ; n51827
g51572 and n51295_not n51827_not ; n51828
g51573 and b[40] n51284_not ; n51829
g51574 and n51282_not n51829 ; n51830
g51575 and n51286_not n51830_not ; n51831
g51576 and n51828_not n51831 ; n51832
g51577 and n51286_not n51832_not ; n51833
g51578 and b[41] n51275_not ; n51834
g51579 and n51273_not n51834 ; n51835
g51580 and n51277_not n51835_not ; n51836
g51581 and n51833_not n51836 ; n51837
g51582 and n51277_not n51837_not ; n51838
g51583 and b[42] n51266_not ; n51839
g51584 and n51264_not n51839 ; n51840
g51585 and n51268_not n51840_not ; n51841
g51586 and n51838_not n51841 ; n51842
g51587 and n51268_not n51842_not ; n51843
g51588 and b[43] n51257_not ; n51844
g51589 and n51255_not n51844 ; n51845
g51590 and n51259_not n51845_not ; n51846
g51591 and n51843_not n51846 ; n51847
g51592 and n51259_not n51847_not ; n51848
g51593 and b[44] n51248_not ; n51849
g51594 and n51246_not n51849 ; n51850
g51595 and n51250_not n51850_not ; n51851
g51596 and n51848_not n51851 ; n51852
g51597 and n51250_not n51852_not ; n51853
g51598 and b[45] n51239_not ; n51854
g51599 and n51237_not n51854 ; n51855
g51600 and n51241_not n51855_not ; n51856
g51601 and n51853_not n51856 ; n51857
g51602 and n51241_not n51857_not ; n51858
g51603 and b[46] n51230_not ; n51859
g51604 and n51228_not n51859 ; n51860
g51605 and n51232_not n51860_not ; n51861
g51606 and n51858_not n51861 ; n51862
g51607 and n51232_not n51862_not ; n51863
g51608 and b[47] n51221_not ; n51864
g51609 and n51219_not n51864 ; n51865
g51610 and n51223_not n51865_not ; n51866
g51611 and n51863_not n51866 ; n51867
g51612 and n51223_not n51867_not ; n51868
g51613 and b[48] n51212_not ; n51869
g51614 and n51210_not n51869 ; n51870
g51615 and n51214_not n51870_not ; n51871
g51616 and n51868_not n51871 ; n51872
g51617 and n51214_not n51872_not ; n51873
g51618 and b[49] n51203_not ; n51874
g51619 and n51201_not n51874 ; n51875
g51620 and n51205_not n51875_not ; n51876
g51621 and n51873_not n51876 ; n51877
g51622 and n51205_not n51877_not ; n51878
g51623 and b[50] n51194_not ; n51879
g51624 and n51192_not n51879 ; n51880
g51625 and n51196_not n51880_not ; n51881
g51626 and n51878_not n51881 ; n51882
g51627 and n51196_not n51882_not ; n51883
g51628 and b[51] n51185_not ; n51884
g51629 and n51183_not n51884 ; n51885
g51630 and n51187_not n51885_not ; n51886
g51631 and n51883_not n51886 ; n51887
g51632 and n51187_not n51887_not ; n51888
g51633 and b[52] n51176_not ; n51889
g51634 and n51174_not n51889 ; n51890
g51635 and n51178_not n51890_not ; n51891
g51636 and n51888_not n51891 ; n51892
g51637 and n51178_not n51892_not ; n51893
g51638 and b[53] n51167_not ; n51894
g51639 and n51165_not n51894 ; n51895
g51640 and n51169_not n51895_not ; n51896
g51641 and n51893_not n51896 ; n51897
g51642 and n51169_not n51897_not ; n51898
g51643 and b[54] n51158_not ; n51899
g51644 and n51156_not n51899 ; n51900
g51645 and n51160_not n51900_not ; n51901
g51646 and n51898_not n51901 ; n51902
g51647 and n51160_not n51902_not ; n51903
g51648 and b[55] n51149_not ; n51904
g51649 and n51147_not n51904 ; n51905
g51650 and n51151_not n51905_not ; n51906
g51651 and n51903_not n51906 ; n51907
g51652 and n51151_not n51907_not ; n51908
g51653 and b[56] n51129_not ; n51909
g51654 and n51127_not n51909 ; n51910
g51655 and n51142_not n51910_not ; n51911
g51656 and n51908_not n51911 ; n51912
g51657 and n51142_not n51912_not ; n51913
g51658 and b[57] n51139_not ; n51914
g51659 and n51137_not n51914 ; n51915
g51660 and n51141_not n51915_not ; n51916
g51661 and n51913_not n51916 ; n51917
g51662 and n51141_not n51917_not ; n51918
g51663 and n23895 n51918_not ; n51919
g51664 and n51130_not n51919_not ; n51920
g51665 and n51151_not n51911 ; n51921
g51666 and n51907_not n51921 ; n51922
g51667 and n51908_not n51911_not ; n51923
g51668 and n51922_not n51923_not ; n51924
g51669 and n23895 n51924_not ; n51925
g51670 and n51918_not n51925 ; n51926
g51671 and n51920_not n51926_not ; n51927
g51672 and b[57]_not n51927_not ; n51928
g51673 and n51150_not n51919_not ; n51929
g51674 and n51160_not n51906 ; n51930
g51675 and n51902_not n51930 ; n51931
g51676 and n51903_not n51906_not ; n51932
g51677 and n51931_not n51932_not ; n51933
g51678 and n23895 n51933_not ; n51934
g51679 and n51918_not n51934 ; n51935
g51680 and n51929_not n51935_not ; n51936
g51681 and b[56]_not n51936_not ; n51937
g51682 and n51159_not n51919_not ; n51938
g51683 and n51169_not n51901 ; n51939
g51684 and n51897_not n51939 ; n51940
g51685 and n51898_not n51901_not ; n51941
g51686 and n51940_not n51941_not ; n51942
g51687 and n23895 n51942_not ; n51943
g51688 and n51918_not n51943 ; n51944
g51689 and n51938_not n51944_not ; n51945
g51690 and b[55]_not n51945_not ; n51946
g51691 and n51168_not n51919_not ; n51947
g51692 and n51178_not n51896 ; n51948
g51693 and n51892_not n51948 ; n51949
g51694 and n51893_not n51896_not ; n51950
g51695 and n51949_not n51950_not ; n51951
g51696 and n23895 n51951_not ; n51952
g51697 and n51918_not n51952 ; n51953
g51698 and n51947_not n51953_not ; n51954
g51699 and b[54]_not n51954_not ; n51955
g51700 and n51177_not n51919_not ; n51956
g51701 and n51187_not n51891 ; n51957
g51702 and n51887_not n51957 ; n51958
g51703 and n51888_not n51891_not ; n51959
g51704 and n51958_not n51959_not ; n51960
g51705 and n23895 n51960_not ; n51961
g51706 and n51918_not n51961 ; n51962
g51707 and n51956_not n51962_not ; n51963
g51708 and b[53]_not n51963_not ; n51964
g51709 and n51186_not n51919_not ; n51965
g51710 and n51196_not n51886 ; n51966
g51711 and n51882_not n51966 ; n51967
g51712 and n51883_not n51886_not ; n51968
g51713 and n51967_not n51968_not ; n51969
g51714 and n23895 n51969_not ; n51970
g51715 and n51918_not n51970 ; n51971
g51716 and n51965_not n51971_not ; n51972
g51717 and b[52]_not n51972_not ; n51973
g51718 and n51195_not n51919_not ; n51974
g51719 and n51205_not n51881 ; n51975
g51720 and n51877_not n51975 ; n51976
g51721 and n51878_not n51881_not ; n51977
g51722 and n51976_not n51977_not ; n51978
g51723 and n23895 n51978_not ; n51979
g51724 and n51918_not n51979 ; n51980
g51725 and n51974_not n51980_not ; n51981
g51726 and b[51]_not n51981_not ; n51982
g51727 and n51204_not n51919_not ; n51983
g51728 and n51214_not n51876 ; n51984
g51729 and n51872_not n51984 ; n51985
g51730 and n51873_not n51876_not ; n51986
g51731 and n51985_not n51986_not ; n51987
g51732 and n23895 n51987_not ; n51988
g51733 and n51918_not n51988 ; n51989
g51734 and n51983_not n51989_not ; n51990
g51735 and b[50]_not n51990_not ; n51991
g51736 and n51213_not n51919_not ; n51992
g51737 and n51223_not n51871 ; n51993
g51738 and n51867_not n51993 ; n51994
g51739 and n51868_not n51871_not ; n51995
g51740 and n51994_not n51995_not ; n51996
g51741 and n23895 n51996_not ; n51997
g51742 and n51918_not n51997 ; n51998
g51743 and n51992_not n51998_not ; n51999
g51744 and b[49]_not n51999_not ; n52000
g51745 and n51222_not n51919_not ; n52001
g51746 and n51232_not n51866 ; n52002
g51747 and n51862_not n52002 ; n52003
g51748 and n51863_not n51866_not ; n52004
g51749 and n52003_not n52004_not ; n52005
g51750 and n23895 n52005_not ; n52006
g51751 and n51918_not n52006 ; n52007
g51752 and n52001_not n52007_not ; n52008
g51753 and b[48]_not n52008_not ; n52009
g51754 and n51231_not n51919_not ; n52010
g51755 and n51241_not n51861 ; n52011
g51756 and n51857_not n52011 ; n52012
g51757 and n51858_not n51861_not ; n52013
g51758 and n52012_not n52013_not ; n52014
g51759 and n23895 n52014_not ; n52015
g51760 and n51918_not n52015 ; n52016
g51761 and n52010_not n52016_not ; n52017
g51762 and b[47]_not n52017_not ; n52018
g51763 and n51240_not n51919_not ; n52019
g51764 and n51250_not n51856 ; n52020
g51765 and n51852_not n52020 ; n52021
g51766 and n51853_not n51856_not ; n52022
g51767 and n52021_not n52022_not ; n52023
g51768 and n23895 n52023_not ; n52024
g51769 and n51918_not n52024 ; n52025
g51770 and n52019_not n52025_not ; n52026
g51771 and b[46]_not n52026_not ; n52027
g51772 and n51249_not n51919_not ; n52028
g51773 and n51259_not n51851 ; n52029
g51774 and n51847_not n52029 ; n52030
g51775 and n51848_not n51851_not ; n52031
g51776 and n52030_not n52031_not ; n52032
g51777 and n23895 n52032_not ; n52033
g51778 and n51918_not n52033 ; n52034
g51779 and n52028_not n52034_not ; n52035
g51780 and b[45]_not n52035_not ; n52036
g51781 and n51258_not n51919_not ; n52037
g51782 and n51268_not n51846 ; n52038
g51783 and n51842_not n52038 ; n52039
g51784 and n51843_not n51846_not ; n52040
g51785 and n52039_not n52040_not ; n52041
g51786 and n23895 n52041_not ; n52042
g51787 and n51918_not n52042 ; n52043
g51788 and n52037_not n52043_not ; n52044
g51789 and b[44]_not n52044_not ; n52045
g51790 and n51267_not n51919_not ; n52046
g51791 and n51277_not n51841 ; n52047
g51792 and n51837_not n52047 ; n52048
g51793 and n51838_not n51841_not ; n52049
g51794 and n52048_not n52049_not ; n52050
g51795 and n23895 n52050_not ; n52051
g51796 and n51918_not n52051 ; n52052
g51797 and n52046_not n52052_not ; n52053
g51798 and b[43]_not n52053_not ; n52054
g51799 and n51276_not n51919_not ; n52055
g51800 and n51286_not n51836 ; n52056
g51801 and n51832_not n52056 ; n52057
g51802 and n51833_not n51836_not ; n52058
g51803 and n52057_not n52058_not ; n52059
g51804 and n23895 n52059_not ; n52060
g51805 and n51918_not n52060 ; n52061
g51806 and n52055_not n52061_not ; n52062
g51807 and b[42]_not n52062_not ; n52063
g51808 and n51285_not n51919_not ; n52064
g51809 and n51295_not n51831 ; n52065
g51810 and n51827_not n52065 ; n52066
g51811 and n51828_not n51831_not ; n52067
g51812 and n52066_not n52067_not ; n52068
g51813 and n23895 n52068_not ; n52069
g51814 and n51918_not n52069 ; n52070
g51815 and n52064_not n52070_not ; n52071
g51816 and b[41]_not n52071_not ; n52072
g51817 and n51294_not n51919_not ; n52073
g51818 and n51304_not n51826 ; n52074
g51819 and n51822_not n52074 ; n52075
g51820 and n51823_not n51826_not ; n52076
g51821 and n52075_not n52076_not ; n52077
g51822 and n23895 n52077_not ; n52078
g51823 and n51918_not n52078 ; n52079
g51824 and n52073_not n52079_not ; n52080
g51825 and b[40]_not n52080_not ; n52081
g51826 and n51303_not n51919_not ; n52082
g51827 and n51313_not n51821 ; n52083
g51828 and n51817_not n52083 ; n52084
g51829 and n51818_not n51821_not ; n52085
g51830 and n52084_not n52085_not ; n52086
g51831 and n23895 n52086_not ; n52087
g51832 and n51918_not n52087 ; n52088
g51833 and n52082_not n52088_not ; n52089
g51834 and b[39]_not n52089_not ; n52090
g51835 and n51312_not n51919_not ; n52091
g51836 and n51322_not n51816 ; n52092
g51837 and n51812_not n52092 ; n52093
g51838 and n51813_not n51816_not ; n52094
g51839 and n52093_not n52094_not ; n52095
g51840 and n23895 n52095_not ; n52096
g51841 and n51918_not n52096 ; n52097
g51842 and n52091_not n52097_not ; n52098
g51843 and b[38]_not n52098_not ; n52099
g51844 and n51321_not n51919_not ; n52100
g51845 and n51331_not n51811 ; n52101
g51846 and n51807_not n52101 ; n52102
g51847 and n51808_not n51811_not ; n52103
g51848 and n52102_not n52103_not ; n52104
g51849 and n23895 n52104_not ; n52105
g51850 and n51918_not n52105 ; n52106
g51851 and n52100_not n52106_not ; n52107
g51852 and b[37]_not n52107_not ; n52108
g51853 and n51330_not n51919_not ; n52109
g51854 and n51340_not n51806 ; n52110
g51855 and n51802_not n52110 ; n52111
g51856 and n51803_not n51806_not ; n52112
g51857 and n52111_not n52112_not ; n52113
g51858 and n23895 n52113_not ; n52114
g51859 and n51918_not n52114 ; n52115
g51860 and n52109_not n52115_not ; n52116
g51861 and b[36]_not n52116_not ; n52117
g51862 and n51339_not n51919_not ; n52118
g51863 and n51349_not n51801 ; n52119
g51864 and n51797_not n52119 ; n52120
g51865 and n51798_not n51801_not ; n52121
g51866 and n52120_not n52121_not ; n52122
g51867 and n23895 n52122_not ; n52123
g51868 and n51918_not n52123 ; n52124
g51869 and n52118_not n52124_not ; n52125
g51870 and b[35]_not n52125_not ; n52126
g51871 and n51348_not n51919_not ; n52127
g51872 and n51358_not n51796 ; n52128
g51873 and n51792_not n52128 ; n52129
g51874 and n51793_not n51796_not ; n52130
g51875 and n52129_not n52130_not ; n52131
g51876 and n23895 n52131_not ; n52132
g51877 and n51918_not n52132 ; n52133
g51878 and n52127_not n52133_not ; n52134
g51879 and b[34]_not n52134_not ; n52135
g51880 and n51357_not n51919_not ; n52136
g51881 and n51367_not n51791 ; n52137
g51882 and n51787_not n52137 ; n52138
g51883 and n51788_not n51791_not ; n52139
g51884 and n52138_not n52139_not ; n52140
g51885 and n23895 n52140_not ; n52141
g51886 and n51918_not n52141 ; n52142
g51887 and n52136_not n52142_not ; n52143
g51888 and b[33]_not n52143_not ; n52144
g51889 and n51366_not n51919_not ; n52145
g51890 and n51376_not n51786 ; n52146
g51891 and n51782_not n52146 ; n52147
g51892 and n51783_not n51786_not ; n52148
g51893 and n52147_not n52148_not ; n52149
g51894 and n23895 n52149_not ; n52150
g51895 and n51918_not n52150 ; n52151
g51896 and n52145_not n52151_not ; n52152
g51897 and b[32]_not n52152_not ; n52153
g51898 and n51375_not n51919_not ; n52154
g51899 and n51385_not n51781 ; n52155
g51900 and n51777_not n52155 ; n52156
g51901 and n51778_not n51781_not ; n52157
g51902 and n52156_not n52157_not ; n52158
g51903 and n23895 n52158_not ; n52159
g51904 and n51918_not n52159 ; n52160
g51905 and n52154_not n52160_not ; n52161
g51906 and b[31]_not n52161_not ; n52162
g51907 and n51384_not n51919_not ; n52163
g51908 and n51394_not n51776 ; n52164
g51909 and n51772_not n52164 ; n52165
g51910 and n51773_not n51776_not ; n52166
g51911 and n52165_not n52166_not ; n52167
g51912 and n23895 n52167_not ; n52168
g51913 and n51918_not n52168 ; n52169
g51914 and n52163_not n52169_not ; n52170
g51915 and b[30]_not n52170_not ; n52171
g51916 and n51393_not n51919_not ; n52172
g51917 and n51403_not n51771 ; n52173
g51918 and n51767_not n52173 ; n52174
g51919 and n51768_not n51771_not ; n52175
g51920 and n52174_not n52175_not ; n52176
g51921 and n23895 n52176_not ; n52177
g51922 and n51918_not n52177 ; n52178
g51923 and n52172_not n52178_not ; n52179
g51924 and b[29]_not n52179_not ; n52180
g51925 and n51402_not n51919_not ; n52181
g51926 and n51412_not n51766 ; n52182
g51927 and n51762_not n52182 ; n52183
g51928 and n51763_not n51766_not ; n52184
g51929 and n52183_not n52184_not ; n52185
g51930 and n23895 n52185_not ; n52186
g51931 and n51918_not n52186 ; n52187
g51932 and n52181_not n52187_not ; n52188
g51933 and b[28]_not n52188_not ; n52189
g51934 and n51411_not n51919_not ; n52190
g51935 and n51421_not n51761 ; n52191
g51936 and n51757_not n52191 ; n52192
g51937 and n51758_not n51761_not ; n52193
g51938 and n52192_not n52193_not ; n52194
g51939 and n23895 n52194_not ; n52195
g51940 and n51918_not n52195 ; n52196
g51941 and n52190_not n52196_not ; n52197
g51942 and b[27]_not n52197_not ; n52198
g51943 and n51420_not n51919_not ; n52199
g51944 and n51430_not n51756 ; n52200
g51945 and n51752_not n52200 ; n52201
g51946 and n51753_not n51756_not ; n52202
g51947 and n52201_not n52202_not ; n52203
g51948 and n23895 n52203_not ; n52204
g51949 and n51918_not n52204 ; n52205
g51950 and n52199_not n52205_not ; n52206
g51951 and b[26]_not n52206_not ; n52207
g51952 and n51429_not n51919_not ; n52208
g51953 and n51439_not n51751 ; n52209
g51954 and n51747_not n52209 ; n52210
g51955 and n51748_not n51751_not ; n52211
g51956 and n52210_not n52211_not ; n52212
g51957 and n23895 n52212_not ; n52213
g51958 and n51918_not n52213 ; n52214
g51959 and n52208_not n52214_not ; n52215
g51960 and b[25]_not n52215_not ; n52216
g51961 and n51438_not n51919_not ; n52217
g51962 and n51448_not n51746 ; n52218
g51963 and n51742_not n52218 ; n52219
g51964 and n51743_not n51746_not ; n52220
g51965 and n52219_not n52220_not ; n52221
g51966 and n23895 n52221_not ; n52222
g51967 and n51918_not n52222 ; n52223
g51968 and n52217_not n52223_not ; n52224
g51969 and b[24]_not n52224_not ; n52225
g51970 and n51447_not n51919_not ; n52226
g51971 and n51457_not n51741 ; n52227
g51972 and n51737_not n52227 ; n52228
g51973 and n51738_not n51741_not ; n52229
g51974 and n52228_not n52229_not ; n52230
g51975 and n23895 n52230_not ; n52231
g51976 and n51918_not n52231 ; n52232
g51977 and n52226_not n52232_not ; n52233
g51978 and b[23]_not n52233_not ; n52234
g51979 and n51456_not n51919_not ; n52235
g51980 and n51466_not n51736 ; n52236
g51981 and n51732_not n52236 ; n52237
g51982 and n51733_not n51736_not ; n52238
g51983 and n52237_not n52238_not ; n52239
g51984 and n23895 n52239_not ; n52240
g51985 and n51918_not n52240 ; n52241
g51986 and n52235_not n52241_not ; n52242
g51987 and b[22]_not n52242_not ; n52243
g51988 and n51465_not n51919_not ; n52244
g51989 and n51475_not n51731 ; n52245
g51990 and n51727_not n52245 ; n52246
g51991 and n51728_not n51731_not ; n52247
g51992 and n52246_not n52247_not ; n52248
g51993 and n23895 n52248_not ; n52249
g51994 and n51918_not n52249 ; n52250
g51995 and n52244_not n52250_not ; n52251
g51996 and b[21]_not n52251_not ; n52252
g51997 and n51474_not n51919_not ; n52253
g51998 and n51484_not n51726 ; n52254
g51999 and n51722_not n52254 ; n52255
g52000 and n51723_not n51726_not ; n52256
g52001 and n52255_not n52256_not ; n52257
g52002 and n23895 n52257_not ; n52258
g52003 and n51918_not n52258 ; n52259
g52004 and n52253_not n52259_not ; n52260
g52005 and b[20]_not n52260_not ; n52261
g52006 and n51483_not n51919_not ; n52262
g52007 and n51493_not n51721 ; n52263
g52008 and n51717_not n52263 ; n52264
g52009 and n51718_not n51721_not ; n52265
g52010 and n52264_not n52265_not ; n52266
g52011 and n23895 n52266_not ; n52267
g52012 and n51918_not n52267 ; n52268
g52013 and n52262_not n52268_not ; n52269
g52014 and b[19]_not n52269_not ; n52270
g52015 and n51492_not n51919_not ; n52271
g52016 and n51502_not n51716 ; n52272
g52017 and n51712_not n52272 ; n52273
g52018 and n51713_not n51716_not ; n52274
g52019 and n52273_not n52274_not ; n52275
g52020 and n23895 n52275_not ; n52276
g52021 and n51918_not n52276 ; n52277
g52022 and n52271_not n52277_not ; n52278
g52023 and b[18]_not n52278_not ; n52279
g52024 and n51501_not n51919_not ; n52280
g52025 and n51511_not n51711 ; n52281
g52026 and n51707_not n52281 ; n52282
g52027 and n51708_not n51711_not ; n52283
g52028 and n52282_not n52283_not ; n52284
g52029 and n23895 n52284_not ; n52285
g52030 and n51918_not n52285 ; n52286
g52031 and n52280_not n52286_not ; n52287
g52032 and b[17]_not n52287_not ; n52288
g52033 and n51510_not n51919_not ; n52289
g52034 and n51520_not n51706 ; n52290
g52035 and n51702_not n52290 ; n52291
g52036 and n51703_not n51706_not ; n52292
g52037 and n52291_not n52292_not ; n52293
g52038 and n23895 n52293_not ; n52294
g52039 and n51918_not n52294 ; n52295
g52040 and n52289_not n52295_not ; n52296
g52041 and b[16]_not n52296_not ; n52297
g52042 and n51519_not n51919_not ; n52298
g52043 and n51529_not n51701 ; n52299
g52044 and n51697_not n52299 ; n52300
g52045 and n51698_not n51701_not ; n52301
g52046 and n52300_not n52301_not ; n52302
g52047 and n23895 n52302_not ; n52303
g52048 and n51918_not n52303 ; n52304
g52049 and n52298_not n52304_not ; n52305
g52050 and b[15]_not n52305_not ; n52306
g52051 and n51528_not n51919_not ; n52307
g52052 and n51538_not n51696 ; n52308
g52053 and n51692_not n52308 ; n52309
g52054 and n51693_not n51696_not ; n52310
g52055 and n52309_not n52310_not ; n52311
g52056 and n23895 n52311_not ; n52312
g52057 and n51918_not n52312 ; n52313
g52058 and n52307_not n52313_not ; n52314
g52059 and b[14]_not n52314_not ; n52315
g52060 and n51537_not n51919_not ; n52316
g52061 and n51547_not n51691 ; n52317
g52062 and n51687_not n52317 ; n52318
g52063 and n51688_not n51691_not ; n52319
g52064 and n52318_not n52319_not ; n52320
g52065 and n23895 n52320_not ; n52321
g52066 and n51918_not n52321 ; n52322
g52067 and n52316_not n52322_not ; n52323
g52068 and b[13]_not n52323_not ; n52324
g52069 and n51546_not n51919_not ; n52325
g52070 and n51556_not n51686 ; n52326
g52071 and n51682_not n52326 ; n52327
g52072 and n51683_not n51686_not ; n52328
g52073 and n52327_not n52328_not ; n52329
g52074 and n23895 n52329_not ; n52330
g52075 and n51918_not n52330 ; n52331
g52076 and n52325_not n52331_not ; n52332
g52077 and b[12]_not n52332_not ; n52333
g52078 and n51555_not n51919_not ; n52334
g52079 and n51565_not n51681 ; n52335
g52080 and n51677_not n52335 ; n52336
g52081 and n51678_not n51681_not ; n52337
g52082 and n52336_not n52337_not ; n52338
g52083 and n23895 n52338_not ; n52339
g52084 and n51918_not n52339 ; n52340
g52085 and n52334_not n52340_not ; n52341
g52086 and b[11]_not n52341_not ; n52342
g52087 and n51564_not n51919_not ; n52343
g52088 and n51574_not n51676 ; n52344
g52089 and n51672_not n52344 ; n52345
g52090 and n51673_not n51676_not ; n52346
g52091 and n52345_not n52346_not ; n52347
g52092 and n23895 n52347_not ; n52348
g52093 and n51918_not n52348 ; n52349
g52094 and n52343_not n52349_not ; n52350
g52095 and b[10]_not n52350_not ; n52351
g52096 and n51573_not n51919_not ; n52352
g52097 and n51583_not n51671 ; n52353
g52098 and n51667_not n52353 ; n52354
g52099 and n51668_not n51671_not ; n52355
g52100 and n52354_not n52355_not ; n52356
g52101 and n23895 n52356_not ; n52357
g52102 and n51918_not n52357 ; n52358
g52103 and n52352_not n52358_not ; n52359
g52104 and b[9]_not n52359_not ; n52360
g52105 and n51582_not n51919_not ; n52361
g52106 and n51592_not n51666 ; n52362
g52107 and n51662_not n52362 ; n52363
g52108 and n51663_not n51666_not ; n52364
g52109 and n52363_not n52364_not ; n52365
g52110 and n23895 n52365_not ; n52366
g52111 and n51918_not n52366 ; n52367
g52112 and n52361_not n52367_not ; n52368
g52113 and b[8]_not n52368_not ; n52369
g52114 and n51591_not n51919_not ; n52370
g52115 and n51601_not n51661 ; n52371
g52116 and n51657_not n52371 ; n52372
g52117 and n51658_not n51661_not ; n52373
g52118 and n52372_not n52373_not ; n52374
g52119 and n23895 n52374_not ; n52375
g52120 and n51918_not n52375 ; n52376
g52121 and n52370_not n52376_not ; n52377
g52122 and b[7]_not n52377_not ; n52378
g52123 and n51600_not n51919_not ; n52379
g52124 and n51610_not n51656 ; n52380
g52125 and n51652_not n52380 ; n52381
g52126 and n51653_not n51656_not ; n52382
g52127 and n52381_not n52382_not ; n52383
g52128 and n23895 n52383_not ; n52384
g52129 and n51918_not n52384 ; n52385
g52130 and n52379_not n52385_not ; n52386
g52131 and b[6]_not n52386_not ; n52387
g52132 and n51609_not n51919_not ; n52388
g52133 and n51619_not n51651 ; n52389
g52134 and n51647_not n52389 ; n52390
g52135 and n51648_not n51651_not ; n52391
g52136 and n52390_not n52391_not ; n52392
g52137 and n23895 n52392_not ; n52393
g52138 and n51918_not n52393 ; n52394
g52139 and n52388_not n52394_not ; n52395
g52140 and b[5]_not n52395_not ; n52396
g52141 and n51618_not n51919_not ; n52397
g52142 and n51627_not n51646 ; n52398
g52143 and n51642_not n52398 ; n52399
g52144 and n51643_not n51646_not ; n52400
g52145 and n52399_not n52400_not ; n52401
g52146 and n23895 n52401_not ; n52402
g52147 and n51918_not n52402 ; n52403
g52148 and n52397_not n52403_not ; n52404
g52149 and b[4]_not n52404_not ; n52405
g52150 and n51626_not n51919_not ; n52406
g52151 and n51637_not n51641 ; n52407
g52152 and n51636_not n52407 ; n52408
g52153 and n51638_not n51641_not ; n52409
g52154 and n52408_not n52409_not ; n52410
g52155 and n23895 n52410_not ; n52411
g52156 and n51918_not n52411 ; n52412
g52157 and n52406_not n52412_not ; n52413
g52158 and b[3]_not n52413_not ; n52414
g52159 and n51631_not n51919_not ; n52415
g52160 and n23611 n51634_not ; n52416
g52161 and n51632_not n52416 ; n52417
g52162 and n23895 n52417_not ; n52418
g52163 and n51636_not n52418 ; n52419
g52164 and n51918_not n52419 ; n52420
g52165 and n52415_not n52420_not ; n52421
g52166 and b[2]_not n52421_not ; n52422
g52167 and n24402 n51918_not ; n52423
g52168 and a[6] n52423_not ; n52424
g52169 and n24406 n51918_not ; n52425
g52170 and n52424_not n52425_not ; n52426
g52171 and b[1] n52426_not ; n52427
g52172 and b[1]_not n52425_not ; n52428
g52173 and n52424_not n52428 ; n52429
g52174 and n52427_not n52429_not ; n52430
g52175 and n24413_not n52430_not ; n52431
g52176 and b[1]_not n52426_not ; n52432
g52177 and n52431_not n52432_not ; n52433
g52178 and b[2] n52420_not ; n52434
g52179 and n52415_not n52434 ; n52435
g52180 and n52422_not n52435_not ; n52436
g52181 and n52433_not n52436 ; n52437
g52182 and n52422_not n52437_not ; n52438
g52183 and b[3] n52412_not ; n52439
g52184 and n52406_not n52439 ; n52440
g52185 and n52414_not n52440_not ; n52441
g52186 and n52438_not n52441 ; n52442
g52187 and n52414_not n52442_not ; n52443
g52188 and b[4] n52403_not ; n52444
g52189 and n52397_not n52444 ; n52445
g52190 and n52405_not n52445_not ; n52446
g52191 and n52443_not n52446 ; n52447
g52192 and n52405_not n52447_not ; n52448
g52193 and b[5] n52394_not ; n52449
g52194 and n52388_not n52449 ; n52450
g52195 and n52396_not n52450_not ; n52451
g52196 and n52448_not n52451 ; n52452
g52197 and n52396_not n52452_not ; n52453
g52198 and b[6] n52385_not ; n52454
g52199 and n52379_not n52454 ; n52455
g52200 and n52387_not n52455_not ; n52456
g52201 and n52453_not n52456 ; n52457
g52202 and n52387_not n52457_not ; n52458
g52203 and b[7] n52376_not ; n52459
g52204 and n52370_not n52459 ; n52460
g52205 and n52378_not n52460_not ; n52461
g52206 and n52458_not n52461 ; n52462
g52207 and n52378_not n52462_not ; n52463
g52208 and b[8] n52367_not ; n52464
g52209 and n52361_not n52464 ; n52465
g52210 and n52369_not n52465_not ; n52466
g52211 and n52463_not n52466 ; n52467
g52212 and n52369_not n52467_not ; n52468
g52213 and b[9] n52358_not ; n52469
g52214 and n52352_not n52469 ; n52470
g52215 and n52360_not n52470_not ; n52471
g52216 and n52468_not n52471 ; n52472
g52217 and n52360_not n52472_not ; n52473
g52218 and b[10] n52349_not ; n52474
g52219 and n52343_not n52474 ; n52475
g52220 and n52351_not n52475_not ; n52476
g52221 and n52473_not n52476 ; n52477
g52222 and n52351_not n52477_not ; n52478
g52223 and b[11] n52340_not ; n52479
g52224 and n52334_not n52479 ; n52480
g52225 and n52342_not n52480_not ; n52481
g52226 and n52478_not n52481 ; n52482
g52227 and n52342_not n52482_not ; n52483
g52228 and b[12] n52331_not ; n52484
g52229 and n52325_not n52484 ; n52485
g52230 and n52333_not n52485_not ; n52486
g52231 and n52483_not n52486 ; n52487
g52232 and n52333_not n52487_not ; n52488
g52233 and b[13] n52322_not ; n52489
g52234 and n52316_not n52489 ; n52490
g52235 and n52324_not n52490_not ; n52491
g52236 and n52488_not n52491 ; n52492
g52237 and n52324_not n52492_not ; n52493
g52238 and b[14] n52313_not ; n52494
g52239 and n52307_not n52494 ; n52495
g52240 and n52315_not n52495_not ; n52496
g52241 and n52493_not n52496 ; n52497
g52242 and n52315_not n52497_not ; n52498
g52243 and b[15] n52304_not ; n52499
g52244 and n52298_not n52499 ; n52500
g52245 and n52306_not n52500_not ; n52501
g52246 and n52498_not n52501 ; n52502
g52247 and n52306_not n52502_not ; n52503
g52248 and b[16] n52295_not ; n52504
g52249 and n52289_not n52504 ; n52505
g52250 and n52297_not n52505_not ; n52506
g52251 and n52503_not n52506 ; n52507
g52252 and n52297_not n52507_not ; n52508
g52253 and b[17] n52286_not ; n52509
g52254 and n52280_not n52509 ; n52510
g52255 and n52288_not n52510_not ; n52511
g52256 and n52508_not n52511 ; n52512
g52257 and n52288_not n52512_not ; n52513
g52258 and b[18] n52277_not ; n52514
g52259 and n52271_not n52514 ; n52515
g52260 and n52279_not n52515_not ; n52516
g52261 and n52513_not n52516 ; n52517
g52262 and n52279_not n52517_not ; n52518
g52263 and b[19] n52268_not ; n52519
g52264 and n52262_not n52519 ; n52520
g52265 and n52270_not n52520_not ; n52521
g52266 and n52518_not n52521 ; n52522
g52267 and n52270_not n52522_not ; n52523
g52268 and b[20] n52259_not ; n52524
g52269 and n52253_not n52524 ; n52525
g52270 and n52261_not n52525_not ; n52526
g52271 and n52523_not n52526 ; n52527
g52272 and n52261_not n52527_not ; n52528
g52273 and b[21] n52250_not ; n52529
g52274 and n52244_not n52529 ; n52530
g52275 and n52252_not n52530_not ; n52531
g52276 and n52528_not n52531 ; n52532
g52277 and n52252_not n52532_not ; n52533
g52278 and b[22] n52241_not ; n52534
g52279 and n52235_not n52534 ; n52535
g52280 and n52243_not n52535_not ; n52536
g52281 and n52533_not n52536 ; n52537
g52282 and n52243_not n52537_not ; n52538
g52283 and b[23] n52232_not ; n52539
g52284 and n52226_not n52539 ; n52540
g52285 and n52234_not n52540_not ; n52541
g52286 and n52538_not n52541 ; n52542
g52287 and n52234_not n52542_not ; n52543
g52288 and b[24] n52223_not ; n52544
g52289 and n52217_not n52544 ; n52545
g52290 and n52225_not n52545_not ; n52546
g52291 and n52543_not n52546 ; n52547
g52292 and n52225_not n52547_not ; n52548
g52293 and b[25] n52214_not ; n52549
g52294 and n52208_not n52549 ; n52550
g52295 and n52216_not n52550_not ; n52551
g52296 and n52548_not n52551 ; n52552
g52297 and n52216_not n52552_not ; n52553
g52298 and b[26] n52205_not ; n52554
g52299 and n52199_not n52554 ; n52555
g52300 and n52207_not n52555_not ; n52556
g52301 and n52553_not n52556 ; n52557
g52302 and n52207_not n52557_not ; n52558
g52303 and b[27] n52196_not ; n52559
g52304 and n52190_not n52559 ; n52560
g52305 and n52198_not n52560_not ; n52561
g52306 and n52558_not n52561 ; n52562
g52307 and n52198_not n52562_not ; n52563
g52308 and b[28] n52187_not ; n52564
g52309 and n52181_not n52564 ; n52565
g52310 and n52189_not n52565_not ; n52566
g52311 and n52563_not n52566 ; n52567
g52312 and n52189_not n52567_not ; n52568
g52313 and b[29] n52178_not ; n52569
g52314 and n52172_not n52569 ; n52570
g52315 and n52180_not n52570_not ; n52571
g52316 and n52568_not n52571 ; n52572
g52317 and n52180_not n52572_not ; n52573
g52318 and b[30] n52169_not ; n52574
g52319 and n52163_not n52574 ; n52575
g52320 and n52171_not n52575_not ; n52576
g52321 and n52573_not n52576 ; n52577
g52322 and n52171_not n52577_not ; n52578
g52323 and b[31] n52160_not ; n52579
g52324 and n52154_not n52579 ; n52580
g52325 and n52162_not n52580_not ; n52581
g52326 and n52578_not n52581 ; n52582
g52327 and n52162_not n52582_not ; n52583
g52328 and b[32] n52151_not ; n52584
g52329 and n52145_not n52584 ; n52585
g52330 and n52153_not n52585_not ; n52586
g52331 and n52583_not n52586 ; n52587
g52332 and n52153_not n52587_not ; n52588
g52333 and b[33] n52142_not ; n52589
g52334 and n52136_not n52589 ; n52590
g52335 and n52144_not n52590_not ; n52591
g52336 and n52588_not n52591 ; n52592
g52337 and n52144_not n52592_not ; n52593
g52338 and b[34] n52133_not ; n52594
g52339 and n52127_not n52594 ; n52595
g52340 and n52135_not n52595_not ; n52596
g52341 and n52593_not n52596 ; n52597
g52342 and n52135_not n52597_not ; n52598
g52343 and b[35] n52124_not ; n52599
g52344 and n52118_not n52599 ; n52600
g52345 and n52126_not n52600_not ; n52601
g52346 and n52598_not n52601 ; n52602
g52347 and n52126_not n52602_not ; n52603
g52348 and b[36] n52115_not ; n52604
g52349 and n52109_not n52604 ; n52605
g52350 and n52117_not n52605_not ; n52606
g52351 and n52603_not n52606 ; n52607
g52352 and n52117_not n52607_not ; n52608
g52353 and b[37] n52106_not ; n52609
g52354 and n52100_not n52609 ; n52610
g52355 and n52108_not n52610_not ; n52611
g52356 and n52608_not n52611 ; n52612
g52357 and n52108_not n52612_not ; n52613
g52358 and b[38] n52097_not ; n52614
g52359 and n52091_not n52614 ; n52615
g52360 and n52099_not n52615_not ; n52616
g52361 and n52613_not n52616 ; n52617
g52362 and n52099_not n52617_not ; n52618
g52363 and b[39] n52088_not ; n52619
g52364 and n52082_not n52619 ; n52620
g52365 and n52090_not n52620_not ; n52621
g52366 and n52618_not n52621 ; n52622
g52367 and n52090_not n52622_not ; n52623
g52368 and b[40] n52079_not ; n52624
g52369 and n52073_not n52624 ; n52625
g52370 and n52081_not n52625_not ; n52626
g52371 and n52623_not n52626 ; n52627
g52372 and n52081_not n52627_not ; n52628
g52373 and b[41] n52070_not ; n52629
g52374 and n52064_not n52629 ; n52630
g52375 and n52072_not n52630_not ; n52631
g52376 and n52628_not n52631 ; n52632
g52377 and n52072_not n52632_not ; n52633
g52378 and b[42] n52061_not ; n52634
g52379 and n52055_not n52634 ; n52635
g52380 and n52063_not n52635_not ; n52636
g52381 and n52633_not n52636 ; n52637
g52382 and n52063_not n52637_not ; n52638
g52383 and b[43] n52052_not ; n52639
g52384 and n52046_not n52639 ; n52640
g52385 and n52054_not n52640_not ; n52641
g52386 and n52638_not n52641 ; n52642
g52387 and n52054_not n52642_not ; n52643
g52388 and b[44] n52043_not ; n52644
g52389 and n52037_not n52644 ; n52645
g52390 and n52045_not n52645_not ; n52646
g52391 and n52643_not n52646 ; n52647
g52392 and n52045_not n52647_not ; n52648
g52393 and b[45] n52034_not ; n52649
g52394 and n52028_not n52649 ; n52650
g52395 and n52036_not n52650_not ; n52651
g52396 and n52648_not n52651 ; n52652
g52397 and n52036_not n52652_not ; n52653
g52398 and b[46] n52025_not ; n52654
g52399 and n52019_not n52654 ; n52655
g52400 and n52027_not n52655_not ; n52656
g52401 and n52653_not n52656 ; n52657
g52402 and n52027_not n52657_not ; n52658
g52403 and b[47] n52016_not ; n52659
g52404 and n52010_not n52659 ; n52660
g52405 and n52018_not n52660_not ; n52661
g52406 and n52658_not n52661 ; n52662
g52407 and n52018_not n52662_not ; n52663
g52408 and b[48] n52007_not ; n52664
g52409 and n52001_not n52664 ; n52665
g52410 and n52009_not n52665_not ; n52666
g52411 and n52663_not n52666 ; n52667
g52412 and n52009_not n52667_not ; n52668
g52413 and b[49] n51998_not ; n52669
g52414 and n51992_not n52669 ; n52670
g52415 and n52000_not n52670_not ; n52671
g52416 and n52668_not n52671 ; n52672
g52417 and n52000_not n52672_not ; n52673
g52418 and b[50] n51989_not ; n52674
g52419 and n51983_not n52674 ; n52675
g52420 and n51991_not n52675_not ; n52676
g52421 and n52673_not n52676 ; n52677
g52422 and n51991_not n52677_not ; n52678
g52423 and b[51] n51980_not ; n52679
g52424 and n51974_not n52679 ; n52680
g52425 and n51982_not n52680_not ; n52681
g52426 and n52678_not n52681 ; n52682
g52427 and n51982_not n52682_not ; n52683
g52428 and b[52] n51971_not ; n52684
g52429 and n51965_not n52684 ; n52685
g52430 and n51973_not n52685_not ; n52686
g52431 and n52683_not n52686 ; n52687
g52432 and n51973_not n52687_not ; n52688
g52433 and b[53] n51962_not ; n52689
g52434 and n51956_not n52689 ; n52690
g52435 and n51964_not n52690_not ; n52691
g52436 and n52688_not n52691 ; n52692
g52437 and n51964_not n52692_not ; n52693
g52438 and b[54] n51953_not ; n52694
g52439 and n51947_not n52694 ; n52695
g52440 and n51955_not n52695_not ; n52696
g52441 and n52693_not n52696 ; n52697
g52442 and n51955_not n52697_not ; n52698
g52443 and b[55] n51944_not ; n52699
g52444 and n51938_not n52699 ; n52700
g52445 and n51946_not n52700_not ; n52701
g52446 and n52698_not n52701 ; n52702
g52447 and n51946_not n52702_not ; n52703
g52448 and b[56] n51935_not ; n52704
g52449 and n51929_not n52704 ; n52705
g52450 and n51937_not n52705_not ; n52706
g52451 and n52703_not n52706 ; n52707
g52452 and n51937_not n52707_not ; n52708
g52453 and b[57] n51926_not ; n52709
g52454 and n51920_not n52709 ; n52710
g52455 and n51928_not n52710_not ; n52711
g52456 and n52708_not n52711 ; n52712
g52457 and n51928_not n52712_not ; n52713
g52458 and n51140_not n51919_not ; n52714
g52459 and n51142_not n51916 ; n52715
g52460 and n51912_not n52715 ; n52716
g52461 and n51913_not n51916_not ; n52717
g52462 and n52716_not n52717_not ; n52718
g52463 and n51919 n52718_not ; n52719
g52464 and n52714_not n52719_not ; n52720
g52465 and b[58]_not n52720_not ; n52721
g52466 and b[58] n52714_not ; n52722
g52467 and n52719_not n52722 ; n52723
g52468 and n24707 n52723_not ; n52724
g52469 and n52721_not n52724 ; n52725
g52470 and n52713_not n52725 ; n52726
g52471 and n23895 n52720_not ; n52727
g52472 and n52726_not n52727_not ; n52728
g52473 and n51937_not n52711 ; n52729
g52474 and n52707_not n52729 ; n52730
g52475 and n52708_not n52711_not ; n52731
g52476 and n52730_not n52731_not ; n52732
g52477 and n52728_not n52732_not ; n52733
g52478 and n51927_not n52727_not ; n52734
g52479 and n52726_not n52734 ; n52735
g52480 and n52733_not n52735_not ; n52736
g52481 and b[58]_not n52736_not ; n52737
g52482 and n51946_not n52706 ; n52738
g52483 and n52702_not n52738 ; n52739
g52484 and n52703_not n52706_not ; n52740
g52485 and n52739_not n52740_not ; n52741
g52486 and n52728_not n52741_not ; n52742
g52487 and n51936_not n52727_not ; n52743
g52488 and n52726_not n52743 ; n52744
g52489 and n52742_not n52744_not ; n52745
g52490 and b[57]_not n52745_not ; n52746
g52491 and n51955_not n52701 ; n52747
g52492 and n52697_not n52747 ; n52748
g52493 and n52698_not n52701_not ; n52749
g52494 and n52748_not n52749_not ; n52750
g52495 and n52728_not n52750_not ; n52751
g52496 and n51945_not n52727_not ; n52752
g52497 and n52726_not n52752 ; n52753
g52498 and n52751_not n52753_not ; n52754
g52499 and b[56]_not n52754_not ; n52755
g52500 and n51964_not n52696 ; n52756
g52501 and n52692_not n52756 ; n52757
g52502 and n52693_not n52696_not ; n52758
g52503 and n52757_not n52758_not ; n52759
g52504 and n52728_not n52759_not ; n52760
g52505 and n51954_not n52727_not ; n52761
g52506 and n52726_not n52761 ; n52762
g52507 and n52760_not n52762_not ; n52763
g52508 and b[55]_not n52763_not ; n52764
g52509 and n51973_not n52691 ; n52765
g52510 and n52687_not n52765 ; n52766
g52511 and n52688_not n52691_not ; n52767
g52512 and n52766_not n52767_not ; n52768
g52513 and n52728_not n52768_not ; n52769
g52514 and n51963_not n52727_not ; n52770
g52515 and n52726_not n52770 ; n52771
g52516 and n52769_not n52771_not ; n52772
g52517 and b[54]_not n52772_not ; n52773
g52518 and n51982_not n52686 ; n52774
g52519 and n52682_not n52774 ; n52775
g52520 and n52683_not n52686_not ; n52776
g52521 and n52775_not n52776_not ; n52777
g52522 and n52728_not n52777_not ; n52778
g52523 and n51972_not n52727_not ; n52779
g52524 and n52726_not n52779 ; n52780
g52525 and n52778_not n52780_not ; n52781
g52526 and b[53]_not n52781_not ; n52782
g52527 and n51991_not n52681 ; n52783
g52528 and n52677_not n52783 ; n52784
g52529 and n52678_not n52681_not ; n52785
g52530 and n52784_not n52785_not ; n52786
g52531 and n52728_not n52786_not ; n52787
g52532 and n51981_not n52727_not ; n52788
g52533 and n52726_not n52788 ; n52789
g52534 and n52787_not n52789_not ; n52790
g52535 and b[52]_not n52790_not ; n52791
g52536 and n52000_not n52676 ; n52792
g52537 and n52672_not n52792 ; n52793
g52538 and n52673_not n52676_not ; n52794
g52539 and n52793_not n52794_not ; n52795
g52540 and n52728_not n52795_not ; n52796
g52541 and n51990_not n52727_not ; n52797
g52542 and n52726_not n52797 ; n52798
g52543 and n52796_not n52798_not ; n52799
g52544 and b[51]_not n52799_not ; n52800
g52545 and n52009_not n52671 ; n52801
g52546 and n52667_not n52801 ; n52802
g52547 and n52668_not n52671_not ; n52803
g52548 and n52802_not n52803_not ; n52804
g52549 and n52728_not n52804_not ; n52805
g52550 and n51999_not n52727_not ; n52806
g52551 and n52726_not n52806 ; n52807
g52552 and n52805_not n52807_not ; n52808
g52553 and b[50]_not n52808_not ; n52809
g52554 and n52018_not n52666 ; n52810
g52555 and n52662_not n52810 ; n52811
g52556 and n52663_not n52666_not ; n52812
g52557 and n52811_not n52812_not ; n52813
g52558 and n52728_not n52813_not ; n52814
g52559 and n52008_not n52727_not ; n52815
g52560 and n52726_not n52815 ; n52816
g52561 and n52814_not n52816_not ; n52817
g52562 and b[49]_not n52817_not ; n52818
g52563 and n52027_not n52661 ; n52819
g52564 and n52657_not n52819 ; n52820
g52565 and n52658_not n52661_not ; n52821
g52566 and n52820_not n52821_not ; n52822
g52567 and n52728_not n52822_not ; n52823
g52568 and n52017_not n52727_not ; n52824
g52569 and n52726_not n52824 ; n52825
g52570 and n52823_not n52825_not ; n52826
g52571 and b[48]_not n52826_not ; n52827
g52572 and n52036_not n52656 ; n52828
g52573 and n52652_not n52828 ; n52829
g52574 and n52653_not n52656_not ; n52830
g52575 and n52829_not n52830_not ; n52831
g52576 and n52728_not n52831_not ; n52832
g52577 and n52026_not n52727_not ; n52833
g52578 and n52726_not n52833 ; n52834
g52579 and n52832_not n52834_not ; n52835
g52580 and b[47]_not n52835_not ; n52836
g52581 and n52045_not n52651 ; n52837
g52582 and n52647_not n52837 ; n52838
g52583 and n52648_not n52651_not ; n52839
g52584 and n52838_not n52839_not ; n52840
g52585 and n52728_not n52840_not ; n52841
g52586 and n52035_not n52727_not ; n52842
g52587 and n52726_not n52842 ; n52843
g52588 and n52841_not n52843_not ; n52844
g52589 and b[46]_not n52844_not ; n52845
g52590 and n52054_not n52646 ; n52846
g52591 and n52642_not n52846 ; n52847
g52592 and n52643_not n52646_not ; n52848
g52593 and n52847_not n52848_not ; n52849
g52594 and n52728_not n52849_not ; n52850
g52595 and n52044_not n52727_not ; n52851
g52596 and n52726_not n52851 ; n52852
g52597 and n52850_not n52852_not ; n52853
g52598 and b[45]_not n52853_not ; n52854
g52599 and n52063_not n52641 ; n52855
g52600 and n52637_not n52855 ; n52856
g52601 and n52638_not n52641_not ; n52857
g52602 and n52856_not n52857_not ; n52858
g52603 and n52728_not n52858_not ; n52859
g52604 and n52053_not n52727_not ; n52860
g52605 and n52726_not n52860 ; n52861
g52606 and n52859_not n52861_not ; n52862
g52607 and b[44]_not n52862_not ; n52863
g52608 and n52072_not n52636 ; n52864
g52609 and n52632_not n52864 ; n52865
g52610 and n52633_not n52636_not ; n52866
g52611 and n52865_not n52866_not ; n52867
g52612 and n52728_not n52867_not ; n52868
g52613 and n52062_not n52727_not ; n52869
g52614 and n52726_not n52869 ; n52870
g52615 and n52868_not n52870_not ; n52871
g52616 and b[43]_not n52871_not ; n52872
g52617 and n52081_not n52631 ; n52873
g52618 and n52627_not n52873 ; n52874
g52619 and n52628_not n52631_not ; n52875
g52620 and n52874_not n52875_not ; n52876
g52621 and n52728_not n52876_not ; n52877
g52622 and n52071_not n52727_not ; n52878
g52623 and n52726_not n52878 ; n52879
g52624 and n52877_not n52879_not ; n52880
g52625 and b[42]_not n52880_not ; n52881
g52626 and n52090_not n52626 ; n52882
g52627 and n52622_not n52882 ; n52883
g52628 and n52623_not n52626_not ; n52884
g52629 and n52883_not n52884_not ; n52885
g52630 and n52728_not n52885_not ; n52886
g52631 and n52080_not n52727_not ; n52887
g52632 and n52726_not n52887 ; n52888
g52633 and n52886_not n52888_not ; n52889
g52634 and b[41]_not n52889_not ; n52890
g52635 and n52099_not n52621 ; n52891
g52636 and n52617_not n52891 ; n52892
g52637 and n52618_not n52621_not ; n52893
g52638 and n52892_not n52893_not ; n52894
g52639 and n52728_not n52894_not ; n52895
g52640 and n52089_not n52727_not ; n52896
g52641 and n52726_not n52896 ; n52897
g52642 and n52895_not n52897_not ; n52898
g52643 and b[40]_not n52898_not ; n52899
g52644 and n52108_not n52616 ; n52900
g52645 and n52612_not n52900 ; n52901
g52646 and n52613_not n52616_not ; n52902
g52647 and n52901_not n52902_not ; n52903
g52648 and n52728_not n52903_not ; n52904
g52649 and n52098_not n52727_not ; n52905
g52650 and n52726_not n52905 ; n52906
g52651 and n52904_not n52906_not ; n52907
g52652 and b[39]_not n52907_not ; n52908
g52653 and n52117_not n52611 ; n52909
g52654 and n52607_not n52909 ; n52910
g52655 and n52608_not n52611_not ; n52911
g52656 and n52910_not n52911_not ; n52912
g52657 and n52728_not n52912_not ; n52913
g52658 and n52107_not n52727_not ; n52914
g52659 and n52726_not n52914 ; n52915
g52660 and n52913_not n52915_not ; n52916
g52661 and b[38]_not n52916_not ; n52917
g52662 and n52126_not n52606 ; n52918
g52663 and n52602_not n52918 ; n52919
g52664 and n52603_not n52606_not ; n52920
g52665 and n52919_not n52920_not ; n52921
g52666 and n52728_not n52921_not ; n52922
g52667 and n52116_not n52727_not ; n52923
g52668 and n52726_not n52923 ; n52924
g52669 and n52922_not n52924_not ; n52925
g52670 and b[37]_not n52925_not ; n52926
g52671 and n52135_not n52601 ; n52927
g52672 and n52597_not n52927 ; n52928
g52673 and n52598_not n52601_not ; n52929
g52674 and n52928_not n52929_not ; n52930
g52675 and n52728_not n52930_not ; n52931
g52676 and n52125_not n52727_not ; n52932
g52677 and n52726_not n52932 ; n52933
g52678 and n52931_not n52933_not ; n52934
g52679 and b[36]_not n52934_not ; n52935
g52680 and n52144_not n52596 ; n52936
g52681 and n52592_not n52936 ; n52937
g52682 and n52593_not n52596_not ; n52938
g52683 and n52937_not n52938_not ; n52939
g52684 and n52728_not n52939_not ; n52940
g52685 and n52134_not n52727_not ; n52941
g52686 and n52726_not n52941 ; n52942
g52687 and n52940_not n52942_not ; n52943
g52688 and b[35]_not n52943_not ; n52944
g52689 and n52153_not n52591 ; n52945
g52690 and n52587_not n52945 ; n52946
g52691 and n52588_not n52591_not ; n52947
g52692 and n52946_not n52947_not ; n52948
g52693 and n52728_not n52948_not ; n52949
g52694 and n52143_not n52727_not ; n52950
g52695 and n52726_not n52950 ; n52951
g52696 and n52949_not n52951_not ; n52952
g52697 and b[34]_not n52952_not ; n52953
g52698 and n52162_not n52586 ; n52954
g52699 and n52582_not n52954 ; n52955
g52700 and n52583_not n52586_not ; n52956
g52701 and n52955_not n52956_not ; n52957
g52702 and n52728_not n52957_not ; n52958
g52703 and n52152_not n52727_not ; n52959
g52704 and n52726_not n52959 ; n52960
g52705 and n52958_not n52960_not ; n52961
g52706 and b[33]_not n52961_not ; n52962
g52707 and n52171_not n52581 ; n52963
g52708 and n52577_not n52963 ; n52964
g52709 and n52578_not n52581_not ; n52965
g52710 and n52964_not n52965_not ; n52966
g52711 and n52728_not n52966_not ; n52967
g52712 and n52161_not n52727_not ; n52968
g52713 and n52726_not n52968 ; n52969
g52714 and n52967_not n52969_not ; n52970
g52715 and b[32]_not n52970_not ; n52971
g52716 and n52180_not n52576 ; n52972
g52717 and n52572_not n52972 ; n52973
g52718 and n52573_not n52576_not ; n52974
g52719 and n52973_not n52974_not ; n52975
g52720 and n52728_not n52975_not ; n52976
g52721 and n52170_not n52727_not ; n52977
g52722 and n52726_not n52977 ; n52978
g52723 and n52976_not n52978_not ; n52979
g52724 and b[31]_not n52979_not ; n52980
g52725 and n52189_not n52571 ; n52981
g52726 and n52567_not n52981 ; n52982
g52727 and n52568_not n52571_not ; n52983
g52728 and n52982_not n52983_not ; n52984
g52729 and n52728_not n52984_not ; n52985
g52730 and n52179_not n52727_not ; n52986
g52731 and n52726_not n52986 ; n52987
g52732 and n52985_not n52987_not ; n52988
g52733 and b[30]_not n52988_not ; n52989
g52734 and n52198_not n52566 ; n52990
g52735 and n52562_not n52990 ; n52991
g52736 and n52563_not n52566_not ; n52992
g52737 and n52991_not n52992_not ; n52993
g52738 and n52728_not n52993_not ; n52994
g52739 and n52188_not n52727_not ; n52995
g52740 and n52726_not n52995 ; n52996
g52741 and n52994_not n52996_not ; n52997
g52742 and b[29]_not n52997_not ; n52998
g52743 and n52207_not n52561 ; n52999
g52744 and n52557_not n52999 ; n53000
g52745 and n52558_not n52561_not ; n53001
g52746 and n53000_not n53001_not ; n53002
g52747 and n52728_not n53002_not ; n53003
g52748 and n52197_not n52727_not ; n53004
g52749 and n52726_not n53004 ; n53005
g52750 and n53003_not n53005_not ; n53006
g52751 and b[28]_not n53006_not ; n53007
g52752 and n52216_not n52556 ; n53008
g52753 and n52552_not n53008 ; n53009
g52754 and n52553_not n52556_not ; n53010
g52755 and n53009_not n53010_not ; n53011
g52756 and n52728_not n53011_not ; n53012
g52757 and n52206_not n52727_not ; n53013
g52758 and n52726_not n53013 ; n53014
g52759 and n53012_not n53014_not ; n53015
g52760 and b[27]_not n53015_not ; n53016
g52761 and n52225_not n52551 ; n53017
g52762 and n52547_not n53017 ; n53018
g52763 and n52548_not n52551_not ; n53019
g52764 and n53018_not n53019_not ; n53020
g52765 and n52728_not n53020_not ; n53021
g52766 and n52215_not n52727_not ; n53022
g52767 and n52726_not n53022 ; n53023
g52768 and n53021_not n53023_not ; n53024
g52769 and b[26]_not n53024_not ; n53025
g52770 and n52234_not n52546 ; n53026
g52771 and n52542_not n53026 ; n53027
g52772 and n52543_not n52546_not ; n53028
g52773 and n53027_not n53028_not ; n53029
g52774 and n52728_not n53029_not ; n53030
g52775 and n52224_not n52727_not ; n53031
g52776 and n52726_not n53031 ; n53032
g52777 and n53030_not n53032_not ; n53033
g52778 and b[25]_not n53033_not ; n53034
g52779 and n52243_not n52541 ; n53035
g52780 and n52537_not n53035 ; n53036
g52781 and n52538_not n52541_not ; n53037
g52782 and n53036_not n53037_not ; n53038
g52783 and n52728_not n53038_not ; n53039
g52784 and n52233_not n52727_not ; n53040
g52785 and n52726_not n53040 ; n53041
g52786 and n53039_not n53041_not ; n53042
g52787 and b[24]_not n53042_not ; n53043
g52788 and n52252_not n52536 ; n53044
g52789 and n52532_not n53044 ; n53045
g52790 and n52533_not n52536_not ; n53046
g52791 and n53045_not n53046_not ; n53047
g52792 and n52728_not n53047_not ; n53048
g52793 and n52242_not n52727_not ; n53049
g52794 and n52726_not n53049 ; n53050
g52795 and n53048_not n53050_not ; n53051
g52796 and b[23]_not n53051_not ; n53052
g52797 and n52261_not n52531 ; n53053
g52798 and n52527_not n53053 ; n53054
g52799 and n52528_not n52531_not ; n53055
g52800 and n53054_not n53055_not ; n53056
g52801 and n52728_not n53056_not ; n53057
g52802 and n52251_not n52727_not ; n53058
g52803 and n52726_not n53058 ; n53059
g52804 and n53057_not n53059_not ; n53060
g52805 and b[22]_not n53060_not ; n53061
g52806 and n52270_not n52526 ; n53062
g52807 and n52522_not n53062 ; n53063
g52808 and n52523_not n52526_not ; n53064
g52809 and n53063_not n53064_not ; n53065
g52810 and n52728_not n53065_not ; n53066
g52811 and n52260_not n52727_not ; n53067
g52812 and n52726_not n53067 ; n53068
g52813 and n53066_not n53068_not ; n53069
g52814 and b[21]_not n53069_not ; n53070
g52815 and n52279_not n52521 ; n53071
g52816 and n52517_not n53071 ; n53072
g52817 and n52518_not n52521_not ; n53073
g52818 and n53072_not n53073_not ; n53074
g52819 and n52728_not n53074_not ; n53075
g52820 and n52269_not n52727_not ; n53076
g52821 and n52726_not n53076 ; n53077
g52822 and n53075_not n53077_not ; n53078
g52823 and b[20]_not n53078_not ; n53079
g52824 and n52288_not n52516 ; n53080
g52825 and n52512_not n53080 ; n53081
g52826 and n52513_not n52516_not ; n53082
g52827 and n53081_not n53082_not ; n53083
g52828 and n52728_not n53083_not ; n53084
g52829 and n52278_not n52727_not ; n53085
g52830 and n52726_not n53085 ; n53086
g52831 and n53084_not n53086_not ; n53087
g52832 and b[19]_not n53087_not ; n53088
g52833 and n52297_not n52511 ; n53089
g52834 and n52507_not n53089 ; n53090
g52835 and n52508_not n52511_not ; n53091
g52836 and n53090_not n53091_not ; n53092
g52837 and n52728_not n53092_not ; n53093
g52838 and n52287_not n52727_not ; n53094
g52839 and n52726_not n53094 ; n53095
g52840 and n53093_not n53095_not ; n53096
g52841 and b[18]_not n53096_not ; n53097
g52842 and n52306_not n52506 ; n53098
g52843 and n52502_not n53098 ; n53099
g52844 and n52503_not n52506_not ; n53100
g52845 and n53099_not n53100_not ; n53101
g52846 and n52728_not n53101_not ; n53102
g52847 and n52296_not n52727_not ; n53103
g52848 and n52726_not n53103 ; n53104
g52849 and n53102_not n53104_not ; n53105
g52850 and b[17]_not n53105_not ; n53106
g52851 and n52315_not n52501 ; n53107
g52852 and n52497_not n53107 ; n53108
g52853 and n52498_not n52501_not ; n53109
g52854 and n53108_not n53109_not ; n53110
g52855 and n52728_not n53110_not ; n53111
g52856 and n52305_not n52727_not ; n53112
g52857 and n52726_not n53112 ; n53113
g52858 and n53111_not n53113_not ; n53114
g52859 and b[16]_not n53114_not ; n53115
g52860 and n52324_not n52496 ; n53116
g52861 and n52492_not n53116 ; n53117
g52862 and n52493_not n52496_not ; n53118
g52863 and n53117_not n53118_not ; n53119
g52864 and n52728_not n53119_not ; n53120
g52865 and n52314_not n52727_not ; n53121
g52866 and n52726_not n53121 ; n53122
g52867 and n53120_not n53122_not ; n53123
g52868 and b[15]_not n53123_not ; n53124
g52869 and n52333_not n52491 ; n53125
g52870 and n52487_not n53125 ; n53126
g52871 and n52488_not n52491_not ; n53127
g52872 and n53126_not n53127_not ; n53128
g52873 and n52728_not n53128_not ; n53129
g52874 and n52323_not n52727_not ; n53130
g52875 and n52726_not n53130 ; n53131
g52876 and n53129_not n53131_not ; n53132
g52877 and b[14]_not n53132_not ; n53133
g52878 and n52342_not n52486 ; n53134
g52879 and n52482_not n53134 ; n53135
g52880 and n52483_not n52486_not ; n53136
g52881 and n53135_not n53136_not ; n53137
g52882 and n52728_not n53137_not ; n53138
g52883 and n52332_not n52727_not ; n53139
g52884 and n52726_not n53139 ; n53140
g52885 and n53138_not n53140_not ; n53141
g52886 and b[13]_not n53141_not ; n53142
g52887 and n52351_not n52481 ; n53143
g52888 and n52477_not n53143 ; n53144
g52889 and n52478_not n52481_not ; n53145
g52890 and n53144_not n53145_not ; n53146
g52891 and n52728_not n53146_not ; n53147
g52892 and n52341_not n52727_not ; n53148
g52893 and n52726_not n53148 ; n53149
g52894 and n53147_not n53149_not ; n53150
g52895 and b[12]_not n53150_not ; n53151
g52896 and n52360_not n52476 ; n53152
g52897 and n52472_not n53152 ; n53153
g52898 and n52473_not n52476_not ; n53154
g52899 and n53153_not n53154_not ; n53155
g52900 and n52728_not n53155_not ; n53156
g52901 and n52350_not n52727_not ; n53157
g52902 and n52726_not n53157 ; n53158
g52903 and n53156_not n53158_not ; n53159
g52904 and b[11]_not n53159_not ; n53160
g52905 and n52369_not n52471 ; n53161
g52906 and n52467_not n53161 ; n53162
g52907 and n52468_not n52471_not ; n53163
g52908 and n53162_not n53163_not ; n53164
g52909 and n52728_not n53164_not ; n53165
g52910 and n52359_not n52727_not ; n53166
g52911 and n52726_not n53166 ; n53167
g52912 and n53165_not n53167_not ; n53168
g52913 and b[10]_not n53168_not ; n53169
g52914 and n52378_not n52466 ; n53170
g52915 and n52462_not n53170 ; n53171
g52916 and n52463_not n52466_not ; n53172
g52917 and n53171_not n53172_not ; n53173
g52918 and n52728_not n53173_not ; n53174
g52919 and n52368_not n52727_not ; n53175
g52920 and n52726_not n53175 ; n53176
g52921 and n53174_not n53176_not ; n53177
g52922 and b[9]_not n53177_not ; n53178
g52923 and n52387_not n52461 ; n53179
g52924 and n52457_not n53179 ; n53180
g52925 and n52458_not n52461_not ; n53181
g52926 and n53180_not n53181_not ; n53182
g52927 and n52728_not n53182_not ; n53183
g52928 and n52377_not n52727_not ; n53184
g52929 and n52726_not n53184 ; n53185
g52930 and n53183_not n53185_not ; n53186
g52931 and b[8]_not n53186_not ; n53187
g52932 and n52396_not n52456 ; n53188
g52933 and n52452_not n53188 ; n53189
g52934 and n52453_not n52456_not ; n53190
g52935 and n53189_not n53190_not ; n53191
g52936 and n52728_not n53191_not ; n53192
g52937 and n52386_not n52727_not ; n53193
g52938 and n52726_not n53193 ; n53194
g52939 and n53192_not n53194_not ; n53195
g52940 and b[7]_not n53195_not ; n53196
g52941 and n52405_not n52451 ; n53197
g52942 and n52447_not n53197 ; n53198
g52943 and n52448_not n52451_not ; n53199
g52944 and n53198_not n53199_not ; n53200
g52945 and n52728_not n53200_not ; n53201
g52946 and n52395_not n52727_not ; n53202
g52947 and n52726_not n53202 ; n53203
g52948 and n53201_not n53203_not ; n53204
g52949 and b[6]_not n53204_not ; n53205
g52950 and n52414_not n52446 ; n53206
g52951 and n52442_not n53206 ; n53207
g52952 and n52443_not n52446_not ; n53208
g52953 and n53207_not n53208_not ; n53209
g52954 and n52728_not n53209_not ; n53210
g52955 and n52404_not n52727_not ; n53211
g52956 and n52726_not n53211 ; n53212
g52957 and n53210_not n53212_not ; n53213
g52958 and b[5]_not n53213_not ; n53214
g52959 and n52422_not n52441 ; n53215
g52960 and n52437_not n53215 ; n53216
g52961 and n52438_not n52441_not ; n53217
g52962 and n53216_not n53217_not ; n53218
g52963 and n52728_not n53218_not ; n53219
g52964 and n52413_not n52727_not ; n53220
g52965 and n52726_not n53220 ; n53221
g52966 and n53219_not n53221_not ; n53222
g52967 and b[4]_not n53222_not ; n53223
g52968 and n52432_not n52436 ; n53224
g52969 and n52431_not n53224 ; n53225
g52970 and n52433_not n52436_not ; n53226
g52971 and n53225_not n53226_not ; n53227
g52972 and n52728_not n53227_not ; n53228
g52973 and n52421_not n52727_not ; n53229
g52974 and n52726_not n53229 ; n53230
g52975 and n53228_not n53230_not ; n53231
g52976 and b[3]_not n53231_not ; n53232
g52977 and n24413 n52429_not ; n53233
g52978 and n52427_not n53233 ; n53234
g52979 and n52431_not n53234_not ; n53235
g52980 and n52728_not n53235 ; n53236
g52981 and n52426_not n52727_not ; n53237
g52982 and n52726_not n53237 ; n53238
g52983 and n53236_not n53238_not ; n53239
g52984 and b[2]_not n53239_not ; n53240
g52985 and b[0] n52728_not ; n53241
g52986 and a[5] n53241_not ; n53242
g52987 and n24413 n52728_not ; n53243
g52988 and n53242_not n53243_not ; n53244
g52989 and b[1] n53244_not ; n53245
g52990 and b[1]_not n53243_not ; n53246
g52991 and n53242_not n53246 ; n53247
g52992 and n53245_not n53247_not ; n53248
g52993 and n25233_not n53248_not ; n53249
g52994 and b[1]_not n53244_not ; n53250
g52995 and n53249_not n53250_not ; n53251
g52996 and b[2] n53238_not ; n53252
g52997 and n53236_not n53252 ; n53253
g52998 and n53240_not n53253_not ; n53254
g52999 and n53251_not n53254 ; n53255
g53000 and n53240_not n53255_not ; n53256
g53001 and b[3] n53230_not ; n53257
g53002 and n53228_not n53257 ; n53258
g53003 and n53232_not n53258_not ; n53259
g53004 and n53256_not n53259 ; n53260
g53005 and n53232_not n53260_not ; n53261
g53006 and b[4] n53221_not ; n53262
g53007 and n53219_not n53262 ; n53263
g53008 and n53223_not n53263_not ; n53264
g53009 and n53261_not n53264 ; n53265
g53010 and n53223_not n53265_not ; n53266
g53011 and b[5] n53212_not ; n53267
g53012 and n53210_not n53267 ; n53268
g53013 and n53214_not n53268_not ; n53269
g53014 and n53266_not n53269 ; n53270
g53015 and n53214_not n53270_not ; n53271
g53016 and b[6] n53203_not ; n53272
g53017 and n53201_not n53272 ; n53273
g53018 and n53205_not n53273_not ; n53274
g53019 and n53271_not n53274 ; n53275
g53020 and n53205_not n53275_not ; n53276
g53021 and b[7] n53194_not ; n53277
g53022 and n53192_not n53277 ; n53278
g53023 and n53196_not n53278_not ; n53279
g53024 and n53276_not n53279 ; n53280
g53025 and n53196_not n53280_not ; n53281
g53026 and b[8] n53185_not ; n53282
g53027 and n53183_not n53282 ; n53283
g53028 and n53187_not n53283_not ; n53284
g53029 and n53281_not n53284 ; n53285
g53030 and n53187_not n53285_not ; n53286
g53031 and b[9] n53176_not ; n53287
g53032 and n53174_not n53287 ; n53288
g53033 and n53178_not n53288_not ; n53289
g53034 and n53286_not n53289 ; n53290
g53035 and n53178_not n53290_not ; n53291
g53036 and b[10] n53167_not ; n53292
g53037 and n53165_not n53292 ; n53293
g53038 and n53169_not n53293_not ; n53294
g53039 and n53291_not n53294 ; n53295
g53040 and n53169_not n53295_not ; n53296
g53041 and b[11] n53158_not ; n53297
g53042 and n53156_not n53297 ; n53298
g53043 and n53160_not n53298_not ; n53299
g53044 and n53296_not n53299 ; n53300
g53045 and n53160_not n53300_not ; n53301
g53046 and b[12] n53149_not ; n53302
g53047 and n53147_not n53302 ; n53303
g53048 and n53151_not n53303_not ; n53304
g53049 and n53301_not n53304 ; n53305
g53050 and n53151_not n53305_not ; n53306
g53051 and b[13] n53140_not ; n53307
g53052 and n53138_not n53307 ; n53308
g53053 and n53142_not n53308_not ; n53309
g53054 and n53306_not n53309 ; n53310
g53055 and n53142_not n53310_not ; n53311
g53056 and b[14] n53131_not ; n53312
g53057 and n53129_not n53312 ; n53313
g53058 and n53133_not n53313_not ; n53314
g53059 and n53311_not n53314 ; n53315
g53060 and n53133_not n53315_not ; n53316
g53061 and b[15] n53122_not ; n53317
g53062 and n53120_not n53317 ; n53318
g53063 and n53124_not n53318_not ; n53319
g53064 and n53316_not n53319 ; n53320
g53065 and n53124_not n53320_not ; n53321
g53066 and b[16] n53113_not ; n53322
g53067 and n53111_not n53322 ; n53323
g53068 and n53115_not n53323_not ; n53324
g53069 and n53321_not n53324 ; n53325
g53070 and n53115_not n53325_not ; n53326
g53071 and b[17] n53104_not ; n53327
g53072 and n53102_not n53327 ; n53328
g53073 and n53106_not n53328_not ; n53329
g53074 and n53326_not n53329 ; n53330
g53075 and n53106_not n53330_not ; n53331
g53076 and b[18] n53095_not ; n53332
g53077 and n53093_not n53332 ; n53333
g53078 and n53097_not n53333_not ; n53334
g53079 and n53331_not n53334 ; n53335
g53080 and n53097_not n53335_not ; n53336
g53081 and b[19] n53086_not ; n53337
g53082 and n53084_not n53337 ; n53338
g53083 and n53088_not n53338_not ; n53339
g53084 and n53336_not n53339 ; n53340
g53085 and n53088_not n53340_not ; n53341
g53086 and b[20] n53077_not ; n53342
g53087 and n53075_not n53342 ; n53343
g53088 and n53079_not n53343_not ; n53344
g53089 and n53341_not n53344 ; n53345
g53090 and n53079_not n53345_not ; n53346
g53091 and b[21] n53068_not ; n53347
g53092 and n53066_not n53347 ; n53348
g53093 and n53070_not n53348_not ; n53349
g53094 and n53346_not n53349 ; n53350
g53095 and n53070_not n53350_not ; n53351
g53096 and b[22] n53059_not ; n53352
g53097 and n53057_not n53352 ; n53353
g53098 and n53061_not n53353_not ; n53354
g53099 and n53351_not n53354 ; n53355
g53100 and n53061_not n53355_not ; n53356
g53101 and b[23] n53050_not ; n53357
g53102 and n53048_not n53357 ; n53358
g53103 and n53052_not n53358_not ; n53359
g53104 and n53356_not n53359 ; n53360
g53105 and n53052_not n53360_not ; n53361
g53106 and b[24] n53041_not ; n53362
g53107 and n53039_not n53362 ; n53363
g53108 and n53043_not n53363_not ; n53364
g53109 and n53361_not n53364 ; n53365
g53110 and n53043_not n53365_not ; n53366
g53111 and b[25] n53032_not ; n53367
g53112 and n53030_not n53367 ; n53368
g53113 and n53034_not n53368_not ; n53369
g53114 and n53366_not n53369 ; n53370
g53115 and n53034_not n53370_not ; n53371
g53116 and b[26] n53023_not ; n53372
g53117 and n53021_not n53372 ; n53373
g53118 and n53025_not n53373_not ; n53374
g53119 and n53371_not n53374 ; n53375
g53120 and n53025_not n53375_not ; n53376
g53121 and b[27] n53014_not ; n53377
g53122 and n53012_not n53377 ; n53378
g53123 and n53016_not n53378_not ; n53379
g53124 and n53376_not n53379 ; n53380
g53125 and n53016_not n53380_not ; n53381
g53126 and b[28] n53005_not ; n53382
g53127 and n53003_not n53382 ; n53383
g53128 and n53007_not n53383_not ; n53384
g53129 and n53381_not n53384 ; n53385
g53130 and n53007_not n53385_not ; n53386
g53131 and b[29] n52996_not ; n53387
g53132 and n52994_not n53387 ; n53388
g53133 and n52998_not n53388_not ; n53389
g53134 and n53386_not n53389 ; n53390
g53135 and n52998_not n53390_not ; n53391
g53136 and b[30] n52987_not ; n53392
g53137 and n52985_not n53392 ; n53393
g53138 and n52989_not n53393_not ; n53394
g53139 and n53391_not n53394 ; n53395
g53140 and n52989_not n53395_not ; n53396
g53141 and b[31] n52978_not ; n53397
g53142 and n52976_not n53397 ; n53398
g53143 and n52980_not n53398_not ; n53399
g53144 and n53396_not n53399 ; n53400
g53145 and n52980_not n53400_not ; n53401
g53146 and b[32] n52969_not ; n53402
g53147 and n52967_not n53402 ; n53403
g53148 and n52971_not n53403_not ; n53404
g53149 and n53401_not n53404 ; n53405
g53150 and n52971_not n53405_not ; n53406
g53151 and b[33] n52960_not ; n53407
g53152 and n52958_not n53407 ; n53408
g53153 and n52962_not n53408_not ; n53409
g53154 and n53406_not n53409 ; n53410
g53155 and n52962_not n53410_not ; n53411
g53156 and b[34] n52951_not ; n53412
g53157 and n52949_not n53412 ; n53413
g53158 and n52953_not n53413_not ; n53414
g53159 and n53411_not n53414 ; n53415
g53160 and n52953_not n53415_not ; n53416
g53161 and b[35] n52942_not ; n53417
g53162 and n52940_not n53417 ; n53418
g53163 and n52944_not n53418_not ; n53419
g53164 and n53416_not n53419 ; n53420
g53165 and n52944_not n53420_not ; n53421
g53166 and b[36] n52933_not ; n53422
g53167 and n52931_not n53422 ; n53423
g53168 and n52935_not n53423_not ; n53424
g53169 and n53421_not n53424 ; n53425
g53170 and n52935_not n53425_not ; n53426
g53171 and b[37] n52924_not ; n53427
g53172 and n52922_not n53427 ; n53428
g53173 and n52926_not n53428_not ; n53429
g53174 and n53426_not n53429 ; n53430
g53175 and n52926_not n53430_not ; n53431
g53176 and b[38] n52915_not ; n53432
g53177 and n52913_not n53432 ; n53433
g53178 and n52917_not n53433_not ; n53434
g53179 and n53431_not n53434 ; n53435
g53180 and n52917_not n53435_not ; n53436
g53181 and b[39] n52906_not ; n53437
g53182 and n52904_not n53437 ; n53438
g53183 and n52908_not n53438_not ; n53439
g53184 and n53436_not n53439 ; n53440
g53185 and n52908_not n53440_not ; n53441
g53186 and b[40] n52897_not ; n53442
g53187 and n52895_not n53442 ; n53443
g53188 and n52899_not n53443_not ; n53444
g53189 and n53441_not n53444 ; n53445
g53190 and n52899_not n53445_not ; n53446
g53191 and b[41] n52888_not ; n53447
g53192 and n52886_not n53447 ; n53448
g53193 and n52890_not n53448_not ; n53449
g53194 and n53446_not n53449 ; n53450
g53195 and n52890_not n53450_not ; n53451
g53196 and b[42] n52879_not ; n53452
g53197 and n52877_not n53452 ; n53453
g53198 and n52881_not n53453_not ; n53454
g53199 and n53451_not n53454 ; n53455
g53200 and n52881_not n53455_not ; n53456
g53201 and b[43] n52870_not ; n53457
g53202 and n52868_not n53457 ; n53458
g53203 and n52872_not n53458_not ; n53459
g53204 and n53456_not n53459 ; n53460
g53205 and n52872_not n53460_not ; n53461
g53206 and b[44] n52861_not ; n53462
g53207 and n52859_not n53462 ; n53463
g53208 and n52863_not n53463_not ; n53464
g53209 and n53461_not n53464 ; n53465
g53210 and n52863_not n53465_not ; n53466
g53211 and b[45] n52852_not ; n53467
g53212 and n52850_not n53467 ; n53468
g53213 and n52854_not n53468_not ; n53469
g53214 and n53466_not n53469 ; n53470
g53215 and n52854_not n53470_not ; n53471
g53216 and b[46] n52843_not ; n53472
g53217 and n52841_not n53472 ; n53473
g53218 and n52845_not n53473_not ; n53474
g53219 and n53471_not n53474 ; n53475
g53220 and n52845_not n53475_not ; n53476
g53221 and b[47] n52834_not ; n53477
g53222 and n52832_not n53477 ; n53478
g53223 and n52836_not n53478_not ; n53479
g53224 and n53476_not n53479 ; n53480
g53225 and n52836_not n53480_not ; n53481
g53226 and b[48] n52825_not ; n53482
g53227 and n52823_not n53482 ; n53483
g53228 and n52827_not n53483_not ; n53484
g53229 and n53481_not n53484 ; n53485
g53230 and n52827_not n53485_not ; n53486
g53231 and b[49] n52816_not ; n53487
g53232 and n52814_not n53487 ; n53488
g53233 and n52818_not n53488_not ; n53489
g53234 and n53486_not n53489 ; n53490
g53235 and n52818_not n53490_not ; n53491
g53236 and b[50] n52807_not ; n53492
g53237 and n52805_not n53492 ; n53493
g53238 and n52809_not n53493_not ; n53494
g53239 and n53491_not n53494 ; n53495
g53240 and n52809_not n53495_not ; n53496
g53241 and b[51] n52798_not ; n53497
g53242 and n52796_not n53497 ; n53498
g53243 and n52800_not n53498_not ; n53499
g53244 and n53496_not n53499 ; n53500
g53245 and n52800_not n53500_not ; n53501
g53246 and b[52] n52789_not ; n53502
g53247 and n52787_not n53502 ; n53503
g53248 and n52791_not n53503_not ; n53504
g53249 and n53501_not n53504 ; n53505
g53250 and n52791_not n53505_not ; n53506
g53251 and b[53] n52780_not ; n53507
g53252 and n52778_not n53507 ; n53508
g53253 and n52782_not n53508_not ; n53509
g53254 and n53506_not n53509 ; n53510
g53255 and n52782_not n53510_not ; n53511
g53256 and b[54] n52771_not ; n53512
g53257 and n52769_not n53512 ; n53513
g53258 and n52773_not n53513_not ; n53514
g53259 and n53511_not n53514 ; n53515
g53260 and n52773_not n53515_not ; n53516
g53261 and b[55] n52762_not ; n53517
g53262 and n52760_not n53517 ; n53518
g53263 and n52764_not n53518_not ; n53519
g53264 and n53516_not n53519 ; n53520
g53265 and n52764_not n53520_not ; n53521
g53266 and b[56] n52753_not ; n53522
g53267 and n52751_not n53522 ; n53523
g53268 and n52755_not n53523_not ; n53524
g53269 and n53521_not n53524 ; n53525
g53270 and n52755_not n53525_not ; n53526
g53271 and b[57] n52744_not ; n53527
g53272 and n52742_not n53527 ; n53528
g53273 and n52746_not n53528_not ; n53529
g53274 and n53526_not n53529 ; n53530
g53275 and n52746_not n53530_not ; n53531
g53276 and b[58] n52735_not ; n53532
g53277 and n52733_not n53532 ; n53533
g53278 and n52737_not n53533_not ; n53534
g53279 and n53531_not n53534 ; n53535
g53280 and n52737_not n53535_not ; n53536
g53281 and n51928_not n52723_not ; n53537
g53282 and n52721_not n53537 ; n53538
g53283 and n52712_not n53538 ; n53539
g53284 and n52721_not n52723_not ; n53540
g53285 and n52713_not n53540_not ; n53541
g53286 and n53539_not n53541_not ; n53542
g53287 and n52728_not n53542_not ; n53543
g53288 and n52720_not n52727_not ; n53544
g53289 and n52726_not n53544 ; n53545
g53290 and n53543_not n53545_not ; n53546
g53291 and b[59]_not n53546_not ; n53547
g53292 and b[59] n53545_not ; n53548
g53293 and n53543_not n53548 ; n53549
g53294 and n280 n53549_not ; n53550
g53295 and n53547_not n53550 ; n53551
g53296 and n53536_not n53551 ; n53552
g53297 and n24707 n53546_not ; n53553
g53298 and n53552_not n53553_not ; n53554
g53299 and n52746_not n53534 ; n53555
g53300 and n53530_not n53555 ; n53556
g53301 and n53531_not n53534_not ; n53557
g53302 and n53556_not n53557_not ; n53558
g53303 and n53554_not n53558_not ; n53559
g53304 and n52736_not n53553_not ; n53560
g53305 and n53552_not n53560 ; n53561
g53306 and n53559_not n53561_not ; n53562
g53307 and b[59]_not n53562_not ; n53563
g53308 and n52755_not n53529 ; n53564
g53309 and n53525_not n53564 ; n53565
g53310 and n53526_not n53529_not ; n53566
g53311 and n53565_not n53566_not ; n53567
g53312 and n53554_not n53567_not ; n53568
g53313 and n52745_not n53553_not ; n53569
g53314 and n53552_not n53569 ; n53570
g53315 and n53568_not n53570_not ; n53571
g53316 and b[58]_not n53571_not ; n53572
g53317 and n52764_not n53524 ; n53573
g53318 and n53520_not n53573 ; n53574
g53319 and n53521_not n53524_not ; n53575
g53320 and n53574_not n53575_not ; n53576
g53321 and n53554_not n53576_not ; n53577
g53322 and n52754_not n53553_not ; n53578
g53323 and n53552_not n53578 ; n53579
g53324 and n53577_not n53579_not ; n53580
g53325 and b[57]_not n53580_not ; n53581
g53326 and n52773_not n53519 ; n53582
g53327 and n53515_not n53582 ; n53583
g53328 and n53516_not n53519_not ; n53584
g53329 and n53583_not n53584_not ; n53585
g53330 and n53554_not n53585_not ; n53586
g53331 and n52763_not n53553_not ; n53587
g53332 and n53552_not n53587 ; n53588
g53333 and n53586_not n53588_not ; n53589
g53334 and b[56]_not n53589_not ; n53590
g53335 and n52782_not n53514 ; n53591
g53336 and n53510_not n53591 ; n53592
g53337 and n53511_not n53514_not ; n53593
g53338 and n53592_not n53593_not ; n53594
g53339 and n53554_not n53594_not ; n53595
g53340 and n52772_not n53553_not ; n53596
g53341 and n53552_not n53596 ; n53597
g53342 and n53595_not n53597_not ; n53598
g53343 and b[55]_not n53598_not ; n53599
g53344 and n52791_not n53509 ; n53600
g53345 and n53505_not n53600 ; n53601
g53346 and n53506_not n53509_not ; n53602
g53347 and n53601_not n53602_not ; n53603
g53348 and n53554_not n53603_not ; n53604
g53349 and n52781_not n53553_not ; n53605
g53350 and n53552_not n53605 ; n53606
g53351 and n53604_not n53606_not ; n53607
g53352 and b[54]_not n53607_not ; n53608
g53353 and n52800_not n53504 ; n53609
g53354 and n53500_not n53609 ; n53610
g53355 and n53501_not n53504_not ; n53611
g53356 and n53610_not n53611_not ; n53612
g53357 and n53554_not n53612_not ; n53613
g53358 and n52790_not n53553_not ; n53614
g53359 and n53552_not n53614 ; n53615
g53360 and n53613_not n53615_not ; n53616
g53361 and b[53]_not n53616_not ; n53617
g53362 and n52809_not n53499 ; n53618
g53363 and n53495_not n53618 ; n53619
g53364 and n53496_not n53499_not ; n53620
g53365 and n53619_not n53620_not ; n53621
g53366 and n53554_not n53621_not ; n53622
g53367 and n52799_not n53553_not ; n53623
g53368 and n53552_not n53623 ; n53624
g53369 and n53622_not n53624_not ; n53625
g53370 and b[52]_not n53625_not ; n53626
g53371 and n52818_not n53494 ; n53627
g53372 and n53490_not n53627 ; n53628
g53373 and n53491_not n53494_not ; n53629
g53374 and n53628_not n53629_not ; n53630
g53375 and n53554_not n53630_not ; n53631
g53376 and n52808_not n53553_not ; n53632
g53377 and n53552_not n53632 ; n53633
g53378 and n53631_not n53633_not ; n53634
g53379 and b[51]_not n53634_not ; n53635
g53380 and n52827_not n53489 ; n53636
g53381 and n53485_not n53636 ; n53637
g53382 and n53486_not n53489_not ; n53638
g53383 and n53637_not n53638_not ; n53639
g53384 and n53554_not n53639_not ; n53640
g53385 and n52817_not n53553_not ; n53641
g53386 and n53552_not n53641 ; n53642
g53387 and n53640_not n53642_not ; n53643
g53388 and b[50]_not n53643_not ; n53644
g53389 and n52836_not n53484 ; n53645
g53390 and n53480_not n53645 ; n53646
g53391 and n53481_not n53484_not ; n53647
g53392 and n53646_not n53647_not ; n53648
g53393 and n53554_not n53648_not ; n53649
g53394 and n52826_not n53553_not ; n53650
g53395 and n53552_not n53650 ; n53651
g53396 and n53649_not n53651_not ; n53652
g53397 and b[49]_not n53652_not ; n53653
g53398 and n52845_not n53479 ; n53654
g53399 and n53475_not n53654 ; n53655
g53400 and n53476_not n53479_not ; n53656
g53401 and n53655_not n53656_not ; n53657
g53402 and n53554_not n53657_not ; n53658
g53403 and n52835_not n53553_not ; n53659
g53404 and n53552_not n53659 ; n53660
g53405 and n53658_not n53660_not ; n53661
g53406 and b[48]_not n53661_not ; n53662
g53407 and n52854_not n53474 ; n53663
g53408 and n53470_not n53663 ; n53664
g53409 and n53471_not n53474_not ; n53665
g53410 and n53664_not n53665_not ; n53666
g53411 and n53554_not n53666_not ; n53667
g53412 and n52844_not n53553_not ; n53668
g53413 and n53552_not n53668 ; n53669
g53414 and n53667_not n53669_not ; n53670
g53415 and b[47]_not n53670_not ; n53671
g53416 and n52863_not n53469 ; n53672
g53417 and n53465_not n53672 ; n53673
g53418 and n53466_not n53469_not ; n53674
g53419 and n53673_not n53674_not ; n53675
g53420 and n53554_not n53675_not ; n53676
g53421 and n52853_not n53553_not ; n53677
g53422 and n53552_not n53677 ; n53678
g53423 and n53676_not n53678_not ; n53679
g53424 and b[46]_not n53679_not ; n53680
g53425 and n52872_not n53464 ; n53681
g53426 and n53460_not n53681 ; n53682
g53427 and n53461_not n53464_not ; n53683
g53428 and n53682_not n53683_not ; n53684
g53429 and n53554_not n53684_not ; n53685
g53430 and n52862_not n53553_not ; n53686
g53431 and n53552_not n53686 ; n53687
g53432 and n53685_not n53687_not ; n53688
g53433 and b[45]_not n53688_not ; n53689
g53434 and n52881_not n53459 ; n53690
g53435 and n53455_not n53690 ; n53691
g53436 and n53456_not n53459_not ; n53692
g53437 and n53691_not n53692_not ; n53693
g53438 and n53554_not n53693_not ; n53694
g53439 and n52871_not n53553_not ; n53695
g53440 and n53552_not n53695 ; n53696
g53441 and n53694_not n53696_not ; n53697
g53442 and b[44]_not n53697_not ; n53698
g53443 and n52890_not n53454 ; n53699
g53444 and n53450_not n53699 ; n53700
g53445 and n53451_not n53454_not ; n53701
g53446 and n53700_not n53701_not ; n53702
g53447 and n53554_not n53702_not ; n53703
g53448 and n52880_not n53553_not ; n53704
g53449 and n53552_not n53704 ; n53705
g53450 and n53703_not n53705_not ; n53706
g53451 and b[43]_not n53706_not ; n53707
g53452 and n52899_not n53449 ; n53708
g53453 and n53445_not n53708 ; n53709
g53454 and n53446_not n53449_not ; n53710
g53455 and n53709_not n53710_not ; n53711
g53456 and n53554_not n53711_not ; n53712
g53457 and n52889_not n53553_not ; n53713
g53458 and n53552_not n53713 ; n53714
g53459 and n53712_not n53714_not ; n53715
g53460 and b[42]_not n53715_not ; n53716
g53461 and n52908_not n53444 ; n53717
g53462 and n53440_not n53717 ; n53718
g53463 and n53441_not n53444_not ; n53719
g53464 and n53718_not n53719_not ; n53720
g53465 and n53554_not n53720_not ; n53721
g53466 and n52898_not n53553_not ; n53722
g53467 and n53552_not n53722 ; n53723
g53468 and n53721_not n53723_not ; n53724
g53469 and b[41]_not n53724_not ; n53725
g53470 and n52917_not n53439 ; n53726
g53471 and n53435_not n53726 ; n53727
g53472 and n53436_not n53439_not ; n53728
g53473 and n53727_not n53728_not ; n53729
g53474 and n53554_not n53729_not ; n53730
g53475 and n52907_not n53553_not ; n53731
g53476 and n53552_not n53731 ; n53732
g53477 and n53730_not n53732_not ; n53733
g53478 and b[40]_not n53733_not ; n53734
g53479 and n52926_not n53434 ; n53735
g53480 and n53430_not n53735 ; n53736
g53481 and n53431_not n53434_not ; n53737
g53482 and n53736_not n53737_not ; n53738
g53483 and n53554_not n53738_not ; n53739
g53484 and n52916_not n53553_not ; n53740
g53485 and n53552_not n53740 ; n53741
g53486 and n53739_not n53741_not ; n53742
g53487 and b[39]_not n53742_not ; n53743
g53488 and n52935_not n53429 ; n53744
g53489 and n53425_not n53744 ; n53745
g53490 and n53426_not n53429_not ; n53746
g53491 and n53745_not n53746_not ; n53747
g53492 and n53554_not n53747_not ; n53748
g53493 and n52925_not n53553_not ; n53749
g53494 and n53552_not n53749 ; n53750
g53495 and n53748_not n53750_not ; n53751
g53496 and b[38]_not n53751_not ; n53752
g53497 and n52944_not n53424 ; n53753
g53498 and n53420_not n53753 ; n53754
g53499 and n53421_not n53424_not ; n53755
g53500 and n53754_not n53755_not ; n53756
g53501 and n53554_not n53756_not ; n53757
g53502 and n52934_not n53553_not ; n53758
g53503 and n53552_not n53758 ; n53759
g53504 and n53757_not n53759_not ; n53760
g53505 and b[37]_not n53760_not ; n53761
g53506 and n52953_not n53419 ; n53762
g53507 and n53415_not n53762 ; n53763
g53508 and n53416_not n53419_not ; n53764
g53509 and n53763_not n53764_not ; n53765
g53510 and n53554_not n53765_not ; n53766
g53511 and n52943_not n53553_not ; n53767
g53512 and n53552_not n53767 ; n53768
g53513 and n53766_not n53768_not ; n53769
g53514 and b[36]_not n53769_not ; n53770
g53515 and n52962_not n53414 ; n53771
g53516 and n53410_not n53771 ; n53772
g53517 and n53411_not n53414_not ; n53773
g53518 and n53772_not n53773_not ; n53774
g53519 and n53554_not n53774_not ; n53775
g53520 and n52952_not n53553_not ; n53776
g53521 and n53552_not n53776 ; n53777
g53522 and n53775_not n53777_not ; n53778
g53523 and b[35]_not n53778_not ; n53779
g53524 and n52971_not n53409 ; n53780
g53525 and n53405_not n53780 ; n53781
g53526 and n53406_not n53409_not ; n53782
g53527 and n53781_not n53782_not ; n53783
g53528 and n53554_not n53783_not ; n53784
g53529 and n52961_not n53553_not ; n53785
g53530 and n53552_not n53785 ; n53786
g53531 and n53784_not n53786_not ; n53787
g53532 and b[34]_not n53787_not ; n53788
g53533 and n52980_not n53404 ; n53789
g53534 and n53400_not n53789 ; n53790
g53535 and n53401_not n53404_not ; n53791
g53536 and n53790_not n53791_not ; n53792
g53537 and n53554_not n53792_not ; n53793
g53538 and n52970_not n53553_not ; n53794
g53539 and n53552_not n53794 ; n53795
g53540 and n53793_not n53795_not ; n53796
g53541 and b[33]_not n53796_not ; n53797
g53542 and n52989_not n53399 ; n53798
g53543 and n53395_not n53798 ; n53799
g53544 and n53396_not n53399_not ; n53800
g53545 and n53799_not n53800_not ; n53801
g53546 and n53554_not n53801_not ; n53802
g53547 and n52979_not n53553_not ; n53803
g53548 and n53552_not n53803 ; n53804
g53549 and n53802_not n53804_not ; n53805
g53550 and b[32]_not n53805_not ; n53806
g53551 and n52998_not n53394 ; n53807
g53552 and n53390_not n53807 ; n53808
g53553 and n53391_not n53394_not ; n53809
g53554 and n53808_not n53809_not ; n53810
g53555 and n53554_not n53810_not ; n53811
g53556 and n52988_not n53553_not ; n53812
g53557 and n53552_not n53812 ; n53813
g53558 and n53811_not n53813_not ; n53814
g53559 and b[31]_not n53814_not ; n53815
g53560 and n53007_not n53389 ; n53816
g53561 and n53385_not n53816 ; n53817
g53562 and n53386_not n53389_not ; n53818
g53563 and n53817_not n53818_not ; n53819
g53564 and n53554_not n53819_not ; n53820
g53565 and n52997_not n53553_not ; n53821
g53566 and n53552_not n53821 ; n53822
g53567 and n53820_not n53822_not ; n53823
g53568 and b[30]_not n53823_not ; n53824
g53569 and n53016_not n53384 ; n53825
g53570 and n53380_not n53825 ; n53826
g53571 and n53381_not n53384_not ; n53827
g53572 and n53826_not n53827_not ; n53828
g53573 and n53554_not n53828_not ; n53829
g53574 and n53006_not n53553_not ; n53830
g53575 and n53552_not n53830 ; n53831
g53576 and n53829_not n53831_not ; n53832
g53577 and b[29]_not n53832_not ; n53833
g53578 and n53025_not n53379 ; n53834
g53579 and n53375_not n53834 ; n53835
g53580 and n53376_not n53379_not ; n53836
g53581 and n53835_not n53836_not ; n53837
g53582 and n53554_not n53837_not ; n53838
g53583 and n53015_not n53553_not ; n53839
g53584 and n53552_not n53839 ; n53840
g53585 and n53838_not n53840_not ; n53841
g53586 and b[28]_not n53841_not ; n53842
g53587 and n53034_not n53374 ; n53843
g53588 and n53370_not n53843 ; n53844
g53589 and n53371_not n53374_not ; n53845
g53590 and n53844_not n53845_not ; n53846
g53591 and n53554_not n53846_not ; n53847
g53592 and n53024_not n53553_not ; n53848
g53593 and n53552_not n53848 ; n53849
g53594 and n53847_not n53849_not ; n53850
g53595 and b[27]_not n53850_not ; n53851
g53596 and n53043_not n53369 ; n53852
g53597 and n53365_not n53852 ; n53853
g53598 and n53366_not n53369_not ; n53854
g53599 and n53853_not n53854_not ; n53855
g53600 and n53554_not n53855_not ; n53856
g53601 and n53033_not n53553_not ; n53857
g53602 and n53552_not n53857 ; n53858
g53603 and n53856_not n53858_not ; n53859
g53604 and b[26]_not n53859_not ; n53860
g53605 and n53052_not n53364 ; n53861
g53606 and n53360_not n53861 ; n53862
g53607 and n53361_not n53364_not ; n53863
g53608 and n53862_not n53863_not ; n53864
g53609 and n53554_not n53864_not ; n53865
g53610 and n53042_not n53553_not ; n53866
g53611 and n53552_not n53866 ; n53867
g53612 and n53865_not n53867_not ; n53868
g53613 and b[25]_not n53868_not ; n53869
g53614 and n53061_not n53359 ; n53870
g53615 and n53355_not n53870 ; n53871
g53616 and n53356_not n53359_not ; n53872
g53617 and n53871_not n53872_not ; n53873
g53618 and n53554_not n53873_not ; n53874
g53619 and n53051_not n53553_not ; n53875
g53620 and n53552_not n53875 ; n53876
g53621 and n53874_not n53876_not ; n53877
g53622 and b[24]_not n53877_not ; n53878
g53623 and n53070_not n53354 ; n53879
g53624 and n53350_not n53879 ; n53880
g53625 and n53351_not n53354_not ; n53881
g53626 and n53880_not n53881_not ; n53882
g53627 and n53554_not n53882_not ; n53883
g53628 and n53060_not n53553_not ; n53884
g53629 and n53552_not n53884 ; n53885
g53630 and n53883_not n53885_not ; n53886
g53631 and b[23]_not n53886_not ; n53887
g53632 and n53079_not n53349 ; n53888
g53633 and n53345_not n53888 ; n53889
g53634 and n53346_not n53349_not ; n53890
g53635 and n53889_not n53890_not ; n53891
g53636 and n53554_not n53891_not ; n53892
g53637 and n53069_not n53553_not ; n53893
g53638 and n53552_not n53893 ; n53894
g53639 and n53892_not n53894_not ; n53895
g53640 and b[22]_not n53895_not ; n53896
g53641 and n53088_not n53344 ; n53897
g53642 and n53340_not n53897 ; n53898
g53643 and n53341_not n53344_not ; n53899
g53644 and n53898_not n53899_not ; n53900
g53645 and n53554_not n53900_not ; n53901
g53646 and n53078_not n53553_not ; n53902
g53647 and n53552_not n53902 ; n53903
g53648 and n53901_not n53903_not ; n53904
g53649 and b[21]_not n53904_not ; n53905
g53650 and n53097_not n53339 ; n53906
g53651 and n53335_not n53906 ; n53907
g53652 and n53336_not n53339_not ; n53908
g53653 and n53907_not n53908_not ; n53909
g53654 and n53554_not n53909_not ; n53910
g53655 and n53087_not n53553_not ; n53911
g53656 and n53552_not n53911 ; n53912
g53657 and n53910_not n53912_not ; n53913
g53658 and b[20]_not n53913_not ; n53914
g53659 and n53106_not n53334 ; n53915
g53660 and n53330_not n53915 ; n53916
g53661 and n53331_not n53334_not ; n53917
g53662 and n53916_not n53917_not ; n53918
g53663 and n53554_not n53918_not ; n53919
g53664 and n53096_not n53553_not ; n53920
g53665 and n53552_not n53920 ; n53921
g53666 and n53919_not n53921_not ; n53922
g53667 and b[19]_not n53922_not ; n53923
g53668 and n53115_not n53329 ; n53924
g53669 and n53325_not n53924 ; n53925
g53670 and n53326_not n53329_not ; n53926
g53671 and n53925_not n53926_not ; n53927
g53672 and n53554_not n53927_not ; n53928
g53673 and n53105_not n53553_not ; n53929
g53674 and n53552_not n53929 ; n53930
g53675 and n53928_not n53930_not ; n53931
g53676 and b[18]_not n53931_not ; n53932
g53677 and n53124_not n53324 ; n53933
g53678 and n53320_not n53933 ; n53934
g53679 and n53321_not n53324_not ; n53935
g53680 and n53934_not n53935_not ; n53936
g53681 and n53554_not n53936_not ; n53937
g53682 and n53114_not n53553_not ; n53938
g53683 and n53552_not n53938 ; n53939
g53684 and n53937_not n53939_not ; n53940
g53685 and b[17]_not n53940_not ; n53941
g53686 and n53133_not n53319 ; n53942
g53687 and n53315_not n53942 ; n53943
g53688 and n53316_not n53319_not ; n53944
g53689 and n53943_not n53944_not ; n53945
g53690 and n53554_not n53945_not ; n53946
g53691 and n53123_not n53553_not ; n53947
g53692 and n53552_not n53947 ; n53948
g53693 and n53946_not n53948_not ; n53949
g53694 and b[16]_not n53949_not ; n53950
g53695 and n53142_not n53314 ; n53951
g53696 and n53310_not n53951 ; n53952
g53697 and n53311_not n53314_not ; n53953
g53698 and n53952_not n53953_not ; n53954
g53699 and n53554_not n53954_not ; n53955
g53700 and n53132_not n53553_not ; n53956
g53701 and n53552_not n53956 ; n53957
g53702 and n53955_not n53957_not ; n53958
g53703 and b[15]_not n53958_not ; n53959
g53704 and n53151_not n53309 ; n53960
g53705 and n53305_not n53960 ; n53961
g53706 and n53306_not n53309_not ; n53962
g53707 and n53961_not n53962_not ; n53963
g53708 and n53554_not n53963_not ; n53964
g53709 and n53141_not n53553_not ; n53965
g53710 and n53552_not n53965 ; n53966
g53711 and n53964_not n53966_not ; n53967
g53712 and b[14]_not n53967_not ; n53968
g53713 and n53160_not n53304 ; n53969
g53714 and n53300_not n53969 ; n53970
g53715 and n53301_not n53304_not ; n53971
g53716 and n53970_not n53971_not ; n53972
g53717 and n53554_not n53972_not ; n53973
g53718 and n53150_not n53553_not ; n53974
g53719 and n53552_not n53974 ; n53975
g53720 and n53973_not n53975_not ; n53976
g53721 and b[13]_not n53976_not ; n53977
g53722 and n53169_not n53299 ; n53978
g53723 and n53295_not n53978 ; n53979
g53724 and n53296_not n53299_not ; n53980
g53725 and n53979_not n53980_not ; n53981
g53726 and n53554_not n53981_not ; n53982
g53727 and n53159_not n53553_not ; n53983
g53728 and n53552_not n53983 ; n53984
g53729 and n53982_not n53984_not ; n53985
g53730 and b[12]_not n53985_not ; n53986
g53731 and n53178_not n53294 ; n53987
g53732 and n53290_not n53987 ; n53988
g53733 and n53291_not n53294_not ; n53989
g53734 and n53988_not n53989_not ; n53990
g53735 and n53554_not n53990_not ; n53991
g53736 and n53168_not n53553_not ; n53992
g53737 and n53552_not n53992 ; n53993
g53738 and n53991_not n53993_not ; n53994
g53739 and b[11]_not n53994_not ; n53995
g53740 and n53187_not n53289 ; n53996
g53741 and n53285_not n53996 ; n53997
g53742 and n53286_not n53289_not ; n53998
g53743 and n53997_not n53998_not ; n53999
g53744 and n53554_not n53999_not ; n54000
g53745 and n53177_not n53553_not ; n54001
g53746 and n53552_not n54001 ; n54002
g53747 and n54000_not n54002_not ; n54003
g53748 and b[10]_not n54003_not ; n54004
g53749 and n53196_not n53284 ; n54005
g53750 and n53280_not n54005 ; n54006
g53751 and n53281_not n53284_not ; n54007
g53752 and n54006_not n54007_not ; n54008
g53753 and n53554_not n54008_not ; n54009
g53754 and n53186_not n53553_not ; n54010
g53755 and n53552_not n54010 ; n54011
g53756 and n54009_not n54011_not ; n54012
g53757 and b[9]_not n54012_not ; n54013
g53758 and n53205_not n53279 ; n54014
g53759 and n53275_not n54014 ; n54015
g53760 and n53276_not n53279_not ; n54016
g53761 and n54015_not n54016_not ; n54017
g53762 and n53554_not n54017_not ; n54018
g53763 and n53195_not n53553_not ; n54019
g53764 and n53552_not n54019 ; n54020
g53765 and n54018_not n54020_not ; n54021
g53766 and b[8]_not n54021_not ; n54022
g53767 and n53214_not n53274 ; n54023
g53768 and n53270_not n54023 ; n54024
g53769 and n53271_not n53274_not ; n54025
g53770 and n54024_not n54025_not ; n54026
g53771 and n53554_not n54026_not ; n54027
g53772 and n53204_not n53553_not ; n54028
g53773 and n53552_not n54028 ; n54029
g53774 and n54027_not n54029_not ; n54030
g53775 and b[7]_not n54030_not ; n54031
g53776 and n53223_not n53269 ; n54032
g53777 and n53265_not n54032 ; n54033
g53778 and n53266_not n53269_not ; n54034
g53779 and n54033_not n54034_not ; n54035
g53780 and n53554_not n54035_not ; n54036
g53781 and n53213_not n53553_not ; n54037
g53782 and n53552_not n54037 ; n54038
g53783 and n54036_not n54038_not ; n54039
g53784 and b[6]_not n54039_not ; n54040
g53785 and n53232_not n53264 ; n54041
g53786 and n53260_not n54041 ; n54042
g53787 and n53261_not n53264_not ; n54043
g53788 and n54042_not n54043_not ; n54044
g53789 and n53554_not n54044_not ; n54045
g53790 and n53222_not n53553_not ; n54046
g53791 and n53552_not n54046 ; n54047
g53792 and n54045_not n54047_not ; n54048
g53793 and b[5]_not n54048_not ; n54049
g53794 and n53240_not n53259 ; n54050
g53795 and n53255_not n54050 ; n54051
g53796 and n53256_not n53259_not ; n54052
g53797 and n54051_not n54052_not ; n54053
g53798 and n53554_not n54053_not ; n54054
g53799 and n53231_not n53553_not ; n54055
g53800 and n53552_not n54055 ; n54056
g53801 and n54054_not n54056_not ; n54057
g53802 and b[4]_not n54057_not ; n54058
g53803 and n53250_not n53254 ; n54059
g53804 and n53249_not n54059 ; n54060
g53805 and n53251_not n53254_not ; n54061
g53806 and n54060_not n54061_not ; n54062
g53807 and n53554_not n54062_not ; n54063
g53808 and n53239_not n53553_not ; n54064
g53809 and n53552_not n54064 ; n54065
g53810 and n54063_not n54065_not ; n54066
g53811 and b[3]_not n54066_not ; n54067
g53812 and n25233 n53247_not ; n54068
g53813 and n53245_not n54068 ; n54069
g53814 and n53249_not n54069_not ; n54070
g53815 and n53554_not n54070 ; n54071
g53816 and n53244_not n53553_not ; n54072
g53817 and n53552_not n54072 ; n54073
g53818 and n54071_not n54073_not ; n54074
g53819 and b[2]_not n54074_not ; n54075
g53820 and b[0] n53554_not ; n54076
g53821 and a[4] n54076_not ; n54077
g53822 and n25233 n53554_not ; n54078
g53823 and n54077_not n54078_not ; n54079
g53824 and b[1] n54079_not ; n54080
g53825 and b[1]_not n54078_not ; n54081
g53826 and n54077_not n54081 ; n54082
g53827 and n54080_not n54082_not ; n54083
g53828 and n26069_not n54083_not ; n54084
g53829 and b[1]_not n54079_not ; n54085
g53830 and n54084_not n54085_not ; n54086
g53831 and b[2] n54073_not ; n54087
g53832 and n54071_not n54087 ; n54088
g53833 and n54075_not n54088_not ; n54089
g53834 and n54086_not n54089 ; n54090
g53835 and n54075_not n54090_not ; n54091
g53836 and b[3] n54065_not ; n54092
g53837 and n54063_not n54092 ; n54093
g53838 and n54067_not n54093_not ; n54094
g53839 and n54091_not n54094 ; n54095
g53840 and n54067_not n54095_not ; n54096
g53841 and b[4] n54056_not ; n54097
g53842 and n54054_not n54097 ; n54098
g53843 and n54058_not n54098_not ; n54099
g53844 and n54096_not n54099 ; n54100
g53845 and n54058_not n54100_not ; n54101
g53846 and b[5] n54047_not ; n54102
g53847 and n54045_not n54102 ; n54103
g53848 and n54049_not n54103_not ; n54104
g53849 and n54101_not n54104 ; n54105
g53850 and n54049_not n54105_not ; n54106
g53851 and b[6] n54038_not ; n54107
g53852 and n54036_not n54107 ; n54108
g53853 and n54040_not n54108_not ; n54109
g53854 and n54106_not n54109 ; n54110
g53855 and n54040_not n54110_not ; n54111
g53856 and b[7] n54029_not ; n54112
g53857 and n54027_not n54112 ; n54113
g53858 and n54031_not n54113_not ; n54114
g53859 and n54111_not n54114 ; n54115
g53860 and n54031_not n54115_not ; n54116
g53861 and b[8] n54020_not ; n54117
g53862 and n54018_not n54117 ; n54118
g53863 and n54022_not n54118_not ; n54119
g53864 and n54116_not n54119 ; n54120
g53865 and n54022_not n54120_not ; n54121
g53866 and b[9] n54011_not ; n54122
g53867 and n54009_not n54122 ; n54123
g53868 and n54013_not n54123_not ; n54124
g53869 and n54121_not n54124 ; n54125
g53870 and n54013_not n54125_not ; n54126
g53871 and b[10] n54002_not ; n54127
g53872 and n54000_not n54127 ; n54128
g53873 and n54004_not n54128_not ; n54129
g53874 and n54126_not n54129 ; n54130
g53875 and n54004_not n54130_not ; n54131
g53876 and b[11] n53993_not ; n54132
g53877 and n53991_not n54132 ; n54133
g53878 and n53995_not n54133_not ; n54134
g53879 and n54131_not n54134 ; n54135
g53880 and n53995_not n54135_not ; n54136
g53881 and b[12] n53984_not ; n54137
g53882 and n53982_not n54137 ; n54138
g53883 and n53986_not n54138_not ; n54139
g53884 and n54136_not n54139 ; n54140
g53885 and n53986_not n54140_not ; n54141
g53886 and b[13] n53975_not ; n54142
g53887 and n53973_not n54142 ; n54143
g53888 and n53977_not n54143_not ; n54144
g53889 and n54141_not n54144 ; n54145
g53890 and n53977_not n54145_not ; n54146
g53891 and b[14] n53966_not ; n54147
g53892 and n53964_not n54147 ; n54148
g53893 and n53968_not n54148_not ; n54149
g53894 and n54146_not n54149 ; n54150
g53895 and n53968_not n54150_not ; n54151
g53896 and b[15] n53957_not ; n54152
g53897 and n53955_not n54152 ; n54153
g53898 and n53959_not n54153_not ; n54154
g53899 and n54151_not n54154 ; n54155
g53900 and n53959_not n54155_not ; n54156
g53901 and b[16] n53948_not ; n54157
g53902 and n53946_not n54157 ; n54158
g53903 and n53950_not n54158_not ; n54159
g53904 and n54156_not n54159 ; n54160
g53905 and n53950_not n54160_not ; n54161
g53906 and b[17] n53939_not ; n54162
g53907 and n53937_not n54162 ; n54163
g53908 and n53941_not n54163_not ; n54164
g53909 and n54161_not n54164 ; n54165
g53910 and n53941_not n54165_not ; n54166
g53911 and b[18] n53930_not ; n54167
g53912 and n53928_not n54167 ; n54168
g53913 and n53932_not n54168_not ; n54169
g53914 and n54166_not n54169 ; n54170
g53915 and n53932_not n54170_not ; n54171
g53916 and b[19] n53921_not ; n54172
g53917 and n53919_not n54172 ; n54173
g53918 and n53923_not n54173_not ; n54174
g53919 and n54171_not n54174 ; n54175
g53920 and n53923_not n54175_not ; n54176
g53921 and b[20] n53912_not ; n54177
g53922 and n53910_not n54177 ; n54178
g53923 and n53914_not n54178_not ; n54179
g53924 and n54176_not n54179 ; n54180
g53925 and n53914_not n54180_not ; n54181
g53926 and b[21] n53903_not ; n54182
g53927 and n53901_not n54182 ; n54183
g53928 and n53905_not n54183_not ; n54184
g53929 and n54181_not n54184 ; n54185
g53930 and n53905_not n54185_not ; n54186
g53931 and b[22] n53894_not ; n54187
g53932 and n53892_not n54187 ; n54188
g53933 and n53896_not n54188_not ; n54189
g53934 and n54186_not n54189 ; n54190
g53935 and n53896_not n54190_not ; n54191
g53936 and b[23] n53885_not ; n54192
g53937 and n53883_not n54192 ; n54193
g53938 and n53887_not n54193_not ; n54194
g53939 and n54191_not n54194 ; n54195
g53940 and n53887_not n54195_not ; n54196
g53941 and b[24] n53876_not ; n54197
g53942 and n53874_not n54197 ; n54198
g53943 and n53878_not n54198_not ; n54199
g53944 and n54196_not n54199 ; n54200
g53945 and n53878_not n54200_not ; n54201
g53946 and b[25] n53867_not ; n54202
g53947 and n53865_not n54202 ; n54203
g53948 and n53869_not n54203_not ; n54204
g53949 and n54201_not n54204 ; n54205
g53950 and n53869_not n54205_not ; n54206
g53951 and b[26] n53858_not ; n54207
g53952 and n53856_not n54207 ; n54208
g53953 and n53860_not n54208_not ; n54209
g53954 and n54206_not n54209 ; n54210
g53955 and n53860_not n54210_not ; n54211
g53956 and b[27] n53849_not ; n54212
g53957 and n53847_not n54212 ; n54213
g53958 and n53851_not n54213_not ; n54214
g53959 and n54211_not n54214 ; n54215
g53960 and n53851_not n54215_not ; n54216
g53961 and b[28] n53840_not ; n54217
g53962 and n53838_not n54217 ; n54218
g53963 and n53842_not n54218_not ; n54219
g53964 and n54216_not n54219 ; n54220
g53965 and n53842_not n54220_not ; n54221
g53966 and b[29] n53831_not ; n54222
g53967 and n53829_not n54222 ; n54223
g53968 and n53833_not n54223_not ; n54224
g53969 and n54221_not n54224 ; n54225
g53970 and n53833_not n54225_not ; n54226
g53971 and b[30] n53822_not ; n54227
g53972 and n53820_not n54227 ; n54228
g53973 and n53824_not n54228_not ; n54229
g53974 and n54226_not n54229 ; n54230
g53975 and n53824_not n54230_not ; n54231
g53976 and b[31] n53813_not ; n54232
g53977 and n53811_not n54232 ; n54233
g53978 and n53815_not n54233_not ; n54234
g53979 and n54231_not n54234 ; n54235
g53980 and n53815_not n54235_not ; n54236
g53981 and b[32] n53804_not ; n54237
g53982 and n53802_not n54237 ; n54238
g53983 and n53806_not n54238_not ; n54239
g53984 and n54236_not n54239 ; n54240
g53985 and n53806_not n54240_not ; n54241
g53986 and b[33] n53795_not ; n54242
g53987 and n53793_not n54242 ; n54243
g53988 and n53797_not n54243_not ; n54244
g53989 and n54241_not n54244 ; n54245
g53990 and n53797_not n54245_not ; n54246
g53991 and b[34] n53786_not ; n54247
g53992 and n53784_not n54247 ; n54248
g53993 and n53788_not n54248_not ; n54249
g53994 and n54246_not n54249 ; n54250
g53995 and n53788_not n54250_not ; n54251
g53996 and b[35] n53777_not ; n54252
g53997 and n53775_not n54252 ; n54253
g53998 and n53779_not n54253_not ; n54254
g53999 and n54251_not n54254 ; n54255
g54000 and n53779_not n54255_not ; n54256
g54001 and b[36] n53768_not ; n54257
g54002 and n53766_not n54257 ; n54258
g54003 and n53770_not n54258_not ; n54259
g54004 and n54256_not n54259 ; n54260
g54005 and n53770_not n54260_not ; n54261
g54006 and b[37] n53759_not ; n54262
g54007 and n53757_not n54262 ; n54263
g54008 and n53761_not n54263_not ; n54264
g54009 and n54261_not n54264 ; n54265
g54010 and n53761_not n54265_not ; n54266
g54011 and b[38] n53750_not ; n54267
g54012 and n53748_not n54267 ; n54268
g54013 and n53752_not n54268_not ; n54269
g54014 and n54266_not n54269 ; n54270
g54015 and n53752_not n54270_not ; n54271
g54016 and b[39] n53741_not ; n54272
g54017 and n53739_not n54272 ; n54273
g54018 and n53743_not n54273_not ; n54274
g54019 and n54271_not n54274 ; n54275
g54020 and n53743_not n54275_not ; n54276
g54021 and b[40] n53732_not ; n54277
g54022 and n53730_not n54277 ; n54278
g54023 and n53734_not n54278_not ; n54279
g54024 and n54276_not n54279 ; n54280
g54025 and n53734_not n54280_not ; n54281
g54026 and b[41] n53723_not ; n54282
g54027 and n53721_not n54282 ; n54283
g54028 and n53725_not n54283_not ; n54284
g54029 and n54281_not n54284 ; n54285
g54030 and n53725_not n54285_not ; n54286
g54031 and b[42] n53714_not ; n54287
g54032 and n53712_not n54287 ; n54288
g54033 and n53716_not n54288_not ; n54289
g54034 and n54286_not n54289 ; n54290
g54035 and n53716_not n54290_not ; n54291
g54036 and b[43] n53705_not ; n54292
g54037 and n53703_not n54292 ; n54293
g54038 and n53707_not n54293_not ; n54294
g54039 and n54291_not n54294 ; n54295
g54040 and n53707_not n54295_not ; n54296
g54041 and b[44] n53696_not ; n54297
g54042 and n53694_not n54297 ; n54298
g54043 and n53698_not n54298_not ; n54299
g54044 and n54296_not n54299 ; n54300
g54045 and n53698_not n54300_not ; n54301
g54046 and b[45] n53687_not ; n54302
g54047 and n53685_not n54302 ; n54303
g54048 and n53689_not n54303_not ; n54304
g54049 and n54301_not n54304 ; n54305
g54050 and n53689_not n54305_not ; n54306
g54051 and b[46] n53678_not ; n54307
g54052 and n53676_not n54307 ; n54308
g54053 and n53680_not n54308_not ; n54309
g54054 and n54306_not n54309 ; n54310
g54055 and n53680_not n54310_not ; n54311
g54056 and b[47] n53669_not ; n54312
g54057 and n53667_not n54312 ; n54313
g54058 and n53671_not n54313_not ; n54314
g54059 and n54311_not n54314 ; n54315
g54060 and n53671_not n54315_not ; n54316
g54061 and b[48] n53660_not ; n54317
g54062 and n53658_not n54317 ; n54318
g54063 and n53662_not n54318_not ; n54319
g54064 and n54316_not n54319 ; n54320
g54065 and n53662_not n54320_not ; n54321
g54066 and b[49] n53651_not ; n54322
g54067 and n53649_not n54322 ; n54323
g54068 and n53653_not n54323_not ; n54324
g54069 and n54321_not n54324 ; n54325
g54070 and n53653_not n54325_not ; n54326
g54071 and b[50] n53642_not ; n54327
g54072 and n53640_not n54327 ; n54328
g54073 and n53644_not n54328_not ; n54329
g54074 and n54326_not n54329 ; n54330
g54075 and n53644_not n54330_not ; n54331
g54076 and b[51] n53633_not ; n54332
g54077 and n53631_not n54332 ; n54333
g54078 and n53635_not n54333_not ; n54334
g54079 and n54331_not n54334 ; n54335
g54080 and n53635_not n54335_not ; n54336
g54081 and b[52] n53624_not ; n54337
g54082 and n53622_not n54337 ; n54338
g54083 and n53626_not n54338_not ; n54339
g54084 and n54336_not n54339 ; n54340
g54085 and n53626_not n54340_not ; n54341
g54086 and b[53] n53615_not ; n54342
g54087 and n53613_not n54342 ; n54343
g54088 and n53617_not n54343_not ; n54344
g54089 and n54341_not n54344 ; n54345
g54090 and n53617_not n54345_not ; n54346
g54091 and b[54] n53606_not ; n54347
g54092 and n53604_not n54347 ; n54348
g54093 and n53608_not n54348_not ; n54349
g54094 and n54346_not n54349 ; n54350
g54095 and n53608_not n54350_not ; n54351
g54096 and b[55] n53597_not ; n54352
g54097 and n53595_not n54352 ; n54353
g54098 and n53599_not n54353_not ; n54354
g54099 and n54351_not n54354 ; n54355
g54100 and n53599_not n54355_not ; n54356
g54101 and b[56] n53588_not ; n54357
g54102 and n53586_not n54357 ; n54358
g54103 and n53590_not n54358_not ; n54359
g54104 and n54356_not n54359 ; n54360
g54105 and n53590_not n54360_not ; n54361
g54106 and b[57] n53579_not ; n54362
g54107 and n53577_not n54362 ; n54363
g54108 and n53581_not n54363_not ; n54364
g54109 and n54361_not n54364 ; n54365
g54110 and n53581_not n54365_not ; n54366
g54111 and b[58] n53570_not ; n54367
g54112 and n53568_not n54367 ; n54368
g54113 and n53572_not n54368_not ; n54369
g54114 and n54366_not n54369 ; n54370
g54115 and n53572_not n54370_not ; n54371
g54116 and b[59] n53561_not ; n54372
g54117 and n53559_not n54372 ; n54373
g54118 and n53563_not n54373_not ; n54374
g54119 and n54371_not n54374 ; n54375
g54120 and n53563_not n54375_not ; n54376
g54121 and n52737_not n53549_not ; n54377
g54122 and n53547_not n54377 ; n54378
g54123 and n53535_not n54378 ; n54379
g54124 and n53547_not n53549_not ; n54380
g54125 and n53536_not n54380_not ; n54381
g54126 and n54379_not n54381_not ; n54382
g54127 and n53554_not n54382_not ; n54383
g54128 and n53546_not n53553_not ; n54384
g54129 and n53552_not n54384 ; n54385
g54130 and n54383_not n54385_not ; n54386
g54131 and b[60]_not n54386_not ; n54387
g54132 and b[60] n54385_not ; n54388
g54133 and n54383_not n54388 ; n54389
g54134 and n403 n54389_not ; n54390
g54135 and n54387_not n54390 ; n54391
g54136 and n54376_not n54391 ; n54392
g54137 and n280 n54386_not ; n54393
g54138 and n54392_not n54393_not ; n54394
g54139 and n53572_not n54374 ; n54395
g54140 and n54370_not n54395 ; n54396
g54141 and n54371_not n54374_not ; n54397
g54142 and n54396_not n54397_not ; n54398
g54143 and n54394_not n54398_not ; n54399
g54144 and n53562_not n54393_not ; n54400
g54145 and n54392_not n54400 ; n54401
g54146 and n54399_not n54401_not ; n54402
g54147 and b[60]_not n54402_not ; n54403
g54148 and n53581_not n54369 ; n54404
g54149 and n54365_not n54404 ; n54405
g54150 and n54366_not n54369_not ; n54406
g54151 and n54405_not n54406_not ; n54407
g54152 and n54394_not n54407_not ; n54408
g54153 and n53571_not n54393_not ; n54409
g54154 and n54392_not n54409 ; n54410
g54155 and n54408_not n54410_not ; n54411
g54156 and b[59]_not n54411_not ; n54412
g54157 and n53590_not n54364 ; n54413
g54158 and n54360_not n54413 ; n54414
g54159 and n54361_not n54364_not ; n54415
g54160 and n54414_not n54415_not ; n54416
g54161 and n54394_not n54416_not ; n54417
g54162 and n53580_not n54393_not ; n54418
g54163 and n54392_not n54418 ; n54419
g54164 and n54417_not n54419_not ; n54420
g54165 and b[58]_not n54420_not ; n54421
g54166 and n53599_not n54359 ; n54422
g54167 and n54355_not n54422 ; n54423
g54168 and n54356_not n54359_not ; n54424
g54169 and n54423_not n54424_not ; n54425
g54170 and n54394_not n54425_not ; n54426
g54171 and n53589_not n54393_not ; n54427
g54172 and n54392_not n54427 ; n54428
g54173 and n54426_not n54428_not ; n54429
g54174 and b[57]_not n54429_not ; n54430
g54175 and n53608_not n54354 ; n54431
g54176 and n54350_not n54431 ; n54432
g54177 and n54351_not n54354_not ; n54433
g54178 and n54432_not n54433_not ; n54434
g54179 and n54394_not n54434_not ; n54435
g54180 and n53598_not n54393_not ; n54436
g54181 and n54392_not n54436 ; n54437
g54182 and n54435_not n54437_not ; n54438
g54183 and b[56]_not n54438_not ; n54439
g54184 and n53617_not n54349 ; n54440
g54185 and n54345_not n54440 ; n54441
g54186 and n54346_not n54349_not ; n54442
g54187 and n54441_not n54442_not ; n54443
g54188 and n54394_not n54443_not ; n54444
g54189 and n53607_not n54393_not ; n54445
g54190 and n54392_not n54445 ; n54446
g54191 and n54444_not n54446_not ; n54447
g54192 and b[55]_not n54447_not ; n54448
g54193 and n53626_not n54344 ; n54449
g54194 and n54340_not n54449 ; n54450
g54195 and n54341_not n54344_not ; n54451
g54196 and n54450_not n54451_not ; n54452
g54197 and n54394_not n54452_not ; n54453
g54198 and n53616_not n54393_not ; n54454
g54199 and n54392_not n54454 ; n54455
g54200 and n54453_not n54455_not ; n54456
g54201 and b[54]_not n54456_not ; n54457
g54202 and n53635_not n54339 ; n54458
g54203 and n54335_not n54458 ; n54459
g54204 and n54336_not n54339_not ; n54460
g54205 and n54459_not n54460_not ; n54461
g54206 and n54394_not n54461_not ; n54462
g54207 and n53625_not n54393_not ; n54463
g54208 and n54392_not n54463 ; n54464
g54209 and n54462_not n54464_not ; n54465
g54210 and b[53]_not n54465_not ; n54466
g54211 and n53644_not n54334 ; n54467
g54212 and n54330_not n54467 ; n54468
g54213 and n54331_not n54334_not ; n54469
g54214 and n54468_not n54469_not ; n54470
g54215 and n54394_not n54470_not ; n54471
g54216 and n53634_not n54393_not ; n54472
g54217 and n54392_not n54472 ; n54473
g54218 and n54471_not n54473_not ; n54474
g54219 and b[52]_not n54474_not ; n54475
g54220 and n53653_not n54329 ; n54476
g54221 and n54325_not n54476 ; n54477
g54222 and n54326_not n54329_not ; n54478
g54223 and n54477_not n54478_not ; n54479
g54224 and n54394_not n54479_not ; n54480
g54225 and n53643_not n54393_not ; n54481
g54226 and n54392_not n54481 ; n54482
g54227 and n54480_not n54482_not ; n54483
g54228 and b[51]_not n54483_not ; n54484
g54229 and n53662_not n54324 ; n54485
g54230 and n54320_not n54485 ; n54486
g54231 and n54321_not n54324_not ; n54487
g54232 and n54486_not n54487_not ; n54488
g54233 and n54394_not n54488_not ; n54489
g54234 and n53652_not n54393_not ; n54490
g54235 and n54392_not n54490 ; n54491
g54236 and n54489_not n54491_not ; n54492
g54237 and b[50]_not n54492_not ; n54493
g54238 and n53671_not n54319 ; n54494
g54239 and n54315_not n54494 ; n54495
g54240 and n54316_not n54319_not ; n54496
g54241 and n54495_not n54496_not ; n54497
g54242 and n54394_not n54497_not ; n54498
g54243 and n53661_not n54393_not ; n54499
g54244 and n54392_not n54499 ; n54500
g54245 and n54498_not n54500_not ; n54501
g54246 and b[49]_not n54501_not ; n54502
g54247 and n53680_not n54314 ; n54503
g54248 and n54310_not n54503 ; n54504
g54249 and n54311_not n54314_not ; n54505
g54250 and n54504_not n54505_not ; n54506
g54251 and n54394_not n54506_not ; n54507
g54252 and n53670_not n54393_not ; n54508
g54253 and n54392_not n54508 ; n54509
g54254 and n54507_not n54509_not ; n54510
g54255 and b[48]_not n54510_not ; n54511
g54256 and n53689_not n54309 ; n54512
g54257 and n54305_not n54512 ; n54513
g54258 and n54306_not n54309_not ; n54514
g54259 and n54513_not n54514_not ; n54515
g54260 and n54394_not n54515_not ; n54516
g54261 and n53679_not n54393_not ; n54517
g54262 and n54392_not n54517 ; n54518
g54263 and n54516_not n54518_not ; n54519
g54264 and b[47]_not n54519_not ; n54520
g54265 and n53698_not n54304 ; n54521
g54266 and n54300_not n54521 ; n54522
g54267 and n54301_not n54304_not ; n54523
g54268 and n54522_not n54523_not ; n54524
g54269 and n54394_not n54524_not ; n54525
g54270 and n53688_not n54393_not ; n54526
g54271 and n54392_not n54526 ; n54527
g54272 and n54525_not n54527_not ; n54528
g54273 and b[46]_not n54528_not ; n54529
g54274 and n53707_not n54299 ; n54530
g54275 and n54295_not n54530 ; n54531
g54276 and n54296_not n54299_not ; n54532
g54277 and n54531_not n54532_not ; n54533
g54278 and n54394_not n54533_not ; n54534
g54279 and n53697_not n54393_not ; n54535
g54280 and n54392_not n54535 ; n54536
g54281 and n54534_not n54536_not ; n54537
g54282 and b[45]_not n54537_not ; n54538
g54283 and n53716_not n54294 ; n54539
g54284 and n54290_not n54539 ; n54540
g54285 and n54291_not n54294_not ; n54541
g54286 and n54540_not n54541_not ; n54542
g54287 and n54394_not n54542_not ; n54543
g54288 and n53706_not n54393_not ; n54544
g54289 and n54392_not n54544 ; n54545
g54290 and n54543_not n54545_not ; n54546
g54291 and b[44]_not n54546_not ; n54547
g54292 and n53725_not n54289 ; n54548
g54293 and n54285_not n54548 ; n54549
g54294 and n54286_not n54289_not ; n54550
g54295 and n54549_not n54550_not ; n54551
g54296 and n54394_not n54551_not ; n54552
g54297 and n53715_not n54393_not ; n54553
g54298 and n54392_not n54553 ; n54554
g54299 and n54552_not n54554_not ; n54555
g54300 and b[43]_not n54555_not ; n54556
g54301 and n53734_not n54284 ; n54557
g54302 and n54280_not n54557 ; n54558
g54303 and n54281_not n54284_not ; n54559
g54304 and n54558_not n54559_not ; n54560
g54305 and n54394_not n54560_not ; n54561
g54306 and n53724_not n54393_not ; n54562
g54307 and n54392_not n54562 ; n54563
g54308 and n54561_not n54563_not ; n54564
g54309 and b[42]_not n54564_not ; n54565
g54310 and n53743_not n54279 ; n54566
g54311 and n54275_not n54566 ; n54567
g54312 and n54276_not n54279_not ; n54568
g54313 and n54567_not n54568_not ; n54569
g54314 and n54394_not n54569_not ; n54570
g54315 and n53733_not n54393_not ; n54571
g54316 and n54392_not n54571 ; n54572
g54317 and n54570_not n54572_not ; n54573
g54318 and b[41]_not n54573_not ; n54574
g54319 and n53752_not n54274 ; n54575
g54320 and n54270_not n54575 ; n54576
g54321 and n54271_not n54274_not ; n54577
g54322 and n54576_not n54577_not ; n54578
g54323 and n54394_not n54578_not ; n54579
g54324 and n53742_not n54393_not ; n54580
g54325 and n54392_not n54580 ; n54581
g54326 and n54579_not n54581_not ; n54582
g54327 and b[40]_not n54582_not ; n54583
g54328 and n53761_not n54269 ; n54584
g54329 and n54265_not n54584 ; n54585
g54330 and n54266_not n54269_not ; n54586
g54331 and n54585_not n54586_not ; n54587
g54332 and n54394_not n54587_not ; n54588
g54333 and n53751_not n54393_not ; n54589
g54334 and n54392_not n54589 ; n54590
g54335 and n54588_not n54590_not ; n54591
g54336 and b[39]_not n54591_not ; n54592
g54337 and n53770_not n54264 ; n54593
g54338 and n54260_not n54593 ; n54594
g54339 and n54261_not n54264_not ; n54595
g54340 and n54594_not n54595_not ; n54596
g54341 and n54394_not n54596_not ; n54597
g54342 and n53760_not n54393_not ; n54598
g54343 and n54392_not n54598 ; n54599
g54344 and n54597_not n54599_not ; n54600
g54345 and b[38]_not n54600_not ; n54601
g54346 and n53779_not n54259 ; n54602
g54347 and n54255_not n54602 ; n54603
g54348 and n54256_not n54259_not ; n54604
g54349 and n54603_not n54604_not ; n54605
g54350 and n54394_not n54605_not ; n54606
g54351 and n53769_not n54393_not ; n54607
g54352 and n54392_not n54607 ; n54608
g54353 and n54606_not n54608_not ; n54609
g54354 and b[37]_not n54609_not ; n54610
g54355 and n53788_not n54254 ; n54611
g54356 and n54250_not n54611 ; n54612
g54357 and n54251_not n54254_not ; n54613
g54358 and n54612_not n54613_not ; n54614
g54359 and n54394_not n54614_not ; n54615
g54360 and n53778_not n54393_not ; n54616
g54361 and n54392_not n54616 ; n54617
g54362 and n54615_not n54617_not ; n54618
g54363 and b[36]_not n54618_not ; n54619
g54364 and n53797_not n54249 ; n54620
g54365 and n54245_not n54620 ; n54621
g54366 and n54246_not n54249_not ; n54622
g54367 and n54621_not n54622_not ; n54623
g54368 and n54394_not n54623_not ; n54624
g54369 and n53787_not n54393_not ; n54625
g54370 and n54392_not n54625 ; n54626
g54371 and n54624_not n54626_not ; n54627
g54372 and b[35]_not n54627_not ; n54628
g54373 and n53806_not n54244 ; n54629
g54374 and n54240_not n54629 ; n54630
g54375 and n54241_not n54244_not ; n54631
g54376 and n54630_not n54631_not ; n54632
g54377 and n54394_not n54632_not ; n54633
g54378 and n53796_not n54393_not ; n54634
g54379 and n54392_not n54634 ; n54635
g54380 and n54633_not n54635_not ; n54636
g54381 and b[34]_not n54636_not ; n54637
g54382 and n53815_not n54239 ; n54638
g54383 and n54235_not n54638 ; n54639
g54384 and n54236_not n54239_not ; n54640
g54385 and n54639_not n54640_not ; n54641
g54386 and n54394_not n54641_not ; n54642
g54387 and n53805_not n54393_not ; n54643
g54388 and n54392_not n54643 ; n54644
g54389 and n54642_not n54644_not ; n54645
g54390 and b[33]_not n54645_not ; n54646
g54391 and n53824_not n54234 ; n54647
g54392 and n54230_not n54647 ; n54648
g54393 and n54231_not n54234_not ; n54649
g54394 and n54648_not n54649_not ; n54650
g54395 and n54394_not n54650_not ; n54651
g54396 and n53814_not n54393_not ; n54652
g54397 and n54392_not n54652 ; n54653
g54398 and n54651_not n54653_not ; n54654
g54399 and b[32]_not n54654_not ; n54655
g54400 and n53833_not n54229 ; n54656
g54401 and n54225_not n54656 ; n54657
g54402 and n54226_not n54229_not ; n54658
g54403 and n54657_not n54658_not ; n54659
g54404 and n54394_not n54659_not ; n54660
g54405 and n53823_not n54393_not ; n54661
g54406 and n54392_not n54661 ; n54662
g54407 and n54660_not n54662_not ; n54663
g54408 and b[31]_not n54663_not ; n54664
g54409 and n53842_not n54224 ; n54665
g54410 and n54220_not n54665 ; n54666
g54411 and n54221_not n54224_not ; n54667
g54412 and n54666_not n54667_not ; n54668
g54413 and n54394_not n54668_not ; n54669
g54414 and n53832_not n54393_not ; n54670
g54415 and n54392_not n54670 ; n54671
g54416 and n54669_not n54671_not ; n54672
g54417 and b[30]_not n54672_not ; n54673
g54418 and n53851_not n54219 ; n54674
g54419 and n54215_not n54674 ; n54675
g54420 and n54216_not n54219_not ; n54676
g54421 and n54675_not n54676_not ; n54677
g54422 and n54394_not n54677_not ; n54678
g54423 and n53841_not n54393_not ; n54679
g54424 and n54392_not n54679 ; n54680
g54425 and n54678_not n54680_not ; n54681
g54426 and b[29]_not n54681_not ; n54682
g54427 and n53860_not n54214 ; n54683
g54428 and n54210_not n54683 ; n54684
g54429 and n54211_not n54214_not ; n54685
g54430 and n54684_not n54685_not ; n54686
g54431 and n54394_not n54686_not ; n54687
g54432 and n53850_not n54393_not ; n54688
g54433 and n54392_not n54688 ; n54689
g54434 and n54687_not n54689_not ; n54690
g54435 and b[28]_not n54690_not ; n54691
g54436 and n53869_not n54209 ; n54692
g54437 and n54205_not n54692 ; n54693
g54438 and n54206_not n54209_not ; n54694
g54439 and n54693_not n54694_not ; n54695
g54440 and n54394_not n54695_not ; n54696
g54441 and n53859_not n54393_not ; n54697
g54442 and n54392_not n54697 ; n54698
g54443 and n54696_not n54698_not ; n54699
g54444 and b[27]_not n54699_not ; n54700
g54445 and n53878_not n54204 ; n54701
g54446 and n54200_not n54701 ; n54702
g54447 and n54201_not n54204_not ; n54703
g54448 and n54702_not n54703_not ; n54704
g54449 and n54394_not n54704_not ; n54705
g54450 and n53868_not n54393_not ; n54706
g54451 and n54392_not n54706 ; n54707
g54452 and n54705_not n54707_not ; n54708
g54453 and b[26]_not n54708_not ; n54709
g54454 and n53887_not n54199 ; n54710
g54455 and n54195_not n54710 ; n54711
g54456 and n54196_not n54199_not ; n54712
g54457 and n54711_not n54712_not ; n54713
g54458 and n54394_not n54713_not ; n54714
g54459 and n53877_not n54393_not ; n54715
g54460 and n54392_not n54715 ; n54716
g54461 and n54714_not n54716_not ; n54717
g54462 and b[25]_not n54717_not ; n54718
g54463 and n53896_not n54194 ; n54719
g54464 and n54190_not n54719 ; n54720
g54465 and n54191_not n54194_not ; n54721
g54466 and n54720_not n54721_not ; n54722
g54467 and n54394_not n54722_not ; n54723
g54468 and n53886_not n54393_not ; n54724
g54469 and n54392_not n54724 ; n54725
g54470 and n54723_not n54725_not ; n54726
g54471 and b[24]_not n54726_not ; n54727
g54472 and n53905_not n54189 ; n54728
g54473 and n54185_not n54728 ; n54729
g54474 and n54186_not n54189_not ; n54730
g54475 and n54729_not n54730_not ; n54731
g54476 and n54394_not n54731_not ; n54732
g54477 and n53895_not n54393_not ; n54733
g54478 and n54392_not n54733 ; n54734
g54479 and n54732_not n54734_not ; n54735
g54480 and b[23]_not n54735_not ; n54736
g54481 and n53914_not n54184 ; n54737
g54482 and n54180_not n54737 ; n54738
g54483 and n54181_not n54184_not ; n54739
g54484 and n54738_not n54739_not ; n54740
g54485 and n54394_not n54740_not ; n54741
g54486 and n53904_not n54393_not ; n54742
g54487 and n54392_not n54742 ; n54743
g54488 and n54741_not n54743_not ; n54744
g54489 and b[22]_not n54744_not ; n54745
g54490 and n53923_not n54179 ; n54746
g54491 and n54175_not n54746 ; n54747
g54492 and n54176_not n54179_not ; n54748
g54493 and n54747_not n54748_not ; n54749
g54494 and n54394_not n54749_not ; n54750
g54495 and n53913_not n54393_not ; n54751
g54496 and n54392_not n54751 ; n54752
g54497 and n54750_not n54752_not ; n54753
g54498 and b[21]_not n54753_not ; n54754
g54499 and n53932_not n54174 ; n54755
g54500 and n54170_not n54755 ; n54756
g54501 and n54171_not n54174_not ; n54757
g54502 and n54756_not n54757_not ; n54758
g54503 and n54394_not n54758_not ; n54759
g54504 and n53922_not n54393_not ; n54760
g54505 and n54392_not n54760 ; n54761
g54506 and n54759_not n54761_not ; n54762
g54507 and b[20]_not n54762_not ; n54763
g54508 and n53941_not n54169 ; n54764
g54509 and n54165_not n54764 ; n54765
g54510 and n54166_not n54169_not ; n54766
g54511 and n54765_not n54766_not ; n54767
g54512 and n54394_not n54767_not ; n54768
g54513 and n53931_not n54393_not ; n54769
g54514 and n54392_not n54769 ; n54770
g54515 and n54768_not n54770_not ; n54771
g54516 and b[19]_not n54771_not ; n54772
g54517 and n53950_not n54164 ; n54773
g54518 and n54160_not n54773 ; n54774
g54519 and n54161_not n54164_not ; n54775
g54520 and n54774_not n54775_not ; n54776
g54521 and n54394_not n54776_not ; n54777
g54522 and n53940_not n54393_not ; n54778
g54523 and n54392_not n54778 ; n54779
g54524 and n54777_not n54779_not ; n54780
g54525 and b[18]_not n54780_not ; n54781
g54526 and n53959_not n54159 ; n54782
g54527 and n54155_not n54782 ; n54783
g54528 and n54156_not n54159_not ; n54784
g54529 and n54783_not n54784_not ; n54785
g54530 and n54394_not n54785_not ; n54786
g54531 and n53949_not n54393_not ; n54787
g54532 and n54392_not n54787 ; n54788
g54533 and n54786_not n54788_not ; n54789
g54534 and b[17]_not n54789_not ; n54790
g54535 and n53968_not n54154 ; n54791
g54536 and n54150_not n54791 ; n54792
g54537 and n54151_not n54154_not ; n54793
g54538 and n54792_not n54793_not ; n54794
g54539 and n54394_not n54794_not ; n54795
g54540 and n53958_not n54393_not ; n54796
g54541 and n54392_not n54796 ; n54797
g54542 and n54795_not n54797_not ; n54798
g54543 and b[16]_not n54798_not ; n54799
g54544 and n53977_not n54149 ; n54800
g54545 and n54145_not n54800 ; n54801
g54546 and n54146_not n54149_not ; n54802
g54547 and n54801_not n54802_not ; n54803
g54548 and n54394_not n54803_not ; n54804
g54549 and n53967_not n54393_not ; n54805
g54550 and n54392_not n54805 ; n54806
g54551 and n54804_not n54806_not ; n54807
g54552 and b[15]_not n54807_not ; n54808
g54553 and n53986_not n54144 ; n54809
g54554 and n54140_not n54809 ; n54810
g54555 and n54141_not n54144_not ; n54811
g54556 and n54810_not n54811_not ; n54812
g54557 and n54394_not n54812_not ; n54813
g54558 and n53976_not n54393_not ; n54814
g54559 and n54392_not n54814 ; n54815
g54560 and n54813_not n54815_not ; n54816
g54561 and b[14]_not n54816_not ; n54817
g54562 and n53995_not n54139 ; n54818
g54563 and n54135_not n54818 ; n54819
g54564 and n54136_not n54139_not ; n54820
g54565 and n54819_not n54820_not ; n54821
g54566 and n54394_not n54821_not ; n54822
g54567 and n53985_not n54393_not ; n54823
g54568 and n54392_not n54823 ; n54824
g54569 and n54822_not n54824_not ; n54825
g54570 and b[13]_not n54825_not ; n54826
g54571 and n54004_not n54134 ; n54827
g54572 and n54130_not n54827 ; n54828
g54573 and n54131_not n54134_not ; n54829
g54574 and n54828_not n54829_not ; n54830
g54575 and n54394_not n54830_not ; n54831
g54576 and n53994_not n54393_not ; n54832
g54577 and n54392_not n54832 ; n54833
g54578 and n54831_not n54833_not ; n54834
g54579 and b[12]_not n54834_not ; n54835
g54580 and n54013_not n54129 ; n54836
g54581 and n54125_not n54836 ; n54837
g54582 and n54126_not n54129_not ; n54838
g54583 and n54837_not n54838_not ; n54839
g54584 and n54394_not n54839_not ; n54840
g54585 and n54003_not n54393_not ; n54841
g54586 and n54392_not n54841 ; n54842
g54587 and n54840_not n54842_not ; n54843
g54588 and b[11]_not n54843_not ; n54844
g54589 and n54022_not n54124 ; n54845
g54590 and n54120_not n54845 ; n54846
g54591 and n54121_not n54124_not ; n54847
g54592 and n54846_not n54847_not ; n54848
g54593 and n54394_not n54848_not ; n54849
g54594 and n54012_not n54393_not ; n54850
g54595 and n54392_not n54850 ; n54851
g54596 and n54849_not n54851_not ; n54852
g54597 and b[10]_not n54852_not ; n54853
g54598 and n54031_not n54119 ; n54854
g54599 and n54115_not n54854 ; n54855
g54600 and n54116_not n54119_not ; n54856
g54601 and n54855_not n54856_not ; n54857
g54602 and n54394_not n54857_not ; n54858
g54603 and n54021_not n54393_not ; n54859
g54604 and n54392_not n54859 ; n54860
g54605 and n54858_not n54860_not ; n54861
g54606 and b[9]_not n54861_not ; n54862
g54607 and n54040_not n54114 ; n54863
g54608 and n54110_not n54863 ; n54864
g54609 and n54111_not n54114_not ; n54865
g54610 and n54864_not n54865_not ; n54866
g54611 and n54394_not n54866_not ; n54867
g54612 and n54030_not n54393_not ; n54868
g54613 and n54392_not n54868 ; n54869
g54614 and n54867_not n54869_not ; n54870
g54615 and b[8]_not n54870_not ; n54871
g54616 and n54049_not n54109 ; n54872
g54617 and n54105_not n54872 ; n54873
g54618 and n54106_not n54109_not ; n54874
g54619 and n54873_not n54874_not ; n54875
g54620 and n54394_not n54875_not ; n54876
g54621 and n54039_not n54393_not ; n54877
g54622 and n54392_not n54877 ; n54878
g54623 and n54876_not n54878_not ; n54879
g54624 and b[7]_not n54879_not ; n54880
g54625 and n54058_not n54104 ; n54881
g54626 and n54100_not n54881 ; n54882
g54627 and n54101_not n54104_not ; n54883
g54628 and n54882_not n54883_not ; n54884
g54629 and n54394_not n54884_not ; n54885
g54630 and n54048_not n54393_not ; n54886
g54631 and n54392_not n54886 ; n54887
g54632 and n54885_not n54887_not ; n54888
g54633 and b[6]_not n54888_not ; n54889
g54634 and n54067_not n54099 ; n54890
g54635 and n54095_not n54890 ; n54891
g54636 and n54096_not n54099_not ; n54892
g54637 and n54891_not n54892_not ; n54893
g54638 and n54394_not n54893_not ; n54894
g54639 and n54057_not n54393_not ; n54895
g54640 and n54392_not n54895 ; n54896
g54641 and n54894_not n54896_not ; n54897
g54642 and b[5]_not n54897_not ; n54898
g54643 and n54075_not n54094 ; n54899
g54644 and n54090_not n54899 ; n54900
g54645 and n54091_not n54094_not ; n54901
g54646 and n54900_not n54901_not ; n54902
g54647 and n54394_not n54902_not ; n54903
g54648 and n54066_not n54393_not ; n54904
g54649 and n54392_not n54904 ; n54905
g54650 and n54903_not n54905_not ; n54906
g54651 and b[4]_not n54906_not ; n54907
g54652 and n54085_not n54089 ; n54908
g54653 and n54084_not n54908 ; n54909
g54654 and n54086_not n54089_not ; n54910
g54655 and n54909_not n54910_not ; n54911
g54656 and n54394_not n54911_not ; n54912
g54657 and n54074_not n54393_not ; n54913
g54658 and n54392_not n54913 ; n54914
g54659 and n54912_not n54914_not ; n54915
g54660 and b[3]_not n54915_not ; n54916
g54661 and n26069 n54082_not ; n54917
g54662 and n54080_not n54917 ; n54918
g54663 and n54084_not n54918_not ; n54919
g54664 and n54394_not n54919 ; n54920
g54665 and n54079_not n54393_not ; n54921
g54666 and n54392_not n54921 ; n54922
g54667 and n54920_not n54922_not ; n54923
g54668 and b[2]_not n54923_not ; n54924
g54669 and b[0] n54394_not ; n54925
g54670 and a[3] n54925_not ; n54926
g54671 and n26069 n54394_not ; n54927
g54672 and n54926_not n54927_not ; n54928
g54673 and b[1] n54928_not ; n54929
g54674 and b[1]_not n54927_not ; n54930
g54675 and n54926_not n54930 ; n54931
g54676 and n54929_not n54931_not ; n54932
g54677 and n26919_not n54932_not ; n54933
g54678 and b[1]_not n54928_not ; n54934
g54679 and n54933_not n54934_not ; n54935
g54680 and b[2] n54922_not ; n54936
g54681 and n54920_not n54936 ; n54937
g54682 and n54924_not n54937_not ; n54938
g54683 and n54935_not n54938 ; n54939
g54684 and n54924_not n54939_not ; n54940
g54685 and b[3] n54914_not ; n54941
g54686 and n54912_not n54941 ; n54942
g54687 and n54916_not n54942_not ; n54943
g54688 and n54940_not n54943 ; n54944
g54689 and n54916_not n54944_not ; n54945
g54690 and b[4] n54905_not ; n54946
g54691 and n54903_not n54946 ; n54947
g54692 and n54907_not n54947_not ; n54948
g54693 and n54945_not n54948 ; n54949
g54694 and n54907_not n54949_not ; n54950
g54695 and b[5] n54896_not ; n54951
g54696 and n54894_not n54951 ; n54952
g54697 and n54898_not n54952_not ; n54953
g54698 and n54950_not n54953 ; n54954
g54699 and n54898_not n54954_not ; n54955
g54700 and b[6] n54887_not ; n54956
g54701 and n54885_not n54956 ; n54957
g54702 and n54889_not n54957_not ; n54958
g54703 and n54955_not n54958 ; n54959
g54704 and n54889_not n54959_not ; n54960
g54705 and b[7] n54878_not ; n54961
g54706 and n54876_not n54961 ; n54962
g54707 and n54880_not n54962_not ; n54963
g54708 and n54960_not n54963 ; n54964
g54709 and n54880_not n54964_not ; n54965
g54710 and b[8] n54869_not ; n54966
g54711 and n54867_not n54966 ; n54967
g54712 and n54871_not n54967_not ; n54968
g54713 and n54965_not n54968 ; n54969
g54714 and n54871_not n54969_not ; n54970
g54715 and b[9] n54860_not ; n54971
g54716 and n54858_not n54971 ; n54972
g54717 and n54862_not n54972_not ; n54973
g54718 and n54970_not n54973 ; n54974
g54719 and n54862_not n54974_not ; n54975
g54720 and b[10] n54851_not ; n54976
g54721 and n54849_not n54976 ; n54977
g54722 and n54853_not n54977_not ; n54978
g54723 and n54975_not n54978 ; n54979
g54724 and n54853_not n54979_not ; n54980
g54725 and b[11] n54842_not ; n54981
g54726 and n54840_not n54981 ; n54982
g54727 and n54844_not n54982_not ; n54983
g54728 and n54980_not n54983 ; n54984
g54729 and n54844_not n54984_not ; n54985
g54730 and b[12] n54833_not ; n54986
g54731 and n54831_not n54986 ; n54987
g54732 and n54835_not n54987_not ; n54988
g54733 and n54985_not n54988 ; n54989
g54734 and n54835_not n54989_not ; n54990
g54735 and b[13] n54824_not ; n54991
g54736 and n54822_not n54991 ; n54992
g54737 and n54826_not n54992_not ; n54993
g54738 and n54990_not n54993 ; n54994
g54739 and n54826_not n54994_not ; n54995
g54740 and b[14] n54815_not ; n54996
g54741 and n54813_not n54996 ; n54997
g54742 and n54817_not n54997_not ; n54998
g54743 and n54995_not n54998 ; n54999
g54744 and n54817_not n54999_not ; n55000
g54745 and b[15] n54806_not ; n55001
g54746 and n54804_not n55001 ; n55002
g54747 and n54808_not n55002_not ; n55003
g54748 and n55000_not n55003 ; n55004
g54749 and n54808_not n55004_not ; n55005
g54750 and b[16] n54797_not ; n55006
g54751 and n54795_not n55006 ; n55007
g54752 and n54799_not n55007_not ; n55008
g54753 and n55005_not n55008 ; n55009
g54754 and n54799_not n55009_not ; n55010
g54755 and b[17] n54788_not ; n55011
g54756 and n54786_not n55011 ; n55012
g54757 and n54790_not n55012_not ; n55013
g54758 and n55010_not n55013 ; n55014
g54759 and n54790_not n55014_not ; n55015
g54760 and b[18] n54779_not ; n55016
g54761 and n54777_not n55016 ; n55017
g54762 and n54781_not n55017_not ; n55018
g54763 and n55015_not n55018 ; n55019
g54764 and n54781_not n55019_not ; n55020
g54765 and b[19] n54770_not ; n55021
g54766 and n54768_not n55021 ; n55022
g54767 and n54772_not n55022_not ; n55023
g54768 and n55020_not n55023 ; n55024
g54769 and n54772_not n55024_not ; n55025
g54770 and b[20] n54761_not ; n55026
g54771 and n54759_not n55026 ; n55027
g54772 and n54763_not n55027_not ; n55028
g54773 and n55025_not n55028 ; n55029
g54774 and n54763_not n55029_not ; n55030
g54775 and b[21] n54752_not ; n55031
g54776 and n54750_not n55031 ; n55032
g54777 and n54754_not n55032_not ; n55033
g54778 and n55030_not n55033 ; n55034
g54779 and n54754_not n55034_not ; n55035
g54780 and b[22] n54743_not ; n55036
g54781 and n54741_not n55036 ; n55037
g54782 and n54745_not n55037_not ; n55038
g54783 and n55035_not n55038 ; n55039
g54784 and n54745_not n55039_not ; n55040
g54785 and b[23] n54734_not ; n55041
g54786 and n54732_not n55041 ; n55042
g54787 and n54736_not n55042_not ; n55043
g54788 and n55040_not n55043 ; n55044
g54789 and n54736_not n55044_not ; n55045
g54790 and b[24] n54725_not ; n55046
g54791 and n54723_not n55046 ; n55047
g54792 and n54727_not n55047_not ; n55048
g54793 and n55045_not n55048 ; n55049
g54794 and n54727_not n55049_not ; n55050
g54795 and b[25] n54716_not ; n55051
g54796 and n54714_not n55051 ; n55052
g54797 and n54718_not n55052_not ; n55053
g54798 and n55050_not n55053 ; n55054
g54799 and n54718_not n55054_not ; n55055
g54800 and b[26] n54707_not ; n55056
g54801 and n54705_not n55056 ; n55057
g54802 and n54709_not n55057_not ; n55058
g54803 and n55055_not n55058 ; n55059
g54804 and n54709_not n55059_not ; n55060
g54805 and b[27] n54698_not ; n55061
g54806 and n54696_not n55061 ; n55062
g54807 and n54700_not n55062_not ; n55063
g54808 and n55060_not n55063 ; n55064
g54809 and n54700_not n55064_not ; n55065
g54810 and b[28] n54689_not ; n55066
g54811 and n54687_not n55066 ; n55067
g54812 and n54691_not n55067_not ; n55068
g54813 and n55065_not n55068 ; n55069
g54814 and n54691_not n55069_not ; n55070
g54815 and b[29] n54680_not ; n55071
g54816 and n54678_not n55071 ; n55072
g54817 and n54682_not n55072_not ; n55073
g54818 and n55070_not n55073 ; n55074
g54819 and n54682_not n55074_not ; n55075
g54820 and b[30] n54671_not ; n55076
g54821 and n54669_not n55076 ; n55077
g54822 and n54673_not n55077_not ; n55078
g54823 and n55075_not n55078 ; n55079
g54824 and n54673_not n55079_not ; n55080
g54825 and b[31] n54662_not ; n55081
g54826 and n54660_not n55081 ; n55082
g54827 and n54664_not n55082_not ; n55083
g54828 and n55080_not n55083 ; n55084
g54829 and n54664_not n55084_not ; n55085
g54830 and b[32] n54653_not ; n55086
g54831 and n54651_not n55086 ; n55087
g54832 and n54655_not n55087_not ; n55088
g54833 and n55085_not n55088 ; n55089
g54834 and n54655_not n55089_not ; n55090
g54835 and b[33] n54644_not ; n55091
g54836 and n54642_not n55091 ; n55092
g54837 and n54646_not n55092_not ; n55093
g54838 and n55090_not n55093 ; n55094
g54839 and n54646_not n55094_not ; n55095
g54840 and b[34] n54635_not ; n55096
g54841 and n54633_not n55096 ; n55097
g54842 and n54637_not n55097_not ; n55098
g54843 and n55095_not n55098 ; n55099
g54844 and n54637_not n55099_not ; n55100
g54845 and b[35] n54626_not ; n55101
g54846 and n54624_not n55101 ; n55102
g54847 and n54628_not n55102_not ; n55103
g54848 and n55100_not n55103 ; n55104
g54849 and n54628_not n55104_not ; n55105
g54850 and b[36] n54617_not ; n55106
g54851 and n54615_not n55106 ; n55107
g54852 and n54619_not n55107_not ; n55108
g54853 and n55105_not n55108 ; n55109
g54854 and n54619_not n55109_not ; n55110
g54855 and b[37] n54608_not ; n55111
g54856 and n54606_not n55111 ; n55112
g54857 and n54610_not n55112_not ; n55113
g54858 and n55110_not n55113 ; n55114
g54859 and n54610_not n55114_not ; n55115
g54860 and b[38] n54599_not ; n55116
g54861 and n54597_not n55116 ; n55117
g54862 and n54601_not n55117_not ; n55118
g54863 and n55115_not n55118 ; n55119
g54864 and n54601_not n55119_not ; n55120
g54865 and b[39] n54590_not ; n55121
g54866 and n54588_not n55121 ; n55122
g54867 and n54592_not n55122_not ; n55123
g54868 and n55120_not n55123 ; n55124
g54869 and n54592_not n55124_not ; n55125
g54870 and b[40] n54581_not ; n55126
g54871 and n54579_not n55126 ; n55127
g54872 and n54583_not n55127_not ; n55128
g54873 and n55125_not n55128 ; n55129
g54874 and n54583_not n55129_not ; n55130
g54875 and b[41] n54572_not ; n55131
g54876 and n54570_not n55131 ; n55132
g54877 and n54574_not n55132_not ; n55133
g54878 and n55130_not n55133 ; n55134
g54879 and n54574_not n55134_not ; n55135
g54880 and b[42] n54563_not ; n55136
g54881 and n54561_not n55136 ; n55137
g54882 and n54565_not n55137_not ; n55138
g54883 and n55135_not n55138 ; n55139
g54884 and n54565_not n55139_not ; n55140
g54885 and b[43] n54554_not ; n55141
g54886 and n54552_not n55141 ; n55142
g54887 and n54556_not n55142_not ; n55143
g54888 and n55140_not n55143 ; n55144
g54889 and n54556_not n55144_not ; n55145
g54890 and b[44] n54545_not ; n55146
g54891 and n54543_not n55146 ; n55147
g54892 and n54547_not n55147_not ; n55148
g54893 and n55145_not n55148 ; n55149
g54894 and n54547_not n55149_not ; n55150
g54895 and b[45] n54536_not ; n55151
g54896 and n54534_not n55151 ; n55152
g54897 and n54538_not n55152_not ; n55153
g54898 and n55150_not n55153 ; n55154
g54899 and n54538_not n55154_not ; n55155
g54900 and b[46] n54527_not ; n55156
g54901 and n54525_not n55156 ; n55157
g54902 and n54529_not n55157_not ; n55158
g54903 and n55155_not n55158 ; n55159
g54904 and n54529_not n55159_not ; n55160
g54905 and b[47] n54518_not ; n55161
g54906 and n54516_not n55161 ; n55162
g54907 and n54520_not n55162_not ; n55163
g54908 and n55160_not n55163 ; n55164
g54909 and n54520_not n55164_not ; n55165
g54910 and b[48] n54509_not ; n55166
g54911 and n54507_not n55166 ; n55167
g54912 and n54511_not n55167_not ; n55168
g54913 and n55165_not n55168 ; n55169
g54914 and n54511_not n55169_not ; n55170
g54915 and b[49] n54500_not ; n55171
g54916 and n54498_not n55171 ; n55172
g54917 and n54502_not n55172_not ; n55173
g54918 and n55170_not n55173 ; n55174
g54919 and n54502_not n55174_not ; n55175
g54920 and b[50] n54491_not ; n55176
g54921 and n54489_not n55176 ; n55177
g54922 and n54493_not n55177_not ; n55178
g54923 and n55175_not n55178 ; n55179
g54924 and n54493_not n55179_not ; n55180
g54925 and b[51] n54482_not ; n55181
g54926 and n54480_not n55181 ; n55182
g54927 and n54484_not n55182_not ; n55183
g54928 and n55180_not n55183 ; n55184
g54929 and n54484_not n55184_not ; n55185
g54930 and b[52] n54473_not ; n55186
g54931 and n54471_not n55186 ; n55187
g54932 and n54475_not n55187_not ; n55188
g54933 and n55185_not n55188 ; n55189
g54934 and n54475_not n55189_not ; n55190
g54935 and b[53] n54464_not ; n55191
g54936 and n54462_not n55191 ; n55192
g54937 and n54466_not n55192_not ; n55193
g54938 and n55190_not n55193 ; n55194
g54939 and n54466_not n55194_not ; n55195
g54940 and b[54] n54455_not ; n55196
g54941 and n54453_not n55196 ; n55197
g54942 and n54457_not n55197_not ; n55198
g54943 and n55195_not n55198 ; n55199
g54944 and n54457_not n55199_not ; n55200
g54945 and b[55] n54446_not ; n55201
g54946 and n54444_not n55201 ; n55202
g54947 and n54448_not n55202_not ; n55203
g54948 and n55200_not n55203 ; n55204
g54949 and n54448_not n55204_not ; n55205
g54950 and b[56] n54437_not ; n55206
g54951 and n54435_not n55206 ; n55207
g54952 and n54439_not n55207_not ; n55208
g54953 and n55205_not n55208 ; n55209
g54954 and n54439_not n55209_not ; n55210
g54955 and b[57] n54428_not ; n55211
g54956 and n54426_not n55211 ; n55212
g54957 and n54430_not n55212_not ; n55213
g54958 and n55210_not n55213 ; n55214
g54959 and n54430_not n55214_not ; n55215
g54960 and b[58] n54419_not ; n55216
g54961 and n54417_not n55216 ; n55217
g54962 and n54421_not n55217_not ; n55218
g54963 and n55215_not n55218 ; n55219
g54964 and n54421_not n55219_not ; n55220
g54965 and b[59] n54410_not ; n55221
g54966 and n54408_not n55221 ; n55222
g54967 and n54412_not n55222_not ; n55223
g54968 and n55220_not n55223 ; n55224
g54969 and n54412_not n55224_not ; n55225
g54970 and b[60] n54401_not ; n55226
g54971 and n54399_not n55226 ; n55227
g54972 and n54403_not n55227_not ; n55228
g54973 and n55225_not n55228 ; n55229
g54974 and n54403_not n55229_not ; n55230
g54975 and n53563_not n54389_not ; n55231
g54976 and n54387_not n55231 ; n55232
g54977 and n54375_not n55232 ; n55233
g54978 and n54387_not n54389_not ; n55234
g54979 and n54376_not n55234_not ; n55235
g54980 and n55233_not n55235_not ; n55236
g54981 and n54394_not n55236_not ; n55237
g54982 and n54386_not n54393_not ; n55238
g54983 and n54392_not n55238 ; n55239
g54984 and n55237_not n55239_not ; n55240
g54985 and b[61]_not n55240_not ; n55241
g54986 and b[61] n55239_not ; n55242
g54987 and n55237_not n55242 ; n55243
g54988 and n279 n55243_not ; n55244
g54989 and n55241_not n55244 ; n55245
g54990 and n55230_not n55245 ; n55246
g54991 and n403 n55240_not ; n55247
g54992 and n55246_not n55247_not ; n55248
g54993 and n54412_not n55228 ; n55249
g54994 and n55224_not n55249 ; n55250
g54995 and n55225_not n55228_not ; n55251
g54996 and n55250_not n55251_not ; n55252
g54997 and n55248_not n55252_not ; n55253
g54998 and n54402_not n55247_not ; n55254
g54999 and n55246_not n55254 ; n55255
g55000 and n55253_not n55255_not ; n55256
g55001 and b[61]_not n55256_not ; n55257
g55002 and n54421_not n55223 ; n55258
g55003 and n55219_not n55258 ; n55259
g55004 and n55220_not n55223_not ; n55260
g55005 and n55259_not n55260_not ; n55261
g55006 and n55248_not n55261_not ; n55262
g55007 and n54411_not n55247_not ; n55263
g55008 and n55246_not n55263 ; n55264
g55009 and n55262_not n55264_not ; n55265
g55010 and b[60]_not n55265_not ; n55266
g55011 and n54430_not n55218 ; n55267
g55012 and n55214_not n55267 ; n55268
g55013 and n55215_not n55218_not ; n55269
g55014 and n55268_not n55269_not ; n55270
g55015 and n55248_not n55270_not ; n55271
g55016 and n54420_not n55247_not ; n55272
g55017 and n55246_not n55272 ; n55273
g55018 and n55271_not n55273_not ; n55274
g55019 and b[59]_not n55274_not ; n55275
g55020 and n54439_not n55213 ; n55276
g55021 and n55209_not n55276 ; n55277
g55022 and n55210_not n55213_not ; n55278
g55023 and n55277_not n55278_not ; n55279
g55024 and n55248_not n55279_not ; n55280
g55025 and n54429_not n55247_not ; n55281
g55026 and n55246_not n55281 ; n55282
g55027 and n55280_not n55282_not ; n55283
g55028 and b[58]_not n55283_not ; n55284
g55029 and n54448_not n55208 ; n55285
g55030 and n55204_not n55285 ; n55286
g55031 and n55205_not n55208_not ; n55287
g55032 and n55286_not n55287_not ; n55288
g55033 and n55248_not n55288_not ; n55289
g55034 and n54438_not n55247_not ; n55290
g55035 and n55246_not n55290 ; n55291
g55036 and n55289_not n55291_not ; n55292
g55037 and b[57]_not n55292_not ; n55293
g55038 and n54457_not n55203 ; n55294
g55039 and n55199_not n55294 ; n55295
g55040 and n55200_not n55203_not ; n55296
g55041 and n55295_not n55296_not ; n55297
g55042 and n55248_not n55297_not ; n55298
g55043 and n54447_not n55247_not ; n55299
g55044 and n55246_not n55299 ; n55300
g55045 and n55298_not n55300_not ; n55301
g55046 and b[56]_not n55301_not ; n55302
g55047 and n54466_not n55198 ; n55303
g55048 and n55194_not n55303 ; n55304
g55049 and n55195_not n55198_not ; n55305
g55050 and n55304_not n55305_not ; n55306
g55051 and n55248_not n55306_not ; n55307
g55052 and n54456_not n55247_not ; n55308
g55053 and n55246_not n55308 ; n55309
g55054 and n55307_not n55309_not ; n55310
g55055 and b[55]_not n55310_not ; n55311
g55056 and n54475_not n55193 ; n55312
g55057 and n55189_not n55312 ; n55313
g55058 and n55190_not n55193_not ; n55314
g55059 and n55313_not n55314_not ; n55315
g55060 and n55248_not n55315_not ; n55316
g55061 and n54465_not n55247_not ; n55317
g55062 and n55246_not n55317 ; n55318
g55063 and n55316_not n55318_not ; n55319
g55064 and b[54]_not n55319_not ; n55320
g55065 and n54484_not n55188 ; n55321
g55066 and n55184_not n55321 ; n55322
g55067 and n55185_not n55188_not ; n55323
g55068 and n55322_not n55323_not ; n55324
g55069 and n55248_not n55324_not ; n55325
g55070 and n54474_not n55247_not ; n55326
g55071 and n55246_not n55326 ; n55327
g55072 and n55325_not n55327_not ; n55328
g55073 and b[53]_not n55328_not ; n55329
g55074 and n54493_not n55183 ; n55330
g55075 and n55179_not n55330 ; n55331
g55076 and n55180_not n55183_not ; n55332
g55077 and n55331_not n55332_not ; n55333
g55078 and n55248_not n55333_not ; n55334
g55079 and n54483_not n55247_not ; n55335
g55080 and n55246_not n55335 ; n55336
g55081 and n55334_not n55336_not ; n55337
g55082 and b[52]_not n55337_not ; n55338
g55083 and n54502_not n55178 ; n55339
g55084 and n55174_not n55339 ; n55340
g55085 and n55175_not n55178_not ; n55341
g55086 and n55340_not n55341_not ; n55342
g55087 and n55248_not n55342_not ; n55343
g55088 and n54492_not n55247_not ; n55344
g55089 and n55246_not n55344 ; n55345
g55090 and n55343_not n55345_not ; n55346
g55091 and b[51]_not n55346_not ; n55347
g55092 and n54511_not n55173 ; n55348
g55093 and n55169_not n55348 ; n55349
g55094 and n55170_not n55173_not ; n55350
g55095 and n55349_not n55350_not ; n55351
g55096 and n55248_not n55351_not ; n55352
g55097 and n54501_not n55247_not ; n55353
g55098 and n55246_not n55353 ; n55354
g55099 and n55352_not n55354_not ; n55355
g55100 and b[50]_not n55355_not ; n55356
g55101 and n54520_not n55168 ; n55357
g55102 and n55164_not n55357 ; n55358
g55103 and n55165_not n55168_not ; n55359
g55104 and n55358_not n55359_not ; n55360
g55105 and n55248_not n55360_not ; n55361
g55106 and n54510_not n55247_not ; n55362
g55107 and n55246_not n55362 ; n55363
g55108 and n55361_not n55363_not ; n55364
g55109 and b[49]_not n55364_not ; n55365
g55110 and n54529_not n55163 ; n55366
g55111 and n55159_not n55366 ; n55367
g55112 and n55160_not n55163_not ; n55368
g55113 and n55367_not n55368_not ; n55369
g55114 and n55248_not n55369_not ; n55370
g55115 and n54519_not n55247_not ; n55371
g55116 and n55246_not n55371 ; n55372
g55117 and n55370_not n55372_not ; n55373
g55118 and b[48]_not n55373_not ; n55374
g55119 and n54538_not n55158 ; n55375
g55120 and n55154_not n55375 ; n55376
g55121 and n55155_not n55158_not ; n55377
g55122 and n55376_not n55377_not ; n55378
g55123 and n55248_not n55378_not ; n55379
g55124 and n54528_not n55247_not ; n55380
g55125 and n55246_not n55380 ; n55381
g55126 and n55379_not n55381_not ; n55382
g55127 and b[47]_not n55382_not ; n55383
g55128 and n54547_not n55153 ; n55384
g55129 and n55149_not n55384 ; n55385
g55130 and n55150_not n55153_not ; n55386
g55131 and n55385_not n55386_not ; n55387
g55132 and n55248_not n55387_not ; n55388
g55133 and n54537_not n55247_not ; n55389
g55134 and n55246_not n55389 ; n55390
g55135 and n55388_not n55390_not ; n55391
g55136 and b[46]_not n55391_not ; n55392
g55137 and n54556_not n55148 ; n55393
g55138 and n55144_not n55393 ; n55394
g55139 and n55145_not n55148_not ; n55395
g55140 and n55394_not n55395_not ; n55396
g55141 and n55248_not n55396_not ; n55397
g55142 and n54546_not n55247_not ; n55398
g55143 and n55246_not n55398 ; n55399
g55144 and n55397_not n55399_not ; n55400
g55145 and b[45]_not n55400_not ; n55401
g55146 and n54565_not n55143 ; n55402
g55147 and n55139_not n55402 ; n55403
g55148 and n55140_not n55143_not ; n55404
g55149 and n55403_not n55404_not ; n55405
g55150 and n55248_not n55405_not ; n55406
g55151 and n54555_not n55247_not ; n55407
g55152 and n55246_not n55407 ; n55408
g55153 and n55406_not n55408_not ; n55409
g55154 and b[44]_not n55409_not ; n55410
g55155 and n54574_not n55138 ; n55411
g55156 and n55134_not n55411 ; n55412
g55157 and n55135_not n55138_not ; n55413
g55158 and n55412_not n55413_not ; n55414
g55159 and n55248_not n55414_not ; n55415
g55160 and n54564_not n55247_not ; n55416
g55161 and n55246_not n55416 ; n55417
g55162 and n55415_not n55417_not ; n55418
g55163 and b[43]_not n55418_not ; n55419
g55164 and n54583_not n55133 ; n55420
g55165 and n55129_not n55420 ; n55421
g55166 and n55130_not n55133_not ; n55422
g55167 and n55421_not n55422_not ; n55423
g55168 and n55248_not n55423_not ; n55424
g55169 and n54573_not n55247_not ; n55425
g55170 and n55246_not n55425 ; n55426
g55171 and n55424_not n55426_not ; n55427
g55172 and b[42]_not n55427_not ; n55428
g55173 and n54592_not n55128 ; n55429
g55174 and n55124_not n55429 ; n55430
g55175 and n55125_not n55128_not ; n55431
g55176 and n55430_not n55431_not ; n55432
g55177 and n55248_not n55432_not ; n55433
g55178 and n54582_not n55247_not ; n55434
g55179 and n55246_not n55434 ; n55435
g55180 and n55433_not n55435_not ; n55436
g55181 and b[41]_not n55436_not ; n55437
g55182 and n54601_not n55123 ; n55438
g55183 and n55119_not n55438 ; n55439
g55184 and n55120_not n55123_not ; n55440
g55185 and n55439_not n55440_not ; n55441
g55186 and n55248_not n55441_not ; n55442
g55187 and n54591_not n55247_not ; n55443
g55188 and n55246_not n55443 ; n55444
g55189 and n55442_not n55444_not ; n55445
g55190 and b[40]_not n55445_not ; n55446
g55191 and n54610_not n55118 ; n55447
g55192 and n55114_not n55447 ; n55448
g55193 and n55115_not n55118_not ; n55449
g55194 and n55448_not n55449_not ; n55450
g55195 and n55248_not n55450_not ; n55451
g55196 and n54600_not n55247_not ; n55452
g55197 and n55246_not n55452 ; n55453
g55198 and n55451_not n55453_not ; n55454
g55199 and b[39]_not n55454_not ; n55455
g55200 and n54619_not n55113 ; n55456
g55201 and n55109_not n55456 ; n55457
g55202 and n55110_not n55113_not ; n55458
g55203 and n55457_not n55458_not ; n55459
g55204 and n55248_not n55459_not ; n55460
g55205 and n54609_not n55247_not ; n55461
g55206 and n55246_not n55461 ; n55462
g55207 and n55460_not n55462_not ; n55463
g55208 and b[38]_not n55463_not ; n55464
g55209 and n54628_not n55108 ; n55465
g55210 and n55104_not n55465 ; n55466
g55211 and n55105_not n55108_not ; n55467
g55212 and n55466_not n55467_not ; n55468
g55213 and n55248_not n55468_not ; n55469
g55214 and n54618_not n55247_not ; n55470
g55215 and n55246_not n55470 ; n55471
g55216 and n55469_not n55471_not ; n55472
g55217 and b[37]_not n55472_not ; n55473
g55218 and n54637_not n55103 ; n55474
g55219 and n55099_not n55474 ; n55475
g55220 and n55100_not n55103_not ; n55476
g55221 and n55475_not n55476_not ; n55477
g55222 and n55248_not n55477_not ; n55478
g55223 and n54627_not n55247_not ; n55479
g55224 and n55246_not n55479 ; n55480
g55225 and n55478_not n55480_not ; n55481
g55226 and b[36]_not n55481_not ; n55482
g55227 and n54646_not n55098 ; n55483
g55228 and n55094_not n55483 ; n55484
g55229 and n55095_not n55098_not ; n55485
g55230 and n55484_not n55485_not ; n55486
g55231 and n55248_not n55486_not ; n55487
g55232 and n54636_not n55247_not ; n55488
g55233 and n55246_not n55488 ; n55489
g55234 and n55487_not n55489_not ; n55490
g55235 and b[35]_not n55490_not ; n55491
g55236 and n54655_not n55093 ; n55492
g55237 and n55089_not n55492 ; n55493
g55238 and n55090_not n55093_not ; n55494
g55239 and n55493_not n55494_not ; n55495
g55240 and n55248_not n55495_not ; n55496
g55241 and n54645_not n55247_not ; n55497
g55242 and n55246_not n55497 ; n55498
g55243 and n55496_not n55498_not ; n55499
g55244 and b[34]_not n55499_not ; n55500
g55245 and n54664_not n55088 ; n55501
g55246 and n55084_not n55501 ; n55502
g55247 and n55085_not n55088_not ; n55503
g55248 and n55502_not n55503_not ; n55504
g55249 and n55248_not n55504_not ; n55505
g55250 and n54654_not n55247_not ; n55506
g55251 and n55246_not n55506 ; n55507
g55252 and n55505_not n55507_not ; n55508
g55253 and b[33]_not n55508_not ; n55509
g55254 and n54673_not n55083 ; n55510
g55255 and n55079_not n55510 ; n55511
g55256 and n55080_not n55083_not ; n55512
g55257 and n55511_not n55512_not ; n55513
g55258 and n55248_not n55513_not ; n55514
g55259 and n54663_not n55247_not ; n55515
g55260 and n55246_not n55515 ; n55516
g55261 and n55514_not n55516_not ; n55517
g55262 and b[32]_not n55517_not ; n55518
g55263 and n54682_not n55078 ; n55519
g55264 and n55074_not n55519 ; n55520
g55265 and n55075_not n55078_not ; n55521
g55266 and n55520_not n55521_not ; n55522
g55267 and n55248_not n55522_not ; n55523
g55268 and n54672_not n55247_not ; n55524
g55269 and n55246_not n55524 ; n55525
g55270 and n55523_not n55525_not ; n55526
g55271 and b[31]_not n55526_not ; n55527
g55272 and n54691_not n55073 ; n55528
g55273 and n55069_not n55528 ; n55529
g55274 and n55070_not n55073_not ; n55530
g55275 and n55529_not n55530_not ; n55531
g55276 and n55248_not n55531_not ; n55532
g55277 and n54681_not n55247_not ; n55533
g55278 and n55246_not n55533 ; n55534
g55279 and n55532_not n55534_not ; n55535
g55280 and b[30]_not n55535_not ; n55536
g55281 and n54700_not n55068 ; n55537
g55282 and n55064_not n55537 ; n55538
g55283 and n55065_not n55068_not ; n55539
g55284 and n55538_not n55539_not ; n55540
g55285 and n55248_not n55540_not ; n55541
g55286 and n54690_not n55247_not ; n55542
g55287 and n55246_not n55542 ; n55543
g55288 and n55541_not n55543_not ; n55544
g55289 and b[29]_not n55544_not ; n55545
g55290 and n54709_not n55063 ; n55546
g55291 and n55059_not n55546 ; n55547
g55292 and n55060_not n55063_not ; n55548
g55293 and n55547_not n55548_not ; n55549
g55294 and n55248_not n55549_not ; n55550
g55295 and n54699_not n55247_not ; n55551
g55296 and n55246_not n55551 ; n55552
g55297 and n55550_not n55552_not ; n55553
g55298 and b[28]_not n55553_not ; n55554
g55299 and n54718_not n55058 ; n55555
g55300 and n55054_not n55555 ; n55556
g55301 and n55055_not n55058_not ; n55557
g55302 and n55556_not n55557_not ; n55558
g55303 and n55248_not n55558_not ; n55559
g55304 and n54708_not n55247_not ; n55560
g55305 and n55246_not n55560 ; n55561
g55306 and n55559_not n55561_not ; n55562
g55307 and b[27]_not n55562_not ; n55563
g55308 and n54727_not n55053 ; n55564
g55309 and n55049_not n55564 ; n55565
g55310 and n55050_not n55053_not ; n55566
g55311 and n55565_not n55566_not ; n55567
g55312 and n55248_not n55567_not ; n55568
g55313 and n54717_not n55247_not ; n55569
g55314 and n55246_not n55569 ; n55570
g55315 and n55568_not n55570_not ; n55571
g55316 and b[26]_not n55571_not ; n55572
g55317 and n54736_not n55048 ; n55573
g55318 and n55044_not n55573 ; n55574
g55319 and n55045_not n55048_not ; n55575
g55320 and n55574_not n55575_not ; n55576
g55321 and n55248_not n55576_not ; n55577
g55322 and n54726_not n55247_not ; n55578
g55323 and n55246_not n55578 ; n55579
g55324 and n55577_not n55579_not ; n55580
g55325 and b[25]_not n55580_not ; n55581
g55326 and n54745_not n55043 ; n55582
g55327 and n55039_not n55582 ; n55583
g55328 and n55040_not n55043_not ; n55584
g55329 and n55583_not n55584_not ; n55585
g55330 and n55248_not n55585_not ; n55586
g55331 and n54735_not n55247_not ; n55587
g55332 and n55246_not n55587 ; n55588
g55333 and n55586_not n55588_not ; n55589
g55334 and b[24]_not n55589_not ; n55590
g55335 and n54754_not n55038 ; n55591
g55336 and n55034_not n55591 ; n55592
g55337 and n55035_not n55038_not ; n55593
g55338 and n55592_not n55593_not ; n55594
g55339 and n55248_not n55594_not ; n55595
g55340 and n54744_not n55247_not ; n55596
g55341 and n55246_not n55596 ; n55597
g55342 and n55595_not n55597_not ; n55598
g55343 and b[23]_not n55598_not ; n55599
g55344 and n54763_not n55033 ; n55600
g55345 and n55029_not n55600 ; n55601
g55346 and n55030_not n55033_not ; n55602
g55347 and n55601_not n55602_not ; n55603
g55348 and n55248_not n55603_not ; n55604
g55349 and n54753_not n55247_not ; n55605
g55350 and n55246_not n55605 ; n55606
g55351 and n55604_not n55606_not ; n55607
g55352 and b[22]_not n55607_not ; n55608
g55353 and n54772_not n55028 ; n55609
g55354 and n55024_not n55609 ; n55610
g55355 and n55025_not n55028_not ; n55611
g55356 and n55610_not n55611_not ; n55612
g55357 and n55248_not n55612_not ; n55613
g55358 and n54762_not n55247_not ; n55614
g55359 and n55246_not n55614 ; n55615
g55360 and n55613_not n55615_not ; n55616
g55361 and b[21]_not n55616_not ; n55617
g55362 and n54781_not n55023 ; n55618
g55363 and n55019_not n55618 ; n55619
g55364 and n55020_not n55023_not ; n55620
g55365 and n55619_not n55620_not ; n55621
g55366 and n55248_not n55621_not ; n55622
g55367 and n54771_not n55247_not ; n55623
g55368 and n55246_not n55623 ; n55624
g55369 and n55622_not n55624_not ; n55625
g55370 and b[20]_not n55625_not ; n55626
g55371 and n54790_not n55018 ; n55627
g55372 and n55014_not n55627 ; n55628
g55373 and n55015_not n55018_not ; n55629
g55374 and n55628_not n55629_not ; n55630
g55375 and n55248_not n55630_not ; n55631
g55376 and n54780_not n55247_not ; n55632
g55377 and n55246_not n55632 ; n55633
g55378 and n55631_not n55633_not ; n55634
g55379 and b[19]_not n55634_not ; n55635
g55380 and n54799_not n55013 ; n55636
g55381 and n55009_not n55636 ; n55637
g55382 and n55010_not n55013_not ; n55638
g55383 and n55637_not n55638_not ; n55639
g55384 and n55248_not n55639_not ; n55640
g55385 and n54789_not n55247_not ; n55641
g55386 and n55246_not n55641 ; n55642
g55387 and n55640_not n55642_not ; n55643
g55388 and b[18]_not n55643_not ; n55644
g55389 and n54808_not n55008 ; n55645
g55390 and n55004_not n55645 ; n55646
g55391 and n55005_not n55008_not ; n55647
g55392 and n55646_not n55647_not ; n55648
g55393 and n55248_not n55648_not ; n55649
g55394 and n54798_not n55247_not ; n55650
g55395 and n55246_not n55650 ; n55651
g55396 and n55649_not n55651_not ; n55652
g55397 and b[17]_not n55652_not ; n55653
g55398 and n54817_not n55003 ; n55654
g55399 and n54999_not n55654 ; n55655
g55400 and n55000_not n55003_not ; n55656
g55401 and n55655_not n55656_not ; n55657
g55402 and n55248_not n55657_not ; n55658
g55403 and n54807_not n55247_not ; n55659
g55404 and n55246_not n55659 ; n55660
g55405 and n55658_not n55660_not ; n55661
g55406 and b[16]_not n55661_not ; n55662
g55407 and n54826_not n54998 ; n55663
g55408 and n54994_not n55663 ; n55664
g55409 and n54995_not n54998_not ; n55665
g55410 and n55664_not n55665_not ; n55666
g55411 and n55248_not n55666_not ; n55667
g55412 and n54816_not n55247_not ; n55668
g55413 and n55246_not n55668 ; n55669
g55414 and n55667_not n55669_not ; n55670
g55415 and b[15]_not n55670_not ; n55671
g55416 and n54835_not n54993 ; n55672
g55417 and n54989_not n55672 ; n55673
g55418 and n54990_not n54993_not ; n55674
g55419 and n55673_not n55674_not ; n55675
g55420 and n55248_not n55675_not ; n55676
g55421 and n54825_not n55247_not ; n55677
g55422 and n55246_not n55677 ; n55678
g55423 and n55676_not n55678_not ; n55679
g55424 and b[14]_not n55679_not ; n55680
g55425 and n54844_not n54988 ; n55681
g55426 and n54984_not n55681 ; n55682
g55427 and n54985_not n54988_not ; n55683
g55428 and n55682_not n55683_not ; n55684
g55429 and n55248_not n55684_not ; n55685
g55430 and n54834_not n55247_not ; n55686
g55431 and n55246_not n55686 ; n55687
g55432 and n55685_not n55687_not ; n55688
g55433 and b[13]_not n55688_not ; n55689
g55434 and n54853_not n54983 ; n55690
g55435 and n54979_not n55690 ; n55691
g55436 and n54980_not n54983_not ; n55692
g55437 and n55691_not n55692_not ; n55693
g55438 and n55248_not n55693_not ; n55694
g55439 and n54843_not n55247_not ; n55695
g55440 and n55246_not n55695 ; n55696
g55441 and n55694_not n55696_not ; n55697
g55442 and b[12]_not n55697_not ; n55698
g55443 and n54862_not n54978 ; n55699
g55444 and n54974_not n55699 ; n55700
g55445 and n54975_not n54978_not ; n55701
g55446 and n55700_not n55701_not ; n55702
g55447 and n55248_not n55702_not ; n55703
g55448 and n54852_not n55247_not ; n55704
g55449 and n55246_not n55704 ; n55705
g55450 and n55703_not n55705_not ; n55706
g55451 and b[11]_not n55706_not ; n55707
g55452 and n54871_not n54973 ; n55708
g55453 and n54969_not n55708 ; n55709
g55454 and n54970_not n54973_not ; n55710
g55455 and n55709_not n55710_not ; n55711
g55456 and n55248_not n55711_not ; n55712
g55457 and n54861_not n55247_not ; n55713
g55458 and n55246_not n55713 ; n55714
g55459 and n55712_not n55714_not ; n55715
g55460 and b[10]_not n55715_not ; n55716
g55461 and n54880_not n54968 ; n55717
g55462 and n54964_not n55717 ; n55718
g55463 and n54965_not n54968_not ; n55719
g55464 and n55718_not n55719_not ; n55720
g55465 and n55248_not n55720_not ; n55721
g55466 and n54870_not n55247_not ; n55722
g55467 and n55246_not n55722 ; n55723
g55468 and n55721_not n55723_not ; n55724
g55469 and b[9]_not n55724_not ; n55725
g55470 and n54889_not n54963 ; n55726
g55471 and n54959_not n55726 ; n55727
g55472 and n54960_not n54963_not ; n55728
g55473 and n55727_not n55728_not ; n55729
g55474 and n55248_not n55729_not ; n55730
g55475 and n54879_not n55247_not ; n55731
g55476 and n55246_not n55731 ; n55732
g55477 and n55730_not n55732_not ; n55733
g55478 and b[8]_not n55733_not ; n55734
g55479 and n54898_not n54958 ; n55735
g55480 and n54954_not n55735 ; n55736
g55481 and n54955_not n54958_not ; n55737
g55482 and n55736_not n55737_not ; n55738
g55483 and n55248_not n55738_not ; n55739
g55484 and n54888_not n55247_not ; n55740
g55485 and n55246_not n55740 ; n55741
g55486 and n55739_not n55741_not ; n55742
g55487 and b[7]_not n55742_not ; n55743
g55488 and n54907_not n54953 ; n55744
g55489 and n54949_not n55744 ; n55745
g55490 and n54950_not n54953_not ; n55746
g55491 and n55745_not n55746_not ; n55747
g55492 and n55248_not n55747_not ; n55748
g55493 and n54897_not n55247_not ; n55749
g55494 and n55246_not n55749 ; n55750
g55495 and n55748_not n55750_not ; n55751
g55496 and b[6]_not n55751_not ; n55752
g55497 and n54916_not n54948 ; n55753
g55498 and n54944_not n55753 ; n55754
g55499 and n54945_not n54948_not ; n55755
g55500 and n55754_not n55755_not ; n55756
g55501 and n55248_not n55756_not ; n55757
g55502 and n54906_not n55247_not ; n55758
g55503 and n55246_not n55758 ; n55759
g55504 and n55757_not n55759_not ; n55760
g55505 and b[5]_not n55760_not ; n55761
g55506 and n54924_not n54943 ; n55762
g55507 and n54939_not n55762 ; n55763
g55508 and n54940_not n54943_not ; n55764
g55509 and n55763_not n55764_not ; n55765
g55510 and n55248_not n55765_not ; n55766
g55511 and n54915_not n55247_not ; n55767
g55512 and n55246_not n55767 ; n55768
g55513 and n55766_not n55768_not ; n55769
g55514 and b[4]_not n55769_not ; n55770
g55515 and n54934_not n54938 ; n55771
g55516 and n54933_not n55771 ; n55772
g55517 and n54935_not n54938_not ; n55773
g55518 and n55772_not n55773_not ; n55774
g55519 and n55248_not n55774_not ; n55775
g55520 and n54923_not n55247_not ; n55776
g55521 and n55246_not n55776 ; n55777
g55522 and n55775_not n55777_not ; n55778
g55523 and b[3]_not n55778_not ; n55779
g55524 and n26919 n54931_not ; n55780
g55525 and n54929_not n55780 ; n55781
g55526 and n54933_not n55781_not ; n55782
g55527 and n55248_not n55782 ; n55783
g55528 and n54928_not n55247_not ; n55784
g55529 and n55246_not n55784 ; n55785
g55530 and n55783_not n55785_not ; n55786
g55531 and b[2]_not n55786_not ; n55787
g55532 and b[0] n55248_not ; n55788
g55533 and a[2] n55788_not ; n55789
g55534 and n26919 n55248_not ; n55790
g55535 and n55789_not n55790_not ; n55791
g55536 and b[1] n55791_not ; n55792
g55537 and b[1]_not n55790_not ; n55793
g55538 and n55789_not n55793 ; n55794
g55539 and n55792_not n55794_not ; n55795
g55540 and n27783_not n55795_not ; n55796
g55541 and b[1]_not n55791_not ; n55797
g55542 and n55796_not n55797_not ; n55798
g55543 and b[2] n55785_not ; n55799
g55544 and n55783_not n55799 ; n55800
g55545 and n55787_not n55800_not ; n55801
g55546 and n55798_not n55801 ; n55802
g55547 and n55787_not n55802_not ; n55803
g55548 and b[3] n55777_not ; n55804
g55549 and n55775_not n55804 ; n55805
g55550 and n55779_not n55805_not ; n55806
g55551 and n55803_not n55806 ; n55807
g55552 and n55779_not n55807_not ; n55808
g55553 and b[4] n55768_not ; n55809
g55554 and n55766_not n55809 ; n55810
g55555 and n55770_not n55810_not ; n55811
g55556 and n55808_not n55811 ; n55812
g55557 and n55770_not n55812_not ; n55813
g55558 and b[5] n55759_not ; n55814
g55559 and n55757_not n55814 ; n55815
g55560 and n55761_not n55815_not ; n55816
g55561 and n55813_not n55816 ; n55817
g55562 and n55761_not n55817_not ; n55818
g55563 and b[6] n55750_not ; n55819
g55564 and n55748_not n55819 ; n55820
g55565 and n55752_not n55820_not ; n55821
g55566 and n55818_not n55821 ; n55822
g55567 and n55752_not n55822_not ; n55823
g55568 and b[7] n55741_not ; n55824
g55569 and n55739_not n55824 ; n55825
g55570 and n55743_not n55825_not ; n55826
g55571 and n55823_not n55826 ; n55827
g55572 and n55743_not n55827_not ; n55828
g55573 and b[8] n55732_not ; n55829
g55574 and n55730_not n55829 ; n55830
g55575 and n55734_not n55830_not ; n55831
g55576 and n55828_not n55831 ; n55832
g55577 and n55734_not n55832_not ; n55833
g55578 and b[9] n55723_not ; n55834
g55579 and n55721_not n55834 ; n55835
g55580 and n55725_not n55835_not ; n55836
g55581 and n55833_not n55836 ; n55837
g55582 and n55725_not n55837_not ; n55838
g55583 and b[10] n55714_not ; n55839
g55584 and n55712_not n55839 ; n55840
g55585 and n55716_not n55840_not ; n55841
g55586 and n55838_not n55841 ; n55842
g55587 and n55716_not n55842_not ; n55843
g55588 and b[11] n55705_not ; n55844
g55589 and n55703_not n55844 ; n55845
g55590 and n55707_not n55845_not ; n55846
g55591 and n55843_not n55846 ; n55847
g55592 and n55707_not n55847_not ; n55848
g55593 and b[12] n55696_not ; n55849
g55594 and n55694_not n55849 ; n55850
g55595 and n55698_not n55850_not ; n55851
g55596 and n55848_not n55851 ; n55852
g55597 and n55698_not n55852_not ; n55853
g55598 and b[13] n55687_not ; n55854
g55599 and n55685_not n55854 ; n55855
g55600 and n55689_not n55855_not ; n55856
g55601 and n55853_not n55856 ; n55857
g55602 and n55689_not n55857_not ; n55858
g55603 and b[14] n55678_not ; n55859
g55604 and n55676_not n55859 ; n55860
g55605 and n55680_not n55860_not ; n55861
g55606 and n55858_not n55861 ; n55862
g55607 and n55680_not n55862_not ; n55863
g55608 and b[15] n55669_not ; n55864
g55609 and n55667_not n55864 ; n55865
g55610 and n55671_not n55865_not ; n55866
g55611 and n55863_not n55866 ; n55867
g55612 and n55671_not n55867_not ; n55868
g55613 and b[16] n55660_not ; n55869
g55614 and n55658_not n55869 ; n55870
g55615 and n55662_not n55870_not ; n55871
g55616 and n55868_not n55871 ; n55872
g55617 and n55662_not n55872_not ; n55873
g55618 and b[17] n55651_not ; n55874
g55619 and n55649_not n55874 ; n55875
g55620 and n55653_not n55875_not ; n55876
g55621 and n55873_not n55876 ; n55877
g55622 and n55653_not n55877_not ; n55878
g55623 and b[18] n55642_not ; n55879
g55624 and n55640_not n55879 ; n55880
g55625 and n55644_not n55880_not ; n55881
g55626 and n55878_not n55881 ; n55882
g55627 and n55644_not n55882_not ; n55883
g55628 and b[19] n55633_not ; n55884
g55629 and n55631_not n55884 ; n55885
g55630 and n55635_not n55885_not ; n55886
g55631 and n55883_not n55886 ; n55887
g55632 and n55635_not n55887_not ; n55888
g55633 and b[20] n55624_not ; n55889
g55634 and n55622_not n55889 ; n55890
g55635 and n55626_not n55890_not ; n55891
g55636 and n55888_not n55891 ; n55892
g55637 and n55626_not n55892_not ; n55893
g55638 and b[21] n55615_not ; n55894
g55639 and n55613_not n55894 ; n55895
g55640 and n55617_not n55895_not ; n55896
g55641 and n55893_not n55896 ; n55897
g55642 and n55617_not n55897_not ; n55898
g55643 and b[22] n55606_not ; n55899
g55644 and n55604_not n55899 ; n55900
g55645 and n55608_not n55900_not ; n55901
g55646 and n55898_not n55901 ; n55902
g55647 and n55608_not n55902_not ; n55903
g55648 and b[23] n55597_not ; n55904
g55649 and n55595_not n55904 ; n55905
g55650 and n55599_not n55905_not ; n55906
g55651 and n55903_not n55906 ; n55907
g55652 and n55599_not n55907_not ; n55908
g55653 and b[24] n55588_not ; n55909
g55654 and n55586_not n55909 ; n55910
g55655 and n55590_not n55910_not ; n55911
g55656 and n55908_not n55911 ; n55912
g55657 and n55590_not n55912_not ; n55913
g55658 and b[25] n55579_not ; n55914
g55659 and n55577_not n55914 ; n55915
g55660 and n55581_not n55915_not ; n55916
g55661 and n55913_not n55916 ; n55917
g55662 and n55581_not n55917_not ; n55918
g55663 and b[26] n55570_not ; n55919
g55664 and n55568_not n55919 ; n55920
g55665 and n55572_not n55920_not ; n55921
g55666 and n55918_not n55921 ; n55922
g55667 and n55572_not n55922_not ; n55923
g55668 and b[27] n55561_not ; n55924
g55669 and n55559_not n55924 ; n55925
g55670 and n55563_not n55925_not ; n55926
g55671 and n55923_not n55926 ; n55927
g55672 and n55563_not n55927_not ; n55928
g55673 and b[28] n55552_not ; n55929
g55674 and n55550_not n55929 ; n55930
g55675 and n55554_not n55930_not ; n55931
g55676 and n55928_not n55931 ; n55932
g55677 and n55554_not n55932_not ; n55933
g55678 and b[29] n55543_not ; n55934
g55679 and n55541_not n55934 ; n55935
g55680 and n55545_not n55935_not ; n55936
g55681 and n55933_not n55936 ; n55937
g55682 and n55545_not n55937_not ; n55938
g55683 and b[30] n55534_not ; n55939
g55684 and n55532_not n55939 ; n55940
g55685 and n55536_not n55940_not ; n55941
g55686 and n55938_not n55941 ; n55942
g55687 and n55536_not n55942_not ; n55943
g55688 and b[31] n55525_not ; n55944
g55689 and n55523_not n55944 ; n55945
g55690 and n55527_not n55945_not ; n55946
g55691 and n55943_not n55946 ; n55947
g55692 and n55527_not n55947_not ; n55948
g55693 and b[32] n55516_not ; n55949
g55694 and n55514_not n55949 ; n55950
g55695 and n55518_not n55950_not ; n55951
g55696 and n55948_not n55951 ; n55952
g55697 and n55518_not n55952_not ; n55953
g55698 and b[33] n55507_not ; n55954
g55699 and n55505_not n55954 ; n55955
g55700 and n55509_not n55955_not ; n55956
g55701 and n55953_not n55956 ; n55957
g55702 and n55509_not n55957_not ; n55958
g55703 and b[34] n55498_not ; n55959
g55704 and n55496_not n55959 ; n55960
g55705 and n55500_not n55960_not ; n55961
g55706 and n55958_not n55961 ; n55962
g55707 and n55500_not n55962_not ; n55963
g55708 and b[35] n55489_not ; n55964
g55709 and n55487_not n55964 ; n55965
g55710 and n55491_not n55965_not ; n55966
g55711 and n55963_not n55966 ; n55967
g55712 and n55491_not n55967_not ; n55968
g55713 and b[36] n55480_not ; n55969
g55714 and n55478_not n55969 ; n55970
g55715 and n55482_not n55970_not ; n55971
g55716 and n55968_not n55971 ; n55972
g55717 and n55482_not n55972_not ; n55973
g55718 and b[37] n55471_not ; n55974
g55719 and n55469_not n55974 ; n55975
g55720 and n55473_not n55975_not ; n55976
g55721 and n55973_not n55976 ; n55977
g55722 and n55473_not n55977_not ; n55978
g55723 and b[38] n55462_not ; n55979
g55724 and n55460_not n55979 ; n55980
g55725 and n55464_not n55980_not ; n55981
g55726 and n55978_not n55981 ; n55982
g55727 and n55464_not n55982_not ; n55983
g55728 and b[39] n55453_not ; n55984
g55729 and n55451_not n55984 ; n55985
g55730 and n55455_not n55985_not ; n55986
g55731 and n55983_not n55986 ; n55987
g55732 and n55455_not n55987_not ; n55988
g55733 and b[40] n55444_not ; n55989
g55734 and n55442_not n55989 ; n55990
g55735 and n55446_not n55990_not ; n55991
g55736 and n55988_not n55991 ; n55992
g55737 and n55446_not n55992_not ; n55993
g55738 and b[41] n55435_not ; n55994
g55739 and n55433_not n55994 ; n55995
g55740 and n55437_not n55995_not ; n55996
g55741 and n55993_not n55996 ; n55997
g55742 and n55437_not n55997_not ; n55998
g55743 and b[42] n55426_not ; n55999
g55744 and n55424_not n55999 ; n56000
g55745 and n55428_not n56000_not ; n56001
g55746 and n55998_not n56001 ; n56002
g55747 and n55428_not n56002_not ; n56003
g55748 and b[43] n55417_not ; n56004
g55749 and n55415_not n56004 ; n56005
g55750 and n55419_not n56005_not ; n56006
g55751 and n56003_not n56006 ; n56007
g55752 and n55419_not n56007_not ; n56008
g55753 and b[44] n55408_not ; n56009
g55754 and n55406_not n56009 ; n56010
g55755 and n55410_not n56010_not ; n56011
g55756 and n56008_not n56011 ; n56012
g55757 and n55410_not n56012_not ; n56013
g55758 and b[45] n55399_not ; n56014
g55759 and n55397_not n56014 ; n56015
g55760 and n55401_not n56015_not ; n56016
g55761 and n56013_not n56016 ; n56017
g55762 and n55401_not n56017_not ; n56018
g55763 and b[46] n55390_not ; n56019
g55764 and n55388_not n56019 ; n56020
g55765 and n55392_not n56020_not ; n56021
g55766 and n56018_not n56021 ; n56022
g55767 and n55392_not n56022_not ; n56023
g55768 and b[47] n55381_not ; n56024
g55769 and n55379_not n56024 ; n56025
g55770 and n55383_not n56025_not ; n56026
g55771 and n56023_not n56026 ; n56027
g55772 and n55383_not n56027_not ; n56028
g55773 and b[48] n55372_not ; n56029
g55774 and n55370_not n56029 ; n56030
g55775 and n55374_not n56030_not ; n56031
g55776 and n56028_not n56031 ; n56032
g55777 and n55374_not n56032_not ; n56033
g55778 and b[49] n55363_not ; n56034
g55779 and n55361_not n56034 ; n56035
g55780 and n55365_not n56035_not ; n56036
g55781 and n56033_not n56036 ; n56037
g55782 and n55365_not n56037_not ; n56038
g55783 and b[50] n55354_not ; n56039
g55784 and n55352_not n56039 ; n56040
g55785 and n55356_not n56040_not ; n56041
g55786 and n56038_not n56041 ; n56042
g55787 and n55356_not n56042_not ; n56043
g55788 and b[51] n55345_not ; n56044
g55789 and n55343_not n56044 ; n56045
g55790 and n55347_not n56045_not ; n56046
g55791 and n56043_not n56046 ; n56047
g55792 and n55347_not n56047_not ; n56048
g55793 and b[52] n55336_not ; n56049
g55794 and n55334_not n56049 ; n56050
g55795 and n55338_not n56050_not ; n56051
g55796 and n56048_not n56051 ; n56052
g55797 and n55338_not n56052_not ; n56053
g55798 and b[53] n55327_not ; n56054
g55799 and n55325_not n56054 ; n56055
g55800 and n55329_not n56055_not ; n56056
g55801 and n56053_not n56056 ; n56057
g55802 and n55329_not n56057_not ; n56058
g55803 and b[54] n55318_not ; n56059
g55804 and n55316_not n56059 ; n56060
g55805 and n55320_not n56060_not ; n56061
g55806 and n56058_not n56061 ; n56062
g55807 and n55320_not n56062_not ; n56063
g55808 and b[55] n55309_not ; n56064
g55809 and n55307_not n56064 ; n56065
g55810 and n55311_not n56065_not ; n56066
g55811 and n56063_not n56066 ; n56067
g55812 and n55311_not n56067_not ; n56068
g55813 and b[56] n55300_not ; n56069
g55814 and n55298_not n56069 ; n56070
g55815 and n55302_not n56070_not ; n56071
g55816 and n56068_not n56071 ; n56072
g55817 and n55302_not n56072_not ; n56073
g55818 and b[57] n55291_not ; n56074
g55819 and n55289_not n56074 ; n56075
g55820 and n55293_not n56075_not ; n56076
g55821 and n56073_not n56076 ; n56077
g55822 and n55293_not n56077_not ; n56078
g55823 and b[58] n55282_not ; n56079
g55824 and n55280_not n56079 ; n56080
g55825 and n55284_not n56080_not ; n56081
g55826 and n56078_not n56081 ; n56082
g55827 and n55284_not n56082_not ; n56083
g55828 and b[59] n55273_not ; n56084
g55829 and n55271_not n56084 ; n56085
g55830 and n55275_not n56085_not ; n56086
g55831 and n56083_not n56086 ; n56087
g55832 and n55275_not n56087_not ; n56088
g55833 and b[60] n55264_not ; n56089
g55834 and n55262_not n56089 ; n56090
g55835 and n55266_not n56090_not ; n56091
g55836 and n56088_not n56091 ; n56092
g55837 and n55266_not n56092_not ; n56093
g55838 and b[61] n55255_not ; n56094
g55839 and n55253_not n56094 ; n56095
g55840 and n55257_not n56095_not ; n56096
g55841 and n56093_not n56096 ; n56097
g55842 and n55257_not n56097_not ; n56098
g55843 and n54403_not n55243_not ; n56099
g55844 and n55241_not n56099 ; n56100
g55845 and n55229_not n56100 ; n56101
g55846 and n55241_not n55243_not ; n56102
g55847 and n55230_not n56102_not ; n56103
g55848 and n56101_not n56103_not ; n56104
g55849 and n55248_not n56104_not ; n56105
g55850 and n55240_not n55247_not ; n56106
g55851 and n55246_not n56106 ; n56107
g55852 and n56105_not n56107_not ; n56108
g55853 and b[62]_not n56108_not ; n56109
g55854 and b[62] n56107_not ; n56110
g55855 and n56105_not n56110 ; n56111
g55856 and b[63]_not n56111_not ; n56112
g55857 and n56109_not n56112 ; n56113
g55858 and n56098_not n56113 ; n56114
g55859 and n279 n56108_not ; n56115
g55860 and n56114_not n56115_not ; n56116
g55861 and n55257_not n56111_not ; n56117
g55862 and n56109_not n56117 ; n56118
g55863 and n56097_not n56118 ; n56119
g55864 and n56109_not n56111_not ; n56120
g55865 and n56098_not n56120_not ; n56121
g55866 and n56119_not n56121_not ; n56122
g55867 and n56116_not n56122_not ; n56123
g55868 and n56108_not n56115_not ; n56124
g55869 and n56114_not n56124 ; n56125
g55870 and n56123_not n56125_not ; n56126
g55871 and b[63]_not n56126_not ; n56127
g55872 and n55266_not n56096 ; n56128
g55873 and n56092_not n56128 ; n56129
g55874 and n56093_not n56096_not ; n56130
g55875 and n56129_not n56130_not ; n56131
g55876 and n56116_not n56131_not ; n56132
g55877 and n55256_not n56115_not ; n56133
g55878 and n56114_not n56133 ; n56134
g55879 and n56132_not n56134_not ; n56135
g55880 and b[62]_not n56135_not ; n56136
g55881 and n55275_not n56091 ; n56137
g55882 and n56087_not n56137 ; n56138
g55883 and n56088_not n56091_not ; n56139
g55884 and n56138_not n56139_not ; n56140
g55885 and n56116_not n56140_not ; n56141
g55886 and n55265_not n56115_not ; n56142
g55887 and n56114_not n56142 ; n56143
g55888 and n56141_not n56143_not ; n56144
g55889 and b[61]_not n56144_not ; n56145
g55890 and n55284_not n56086 ; n56146
g55891 and n56082_not n56146 ; n56147
g55892 and n56083_not n56086_not ; n56148
g55893 and n56147_not n56148_not ; n56149
g55894 and n56116_not n56149_not ; n56150
g55895 and n55274_not n56115_not ; n56151
g55896 and n56114_not n56151 ; n56152
g55897 and n56150_not n56152_not ; n56153
g55898 and b[60]_not n56153_not ; n56154
g55899 and n55293_not n56081 ; n56155
g55900 and n56077_not n56155 ; n56156
g55901 and n56078_not n56081_not ; n56157
g55902 and n56156_not n56157_not ; n56158
g55903 and n56116_not n56158_not ; n56159
g55904 and n55283_not n56115_not ; n56160
g55905 and n56114_not n56160 ; n56161
g55906 and n56159_not n56161_not ; n56162
g55907 and b[59]_not n56162_not ; n56163
g55908 and n55302_not n56076 ; n56164
g55909 and n56072_not n56164 ; n56165
g55910 and n56073_not n56076_not ; n56166
g55911 and n56165_not n56166_not ; n56167
g55912 and n56116_not n56167_not ; n56168
g55913 and n55292_not n56115_not ; n56169
g55914 and n56114_not n56169 ; n56170
g55915 and n56168_not n56170_not ; n56171
g55916 and b[58]_not n56171_not ; n56172
g55917 and n55311_not n56071 ; n56173
g55918 and n56067_not n56173 ; n56174
g55919 and n56068_not n56071_not ; n56175
g55920 and n56174_not n56175_not ; n56176
g55921 and n56116_not n56176_not ; n56177
g55922 and n55301_not n56115_not ; n56178
g55923 and n56114_not n56178 ; n56179
g55924 and n56177_not n56179_not ; n56180
g55925 and b[57]_not n56180_not ; n56181
g55926 and n55320_not n56066 ; n56182
g55927 and n56062_not n56182 ; n56183
g55928 and n56063_not n56066_not ; n56184
g55929 and n56183_not n56184_not ; n56185
g55930 and n56116_not n56185_not ; n56186
g55931 and n55310_not n56115_not ; n56187
g55932 and n56114_not n56187 ; n56188
g55933 and n56186_not n56188_not ; n56189
g55934 and b[56]_not n56189_not ; n56190
g55935 and n55329_not n56061 ; n56191
g55936 and n56057_not n56191 ; n56192
g55937 and n56058_not n56061_not ; n56193
g55938 and n56192_not n56193_not ; n56194
g55939 and n56116_not n56194_not ; n56195
g55940 and n55319_not n56115_not ; n56196
g55941 and n56114_not n56196 ; n56197
g55942 and n56195_not n56197_not ; n56198
g55943 and b[55]_not n56198_not ; n56199
g55944 and n55338_not n56056 ; n56200
g55945 and n56052_not n56200 ; n56201
g55946 and n56053_not n56056_not ; n56202
g55947 and n56201_not n56202_not ; n56203
g55948 and n56116_not n56203_not ; n56204
g55949 and n55328_not n56115_not ; n56205
g55950 and n56114_not n56205 ; n56206
g55951 and n56204_not n56206_not ; n56207
g55952 and b[54]_not n56207_not ; n56208
g55953 and n55347_not n56051 ; n56209
g55954 and n56047_not n56209 ; n56210
g55955 and n56048_not n56051_not ; n56211
g55956 and n56210_not n56211_not ; n56212
g55957 and n56116_not n56212_not ; n56213
g55958 and n55337_not n56115_not ; n56214
g55959 and n56114_not n56214 ; n56215
g55960 and n56213_not n56215_not ; n56216
g55961 and b[53]_not n56216_not ; n56217
g55962 and n55356_not n56046 ; n56218
g55963 and n56042_not n56218 ; n56219
g55964 and n56043_not n56046_not ; n56220
g55965 and n56219_not n56220_not ; n56221
g55966 and n56116_not n56221_not ; n56222
g55967 and n55346_not n56115_not ; n56223
g55968 and n56114_not n56223 ; n56224
g55969 and n56222_not n56224_not ; n56225
g55970 and b[52]_not n56225_not ; n56226
g55971 and n55365_not n56041 ; n56227
g55972 and n56037_not n56227 ; n56228
g55973 and n56038_not n56041_not ; n56229
g55974 and n56228_not n56229_not ; n56230
g55975 and n56116_not n56230_not ; n56231
g55976 and n55355_not n56115_not ; n56232
g55977 and n56114_not n56232 ; n56233
g55978 and n56231_not n56233_not ; n56234
g55979 and b[51]_not n56234_not ; n56235
g55980 and n55374_not n56036 ; n56236
g55981 and n56032_not n56236 ; n56237
g55982 and n56033_not n56036_not ; n56238
g55983 and n56237_not n56238_not ; n56239
g55984 and n56116_not n56239_not ; n56240
g55985 and n55364_not n56115_not ; n56241
g55986 and n56114_not n56241 ; n56242
g55987 and n56240_not n56242_not ; n56243
g55988 and b[50]_not n56243_not ; n56244
g55989 and n55383_not n56031 ; n56245
g55990 and n56027_not n56245 ; n56246
g55991 and n56028_not n56031_not ; n56247
g55992 and n56246_not n56247_not ; n56248
g55993 and n56116_not n56248_not ; n56249
g55994 and n55373_not n56115_not ; n56250
g55995 and n56114_not n56250 ; n56251
g55996 and n56249_not n56251_not ; n56252
g55997 and b[49]_not n56252_not ; n56253
g55998 and n55392_not n56026 ; n56254
g55999 and n56022_not n56254 ; n56255
g56000 and n56023_not n56026_not ; n56256
g56001 and n56255_not n56256_not ; n56257
g56002 and n56116_not n56257_not ; n56258
g56003 and n55382_not n56115_not ; n56259
g56004 and n56114_not n56259 ; n56260
g56005 and n56258_not n56260_not ; n56261
g56006 and b[48]_not n56261_not ; n56262
g56007 and n55401_not n56021 ; n56263
g56008 and n56017_not n56263 ; n56264
g56009 and n56018_not n56021_not ; n56265
g56010 and n56264_not n56265_not ; n56266
g56011 and n56116_not n56266_not ; n56267
g56012 and n55391_not n56115_not ; n56268
g56013 and n56114_not n56268 ; n56269
g56014 and n56267_not n56269_not ; n56270
g56015 and b[47]_not n56270_not ; n56271
g56016 and n55410_not n56016 ; n56272
g56017 and n56012_not n56272 ; n56273
g56018 and n56013_not n56016_not ; n56274
g56019 and n56273_not n56274_not ; n56275
g56020 and n56116_not n56275_not ; n56276
g56021 and n55400_not n56115_not ; n56277
g56022 and n56114_not n56277 ; n56278
g56023 and n56276_not n56278_not ; n56279
g56024 and b[46]_not n56279_not ; n56280
g56025 and n55419_not n56011 ; n56281
g56026 and n56007_not n56281 ; n56282
g56027 and n56008_not n56011_not ; n56283
g56028 and n56282_not n56283_not ; n56284
g56029 and n56116_not n56284_not ; n56285
g56030 and n55409_not n56115_not ; n56286
g56031 and n56114_not n56286 ; n56287
g56032 and n56285_not n56287_not ; n56288
g56033 and b[45]_not n56288_not ; n56289
g56034 and n55428_not n56006 ; n56290
g56035 and n56002_not n56290 ; n56291
g56036 and n56003_not n56006_not ; n56292
g56037 and n56291_not n56292_not ; n56293
g56038 and n56116_not n56293_not ; n56294
g56039 and n55418_not n56115_not ; n56295
g56040 and n56114_not n56295 ; n56296
g56041 and n56294_not n56296_not ; n56297
g56042 and b[44]_not n56297_not ; n56298
g56043 and n55437_not n56001 ; n56299
g56044 and n55997_not n56299 ; n56300
g56045 and n55998_not n56001_not ; n56301
g56046 and n56300_not n56301_not ; n56302
g56047 and n56116_not n56302_not ; n56303
g56048 and n55427_not n56115_not ; n56304
g56049 and n56114_not n56304 ; n56305
g56050 and n56303_not n56305_not ; n56306
g56051 and b[43]_not n56306_not ; n56307
g56052 and n55446_not n55996 ; n56308
g56053 and n55992_not n56308 ; n56309
g56054 and n55993_not n55996_not ; n56310
g56055 and n56309_not n56310_not ; n56311
g56056 and n56116_not n56311_not ; n56312
g56057 and n55436_not n56115_not ; n56313
g56058 and n56114_not n56313 ; n56314
g56059 and n56312_not n56314_not ; n56315
g56060 and b[42]_not n56315_not ; n56316
g56061 and n55455_not n55991 ; n56317
g56062 and n55987_not n56317 ; n56318
g56063 and n55988_not n55991_not ; n56319
g56064 and n56318_not n56319_not ; n56320
g56065 and n56116_not n56320_not ; n56321
g56066 and n55445_not n56115_not ; n56322
g56067 and n56114_not n56322 ; n56323
g56068 and n56321_not n56323_not ; n56324
g56069 and b[41]_not n56324_not ; n56325
g56070 and n55464_not n55986 ; n56326
g56071 and n55982_not n56326 ; n56327
g56072 and n55983_not n55986_not ; n56328
g56073 and n56327_not n56328_not ; n56329
g56074 and n56116_not n56329_not ; n56330
g56075 and n55454_not n56115_not ; n56331
g56076 and n56114_not n56331 ; n56332
g56077 and n56330_not n56332_not ; n56333
g56078 and b[40]_not n56333_not ; n56334
g56079 and n55473_not n55981 ; n56335
g56080 and n55977_not n56335 ; n56336
g56081 and n55978_not n55981_not ; n56337
g56082 and n56336_not n56337_not ; n56338
g56083 and n56116_not n56338_not ; n56339
g56084 and n55463_not n56115_not ; n56340
g56085 and n56114_not n56340 ; n56341
g56086 and n56339_not n56341_not ; n56342
g56087 and b[39]_not n56342_not ; n56343
g56088 and n55482_not n55976 ; n56344
g56089 and n55972_not n56344 ; n56345
g56090 and n55973_not n55976_not ; n56346
g56091 and n56345_not n56346_not ; n56347
g56092 and n56116_not n56347_not ; n56348
g56093 and n55472_not n56115_not ; n56349
g56094 and n56114_not n56349 ; n56350
g56095 and n56348_not n56350_not ; n56351
g56096 and b[38]_not n56351_not ; n56352
g56097 and n55491_not n55971 ; n56353
g56098 and n55967_not n56353 ; n56354
g56099 and n55968_not n55971_not ; n56355
g56100 and n56354_not n56355_not ; n56356
g56101 and n56116_not n56356_not ; n56357
g56102 and n55481_not n56115_not ; n56358
g56103 and n56114_not n56358 ; n56359
g56104 and n56357_not n56359_not ; n56360
g56105 and b[37]_not n56360_not ; n56361
g56106 and n55500_not n55966 ; n56362
g56107 and n55962_not n56362 ; n56363
g56108 and n55963_not n55966_not ; n56364
g56109 and n56363_not n56364_not ; n56365
g56110 and n56116_not n56365_not ; n56366
g56111 and n55490_not n56115_not ; n56367
g56112 and n56114_not n56367 ; n56368
g56113 and n56366_not n56368_not ; n56369
g56114 and b[36]_not n56369_not ; n56370
g56115 and n55509_not n55961 ; n56371
g56116 and n55957_not n56371 ; n56372
g56117 and n55958_not n55961_not ; n56373
g56118 and n56372_not n56373_not ; n56374
g56119 and n56116_not n56374_not ; n56375
g56120 and n55499_not n56115_not ; n56376
g56121 and n56114_not n56376 ; n56377
g56122 and n56375_not n56377_not ; n56378
g56123 and b[35]_not n56378_not ; n56379
g56124 and n55518_not n55956 ; n56380
g56125 and n55952_not n56380 ; n56381
g56126 and n55953_not n55956_not ; n56382
g56127 and n56381_not n56382_not ; n56383
g56128 and n56116_not n56383_not ; n56384
g56129 and n55508_not n56115_not ; n56385
g56130 and n56114_not n56385 ; n56386
g56131 and n56384_not n56386_not ; n56387
g56132 and b[34]_not n56387_not ; n56388
g56133 and n55527_not n55951 ; n56389
g56134 and n55947_not n56389 ; n56390
g56135 and n55948_not n55951_not ; n56391
g56136 and n56390_not n56391_not ; n56392
g56137 and n56116_not n56392_not ; n56393
g56138 and n55517_not n56115_not ; n56394
g56139 and n56114_not n56394 ; n56395
g56140 and n56393_not n56395_not ; n56396
g56141 and b[33]_not n56396_not ; n56397
g56142 and n55536_not n55946 ; n56398
g56143 and n55942_not n56398 ; n56399
g56144 and n55943_not n55946_not ; n56400
g56145 and n56399_not n56400_not ; n56401
g56146 and n56116_not n56401_not ; n56402
g56147 and n55526_not n56115_not ; n56403
g56148 and n56114_not n56403 ; n56404
g56149 and n56402_not n56404_not ; n56405
g56150 and b[32]_not n56405_not ; n56406
g56151 and n55545_not n55941 ; n56407
g56152 and n55937_not n56407 ; n56408
g56153 and n55938_not n55941_not ; n56409
g56154 and n56408_not n56409_not ; n56410
g56155 and n56116_not n56410_not ; n56411
g56156 and n55535_not n56115_not ; n56412
g56157 and n56114_not n56412 ; n56413
g56158 and n56411_not n56413_not ; n56414
g56159 and b[31]_not n56414_not ; n56415
g56160 and n55554_not n55936 ; n56416
g56161 and n55932_not n56416 ; n56417
g56162 and n55933_not n55936_not ; n56418
g56163 and n56417_not n56418_not ; n56419
g56164 and n56116_not n56419_not ; n56420
g56165 and n55544_not n56115_not ; n56421
g56166 and n56114_not n56421 ; n56422
g56167 and n56420_not n56422_not ; n56423
g56168 and b[30]_not n56423_not ; n56424
g56169 and n55563_not n55931 ; n56425
g56170 and n55927_not n56425 ; n56426
g56171 and n55928_not n55931_not ; n56427
g56172 and n56426_not n56427_not ; n56428
g56173 and n56116_not n56428_not ; n56429
g56174 and n55553_not n56115_not ; n56430
g56175 and n56114_not n56430 ; n56431
g56176 and n56429_not n56431_not ; n56432
g56177 and b[29]_not n56432_not ; n56433
g56178 and n55572_not n55926 ; n56434
g56179 and n55922_not n56434 ; n56435
g56180 and n55923_not n55926_not ; n56436
g56181 and n56435_not n56436_not ; n56437
g56182 and n56116_not n56437_not ; n56438
g56183 and n55562_not n56115_not ; n56439
g56184 and n56114_not n56439 ; n56440
g56185 and n56438_not n56440_not ; n56441
g56186 and b[28]_not n56441_not ; n56442
g56187 and n55581_not n55921 ; n56443
g56188 and n55917_not n56443 ; n56444
g56189 and n55918_not n55921_not ; n56445
g56190 and n56444_not n56445_not ; n56446
g56191 and n56116_not n56446_not ; n56447
g56192 and n55571_not n56115_not ; n56448
g56193 and n56114_not n56448 ; n56449
g56194 and n56447_not n56449_not ; n56450
g56195 and b[27]_not n56450_not ; n56451
g56196 and n55590_not n55916 ; n56452
g56197 and n55912_not n56452 ; n56453
g56198 and n55913_not n55916_not ; n56454
g56199 and n56453_not n56454_not ; n56455
g56200 and n56116_not n56455_not ; n56456
g56201 and n55580_not n56115_not ; n56457
g56202 and n56114_not n56457 ; n56458
g56203 and n56456_not n56458_not ; n56459
g56204 and b[26]_not n56459_not ; n56460
g56205 and n55599_not n55911 ; n56461
g56206 and n55907_not n56461 ; n56462
g56207 and n55908_not n55911_not ; n56463
g56208 and n56462_not n56463_not ; n56464
g56209 and n56116_not n56464_not ; n56465
g56210 and n55589_not n56115_not ; n56466
g56211 and n56114_not n56466 ; n56467
g56212 and n56465_not n56467_not ; n56468
g56213 and b[25]_not n56468_not ; n56469
g56214 and n55608_not n55906 ; n56470
g56215 and n55902_not n56470 ; n56471
g56216 and n55903_not n55906_not ; n56472
g56217 and n56471_not n56472_not ; n56473
g56218 and n56116_not n56473_not ; n56474
g56219 and n55598_not n56115_not ; n56475
g56220 and n56114_not n56475 ; n56476
g56221 and n56474_not n56476_not ; n56477
g56222 and b[24]_not n56477_not ; n56478
g56223 and n55617_not n55901 ; n56479
g56224 and n55897_not n56479 ; n56480
g56225 and n55898_not n55901_not ; n56481
g56226 and n56480_not n56481_not ; n56482
g56227 and n56116_not n56482_not ; n56483
g56228 and n55607_not n56115_not ; n56484
g56229 and n56114_not n56484 ; n56485
g56230 and n56483_not n56485_not ; n56486
g56231 and b[23]_not n56486_not ; n56487
g56232 and n55626_not n55896 ; n56488
g56233 and n55892_not n56488 ; n56489
g56234 and n55893_not n55896_not ; n56490
g56235 and n56489_not n56490_not ; n56491
g56236 and n56116_not n56491_not ; n56492
g56237 and n55616_not n56115_not ; n56493
g56238 and n56114_not n56493 ; n56494
g56239 and n56492_not n56494_not ; n56495
g56240 and b[22]_not n56495_not ; n56496
g56241 and n55635_not n55891 ; n56497
g56242 and n55887_not n56497 ; n56498
g56243 and n55888_not n55891_not ; n56499
g56244 and n56498_not n56499_not ; n56500
g56245 and n56116_not n56500_not ; n56501
g56246 and n55625_not n56115_not ; n56502
g56247 and n56114_not n56502 ; n56503
g56248 and n56501_not n56503_not ; n56504
g56249 and b[21]_not n56504_not ; n56505
g56250 and n55644_not n55886 ; n56506
g56251 and n55882_not n56506 ; n56507
g56252 and n55883_not n55886_not ; n56508
g56253 and n56507_not n56508_not ; n56509
g56254 and n56116_not n56509_not ; n56510
g56255 and n55634_not n56115_not ; n56511
g56256 and n56114_not n56511 ; n56512
g56257 and n56510_not n56512_not ; n56513
g56258 and b[20]_not n56513_not ; n56514
g56259 and n55653_not n55881 ; n56515
g56260 and n55877_not n56515 ; n56516
g56261 and n55878_not n55881_not ; n56517
g56262 and n56516_not n56517_not ; n56518
g56263 and n56116_not n56518_not ; n56519
g56264 and n55643_not n56115_not ; n56520
g56265 and n56114_not n56520 ; n56521
g56266 and n56519_not n56521_not ; n56522
g56267 and b[19]_not n56522_not ; n56523
g56268 and n55662_not n55876 ; n56524
g56269 and n55872_not n56524 ; n56525
g56270 and n55873_not n55876_not ; n56526
g56271 and n56525_not n56526_not ; n56527
g56272 and n56116_not n56527_not ; n56528
g56273 and n55652_not n56115_not ; n56529
g56274 and n56114_not n56529 ; n56530
g56275 and n56528_not n56530_not ; n56531
g56276 and b[18]_not n56531_not ; n56532
g56277 and n55671_not n55871 ; n56533
g56278 and n55867_not n56533 ; n56534
g56279 and n55868_not n55871_not ; n56535
g56280 and n56534_not n56535_not ; n56536
g56281 and n56116_not n56536_not ; n56537
g56282 and n55661_not n56115_not ; n56538
g56283 and n56114_not n56538 ; n56539
g56284 and n56537_not n56539_not ; n56540
g56285 and b[17]_not n56540_not ; n56541
g56286 and n55680_not n55866 ; n56542
g56287 and n55862_not n56542 ; n56543
g56288 and n55863_not n55866_not ; n56544
g56289 and n56543_not n56544_not ; n56545
g56290 and n56116_not n56545_not ; n56546
g56291 and n55670_not n56115_not ; n56547
g56292 and n56114_not n56547 ; n56548
g56293 and n56546_not n56548_not ; n56549
g56294 and b[16]_not n56549_not ; n56550
g56295 and n55689_not n55861 ; n56551
g56296 and n55857_not n56551 ; n56552
g56297 and n55858_not n55861_not ; n56553
g56298 and n56552_not n56553_not ; n56554
g56299 and n56116_not n56554_not ; n56555
g56300 and n55679_not n56115_not ; n56556
g56301 and n56114_not n56556 ; n56557
g56302 and n56555_not n56557_not ; n56558
g56303 and b[15]_not n56558_not ; n56559
g56304 and n55698_not n55856 ; n56560
g56305 and n55852_not n56560 ; n56561
g56306 and n55853_not n55856_not ; n56562
g56307 and n56561_not n56562_not ; n56563
g56308 and n56116_not n56563_not ; n56564
g56309 and n55688_not n56115_not ; n56565
g56310 and n56114_not n56565 ; n56566
g56311 and n56564_not n56566_not ; n56567
g56312 and b[14]_not n56567_not ; n56568
g56313 and n55707_not n55851 ; n56569
g56314 and n55847_not n56569 ; n56570
g56315 and n55848_not n55851_not ; n56571
g56316 and n56570_not n56571_not ; n56572
g56317 and n56116_not n56572_not ; n56573
g56318 and n55697_not n56115_not ; n56574
g56319 and n56114_not n56574 ; n56575
g56320 and n56573_not n56575_not ; n56576
g56321 and b[13]_not n56576_not ; n56577
g56322 and n55716_not n55846 ; n56578
g56323 and n55842_not n56578 ; n56579
g56324 and n55843_not n55846_not ; n56580
g56325 and n56579_not n56580_not ; n56581
g56326 and n56116_not n56581_not ; n56582
g56327 and n55706_not n56115_not ; n56583
g56328 and n56114_not n56583 ; n56584
g56329 and n56582_not n56584_not ; n56585
g56330 and b[12]_not n56585_not ; n56586
g56331 and n55725_not n55841 ; n56587
g56332 and n55837_not n56587 ; n56588
g56333 and n55838_not n55841_not ; n56589
g56334 and n56588_not n56589_not ; n56590
g56335 and n56116_not n56590_not ; n56591
g56336 and n55715_not n56115_not ; n56592
g56337 and n56114_not n56592 ; n56593
g56338 and n56591_not n56593_not ; n56594
g56339 and b[11]_not n56594_not ; n56595
g56340 and n55734_not n55836 ; n56596
g56341 and n55832_not n56596 ; n56597
g56342 and n55833_not n55836_not ; n56598
g56343 and n56597_not n56598_not ; n56599
g56344 and n56116_not n56599_not ; n56600
g56345 and n55724_not n56115_not ; n56601
g56346 and n56114_not n56601 ; n56602
g56347 and n56600_not n56602_not ; n56603
g56348 and b[10]_not n56603_not ; n56604
g56349 and n55743_not n55831 ; n56605
g56350 and n55827_not n56605 ; n56606
g56351 and n55828_not n55831_not ; n56607
g56352 and n56606_not n56607_not ; n56608
g56353 and n56116_not n56608_not ; n56609
g56354 and n55733_not n56115_not ; n56610
g56355 and n56114_not n56610 ; n56611
g56356 and n56609_not n56611_not ; n56612
g56357 and b[9]_not n56612_not ; n56613
g56358 and n55752_not n55826 ; n56614
g56359 and n55822_not n56614 ; n56615
g56360 and n55823_not n55826_not ; n56616
g56361 and n56615_not n56616_not ; n56617
g56362 and n56116_not n56617_not ; n56618
g56363 and n55742_not n56115_not ; n56619
g56364 and n56114_not n56619 ; n56620
g56365 and n56618_not n56620_not ; n56621
g56366 and b[8]_not n56621_not ; n56622
g56367 and n55761_not n55821 ; n56623
g56368 and n55817_not n56623 ; n56624
g56369 and n55818_not n55821_not ; n56625
g56370 and n56624_not n56625_not ; n56626
g56371 and n56116_not n56626_not ; n56627
g56372 and n55751_not n56115_not ; n56628
g56373 and n56114_not n56628 ; n56629
g56374 and n56627_not n56629_not ; n56630
g56375 and b[7]_not n56630_not ; n56631
g56376 and n55770_not n55816 ; n56632
g56377 and n55812_not n56632 ; n56633
g56378 and n55813_not n55816_not ; n56634
g56379 and n56633_not n56634_not ; n56635
g56380 and n56116_not n56635_not ; n56636
g56381 and n55760_not n56115_not ; n56637
g56382 and n56114_not n56637 ; n56638
g56383 and n56636_not n56638_not ; n56639
g56384 and b[6]_not n56639_not ; n56640
g56385 and n55779_not n55811 ; n56641
g56386 and n55807_not n56641 ; n56642
g56387 and n55808_not n55811_not ; n56643
g56388 and n56642_not n56643_not ; n56644
g56389 and n56116_not n56644_not ; n56645
g56390 and n55769_not n56115_not ; n56646
g56391 and n56114_not n56646 ; n56647
g56392 and n56645_not n56647_not ; n56648
g56393 and b[5]_not n56648_not ; n56649
g56394 and n55787_not n55806 ; n56650
g56395 and n55802_not n56650 ; n56651
g56396 and n55803_not n55806_not ; n56652
g56397 and n56651_not n56652_not ; n56653
g56398 and n56116_not n56653_not ; n56654
g56399 and n55778_not n56115_not ; n56655
g56400 and n56114_not n56655 ; n56656
g56401 and n56654_not n56656_not ; n56657
g56402 and b[4]_not n56657_not ; n56658
g56403 and n55797_not n55801 ; n56659
g56404 and n55796_not n56659 ; n56660
g56405 and n55798_not n55801_not ; n56661
g56406 and n56660_not n56661_not ; n56662
g56407 and n56116_not n56662_not ; n56663
g56408 and n55786_not n56115_not ; n56664
g56409 and n56114_not n56664 ; n56665
g56410 and n56663_not n56665_not ; n56666
g56411 and b[3]_not n56666_not ; n56667
g56412 and n27783 n55794_not ; n56668
g56413 and n55792_not n56668 ; n56669
g56414 and n55796_not n56669_not ; n56670
g56415 and n56116_not n56670 ; n56671
g56416 and n55791_not n56115_not ; n56672
g56417 and n56114_not n56672 ; n56673
g56418 and n56671_not n56673_not ; n56674
g56419 and b[2]_not n56674_not ; n56675
g56420 and b[0] n56116_not ; n56676
g56421 and a[1] n56676_not ; n56677
g56422 and n27783 n56116_not ; n56678
g56423 and n56677_not n56678_not ; n56679
g56424 and b[1] n56679_not ; n56680
g56425 and b[1]_not n56678_not ; n56681
g56426 and n56677_not n56681 ; n56682
g56427 and n56680_not n56682_not ; n56683
g56428 and n28345_not n56683_not ; n56684
g56429 and b[1]_not n56679_not ; n56685
g56430 and n56684_not n56685_not ; n56686
g56431 and b[2] n56673_not ; n56687
g56432 and n56671_not n56687 ; n56688
g56433 and n56675_not n56688_not ; n56689
g56434 and n56686_not n56689 ; n56690
g56435 and n56675_not n56690_not ; n56691
g56436 and b[3] n56665_not ; n56692
g56437 and n56663_not n56692 ; n56693
g56438 and n56667_not n56693_not ; n56694
g56439 and n56691_not n56694 ; n56695
g56440 and n56667_not n56695_not ; n56696
g56441 and b[4] n56656_not ; n56697
g56442 and n56654_not n56697 ; n56698
g56443 and n56658_not n56698_not ; n56699
g56444 and n56696_not n56699 ; n56700
g56445 and n56658_not n56700_not ; n56701
g56446 and b[5] n56647_not ; n56702
g56447 and n56645_not n56702 ; n56703
g56448 and n56649_not n56703_not ; n56704
g56449 and n56701_not n56704 ; n56705
g56450 and n56649_not n56705_not ; n56706
g56451 and b[6] n56638_not ; n56707
g56452 and n56636_not n56707 ; n56708
g56453 and n56640_not n56708_not ; n56709
g56454 and n56706_not n56709 ; n56710
g56455 and n56640_not n56710_not ; n56711
g56456 and b[7] n56629_not ; n56712
g56457 and n56627_not n56712 ; n56713
g56458 and n56631_not n56713_not ; n56714
g56459 and n56711_not n56714 ; n56715
g56460 and n56631_not n56715_not ; n56716
g56461 and b[8] n56620_not ; n56717
g56462 and n56618_not n56717 ; n56718
g56463 and n56622_not n56718_not ; n56719
g56464 and n56716_not n56719 ; n56720
g56465 and n56622_not n56720_not ; n56721
g56466 and b[9] n56611_not ; n56722
g56467 and n56609_not n56722 ; n56723
g56468 and n56613_not n56723_not ; n56724
g56469 and n56721_not n56724 ; n56725
g56470 and n56613_not n56725_not ; n56726
g56471 and b[10] n56602_not ; n56727
g56472 and n56600_not n56727 ; n56728
g56473 and n56604_not n56728_not ; n56729
g56474 and n56726_not n56729 ; n56730
g56475 and n56604_not n56730_not ; n56731
g56476 and b[11] n56593_not ; n56732
g56477 and n56591_not n56732 ; n56733
g56478 and n56595_not n56733_not ; n56734
g56479 and n56731_not n56734 ; n56735
g56480 and n56595_not n56735_not ; n56736
g56481 and b[12] n56584_not ; n56737
g56482 and n56582_not n56737 ; n56738
g56483 and n56586_not n56738_not ; n56739
g56484 and n56736_not n56739 ; n56740
g56485 and n56586_not n56740_not ; n56741
g56486 and b[13] n56575_not ; n56742
g56487 and n56573_not n56742 ; n56743
g56488 and n56577_not n56743_not ; n56744
g56489 and n56741_not n56744 ; n56745
g56490 and n56577_not n56745_not ; n56746
g56491 and b[14] n56566_not ; n56747
g56492 and n56564_not n56747 ; n56748
g56493 and n56568_not n56748_not ; n56749
g56494 and n56746_not n56749 ; n56750
g56495 and n56568_not n56750_not ; n56751
g56496 and b[15] n56557_not ; n56752
g56497 and n56555_not n56752 ; n56753
g56498 and n56559_not n56753_not ; n56754
g56499 and n56751_not n56754 ; n56755
g56500 and n56559_not n56755_not ; n56756
g56501 and b[16] n56548_not ; n56757
g56502 and n56546_not n56757 ; n56758
g56503 and n56550_not n56758_not ; n56759
g56504 and n56756_not n56759 ; n56760
g56505 and n56550_not n56760_not ; n56761
g56506 and b[17] n56539_not ; n56762
g56507 and n56537_not n56762 ; n56763
g56508 and n56541_not n56763_not ; n56764
g56509 and n56761_not n56764 ; n56765
g56510 and n56541_not n56765_not ; n56766
g56511 and b[18] n56530_not ; n56767
g56512 and n56528_not n56767 ; n56768
g56513 and n56532_not n56768_not ; n56769
g56514 and n56766_not n56769 ; n56770
g56515 and n56532_not n56770_not ; n56771
g56516 and b[19] n56521_not ; n56772
g56517 and n56519_not n56772 ; n56773
g56518 and n56523_not n56773_not ; n56774
g56519 and n56771_not n56774 ; n56775
g56520 and n56523_not n56775_not ; n56776
g56521 and b[20] n56512_not ; n56777
g56522 and n56510_not n56777 ; n56778
g56523 and n56514_not n56778_not ; n56779
g56524 and n56776_not n56779 ; n56780
g56525 and n56514_not n56780_not ; n56781
g56526 and b[21] n56503_not ; n56782
g56527 and n56501_not n56782 ; n56783
g56528 and n56505_not n56783_not ; n56784
g56529 and n56781_not n56784 ; n56785
g56530 and n56505_not n56785_not ; n56786
g56531 and b[22] n56494_not ; n56787
g56532 and n56492_not n56787 ; n56788
g56533 and n56496_not n56788_not ; n56789
g56534 and n56786_not n56789 ; n56790
g56535 and n56496_not n56790_not ; n56791
g56536 and b[23] n56485_not ; n56792
g56537 and n56483_not n56792 ; n56793
g56538 and n56487_not n56793_not ; n56794
g56539 and n56791_not n56794 ; n56795
g56540 and n56487_not n56795_not ; n56796
g56541 and b[24] n56476_not ; n56797
g56542 and n56474_not n56797 ; n56798
g56543 and n56478_not n56798_not ; n56799
g56544 and n56796_not n56799 ; n56800
g56545 and n56478_not n56800_not ; n56801
g56546 and b[25] n56467_not ; n56802
g56547 and n56465_not n56802 ; n56803
g56548 and n56469_not n56803_not ; n56804
g56549 and n56801_not n56804 ; n56805
g56550 and n56469_not n56805_not ; n56806
g56551 and b[26] n56458_not ; n56807
g56552 and n56456_not n56807 ; n56808
g56553 and n56460_not n56808_not ; n56809
g56554 and n56806_not n56809 ; n56810
g56555 and n56460_not n56810_not ; n56811
g56556 and b[27] n56449_not ; n56812
g56557 and n56447_not n56812 ; n56813
g56558 and n56451_not n56813_not ; n56814
g56559 and n56811_not n56814 ; n56815
g56560 and n56451_not n56815_not ; n56816
g56561 and b[28] n56440_not ; n56817
g56562 and n56438_not n56817 ; n56818
g56563 and n56442_not n56818_not ; n56819
g56564 and n56816_not n56819 ; n56820
g56565 and n56442_not n56820_not ; n56821
g56566 and b[29] n56431_not ; n56822
g56567 and n56429_not n56822 ; n56823
g56568 and n56433_not n56823_not ; n56824
g56569 and n56821_not n56824 ; n56825
g56570 and n56433_not n56825_not ; n56826
g56571 and b[30] n56422_not ; n56827
g56572 and n56420_not n56827 ; n56828
g56573 and n56424_not n56828_not ; n56829
g56574 and n56826_not n56829 ; n56830
g56575 and n56424_not n56830_not ; n56831
g56576 and b[31] n56413_not ; n56832
g56577 and n56411_not n56832 ; n56833
g56578 and n56415_not n56833_not ; n56834
g56579 and n56831_not n56834 ; n56835
g56580 and n56415_not n56835_not ; n56836
g56581 and b[32] n56404_not ; n56837
g56582 and n56402_not n56837 ; n56838
g56583 and n56406_not n56838_not ; n56839
g56584 and n56836_not n56839 ; n56840
g56585 and n56406_not n56840_not ; n56841
g56586 and b[33] n56395_not ; n56842
g56587 and n56393_not n56842 ; n56843
g56588 and n56397_not n56843_not ; n56844
g56589 and n56841_not n56844 ; n56845
g56590 and n56397_not n56845_not ; n56846
g56591 and b[34] n56386_not ; n56847
g56592 and n56384_not n56847 ; n56848
g56593 and n56388_not n56848_not ; n56849
g56594 and n56846_not n56849 ; n56850
g56595 and n56388_not n56850_not ; n56851
g56596 and b[35] n56377_not ; n56852
g56597 and n56375_not n56852 ; n56853
g56598 and n56379_not n56853_not ; n56854
g56599 and n56851_not n56854 ; n56855
g56600 and n56379_not n56855_not ; n56856
g56601 and b[36] n56368_not ; n56857
g56602 and n56366_not n56857 ; n56858
g56603 and n56370_not n56858_not ; n56859
g56604 and n56856_not n56859 ; n56860
g56605 and n56370_not n56860_not ; n56861
g56606 and b[37] n56359_not ; n56862
g56607 and n56357_not n56862 ; n56863
g56608 and n56361_not n56863_not ; n56864
g56609 and n56861_not n56864 ; n56865
g56610 and n56361_not n56865_not ; n56866
g56611 and b[38] n56350_not ; n56867
g56612 and n56348_not n56867 ; n56868
g56613 and n56352_not n56868_not ; n56869
g56614 and n56866_not n56869 ; n56870
g56615 and n56352_not n56870_not ; n56871
g56616 and b[39] n56341_not ; n56872
g56617 and n56339_not n56872 ; n56873
g56618 and n56343_not n56873_not ; n56874
g56619 and n56871_not n56874 ; n56875
g56620 and n56343_not n56875_not ; n56876
g56621 and b[40] n56332_not ; n56877
g56622 and n56330_not n56877 ; n56878
g56623 and n56334_not n56878_not ; n56879
g56624 and n56876_not n56879 ; n56880
g56625 and n56334_not n56880_not ; n56881
g56626 and b[41] n56323_not ; n56882
g56627 and n56321_not n56882 ; n56883
g56628 and n56325_not n56883_not ; n56884
g56629 and n56881_not n56884 ; n56885
g56630 and n56325_not n56885_not ; n56886
g56631 and b[42] n56314_not ; n56887
g56632 and n56312_not n56887 ; n56888
g56633 and n56316_not n56888_not ; n56889
g56634 and n56886_not n56889 ; n56890
g56635 and n56316_not n56890_not ; n56891
g56636 and b[43] n56305_not ; n56892
g56637 and n56303_not n56892 ; n56893
g56638 and n56307_not n56893_not ; n56894
g56639 and n56891_not n56894 ; n56895
g56640 and n56307_not n56895_not ; n56896
g56641 and b[44] n56296_not ; n56897
g56642 and n56294_not n56897 ; n56898
g56643 and n56298_not n56898_not ; n56899
g56644 and n56896_not n56899 ; n56900
g56645 and n56298_not n56900_not ; n56901
g56646 and b[45] n56287_not ; n56902
g56647 and n56285_not n56902 ; n56903
g56648 and n56289_not n56903_not ; n56904
g56649 and n56901_not n56904 ; n56905
g56650 and n56289_not n56905_not ; n56906
g56651 and b[46] n56278_not ; n56907
g56652 and n56276_not n56907 ; n56908
g56653 and n56280_not n56908_not ; n56909
g56654 and n56906_not n56909 ; n56910
g56655 and n56280_not n56910_not ; n56911
g56656 and b[47] n56269_not ; n56912
g56657 and n56267_not n56912 ; n56913
g56658 and n56271_not n56913_not ; n56914
g56659 and n56911_not n56914 ; n56915
g56660 and n56271_not n56915_not ; n56916
g56661 and b[48] n56260_not ; n56917
g56662 and n56258_not n56917 ; n56918
g56663 and n56262_not n56918_not ; n56919
g56664 and n56916_not n56919 ; n56920
g56665 and n56262_not n56920_not ; n56921
g56666 and b[49] n56251_not ; n56922
g56667 and n56249_not n56922 ; n56923
g56668 and n56253_not n56923_not ; n56924
g56669 and n56921_not n56924 ; n56925
g56670 and n56253_not n56925_not ; n56926
g56671 and b[50] n56242_not ; n56927
g56672 and n56240_not n56927 ; n56928
g56673 and n56244_not n56928_not ; n56929
g56674 and n56926_not n56929 ; n56930
g56675 and n56244_not n56930_not ; n56931
g56676 and b[51] n56233_not ; n56932
g56677 and n56231_not n56932 ; n56933
g56678 and n56235_not n56933_not ; n56934
g56679 and n56931_not n56934 ; n56935
g56680 and n56235_not n56935_not ; n56936
g56681 and b[52] n56224_not ; n56937
g56682 and n56222_not n56937 ; n56938
g56683 and n56226_not n56938_not ; n56939
g56684 and n56936_not n56939 ; n56940
g56685 and n56226_not n56940_not ; n56941
g56686 and b[53] n56215_not ; n56942
g56687 and n56213_not n56942 ; n56943
g56688 and n56217_not n56943_not ; n56944
g56689 and n56941_not n56944 ; n56945
g56690 and n56217_not n56945_not ; n56946
g56691 and b[54] n56206_not ; n56947
g56692 and n56204_not n56947 ; n56948
g56693 and n56208_not n56948_not ; n56949
g56694 and n56946_not n56949 ; n56950
g56695 and n56208_not n56950_not ; n56951
g56696 and b[55] n56197_not ; n56952
g56697 and n56195_not n56952 ; n56953
g56698 and n56199_not n56953_not ; n56954
g56699 and n56951_not n56954 ; n56955
g56700 and n56199_not n56955_not ; n56956
g56701 and b[56] n56188_not ; n56957
g56702 and n56186_not n56957 ; n56958
g56703 and n56190_not n56958_not ; n56959
g56704 and n56956_not n56959 ; n56960
g56705 and n56190_not n56960_not ; n56961
g56706 and b[57] n56179_not ; n56962
g56707 and n56177_not n56962 ; n56963
g56708 and n56181_not n56963_not ; n56964
g56709 and n56961_not n56964 ; n56965
g56710 and n56181_not n56965_not ; n56966
g56711 and b[58] n56170_not ; n56967
g56712 and n56168_not n56967 ; n56968
g56713 and n56172_not n56968_not ; n56969
g56714 and n56966_not n56969 ; n56970
g56715 and n56172_not n56970_not ; n56971
g56716 and b[59] n56161_not ; n56972
g56717 and n56159_not n56972 ; n56973
g56718 and n56163_not n56973_not ; n56974
g56719 and n56971_not n56974 ; n56975
g56720 and n56163_not n56975_not ; n56976
g56721 and b[60] n56152_not ; n56977
g56722 and n56150_not n56977 ; n56978
g56723 and n56154_not n56978_not ; n56979
g56724 and n56976_not n56979 ; n56980
g56725 and n56154_not n56980_not ; n56981
g56726 and b[61] n56143_not ; n56982
g56727 and n56141_not n56982 ; n56983
g56728 and n56145_not n56983_not ; n56984
g56729 and n56981_not n56984 ; n56985
g56730 and n56145_not n56985_not ; n56986
g56731 and b[62] n56134_not ; n56987
g56732 and n56132_not n56987 ; n56988
g56733 and n56136_not n56988_not ; n56989
g56734 and n56986_not n56989 ; n56990
g56735 and n56136_not n56990_not ; n56991
g56736 and b[63] n56125_not ; n56992
g56737 and n56123_not n56992 ; n56993
g56738 and n56127_not n56993_not ; n56994
g56739 and n56991_not n56994 ; n56995
g56740 and n56127_not n56995_not ; n56996
g56741 and b[0] n56996_not ; n56997
g56742 and a[0] n56997_not ; n56998
g56743 and n28345 n56996_not ; n56999
g56744 and n56998_not n56999_not ; remainder[0]
g56745 and n28345 n56682_not ; n57001
g56746 and n56680_not n57001 ; n57002
g56747 and n56684_not n57002_not ; n57003
g56748 and n56996_not n57003 ; n57004
g56749 and n56127_not n56679_not ; n57005
g56750 and n56995_not n57005 ; n57006
g56751 and n57004_not n57006_not ; remainder[1]
g56752 and n56685_not n56689 ; n57008
g56753 and n56684_not n57008 ; n57009
g56754 and n56686_not n56689_not ; n57010
g56755 and n57009_not n57010_not ; n57011
g56756 and n56996_not n57011_not ; n57012
g56757 and n56127_not n56674_not ; n57013
g56758 and n56995_not n57013 ; n57014
g56759 and n57012_not n57014_not ; remainder[2]
g56760 and n56675_not n56694 ; n57016
g56761 and n56690_not n57016 ; n57017
g56762 and n56691_not n56694_not ; n57018
g56763 and n57017_not n57018_not ; n57019
g56764 and n56996_not n57019_not ; n57020
g56765 and n56127_not n56666_not ; n57021
g56766 and n56995_not n57021 ; n57022
g56767 and n57020_not n57022_not ; remainder[3]
g56768 and n56667_not n56699 ; n57024
g56769 and n56695_not n57024 ; n57025
g56770 and n56696_not n56699_not ; n57026
g56771 and n57025_not n57026_not ; n57027
g56772 and n56996_not n57027_not ; n57028
g56773 and n56127_not n56657_not ; n57029
g56774 and n56995_not n57029 ; n57030
g56775 and n57028_not n57030_not ; remainder[4]
g56776 and n56658_not n56704 ; n57032
g56777 and n56700_not n57032 ; n57033
g56778 and n56701_not n56704_not ; n57034
g56779 and n57033_not n57034_not ; n57035
g56780 and n56996_not n57035_not ; n57036
g56781 and n56127_not n56648_not ; n57037
g56782 and n56995_not n57037 ; n57038
g56783 and n57036_not n57038_not ; remainder[5]
g56784 and n56649_not n56709 ; n57040
g56785 and n56705_not n57040 ; n57041
g56786 and n56706_not n56709_not ; n57042
g56787 and n57041_not n57042_not ; n57043
g56788 and n56996_not n57043_not ; n57044
g56789 and n56127_not n56639_not ; n57045
g56790 and n56995_not n57045 ; n57046
g56791 and n57044_not n57046_not ; remainder[6]
g56792 and n56640_not n56714 ; n57048
g56793 and n56710_not n57048 ; n57049
g56794 and n56711_not n56714_not ; n57050
g56795 and n57049_not n57050_not ; n57051
g56796 and n56996_not n57051_not ; n57052
g56797 and n56127_not n56630_not ; n57053
g56798 and n56995_not n57053 ; n57054
g56799 and n57052_not n57054_not ; remainder[7]
g56800 and n56631_not n56719 ; n57056
g56801 and n56715_not n57056 ; n57057
g56802 and n56716_not n56719_not ; n57058
g56803 and n57057_not n57058_not ; n57059
g56804 and n56996_not n57059_not ; n57060
g56805 and n56127_not n56621_not ; n57061
g56806 and n56995_not n57061 ; n57062
g56807 and n57060_not n57062_not ; remainder[8]
g56808 and n56622_not n56724 ; n57064
g56809 and n56720_not n57064 ; n57065
g56810 and n56721_not n56724_not ; n57066
g56811 and n57065_not n57066_not ; n57067
g56812 and n56996_not n57067_not ; n57068
g56813 and n56127_not n56612_not ; n57069
g56814 and n56995_not n57069 ; n57070
g56815 and n57068_not n57070_not ; remainder[9]
g56816 and n56613_not n56729 ; n57072
g56817 and n56725_not n57072 ; n57073
g56818 and n56726_not n56729_not ; n57074
g56819 and n57073_not n57074_not ; n57075
g56820 and n56996_not n57075_not ; n57076
g56821 and n56127_not n56603_not ; n57077
g56822 and n56995_not n57077 ; n57078
g56823 and n57076_not n57078_not ; remainder[10]
g56824 and n56604_not n56734 ; n57080
g56825 and n56730_not n57080 ; n57081
g56826 and n56731_not n56734_not ; n57082
g56827 and n57081_not n57082_not ; n57083
g56828 and n56996_not n57083_not ; n57084
g56829 and n56127_not n56594_not ; n57085
g56830 and n56995_not n57085 ; n57086
g56831 and n57084_not n57086_not ; remainder[11]
g56832 and n56595_not n56739 ; n57088
g56833 and n56735_not n57088 ; n57089
g56834 and n56736_not n56739_not ; n57090
g56835 and n57089_not n57090_not ; n57091
g56836 and n56996_not n57091_not ; n57092
g56837 and n56127_not n56585_not ; n57093
g56838 and n56995_not n57093 ; n57094
g56839 and n57092_not n57094_not ; remainder[12]
g56840 and n56586_not n56744 ; n57096
g56841 and n56740_not n57096 ; n57097
g56842 and n56741_not n56744_not ; n57098
g56843 and n57097_not n57098_not ; n57099
g56844 and n56996_not n57099_not ; n57100
g56845 and n56127_not n56576_not ; n57101
g56846 and n56995_not n57101 ; n57102
g56847 and n57100_not n57102_not ; remainder[13]
g56848 and n56577_not n56749 ; n57104
g56849 and n56745_not n57104 ; n57105
g56850 and n56746_not n56749_not ; n57106
g56851 and n57105_not n57106_not ; n57107
g56852 and n56996_not n57107_not ; n57108
g56853 and n56127_not n56567_not ; n57109
g56854 and n56995_not n57109 ; n57110
g56855 and n57108_not n57110_not ; remainder[14]
g56856 and n56568_not n56754 ; n57112
g56857 and n56750_not n57112 ; n57113
g56858 and n56751_not n56754_not ; n57114
g56859 and n57113_not n57114_not ; n57115
g56860 and n56996_not n57115_not ; n57116
g56861 and n56127_not n56558_not ; n57117
g56862 and n56995_not n57117 ; n57118
g56863 and n57116_not n57118_not ; remainder[15]
g56864 and n56559_not n56759 ; n57120
g56865 and n56755_not n57120 ; n57121
g56866 and n56756_not n56759_not ; n57122
g56867 and n57121_not n57122_not ; n57123
g56868 and n56996_not n57123_not ; n57124
g56869 and n56127_not n56549_not ; n57125
g56870 and n56995_not n57125 ; n57126
g56871 and n57124_not n57126_not ; remainder[16]
g56872 and n56550_not n56764 ; n57128
g56873 and n56760_not n57128 ; n57129
g56874 and n56761_not n56764_not ; n57130
g56875 and n57129_not n57130_not ; n57131
g56876 and n56996_not n57131_not ; n57132
g56877 and n56127_not n56540_not ; n57133
g56878 and n56995_not n57133 ; n57134
g56879 and n57132_not n57134_not ; remainder[17]
g56880 and n56541_not n56769 ; n57136
g56881 and n56765_not n57136 ; n57137
g56882 and n56766_not n56769_not ; n57138
g56883 and n57137_not n57138_not ; n57139
g56884 and n56996_not n57139_not ; n57140
g56885 and n56127_not n56531_not ; n57141
g56886 and n56995_not n57141 ; n57142
g56887 and n57140_not n57142_not ; remainder[18]
g56888 and n56532_not n56774 ; n57144
g56889 and n56770_not n57144 ; n57145
g56890 and n56771_not n56774_not ; n57146
g56891 and n57145_not n57146_not ; n57147
g56892 and n56996_not n57147_not ; n57148
g56893 and n56127_not n56522_not ; n57149
g56894 and n56995_not n57149 ; n57150
g56895 and n57148_not n57150_not ; remainder[19]
g56896 and n56523_not n56779 ; n57152
g56897 and n56775_not n57152 ; n57153
g56898 and n56776_not n56779_not ; n57154
g56899 and n57153_not n57154_not ; n57155
g56900 and n56996_not n57155_not ; n57156
g56901 and n56127_not n56513_not ; n57157
g56902 and n56995_not n57157 ; n57158
g56903 and n57156_not n57158_not ; remainder[20]
g56904 and n56514_not n56784 ; n57160
g56905 and n56780_not n57160 ; n57161
g56906 and n56781_not n56784_not ; n57162
g56907 and n57161_not n57162_not ; n57163
g56908 and n56996_not n57163_not ; n57164
g56909 and n56127_not n56504_not ; n57165
g56910 and n56995_not n57165 ; n57166
g56911 and n57164_not n57166_not ; remainder[21]
g56912 and n56505_not n56789 ; n57168
g56913 and n56785_not n57168 ; n57169
g56914 and n56786_not n56789_not ; n57170
g56915 and n57169_not n57170_not ; n57171
g56916 and n56996_not n57171_not ; n57172
g56917 and n56127_not n56495_not ; n57173
g56918 and n56995_not n57173 ; n57174
g56919 and n57172_not n57174_not ; remainder[22]
g56920 and n56496_not n56794 ; n57176
g56921 and n56790_not n57176 ; n57177
g56922 and n56791_not n56794_not ; n57178
g56923 and n57177_not n57178_not ; n57179
g56924 and n56996_not n57179_not ; n57180
g56925 and n56127_not n56486_not ; n57181
g56926 and n56995_not n57181 ; n57182
g56927 and n57180_not n57182_not ; remainder[23]
g56928 and n56487_not n56799 ; n57184
g56929 and n56795_not n57184 ; n57185
g56930 and n56796_not n56799_not ; n57186
g56931 and n57185_not n57186_not ; n57187
g56932 and n56996_not n57187_not ; n57188
g56933 and n56127_not n56477_not ; n57189
g56934 and n56995_not n57189 ; n57190
g56935 and n57188_not n57190_not ; remainder[24]
g56936 and n56478_not n56804 ; n57192
g56937 and n56800_not n57192 ; n57193
g56938 and n56801_not n56804_not ; n57194
g56939 and n57193_not n57194_not ; n57195
g56940 and n56996_not n57195_not ; n57196
g56941 and n56127_not n56468_not ; n57197
g56942 and n56995_not n57197 ; n57198
g56943 and n57196_not n57198_not ; remainder[25]
g56944 and n56469_not n56809 ; n57200
g56945 and n56805_not n57200 ; n57201
g56946 and n56806_not n56809_not ; n57202
g56947 and n57201_not n57202_not ; n57203
g56948 and n56996_not n57203_not ; n57204
g56949 and n56127_not n56459_not ; n57205
g56950 and n56995_not n57205 ; n57206
g56951 and n57204_not n57206_not ; remainder[26]
g56952 and n56460_not n56814 ; n57208
g56953 and n56810_not n57208 ; n57209
g56954 and n56811_not n56814_not ; n57210
g56955 and n57209_not n57210_not ; n57211
g56956 and n56996_not n57211_not ; n57212
g56957 and n56127_not n56450_not ; n57213
g56958 and n56995_not n57213 ; n57214
g56959 and n57212_not n57214_not ; remainder[27]
g56960 and n56451_not n56819 ; n57216
g56961 and n56815_not n57216 ; n57217
g56962 and n56816_not n56819_not ; n57218
g56963 and n57217_not n57218_not ; n57219
g56964 and n56996_not n57219_not ; n57220
g56965 and n56127_not n56441_not ; n57221
g56966 and n56995_not n57221 ; n57222
g56967 and n57220_not n57222_not ; remainder[28]
g56968 and n56442_not n56824 ; n57224
g56969 and n56820_not n57224 ; n57225
g56970 and n56821_not n56824_not ; n57226
g56971 and n57225_not n57226_not ; n57227
g56972 and n56996_not n57227_not ; n57228
g56973 and n56127_not n56432_not ; n57229
g56974 and n56995_not n57229 ; n57230
g56975 and n57228_not n57230_not ; remainder[29]
g56976 and n56433_not n56829 ; n57232
g56977 and n56825_not n57232 ; n57233
g56978 and n56826_not n56829_not ; n57234
g56979 and n57233_not n57234_not ; n57235
g56980 and n56996_not n57235_not ; n57236
g56981 and n56127_not n56423_not ; n57237
g56982 and n56995_not n57237 ; n57238
g56983 and n57236_not n57238_not ; remainder[30]
g56984 and n56424_not n56834 ; n57240
g56985 and n56830_not n57240 ; n57241
g56986 and n56831_not n56834_not ; n57242
g56987 and n57241_not n57242_not ; n57243
g56988 and n56996_not n57243_not ; n57244
g56989 and n56127_not n56414_not ; n57245
g56990 and n56995_not n57245 ; n57246
g56991 and n57244_not n57246_not ; remainder[31]
g56992 and n56415_not n56839 ; n57248
g56993 and n56835_not n57248 ; n57249
g56994 and n56836_not n56839_not ; n57250
g56995 and n57249_not n57250_not ; n57251
g56996 and n56996_not n57251_not ; n57252
g56997 and n56127_not n56405_not ; n57253
g56998 and n56995_not n57253 ; n57254
g56999 and n57252_not n57254_not ; remainder[32]
g57000 and n56406_not n56844 ; n57256
g57001 and n56840_not n57256 ; n57257
g57002 and n56841_not n56844_not ; n57258
g57003 and n57257_not n57258_not ; n57259
g57004 and n56996_not n57259_not ; n57260
g57005 and n56127_not n56396_not ; n57261
g57006 and n56995_not n57261 ; n57262
g57007 and n57260_not n57262_not ; remainder[33]
g57008 and n56397_not n56849 ; n57264
g57009 and n56845_not n57264 ; n57265
g57010 and n56846_not n56849_not ; n57266
g57011 and n57265_not n57266_not ; n57267
g57012 and n56996_not n57267_not ; n57268
g57013 and n56127_not n56387_not ; n57269
g57014 and n56995_not n57269 ; n57270
g57015 and n57268_not n57270_not ; remainder[34]
g57016 and n56388_not n56854 ; n57272
g57017 and n56850_not n57272 ; n57273
g57018 and n56851_not n56854_not ; n57274
g57019 and n57273_not n57274_not ; n57275
g57020 and n56996_not n57275_not ; n57276
g57021 and n56127_not n56378_not ; n57277
g57022 and n56995_not n57277 ; n57278
g57023 and n57276_not n57278_not ; remainder[35]
g57024 and n56379_not n56859 ; n57280
g57025 and n56855_not n57280 ; n57281
g57026 and n56856_not n56859_not ; n57282
g57027 and n57281_not n57282_not ; n57283
g57028 and n56996_not n57283_not ; n57284
g57029 and n56127_not n56369_not ; n57285
g57030 and n56995_not n57285 ; n57286
g57031 and n57284_not n57286_not ; remainder[36]
g57032 and n56370_not n56864 ; n57288
g57033 and n56860_not n57288 ; n57289
g57034 and n56861_not n56864_not ; n57290
g57035 and n57289_not n57290_not ; n57291
g57036 and n56996_not n57291_not ; n57292
g57037 and n56127_not n56360_not ; n57293
g57038 and n56995_not n57293 ; n57294
g57039 and n57292_not n57294_not ; remainder[37]
g57040 and n56361_not n56869 ; n57296
g57041 and n56865_not n57296 ; n57297
g57042 and n56866_not n56869_not ; n57298
g57043 and n57297_not n57298_not ; n57299
g57044 and n56996_not n57299_not ; n57300
g57045 and n56127_not n56351_not ; n57301
g57046 and n56995_not n57301 ; n57302
g57047 and n57300_not n57302_not ; remainder[38]
g57048 and n56352_not n56874 ; n57304
g57049 and n56870_not n57304 ; n57305
g57050 and n56871_not n56874_not ; n57306
g57051 and n57305_not n57306_not ; n57307
g57052 and n56996_not n57307_not ; n57308
g57053 and n56127_not n56342_not ; n57309
g57054 and n56995_not n57309 ; n57310
g57055 and n57308_not n57310_not ; remainder[39]
g57056 and n56343_not n56879 ; n57312
g57057 and n56875_not n57312 ; n57313
g57058 and n56876_not n56879_not ; n57314
g57059 and n57313_not n57314_not ; n57315
g57060 and n56996_not n57315_not ; n57316
g57061 and n56127_not n56333_not ; n57317
g57062 and n56995_not n57317 ; n57318
g57063 and n57316_not n57318_not ; remainder[40]
g57064 and n56334_not n56884 ; n57320
g57065 and n56880_not n57320 ; n57321
g57066 and n56881_not n56884_not ; n57322
g57067 and n57321_not n57322_not ; n57323
g57068 and n56996_not n57323_not ; n57324
g57069 and n56127_not n56324_not ; n57325
g57070 and n56995_not n57325 ; n57326
g57071 and n57324_not n57326_not ; remainder[41]
g57072 and n56325_not n56889 ; n57328
g57073 and n56885_not n57328 ; n57329
g57074 and n56886_not n56889_not ; n57330
g57075 and n57329_not n57330_not ; n57331
g57076 and n56996_not n57331_not ; n57332
g57077 and n56127_not n56315_not ; n57333
g57078 and n56995_not n57333 ; n57334
g57079 and n57332_not n57334_not ; remainder[42]
g57080 and n56316_not n56894 ; n57336
g57081 and n56890_not n57336 ; n57337
g57082 and n56891_not n56894_not ; n57338
g57083 and n57337_not n57338_not ; n57339
g57084 and n56996_not n57339_not ; n57340
g57085 and n56127_not n56306_not ; n57341
g57086 and n56995_not n57341 ; n57342
g57087 and n57340_not n57342_not ; remainder[43]
g57088 and n56307_not n56899 ; n57344
g57089 and n56895_not n57344 ; n57345
g57090 and n56896_not n56899_not ; n57346
g57091 and n57345_not n57346_not ; n57347
g57092 and n56996_not n57347_not ; n57348
g57093 and n56127_not n56297_not ; n57349
g57094 and n56995_not n57349 ; n57350
g57095 and n57348_not n57350_not ; remainder[44]
g57096 and n56298_not n56904 ; n57352
g57097 and n56900_not n57352 ; n57353
g57098 and n56901_not n56904_not ; n57354
g57099 and n57353_not n57354_not ; n57355
g57100 and n56996_not n57355_not ; n57356
g57101 and n56127_not n56288_not ; n57357
g57102 and n56995_not n57357 ; n57358
g57103 and n57356_not n57358_not ; remainder[45]
g57104 and n56289_not n56909 ; n57360
g57105 and n56905_not n57360 ; n57361
g57106 and n56906_not n56909_not ; n57362
g57107 and n57361_not n57362_not ; n57363
g57108 and n56996_not n57363_not ; n57364
g57109 and n56127_not n56279_not ; n57365
g57110 and n56995_not n57365 ; n57366
g57111 and n57364_not n57366_not ; remainder[46]
g57112 and n56280_not n56914 ; n57368
g57113 and n56910_not n57368 ; n57369
g57114 and n56911_not n56914_not ; n57370
g57115 and n57369_not n57370_not ; n57371
g57116 and n56996_not n57371_not ; n57372
g57117 and n56127_not n56270_not ; n57373
g57118 and n56995_not n57373 ; n57374
g57119 and n57372_not n57374_not ; remainder[47]
g57120 and n56271_not n56919 ; n57376
g57121 and n56915_not n57376 ; n57377
g57122 and n56916_not n56919_not ; n57378
g57123 and n57377_not n57378_not ; n57379
g57124 and n56996_not n57379_not ; n57380
g57125 and n56127_not n56261_not ; n57381
g57126 and n56995_not n57381 ; n57382
g57127 and n57380_not n57382_not ; remainder[48]
g57128 and n56262_not n56924 ; n57384
g57129 and n56920_not n57384 ; n57385
g57130 and n56921_not n56924_not ; n57386
g57131 and n57385_not n57386_not ; n57387
g57132 and n56996_not n57387_not ; n57388
g57133 and n56127_not n56252_not ; n57389
g57134 and n56995_not n57389 ; n57390
g57135 and n57388_not n57390_not ; remainder[49]
g57136 and n56253_not n56929 ; n57392
g57137 and n56925_not n57392 ; n57393
g57138 and n56926_not n56929_not ; n57394
g57139 and n57393_not n57394_not ; n57395
g57140 and n56996_not n57395_not ; n57396
g57141 and n56127_not n56243_not ; n57397
g57142 and n56995_not n57397 ; n57398
g57143 and n57396_not n57398_not ; remainder[50]
g57144 and n56244_not n56934 ; n57400
g57145 and n56930_not n57400 ; n57401
g57146 and n56931_not n56934_not ; n57402
g57147 and n57401_not n57402_not ; n57403
g57148 and n56996_not n57403_not ; n57404
g57149 and n56127_not n56234_not ; n57405
g57150 and n56995_not n57405 ; n57406
g57151 and n57404_not n57406_not ; remainder[51]
g57152 and n56235_not n56939 ; n57408
g57153 and n56935_not n57408 ; n57409
g57154 and n56936_not n56939_not ; n57410
g57155 and n57409_not n57410_not ; n57411
g57156 and n56996_not n57411_not ; n57412
g57157 and n56127_not n56225_not ; n57413
g57158 and n56995_not n57413 ; n57414
g57159 and n57412_not n57414_not ; remainder[52]
g57160 and n56226_not n56944 ; n57416
g57161 and n56940_not n57416 ; n57417
g57162 and n56941_not n56944_not ; n57418
g57163 and n57417_not n57418_not ; n57419
g57164 and n56996_not n57419_not ; n57420
g57165 and n56127_not n56216_not ; n57421
g57166 and n56995_not n57421 ; n57422
g57167 and n57420_not n57422_not ; remainder[53]
g57168 and n56217_not n56949 ; n57424
g57169 and n56945_not n57424 ; n57425
g57170 and n56946_not n56949_not ; n57426
g57171 and n57425_not n57426_not ; n57427
g57172 and n56996_not n57427_not ; n57428
g57173 and n56127_not n56207_not ; n57429
g57174 and n56995_not n57429 ; n57430
g57175 and n57428_not n57430_not ; remainder[54]
g57176 and n56208_not n56954 ; n57432
g57177 and n56950_not n57432 ; n57433
g57178 and n56951_not n56954_not ; n57434
g57179 and n57433_not n57434_not ; n57435
g57180 and n56996_not n57435_not ; n57436
g57181 and n56127_not n56198_not ; n57437
g57182 and n56995_not n57437 ; n57438
g57183 and n57436_not n57438_not ; remainder[55]
g57184 and n56199_not n56959 ; n57440
g57185 and n56955_not n57440 ; n57441
g57186 and n56956_not n56959_not ; n57442
g57187 and n57441_not n57442_not ; n57443
g57188 and n56996_not n57443_not ; n57444
g57189 and n56127_not n56189_not ; n57445
g57190 and n56995_not n57445 ; n57446
g57191 and n57444_not n57446_not ; remainder[56]
g57192 and n56190_not n56964 ; n57448
g57193 and n56960_not n57448 ; n57449
g57194 and n56961_not n56964_not ; n57450
g57195 and n57449_not n57450_not ; n57451
g57196 and n56996_not n57451_not ; n57452
g57197 and n56127_not n56180_not ; n57453
g57198 and n56995_not n57453 ; n57454
g57199 and n57452_not n57454_not ; remainder[57]
g57200 and n56181_not n56969 ; n57456
g57201 and n56965_not n57456 ; n57457
g57202 and n56966_not n56969_not ; n57458
g57203 and n57457_not n57458_not ; n57459
g57204 and n56996_not n57459_not ; n57460
g57205 and n56127_not n56171_not ; n57461
g57206 and n56995_not n57461 ; n57462
g57207 and n57460_not n57462_not ; remainder[58]
g57208 and n56172_not n56974 ; n57464
g57209 and n56970_not n57464 ; n57465
g57210 and n56971_not n56974_not ; n57466
g57211 and n57465_not n57466_not ; n57467
g57212 and n56996_not n57467_not ; n57468
g57213 and n56127_not n56162_not ; n57469
g57214 and n56995_not n57469 ; n57470
g57215 and n57468_not n57470_not ; remainder[59]
g57216 and n56163_not n56979 ; n57472
g57217 and n56975_not n57472 ; n57473
g57218 and n56976_not n56979_not ; n57474
g57219 and n57473_not n57474_not ; n57475
g57220 and n56996_not n57475_not ; n57476
g57221 and n56127_not n56153_not ; n57477
g57222 and n56995_not n57477 ; n57478
g57223 and n57476_not n57478_not ; remainder[60]
g57224 and n56154_not n56984 ; n57480
g57225 and n56980_not n57480 ; n57481
g57226 and n56981_not n56984_not ; n57482
g57227 and n57481_not n57482_not ; n57483
g57228 and n56996_not n57483_not ; n57484
g57229 and n56127_not n56144_not ; n57485
g57230 and n56995_not n57485 ; n57486
g57231 and n57484_not n57486_not ; remainder[61]
g57232 and n56145_not n56989 ; n57488
g57233 and n56985_not n57488 ; n57489
g57234 and n56986_not n56989_not ; n57490
g57235 and n57489_not n57490_not ; n57491
g57236 and n56996_not n57491_not ; n57492
g57237 and n56127_not n56135_not ; n57493
g57238 and n56995_not n57493 ; n57494
g57239 and n57492_not n57494_not ; remainder[62]
g57240 and n56136_not n56994 ; n57496
g57241 and n56990_not n57496 ; n57497
g57242 and n56991_not n56994_not ; n57498
g57243 and n57497_not n57498_not ; n57499
g57244 and n56996_not n57499_not ; n57500
g57245 and n56126_not n56127_not ; n57501
g57246 and n56995_not n57501 ; n57502
g57247 and n57500_not n57502_not ; remainder[63]
g57248 not n500 ; n500_not
g57249 not n501 ; n501_not
g57250 not n510 ; n510_not
g57251 not n321 ; n321_not
g57252 not n330 ; n330_not
g57253 not n502 ; n502_not
g57254 not n322 ; n322_not
g57255 not n331 ; n331_not
g57256 not n521 ; n521_not
g57257 not n440 ; n440_not
g57258 not n800 ; n800_not
g57259 not n620 ; n620_not
g57260 not n611 ; n611_not
g57261 not n323 ; n323_not
g57262 not n503 ; n503_not
g57263 not n530 ; n530_not
g57264 not n504 ; n504_not
g57265 not n522 ; n522_not
g57266 not n360 ; n360_not
g57267 not n441 ; n441_not
g57268 not n621 ; n621_not
g57269 not n612 ; n612_not
g57270 not n720 ; n720_not
g57271 not n711 ; n711_not
g57272 not n531 ; n531_not
g57273 not n900 ; n900_not
g57274 not n810 ; n810_not
g57275 not n801 ; n801_not
g57276 not n603 ; n603_not
g57277 not n361 ; n361_not
g57278 not n910 ; n910_not
g57279 not n901 ; n901_not
g57280 not n532 ; n532_not
g57281 not n703 ; n703_not
g57282 not n811 ; n811_not
g57283 not n325 ; n325_not
g57284 not n640 ; n640_not
g57285 not n523 ; n523_not
g57286 not n730 ; n730_not
g57287 not n820 ; n820_not
g57288 not n622 ; n622_not
g57289 not n613 ; n613_not
g57290 not n514 ; n514_not
g57291 not n712 ; n712_not
g57292 not n721 ; n721_not
g57293 not n442 ; n442_not
g57294 not n802 ; n802_not
g57295 not n604 ; n604_not
g57296 not n505 ; n505_not
g57297 not n623 ; n623_not
g57298 not n614 ; n614_not
g57299 not n434 ; n434_not
g57300 not n326 ; n326_not
g57301 not n506 ; n506_not
g57302 not n803 ; n803_not
g57303 not n722 ; n722_not
g57304 not n362 ; n362_not
g57305 not n470 ; n470_not
g57306 not n443 ; n443_not
g57307 not n452 ; n452_not
g57308 not n704 ; n704_not
g57309 not n713 ; n713_not
g57310 not n471 ; n471_not
g57311 not n480 ; n480_not
g57312 not n363 ; n363_not
g57313 not n453 ; n453_not
g57314 not n813 ; n813_not
g57315 not n921 ; n921_not
g57316 not n435 ; n435_not
g57317 not n327 ; n327_not
g57318 not n426 ; n426_not
g57319 not n507 ; n507_not
g57320 not n444 ; n444_not
g57321 not n903 ; n903_not
g57322 not n840 ; n840_not
g57323 not n804 ; n804_not
g57324 not n912 ; n912_not
g57325 not n534 ; n534_not
g57326 not n606 ; n606_not
g57327 not n930 ; n930_not
g57328 not n750 ; n750_not
g57329 not n822 ; n822_not
g57330 not n741 ; n741_not
g57331 not n732 ; n732_not
g57332 not n831 ; n831_not
g57333 not n841 ; n841_not
g57334 not n508 ; n508_not
g57335 not n490 ; n490_not
g57336 not n733 ; n733_not
g57337 not n751 ; n751_not
g57338 not n481 ; n481_not
g57339 not n832 ; n832_not
g57340 not n814 ; n814_not
g57341 not n904 ; n904_not
g57342 not n823 ; n823_not
g57343 not n931 ; n931_not
g57344 not n553 ; n553_not
g57345 not n913 ; n913_not
g57346 not n544 ; n544_not
g57347 not n526 ; n526_not
g57348 not n571 ; n571_not
g57349 not n517 ; n517_not
g57350 not n580 ; n580_not
g57351 not n607 ; n607_not
g57352 not n922 ; n922_not
g57353 not n625 ; n625_not
g57354 not n670 ; n670_not
g57355 not n715 ; n715_not
g57356 not n724 ; n724_not
g57357 not n427 ; n427_not
g57358 not n436 ; n436_not
g57359 not n940 ; n940_not
g57360 not n445 ; n445_not
g57361 not n805 ; n805_not
g57362 not n472 ; n472_not
g57363 not n328 ; n328_not
g57364 not n743 ; n743_not
g57365 not n626 ; n626_not
g57366 not n572 ; n572_not
g57367 not n923 ; n923_not
g57368 not n941 ; n941_not
g57369 not n752 ; n752_not
g57370 not n554 ; n554_not
g57371 not n671 ; n671_not
g57372 not n545 ; n545_not
g57373 not n437 ; n437_not
g57374 not n761 ; n761_not
g57375 not n581 ; n581_not
g57376 not n932 ; n932_not
g57377 not n617 ; n617_not
g57378 not n824 ; n824_not
g57379 not n680 ; n680_not
g57380 not n608 ; n608_not
g57381 not n860 ; n860_not
g57382 not n815 ; n815_not
g57383 not n257 ; n257_not
g57384 not n707 ; n707_not
g57385 not n734 ; n734_not
g57386 not n329 ; n329_not
g57387 not n914 ; n914_not
g57388 not n662 ; n662_not
g57389 not n833 ; n833_not
g57390 not n806 ; n806_not
g57391 not n905 ; n905_not
g57392 not n446 ; n446_not
g57393 not n509 ; n509_not
g57394 not n527 ; n527_not
g57395 not n456 ; n456_not
g57396 not n816 ; n816_not
g57397 not n861 ; n861_not
g57398 not n609 ; n609_not
g57399 not n825 ; n825_not
g57400 not n906 ; n906_not
g57401 not n717 ; n717_not
g57402 not n807 ; n807_not
g57403 not n582 ; n582_not
g57404 not n636 ; n636_not
g57405 not n555 ; n555_not
g57406 not n942 ; n942_not
g57407 not n681 ; n681_not
g57408 not n483 ; n483_not
g57409 not n618 ; n618_not
g57410 not n834 ; n834_not
g57411 not n933 ; n933_not
g57412 not n870 ; n870_not
g57413 not n924 ; n924_not
g57414 not n771 ; n771_not
g57415 not n546 ; n546_not
g57416 not n663 ; n663_not
g57417 not n726 ; n726_not
g57418 not n735 ; n735_not
g57419 not n915 ; n915_not
g57420 not n762 ; n762_not
g57421 not n519 ; n519_not
g57422 not n438 ; n438_not
g57423 not n573 ; n573_not
g57424 not n637 ; n637_not
g57425 not n673 ; n673_not
g57426 not n349 ; n349_not
g57427 not n664 ; n664_not
g57428 not n583 ; n583_not
g57429 not n763 ; n763_not
g57430 not n772 ; n772_not
g57431 not n790 ; n790_not
g57432 not n781 ; n781_not
g57433 not n709 ; n709_not
g57434 not n745 ; n745_not
g57435 not n754 ; n754_not
g57436 not n970 ; n970_not
g57437 not n574 ; n574_not
g57438 not n961 ; n961_not
g57439 not n682 ; n682_not
g57440 not n691 ; n691_not
g57441 not n547 ; n547_not
g57442 not n880 ; n880_not
g57443 not n529 ; n529_not
g57444 not n871 ; n871_not
g57445 not n862 ; n862_not
g57446 not n565 ; n565_not
g57447 not n692 ; n692_not
g57448 not n980 ; n980_not
g57449 not n548 ; n548_not
g57450 not n890 ; n890_not
g57451 not n674 ; n674_not
g57452 not n728 ; n728_not
g57453 not n764 ; n764_not
g57454 not n737 ; n737_not
g57455 not n863 ; n863_not
g57456 not n584 ; n584_not
g57457 not n962 ; n962_not
g57458 not n557 ; n557_not
g57459 not n854 ; n854_not
g57460 not n827 ; n827_not
g57461 not n755 ; n755_not
g57462 not n575 ; n575_not
g57463 not n935 ; n935_not
g57464 not n836 ; n836_not
g57465 not n719 ; n719_not
g57466 not n926 ; n926_not
g57467 not n566 ; n566_not
g57468 not n746 ; n746_not
g57469 not n656 ; n656_not
g57470 not n908 ; n908_not
g57471 not n647 ; n647_not
g57472 not n809 ; n809_not
g57473 not n872 ; n872_not
g57474 not n818 ; n818_not
g57475 not n458 ; n458_not
g57476 not n782 ; n782_not
g57477 not n917 ; n917_not
g57478 not n638 ; n638_not
g57479 not n683 ; n683_not
g57480 not n359 ; n359_not
g57481 not n944 ; n944_not
g57482 not n881 ; n881_not
g57483 not n773 ; n773_not
g57484 not n756 ; n756_not
g57485 not n738 ; n738_not
g57486 not n873 ; n873_not
g57487 not n774 ; n774_not
g57488 not n972 ; n972_not
g57489 not n648 ; n648_not
g57490 not n747 ; n747_not
g57491 not n990 ; n990_not
g57492 not n666 ; n666_not
g57493 not n576 ; n576_not
g57494 not n963 ; n963_not
g57495 not n819 ; n819_not
g57496 not n729 ; n729_not
g57497 not n558 ; n558_not
g57498 not n927 ; n927_not
g57499 not n783 ; n783_not
g57500 not n855 ; n855_not
g57501 not n468 ; n468_not
g57502 not n828 ; n828_not
g57503 not n792 ; n792_not
g57504 not n918 ; n918_not
g57505 not n936 ; n936_not
g57506 not n882 ; n882_not
g57507 not n693 ; n693_not
g57508 not n675 ; n675_not
g57509 not n657 ; n657_not
g57510 not n909 ; n909_not
g57511 not n891 ; n891_not
g57512 not n639 ; n639_not
g57513 not n847 ; n847_not
g57514 not n694 ; n694_not
g57515 not n496 ; n496_not
g57516 not n919 ; n919_not
g57517 not n739 ; n739_not
g57518 not n883 ; n883_not
g57519 not n766 ; n766_not
g57520 not n757 ; n757_not
g57521 not n856 ; n856_not
g57522 not n982 ; n982_not
g57523 not n469 ; n469_not
g57524 not n685 ; n685_not
g57525 not n784 ; n784_not
g57526 not n649 ; n649_not
g57527 not n973 ; n973_not
g57528 not n955 ; n955_not
g57529 not n559 ; n559_not
g57530 not n577 ; n577_not
g57531 not n928 ; n928_not
g57532 not n586 ; n586_not
g57533 not n829 ; n829_not
g57534 not n748 ; n748_not
g57535 not n793 ; n793_not
g57536 not n937 ; n937_not
g57537 not n676 ; n676_not
g57538 not n667 ; n667_not
g57539 not n865 ; n865_not
g57540 not n892 ; n892_not
g57541 not n974 ; n974_not
g57542 not n839 ; n839_not
g57543 not n479 ; n479_not
g57544 not n992 ; n992_not
g57545 not n893 ; n893_not
g57546 not n497 ; n497_not
g57547 not n668 ; n668_not
g57548 not n848 ; n848_not
g57549 not n767 ; n767_not
g57550 not n875 ; n875_not
g57551 not n758 ; n758_not
g57552 not n677 ; n677_not
g57553 not n956 ; n956_not
g57554 not n866 ; n866_not
g57555 not n749 ; n749_not
g57556 not n965 ; n965_not
g57557 not n578 ; n578_not
g57558 not n947 ; n947_not
g57559 not n794 ; n794_not
g57560 not n776 ; n776_not
g57561 not n983 ; n983_not
g57562 not n759 ; n759_not
g57563 not n858 ; n858_not
g57564 not n867 ; n867_not
g57565 not n498 ; n498_not
g57566 not n939 ; n939_not
g57567 not n669 ; n669_not
g57568 not n993 ; n993_not
g57569 not n579 ; n579_not
g57570 not n966 ; n966_not
g57571 not n489 ; n489_not
g57572 not n678 ; n678_not
g57573 not n696 ; n696_not
g57574 not n984 ; n984_not
g57575 not n948 ; n948_not
g57576 not n975 ; n975_not
g57577 not n768 ; n768_not
g57578 not n777 ; n777_not
g57579 not n885 ; n885_not
g57580 not n876 ; n876_not
g57581 not n499 ; n499_not
g57582 not n985 ; n985_not
g57583 not n967 ; n967_not
g57584 not n994 ; n994_not
g57585 not n949 ; n949_not
g57586 not n877 ; n877_not
g57587 not n868 ; n868_not
g57588 not n859 ; n859_not
g57589 not n769 ; n769_not
g57590 not n778 ; n778_not
g57591 not n796 ; n796_not
g57592 not n886 ; n886_not
g57593 not n697 ; n697_not
g57594 not n688 ; n688_not
g57595 not n679 ; n679_not
g57596 not n797 ; n797_not
g57597 not n878 ; n878_not
g57598 not n887 ; n887_not
g57599 not n995 ; n995_not
g57600 not n977 ; n977_not
g57601 not n968 ; n968_not
g57602 not n689 ; n689_not
g57603 not n779 ; n779_not
g57604 not n897 ; n897_not
g57605 not n987 ; n987_not
g57606 not n969 ; n969_not
g57607 not n888 ; n888_not
g57608 not n798 ; n798_not
g57609 not n978 ; n978_not
g57610 not n979 ; n979_not
g57611 not n997 ; n997_not
g57612 not n988 ; n988_not
g57613 not n989 ; n989_not
g57614 not n899 ; n899_not
g57615 not n998 ; n998_not
g57616 not n999 ; n999_not
g57617 not n1000 ; n1000_not
g57618 not n1010 ; n1010_not
g57619 not n1001 ; n1001_not
g57620 not n2000 ; n2000_not
g57621 not n1100 ; n1100_not
g57622 not n1020 ; n1020_not
g57623 not n1101 ; n1101_not
g57624 not n1110 ; n1110_not
g57625 not n3000 ; n3000_not
g57626 not n1200 ; n1200_not
g57627 not n2010 ; n2010_not
g57628 not n2100 ; n2100_not
g57629 not n2200 ; n2200_not
g57630 not n1111 ; n1111_not
g57631 not n3100 ; n3100_not
g57632 not n1120 ; n1120_not
g57633 not n2011 ; n2011_not
g57634 not n3001 ; n3001_not
g57635 not n1021 ; n1021_not
g57636 not n1102 ; n1102_not
g57637 not n3010 ; n3010_not
g57638 not n2002 ; n2002_not
g57639 not n1030 ; n1030_not
g57640 not n2110 ; n2110_not
g57641 not n2101 ; n2101_not
g57642 not n1300 ; n1300_not
g57643 not n1003 ; n1003_not
g57644 not n2300 ; n2300_not
g57645 not n3101 ; n3101_not
g57646 not n2021 ; n2021_not
g57647 not n2111 ; n2111_not
g57648 not n1121 ; n1121_not
g57649 not n1130 ; n1130_not
g57650 not n2012 ; n2012_not
g57651 not n2102 ; n2102_not
g57652 not n2201 ; n2201_not
g57653 not n5000 ; n5000_not
g57654 not n1004 ; n1004_not
g57655 not n4001 ; n4001_not
g57656 not n3020 ; n3020_not
g57657 not n2030 ; n2030_not
g57658 not n2120 ; n2120_not
g57659 not n3011 ; n3011_not
g57660 not n1220 ; n1220_not
g57661 not n1211 ; n1211_not
g57662 not n1202 ; n1202_not
g57663 not n3110 ; n3110_not
g57664 not n2210 ; n2210_not
g57665 not n1112 ; n1112_not
g57666 not n3200 ; n3200_not
g57667 not n3002 ; n3002_not
g57668 not n1040 ; n1040_not
g57669 not n4010 ; n4010_not
g57670 not n1400 ; n1400_not
g57671 not n1022 ; n1022_not
g57672 not n1031 ; n1031_not
g57673 not n2003 ; n2003_not
g57674 not n2211 ; n2211_not
g57675 not n2004 ; n2004_not
g57676 not n2013 ; n2013_not
g57677 not n2220 ; n2220_not
g57678 not n1050 ; n1050_not
g57679 not n2022 ; n2022_not
g57680 not n3300 ; n3300_not
g57681 not n1320 ; n1320_not
g57682 not n2031 ; n2031_not
g57683 not n2040 ; n2040_not
g57684 not n1041 ; n1041_not
g57685 not n1311 ; n1311_not
g57686 not n5010 ; n5010_not
g57687 not n1302 ; n1302_not
g57688 not n1032 ; n1032_not
g57689 not n2202 ; n2202_not
g57690 not n2400 ; n2400_not
g57691 not n5001 ; n5001_not
g57692 not n1140 ; n1140_not
g57693 not n1131 ; n1131_not
g57694 not n1410 ; n1410_not
g57695 not n1122 ; n1122_not
g57696 not n1104 ; n1104_not
g57697 not n1203 ; n1203_not
g57698 not n1212 ; n1212_not
g57699 not n3201 ; n3201_not
g57700 not n1500 ; n1500_not
g57701 not n4011 ; n4011_not
g57702 not n4002 ; n4002_not
g57703 not n4101 ; n4101_not
g57704 not n3210 ; n3210_not
g57705 not n1005 ; n1005_not
g57706 not n4300 ; n4300_not
g57707 not n5011 ; n5011_not
g57708 not n1141 ; n1141_not
g57709 not n1132 ; n1132_not
g57710 not n2320 ; n2320_not
g57711 not n1150 ; n1150_not
g57712 not n5020 ; n5020_not
g57713 not n1402 ; n1402_not
g57714 not n3211 ; n3211_not
g57715 not n2050 ; n2050_not
g57716 not n2410 ; n2410_not
g57717 not n2311 ; n2311_not
g57718 not n3301 ; n3301_not
g57719 not n1015 ; n1015_not
g57720 not n3103 ; n3103_not
g57721 not n3040 ; n3040_not
g57722 not n3202 ; n3202_not
g57723 not n4003 ; n4003_not
g57724 not n3310 ; n3310_not
g57725 not n3400 ; n3400_not
g57726 not n2500 ; n2500_not
g57727 not n4210 ; n4210_not
g57728 not n5200 ; n5200_not
g57729 not n5002 ; n5002_not
g57730 not n1114 ; n1114_not
g57731 not n1420 ; n1420_not
g57732 not n1060 ; n1060_not
g57733 not n1051 ; n1051_not
g57734 not n1042 ; n1042_not
g57735 not n1024 ; n1024_not
g57736 not n2140 ; n2140_not
g57737 not n2230 ; n2230_not
g57738 not n1330 ; n1330_not
g57739 not n2041 ; n2041_not
g57740 not n2131 ; n2131_not
g57741 not n2221 ; n2221_not
g57742 not n1321 ; n1321_not
g57743 not n6001 ; n6001_not
g57744 not n2122 ; n2122_not
g57745 not n1312 ; n1312_not
g57746 not n2113 ; n2113_not
g57747 not n2212 ; n2212_not
g57748 not n2104 ; n2104_not
g57749 not n1303 ; n1303_not
g57750 not n6100 ; n6100_not
g57751 not n3022 ; n3022_not
g57752 not n2302 ; n2302_not
g57753 not n7000 ; n7000_not
g57754 not n3004 ; n3004_not
g57755 not n3112 ; n3112_not
g57756 not n4030 ; n4030_not
g57757 not n6010 ; n6010_not
g57758 not n1204 ; n1204_not
g57759 not n3121 ; n3121_not
g57760 not n1105 ; n1105_not
g57761 not n1213 ; n1213_not
g57762 not n1231 ; n1231_not
g57763 not n3013 ; n3013_not
g57764 not n3031 ; n3031_not
g57765 not n4102 ; n4102_not
g57766 not n3220 ; n3220_not
g57767 not n2005 ; n2005_not
g57768 not n4201 ; n4201_not
g57769 not n4111 ; n4111_not
g57770 not n1006 ; n1006_not
g57771 not n5101 ; n5101_not
g57772 not n7001 ; n7001_not
g57773 not n1142 ; n1142_not
g57774 not n2420 ; n2420_not
g57775 not n3113 ; n3113_not
g57776 not n1034 ; n1034_not
g57777 not n2123 ; n2123_not
g57778 not n4031 ; n4031_not
g57779 not n1106 ; n1106_not
g57780 not n1502 ; n1502_not
g57781 not n5300 ; n5300_not
g57782 not n2402 ; n2402_not
g57783 not n4310 ; n4310_not
g57784 not n2132 ; n2132_not
g57785 not n5021 ; n5021_not
g57786 not n1025 ; n1025_not
g57787 not n2303 ; n2303_not
g57788 not n3041 ; n3041_not
g57789 not n4202 ; n4202_not
g57790 not n3320 ; n3320_not
g57791 not n2015 ; n2015_not
g57792 not n5102 ; n5102_not
g57793 not n2105 ; n2105_not
g57794 not n6020 ; n6020_not
g57795 not n1016 ; n1016_not
g57796 not n2114 ; n2114_not
g57797 not n3311 ; n3311_not
g57798 not n6200 ; n6200_not
g57799 not n3005 ; n3005_not
g57800 not n1241 ; n1241_not
g57801 not n6011 ; n6011_not
g57802 not n3302 ; n3302_not
g57803 not n1511 ; n1511_not
g57804 not n1115 ; n1115_not
g57805 not n6110 ; n6110_not
g57806 not n2222 ; n2222_not
g57807 not n6002 ; n6002_not
g57808 not n2231 ; n2231_not
g57809 not n2042 ; n2042_not
g57810 not n4004 ; n4004_not
g57811 not n3500 ; n3500_not
g57812 not n2006 ; n2006_not
g57813 not n1331 ; n1331_not
g57814 not n1322 ; n1322_not
g57815 not n3140 ; n3140_not
g57816 not n7010 ; n7010_not
g57817 not n6101 ; n6101_not
g57818 not n5003 ; n5003_not
g57819 not n1007 ; n1007_not
g57820 not n3023 ; n3023_not
g57821 not n1160 ; n1160_not
g57822 not n1430 ; n1430_not
g57823 not n2204 ; n2204_not
g57824 not n4220 ; n4220_not
g57825 not n3230 ; n3230_not
g57826 not n1250 ; n1250_not
g57827 not n2141 ; n2141_not
g57828 not n8000 ; n8000_not
g57829 not n1223 ; n1223_not
g57830 not n5012 ; n5012_not
g57831 not n5111 ; n5111_not
g57832 not n1232 ; n1232_not
g57833 not n2060 ; n2060_not
g57834 not n3032 ; n3032_not
g57835 not n2150 ; n2150_not
g57836 not n2051 ; n2051_not
g57837 not n3014 ; n3014_not
g57838 not n1340 ; n1340_not
g57839 not n2240 ; n2240_not
g57840 not n3212 ; n3212_not
g57841 not n3203 ; n3203_not
g57842 not n1520 ; n1520_not
g57843 not n4121 ; n4121_not
g57844 not n1403 ; n1403_not
g57845 not n4211 ; n4211_not
g57846 not n1124 ; n1124_not
g57847 not n1601 ; n1601_not
g57848 not n4112 ; n4112_not
g57849 not n2330 ; n2330_not
g57850 not n2312 ; n2312_not
g57851 not n1412 ; n1412_not
g57852 not n1304 ; n1304_not
g57853 not n3221 ; n3221_not
g57854 not n1313 ; n1313_not
g57855 not n4301 ; n4301_not
g57856 not n5201 ; n5201_not
g57857 not n5210 ; n5210_not
g57858 not n4103 ; n4103_not
g57859 not n3050 ; n3050_not
g57860 not n2501 ; n2501_not
g57861 not n2510 ; n2510_not
g57862 not n2321 ; n2321_not
g57863 not n1151 ; n1151_not
g57864 not n3104 ; n3104_not
g57865 not n5112 ; n5112_not
g57866 not n7101 ; n7101_not
g57867 not n1305 ; n1305_not
g57868 not n1701 ; n1701_not
g57869 not n1350 ; n1350_not
g57870 not n6021 ; n6021_not
g57871 not n1521 ; n1521_not
g57872 not n1161 ; n1161_not
g57873 not n2124 ; n2124_not
g57874 not n5040 ; n5040_not
g57875 not n3510 ; n3510_not
g57876 not n6300 ; n6300_not
g57877 not n3303 ; n3303_not
g57878 not n3501 ; n3501_not
g57879 not n1611 ; n1611_not
g57880 not n2133 ; n2133_not
g57881 not n1503 ; n1503_not
g57882 not n1314 ; n1314_not
g57883 not n1224 ; n1224_not
g57884 not n1530 ; n1530_not
g57885 not n6030 ; n6030_not
g57886 not n4032 ; n4032_not
g57887 not n5103 ; n5103_not
g57888 not n4113 ; n4113_not
g57889 not n5400 ; n5400_not
g57890 not n3240 ; n3240_not
g57891 not n1440 ; n1440_not
g57892 not n3312 ; n3312_not
g57893 not n1341 ; n1341_not
g57894 not n2106 ; n2106_not
g57895 not n1413 ; n1413_not
g57896 not n4104 ; n4104_not
g57897 not n3420 ; n3420_not
g57898 not n9000 ; n9000_not
g57899 not n6210 ; n6210_not
g57900 not n3222 ; n3222_not
g57901 not n3321 ; n3321_not
g57902 not n7002 ; n7002_not
g57903 not n2115 ; n2115_not
g57904 not n2160 ; n2160_not
g57905 not n1332 ; n1332_not
g57906 not n3330 ; n3330_not
g57907 not n5121 ; n5121_not
g57908 not n1422 ; n1422_not
g57909 not n4401 ; n4401_not
g57910 not n3141 ; n3141_not
g57911 not n1323 ; n1323_not
g57912 not n4122 ; n4122_not
g57913 not n2151 ; n2151_not
g57914 not n1251 ; n1251_not
g57915 not n4041 ; n4041_not
g57916 not n1512 ; n1512_not
g57917 not n2034 ; n2034_not
g57918 not n1404 ; n1404_not
g57919 not n4131 ; n4131_not
g57920 not n6201 ; n6201_not
g57921 not n1602 ; n1602_not
g57922 not n1800 ; n1800_not
g57923 not n6003 ; n6003_not
g57924 not n3213 ; n3213_not
g57925 not n2142 ; n2142_not
g57926 not n4500 ; n4500_not
g57927 not n8010 ; n8010_not
g57928 not n3015 ; n3015_not
g57929 not n1710 ; n1710_not
g57930 not n3006 ; n3006_not
g57931 not n2025 ; n2025_not
g57932 not n1260 ; n1260_not
g57933 not n6012 ; n6012_not
g57934 not n2340 ; n2340_not
g57935 not n2331 ; n2331_not
g57936 not n1206 ; n1206_not
g57937 not n1107 ; n1107_not
g57938 not n4212 ; n4212_not
g57939 not n2430 ; n2430_not
g57940 not n4203 ; n4203_not
g57941 not n2322 ; n2322_not
g57942 not n2232 ; n2232_not
g57943 not n1080 ; n1080_not
g57944 not n6111 ; n6111_not
g57945 not n2502 ; n2502_not
g57946 not n2205 ; n2205_not
g57947 not n3600 ; n3600_not
g57948 not n3033 ; n3033_not
g57949 not n2070 ; n2070_not
g57950 not n2304 ; n2304_not
g57951 not n2403 ; n2403_not
g57952 not n1134 ; n1134_not
g57953 not n1215 ; n1215_not
g57954 not n1071 ; n1071_not
g57955 not n4302 ; n4302_not
g57956 not n3105 ; n3105_not
g57957 not n1125 ; n1125_not
g57958 not n1170 ; n1170_not
g57959 not n3042 ; n3042_not
g57960 not n2241 ; n2241_not
g57961 not n4221 ; n4221_not
g57962 not n2250 ; n2250_not
g57963 not n2511 ; n2511_not
g57964 not n3051 ; n3051_not
g57965 not n4230 ; n4230_not
g57966 not n2520 ; n2520_not
g57967 not n1116 ; n1116_not
g57968 not n6120 ; n6120_not
g57969 not n3231 ; n3231_not
g57970 not n2313 ; n2313_not
g57971 not n1035 ; n1035_not
g57972 not n3132 ; n3132_not
g57973 not n2052 ; n2052_not
g57974 not n1062 ; n1062_not
g57975 not n2043 ; n2043_not
g57976 not n1008 ; n1008_not
g57977 not n6102 ; n6102_not
g57978 not n7011 ; n7011_not
g57979 not n2412 ; n2412_not
g57980 not n8100 ; n8100_not
g57981 not n3060 ; n3060_not
g57982 not n3024 ; n3024_not
g57983 not n2061 ; n2061_not
g57984 not n2214 ; n2214_not
g57985 not n4311 ; n4311_not
g57986 not n1053 ; n1053_not
g57987 not n1242 ; n1242_not
g57988 not n3150 ; n3150_not
g57989 not n3114 ; n3114_not
g57990 not n1044 ; n1044_not
g57991 not n4320 ; n4320_not
g57992 not n9001 ; n9001_not
g57993 not n5212 ; n5212_not
g57994 not n3412 ; n3412_not
g57995 not n5203 ; n5203_not
g57996 not n7300 ; n7300_not
g57997 not n5131 ; n5131_not
g57998 not n4132 ; n4132_not
g57999 not n2422 ; n2422_not
g58000 not n3223 ; n3223_not
g58001 not n5113 ; n5113_not
g58002 not n1414 ; n1414_not
g58003 not n4123 ; n4123_not
g58004 not n2305 ; n2305_not
g58005 not n1423 ; n1423_not
g58006 not n5104 ; n5104_not
g58007 not n2800 ; n2800_not
g58008 not n2008 ; n2008_not
g58009 not n2314 ; n2314_not
g58010 not n3160 ; n3160_not
g58011 not n4411 ; n4411_not
g58012 not n4114 ; n4114_not
g58013 not n7111 ; n7111_not
g58014 not n2242 ; n2242_not
g58015 not n8110 ; n8110_not
g58016 not n3151 ; n3151_not
g58017 not n1405 ; n1405_not
g58018 not n2701 ; n2701_not
g58019 not n2251 ; n2251_not
g58020 not n3430 ; n3430_not
g58021 not n2440 ; n2440_not
g58022 not n4042 ; n4042_not
g58023 not n2260 ; n2260_not
g58024 not n1720 ; n1720_not
g58025 not n1603 ; n1603_not
g58026 not n1504 ; n1504_not
g58027 not n8101 ; n8101_not
g58028 not n5311 ; n5311_not
g58029 not n4051 ; n4051_not
g58030 not n1612 ; n1612_not
g58031 not n5302 ; n5302_not
g58032 not n5041 ; n5041_not
g58033 not n7021 ; n7021_not
g58034 not n8200 ; n8200_not
g58035 not n3232 ; n3232_not
g58036 not n4510 ; n4510_not
g58037 not n1630 ; n1630_not
g58038 not n5401 ; n5401_not
g58039 not n4501 ; n4501_not
g58040 not n2404 ; n2404_not
g58041 not n1540 ; n1540_not
g58042 not n3133 ; n3133_not
g58043 not n1531 ; n1531_not
g58044 not n2620 ; n2620_not
g58045 not n4600 ; n4600_not
g58046 not n1702 ; n1702_not
g58047 not n7201 ; n7201_not
g58048 not n7012 ; n7012_not
g58049 not n7003 ; n7003_not
g58050 not n2611 ; n2611_not
g58051 not n1522 ; n1522_not
g58052 not n3124 ; n3124_not
g58053 not n2602 ; n2602_not
g58054 not n1711 ; n1711_not
g58055 not n4033 ; n4033_not
g58056 not n1513 ; n1513_not
g58057 not n5320 ; n5320_not
g58058 not n7210 ; n7210_not
g58059 not n5122 ; n5122_not
g58060 not n3421 ; n3421_not
g58061 not n6211 ; n6211_not
g58062 not n5230 ; n5230_not
g58063 not n3511 ; n3511_not
g58064 not n4006 ; n4006_not
g58065 not n5221 ; n5221_not
g58066 not n6202 ; n6202_not
g58067 not n6310 ; n6310_not
g58068 not n1621 ; n1621_not
g58069 not n2413 ; n2413_not
g58070 not n9010 ; n9010_not
g58071 not n1810 ; n1810_not
g58072 not n6301 ; n6301_not
g58073 not n8020 ; n8020_not
g58074 not n1801 ; n1801_not
g58075 not n3205 ; n3205_not
g58076 not n1243 ; n1243_not
g58077 not n1045 ; n1045_not
g58078 not n1126 ; n1126_not
g58079 not n1171 ; n1171_not
g58080 not n1054 ; n1054_not
g58081 not n1180 ; n1180_not
g58082 not n1063 ; n1063_not
g58083 not n1117 ; n1117_not
g58084 not n1072 ; n1072_not
g58085 not n4402 ; n4402_not
g58086 not n1081 ; n1081_not
g58087 not n1090 ; n1090_not
g58088 not n2206 ; n2206_not
g58089 not n2350 ; n2350_not
g58090 not n6400 ; n6400_not
g58091 not n2161 ; n2161_not
g58092 not n1432 ; n1432_not
g58093 not n2341 ; n2341_not
g58094 not n2170 ; n2170_not
g58095 not n2332 ; n2332_not
g58096 not n2323 ; n2323_not
g58097 not n1036 ; n1036_not
g58098 not n1135 ; n1135_not
g58099 not n1153 ; n1153_not
g58100 not n1225 ; n1225_not
g58101 not n5014 ; n5014_not
g58102 not n4330 ; n4330_not
g58103 not n1261 ; n1261_not
g58104 not n2224 ; n2224_not
g58105 not n1270 ; n1270_not
g58106 not n1162 ; n1162_not
g58107 not n5005 ; n5005_not
g58108 not n1207 ; n1207_not
g58109 not n5023 ; n5023_not
g58110 not n2215 ; n2215_not
g58111 not n1216 ; n1216_not
g58112 not n2152 ; n2152_not
g58113 not n9100 ; n9100_not
g58114 not n1450 ; n1450_not
g58115 not n2026 ; n2026_not
g58116 not n2035 ; n2035_not
g58117 not n1441 ; n1441_not
g58118 not n6220 ; n6220_not
g58119 not n8002 ; n8002_not
g58120 not n7102 ; n7102_not
g58121 not n8210 ; n8210_not
g58122 not n2162 ; n2162_not
g58123 not n8102 ; n8102_not
g58124 not n5303 ; n5303_not
g58125 not n8030 ; n8030_not
g58126 not n3251 ; n3251_not
g58127 not n2522 ; n2522_not
g58128 not n6104 ; n6104_not
g58129 not n8201 ; n8201_not
g58130 not n2216 ; n2216_not
g58131 not n4061 ; n4061_not
g58132 not n3161 ; n3161_not
g58133 not n2405 ; n2405_not
g58134 not n2036 ; n2036_not
g58135 not n5123 ; n5123_not
g58136 not n8120 ; n8120_not
g58137 not n6023 ; n6023_not
g58138 not n2144 ; n2144_not
g58139 not n6311 ; n6311_not
g58140 not n2504 ; n2504_not
g58141 not n8111 ; n8111_not
g58142 not n4151 ; n4151_not
g58143 not n2153 ; n2153_not
g58144 not n6014 ; n6014_not
g58145 not n5114 ; n5114_not
g58146 not n2513 ; n2513_not
g58147 not n6221 ; n6221_not
g58148 not n8300 ; n8300_not
g58149 not n4133 ; n4133_not
g58150 not n4412 ; n4412_not
g58151 not n2603 ; n2603_not
g58152 not n2612 ; n2612_not
g58153 not n4232 ; n4232_not
g58154 not n1703 ; n1703_not
g58155 not n3332 ; n3332_not
g58156 not n1811 ; n1811_not
g58157 not n2207 ; n2207_not
g58158 not n2009 ; n2009_not
g58159 not n5006 ; n5006_not
g58160 not n4700 ; n4700_not
g58161 not n2621 ; n2621_not
g58162 not n2540 ; n2540_not
g58163 not n5330 ; n5330_not
g58164 not n2900 ; n2900_not
g58165 not n7004 ; n7004_not
g58166 not n2630 ; n2630_not
g58167 not n5312 ; n5312_not
g58168 not n3035 ; n3035_not
g58169 not n2801 ; n2801_not
g58170 not n2027 ; n2027_not
g58171 not n5015 ; n5015_not
g58172 not n1721 ; n1721_not
g58173 not n4214 ; n4214_not
g58174 not n2234 ; n2234_not
g58175 not n2171 ; n2171_not
g58176 not n6005 ; n6005_not
g58177 not n2225 ; n2225_not
g58178 not n7013 ; n7013_not
g58179 not n2414 ; n2414_not
g58180 not n4124 ; n4124_not
g58181 not n6302 ; n6302_not
g58182 not n4241 ; n4241_not
g58183 not n4043 ; n4043_not
g58184 not n5321 ; n5321_not
g58185 not n1712 ; n1712_not
g58186 not n2531 ; n2531_not
g58187 not n4106 ; n4106_not
g58188 not n3413 ; n3413_not
g58189 not n2072 ; n2072_not
g58190 not n5222 ; n5222_not
g58191 not n2450 ; n2450_not
g58192 not n4403 ; n4403_not
g58193 not n6131 ; n6131_not
g58194 not n5132 ; n5132_not
g58195 not n3350 ; n3350_not
g58196 not n5231 ; n5231_not
g58197 not n6041 ; n6041_not
g58198 not n2180 ; n2180_not
g58199 not n6122 ; n6122_not
g58200 not n7031 ; n7031_not
g58201 not n3143 ; n3143_not
g58202 not n6320 ; n6320_not
g58203 not n5240 ; n5240_not
g58204 not n3017 ; n3017_not
g58205 not n2081 ; n2081_not
g58206 not n3431 ; n3431_not
g58207 not n6050 ; n6050_not
g58208 not n2063 ; n2063_not
g58209 not n1910 ; n1910_not
g58210 not n4160 ; n4160_not
g58211 not n3008 ; n3008_not
g58212 not n3206 ; n3206_not
g58213 not n3215 ; n3215_not
g58214 not n5204 ; n5204_not
g58215 not n1901 ; n1901_not
g58216 not n6140 ; n6140_not
g58217 not n5213 ; n5213_not
g58218 not n8012 ; n8012_not
g58219 not n7121 ; n7121_not
g58220 not n3314 ; n3314_not
g58221 not n4205 ; n4205_not
g58222 not n2054 ; n2054_not
g58223 not n4331 ; n4331_not
g58224 not n3323 ; n3323_not
g58225 not n1820 ; n1820_not
g58226 not n1802 ; n1802_not
g58227 not n2810 ; n2810_not
g58228 not n3233 ; n3233_not
g58229 not n3026 ; n3026_not
g58230 not n2126 ; n2126_not
g58231 not n3152 ; n3152_not
g58232 not n6032 ; n6032_not
g58233 not n5141 ; n5141_not
g58234 not n6113 ; n6113_not
g58235 not n3260 ; n3260_not
g58236 not n2432 ; n2432_not
g58237 not n2135 ; n2135_not
g58238 not n2090 ; n2090_not
g58239 not n3242 ; n3242_not
g58240 not n5051 ; n5051_not
g58241 not n3440 ; n3440_not
g58242 not n3125 ; n3125_not
g58243 not n4223 ; n4223_not
g58244 not n3341 ; n3341_not
g58245 not n2045 ; n2045_not
g58246 not n3305 ; n3305_not
g58247 not n6212 ; n6212_not
g58248 not n2108 ; n2108_not
g58249 not n5042 ; n5042_not
g58250 not n7103 ; n7103_not
g58251 not n2423 ; n2423_not
g58252 not n2117 ; n2117_not
g58253 not n1208 ; n1208_not
g58254 not n1154 ; n1154_not
g58255 not n1343 ; n1343_not
g58256 not n5402 ; n5402_not
g58257 not n3107 ; n3107_not
g58258 not n1163 ; n1163_not
g58259 not n7310 ; n7310_not
g58260 not n4313 ; n4313_not
g58261 not n3170 ; n3170_not
g58262 not n1325 ; n1325_not
g58263 not n1613 ; n1613_not
g58264 not n4025 ; n4025_not
g58265 not n3512 ; n3512_not
g58266 not n4421 ; n4421_not
g58267 not n3710 ; n3710_not
g58268 not n1091 ; n1091_not
g58269 not n1082 ; n1082_not
g58270 not n1640 ; n1640_not
g58271 not n1217 ; n1217_not
g58272 not n1622 ; n1622_not
g58273 not n1172 ; n1172_not
g58274 not n1415 ; n1415_not
g58275 not n3071 ; n3071_not
g58276 not n6401 ; n6401_not
g58277 not n1424 ; n1424_not
g58278 not n4322 ; n4322_not
g58279 not n1631 ; n1631_not
g58280 not n4304 ; n4304_not
g58281 not n4250 ; n4250_not
g58282 not n3521 ; n3521_not
g58283 not n3701 ; n3701_not
g58284 not n5501 ; n5501_not
g58285 not n3053 ; n3053_not
g58286 not n1280 ; n1280_not
g58287 not n4034 ; n4034_not
g58288 not n1181 ; n1181_not
g58289 not n1019 ; n1019_not
g58290 not n3530 ; n3530_not
g58291 not n6500 ; n6500_not
g58292 not n1064 ; n1064_not
g58293 not n1433 ; n1433_not
g58294 not n7211 ; n7211_not
g58295 not n1028 ; n1028_not
g58296 not n1271 ; n1271_not
g58297 not n1334 ; n1334_not
g58298 not n3062 ; n3062_not
g58299 not n4052 ; n4052_not
g58300 not n5411 ; n5411_not
g58301 not n1055 ; n1055_not
g58302 not n1604 ; n1604_not
g58303 not n1190 ; n1190_not
g58304 not n1127 ; n1127_not
g58305 not n1460 ; n1460_not
g58306 not n3116 ; n3116_not
g58307 not n6410 ; n6410_not
g58308 not n3620 ; n3620_not
g58309 not n1370 ; n1370_not
g58310 not n1244 ; n1244_not
g58311 not n8003 ; n8003_not
g58312 not n1136 ; n1136_not
g58313 not n7022 ; n7022_not
g58314 not n7220 ; n7220_not
g58315 not n1037 ; n1037_not
g58316 not n1046 ; n1046_not
g58317 not n3602 ; n3602_not
g58318 not n1316 ; n1316_not
g58319 not n3080 ; n3080_not
g58320 not n1073 ; n1073_not
g58321 not n1307 ; n1307_not
g58322 not n3044 ; n3044_not
g58323 not n6230 ; n6230_not
g58324 not n1361 ; n1361_not
g58325 not n7202 ; n7202_not
g58326 not n1352 ; n1352_not
g58327 not n3503 ; n3503_not
g58328 not n7301 ; n7301_not
g58329 not n3611 ; n3611_not
g58330 not n1109 ; n1109_not
g58331 not n7400 ; n7400_not
g58332 not n7112 ; n7112_not
g58333 not n1253 ; n1253_not
g58334 not n3333 ; n3333_not
g58335 not n3153 ; n3153_not
g58336 not n2613 ; n2613_not
g58337 not n5601 ; n5601_not
g58338 not n6222 ; n6222_not
g58339 not n7032 ; n7032_not
g58340 not n3162 ; n3162_not
g58341 not n3072 ; n3072_not
g58342 not n2181 ; n2181_not
g58343 not n7023 ; n7023_not
g58344 not n4224 ; n4224_not
g58345 not n6042 ; n6042_not
g58346 not n3252 ; n3252_not
g58347 not n3126 ; n3126_not
g58348 not n4233 ; n4233_not
g58349 not n3018 ; n3018_not
g58350 not n2820 ; n2820_not
g58351 not n5106 ; n5106_not
g58352 not n2730 ; n2730_not
g58353 not n2631 ; n2631_not
g58354 not n3063 ; n3063_not
g58355 not n3117 ; n3117_not
g58356 not n2442 ; n2442_not
g58357 not n2172 ; n2172_not
g58358 not n1515 ; n1515_not
g58359 not n6150 ; n6150_not
g58360 not n8040 ; n8040_not
g58361 not n1029 ; n1029_not
g58362 not n5133 ; n5133_not
g58363 not n3036 ; n3036_not
g58364 not n5124 ; n5124_not
g58365 not n7104 ; n7104_not
g58366 not n2550 ; n2550_not
g58367 not n4314 ; n4314_not
g58368 not n6105 ; n6105_not
g58369 not n5151 ; n5151_not
g58370 not n6330 ; n6330_not
g58371 not n1506 ; n1506_not
g58372 not n1317 ; n1317_not
g58373 not n5700 ; n5700_not
g58374 not n2802 ; n2802_not
g58375 not n3108 ; n3108_not
g58376 not n3225 ; n3225_not
g58377 not n2415 ; n2415_not
g58378 not n4404 ; n4404_not
g58379 not n2901 ; n2901_not
g58380 not n4413 ; n4413_not
g58381 not n4134 ; n4134_not
g58382 not n2712 ; n2712_not
g58383 not n6312 ; n6312_not
g58384 not n2424 ; n2424_not
g58385 not n4422 ; n4422_not
g58386 not n3360 ; n3360_not
g58387 not n4251 ; n4251_not
g58388 not n2640 ; n2640_not
g58389 not n1326 ; n1326_not
g58390 not n4215 ; n4215_not
g58391 not n1524 ; n1524_not
g58392 not n9300 ; n9300_not
g58393 not n5610 ; n5610_not
g58394 not n4152 ; n4152_not
g58395 not n4260 ; n4260_not
g58396 not n6060 ; n6060_not
g58397 not n9111 ; n9111_not
g58398 not n3081 ; n3081_not
g58399 not n1119 ; n1119_not
g58400 not n3315 ; n3315_not
g58401 not n2091 ; n2091_not
g58402 not n6402 ; n6402_not
g58403 not n2343 ; n2343_not
g58404 not n3612 ; n3612_not
g58405 not n7230 ; n7230_not
g58406 not n4242 ; n4242_not
g58407 not n2532 ; n2532_not
g58408 not n4026 ; n4026_not
g58409 not n6132 ; n6132_not
g58410 not n2811 ; n2811_not
g58411 not n2082 ; n2082_not
g58412 not n4332 ; n4332_not
g58413 not n2910 ; n2910_not
g58414 not n1407 ; n1407_not
g58415 not n5061 ; n5061_not
g58416 not n4323 ; n4323_not
g58417 not n2307 ; n2307_not
g58418 not n2352 ; n2352_not
g58419 not n6510 ; n6510_not
g58420 not n2190 ; n2190_not
g58421 not n6123 ; n6123_not
g58422 not n2073 ; n2073_not
g58423 not n6141 ; n6141_not
g58424 not n2316 ; n2316_not
g58425 not n1137 ; n1137_not
g58426 not n1245 ; n1245_not
g58427 not n2523 ; n2523_not
g58428 not n2136 ; n2136_not
g58429 not n2127 ; n2127_not
g58430 not n5034 ; n5034_not
g58431 not n1362 ; n1362_not
g58432 not n1353 ; n1353_not
g58433 not n3009 ; n3009_not
g58434 not n2118 ; n2118_not
g58435 not n3045 ; n3045_not
g58436 not n1254 ; n1254_not
g58437 not n6600 ; n6600_not
g58438 not n2325 ; n2325_not
g58439 not n3603 ; n3603_not
g58440 not n1155 ; n1155_not
g58441 not n1380 ; n1380_not
g58442 not n3243 ; n3243_not
g58443 not n2109 ; n2109_not
g58444 not n4170 ; n4170_not
g58445 not n2334 ; n2334_not
g58446 not n3342 ; n3342_not
g58447 not n8004 ; n8004_not
g58448 not n4305 ; n4305_not
g58449 not n7113 ; n7113_not
g58450 not n3306 ; n3306_not
g58451 not n2541 ; n2541_not
g58452 not n1461 ; n1461_not
g58453 not n6015 ; n6015_not
g58454 not n2037 ; n2037_not
g58455 not n2721 ; n2721_not
g58456 not n9030 ; n9030_not
g58457 not n4107 ; n4107_not
g58458 not n5016 ; n5016_not
g58459 not n3441 ; n3441_not
g58460 not n1470 ; n1470_not
g58461 not n2154 ; n2154_not
g58462 not n2028 ; n2028_not
g58463 not n6501 ; n6501_not
g58464 not n1164 ; n1164_not
g58465 not n3054 ; n3054_not
g58466 not n1335 ; n1335_not
g58467 not n6006 ; n6006_not
g58468 not n6051 ; n6051_not
g58469 not n1425 ; n1425_not
g58470 not n1173 ; n1173_not
g58471 not n6114 ; n6114_not
g58472 not n7041 ; n7041_not
g58473 not n3090 ; n3090_not
g58474 not n6321 ; n6321_not
g58475 not n1434 ; n1434_not
g58476 not n1092 ; n1092_not
g58477 not n1344 ; n1344_not
g58478 not n2064 ; n2064_not
g58479 not n4161 ; n4161_not
g58480 not n9120 ; n9120_not
g58481 not n5511 ; n5511_not
g58482 not n1443 ; n1443_not
g58483 not n2361 ; n2361_not
g58484 not n2055 ; n2055_not
g58485 not n3171 ; n3171_not
g58486 not n7122 ; n7122_not
g58487 not n3351 ; n3351_not
g58488 not n9102 ; n9102_not
g58489 not n2046 ; n2046_not
g58490 not n3180 ; n3180_not
g58491 not n9021 ; n9021_not
g58492 not n4512 ; n4512_not
g58493 not n2460 ; n2460_not
g58494 not n3207 ; n3207_not
g58495 not n1623 ; n1623_not
g58496 not n4521 ; n4521_not
g58497 not n3711 ; n3711_not
g58498 not n9012 ; n9012_not
g58499 not n6024 ; n6024_not
g58500 not n1614 ; n1614_not
g58501 not n1632 ; n1632_not
g58502 not n4530 ; n4530_not
g58503 not n1731 ; n1731_not
g58504 not n5304 ; n5304_not
g58505 not n5052 ; n5052_not
g58506 not n4053 ; n4053_not
g58507 not n1641 ; n1641_not
g58508 not n4710 ; n4710_not
g58509 not n4062 ; n4062_not
g58510 not n4611 ; n4611_not
g58511 not n8022 ; n8022_not
g58512 not n4503 ; n4503_not
g58513 not n2271 ; n2271_not
g58514 not n1821 ; n1821_not
g58515 not n1803 ; n1803_not
g58516 not n3450 ; n3450_not
g58517 not n3261 ; n3261_not
g58518 not n2226 ; n2226_not
g58519 not n1812 ; n1812_not
g58520 not n1191 ; n1191_not
g58521 not n7401 ; n7401_not
g58522 not n1263 ; n1263_not
g58523 not n4071 ; n4071_not
g58524 not n6240 ; n6240_not
g58525 not n3027 ; n3027_not
g58526 not n1182 ; n1182_not
g58527 not n6033 ; n6033_not
g58528 not n8400 ; n8400_not
g58529 not n9210 ; n9210_not
g58530 not n4602 ; n4602_not
g58531 not n5502 ; n5502_not
g58532 not n5322 ; n5322_not
g58533 not n7203 ; n7203_not
g58534 not n2217 ; n2217_not
g58535 not n4620 ; n4620_not
g58536 not n3900 ; n3900_not
g58537 not n7410 ; n7410_not
g58538 not n7005 ; n7005_not
g58539 not n5340 ; n5340_not
g58540 not n3630 ; n3630_not
g58541 not n9201 ; n9201_not
g58542 not n5331 ; n5331_not
g58543 not n3144 ; n3144_not
g58544 not n1218 ; n1218_not
g58545 not n2253 ; n2253_not
g58546 not n5313 ; n5313_not
g58547 not n3270 ; n3270_not
g58548 not n2505 ; n2505_not
g58549 not n1209 ; n1209_not
g58550 not n1740 ; n1740_not
g58551 not n2244 ; n2244_not
g58552 not n6231 ; n6231_not
g58553 not n7014 ; n7014_not
g58554 not n2262 ; n2262_not
g58555 not n6420 ; n6420_not
g58556 not n4044 ; n4044_not
g58557 not n3216 ; n3216_not
g58558 not n1281 ; n1281_not
g58559 not n7302 ; n7302_not
g58560 not n3531 ; n3531_not
g58561 not n1551 ; n1551_not
g58562 not n4701 ; n4701_not
g58563 not n6204 ; n6204_not
g58564 not n5142 ; n5142_not
g58565 not n3540 ; n3540_not
g58566 not n5214 ; n5214_not
g58567 not n3414 ; n3414_not
g58568 not n2280 ; n2280_not
g58569 not n1290 ; n1290_not
g58570 not n7311 ; n7311_not
g58571 not n1560 ; n1560_not
g58572 not n7131 ; n7131_not
g58573 not n5223 ; n5223_not
g58574 not n4800 ; n4800_not
g58575 not n1308 ; n1308_not
g58576 not n7221 ; n7221_not
g58577 not n1533 ; n1533_not
g58578 not n4206 ; n4206_not
g58579 not n8013 ; n8013_not
g58580 not n7500 ; n7500_not
g58581 not n2514 ; n2514_not
g58582 not n4350 ; n4350_not
g58583 not n3504 ; n3504_not
g58584 not n5007 ; n5007_not
g58585 not n1542 ; n1542_not
g58586 not n4116 ; n4116_not
g58587 not n1911 ; n1911_not
g58588 not n3621 ; n3621_not
g58589 not n5205 ; n5205_not
g58590 not n1902 ; n1902_not
g58591 not n4431 ; n4431_not
g58592 not n5241 ; n5241_not
g58593 not n7212 ; n7212_not
g58594 not n3324 ; n3324_not
g58595 not n5421 ; n5421_not
g58596 not n5250 ; n5250_not
g58597 not n7320 ; n7320_not
g58598 not n2433 ; n2433_not
g58599 not n6411 ; n6411_not
g58600 not n5412 ; n5412_not
g58601 not n5232 ; n5232_not
g58602 not n1830 ; n1830_not
g58603 not n3423 ; n3423_not
g58604 not n3801 ; n3801_not
g58605 not n4612 ; n4612_not
g58606 not n2272 ; n2272_not
g58607 not n2290 ; n2290_not
g58608 not n8212 ; n8212_not
g58609 not n8410 ; n8410_not
g58610 not n3073 ; n3073_not
g58611 not n1237 ; n1237_not
g58612 not n2506 ; n2506_not
g58613 not n3451 ; n3451_not
g58614 not n6322 ; n6322_not
g58615 not n9112 ; n9112_not
g58616 not n4720 ; n4720_not
g58617 not n2308 ; n2308_not
g58618 not n2191 ; n2191_not
g58619 not n4711 ; n4711_not
g58620 not n3325 ; n3325_not
g58621 not n4315 ; n4315_not
g58622 not n6007 ; n6007_not
g58623 not n2515 ; n2515_not
g58624 not n5620 ; n5620_not
g58625 not n6160 ; n6160_not
g58626 not n9130 ; n9130_not
g58627 not n4621 ; n4621_not
g58628 not n2281 ; n2281_not
g58629 not n8401 ; n8401_not
g58630 not n4630 ; n4630_not
g58631 not n2263 ; n2263_not
g58632 not n4027 ; n4027_not
g58633 not n4306 ; n4306_not
g58634 not n5611 ; n5611_not
g58635 not n3640 ; n3640_not
g58636 not n4108 ; n4108_not
g58637 not n3631 ; n3631_not
g58638 not n9211 ; n9211_not
g58639 not n8005 ; n8005_not
g58640 not n2425 ; n2425_not
g58641 not n6124 ; n6124_not
g58642 not n3118 ; n3118_not
g58643 not n4810 ; n4810_not
g58644 not n6214 ; n6214_not
g58645 not n8122 ; n8122_not
g58646 not n5413 ; n5413_not
g58647 not n3280 ; n3280_not
g58648 not n4801 ; n4801_not
g58649 not n4054 ; n4054_not
g58650 not n3703 ; n3703_not
g58651 not n9220 ; n9220_not
g58652 not n6070 ; n6070_not
g58653 not n5404 ; n5404_not
g58654 not n3712 ; n3712_not
g58655 not n9400 ; n9400_not
g58656 not n6151 ; n6151_not
g58657 not n2470 ; n2470_not
g58658 not n4513 ; n4513_not
g58659 not n6034 ; n6034_not
g58660 not n6142 ; n6142_not
g58661 not n2443 ; n2443_not
g58662 not n3217 ; n3217_not
g58663 not n4504 ; n4504_not
g58664 not n6061 ; n6061_not
g58665 not n3037 ; n3037_not
g58666 not n7033 ; n7033_not
g58667 not n2434 ; n2434_not
g58668 not n6133 ; n6133_not
g58669 not n3424 ; n3424_not
g58670 not n4072 ; n4072_not
g58671 not n5422 ; n5422_not
g58672 not n3271 ; n3271_not
g58673 not n2533 ; n2533_not
g58674 not n6232 ; n6232_not
g58675 not n4063 ; n4063_not
g58676 not n2650 ; n2650_not
g58677 not n2542 ; n2542_not
g58678 not n2614 ; n2614_not
g58679 not n8140 ; n8140_not
g58680 not n7006 ; n7006_not
g58681 not n3019 ; n3019_not
g58682 not n8131 ; n8131_not
g58683 not n2623 ; n2623_not
g58684 not n2551 ; n2551_not
g58685 not n6241 ; n6241_not
g58686 not n2641 ; n2641_not
g58687 not n3145 ; n3145_not
g58688 not n2560 ; n2560_not
g58689 not n6043 ; n6043_not
g58690 not n7024 ; n7024_not
g58691 not n6115 ; n6115_not
g58692 not n3208 ; n3208_not
g58693 not n7510 ; n7510_not
g58694 not n7501 ; n7501_not
g58695 not n3028 ; n3028_not
g58696 not n3262 ; n3262_not
g58697 not n2524 ; n2524_not
g58698 not n9040 ; n9040_not
g58699 not n6106 ; n6106_not
g58700 not n3721 ; n3721_not
g58701 not n8500 ; n8500_not
g58702 not n2380 ; n2380_not
g58703 not n4603 ; n4603_not
g58704 not n1093 ; n1093_not
g58705 not n2155 ; n2155_not
g58706 not n2371 ; n2371_not
g58707 not n8203 ; n8203_not
g58708 not n1084 ; n1084_not
g58709 not n9013 ; n9013_not
g58710 not n3307 ; n3307_not
g58711 not n2722 ; n2722_not
g58712 not n1075 ; n1075_not
g58713 not n3055 ; n3055_not
g58714 not n1066 ; n1066_not
g58715 not n3802 ; n3802_not
g58716 not n3226 ; n3226_not
g58717 not n1057 ; n1057_not
g58718 not n2182 ; n2182_not
g58719 not n6016 ; n6016_not
g58720 not n2317 ; n2317_not
g58721 not n4324 ; n4324_not
g58722 not n1147 ; n1147_not
g58723 not n7051 ; n7051_not
g58724 not n3163 ; n3163_not
g58725 not n2326 ; n2326_not
g58726 not n3244 ; n3244_not
g58727 not n1129 ; n1129_not
g58728 not n3316 ; n3316_not
g58729 not n2335 ; n2335_not
g58730 not n2344 ; n2344_not
g58731 not n2911 ; n2911_not
g58732 not n6025 ; n6025_not
g58733 not n2353 ; n2353_not
g58734 not n3064 ; n3064_not
g58735 not n4540 ; n4540_not
g58736 not n3109 ; n3109_not
g58737 not n6052 ; n6052_not
g58738 not n5710 ; n5710_not
g58739 not n6601 ; n6601_not
g58740 not n2452 ; n2452_not
g58741 not n4531 ; n4531_not
g58742 not n7042 ; n7042_not
g58743 not n3541 ; n3541_not
g58744 not n8113 ; n8113_not
g58745 not n4522 ; n4522_not
g58746 not n9121 ; n9121_not
g58747 not n1750 ; n1750_not
g58748 not n3811 ; n3811_not
g58749 not n1048 ; n1048_not
g58750 not n8023 ; n8023_not
g58751 not n1039 ; n1039_not
g58752 not n2407 ; n2407_not
g58753 not n8014 ; n8014_not
g58754 not n8104 ; n8104_not
g58755 not n9301 ; n9301_not
g58756 not n9202 ; n9202_not
g58757 not n2713 ; n2713_not
g58758 not n3046 ; n3046_not
g58759 not n3253 ; n3253_not
g58760 not n5701 ; n5701_not
g58761 not n4216 ; n4216_not
g58762 not n7123 ; n7123_not
g58763 not n1813 ; n1813_not
g58764 not n4225 ; n4225_not
g58765 not n4414 ; n4414_not
g58766 not n4207 ; n4207_not
g58767 not n4432 ; n4432_not
g58768 not n7114 ; n7114_not
g58769 not n1390 ; n1390_not
g58770 not n1903 ; n1903_not
g58771 not n3406 ; n3406_not
g58772 not n1732 ; n1732_not
g58773 not n5143 ; n5143_not
g58774 not n1912 ; n1912_not
g58775 not n1543 ; n1543_not
g58776 not n4234 ; n4234_not
g58777 not n5152 ; n5152_not
g58778 not n8320 ; n8320_not
g58779 not n7141 ; n7141_not
g58780 not n5431 ; n5431_not
g58781 not n4009 ; n4009_not
g58782 not n1561 ; n1561_not
g58783 not n4423 ; n4423_not
g58784 not n5134 ; n5134_not
g58785 not n8311 ; n8311_not
g58786 not n4243 ; n4243_not
g58787 not n1516 ; n1516_not
g58788 not n3370 ; n3370_not
g58789 not n4252 ; n4252_not
g58790 not n8050 ; n8050_not
g58791 not n9103 ; n9103_not
g58792 not n1507 ; n1507_not
g58793 not n6250 ; n6250_not
g58794 not n5116 ; n5116_not
g58795 not n3361 ; n3361_not
g58796 not n4261 ; n4261_not
g58797 not n3550 ; n3550_not
g58798 not n1930 ; n1930_not
g58799 not n1534 ; n1534_not
g58800 not n5602 ; n5602_not
g58801 not n6610 ; n6610_not
g58802 not n4126 ; n4126_not
g58803 not n1525 ; n1525_not
g58804 not n5161 ; n5161_not
g58805 not n1408 ; n1408_not
g58806 not n6700 ; n6700_not
g58807 not n1624 ; n1624_not
g58808 not n5053 ; n5053_not
g58809 not n4162 ; n4162_not
g58810 not n1651 ; n1651_not
g58811 not n8032 ; n8032_not
g58812 not n8041 ; n8041_not
g58813 not n9022 ; n9022_not
g58814 not n1723 ; n1723_not
g58815 not n1642 ; n1642_not
g58816 not n1714 ; n1714_not
g58817 not n5044 ; n5044_not
g58818 not n1705 ; n1705_not
g58819 not n4153 ; n4153_not
g58820 not n4351 ; n4351_not
g58821 not n4036 ; n4036_not
g58822 not n5062 ; n5062_not
g58823 not n1660 ; n1660_not
g58824 not n3505 ; n3505_not
g58825 not n1606 ; n1606_not
g58826 not n4081 ; n4081_not
g58827 not n1822 ; n1822_not
g58828 not n4441 ; n4441_not
g58829 not n4180 ; n4180_not
g58830 not n1831 ; n1831_not
g58831 not n4018 ; n4018_not
g58832 not n7132 ; n7132_not
g58833 not n8302 ; n8302_not
g58834 not n1840 ; n1840_not
g58835 not n3433 ; n3433_not
g58836 not n4171 ; n4171_not
g58837 not n3514 ; n3514_not
g58838 not n2920 ; n2920_not
g58839 not n5107 ; n5107_not
g58840 not n9031 ; n9031_not
g58841 not n3460 ; n3460_not
g58842 not n1462 ; n1462_not
g58843 not n3190 ; n3190_not
g58844 not n1291 ; n1291_not
g58845 not n3343 ; n3343_not
g58846 not n5026 ; n5026_not
g58847 not n5530 ; n5530_not
g58848 not n1309 ; n1309_not
g58849 not n1381 ; n1381_not
g58850 not n5071 ; n5071_not
g58851 not n8221 ; n8221_not
g58852 not n2074 ; n2074_not
g58853 not n5512 ; n5512_not
g58854 not n1417 ; n1417_not
g58855 not n5521 ; n5521_not
g58856 not n2083 ; n2083_not
g58857 not n3082 ; n3082_not
g58858 not n6205 ; n6205_not
g58859 not n3622 ; n3622_not
g58860 not n2092 ; n2092_not
g58861 not n3181 ; n3181_not
g58862 not n2164 ; n2164_not
g58863 not n2146 ; n2146_not
g58864 not n1354 ; n1354_not
g58865 not n2137 ; n2137_not
g58866 not n3091 ; n3091_not
g58867 not n4270 ; n4270_not
g58868 not n1336 ; n1336_not
g58869 not n3172 ; n3172_not
g58870 not n8230 ; n8230_not
g58871 not n3613 ; n3613_not
g58872 not n1345 ; n1345_not
g58873 not n1255 ; n1255_not
g58874 not n3604 ; n3604_not
g58875 not n5035 ; n5035_not
g58876 not n1318 ; n1318_not
g58877 not n1327 ; n1327_not
g58878 not n2119 ; n2119_not
g58879 not n1363 ; n1363_not
g58880 not n3334 ; n3334_not
g58881 not n1246 ; n1246_not
g58882 not n2128 ; n2128_not
g58883 not n1264 ; n1264_not
g58884 not n4117 ; n4117_not
g58885 not n1471 ; n1471_not
g58886 not n2236 ; n2236_not
g58887 not n5503 ; n5503_not
g58888 not n2227 ; n2227_not
g58889 not n2038 ; n2038_not
g58890 not n1435 ; n1435_not
g58891 not n2047 ; n2047_not
g58892 not n3352 ; n3352_not
g58893 not n3235 ; n3235_not
g58894 not n2254 ; n2254_not
g58895 not n7600 ; n7600_not
g58896 not n1480 ; n1480_not
g58897 not n2245 ; n2245_not
g58898 not n6304 ; n6304_not
g58899 not n2056 ; n2056_not
g58900 not n1444 ; n1444_not
g58901 not n1273 ; n1273_not
g58902 not n2209 ; n2209_not
g58903 not n2065 ; n2065_not
g58904 not n4271 ; n4271_not
g58905 not n9140 ; n9140_not
g58906 not n2534 ; n2534_not
g58907 not n9032 ; n9032_not
g58908 not n4631 ; n4631_not
g58909 not n3029 ; n3029_not
g58910 not n2660 ; n2660_not
g58911 not n9500 ; n9500_not
g58912 not n2921 ; n2921_not
g58913 not n3038 ; n3038_not
g58914 not n4163 ; n4163_not
g58915 not n4721 ; n4721_not
g58916 not n3146 ; n3146_not
g58917 not n9014 ; n9014_not
g58918 not n6350 ; n6350_not
g58919 not n6620 ; n6620_not
g58920 not n8510 ; n8510_not
g58921 not n7601 ; n7601_not
g58922 not n4262 ; n4262_not
g58923 not n7223 ; n7223_not
g58924 not n2543 ; n2543_not
g58925 not n2903 ; n2903_not
g58926 not n4145 ; n4145_not
g58927 not n6800 ; n6800_not
g58928 not n4064 ; n4064_not
g58929 not n4253 ; n4253_not
g58930 not n7700 ; n7700_not
g58931 not n6422 ; n6422_not
g58932 not n4451 ; n4451_not
g58933 not n6062 ; n6062_not
g58934 not n3227 ; n3227_not
g58935 not n6404 ; n6404_not
g58936 not n6710 ; n6710_not
g58937 not n4730 ; n4730_not
g58938 not n4235 ; n4235_not
g58939 not n4154 ; n4154_not
g58940 not n4325 ; n4325_not
g58941 not n3083 ; n3083_not
g58942 not n2516 ; n2516_not
g58943 not n2750 ; n2750_not
g58944 not n4226 ; n4226_not
g58945 not n2651 ; n2651_not
g58946 not n3119 ; n3119_not
g58947 not n4640 ; n4640_not
g58948 not n4244 ; n4244_not
g58949 not n2525 ; n2525_not
g58950 not n4460 ; n4460_not
g58951 not n2507 ; n2507_not
g58952 not n4352 ; n4352_not
g58953 not n7214 ; n7214_not
g58954 not n9122 ; n9122_not
g58955 not n2723 ; n2723_not
g58956 not n4082 ; n4082_not
g58957 not n6035 ; n6035_not
g58958 not n2822 ; n2822_not
g58959 not n6332 ; n6332_not
g58960 not n4424 ; n4424_not
g58961 not n9023 ; n9023_not
g58962 not n3074 ; n3074_not
g58963 not n6017 ; n6017_not
g58964 not n6044 ; n6044_not
g58965 not n7250 ; n7250_not
g58966 not n4217 ; n4217_not
g58967 not n3065 ; n3065_not
g58968 not n3047 ; n3047_not
g58969 not n6251 ; n6251_not
g58970 not n2831 ; n2831_not
g58971 not n7205 ; n7205_not
g58972 not n4703 ; n4703_not
g58973 not n7304 ; n7304_not
g58974 not n9230 ; n9230_not
g58975 not n9113 ; n9113_not
g58976 not n6701 ; n6701_not
g58977 not n2462 ; n2462_not
g58978 not n4037 ; n4037_not
g58979 not n3056 ; n3056_not
g58980 not n2804 ; n2804_not
g58981 not n4316 ; n4316_not
g58982 not n6026 ; n6026_not
g58983 not n4307 ; n4307_not
g58984 not n3182 ; n3182_not
g58985 not n3092 ; n3092_not
g58986 not n2714 ; n2714_not
g58987 not n4406 ; n4406_not
g58988 not n4280 ; n4280_not
g58989 not n3218 ; n3218_not
g58990 not n2813 ; n2813_not
g58991 not n4073 ; n4073_not
g58992 not n7610 ; n7610_not
g58993 not n6341 ; n6341_not
g58994 not n2930 ; n2930_not
g58995 not n4433 ; n4433_not
g58996 not n6413 ; n6413_not
g58997 not n3155 ; n3155_not
g58998 not n6611 ; n6611_not
g58999 not n2480 ; n2480_not
g59000 not n3173 ; n3173_not
g59001 not n4181 ; n4181_not
g59002 not n6242 ; n6242_not
g59003 not n7430 ; n7430_not
g59004 not n7511 ; n7511_not
g59005 not n4172 ; n4172_not
g59006 not n6314 ; n6314_not
g59007 not n8060 ; n8060_not
g59008 not n2741 ; n2741_not
g59009 not n7232 ; n7232_not
g59010 not n7322 ; n7322_not
g59011 not n6305 ; n6305_not
g59012 not n6602 ; n6602_not
g59013 not n2732 ; n2732_not
g59014 not n7520 ; n7520_not
g59015 not n4208 ; n4208_not
g59016 not n8501 ; n8501_not
g59017 not n7241 ; n7241_not
g59018 not n6008 ; n6008_not
g59019 not n6053 ; n6053_not
g59020 not n4361 ; n4361_not
g59021 not n8600 ; n8600_not
g59022 not n2624 ; n2624_not
g59023 not n2471 ; n2471_not
g59024 not n2840 ; n2840_not
g59025 not n7313 ; n7313_not
g59026 not n4190 ; n4190_not
g59027 not n2615 ; n2615_not
g59028 not n4442 ; n4442_not
g59029 not n5342 ; n5342_not
g59030 not n5063 ; n5063_not
g59031 not n3524 ; n3524_not
g59032 not n5351 ; n5351_not
g59033 not n1670 ; n1670_not
g59034 not n5360 ; n5360_not
g59035 not n1661 ; n1661_not
g59036 not n1607 ; n1607_not
g59037 not n1652 ; n1652_not
g59038 not n5054 ; n5054_not
g59039 not n5630 ; n5630_not
g59040 not n3506 ; n3506_not
g59041 not n5027 ; n5027_not
g59042 not n5432 ; n5432_not
g59043 not n3236 ; n3236_not
g59044 not n1634 ; n1634_not
g59045 not n1562 ; n1562_not
g59046 not n4046 ; n4046_not
g59047 not n1724 ; n1724_not
g59048 not n5423 ; n5423_not
g59049 not n1715 ; n1715_not
g59050 not n5324 ; n5324_not
g59051 not n1706 ; n1706_not
g59052 not n7142 ; n7142_not
g59053 not n5333 ; n5333_not
g59054 not n7412 ; n7412_not
g59055 not n3533 ; n3533_not
g59056 not n5072 ; n5072_not
g59057 not n7133 ; n7133_not
g59058 not n3425 ; n3425_not
g59059 not n1571 ; n1571_not
g59060 not n1553 ; n1553_not
g59061 not n9104 ; n9104_not
g59062 not n5441 ; n5441_not
g59063 not n7124 ; n7124_not
g59064 not n5315 ; n5315_not
g59065 not n3812 ; n3812_not
g59066 not n3434 ; n3434_not
g59067 not n3515 ; n3515_not
g59068 not n5621 ; n5621_not
g59069 not n1472 ; n1472_not
g59070 not n5405 ; n5405_not
g59071 not n1616 ; n1616_not
g59072 not n4019 ; n4019_not
g59073 not n5414 ; n5414_not
g59074 not n8114 ; n8114_not
g59075 not n3902 ; n3902_not
g59076 not n7151 ; n7151_not
g59077 not n9203 ; n9203_not
g59078 not n5252 ; n5252_not
g59079 not n8303 ; n8303_not
g59080 not n4091 ; n4091_not
g59081 not n3911 ; n3911_not
g59082 not n9212 ; n9212_not
g59083 not n5117 ; n5117_not
g59084 not n3443 ; n3443_not
g59085 not n7007 ; n7007_not
g59086 not n5261 ; n5261_not
g59087 not n3416 ; n3416_not
g59088 not n5216 ; n5216_not
g59089 not n8015 ; n8015_not
g59090 not n5225 ; n5225_not
g59091 not n5234 ; n5234_not
g59092 not n5243 ; n5243_not
g59093 not n8123 ; n8123_not
g59094 not n7421 ; n7421_not
g59095 not n8024 ; n8024_not
g59096 not n3470 ; n3470_not
g59097 not n3803 ; n3803_not
g59098 not n1760 ; n1760_not
g59099 not n1733 ; n1733_not
g59100 not n1751 ; n1751_not
g59101 not n5306 ; n5306_not
g59102 not n3551 ; n3551_not
g59103 not n3920 ; n3920_not
g59104 not n1643 ; n1643_not
g59105 not n9221 ; n9221_not
g59106 not n1805 ; n1805_not
g59107 not n5108 ; n5108_not
g59108 not n3560 ; n3560_not
g59109 not n5270 ; n5270_not
g59110 not n3461 ; n3461_not
g59111 not n5603 ; n5603_not
g59112 not n3614 ; n3614_not
g59113 not n1265 ; n1265_not
g59114 not n5513 ; n5513_not
g59115 not n1274 ; n1274_not
g59116 not n8222 ; n8222_not
g59117 not n1283 ; n1283_not
g59118 not n3623 ; n3623_not
g59119 not n5504 ; n5504_not
g59120 not n1373 ; n1373_not
g59121 not n5612 ; n5612_not
g59122 not n1238 ; n1238_not
g59123 not n3605 ; n3605_not
g59124 not n6521 ; n6521_not
g59125 not n8231 ; n8231_not
g59126 not n7403 ; n7403_not
g59127 not n1256 ; n1256_not
g59128 not n8033 ; n8033_not
g59129 not n5522 ; n5522_not
g59130 not n1058 ; n1058_not
g59131 not n3641 ; n3641_not
g59132 not n1166 ; n1166_not
g59133 not n1067 ; n1067_not
g59134 not n1157 ; n1157_not
g59135 not n1139 ; n1139_not
g59136 not n1076 ; n1076_not
g59137 not n1094 ; n1094_not
g59138 not n8204 ; n8204_not
g59139 not n3650 ; n3650_not
g59140 not n6440 ; n6440_not
g59141 not n6530 ; n6530_not
g59142 not n8213 ; n8213_not
g59143 not n1049 ; n1049_not
g59144 not n3632 ; n3632_not
g59145 not n1193 ; n1193_not
g59146 not n1184 ; n1184_not
g59147 not n6431 ; n6431_not
g59148 not n1175 ; n1175_not
g59149 not n1508 ; n1508_not
g59150 not n1418 ; n1418_not
g59151 not n8240 ; n8240_not
g59152 not n8420 ; n8420_not
g59153 not n1490 ; n1490_not
g59154 not n9320 ; n9320_not
g59155 not n1544 ; n1544_not
g59156 not n1535 ; n1535_not
g59157 not n7034 ; n7034_not
g59158 not n3722 ; n3722_not
g59159 not n1526 ; n1526_not
g59160 not n9131 ; n9131_not
g59161 not n1517 ; n1517_not
g59162 not n1409 ; n1409_not
g59163 not n6215 ; n6215_not
g59164 not n1427 ; n1427_not
g59165 not n6512 ; n6512_not
g59166 not n5180 ; n5180_not
g59167 not n6206 ; n6206_not
g59168 not n1391 ; n1391_not
g59169 not n1481 ; n1481_not
g59170 not n9401 ; n9401_not
g59171 not n6503 ; n6503_not
g59172 not n8105 ; n8105_not
g59173 not n9050 ; n9050_not
g59174 not n8411 ; n8411_not
g59175 not n5207 ; n5207_not
g59176 not n1445 ; n1445_not
g59177 not n6152 ; n6152_not
g59178 not n4811 ; n4811_not
g59179 not n7052 ; n7052_not
g59180 not n6143 ; n6143_not
g59181 not n2417 ; n2417_not
g59182 not n5720 ; n5720_not
g59183 not n4901 ; n4901_not
g59184 not n2390 ; n2390_not
g59185 not n4910 ; n4910_not
g59186 not n7043 ; n7043_not
g59187 not n6134 ; n6134_not
g59188 not n2381 ; n2381_not
g59189 not n4532 ; n4532_not
g59190 not n9041 ; n9041_not
g59191 not n4541 ; n4541_not
g59192 not n6161 ; n6161_not
g59193 not n2444 ; n2444_not
g59194 not n4550 ; n4550_not
g59195 not n2435 ; n2435_not
g59196 not n3191 ; n3191_not
g59197 not n4622 ; n4622_not
g59198 not n2336 ; n2336_not
g59199 not n2327 ; n2327_not
g59200 not n2318 ; n2318_not
g59201 not n5801 ; n5801_not
g59202 not n2309 ; n2309_not
g59203 not n4109 ; n4109_not
g59204 not n6116 ; n6116_not
g59205 not n2192 ; n2192_not
g59206 not n2372 ; n2372_not
g59207 not n4604 ; n4604_not
g59208 not n3731 ; n3731_not
g59209 not n9410 ; n9410_not
g59210 not n4613 ; n4613_not
g59211 not n8141 ; n8141_not
g59212 not n2354 ; n2354_not
g59213 not n2165 ; n2165_not
g59214 not n6125 ; n6125_not
g59215 not n2345 ; n2345_not
g59216 not n7016 ; n7016_not
g59217 not n6224 ; n6224_not
g59218 not n2570 ; n2570_not
g59219 not n7331 ; n7331_not
g59220 not n2561 ; n2561_not
g59221 not n4523 ; n4523_not
g59222 not n2552 ; n2552_not
g59223 not n4514 ; n4514_not
g59224 not n2633 ; n2633_not
g59225 not n6260 ; n6260_not
g59226 not n6071 ; n6071_not
g59227 not n6080 ; n6080_not
g59228 not n2453 ; n2453_not
g59229 not n4505 ; n4505_not
g59230 not n2408 ; n2408_not
g59231 not n6107 ; n6107_not
g59232 not n7340 ; n7340_not
g59233 not n8132 ; n8132_not
g59234 not n4127 ; n4127_not
g59235 not n5126 ; n5126_not
g59236 not n8150 ; n8150_not
g59237 not n8330 ; n8330_not
g59238 not n5144 ; n5144_not
g59239 not n2084 ; n2084_not
g59240 not n5009 ; n5009_not
g59241 not n2075 ; n2075_not
g59242 not n4118 ; n4118_not
g59243 not n2066 ; n2066_not
g59244 not n2057 ; n2057_not
g59245 not n5081 ; n5081_not
g59246 not n2048 ; n2048_not
g59247 not n5711 ; n5711_not
g59248 not n1931 ; n1931_not
g59249 not n1922 ; n1922_not
g59250 not n8321 ; n8321_not
g59251 not n3407 ; n3407_not
g59252 not n8312 ; n8312_not
g59253 not n5702 ; n5702_not
g59254 not n5153 ; n5153_not
g59255 not n4136 ; n4136_not
g59256 not n7106 ; n7106_not
g59257 not n5162 ; n5162_not
g59258 not n1940 ; n1940_not
g59259 not n2255 ; n2255_not
g59260 not n7061 ; n7061_not
g59261 not n2246 ; n2246_not
g59262 not n2237 ; n2237_not
g59263 not n2219 ; n2219_not
g59264 not n2093 ; n2093_not
g59265 not n2291 ; n2291_not
g59266 not n2282 ; n2282_not
g59267 not n2273 ; n2273_not
g59268 not n2264 ; n2264_not
g59269 not n2138 ; n2138_not
g59270 not n2129 ; n2129_not
g59271 not n5045 ; n5045_not
g59272 not n5018 ; n5018_not
g59273 not n2174 ; n2174_not
g59274 not n3705 ; n3705_not
g59275 not n3147 ; n3147_not
g59276 not n3525 ; n3525_not
g59277 not n3534 ; n3534_not
g59278 not n3804 ; n3804_not
g59279 not n3741 ; n3741_not
g59280 not n3444 ; n3444_not
g59281 not n3831 ; n3831_not
g59282 not n3435 ; n3435_not
g59283 not n7350 ; n7350_not
g59284 not n3165 ; n3165_not
g59285 not n7332 ; n7332_not
g59286 not n3813 ; n3813_not
g59287 not n6621 ; n6621_not
g59288 not n3426 ; n3426_not
g59289 not n7341 ; n7341_not
g59290 not n3543 ; n3543_not
g59291 not n3723 ; n3723_not
g59292 not n3714 ; n3714_not
g59293 not n6612 ; n6612_not
g59294 not n3354 ; n3354_not
g59295 not n6702 ; n6702_not
g59296 not n6333 ; n6333_not
g59297 not n3363 ; n3363_not
g59298 not n6720 ; n6720_not
g59299 not n6360 ; n6360_not
g59300 not n4128 ; n4128_not
g59301 not n3372 ; n3372_not
g59302 not n3840 ; n3840_not
g59303 not n3156 ; n3156_not
g59304 not n3381 ; n3381_not
g59305 not n3390 ; n3390_not
g59306 not n4119 ; n4119_not
g59307 not n6450 ; n6450_not
g59308 not n3417 ; n3417_not
g59309 not n7413 ; n7413_not
g59310 not n4083 ; n4083_not
g59311 not n3345 ; n3345_not
g59312 not n4074 ; n4074_not
g59313 not n3453 ; n3453_not
g59314 not n3336 ; n3336_not
g59315 not n3264 ; n3264_not
g59316 not n4092 ; n4092_not
g59317 not n3912 ; n3912_not
g59318 not n3273 ; n3273_not
g59319 not n6342 ; n6342_not
g59320 not n3282 ; n3282_not
g59321 not n3903 ; n3903_not
g59322 not n6711 ; n6711_not
g59323 not n3291 ; n3291_not
g59324 not n3255 ; n3255_not
g59325 not n8601 ; n8601_not
g59326 not n7530 ; n7530_not
g59327 not n6432 ; n6432_not
g59328 not n3192 ; n3192_not
g59329 not n3309 ; n3309_not
g59330 not n3921 ; n3921_not
g59331 not n3930 ; n3930_not
g59332 not n6441 ; n6441_not
g59333 not n3228 ; n3228_not
g59334 not n3327 ; n3327_not
g59335 not n8610 ; n8610_not
g59336 not n3183 ; n3183_not
g59337 not n3237 ; n3237_not
g59338 not n6351 ; n6351_not
g59339 not n8700 ; n8700_not
g59340 not n3318 ; n3318_not
g59341 not n3246 ; n3246_not
g59342 not n6252 ; n6252_not
g59343 not n8421 ; n8421_not
g59344 not n3732 ; n3732_not
g59345 not n7305 ; n7305_not
g59346 not n6216 ; n6216_not
g59347 not n7521 ; n7521_not
g59348 not n7314 ; n7314_not
g59349 not n6504 ; n6504_not
g59350 not n3480 ; n3480_not
g59351 not n6513 ; n6513_not
g59352 not n6207 ; n6207_not
g59353 not n3471 ; n3471_not
g59354 not n6522 ; n6522_not
g59355 not n6531 ; n6531_not
g59356 not n6540 ; n6540_not
g59357 not n7323 ; n7323_not
g59358 not n6180 ; n6180_not
g59359 not n7260 ; n7260_not
g59360 not n4056 ; n4056_not
g59361 not n8430 ; n8430_not
g59362 not n4038 ; n4038_not
g59363 not n6225 ; n6225_not
g59364 not n9420 ; n9420_not
g59365 not n7404 ; n7404_not
g59366 not n3516 ; n3516_not
g59367 not n4029 ; n4029_not
g59368 not n1770 ; n1770_not
g59369 not n1707 ; n1707_not
g59370 not n7620 ; n7620_not
g59371 not n1716 ; n1716_not
g59372 not n1725 ; n1725_not
g59373 not n1752 ; n1752_not
g59374 not n7017 ; n7017_not
g59375 not n7143 ; n7143_not
g59376 not n5307 ; n5307_not
g59377 not n8034 ; n8034_not
g59378 not n5316 ; n5316_not
g59379 not n1572 ; n1572_not
g59380 not n5082 ; n5082_not
g59381 not n9060 ; n9060_not
g59382 not n4920 ; n4920_not
g59383 not n1644 ; n1644_not
g59384 not n1653 ; n1653_not
g59385 not n7422 ; n7422_not
g59386 not n5109 ; n5109_not
g59387 not n1662 ; n1662_not
g59388 not n7152 ; n7152_not
g59389 not n1671 ; n1671_not
g59390 not n5271 ; n5271_not
g59391 not n1680 ; n1680_not
g59392 not n7170 ; n7170_not
g59393 not n5280 ; n5280_not
g59394 not n8025 ; n8025_not
g59395 not n1635 ; n1635_not
g59396 not n1617 ; n1617_not
g59397 not n5406 ; n5406_not
g59398 not n1464 ; n1464_not
g59399 not n8250 ; n8250_not
g59400 not n1482 ; n1482_not
g59401 not n1608 ; n1608_not
g59402 not n1491 ; n1491_not
g59403 not n1509 ; n1509_not
g59404 not n7800 ; n7800_not
g59405 not n9213 ; n9213_not
g59406 not n1518 ; n1518_not
g59407 not n1527 ; n1527_not
g59408 not n1581 ; n1581_not
g59409 not n1536 ; n1536_not
g59410 not n5424 ; n5424_not
g59411 not n5325 ; n5325_not
g59412 not n2382 ; n2382_not
g59413 not n5073 ; n5073_not
g59414 not n5334 ; n5334_not
g59415 not n7611 ; n7611_not
g59416 not n7134 ; n7134_not
g59417 not n5343 ; n5343_not
g59418 not n5064 ; n5064_not
g59419 not n8043 ; n8043_not
g59420 not n5352 ; n5352_not
g59421 not n9204 ; n9204_not
g59422 not n7206 ; n7206_not
g59423 not n5361 ; n5361_not
g59424 not n5019 ; n5019_not
g59425 not n5028 ; n5028_not
g59426 not n5370 ; n5370_not
g59427 not n5046 ; n5046_not
g59428 not n9132 ; n9132_not
g59429 not n7431 ; n7431_not
g59430 not n5154 ; n5154_not
g59431 not n4821 ; n4821_not
g59432 not n1905 ; n1905_not
g59433 not n5163 ; n5163_not
g59434 not n1950 ; n1950_not
g59435 not n4830 ; n4830_not
g59436 not n1914 ; n1914_not
g59437 not n5181 ; n5181_not
g59438 not n1941 ; n1941_not
g59439 not n9141 ; n9141_not
g59440 not n1923 ; n1923_not
g59441 not n8322 ; n8322_not
g59442 not n5190 ; n5190_not
g59443 not n9114 ; n9114_not
g59444 not n5091 ; n5091_not
g59445 not n8340 ; n8340_not
g59446 not n8007 ; n8007_not
g59447 not n9123 ; n9123_not
g59448 not n1824 ; n1824_not
g59449 not n9042 ; n9042_not
g59450 not n1833 ; n1833_not
g59451 not n5118 ; n5118_not
g59452 not n1842 ; n1842_not
g59453 not n1851 ; n1851_not
g59454 not n1860 ; n1860_not
g59455 not n5136 ; n5136_not
g59456 not n8331 ; n8331_not
g59457 not n9051 ; n9051_not
g59458 not n5244 ; n5244_not
g59459 not n4902 ; n4902_not
g59460 not n8304 ; n8304_not
g59461 not n5253 ; n5253_not
g59462 not n4911 ; n4911_not
g59463 not n5262 ; n5262_not
g59464 not n1806 ; n1806_not
g59465 not n1761 ; n1761_not
g59466 not n7116 ; n7116_not
g59467 not n5208 ; n5208_not
g59468 not n8313 ; n8313_not
g59469 not n6810 ; n6810_not
g59470 not n9150 ; n9150_not
g59471 not n5217 ; n5217_not
g59472 not n6801 ; n6801_not
g59473 not n5226 ; n5226_not
g59474 not n5235 ; n5235_not
g59475 not n5127 ; n5127_not
g59476 not n1077 ; n1077_not
g59477 not n1068 ; n1068_not
g59478 not n1059 ; n1059_not
g59479 not n7107 ; n7107_not
g59480 not n5901 ; n5901_not
g59481 not n9312 ; n9312_not
g59482 not n8106 ; n8106_not
g59483 not n9321 ; n9321_not
g59484 not n9330 ; n9330_not
g59485 not n5442 ; n5442_not
g59486 not n5433 ; n5433_not
g59487 not n1239 ; n1239_not
g59488 not n1095 ; n1095_not
g59489 not n1194 ; n1194_not
g59490 not n1185 ; n1185_not
g59491 not n1176 ; n1176_not
g59492 not n1167 ; n1167_not
g59493 not n7251 ; n7251_not
g59494 not n1158 ; n1158_not
g59495 not n1149 ; n1149_not
g59496 not n8205 ; n8205_not
g59497 not n1086 ; n1086_not
g59498 not n7710 ; n7710_not
g59499 not n8151 ; n8151_not
g59500 not n7053 ; n7053_not
g59501 not n7701 ; n7701_not
g59502 not n9411 ; n9411_not
g59503 not n8142 ; n8142_not
g59504 not n9105 ; n9105_not
g59505 not n5811 ; n5811_not
g59506 not n9600 ; n9600_not
g59507 not n8133 ; n8133_not
g59508 not n8115 ; n8115_not
g59509 not n9240 ; n9240_not
g59510 not n9231 ; n9231_not
g59511 not n9222 ; n9222_not
g59512 not n7044 ; n7044_not
g59513 not n8124 ; n8124_not
g59514 not n8160 ; n8160_not
g59515 not n7062 ; n7062_not
g59516 not n1419 ; n1419_not
g59517 not n1455 ; n1455_not
g59518 not n7224 ; n7224_not
g59519 not n1428 ; n1428_not
g59520 not n1446 ; n1446_not
g59521 not n1437 ; n1437_not
g59522 not n1329 ; n1329_not
g59523 not n1338 ; n1338_not
g59524 not n1545 ; n1545_not
g59525 not n7215 ; n7215_not
g59526 not n1374 ; n1374_not
g59527 not n5451 ; n5451_not
g59528 not n8241 ; n8241_not
g59529 not n1356 ; n1356_not
g59530 not n1347 ; n1347_not
g59531 not n1266 ; n1266_not
g59532 not n5514 ; n5514_not
g59533 not n1275 ; n1275_not
g59534 not n8223 ; n8223_not
g59535 not n1284 ; n1284_not
g59536 not n7242 ; n7242_not
g59537 not n1248 ; n1248_not
g59538 not n8214 ; n8214_not
g59539 not n5523 ; n5523_not
g59540 not n1365 ; n1365_not
g59541 not n5532 ; n5532_not
g59542 not n1392 ; n1392_not
g59543 not n8070 ; n8070_not
g59544 not n8232 ; n8232_not
g59545 not n5550 ; n5550_not
g59546 not n7233 ; n7233_not
g59547 not n2850 ; n2850_not
g59548 not n2724 ; n2724_not
g59549 not n5802 ; n5802_not
g59550 not n4443 ; n4443_not
g59551 not n2940 ; n2940_not
g59552 not n9006 ; n9006_not
g59553 not n2409 ; n2409_not
g59554 not n4452 ; n4452_not
g59555 not n2427 ; n2427_not
g59556 not n2715 ; n2715_not
g59557 not n4371 ; n4371_not
g59558 not n6261 ; n6261_not
g59559 not n2445 ; n2445_not
g59560 not n2454 ; n2454_not
g59561 not n2247 ; n2247_not
g59562 not n2832 ; n2832_not
g59563 not n6405 ; n6405_not
g59564 not n2733 ; n2733_not
g59565 not n4740 ; n4740_not
g59566 not n4362 ; n4362_not
g59567 not n2157 ; n2157_not
g59568 not n2364 ; n2364_not
g59569 not n4434 ; n4434_not
g59570 not n4353 ; n4353_not
g59571 not n2931 ; n2931_not
g59572 not n2841 ; n2841_not
g59573 not n9033 ; n9033_not
g59574 not n2616 ; n2616_not
g59575 not n7026 ; n7026_not
g59576 not n7503 ; n7503_not
g59577 not n4713 ; n4713_not
g59578 not n6630 ; n6630_not
g59579 not n2670 ; n2670_not
g59580 not n2913 ; n2913_not
g59581 not n6234 ; n6234_not
g59582 not n2661 ; n2661_not
g59583 not n2607 ; n2607_not
g59584 not n2643 ; n2643_not
g59585 not n4137 ; n4137_not
g59586 not n9024 ; n9024_not
g59587 not n2625 ; n2625_not
g59588 not n4731 ; n4731_not
g59589 not n8511 ; n8511_not
g59590 not n6900 ; n6900_not
g59591 not n4416 ; n4416_not
g59592 not n2418 ; n2418_not
g59593 not n4803 ; n4803_not
g59594 not n2148 ; n2148_not
g59595 not n6414 ; n6414_not
g59596 not n6315 ; n6315_not
g59597 not n2166 ; n2166_not
g59598 not n2184 ; n2184_not
g59599 not n2751 ; n2751_not
g59600 not n6270 ; n6270_not
g59601 not n4704 ; n4704_not
g59602 not n4047 ; n4047_not
g59603 not n2229 ; n2229_not
g59604 not n2238 ; n2238_not
g59605 not n6306 ; n6306_not
g59606 not n6423 ; n6423_not
g59607 not n9015 ; n9015_not
g59608 not n7071 ; n7071_not
g59609 not n4407 ; n4407_not
g59610 not n2805 ; n2805_not
g59611 not n2760 ; n2760_not
g59612 not n2742 ; n2742_not
g59613 not n8403 ; n8403_not
g59614 not n2634 ; n2634_not
g59615 not n2823 ; n2823_not
g59616 not n2904 ; n2904_not
g59617 not n2175 ; n2175_not
g59618 not n2814 ; n2814_not
g59619 not n4507 ; n4507_not
g59620 not n4444 ; n4444_not
g59621 not n4561 ; n4561_not
g59622 not n5605 ; n5605_not
g59623 not n4462 ; n4462_not
g59624 not n8053 ; n8053_not
g59625 not n5551 ; n5551_not
g59626 not n6307 ; n6307_not
g59627 not n5164 ; n5164_not
g59628 not n5533 ; n5533_not
g59629 not n5227 ; n5227_not
g59630 not n5245 ; n5245_not
g59631 not n5209 ; n5209_not
g59632 not n5614 ; n5614_not
g59633 not n6316 ; n6316_not
g59634 not n8404 ; n8404_not
g59635 not n4525 ; n4525_not
g59636 not n4534 ; n4534_not
g59637 not n5560 ; n5560_not
g59638 not n4417 ; n4417_not
g59639 not n5254 ; n5254_not
g59640 not n5182 ; n5182_not
g59641 not n5218 ; n5218_not
g59642 not n5524 ; n5524_not
g59643 not n8080 ; n8080_not
g59644 not n4552 ; n4552_not
g59645 not n7810 ; n7810_not
g59646 not n4480 ; n4480_not
g59647 not n5191 ; n5191_not
g59648 not n4453 ; n4453_not
g59649 not n8215 ; n8215_not
g59650 not n4516 ; n4516_not
g59651 not n4237 ; n4237_not
g59652 not n3940 ; n3940_not
g59653 not n4408 ; n4408_not
g59654 not n4543 ; n4543_not
g59655 not n4570 ; n4570_not
g59656 not n4831 ; n4831_not
g59657 not n5236 ; n5236_not
g59658 not n8224 ; n8224_not
g59659 not n6532 ; n6532_not
g59660 not n5407 ; n5407_not
g59661 not n8125 ; n8125_not
g59662 not n3580 ; n3580_not
g59663 not n3571 ; n3571_not
g59664 not n6541 ; n6541_not
g59665 not n4039 ; n4039_not
g59666 not n4309 ; n4309_not
g59667 not n8161 ; n8161_not
g59668 not n8008 ; n8008_not
g59669 not n6604 ; n6604_not
g59670 not n3562 ; n3562_not
g59671 not n4318 ; n4318_not
g59672 not n5380 ; n5380_not
g59673 not n3553 ; n3553_not
g59674 not n4327 ; n4327_not
g59675 not n5740 ; n5740_not
g59676 not n5371 ; n5371_not
g59677 not n8116 ; n8116_not
g59678 not n4345 ; n4345_not
g59679 not n5821 ; n5821_not
g59680 not n3661 ; n3661_not
g59681 not n6514 ; n6514_not
g59682 not n3652 ; n3652_not
g59683 not n3751 ; n3751_not
g59684 not n3643 ; n3643_not
g59685 not n8134 ; n8134_not
g59686 not n4264 ; n4264_not
g59687 not n3634 ; n3634_not
g59688 not n5803 ; n5803_not
g59689 not n3625 ; n3625_not
g59690 not n6262 ; n6262_not
g59691 not n4255 ; n4255_not
g59692 not n3616 ; n3616_not
g59693 not n4273 ; n4273_not
g59694 not n6523 ; n6523_not
g59695 not n8143 ; n8143_not
g59696 not n3607 ; n3607_not
g59697 not n4057 ; n4057_not
g59698 not n4282 ; n4282_not
g59699 not n4048 ; n4048_not
g59700 not n4291 ; n4291_not
g59701 not n8152 ; n8152_not
g59702 not n3832 ; n3832_not
g59703 not n5317 ; n5317_not
g59704 not n5308 ; n5308_not
g59705 not n4381 ; n4381_not
g59706 not n6280 ; n6280_not
g59707 not n5290 ; n5290_not
g59708 not n5650 ; n5650_not
g59709 not n5281 ; n5281_not
g59710 not n5911 ; n5911_not
g59711 not n4426 ; n4426_not
g59712 not n5641 ; n5641_not
g59713 not n7450 ; n7450_not
g59714 not n6190 ; n6190_not
g59715 not n7801 ; n7801_not
g59716 not n5272 ; n5272_not
g59717 not n5632 ; n5632_not
g59718 not n5263 ; n5263_not
g59719 not n3841 ; n3841_not
g59720 not n5623 ; n5623_not
g59721 not n8206 ; n8206_not
g59722 not n5731 ; n5731_not
g59723 not n5362 ; n5362_not
g59724 not n8170 ; n8170_not
g59725 not n5722 ; n5722_not
g59726 not n5434 ; n5434_not
g59727 not n3814 ; n3814_not
g59728 not n5353 ; n5353_not
g59729 not n5713 ; n5713_not
g59730 not n5344 ; n5344_not
g59731 not n6550 ; n6550_not
g59732 not n4246 ; n4246_not
g59733 not n5704 ; n5704_not
g59734 not n7504 ; n7504_not
g59735 not n4354 ; n4354_not
g59736 not n8107 ; n8107_not
g59737 not n5443 ; n5443_not
g59738 not n5335 ; n5335_not
g59739 not n3544 ; n3544_not
g59740 not n4363 ; n4363_not
g59741 not n5452 ; n5452_not
g59742 not n5326 ; n5326_not
g59743 not n7360 ; n7360_not
g59744 not n6271 ; n6271_not
g59745 not n4750 ; n4750_not
g59746 not n3913 ; n3913_not
g59747 not n6136 ; n6136_not
g59748 not n4093 ; n4093_not
g59749 not n5119 ; n5119_not
g59750 not n4912 ; n4912_not
g59751 not n3904 ; n3904_not
g59752 not n7711 ; n7711_not
g59753 not n4903 ; n4903_not
g59754 not n4741 ; n4741_not
g59755 not n8305 ; n8305_not
g59756 not n4183 ; n4183_not
g59757 not n5128 ; n5128_not
g59758 not n5137 ; n5137_not
g59759 not n8017 ; n8017_not
g59760 not n6127 ; n6127_not
g59761 not n7900 ; n7900_not
g59762 not n5812 ; n5812_not
g59763 not n6046 ; n6046_not
g59764 not n8233 ; n8233_not
g59765 not n8413 ; n8413_not
g59766 not n6118 ; n6118_not
g59767 not n8242 ; n8242_not
g59768 not n7621 ; n7621_not
g59769 not n6028 ; n6028_not
g59770 not n4066 ; n4066_not
g59771 not n8440 ; n8440_not
g59772 not n6163 ; n6163_not
g59773 not n6154 ; n6154_not
g59774 not n8431 ; n8431_not
g59775 not n4930 ; n4930_not
g59776 not n6145 ; n6145_not
g59777 not n3931 ; n3931_not
g59778 not n7720 ; n7720_not
g59779 not n4192 ; n4192_not
g59780 not n3922 ; n3922_not
g59781 not n4084 ; n4084_not
g59782 not n7630 ; n7630_not
g59783 not n6037 ; n6037_not
g59784 not n4921 ; n4921_not
g59785 not n6064 ; n6064_not
g59786 not n3850 ; n3850_not
g59787 not n4129 ; n4129_not
g59788 not n6091 ; n6091_not
g59789 not n4147 ; n4147_not
g59790 not n1942 ; n1942_not
g59791 not n5047 ; n5047_not
g59792 not n4156 ; n4156_not
g59793 not n4165 ; n4165_not
g59794 not n6073 ; n6073_not
g59795 not n5056 ; n5056_not
g59796 not n8332 ; n8332_not
g59797 not n5083 ; n5083_not
g59798 not n5074 ; n5074_not
g59799 not n8323 ; n8323_not
g59800 not n8314 ; n8314_not
g59801 not n6082 ; n6082_not
g59802 not n7423 ; n7423_not
g59803 not n9700 ; n9700_not
g59804 not n6109 ; n6109_not
g59805 not n8251 ; n8251_not
g59806 not n7702 ; n7702_not
g59807 not n4714 ; n4714_not
g59808 not n8260 ; n8260_not
g59809 not n6055 ; n6055_not
g59810 not n4840 ; n4840_not
g59811 not n4822 ; n4822_not
g59812 not n4174 ; n4174_not
g59813 not n4705 ; n4705_not
g59814 not n5146 ; n5146_not
g59815 not n4138 ; n4138_not
g59816 not n4372 ; n4372_not
g59817 not n4642 ; n4642_not
g59818 not n3706 ; n3706_not
g59819 not n4651 ; n4651_not
g59820 not n5461 ; n5461_not
g59821 not n6226 ; n6226_not
g59822 not n4660 ; n4660_not
g59823 not n8062 ; n8062_not
g59824 not n5506 ; n5506_not
g59825 not n3742 ; n3742_not
g59826 not n7405 ; n7405_not
g59827 not n3733 ; n3733_not
g59828 not n4606 ; n4606_not
g59829 not n6217 ; n6217_not
g59830 not n4615 ; n4615_not
g59831 not n4624 ; n4624_not
g59832 not n5902 ; n5902_not
g59833 not n4633 ; n4633_not
g59834 not n4228 ; n4228_not
g59835 not n3724 ; n3724_not
g59836 not n7180 ; n7180_not
g59837 not n8503 ; n8503_not
g59838 not n8035 ; n8035_not
g59839 not n7603 ; n7603_not
g59840 not n6235 ; n6235_not
g59841 not n4804 ; n4804_not
g59842 not n9421 ; n9421_not
g59843 not n5092 ; n5092_not
g59844 not n7612 ; n7612_not
g59845 not n6019 ; n6019_not
g59846 not n8521 ; n8521_not
g59847 not n7414 ; n7414_not
g59848 not n5416 ; n5416_not
g59849 not n6244 ; n6244_not
g59850 not n4723 ; n4723_not
g59851 not n4219 ; n4219_not
g59852 not n8044 ; n8044_not
g59853 not n1366 ; n1366_not
g59854 not n7063 ; n7063_not
g59855 not n2518 ; n2518_not
g59856 not n6370 ; n6370_not
g59857 not n3238 ; n3238_not
g59858 not n1276 ; n1276_not
g59859 not n2482 ; n2482_not
g59860 not n2347 ; n2347_not
g59861 not n3265 ; n3265_not
g59862 not n1456 ; n1456_not
g59863 not n7108 ; n7108_not
g59864 not n7252 ; n7252_not
g59865 not n3274 ; n3274_not
g59866 not n1924 ; n1924_not
g59867 not n9313 ; n9313_not
g59868 not n1393 ; n1393_not
g59869 not n3292 ; n3292_not
g59870 not n2626 ; n2626_not
g59871 not n2149 ; n2149_not
g59872 not n2608 ; n2608_not
g59873 not n1285 ; n1285_not
g59874 not n7531 ; n7531_not
g59875 not n2833 ; n2833_not
g59876 not n3490 ; n3490_not
g59877 not n6640 ; n6640_not
g59878 not n6352 ; n6352_not
g59879 not n1906 ; n1906_not
g59880 not n7207 ; n7207_not
g59881 not n3517 ; n3517_not
g59882 not n1348 ; n1348_not
g59883 not n1357 ; n1357_not
g59884 not n2950 ; n2950_not
g59885 not n1753 ; n1753_not
g59886 not n2851 ; n2851_not
g59887 not n2257 ; n2257_not
g59888 not n1780 ; n1780_not
g59889 not n3247 ; n3247_not
g59890 not n7243 ; n7243_not
g59891 not n1339 ; n1339_not
g59892 not n2167 ; n2167_not
g59893 not n7117 ; n7117_not
g59894 not n1375 ; n1375_not
g59895 not n1681 ; n1681_not
g59896 not n2842 ; n2842_not
g59897 not n2725 ; n2725_not
g59898 not n3256 ; n3256_not
g59899 not n6361 ; n6361_not
g59900 not n2248 ; n2248_not
g59901 not n3193 ; n3193_not
g59902 not n1915 ; n1915_not
g59903 not n2419 ; n2419_not
g59904 not n2365 ; n2365_not
g59905 not n6406 ; n6406_not
g59906 not n2815 ; n2815_not
g59907 not n1195 ; n1195_not
g59908 not n2635 ; n2635_not
g59909 not n1555 ; n1555_not
g59910 not n6415 ; n6415_not
g59911 not n1186 ; n1186_not
g59912 not n1168 ; n1168_not
g59913 not n7171 ; n7171_not
g59914 not n2077 ; n2077_not
g59915 not n7333 ; n7333_not
g59916 not n1564 ; n1564_not
g59917 not n2644 ; n2644_not
g59918 not n1177 ; n1177_not
g59919 not n2806 ; n2806_not
g59920 not n1960 ; n1960_not
g59921 not n6424 ; n6424_not
g59922 not n7315 ; n7315_not
g59923 not n7036 ; n7036_not
g59924 not n7153 ; n7153_not
g59925 not n6712 ; n6712_not
g59926 not n2356 ; n2356_not
g59927 not n1258 ; n1258_not
g59928 not n3283 ; n3283_not
g59929 not n9340 ; n9340_not
g59930 not n7009 ; n7009_not
g59931 not n1690 ; n1690_not
g59932 not n2068 ; n2068_not
g59933 not n2473 ; n2473_not
g59934 not n7324 ; n7324_not
g59935 not n7018 ; n7018_not
g59936 not n3481 ; n3481_not
g59937 not n2059 ; n2059_not
g59938 not n2824 ; n2824_not
g59939 not n1843 ; n1843_not
g59940 not n6721 ; n6721_not
g59941 not n1645 ; n1645_not
g59942 not n1447 ; n1447_not
g59943 not n6334 ; n6334_not
g59944 not n3418 ; n3418_not
g59945 not n7225 ; n7225_not
g59946 not n3364 ; n3364_not
g59947 not n2905 ; n2905_not
g59948 not n7351 ; n7351_not
g59949 not n1852 ; n1852_not
g59950 not n7216 ; n7216_not
g59951 not n3436 ; n3436_not
g59952 not n6622 ; n6622_not
g59953 not n3355 ; n3355_not
g59954 not n9520 ; n9520_not
g59955 not n3166 ; n3166_not
g59956 not n1654 ; n1654_not
g59957 not n2428 ; n2428_not
g59958 not n2581 ; n2581_not
g59959 not n1429 ; n1429_not
g59960 not n6343 ; n6343_not
g59961 not n3373 ; n3373_not
g59962 not n6730 ; n6730_not
g59963 not n1636 ; n1636_not
g59964 not n1825 ; n1825_not
g59965 not n1807 ; n1807_not
g59966 not n9601 ; n9601_not
g59967 not n1474 ; n1474_not
g59968 not n3382 ; n3382_not
g59969 not n7306 ; n7306_not
g59970 not n3148 ; n3148_not
g59971 not n1465 ; n1465_not
g59972 not n3157 ; n3157_not
g59973 not n1438 ; n1438_not
g59974 not n1834 ; n1834_not
g59975 not n3391 ; n3391_not
g59976 not n2383 ; n2383_not
g59977 not n2923 ; n2923_not
g59978 not n6505 ; n6505_not
g59979 not n7126 ; n7126_not
g59980 not n3328 ; n3328_not
g59981 not n1771 ; n1771_not
g59982 not n2338 ; n2338_not
g59983 not n2491 ; n2491_not
g59984 not n7234 ; n7234_not
g59985 not n6631 ; n6631_not
g59986 not n1762 ; n1762_not
g59987 not n2941 ; n2941_not
g59988 not n3508 ; n3508_not
g59989 not n3319 ; n3319_not
g59990 not n2860 ; n2860_not
g59991 not n2266 ; n2266_not
g59992 not n2185 ; n2185_not
g59993 not n2284 ; n2284_not
g59994 not n1249 ; n1249_not
g59995 not n3445 ; n3445_not
g59996 not n7144 ; n7144_not
g59997 not n2509 ; n2509_not
g59998 not n2275 ; n2275_not
g59999 not n1861 ; n1861_not
g60000 not n2176 ; n2176_not
g60001 not n1663 ; n1663_not
g60002 not n3346 ; n3346_not
g60003 not n2329 ; n2329_not
g60004 not n2590 ; n2590_not
g60005 not n1870 ; n1870_not
g60006 not n3463 ; n3463_not
g60007 not n3337 ; n3337_not
g60008 not n1672 ; n1672_not
g60009 not n7540 ; n7540_not
g60010 not n9610 ; n9610_not
g60011 not n7513 ; n7513_not
g60012 not n7054 ; n7054_not
g60013 not n2554 ; n2554_not
g60014 not n2734 ; n2734_not
g60015 not n1609 ; n1609_not
g60016 not n2680 ; n2680_not
g60017 not n2671 ; n2671_not
g60018 not n7342 ; n7342_not
g60019 not n3094 ; n3094_not
g60020 not n9331 ; n9331_not
g60021 not n9430 ; n9430_not
g60022 not n2752 ; n2752_not
g60023 not n2545 ; n2545_not
g60024 not n1708 ; n1708_not
g60025 not n6451 ; n6451_not
g60026 not n2392 ; n2392_not
g60027 not n1573 ; n1573_not
g60028 not n6442 ; n6442_not
g60029 not n1582 ; n1582_not
g60030 not n1618 ; n1618_not
g60031 not n6460 ; n6460_not
g60032 not n3670 ; n3670_not
g60033 not n2743 ; n2743_not
g60034 not n7270 ; n7270_not
g60035 not n3058 ; n3058_not
g60036 not n3076 ; n3076_not
g60037 not n2158 ; n2158_not
g60038 not n2455 ; n2455_not
g60039 not n2563 ; n2563_not
g60040 not n2293 ; n2293_not
g60041 not n3067 ; n3067_not
g60042 not n7072 ; n7072_not
g60043 not n2437 ; n2437_not
g60044 not n3715 ; n3715_not
g60045 not n2086 ; n2086_not
g60046 not n7081 ; n7081_not
g60047 not n6433 ; n6433_not
g60048 not n2914 ; n2914_not
g60049 not n2095 ; n2095_not
g60050 not n3049 ; n3049_not
g60051 not n3085 ; n3085_not
g60052 not n9403 ; n9403_not
g60053 not n1726 ; n1726_not
g60054 not n2653 ; n2653_not
g60055 not n3454 ; n3454_not
g60056 not n1078 ; n1078_not
g60057 not n3175 ; n3175_not
g60058 not n1591 ; n1591_not
g60059 not n1069 ; n1069_not
g60060 not n2770 ; n2770_not
g60061 not n1744 ; n1744_not
g60062 not n7261 ; n7261_not
g60063 not n2536 ; n2536_not
g60064 not n2761 ; n2761_not
g60065 not n2527 ; n2527_not
g60066 not n2464 ; n2464_not
g60067 not n1159 ; n1159_not
g60068 not n7027 ; n7027_not
g60069 not n1717 ; n1717_not
g60070 not n2572 ; n2572_not
g60071 not n3139 ; n3139_not
g60072 not n2194 ; n2194_not
g60073 not n8054 ; n8054_not
g60074 not n2906 ; n2906_not
g60075 not n7181 ; n7181_not
g60076 not n4319 ; n4319_not
g60077 not n4346 ; n4346_not
g60078 not n2366 ; n2366_not
g60079 not n5093 ; n5093_not
g60080 not n4409 ; n4409_not
g60081 not n6371 ; n6371_not
g60082 not n4139 ; n4139_not
g60083 not n6902 ; n6902_not
g60084 not n9206 ; n9206_not
g60085 not n2762 ; n2762_not
g60086 not n8027 ; n8027_not
g60087 not n7415 ; n7415_not
g60088 not n1556 ; n1556_not
g60089 not n5345 ; n5345_not
g60090 not n5291 ; n5291_not
g60091 not n6380 ; n6380_not
g60092 not n2951 ; n2951_not
g60093 not n4391 ; n4391_not
g60094 not n2393 ; n2393_not
g60095 not n1574 ; n1574_not
g60096 not n6641 ; n6641_not
g60097 not n2087 ; n2087_not
g60098 not n7172 ; n7172_not
g60099 not n5318 ; n5318_not
g60100 not n2285 ; n2285_not
g60101 not n2564 ; n2564_not
g60102 not n6911 ; n6911_not
g60103 not n1628 ; n1628_not
g60104 not n2717 ; n2717_not
g60105 not n3059 ; n3059_not
g60106 not n9800 ; n9800_not
g60107 not n1763 ; n1763_not
g60108 not n7190 ; n7190_not
g60109 not n2573 ; n2573_not
g60110 not n5336 ; n5336_not
g60111 not n2384 ; n2384_not
g60112 not n2960 ; n2960_not
g60113 not n6632 ; n6632_not
g60114 not n4724 ; n4724_not
g60115 not n5084 ; n5084_not
g60116 not n7154 ; n7154_not
g60117 not n5309 ; n5309_not
g60118 not n2924 ; n2924_not
g60119 not n7910 ; n7910_not
g60120 not n1583 ; n1583_not
g60121 not n7505 ; n7505_not
g60122 not n2744 ; n2744_not
g60123 not n1745 ; n1745_not
g60124 not n6029 ; n6029_not
g60125 not n7406 ; n7406_not
g60126 not n4364 ; n4364_not
g60127 not n4418 ; n4418_not
g60128 not n1772 ; n1772_not
g60129 not n7208 ; n7208_not
g60130 not n2357 ; n2357_not
g60131 not n2735 ; n2735_not
g60132 not n5282 ; n5282_not
g60133 not n7325 ; n7325_not
g60134 not n6650 ; n6650_not
g60135 not n5327 ; n5327_not
g60136 not n6281 ; n6281_not
g60137 not n3716 ; n3716_not
g60138 not n5273 ; n5273_not
g60139 not n2933 ; n2933_not
g60140 not n5813 ; n5813_not
g60141 not n5264 ; n5264_not
g60142 not n6272 ; n6272_not
g60143 not n1592 ; n1592_not
g60144 not n7019 ; n7019_not
g60145 not n1790 ; n1790_not
g60146 not n2915 ; n2915_not
g60147 not n4373 ; n4373_not
g60148 not n2753 ; n2753_not
g60149 not n1844 ; n1844_not
g60150 not n2708 ; n2708_not
g60151 not n4607 ; n4607_not
g60152 not n4904 ; n4904_not
g60153 not n7091 ; n7091_not
g60154 not n1835 ; n1835_not
g60155 not n7253 ; n7253_not
g60156 not n4913 ; n4913_not
g60157 not n1826 ; n1826_not
g60158 not n9035 ; n9035_not
g60159 not n4616 ; n4616_not
g60160 not n7460 ; n7460_not
g60161 not n8342 ; n8342_not
g60162 not n4940 ; n4940_not
g60163 not n9125 ; n9125_not
g60164 not n2663 ; n2663_not
g60165 not n4931 ; n4931_not
g60166 not n4625 ; n4625_not
g60167 not n4382 ; n4382_not
g60168 not n8351 ; n8351_not
g60169 not n4922 ; n4922_not
g60170 not n1808 ; n1808_not
g60171 not n7550 ; n7550_not
g60172 not n1970 ; n1970_not
g60173 not n9431 ; n9431_not
g60174 not n4580 ; n4580_not
g60175 not n1880 ; n1880_not
g60176 not n9026 ; n9026_not
g60177 not n6317 ; n6317_not
g60178 not n5138 ; n5138_not
g60179 not n4733 ; n4733_not
g60180 not n2654 ; n2654_not
g60181 not n2636 ; n2636_not
g60182 not n1871 ; n1871_not
g60183 not n9134 ; n9134_not
g60184 not n2780 ; n2780_not
g60185 not n6605 ; n6605_not
g60186 not n1853 ; n1853_not
g60187 not n8531 ; n8531_not
g60188 not n2771 ; n2771_not
g60189 not n1862 ; n1862_not
g60190 not n6065 ; n6065_not
g60191 not n2645 ; n2645_not
g60192 not n7451 ; n7451_not
g60193 not n5129 ; n5129_not
g60194 not n4670 ; n4670_not
g60195 not n2690 ; n2690_not
g60196 not n7280 ; n7280_not
g60197 not n9116 ; n9116_not
g60198 not n4715 ; n4715_not
g60199 not n2096 ; n2096_not
g60200 not n7307 ; n7307_not
g60201 not n5048 ; n5048_not
g60202 not n1907 ; n1907_not
g60203 not n8063 ; n8063_not
g60204 not n4706 ; n4706_not
g60205 not n1943 ; n1943_not
g60206 not n2681 ; n2681_not
g60207 not n7064 ; n7064_not
g60208 not n8072 ; n8072_not
g60209 not n8513 ; n8513_not
g60210 not n7523 ; n7523_not
g60211 not n9602 ; n9602_not
g60212 not n7073 ; n7073_not
g60213 not n1916 ; n1916_not
g60214 not n9107 ; n9107_not
g60215 not n6254 ; n6254_not
g60216 not n9044 ; n9044_not
g60217 not n2159 ; n2159_not
g60218 not n7262 ; n7262_not
g60219 not n4643 ; n4643_not
g60220 not n7316 ; n7316_not
g60221 not n8360 ; n8360_not
g60222 not n7541 ; n7541_not
g60223 not n6074 ; n6074_not
g60224 not n4634 ; n4634_not
g60225 not n2078 ; n2078_not
g60226 not n5066 ; n5066_not
g60227 not n6092 ; n6092_not
g60228 not n4661 ; n4661_not
g60229 not n2177 ; n2177_not
g60230 not n6083 ; n6083_not
g60231 not n2069 ; n2069_not
g60232 not n4652 ; n4652_not
g60233 not n7271 ; n7271_not
g60234 not n2186 ; n2186_not
g60235 not n2843 ; n2843_not
g60236 not n5228 ; n5228_not
g60237 not n4454 ; n4454_not
g60238 not n7136 ; n7136_not
g60239 not n4760 ; n4760_not
g60240 not n7442 ; n7442_not
g60241 not n6353 ; n6353_not
g60242 not n4481 ; n4481_not
g60243 not n8405 ; n8405_not
g60244 not n2852 ; n2852_not
g60245 not n5822 ; n5822_not
g60246 not n9161 ; n9161_not
g60247 not n5219 ; n5219_not
g60248 not n2609 ; n2609_not
g60249 not n9152 ; n9152_not
g60250 not n6920 ; n6920_not
g60251 not n6047 ; n6047_not
g60252 not n7118 ; n7118_not
g60253 not n2267 ; n2267_not
g60254 not n7226 ; n7226_not
g60255 not n6812 ; n6812_not
g60256 not n4751 ; n4751_not
g60257 not n9008 ; n9008_not
g60258 not n6344 ; n6344_not
g60259 not n6803 ; n6803_not
g60260 not n4490 ; n4490_not
g60261 not n4436 ; n4436_not
g60262 not n6290 ; n6290_not
g60263 not n5255 ; n5255_not
g60264 not n5246 ; n5246_not
g60265 not n6038 ; n6038_not
g60266 not n2807 ; n2807_not
g60267 not n9170 ; n9170_not
g60268 not n2816 ; n2816_not
g60269 not n1781 ; n1781_not
g60270 not n6227 ; n6227_not
g60271 not n2582 ; n2582_not
g60272 not n5237 ; n5237_not
g60273 not n8900 ; n8900_not
g60274 not n2834 ; n2834_not
g60275 not n2276 ; n2276_not
g60276 not n4463 ; n4463_not
g60277 not n7424 ; n7424_not
g60278 not n2825 ; n2825_not
g60279 not n6362 ; n6362_not
g60280 not n7217 ; n7217_not
g60281 not n4544 ; n4544_not
g60282 not n2618 ; n2618_not
g60283 not n1952 ; n1952_not
g60284 not n4823 ; n4823_not
g60285 not n6326 ; n6326_not
g60286 not n8540 ; n8540_not
g60287 not n9017 ; n9017_not
g60288 not n4553 ; n4553_not
g60289 not n9143 ; n9143_not
g60290 not n4850 ; n4850_not
g60291 not n4571 ; n4571_not
g60292 not n4841 ; n4841_not
g60293 not n8009 ; n8009_not
g60294 not n4832 ; n4832_not
g60295 not n4562 ; n4562_not
g60296 not n7244 ; n7244_not
g60297 not n8504 ; n8504_not
g60298 not n5156 ; n5156_not
g60299 not n5183 ; n5183_not
g60300 not n7235 ; n7235_not
g60301 not n7109 ; n7109_not
g60302 not n6335 ; n6335_not
g60303 not n6821 ; n6821_not
g60304 not n4517 ; n4517_not
g60305 not n5192 ; n5192_not
g60306 not n6236 ; n6236_not
g60307 not n5147 ; n5147_not
g60308 not n2258 ; n2258_not
g60309 not n4508 ; n4508_not
g60310 not n4427 ; n4427_not
g60311 not n9521 ; n9521_not
g60312 not n6056 ; n6056_not
g60313 not n4535 ; n4535_not
g60314 not n5174 ; n5174_not
g60315 not n6830 ; n6830_not
g60316 not n9053 ; n9053_not
g60317 not n4526 ; n4526_not
g60318 not n3626 ; n3626_not
g60319 not n6416 ; n6416_not
g60320 not n7361 ; n7361_not
g60321 not n7046 ; n7046_not
g60322 not n3914 ; n3914_not
g60323 not n3329 ; n3329_not
g60324 not n3635 ; n3635_not
g60325 not n3608 ; n3608_not
g60326 not n8711 ; n8711_not
g60327 not n2465 ; n2465_not
g60328 not n5633 ; n5633_not
g60329 not n6515 ; n6515_not
g60330 not n5552 ; n5552_not
g60331 not n3923 ; n3923_not
g60332 not n3941 ; n3941_not
g60333 not n3590 ; n3590_not
g60334 not n5921 ; n5921_not
g60335 not n3752 ; n3752_not
g60336 not n6506 ; n6506_not
g60337 not n3653 ; n3653_not
g60338 not n9314 ; n9314_not
g60339 not n3932 ; n3932_not
g60340 not n6407 ; n6407_not
g60341 not n5624 ; n5624_not
g60342 not n5804 ; n5804_not
g60343 not n9260 ; n9260_not
g60344 not n3644 ; n3644_not
g60345 not n1097 ; n1097_not
g60346 not n8720 ; n8720_not
g60347 not n7352 ; n7352_not
g60348 not n1088 ; n1088_not
g60349 not n3356 ; n3356_not
g60350 not n2249 ; n2249_not
g60351 not n5903 ; n5903_not
g60352 not n6425 ; n6425_not
g60353 not n6533 ; n6533_not
g60354 not n5660 ; n5660_not
g60355 not n6191 ; n6191_not
g60356 not n3617 ; n3617_not
g60357 not n3338 ; n3338_not
g60358 not n3464 ; n3464_not
g60359 not n3905 ; n3905_not
g60360 not n5642 ; n5642_not
g60361 not n6137 ; n6137_not
g60362 not n6524 ; n6524_not
g60363 not n3347 ; n3347_not
g60364 not n3455 ; n3455_not
g60365 not n9440 ; n9440_not
g60366 not n5651 ; n5651_not
g60367 not n3284 ; n3284_not
g60368 not n3563 ; n3563_not
g60369 not n9512 ; n9512_not
g60370 not n3707 ; n3707_not
g60371 not n2483 ; n2483_not
g60372 not n9611 ; n9611_not
g60373 not n3275 ; n3275_not
g60374 not n3554 ; n3554_not
g60375 not n7343 ; n7343_not
g60376 not n9080 ; n9080_not
g60377 not n3518 ; n3518_not
g60378 not n5561 ; n5561_not
g60379 not n3257 ; n3257_not
g60380 not n6470 ; n6470_not
g60381 not n3509 ; n3509_not
g60382 not n1259 ; n1259_not
g60383 not n8423 ; n8423_not
g60384 not n3248 ; n3248_not
g60385 not n9242 ; n9242_not
g60386 not n2339 ; n2339_not
g60387 not n5570 ; n5570_not
g60388 not n3266 ; n3266_not
g60389 not n6704 ; n6704_not
g60390 not n9251 ; n9251_not
g60391 not n2474 ; n2474_not
g60392 not n3581 ; n3581_not
g60393 not n3671 ; n3671_not
g60394 not n8414 ; n8414_not
g60395 not n8702 ; n8702_not
g60396 not n3950 ; n3950_not
g60397 not n5606 ; n5606_not
g60398 not n3743 ; n3743_not
g60399 not n7370 ; n7370_not
g60400 not n3662 ; n3662_not
g60401 not n5615 ; n5615_not
g60402 not n2348 ; n2348_not
g60403 not n1286 ; n1286_not
g60404 not n3491 ; n3491_not
g60405 not n9701 ; n9701_not
g60406 not n1268 ; n1268_not
g60407 not n5507 ; n5507_not
g60408 not n3734 ; n3734_not
g60409 not n3572 ; n3572_not
g60410 not n3293 ; n3293_not
g60411 not n3680 ; n3680_not
g60412 not n5930 ; n5930_not
g60413 not n8801 ; n8801_not
g60414 not n6155 ; n6155_not
g60415 not n9503 ; n9503_not
g60416 not n5408 ; n5408_not
g60417 not n5417 ; n5417_not
g60418 not n5750 ; n5750_not
g60419 not n6182 ; n6182_not
g60420 not n3419 ; n3419_not
g60421 not n5741 ; n5741_not
g60422 not n6461 ; n6461_not
g60423 not n7082 ; n7082_not
g60424 not n5732 ; n5732_not
g60425 not n8810 ; n8810_not
g60426 not n9350 ; n9350_not
g60427 not n3806 ; n3806_not
g60428 not n8441 ; n8441_not
g60429 not n9620 ; n9620_not
g60430 not n5831 ; n5831_not
g60431 not n6614 ; n6614_not
g60432 not n8450 ; n8450_not
g60433 not n2429 ; n2429_not
g60434 not n7334 ; n7334_not
g60435 not n6173 ; n6173_not
g60436 not n9530 ; n9530_not
g60437 not n3761 ; n3761_not
g60438 not n9413 ; n9413_not
g60439 not n9710 ; n9710_not
g60440 not n6434 ; n6434_not
g60441 not n3860 ; n3860_not
g60442 not n6560 ; n6560_not
g60443 not n3374 ; n3374_not
g60444 not n3851 ; n3851_not
g60445 not n9323 ; n9323_not
g60446 not n6542 ; n6542_not
g60447 not n3365 ; n3365_not
g60448 not n5462 ; n5462_not
g60449 not n3446 ; n3446_not
g60450 not n6551 ; n6551_not
g60451 not n7028 ; n7028_not
g60452 not n5453 ; n5453_not
g60453 not n8018 ; n8018_not
g60454 not n3833 ; n3833_not
g60455 not n5714 ; n5714_not
g60456 not n3392 ; n3392_not
g60457 not n7514 ; n7514_not
g60458 not n6452 ; n6452_not
g60459 not n5723 ; n5723_not
g60460 not n6146 ; n6146_not
g60461 not n9341 ; n9341_not
g60462 not n3545 ; n3545_not
g60463 not n7037 ; n7037_not
g60464 not n3842 ; n3842_not
g60465 not n5444 ; n5444_not
g60466 not n5705 ; n5705_not
g60467 not n3383 ; n3383_not
g60468 not n2447 ; n2447_not
g60469 not n6443 ; n6443_not
g60470 not n4094 ; n4094_not
g60471 not n1547 ; n1547_not
g60472 not n7127 ; n7127_not
g60473 not n4805 ; n4805_not
g60474 not n9062 ; n9062_not
g60475 not n1565 ; n1565_not
g60476 not n2528 ; n2528_not
g60477 not n4229 ; n4229_not
g60478 not n1529 ; n1529_not
g60479 not n3185 ; n3185_not
g60480 not n8603 ; n8603_not
g60481 not n1538 ; n1538_not
g60482 not n5354 ; n5354_not
g60483 not n5426 ; n5426_not
g60484 not n4238 ; n4238_not
g60485 not n4184 ; n4184_not
g60486 not n6722 ; n6722_not
g60487 not n5471 ; n5471_not
g60488 not n1358 ; n1358_not
g60489 not n4175 ; n4175_not
g60490 not n3176 ; n3176_not
g60491 not n1349 ; n1349_not
g60492 not n4166 ; n4166_not
g60493 not n8621 ; n8621_not
g60494 not n2519 ; n2519_not
g60495 not n1394 ; n1394_not
g60496 not n8612 ; n8612_not
g60497 not n4193 ; n4193_not
g60498 not n9224 ; n9224_not
g60499 not n1367 ; n1367_not
g60500 not n5372 ; n5372_not
g60501 not n4283 ; n4283_not
g60502 not n2195 ; n2195_not
g60503 not n3095 ; n3095_not
g60504 not n2555 ; n2555_not
g60505 not n4049 ; n4049_not
g60506 not n4292 ; n4292_not
g60507 not n3068 ; n3068_not
g60508 not n2294 ; n2294_not
g60509 not n8045 ; n8045_not
g60510 not n3077 ; n3077_not
g60511 not n6119 ; n6119_not
g60512 not n3086 ; n3086_not
g60513 not n5057 ; n5057_not
g60514 not n5363 ; n5363_not
g60515 not n5381 ; n5381_not
g60516 not n1484 ; n1484_not
g60517 not n2537 ; n2537_not
g60518 not n4256 ; n4256_not
g60519 not n3158 ; n3158_not
g60520 not n1493 ; n1493_not
g60521 not n3167 ; n3167_not
g60522 not n4247 ; n4247_not
g60523 not n1619 ; n1619_not
g60524 not n4274 ; n4274_not
g60525 not n9215 ; n9215_not
g60526 not n1475 ; n1475_not
g60527 not n4058 ; n4058_not
g60528 not n2546 ; n2546_not
g60529 not n4265 ; n4265_not
g60530 not n4067 ; n4067_not
g60531 not n4076 ; n4076_not
g60532 not n9071 ; n9071_not
g60533 not n9404 ; n9404_not
g60534 not n5912 ; n5912_not
g60535 not n2438 ; n2438_not
g60536 not n9233 ; n9233_not
g60537 not n5534 ; n5534_not
g60538 not n2492 ; n2492_not
g60539 not n3473 ; n3473_not
g60540 not n6128 ; n6128_not
g60541 not n6209 ; n6209_not
g60542 not n4148 ; n4148_not
g60543 not n1448 ; n1448_not
g60544 not n8630 ; n8630_not
g60545 not n1439 ; n1439_not
g60546 not n4157 ; n4157_not
g60547 not n5516 ; n5516_not
g60548 not n3428 ; n3428_not
g60549 not n6245 ; n6245_not
g60550 not n8262 ; n8262_not
g60551 not n2295 ; n2295_not
g60552 not n9090 ; n9090_not
g60553 not n2286 ; n2286_not
g60554 not n2088 ; n2088_not
g60555 not n8271 ; n8271_not
g60556 not n2097 ; n2097_not
g60557 not n8406 ; n8406_not
g60558 not n6138 ; n6138_not
g60559 not n6156 ; n6156_not
g60560 not n2196 ; n2196_not
g60561 not n8190 ; n8190_not
g60562 not n8415 ; n8415_not
g60563 not n5823 ; n5823_not
g60564 not n6129 ; n6129_not
g60565 not n5814 ; n5814_not
g60566 not n8226 ; n8226_not
g60567 not n2349 ; n2349_not
g60568 not n8253 ; n8253_not
g60569 not n2079 ; n2079_not
g60570 not n2376 ; n2376_not
g60571 not n8217 ; n8217_not
g60572 not n2358 ; n2358_not
g60573 not n2394 ; n2394_not
g60574 not n2187 ; n2187_not
g60575 not n8208 ; n8208_not
g60576 not n8244 ; n8244_not
g60577 not n8280 ; n8280_not
g60578 not n2169 ; n2169_not
g60579 not n4734 ; n4734_not
g60580 not n4725 ; n4725_not
g60581 not n2385 ; n2385_not
g60582 not n9081 ; n9081_not
g60583 not n7056 ; n7056_not
g60584 not n4761 ; n4761_not
g60585 not n9414 ; n9414_not
g60586 not n4716 ; n4716_not
g60587 not n8433 ; n8433_not
g60588 not n6147 ; n6147_not
g60589 not n8235 ; n8235_not
g60590 not n6093 ; n6093_not
g60591 not n1386 ; n1386_not
g60592 not n1368 ; n1368_not
g60593 not n1359 ; n1359_not
g60594 not n8073 ; n8073_not
g60595 not n6822 ; n6822_not
g60596 not n5562 ; n5562_not
g60597 not n5940 ; n5940_not
g60598 not n9243 ; n9243_not
g60599 not n5571 ; n5571_not
g60600 not n1269 ; n1269_not
g60601 not n5922 ; n5922_not
g60602 not n5517 ; n5517_not
g60603 not n5580 ; n5580_not
g60604 not n8082 ; n8082_not
g60605 not n1296 ; n1296_not
g60606 not n5508 ; n5508_not
g60607 not n5931 ; n5931_not
g60608 not n1278 ; n1278_not
g60609 not n1179 ; n1179_not
g60610 not n1188 ; n1188_not
g60611 not n6831 ; n6831_not
g60612 not n1197 ; n1197_not
g60613 not n9252 ; n9252_not
g60614 not n5607 ; n5607_not
g60615 not n1089 ; n1089_not
g60616 not n5913 ; n5913_not
g60617 not n9441 ; n9441_not
g60618 not n8028 ; n8028_not
g60619 not n5616 ; n5616_not
g60620 not n5418 ; n5418_not
g60621 not n1593 ; n1593_not
g60622 not n1584 ; n1584_not
g60623 not n1557 ; n1557_not
g60624 not n5436 ; n5436_not
g60625 not n1566 ; n1566_not
g60626 not n6804 ; n6804_not
g60627 not n1548 ; n1548_not
g60628 not n1395 ; n1395_not
g60629 not n1539 ; n1539_not
g60630 not n5454 ; n5454_not
g60631 not n5463 ; n5463_not
g60632 not n9225 ; n9225_not
g60633 not n5481 ; n5481_not
g60634 not n1494 ; n1494_not
g60635 not n6813 ; n6813_not
g60636 not n1485 ; n1485_not
g60637 not n7119 ; n7119_not
g60638 not n5526 ; n5526_not
g60639 not n5535 ; n5535_not
g60640 not n5904 ; n5904_not
g60641 not n9234 ; n9234_not
g60642 not n7083 ; n7083_not
g60643 not n8172 ; n8172_not
g60644 not n5724 ; n5724_not
g60645 not n7038 ; n7038_not
g60646 not n5733 ; n5733_not
g60647 not n9351 ; n9351_not
g60648 not n7074 ; n7074_not
g60649 not n5427 ; n5427_not
g60650 not n5742 ; n5742_not
g60651 not n8118 ; n8118_not
g60652 not n9360 ; n9360_not
g60653 not n6903 ; n6903_not
g60654 not n5751 ; n5751_not
g60655 not n7047 ; n7047_not
g60656 not n8163 ; n8163_not
g60657 not n5760 ; n5760_not
g60658 not n6912 ; n6912_not
g60659 not n5409 ; n5409_not
g60660 not n8127 ; n8127_not
g60661 not n6921 ; n6921_not
g60662 not n5841 ; n5841_not
g60663 not n8154 ; n8154_not
g60664 not n9405 ; n9405_not
g60665 not n6930 ; n6930_not
g60666 not n8145 ; n8145_not
g60667 not n9423 ; n9423_not
g60668 not n8136 ; n8136_not
g60669 not n5625 ; n5625_not
g60670 not n9261 ; n9261_not
g60671 not n5634 ; n5634_not
g60672 not n8091 ; n8091_not
g60673 not n6840 ; n6840_not
g60674 not n5643 ; n5643_not
g60675 not n8019 ; n8019_not
g60676 not n1098 ; n1098_not
g60677 not n5652 ; n5652_not
g60678 not n9270 ; n9270_not
g60679 not n5472 ; n5472_not
g60680 not n5661 ; n5661_not
g60681 not n5670 ; n5670_not
g60682 not n7029 ; n7029_not
g60683 not n9306 ; n9306_not
g60684 not n8181 ; n8181_not
g60685 not n7092 ; n7092_not
g60686 not n5706 ; n5706_not
g60687 not n8109 ; n8109_not
g60688 not n9333 ; n9333_not
g60689 not n5715 ; n5715_not
g60690 not n8334 ; n8334_not
g60691 not n1863 ; n1863_not
g60692 not n9135 ; n9135_not
g60693 not n5139 ; n5139_not
g60694 not n1872 ; n1872_not
g60695 not n1881 ; n1881_not
g60696 not n5148 ; n5148_not
g60697 not n1962 ; n1962_not
g60698 not n8325 ; n8325_not
g60699 not n1890 ; n1890_not
g60700 not n4815 ; n4815_not
g60701 not n9144 ; n9144_not
g60702 not n5166 ; n5166_not
g60703 not n1908 ; n1908_not
g60704 not n6057 ; n6057_not
g60705 not n1917 ; n1917_not
g60706 not n1944 ; n1944_not
g60707 not n5157 ; n5157_not
g60708 not n7443 ; n7443_not
g60709 not n1746 ; n1746_not
g60710 not n8316 ; n8316_not
g60711 not n8910 ; n8910_not
g60712 not n6048 ; n6048_not
g60713 not n9153 ; n9153_not
g60714 not n5832 ; n5832_not
g60715 not n8307 ; n8307_not
g60716 not n1953 ; n1953_not
g60717 not n9108 ; n9108_not
g60718 not n7470 ; n7470_not
g60719 not n5049 ; n5049_not
g60720 not n5058 ; n5058_not
g60721 not n9117 ; n9117_not
g60722 not n6084 ; n6084_not
g60723 not n7461 ; n7461_not
g60724 not n1980 ; n1980_not
g60725 not n8370 ; n8370_not
g60726 not n5076 ; n5076_not
g60727 not n8361 ; n8361_not
g60728 not n6075 ; n6075_not
g60729 not n5094 ; n5094_not
g60730 not n9126 ; n9126_not
g60731 not n8352 ; n8352_not
g60732 not n1818 ; n1818_not
g60733 not n1827 ; n1827_not
g60734 not n1836 ; n1836_not
g60735 not n1845 ; n1845_not
g60736 not n6066 ; n6066_not
g60737 not n8343 ; n8343_not
g60738 not n1854 ; n1854_not
g60739 not n1719 ; n1719_not
g60740 not n1692 ; n1692_not
g60741 not n8037 ; n8037_not
g60742 not n1683 ; n1683_not
g60743 not n7137 ; n7137_not
g60744 not n9207 ; n9207_not
g60745 not n5067 ; n5067_not
g60746 not n1674 ; n1674_not
g60747 not n1665 ; n1665_not
g60748 not n9450 ; n9450_not
g60749 not n1656 ; n1656_not
g60750 not n8046 ; n8046_not
g60751 not n1647 ; n1647_not
g60752 not n7128 ; n7128_not
g60753 not n1638 ; n1638_not
g60754 not n9216 ; n9216_not
g60755 not n1476 ; n1476_not
g60756 not n1773 ; n1773_not
g60757 not n9162 ; n9162_not
g60758 not n1782 ; n1782_not
g60759 not n7146 ; n7146_not
g60760 not n1791 ; n1791_not
g60761 not n8901 ; n8901_not
g60762 not n6039 ; n6039_not
g60763 not n9171 ; n9171_not
g60764 not n7164 ; n7164_not
g60765 not n9180 ; n9180_not
g60766 not n1755 ; n1755_not
g60767 not n7920 ; n7920_not
g60768 not n1728 ; n1728_not
g60769 not n2961 ; n2961_not
g60770 not n2916 ; n2916_not
g60771 not n7641 ; n7641_not
g60772 not n3069 ; n3069_not
g60773 not n3078 ; n3078_not
g60774 not n7650 ; n7650_not
g60775 not n3087 ; n3087_not
g60776 not n4293 ; n4293_not
g60777 not n3096 ; n3096_not
g60778 not n6642 ; n6642_not
g60779 not n4383 ; n4383_not
g60780 not n7605 ; n7605_not
g60781 not n7614 ; n7614_not
g60782 not n4374 ; n4374_not
g60783 not n6651 ; n6651_not
g60784 not n6660 ; n6660_not
g60785 not n7623 ; n7623_not
g60786 not n4356 ; n4356_not
g60787 not n2934 ; n2934_not
g60788 not n2925 ; n2925_not
g60789 not n7632 ; n7632_not
g60790 not n4347 ; n4347_not
g60791 not n4338 ; n4338_not
g60792 not n4248 ; n4248_not
g60793 not n4077 ; n4077_not
g60794 not n3177 ; n3177_not
g60795 not n8604 ; n8604_not
g60796 not n3195 ; n3195_not
g60797 not n4239 ; n4239_not
g60798 not n6705 ; n6705_not
g60799 not n3249 ; n3249_not
g60800 not n3258 ; n3258_not
g60801 not n7704 ; n7704_not
g60802 not n3267 ; n3267_not
g60803 not n3276 ; n3276_not
g60804 not n8460 ; n8460_not
g60805 not n3285 ; n3285_not
g60806 not n7713 ; n7713_not
g60807 not n3294 ; n3294_not
g60808 not n4194 ; n4194_not
g60809 not n7560 ; n7560_not
g60810 not n4284 ; n4284_not
g60811 not n2880 ; n2880_not
g60812 not n4275 ; n4275_not
g60813 not n4059 ; n4059_not
g60814 not n4266 ; n4266_not
g60815 not n2871 ; n2871_not
g60816 not n4257 ; n4257_not
g60817 not n4068 ; n4068_not
g60818 not n7551 ; n7551_not
g60819 not n3168 ; n3168_not
g60820 not n9027 ; n9027_not
g60821 not n4581 ; n4581_not
g60822 not n2709 ; n2709_not
g60823 not n2646 ; n2646_not
g60824 not n4572 ; n4572_not
g60825 not n9018 ; n9018_not
g60826 not n4563 ; n4563_not
g60827 not n4554 ; n4554_not
g60828 not n4419 ; n4419_not
g60829 not n6606 ; n6606_not
g60830 not n4545 ; n4545_not
g60831 not n4536 ; n4536_not
g60832 not n4428 ; n4428_not
g60833 not n6282 ; n6282_not
g60834 not n4626 ; n4626_not
g60835 not n6291 ; n6291_not
g60836 not n4617 ; n4617_not
g60837 not n7902 ; n7902_not
g60838 not n4608 ; n4608_not
g60839 not n4392 ; n4392_not
g60840 not n8514 ; n8514_not
g60841 not n2664 ; n2664_not
g60842 not n8532 ; n8532_not
g60843 not n6309 ; n6309_not
g60844 not n2655 ; n2655_not
g60845 not n4590 ; n4590_not
g60846 not n4464 ; n4464_not
g60847 not n4446 ; n4446_not
g60848 not n2943 ; n2943_not
g60849 not n2727 ; n2727_not
g60850 not n2718 ; n2718_not
g60851 not n2970 ; n2970_not
g60852 not n4527 ; n4527_not
g60853 not n4437 ; n4437_not
g60854 not n4518 ; n4518_not
g60855 not n2619 ; n2619_not
g60856 not n6615 ; n6615_not
g60857 not n8541 ; n8541_not
g60858 not n4509 ; n4509_not
g60859 not n2862 ; n2862_not
g60860 not n9009 ; n9009_not
g60861 not n4491 ; n4491_not
g60862 not n8550 ; n8550_not
g60863 not n3807 ; n3807_not
g60864 not n3564 ; n3564_not
g60865 not n3546 ; n3546_not
g60866 not n3825 ; n3825_not
g60867 not n3555 ; n3555_not
g60868 not n3816 ; n3816_not
g60869 not n3429 ; n3429_not
g60870 not n7506 ; n7506_not
g60871 not n3573 ; n3573_not
g60872 not n3474 ; n3474_not
g60873 not n3762 ; n3762_not
g60874 not n3645 ; n3645_not
g60875 not n8712 ; n8712_not
g60876 not n3465 ; n3465_not
g60877 not n3636 ; n3636_not
g60878 not n3627 ; n3627_not
g60879 not n3456 ; n3456_not
g60880 not n3618 ; n3618_not
g60881 not n8721 ; n8721_not
g60882 not n3609 ; n3609_not
g60883 not n7812 ; n7812_not
g60884 not n8730 ; n8730_not
g60885 not n6192 ; n6192_not
g60886 not n3591 ; n3591_not
g60887 not n7803 ; n7803_not
g60888 not n3582 ; n3582_not
g60889 not n3690 ; n3690_not
g60890 not n6624 ; n6624_not
g60891 not n3753 ; n3753_not
g60892 not n3654 ; n3654_not
g60893 not n3681 ; n3681_not
g60894 not n3663 ; n3663_not
g60895 not n3744 ; n3744_not
g60896 not n3672 ; n3672_not
g60897 not n9504 ; n9504_not
g60898 not n3708 ; n3708_not
g60899 not n8802 ; n8802_not
g60900 not n3717 ; n3717_not
g60901 not n3771 ; n3771_not
g60902 not n3726 ; n3726_not
g60903 not n6732 ; n6732_not
g60904 not n3375 ; n3375_not
g60905 not n6723 ; n6723_not
g60906 not n3384 ; n3384_not
g60907 not n3393 ; n3393_not
g60908 not n8451 ; n8451_not
g60909 not n8631 ; n8631_not
g60910 not n8640 ; n8640_not
g60911 not n3366 ; n3366_not
g60912 not n3438 ; n3438_not
g60913 not n3357 ; n3357_not
g60914 not n4086 ; n4086_not
g60915 not n3348 ; n3348_not
g60916 not n3339 ; n3339_not
g60917 not n8613 ; n8613_not
g60918 not n6255 ; n6255_not
g60919 not n4185 ; n4185_not
g60920 not n3186 ; n3186_not
g60921 not n4176 ; n4176_not
g60922 not n4167 ; n4167_not
g60923 not n8622 ; n8622_not
g60924 not n4158 ; n4158_not
g60925 not n6246 ; n6246_not
g60926 not n4149 ; n4149_not
g60927 not n7722 ; n7722_not
g60928 not n8424 ; n8424_not
g60929 not n7821 ; n7821_not
g60930 not n9513 ; n9513_not
g60931 not n7524 ; n7524_not
g60932 not n7731 ; n7731_not
g60933 not n7515 ; n7515_not
g60934 not n8703 ; n8703_not
g60935 not n7740 ; n7740_not
g60936 not n6237 ; n6237_not
g60937 not n7830 ; n7830_not
g60938 not n6714 ; n6714_not
g60939 not n3483 ; n3483_not
g60940 not n3519 ; n3519_not
g60941 not n3528 ; n3528_not
g60942 not n3537 ; n3537_not
g60943 not n2466 ; n2466_not
g60944 not n8523 ; n8523_not
g60945 not n8505 ; n8505_not
g60946 not n2268 ; n2268_not
g60947 not n2448 ; n2448_not
g60948 not n2475 ; n2475_not
g60949 not n2691 ; n2691_not
g60950 not n2277 ; n2277_not
g60951 not n9045 ; n9045_not
g60952 not n2439 ; n2439_not
g60953 not n2484 ; n2484_not
g60954 not n9072 ; n9072_not
g60955 not n4806 ; n4806_not
g60956 not n4680 ; n4680_not
g60957 not n2259 ; n2259_not
g60958 not n4662 ; n4662_not
g60959 not n2457 ; n2457_not
g60960 not n7533 ; n7533_not
g60961 not n4671 ; n4671_not
g60962 not n6264 ; n6264_not
g60963 not n2565 ; n2565_not
g60964 not n2574 ; n2574_not
g60965 not n9324 ; n9324_not
g60966 not n4770 ; n4770_not
g60967 not n2628 ; n2628_not
g60968 not n2583 ; n2583_not
g60969 not n4743 ; n4743_not
g60970 not n9054 ; n9054_not
g60971 not n2493 ; n2493_not
g60972 not n9063 ; n9063_not
g60973 not n2529 ; n2529_not
g60974 not n2538 ; n2538_not
g60975 not n2547 ; n2547_not
g60976 not n2673 ; n2673_not
g60977 not n2556 ; n2556_not
g60978 not n6219 ; n6219_not
g60979 not n6174 ; n6174_not
g60980 not n4653 ; n4653_not
g60981 not n9036 ; n9036_not
g60982 not n6183 ; n6183_not
g60983 not n4635 ; n4635_not
g60984 not n4644 ; n4644_not
g60985 not n8209 ; n8209_not
g60986 not n6940 ; n6940_not
g60987 not n5527 ; n5527_not
g60988 not n6472 ; n6472_not
g60989 not n9235 ; n9235_not
g60990 not n5545 ; n5545_not
g60991 not n3493 ; n3493_not
g60992 not n5554 ; n5554_not
g60993 not n8029 ; n8029_not
g60994 not n8434 ; n8434_not
g60995 not n6706 ; n6706_not
g60996 not n6832 ; n6832_not
g60997 not n9064 ; n9064_not
g60998 not n5536 ; n5536_not
g60999 not n3529 ; n3529_not
g61000 not n5833 ; n5833_not
g61001 not n8047 ; n8047_not
g61002 not n8191 ; n8191_not
g61003 not n2296 ; n2296_not
g61004 not n7480 ; n7480_not
g61005 not n6463 ; n6463_not
g61006 not n8650 ; n8650_not
g61007 not n5167 ; n5167_not
g61008 not n1387 ; n1387_not
g61009 not n9640 ; n9640_not
g61010 not n8416 ; n8416_not
g61011 not n6184 ; n6184_not
g61012 not n7345 ; n7345_not
g61013 not n8353 ; n8353_not
g61014 not n7831 ; n7831_not
g61015 not n3466 ; n3466_not
g61016 not n3475 ; n3475_not
g61017 not n4483 ; n4483_not
g61018 not n5707 ; n5707_not
g61019 not n9415 ; n9415_not
g61020 not n4951 ; n4951_not
g61021 not n8083 ; n8083_not
g61022 not n3727 ; n3727_not
g61023 not n4942 ; n4942_not
g61024 not n6490 ; n6490_not
g61025 not n5509 ; n5509_not
g61026 not n1288 ; n1288_not
g61027 not n7822 ; n7822_not
g61028 not n8218 ; n8218_not
g61029 not n9406 ; n9406_not
g61030 not n5590 ; n5590_not
g61031 not n5932 ; n5932_not
g61032 not n7471 ; n7471_not
g61033 not n4825 ; n4825_not
g61034 not n8236 ; n8236_not
g61035 not n4735 ; n4735_not
g61036 not n3970 ; n3970_not
g61037 not n3763 ; n3763_not
g61038 not n8245 ; n8245_not
g61039 not n9073 ; n9073_not
g61040 not n8146 ; n8146_not
g61041 not n8227 ; n8227_not
g61042 not n2287 ; n2287_not
g61043 not n5941 ; n5941_not
g61044 not n3538 ; n3538_not
g61045 not n5518 ; n5518_not
g61046 not n7057 ; n7057_not
g61047 not n1198 ; n1198_not
g61048 not n9082 ; n9082_not
g61049 not n6481 ; n6481_not
g61050 not n8425 ; n8425_not
g61051 not n5572 ; n5572_not
g61052 not n9244 ; n9244_not
g61053 not n3718 ; n3718_not
g61054 not n1189 ; n1189_not
g61055 not n1279 ; n1279_not
g61056 not n9370 ; n9370_not
g61057 not n9514 ; n9514_not
g61058 not n7723 ; n7723_not
g61059 not n7237 ; n7237_not
g61060 not n5581 ; n5581_not
g61061 not n5725 ; n5725_not
g61062 not n6751 ; n6751_not
g61063 not n3196 ; n3196_not
g61064 not n4564 ; n4564_not
g61065 not n8614 ; n8614_not
g61066 not n9433 ; n9433_not
g61067 not n6229 ; n6229_not
g61068 not n2269 ; n2269_not
g61069 not n5743 ; n5743_not
g61070 not n5464 ; n5464_not
g61071 not n3187 ; n3187_not
g61072 not n5824 ; n5824_not
g61073 not n6931 ; n6931_not
g61074 not n6436 ; n6436_not
g61075 not n8164 ; n8164_not
g61076 not n5473 ; n5473_not
g61077 not n2278 ; n2278_not
g61078 not n4555 ; n4555_not
g61079 not n9226 ; n9226_not
g61080 not n3178 ; n3178_not
g61081 not n3736 ; n3736_not
g61082 not n4546 ; n4546_not
g61083 not n8623 ; n8623_not
g61084 not n9361 ; n9361_not
g61085 not n4087 ; n4087_not
g61086 not n8911 ; n8911_not
g61087 not n6814 ; n6814_not
g61088 not n1558 ; n1558_not
g61089 not n9055 ; n9055_not
g61090 not n4582 ; n4582_not
g61091 not n2593 ; n2593_not
g61092 not n6427 ; n6427_not
g61093 not n7705 ; n7705_not
g61094 not n5446 ; n5446_not
g61095 not n4753 ; n4753_not
g61096 not n8155 ; n8155_not
g61097 not n6715 ; n6715_not
g61098 not n7219 ; n7219_not
g61099 not n2377 ; n2377_not
g61100 not n4573 ; n4573_not
g61101 not n7534 ; n7534_not
g61102 not n8461 ; n8461_not
g61103 not n5734 ; n5734_not
g61104 not n9622 ; n9622_not
g61105 not n8344 ; n8344_not
g61106 not n7714 ; n7714_not
g61107 not n5716 ; n5716_not
g61108 not n9613 ; n9613_not
g61109 not n5806 ; n5806_not
g61110 not n8335 ; n8335_not
g61111 not n8632 ; n8632_not
g61112 not n9424 ; n9424_not
g61113 not n7228 ; n7228_not
g61114 not n8182 ; n8182_not
g61115 not n5761 ; n5761_not
g61116 not n7048 ; n7048_not
g61117 not n6454 ; n6454_not
g61118 not n9820 ; n9820_not
g61119 not n4096 ; n4096_not
g61120 not n8641 ; n8641_not
g61121 not n4960 ; n4960_not
g61122 not n4771 ; n4771_not
g61123 not n3754 ; n3754_not
g61124 not n4726 ; n4726_not
g61125 not n5770 ; n5770_not
g61126 not n3448 ; n3448_not
g61127 not n4078 ; n4078_not
g61128 not n4069 ; n4069_not
g61129 not n6166 ; n6166_not
g61130 not n9091 ; n9091_not
g61131 not n7354 ; n7354_not
g61132 not n6247 ; n6247_not
g61133 not n4537 ; n4537_not
g61134 not n6823 ; n6823_not
g61135 not n6742 ; n6742_not
g61136 not n9802 ; n9802_not
g61137 not n5491 ; n5491_not
g61138 not n9730 ; n9730_not
g61139 not n4780 ; n4780_not
g61140 not n6445 ; n6445_not
g61141 not n2197 ; n2197_not
g61142 not n4528 ; n4528_not
g61143 not n8137 ; n8137_not
g61144 not n5752 ; n5752_not
g61145 not n7525 ; n7525_not
g61146 not n1468 ; n1468_not
g61147 not n2395 ; n2395_not
g61148 not n8173 ; n8173_not
g61149 not n4519 ; n4519_not
g61150 not n8443 ; n8443_not
g61151 not n1459 ; n1459_not
g61152 not n8326 ; n8326_not
g61153 not n6580 ; n6580_not
g61154 not n7282 ; n7282_not
g61155 not n3844 ; n3844_not
g61156 not n3781 ; n3781_not
g61157 not n8821 ; n8821_not
g61158 not n3709 ; n3709_not
g61159 not n6607 ; n6607_not
g61160 not n5635 ; n5635_not
g61161 not n5680 ; n5680_not
g61162 not n3439 ; n3439_not
g61163 not n9901 ; n9901_not
g61164 not n3835 ; n3835_not
g61165 not n3817 ; n3817_not
g61166 not n8308 ; n8308_not
g61167 not n4915 ; n4915_not
g61168 not n7084 ; n7084_not
g61169 not n3808 ; n3808_not
g61170 not n8740 ; n8740_not
g61171 not n9307 ; n9307_not
g61172 not n7273 ; n7273_not
g61173 not n7804 ; n7804_not
g61174 not n8290 ; n8290_not
g61175 not n9703 ; n9703_not
g61176 not n9316 ; n9316_not
g61177 not n5617 ; n5617_not
g61178 not n3862 ; n3862_not
g61179 not n6562 ; n6562_not
g61180 not n7381 ; n7381_not
g61181 not n3853 ; n3853_not
g61182 not n6652 ; n6652_not
g61183 not n5626 ; n5626_not
g61184 not n8380 ; n8380_not
g61185 not n2449 ; n2449_not
g61186 not n7327 ; n7327_not
g61187 not n9325 ; n9325_not
g61188 not n8371 ; n8371_not
g61189 not n6634 ; n6634_not
g61190 not n4861 ; n4861_not
g61191 not n7039 ; n7039_not
g61192 not n7363 ; n7363_not
g61193 not n4906 ; n4906_not
g61194 not n5662 ; n5662_not
g61195 not n8803 ; n8803_not
g61196 not n5419 ; n5419_not
g61197 not n8119 ; n8119_not
g61198 not n8317 ; n8317_not
g61199 not n7930 ; n7930_not
g61200 not n6913 ; n6913_not
g61201 not n5671 ; n5671_not
g61202 not n7318 ; n7318_not
g61203 not n5644 ; n5644_not
g61204 not n7291 ; n7291_not
g61205 not n7372 ; n7372_not
g61206 not n5437 ; n5437_not
g61207 not n9505 ; n9505_not
g61208 not n7750 ; n7750_not
g61209 not n9343 ; n9343_not
g61210 not n6922 ; n6922_not
g61211 not n4852 ; n4852_not
g61212 not n5428 ; n5428_not
g61213 not n2359 ; n2359_not
g61214 not n5851 ; n5851_not
g61215 not n5653 ; n5653_not
g61216 not n6904 ; n6904_not
g61217 not n7309 ; n7309_not
g61218 not n8254 ; n8254_not
g61219 not n7741 ; n7741_not
g61220 not n3934 ; n3934_not
g61221 not n4744 ; n4744_not
g61222 not n6517 ; n6517_not
g61223 not n5914 ; n5914_not
g61224 not n9811 ; n9811_not
g61225 not n9262 ; n9262_not
g61226 not n3925 ; n3925_not
g61227 not n9541 ; n9541_not
g61228 not n7336 ; n7336_not
g61229 not n3916 ; n3916_not
g61230 not n8713 ; n8713_not
g61231 not n5482 ; n5482_not
g61232 not n7732 ; n7732_not
g61233 not n6841 ; n6841_not
g61234 not n3961 ; n3961_not
g61235 not n9253 ; n9253_not
g61236 not n8128 ; n8128_not
g61237 not n3484 ; n3484_not
g61238 not n3952 ; n3952_not
g61239 not n6616 ; n6616_not
g61240 not n5608 ; n5608_not
g61241 not n8704 ; n8704_not
g61242 not n7246 ; n7246_not
g61243 not n6508 ; n6508_not
g61244 not n7516 ; n7516_not
g61245 not n5923 ; n5923_not
g61246 not n3943 ; n3943_not
g61247 not n4834 ; n4834_not
g61248 not n4933 ; n4933_not
g61249 not n7255 ; n7255_not
g61250 not n4870 ; n4870_not
g61251 not n8731 ; n8731_not
g61252 not n6661 ; n6661_not
g61253 not n6544 ; n6544_not
g61254 not n1099 ; n1099_not
g61255 not n9280 ; n9280_not
g61256 not n3880 ; n3880_not
g61257 not n7264 ; n7264_not
g61258 not n7390 ; n7390_not
g61259 not n8281 ; n8281_not
g61260 not n6553 ; n6553_not
g61261 not n3871 ; n3871_not
g61262 not n7093 ; n7093_not
g61263 not n6526 ; n6526_not
g61264 not n3907 ; n3907_not
g61265 not n6850 ; n6850_not
g61266 not n8092 ; n8092_not
g61267 not n3772 ; n3772_not
g61268 not n8263 ; n8263_not
g61269 not n8470 ; n8470_not
g61270 not n9451 ; n9451_not
g61271 not n8722 ; n8722_not
g61272 not n7813 ; n7813_not
g61273 not n6535 ; n6535_not
g61274 not n8272 ; n8272_not
g61275 not n9271 ; n9271_not
g61276 not n4924 ; n4924_not
g61277 not n4843 ; n4843_not
g61278 not n4474 ; n4474_not
g61279 not n8551 ; n8551_not
g61280 not n6355 ; n6355_not
g61281 not n2854 ; n2854_not
g61282 not n9163 ; n9163_not
g61283 not n7561 ; n7561_not
g61284 not n2881 ; n2881_not
g61285 not n7444 ; n7444_not
g61286 not n2845 ; n2845_not
g61287 not n6625 ; n6625_not
g61288 not n7138 ; n7138_not
g61289 not n6292 ; n6292_not
g61290 not n1783 ; n1783_not
g61291 not n5239 ; n5239_not
g61292 not n6364 ; n6364_not
g61293 not n4465 ; n4465_not
g61294 not n2890 ; n2890_not
g61295 not n2836 ; n2836_not
g61296 not n8524 ; n8524_not
g61297 not n6760 ; n6760_not
g61298 not n2827 ; n2827_not
g61299 not n4456 ; n4456_not
g61300 not n5248 ; n5248_not
g61301 not n5059 ; n5059_not
g61302 not n4357 ; n4357_not
g61303 not n4447 ; n4447_not
g61304 not n8542 ; n8542_not
g61305 not n9154 ; n9154_not
g61306 not n2863 ; n2863_not
g61307 not n4672 ; n4672_not
g61308 not n6346 ; n6346_not
g61309 not n2872 ; n2872_not
g61310 not n7903 ; n7903_not
g61311 not n6805 ; n6805_not
g61312 not n7129 ; n7129_not
g61313 not n5275 ; n5275_not
g61314 not n9109 ; n9109_not
g61315 not n6256 ; n6256_not
g61316 not n9181 ; n9181_not
g61317 not n2737 ; n2737_not
g61318 not n2953 ; n2953_not
g61319 not n8560 ; n8560_not
g61320 not n1963 ; n1963_not
g61321 not n2692 ; n2692_not
g61322 not n5284 ; n5284_not
g61323 not n9046 ; n9046_not
g61324 not n1954 ; n1954_not
g61325 not n7174 ; n7174_not
g61326 not n2971 ; n2971_not
g61327 not n6382 ; n6382_not
g61328 not n4393 ; n4393_not
g61329 not n8515 ; n8515_not
g61330 not n5293 ; n5293_not
g61331 not n2728 ; n2728_not
g61332 not n4384 ; n4384_not
g61333 not n2980 ; n2980_not
g61334 not n8074 ; n8074_not
g61335 not n2818 ; n2818_not
g61336 not n2809 ; n2809_not
g61337 not n2908 ; n2908_not
g61338 not n2791 ; n2791_not
g61339 not n7570 ; n7570_not
g61340 not n8506 ; n8506_not
g61341 not n9172 ; n9172_not
g61342 not n1792 ; n1792_not
g61343 not n2782 ; n2782_not
g61344 not n7426 ; n7426_not
g61345 not n5257 ; n5257_not
g61346 not n7156 ; n7156_not
g61347 not n2773 ; n2773_not
g61348 not n4438 ; n4438_not
g61349 not n6373 ; n6373_not
g61350 not n9604 ; n9604_not
g61351 not n2926 ; n2926_not
g61352 not n4429 ; n4429_not
g61353 not n2764 ; n2764_not
g61354 not n5266 ; n5266_not
g61355 not n2935 ; n2935_not
g61356 not n2755 ; n2755_not
g61357 not n2746 ; n2746_not
g61358 not n8533 ; n8533_not
g61359 not n2656 ; n2656_not
g61360 not n4591 ; n4591_not
g61361 not n9028 ; n9028_not
g61362 not n7543 ; n7543_not
g61363 not n6319 ; n6319_not
g61364 not n7453 ; n7453_not
g61365 not n4645 ; n4645_not
g61366 not n9037 ; n9037_not
g61367 not n1972 ; n1972_not
g61368 not n6274 ; n6274_not
g61369 not n9136 ; n9136_not
g61370 not n9019 ; n9019_not
g61371 not n5842 ; n5842_not
g61372 not n2674 ; n2674_not
g61373 not n4627 ; n4627_not
g61374 not n9127 ; n9127_not
g61375 not n9631 ; n9631_not
g61376 not n7912 ; n7912_not
g61377 not n4618 ; n4618_not
g61378 not n2665 ; n2665_not
g61379 not n4636 ; n4636_not
g61380 not n4609 ; n4609_not
g61381 not n5086 ; n5086_not
g61382 not n1990 ; n1990_not
g61383 not n8920 ; n8920_not
g61384 not n5068 ; n5068_not
g61385 not n2629 ; n2629_not
g61386 not n1936 ; n1936_not
g61387 not n6337 ; n6337_not
g61388 not n5185 ; n5185_not
g61389 not n9460 ; n9460_not
g61390 not n4663 ; n4663_not
g61391 not n9712 ; n9712_not
g61392 not n5149 ; n5149_not
g61393 not n5194 ; n5194_not
g61394 not n9532 ; n9532_not
g61395 not n1756 ; n1756_not
g61396 not n6328 ; n6328_not
g61397 not n5158 ; n5158_not
g61398 not n4654 ; n4654_not
g61399 not n9145 ; n9145_not
g61400 not n1945 ; n1945_not
g61401 not n5176 ; n5176_not
g61402 not n9118 ; n9118_not
g61403 not n5356 ; n5356_not
g61404 not n1666 ; n1666_not
g61405 not n2179 ; n2179_not
g61406 not n1657 ; n1657_not
g61407 not n7066 ; n7066_not
g61408 not n7651 ; n7651_not
g61409 not n6409 ; n6409_not
g61410 not n5365 ; n5365_not
g61411 not n9721 ; n9721_not
g61412 not n1648 ; n1648_not
g61413 not n1495 ; n1495_not
g61414 not n5374 ; n5374_not
g61415 not n7840 ; n7840_not
g61416 not n4339 ; n4339_not
g61417 not n1693 ; n1693_not
g61418 not n7633 ; n7633_not
g61419 not n9523 ; n9523_not
g61420 not n5338 ; n5338_not
g61421 not n2683 ; n2683_not
g61422 not n1684 ; n1684_not
g61423 not n6670 ; n6670_not
g61424 not n5347 ; n5347_not
g61425 not n9208 ; n9208_not
g61426 not n7642 ; n7642_not
g61427 not n1675 ; n1675_not
g61428 not n1594 ; n1594_not
g61429 not n7408 ; n7408_not
g61430 not n9217 ; n9217_not
g61431 not n9550 ; n9550_not
g61432 not n1549 ; n1549_not
g61433 not n8605 ; n8605_not
g61434 not n1576 ; n1576_not
g61435 not n1567 ; n1567_not
g61436 not n1639 ; n1639_not
g61437 not n5383 ; n5383_not
g61438 not n7660 ; n7660_not
g61439 not n1477 ; n1477_not
g61440 not n2638 ; n2638_not
g61441 not n1486 ; n1486_not
g61442 not n6265 ; n6265_not
g61443 not n6418 ; n6418_not
g61444 not n8038 ; n8038_not
g61445 not n7606 ; n7606_not
g61446 not n5329 ; n5329_not
g61447 not n5077 ; n5077_not
g61448 not n7192 ; n7192_not
g61449 not n7615 ; n7615_not
g61450 not n2458 ; n2458_not
g61451 not n9334 ; n9334_not
g61452 not n9190 ; n9190_not
g61453 not n4708 ; n4708_not
g61454 not n1765 ; n1765_not
g61455 not n2944 ; n2944_not
g61456 not n7183 ; n7183_not
g61457 not n6391 ; n6391_not
g61458 not n7147 ; n7147_not
g61459 not n7417 ; n7417_not
g61460 not n7624 ; n7624_not
g61461 not n4366 ; n4366_not
g61462 not n7184 ; n7184_not
g61463 not n7067 ; n7067_not
g61464 not n7580 ; n7580_not
g61465 not n7661 ; n7661_not
g61466 not n6275 ; n6275_not
g61467 not n9641 ; n9641_not
g61468 not n8066 ; n8066_not
g61469 not n5834 ; n5834_not
g61470 not n7328 ; n7328_not
g61471 not n7670 ; n7670_not
g61472 not n8039 ; n8039_not
g61473 not n8057 ; n8057_not
g61474 not n5924 ; n5924_not
g61475 not n6752 ; n6752_not
g61476 not n6743 ; n6743_not
g61477 not n7508 ; n7508_not
g61478 not n6086 ; n6086_not
g61479 not n7715 ; n7715_not
g61480 not n6509 ; n6509_not
g61481 not n9605 ; n9605_not
g61482 not n6329 ; n6329_not
g61483 not n7463 ; n7463_not
g61484 not n9425 ; n9425_not
g61485 not n5843 ; n5843_not
g61486 not n9416 ; n9416_not
g61487 not n7319 ; n7319_not
g61488 not n5555 ; n5555_not
g61489 not n7724 ; n7724_not
g61490 not n6437 ; n6437_not
g61491 not n6419 ; n6419_not
g61492 not n7247 ; n7247_not
g61493 not n6095 ; n6095_not
g61494 not n7823 ; n7823_not
g61495 not n8048 ; n8048_not
g61496 not n6185 ; n6185_not
g61497 not n7058 ; n7058_not
g61498 not n7706 ; n7706_not
g61499 not n6428 ; n6428_not
g61500 not n6617 ; n6617_not
g61501 not n6068 ; n6068_not
g61502 not n6167 ; n6167_not
g61503 not n9650 ; n9650_not
g61504 not n7904 ; n7904_not
g61505 not n7049 ; n7049_not
g61506 not n6383 ; n6383_not
g61507 not n7418 ; n7418_not
g61508 not n6077 ; n6077_not
g61509 not n6392 ; n6392_not
g61510 not n7922 ; n7922_not
g61511 not n6257 ; n6257_not
g61512 not n6707 ; n6707_not
g61513 not n6158 ; n6158_not
g61514 not n9632 ; n9632_not
g61515 not n7940 ; n7940_not
g61516 not n7544 ; n7544_not
g61517 not n7535 ; n7535_not
g61518 not n6284 ; n6284_not
g61519 not n7355 ; n7355_not
g61520 not n7157 ; n7157_not
g61521 not n7337 ; n7337_not
g61522 not n7238 ; n7238_not
g61523 not n6626 ; n6626_not
g61524 not n6149 ; n6149_not
g61525 not n7094 ; n7094_not
g61526 not n7616 ; n7616_not
g61527 not n6239 ; n6239_not
g61528 not n5951 ; n5951_not
g61529 not n9623 ; n9623_not
g61530 not n9560 ; n9560_not
g61531 not n7175 ; n7175_not
g61532 not n7733 ; n7733_not
g61533 not n6491 ; n6491_not
g61534 not n7346 ; n7346_not
g61535 not n5960 ; n5960_not
g61536 not n7607 ; n7607_not
g61537 not n6554 ; n6554_not
g61538 not n6464 ; n6464_not
g61539 not n7571 ; n7571_not
g61540 not n6473 ; n6473_not
g61541 not n9614 ; n9614_not
g61542 not n7805 ; n7805_not
g61543 not n7454 ; n7454_not
g61544 not n7841 ; n7841_not
g61545 not n7526 ; n7526_not
g61546 not n7139 ; n7139_not
g61547 not n7076 ; n7076_not
g61548 not n6527 ; n6527_not
g61549 not n6716 ; n6716_not
g61550 not n6347 ; n6347_not
g61551 not n7274 ; n7274_not
g61552 not n7382 ; n7382_not
g61553 not n7643 ; n7643_not
g61554 not n5807 ; n5807_not
g61555 not n7481 ; n7481_not
g61556 not n6671 ; n6671_not
g61557 not n7832 ; n7832_not
g61558 not n9461 ; n9461_not
g61559 not n6536 ; n6536_not
g61560 not n6365 ; n6365_not
g61561 not n7193 ; n7193_not
g61562 not n7634 ; n7634_not
g61563 not n7256 ; n7256_not
g61564 not n7436 ; n7436_not
g61565 not n7148 ; n7148_not
g61566 not n5906 ; n5906_not
g61567 not n7409 ; n7409_not
g61568 not n7814 ; n7814_not
g61569 not n6545 ; n6545_not
g61570 not n9434 ; n9434_not
g61571 not n6662 ; n6662_not
g61572 not n6059 ; n6059_not
g61573 not n7265 ; n7265_not
g61574 not n7391 ; n7391_not
g61575 not n6356 ; n6356_not
g61576 not n9551 ; n9551_not
g61577 not n6725 ; n6725_not
g61578 not n6446 ; n6446_not
g61579 not n7166 ; n7166_not
g61580 not n7751 ; n7751_not
g61581 not n9506 ; n9506_not
g61582 not n5852 ; n5852_not
g61583 not n6644 ; n6644_not
g61584 not n7490 ; n7490_not
g61585 not n6482 ; n6482_not
g61586 not n5564 ; n5564_not
g61587 not n7364 ; n7364_not
g61588 not n7850 ; n7850_not
g61589 not n7553 ; n7553_not
g61590 not n7760 ; n7760_not
g61591 not n6635 ; n6635_not
g61592 not n5861 ; n5861_not
g61593 not n6680 ; n6680_not
g61594 not n5942 ; n5942_not
g61595 not n7283 ; n7283_not
g61596 not n6455 ; n6455_not
g61597 not n6266 ; n6266_not
g61598 not n7229 ; n7229_not
g61599 not n6590 ; n6590_not
g61600 not n6194 ; n6194_not
g61601 not n6374 ; n6374_not
g61602 not n7373 ; n7373_not
g61603 not n7652 ; n7652_not
g61604 not n6338 ; n6338_not
g61605 not n6518 ; n6518_not
g61606 not n7292 ; n7292_not
g61607 not n7625 ; n7625_not
g61608 not n7742 ; n7742_not
g61609 not n2594 ; n2594_not
g61610 not n1757 ; n1757_not
g61611 not n2378 ; n2378_not
g61612 not n3845 ; n3845_not
g61613 not n8183 ; n8183_not
g61614 not n2585 ; n2585_not
g61615 not n4880 ; n4880_not
g61616 not n8516 ; n8516_not
g61617 not n8174 ; n8174_not
g61618 not n8453 ; n8453_not
g61619 not n1775 ; n1775_not
g61620 not n4871 ; n4871_not
g61621 not n8381 ; n8381_not
g61622 not n2576 ; n2576_not
g61623 not n8165 ; n8165_not
g61624 not n8309 ; n8309_not
g61625 not n3854 ; n3854_not
g61626 not n4862 ; n4862_not
g61627 not n4781 ; n4781_not
g61628 not n8219 ; n8219_not
g61629 not n8327 ; n8327_not
g61630 not n3791 ; n3791_not
g61631 not n2558 ; n2558_not
g61632 not n8318 ; n8318_not
g61633 not n3809 ; n3809_not
g61634 not n1577 ; n1577_not
g61635 not n4907 ; n4907_not
g61636 not n3818 ; n3818_not
g61637 not n1568 ; n1568_not
g61638 not n8435 ; n8435_not
g61639 not n3827 ; n3827_not
g61640 not n2567 ; n2567_not
g61641 not n3836 ; n3836_not
g61642 not n8192 ; n8192_not
g61643 not n1739 ; n1739_not
g61644 not n1748 ; n1748_not
g61645 not n4484 ; n4484_not
g61646 not n9470 ; n9470_not
g61647 not n4808 ; n4808_not
g61648 not n1793 ; n1793_not
g61649 not n4493 ; n4493_not
g61650 not n8291 ; n8291_not
g61651 not n4790 ; n4790_not
g61652 not n8093 ; n8093_not
g61653 not n3881 ; n3881_not
g61654 not n4763 ; n4763_not
g61655 not n1829 ; n1829_not
g61656 not n8084 ; n8084_not
g61657 not n8282 ; n8282_not
g61658 not n2549 ; n2549_not
g61659 not n3782 ; n3782_not
g61660 not n9803 ; n9803_not
g61661 not n8156 ; n8156_not
g61662 not n4853 ; n4853_not
g61663 not n8147 ; n8147_not
g61664 not n3863 ; n3863_not
g61665 not n4844 ; n4844_not
g61666 not n8138 ; n8138_not
g61667 not n4835 ; n4835_not
g61668 not n8471 ; n8471_not
g61669 not n8129 ; n8129_not
g61670 not n3872 ; n3872_not
g61671 not n4826 ; n4826_not
g61672 not n8480 ; n8480_not
g61673 not n8390 ; n8390_not
g61674 not n4817 ; n4817_not
g61675 not n3683 ; n3683_not
g61676 not n8354 ; n8354_not
g61677 not n2477 ; n2477_not
g61678 not n3692 ; n3692_not
g61679 not n4691 ; n4691_not
g61680 not n1586 ; n1586_not
g61681 not n2486 ; n2486_not
g61682 not n1649 ; n1649_not
g61683 not n1658 ; n1658_not
g61684 not n1667 ; n1667_not
g61685 not n4709 ; n4709_not
g61686 not n8822 ; n8822_not
g61687 not n8345 ; n8345_not
g61688 not n3656 ; n3656_not
g61689 not n3665 ; n3665_not
g61690 not n5096 ; n5096_not
g61691 not n3674 ; n3674_not
g61692 not n1388 ; n1388_not
g61693 not n2468 ; n2468_not
g61694 not n8336 ; n8336_not
g61695 not n8363 ; n8363_not
g61696 not n1559 ; n1559_not
g61697 not n5078 ; n5078_not
g61698 not n8813 ; n8813_not
g61699 not n5069 ; n5069_not
g61700 not n3764 ; n3764_not
g61701 not n4952 ; n4952_not
g61702 not n8237 ; n8237_not
g61703 not n3773 ; n3773_not
g61704 not n1694 ; n1694_not
g61705 not n4943 ; n4943_not
g61706 not n8228 ; n8228_not
g61707 not n4736 ; n4736_not
g61708 not n4934 ; n4934_not
g61709 not n4925 ; n4925_not
g61710 not n2648 ; n2648_not
g61711 not n4745 ; n4745_not
g61712 not n9704 ; n9704_not
g61713 not n8426 ; n8426_not
g61714 not n4916 ; n4916_not
g61715 not n4754 ; n4754_not
g61716 not n3719 ; n3719_not
g61717 not n8273 ; n8273_not
g61718 not n8264 ; n8264_not
g61719 not n1676 ; n1676_not
g61720 not n2675 ; n2675_not
g61721 not n8255 ; n8255_not
g61722 not n8408 ; n8408_not
g61723 not n3728 ; n3728_not
g61724 not n1685 ; n1685_not
g61725 not n4970 ; n4970_not
g61726 not n8246 ; n8246_not
g61727 not n3746 ; n3746_not
g61728 not n2495 ; n2495_not
g61729 not n4961 ; n4961_not
g61730 not n2666 ; n2666_not
g61731 not n4466 ; n4466_not
g61732 not n1964 ; n1964_not
g61733 not n4079 ; n4079_not
g61734 not n4088 ; n4088_not
g61735 not n4448 ; n4448_not
g61736 not n4169 ; n4169_not
g61737 not n4439 ; n4439_not
g61738 not n4178 ; n4178_not
g61739 not n1982 ; n1982_not
g61740 not n9821 ; n9821_not
g61741 not n4187 ; n4187_not
g61742 not n9902 ; n9902_not
g61743 not n8921 ; n8921_not
g61744 not n4196 ; n4196_not
g61745 not n4394 ; n4394_not
g61746 not n4475 ; n4475_not
g61747 not n9731 ; n9731_not
g61748 not n1937 ; n1937_not
g61749 not n1955 ; n1955_not
g61750 not n8444 ; n8444_not
g61751 not n4457 ; n4457_not
g61752 not n4097 ; n4097_not
g61753 not n4295 ; n4295_not
g61754 not n9722 ; n9722_not
g61755 not n4286 ; n4286_not
g61756 not n4277 ; n4277_not
g61757 not n4259 ; n4259_not
g61758 not n4268 ; n4268_not
g61759 not n2099 ; n2099_not
g61760 not n2189 ; n2189_not
g61761 not n8930 ; n8930_not
g61762 not n1973 ; n1973_not
g61763 not n4376 ; n4376_not
g61764 not n9524 ; n9524_not
g61765 not n4358 ; n4358_not
g61766 not n4349 ; n4349_not
g61767 not n3917 ; n3917_not
g61768 not n1856 ; n1856_not
g61769 not n3926 ; n3926_not
g61770 not n9713 ; n9713_not
g61771 not n4367 ; n4367_not
g61772 not n3935 ; n3935_not
g61773 not n9740 ; n9740_not
g61774 not n3944 ; n3944_not
g61775 not n1838 ; n1838_not
g61776 not n3890 ; n3890_not
g61777 not n4718 ; n4718_not
g61778 not n8075 ; n8075_not
g61779 not n1847 ; n1847_not
g61780 not n4682 ; n4682_not
g61781 not n3908 ; n3908_not
g61782 not n9371 ; n9371_not
g61783 not n8525 ; n8525_not
g61784 not n1892 ; n1892_not
g61785 not n2387 ; n2387_not
g61786 not n9515 ; n9515_not
g61787 not n1919 ; n1919_not
g61788 not n3953 ; n3953_not
g61789 not n1865 ; n1865_not
g61790 not n3962 ; n3962_not
g61791 not n1874 ; n1874_not
g61792 not n2459 ; n2459_not
g61793 not n3737 ; n3737_not
g61794 not n3971 ; n3971_not
g61795 not n8534 ; n8534_not
g61796 not n1883 ; n1883_not
g61797 not n3980 ; n3980_not
g61798 not n1766 ; n1766_not
g61799 not n3287 ; n3287_not
g61800 not n5519 ; n5519_not
g61801 not n5528 ; n5528_not
g61802 not n3278 ; n3278_not
g61803 not n5537 ; n5537_not
g61804 not n5546 ; n5546_not
g61805 not n3269 ; n3269_not
g61806 not n9344 ; n9344_not
g61807 not n9326 ; n9326_not
g61808 not n9335 ; n9335_not
g61809 not n2891 ; n2891_not
g61810 not n2918 ; n2918_not
g61811 not n2990 ; n2990_not
g61812 not n3197 ; n3197_not
g61813 not n5492 ; n5492_not
g61814 not n3188 ; n3188_not
g61815 not n5339 ; n5339_not
g61816 not n3395 ; n3395_not
g61817 not n5348 ; n5348_not
g61818 not n2828 ; n2828_not
g61819 not n5357 ; n5357_not
g61820 not n5366 ; n5366_not
g61821 not n3386 ; n3386_not
g61822 not n2837 ; n2837_not
g61823 not n8840 ; n8840_not
g61824 not n5375 ; n5375_not
g61825 not n3377 ; n3377_not
g61826 not n2846 ; n2846_not
g61827 not n3368 ; n3368_not
g61828 not n2864 ; n2864_not
g61829 not n5483 ; n5483_not
g61830 not n3296 ; n3296_not
g61831 not n5474 ; n5474_not
g61832 not n9317 ; n9317_not
g61833 not n8903 ; n8903_not
g61834 not n2873 ; n2873_not
g61835 not n5456 ; n5456_not
g61836 not n5438 ; n5438_not
g61837 not n5429 ; n5429_not
g61838 not n8831 ; n8831_not
g61839 not n2855 ; n2855_not
g61840 not n3359 ; n3359_not
g61841 not n2954 ; n2954_not
g61842 not n2819 ; n2819_not
g61843 not n2909 ; n2909_not
g61844 not n2981 ; n2981_not
g61845 not n2792 ; n2792_not
g61846 not n2738 ; n2738_not
g61847 not n2783 ; n2783_not
g61848 not n5780 ; n5780_not
g61849 not n2774 ; n2774_not
g61850 not n9542 ; n9542_not
g61851 not n2765 ; n2765_not
g61852 not n2945 ; n2945_not
g61853 not n2936 ; n2936_not
g61854 not n2756 ; n2756_not
g61855 not n5816 ; n5816_not
g61856 not n2747 ; n2747_not
g61857 not n3089 ; n3089_not
g61858 not n3098 ; n3098_not
g61859 not n9353 ; n9353_not
g61860 not n9911 ; n9911_not
g61861 not n5447 ; n5447_not
g61862 not n2729 ; n2729_not
g61863 not n9380 ; n9380_not
g61864 not n1289 ; n1289_not
g61865 not n1298 ; n1298_not
g61866 not n3593 ; n3593_not
g61867 not n3494 ; n3494_not
g61868 not n5177 ; n5177_not
g61869 not n5087 ; n5087_not
g61870 not n5159 ; n5159_not
g61871 not n3638 ; n3638_not
g61872 not n5168 ; n5168_not
g61873 not n5267 ; n5267_not
g61874 not n3575 ; n3575_not
g61875 not n1469 ; n1469_not
g61876 not n9443 ; n9443_not
g61877 not n5186 ; n5186_not
g61878 not n5294 ; n5294_not
g61879 not n3476 ; n3476_not
g61880 not n2684 ; n2684_not
g61881 not n3548 ; n3548_not
g61882 not n3539 ; n3539_not
g61883 not n5276 ; n5276_not
g61884 not n3485 ; n3485_not
g61885 not n9533 ; n9533_not
g61886 not n3557 ; n3557_not
g61887 not n3629 ; n3629_not
g61888 not n5285 ; n5285_not
g61889 not n3458 ; n3458_not
g61890 not n2639 ; n2639_not
g61891 not n1199 ; n1199_not
g61892 not n7913 ; n7913_not
g61893 not n5258 ; n5258_not
g61894 not n3584 ; n3584_not
g61895 not n3449 ; n3449_not
g61896 not n1397 ; n1397_not
g61897 not n3647 ; n3647_not
g61898 not n5195 ; n5195_not
g61899 not n5249 ; n5249_not
g61900 not n3566 ; n3566_not
g61901 not n7581 ; n7581_not
g61902 not n8931 ; n8931_not
g61903 not n9516 ; n9516_not
g61904 not n8436 ; n8436_not
g61905 not n6087 ; n6087_not
g61906 not n6474 ; n6474_not
g61907 not n2739 ; n2739_not
g61908 not n8805 ; n8805_not
g61909 not n8652 ; n8652_not
g61910 not n6681 ; n6681_not
g61911 not n3594 ; n3594_not
g61912 not n7518 ; n7518_not
g61913 not n3693 ; n3693_not
g61914 not n9084 ; n9084_not
g61915 not n6816 ; n6816_not
g61916 not n2856 ; n2856_not
g61917 not n9813 ; n9813_not
g61918 not n8634 ; n8634_not
g61919 not n6636 ; n6636_not
g61920 not n8661 ; n8661_not
g61921 not n6672 ; n6672_not
g61922 not n9039 ; n9039_not
g61923 not n2874 ; n2874_not
g61924 not n3585 ; n3585_not
g61925 not n3819 ; n3819_not
g61926 not n3990 ; n3990_not
g61927 not n2748 ; n2748_not
g61928 not n2757 ; n2757_not
g61929 not n2397 ; n2397_not
g61930 not n3981 ; n3981_not
g61931 not n6492 ; n6492_not
g61932 not n7509 ; n7509_not
g61933 not n3729 ; n3729_not
g61934 not n6906 ; n6906_not
g61935 not n7536 ; n7536_not
g61936 not n3972 ; n3972_not
g61937 not n3099 ; n3099_not
g61938 not n8670 ; n8670_not
g61939 not n6096 ; n6096_not
g61940 not n9732 ; n9732_not
g61941 not n9606 ; n9606_not
g61942 not n8841 ; n8841_not
g61943 not n2676 ; n2676_not
g61944 not n2478 ; n2478_not
g61945 not n2955 ; n2955_not
g61946 not n8643 ; n8643_not
g61947 not n6483 ; n6483_not
g61948 not n6807 ; n6807_not
g61949 not n6690 ; n6690_not
g61950 not n2946 ; n2946_not
g61951 not n6852 ; n6852_not
g61952 not n9822 ; n9822_not
g61953 not n3666 ; n3666_not
g61954 not n9318 ; n9318_not
g61955 not n4098 ; n4098_not
g61956 not n1938 ; n1938_not
g61957 not n9048 ; n9048_not
g61958 not n4197 ; n4197_not
g61959 not n2784 ; n2784_not
g61960 not n4188 ; n4188_not
g61961 not n2793 ; n2793_not
g61962 not n3675 ; n3675_not
g61963 not n8616 ; n8616_not
g61964 not n7068 ; n7068_not
g61965 not n6438 ; n6438_not
g61966 not n4179 ; n4179_not
g61967 not n6843 ; n6843_not
g61968 not n8607 ; n8607_not
g61969 not n2919 ; n2919_not
g61970 not n2199 ; n2199_not
g61971 not n2991 ; n2991_not
g61972 not n3648 ; n3648_not
g61973 not n8535 ; n8535_not
g61974 not n7464 ; n7464_not
g61975 not n8571 ; n8571_not
g61976 not n6861 ; n6861_not
g61977 not n8580 ; n8580_not
g61978 not n6870 ; n6870_not
g61979 not n8562 ; n8562_not
g61980 not n4089 ; n4089_not
g61981 not n2766 ; n2766_not
g61982 not n3657 ; n3657_not
g61983 not n6429 ; n6429_not
g61984 not n2694 ; n2694_not
g61985 not n6654 ; n6654_not
g61986 not n3639 ; n3639_not
g61987 not n2775 ; n2775_not
g61988 not n2973 ; n2973_not
g61989 not n2685 ; n2685_not
g61990 not n2469 ; n2469_not
g61991 not n8445 ; n8445_not
g61992 not n9093 ; n9093_not
g61993 not n6456 ; n6456_not
g61994 not n2289 ; n2289_not
g61995 not n8940 ; n8940_not
g61996 not n2298 ; n2298_not
g61997 not n2847 ; n2847_not
g61998 not n6078 ; n6078_not
g61999 not n6825 ; n6825_not
g62000 not n9471 ; n9471_not
g62001 not n7590 ; n7590_not
g62002 not n6591 ; n6591_not
g62003 not n9336 ; n9336_not
g62004 not n3684 ; n3684_not
g62005 not n6465 ; n6465_not
g62006 not n8814 ; n8814_not
g62007 not n8625 ; n8625_not
g62008 not n3459 ; n3459_not
g62009 not n7059 ; n7059_not
g62010 not n8553 ; n8553_not
g62011 not n6447 ; n6447_not
g62012 not n2829 ; n2829_not
g62013 not n8454 ; n8454_not
g62014 not n8544 ; n8544_not
g62015 not n6834 ; n6834_not
g62016 not n2838 ; n2838_not
g62017 not n6069 ; n6069_not
g62018 not n8832 ; n8832_not
g62019 not n6645 ; n6645_not
g62020 not n3873 ; n3873_not
g62021 not n3297 ; n3297_not
g62022 not n3549 ; n3549_not
g62023 not n3792 ; n3792_not
g62024 not n6933 ; n6933_not
g62025 not n6753 ; n6753_not
g62026 not n9345 ; n9345_not
g62027 not n8742 ; n8742_not
g62028 not n2658 ; n2658_not
g62029 not n3864 ; n3864_not
g62030 not n3783 ; n3783_not
g62031 not n8706 ; n8706_not
g62032 not n9480 ; n9480_not
g62033 not n2865 ; n2865_not
g62034 not n8751 ; n8751_not
g62035 not n8715 ; n8715_not
g62036 not n2568 ; n2568_not
g62037 not n3882 ; n3882_not
g62038 not n3279 ; n3279_not
g62039 not n6546 ; n6546_not
g62040 not n2883 ; n2883_not
g62041 not n6762 ; n6762_not
g62042 not n9615 ; n9615_not
g62043 not n9804 ; n9804_not
g62044 not n3558 ; n3558_not
g62045 not n2559 ; n2559_not
g62046 not n6186 ; n6186_not
g62047 not n7563 ; n7563_not
g62048 not n6960 ; n6960_not
g62049 not n3288 ; n3288_not
g62050 not n3495 ; n3495_not
g62051 not n3774 ; n3774_not
g62052 not n8391 ; n8391_not
g62053 not n3198 ; n3198_not
g62054 not n6555 ; n6555_not
g62055 not n3846 ; n3846_not
g62056 not n7491 ; n7491_not
g62057 not n3468 ; n3468_not
g62058 not n3387 ; n3387_not
g62059 not n8760 ; n8760_not
g62060 not n2577 ; n2577_not
g62061 not n6726 ; n6726_not
g62062 not n8733 ; n8733_not
g62063 not n2595 ; n2595_not
g62064 not n9354 ; n9354_not
g62065 not n3837 ; n3837_not
g62066 not n6717 ; n6717_not
g62067 not n6951 ; n6951_not
g62068 not n3828 ; n3828_not
g62069 not n3855 ; n3855_not
g62070 not n6609 ; n6609_not
g62071 not n6744 ; n6744_not
g62072 not n6573 ; n6573_not
g62073 not n3369 ; n3369_not
g62074 not n6942 ; n6942_not
g62075 not n8724 ; n8724_not
g62076 not n9561 ; n9561_not
g62077 not n3486 ; n3486_not
g62078 not n2586 ; n2586_not
g62079 not n2388 ; n2388_not
g62080 not n2649 ; n2649_not
g62081 not n9057 ; n9057_not
g62082 not n3378 ; n3378_not
g62083 not n6582 ; n6582_not
g62084 not n9570 ; n9570_not
g62085 not n9075 ; n9075_not
g62086 not n6627 ; n6627_not
g62087 not n3936 ; n3936_not
g62088 not n9741 ; n9741_not
g62089 not n7545 ; n7545_not
g62090 not n6915 ; n6915_not
g62091 not n6519 ; n6519_not
g62092 not n3927 ; n3927_not
g62093 not n8409 ; n8409_not
g62094 not n2487 ; n2487_not
g62095 not n2928 ; n2928_not
g62096 not n8850 ; n8850_not
g62097 not n3963 ; n3963_not
g62098 not n9750 ; n9750_not
g62099 not n3576 ; n3576_not
g62100 not n3738 ; n3738_not
g62101 not n9912 ; n9912_not
g62102 not n7554 ; n7554_not
g62103 not n3954 ; n3954_not
g62104 not n3747 ; n3747_not
g62105 not n3945 ; n3945_not
g62106 not n6771 ; n6771_not
g62107 not n8364 ; n8364_not
g62108 not n8913 ; n8913_not
g62109 not n9066 ; n9066_not
g62110 not n3891 ; n3891_not
g62111 not n9426 ; n9426_not
g62112 not n6537 ; n6537_not
g62113 not n3756 ; n3756_not
g62114 not n6159 ; n6159_not
g62115 not n6168 ; n6168_not
g62116 not n6195 ; n6195_not
g62117 not n8355 ; n8355_not
g62118 not n3918 ; n3918_not
g62119 not n6780 ; n6780_not
g62120 not n2496 ; n2496_not
g62121 not n2982 ; n2982_not
g62122 not n3909 ; n3909_not
g62123 not n3567 ; n3567_not
g62124 not n6528 ; n6528_not
g62125 not n6924 ; n6924_not
g62126 not n5097 ; n5097_not
g62127 not n7914 ; n7914_not
g62128 not n9255 ; n9255_not
g62129 not n5169 ; n5169_not
g62130 not n5286 ; n5286_not
g62131 not n1299 ; n1299_not
g62132 not n7239 ; n7239_not
g62133 not n5277 ; n5277_not
g62134 not n5268 ; n5268_not
g62135 not n9246 ; n9246_not
g62136 not n7905 ; n7905_not
g62137 not n5259 ; n5259_not
g62138 not n5862 ; n5862_not
g62139 not n9534 ; n9534_not
g62140 not n5853 ; n5853_not
g62141 not n9237 ; n9237_not
g62142 not n5196 ; n5196_not
g62143 not n5187 ; n5187_not
g62144 not n7392 ; n7392_not
g62145 not n5376 ; n5376_not
g62146 not n9282 ; n9282_not
g62147 not n5367 ; n5367_not
g62148 not n5358 ; n5358_not
g62149 not n5349 ; n5349_not
g62150 not n7257 ; n7257_not
g62151 not n9273 ; n9273_not
g62152 not n5079 ; n5079_not
g62153 not n9264 ; n9264_not
g62154 not n9651 ; n9651_not
g62155 not n7923 ; n7923_not
g62156 not n5088 ; n5088_not
g62157 not n7248 ; n7248_not
g62158 not n5295 ; n5295_not
g62159 not n4971 ; n4971_not
g62160 not n5817 ; n5817_not
g62161 not n4962 ; n4962_not
g62162 not n8418 ; n8418_not
g62163 not n4953 ; n4953_not
g62164 not n1587 ; n1587_not
g62165 not n5808 ; n5808_not
g62166 not n4944 ; n4944_not
g62167 not n4935 ; n4935_not
g62168 not n4926 ; n4926_not
g62169 not n4746 ; n4746_not
g62170 not n7194 ; n7194_not
g62171 not n4917 ; n4917_not
g62172 not n9903 ; n9903_not
g62173 not n1578 ; n1578_not
g62174 not n4908 ; n4908_not
g62175 not n4755 ; n4755_not
g62176 not n9705 ; n9705_not
g62177 not n4764 ; n4764_not
g62178 not n9552 ; n9552_not
g62179 not n1569 ; n1569_not
g62180 not n5781 ; n5781_not
g62181 not n7185 ; n7185_not
g62182 not n7950 ; n7950_not
g62183 not n9192 ; n9192_not
g62184 not n4890 ; n4890_not
g62185 not n1749 ; n1749_not
g62186 not n5178 ; n5178_not
g62187 not n1479 ; n1479_not
g62188 not n5844 ; n5844_not
g62189 not n1488 ; n1488_not
g62190 not n8346 ; n8346_not
g62191 not n9228 ; n9228_not
g62192 not n1497 ; n1497_not
g62193 not n1398 ; n1398_not
g62194 not n9219 ; n9219_not
g62195 not n9435 ; n9435_not
g62196 not n8373 ; n8373_not
g62197 not n9381 ; n9381_not
g62198 not n4683 ; n4683_not
g62199 not n1596 ; n1596_not
g62200 not n4980 ; n4980_not
g62201 not n4719 ; n4719_not
g62202 not n9642 ; n9642_not
g62203 not n9156 ; n9156_not
g62204 not n5664 ; n5664_not
g62205 not n5745 ; n5745_not
g62206 not n5736 ; n5736_not
g62207 not n5655 ; n5655_not
g62208 not n9165 ; n9165_not
g62209 not n5727 ; n5727_not
g62210 not n5646 ; n5646_not
g62211 not n9174 ; n9174_not
g62212 not n5718 ; n5718_not
g62213 not n5871 ; n5871_not
g62214 not n5439 ; n5439_not
g62215 not n5637 ; n5637_not
g62216 not n5709 ; n5709_not
g62217 not n9390 ; n9390_not
g62218 not n7329 ; n7329_not
g62219 not n5628 ; n5628_not
g62220 not n9183 ; n9183_not
g62221 not n5448 ; n5448_not
g62222 not n9444 ; n9444_not
g62223 not n5619 ; n5619_not
g62224 not n5691 ; n5691_not
g62225 not n5457 ; n5457_not
g62226 not n5682 ; n5682_not
g62227 not n9921 ; n9921_not
g62228 not n5673 ; n5673_not
g62229 not n5826 ; n5826_not
g62230 not n5754 ; n5754_not
g62231 not n9543 ; n9543_not
g62232 not n5763 ; n5763_not
g62233 not n5772 ; n5772_not
g62234 not n7356 ; n7356_not
g62235 not n5790 ; n5790_not
g62236 not n7347 ; n7347_not
g62237 not n9129 ; n9129_not
g62238 not n9138 ; n9138_not
g62239 not n9408 ; n9408_not
g62240 not n9147 ; n9147_not
g62241 not n7338 ; n7338_not
g62242 not n9660 ; n9660_not
g62243 not n5565 ; n5565_not
g62244 not n7374 ; n7374_not
g62245 not n5529 ; n5529_not
g62246 not n7284 ; n7284_not
g62247 not n5952 ; n5952_not
g62248 not n5907 ; n5907_not
g62249 not n9291 ; n9291_not
g62250 not n5493 ; n5493_not
g62251 not n5961 ; n5961_not
g62252 not n7383 ; n7383_not
g62253 not n5484 ; n5484_not
g62254 not n8067 ; n8067_not
g62255 not n7275 ; n7275_not
g62256 not n5466 ; n5466_not
g62257 not n5970 ; n5970_not
g62258 not n8058 ; n8058_not
g62259 not n7266 ; n7266_not
g62260 not n5394 ; n5394_not
g62261 not n9363 ; n9363_not
g62262 not n5592 ; n5592_not
g62263 not n5583 ; n5583_not
g62264 not n7077 ; n7077_not
g62265 not n5574 ; n5574_not
g62266 not n7365 ; n7365_not
g62267 not n5916 ; n5916_not
g62268 not n5934 ; n5934_not
g62269 not n7293 ; n7293_not
g62270 not n4287 ; n4287_not
g62271 not n1866 ; n1866_not
g62272 not n7437 ; n7437_not
g62273 not n6294 ; n6294_not
g62274 not n9831 ; n9831_not
g62275 not n1776 ; n1776_not
g62276 not n1875 ; n1875_not
g62277 not n4278 ; n4278_not
g62278 not n7446 ; n7446_not
g62279 not n4269 ; n4269_not
g62280 not n1767 ; n1767_not
g62281 not n1884 ; n1884_not
g62282 not n4593 ; n4593_not
g62283 not n1893 ; n1893_not
g62284 not n5943 ; n5943_not
g62285 not n4584 ; n4584_not
g62286 not n4575 ; n4575_not
g62287 not n1758 ; n1758_not
g62288 not n4566 ; n4566_not
g62289 not n4557 ; n4557_not
g62290 not n4548 ; n4548_not
g62291 not n7149 ; n7149_not
g62292 not n4728 ; n4728_not
g62293 not n4629 ; n4629_not
g62294 not n4638 ; n4638_not
g62295 not n4647 ; n4647_not
g62296 not n8508 ; n8508_not
g62297 not n4656 ; n4656_not
g62298 not n4665 ; n4665_not
g62299 not n6249 ; n6249_not
g62300 not n4674 ; n4674_not
g62301 not n8904 ; n8904_not
g62302 not n4692 ; n4692_not
g62303 not n1848 ; n1848_not
g62304 not n4359 ; n4359_not
g62305 not n6267 ; n6267_not
g62306 not n1857 ; n1857_not
g62307 not n9714 ; n9714_not
g62308 not n6276 ; n6276_not
g62309 not n4368 ; n4368_not
g62310 not n4296 ; n4296_not
g62311 not n9633 ; n9633_not
g62312 not n4377 ; n4377_not
g62313 not n6375 ; n6375_not
g62314 not n7455 ; n7455_not
g62315 not n1992 ; n1992_not
g62316 not n6285 ; n6285_not
g62317 not n6384 ; n6384_not
g62318 not n9525 ; n9525_not
g62319 not n4386 ; n4386_not
g62320 not n7086 ; n7086_not
g62321 not n1983 ; n1983_not
g62322 not n6393 ; n6393_not
g62323 not n1974 ; n1974_not
g62324 not n8481 ; n8481_not
g62325 not n1965 ; n1965_not
g62326 not n9624 ; n9624_not
g62327 not n9723 ; n9723_not
g62328 not n7473 ; n7473_not
g62329 not n4539 ; n4539_not
g62330 not n6339 ; n6339_not
g62331 not n1947 ; n1947_not
g62332 not n4449 ; n4449_not
g62333 not n6348 ; n6348_not
g62334 not n4494 ; n4494_not
g62335 not n4467 ; n4467_not
g62336 not n4458 ; n4458_not
g62337 not n6357 ; n6357_not
g62338 not n6366 ; n6366_not
g62339 not n8490 ; n8490_not
g62340 not n4791 ; n4791_not
g62341 not n4836 ; n4836_not
g62342 not n4827 ; n4827_not
g62343 not n4809 ; n4809_not
g62344 not n7167 ; n7167_not
g62345 not n4818 ; n4818_not
g62346 not n4773 ; n4773_not
g62347 not n7158 ; n7158_not
g62348 not n7419 ; n7419_not
g62349 not n4881 ; n4881_not
g62350 not n7176 ; n7176_not
g62351 not n4872 ; n4872_not
g62352 not n9453 ; n9453_not
g62353 not n7932 ; n7932_not
g62354 not n4863 ; n4863_not
g62355 not n8463 ; n8463_not
g62356 not n4854 ; n4854_not
g62357 not n1785 ; n1785_not
g62358 not n4845 ; n4845_not
g62359 not n1839 ; n1839_not
g62360 not n7159 ; n7159_not
g62361 not n1696 ; n1696_not
g62362 not n2389 ; n2389_not
g62363 not n7528 ; n7528_not
g62364 not n2956 ; n2956_not
g62365 not n9643 ; n9643_not
g62366 not n8581 ; n8581_not
g62367 not n9373 ; n9373_not
g62368 not n9067 ; n9067_not
g62369 not n9139 ; n9139_not
g62370 not n9652 ; n9652_not
g62371 not n7069 ; n7069_not
g62372 not n9805 ; n9805_not
g62373 not n2686 ; n2686_not
g62374 not n6637 ; n6637_not
g62375 not n9094 ; n9094_not
g62376 not n1975 ; n1975_not
g62377 not n7096 ; n7096_not
g62378 not n8527 ; n8527_not
g62379 not n8626 ; n8626_not
g62380 not n8770 ; n8770_not
g62381 not n1687 ; n1687_not
g62382 not n1984 ; n1984_not
g62383 not n1777 ; n1777_not
g62384 not n7456 ; n7456_not
g62385 not n9904 ; n9904_not
g62386 not n9346 ; n9346_not
g62387 not n9436 ; n9436_not
g62388 not n9508 ; n9508_not
g62389 not n9049 ; n9049_not
g62390 not n6970 ; n6970_not
g62391 not n8734 ; n8734_not
g62392 not n1957 ; n1957_not
g62393 not n8761 ; n8761_not
g62394 not n9670 ; n9670_not
g62395 not n7429 ; n7429_not
g62396 not n7573 ; n7573_not
g62397 not n9355 ; n9355_not
g62398 not n2938 ; n2938_not
g62399 not n6907 ; n6907_not
g62400 not n9085 ; n9085_not
g62401 not n8671 ; n8671_not
g62402 not n1678 ; n1678_not
g62403 not n9913 ; n9913_not
g62404 not n9661 ; n9661_not
g62405 not n8860 ; n8860_not
g62406 not n8617 ; n8617_not
g62407 not n9292 ; n9292_not
g62408 not n2668 ; n2668_not
g62409 not n2299 ; n2299_not
g62410 not n9283 ; n9283_not
g62411 not n2974 ; n2974_not
g62412 not n7465 ; n7465_not
g62413 not n7078 ; n7078_not
g62414 not n6646 ; n6646_not
g62415 not n9418 ; n9418_not
g62416 not n8644 ; n8644_not
g62417 not n9607 ; n9607_not
g62418 not n2578 ; n2578_not
g62419 not n7609 ; n7609_not
g62420 not n9193 ; n9193_not
g62421 not n9616 ; n9616_not
g62422 not n1948 ; n1948_not
g62423 not n2587 ; n2587_not
g62424 not n6871 ; n6871_not
g62425 not n9319 ; n9319_not
g62426 not n6655 ; n6655_not
g62427 not n8716 ; n8716_not
g62428 not n8635 ; n8635_not
g62429 not n6592 ; n6592_not
g62430 not n9571 ; n9571_not
g62431 not n8662 ; n8662_not
g62432 not n1579 ; n1579_not
g62433 not n9481 ; n9481_not
g62434 not n9391 ; n9391_not
g62435 not n2569 ; n2569_not
g62436 not n2488 ; n2488_not
g62437 not n9634 ; n9634_not
g62438 not n8941 ; n8941_not
g62439 not n7591 ; n7591_not
g62440 not n9580 ; n9580_not
g62441 not n9832 ; n9832_not
g62442 not n1399 ; n1399_not
g62443 not n8653 ; n8653_not
g62444 not n8725 ; n8725_not
g62445 not n1993 ; n1993_not
g62446 not n9931 ; n9931_not
g62447 not n7177 ; n7177_not
g62448 not n9463 ; n9463_not
g62449 not n9184 ; n9184_not
g62450 not n9238 ; n9238_not
g62451 not n9625 ; n9625_not
g62452 not n1768 ; n1768_not
g62453 not n6880 ; n6880_not
g62454 not n9274 ; n9274_not
g62455 not n8806 ; n8806_not
g62456 not n9742 ; n9742_not
g62457 not n9058 ; n9058_not
g62458 not n8752 ; n8752_not
g62459 not n1867 ; n1867_not
g62460 not n7555 ; n7555_not
g62461 not n8815 ; n8815_not
g62462 not n9229 ; n9229_not
g62463 not n8833 ; n8833_not
g62464 not n5791 ; n5791_not
g62465 not n1849 ; n1849_not
g62466 not n6943 ; n6943_not
g62467 not n1795 ; n1795_not
g62468 not n2479 ; n2479_not
g62469 not n9076 ; n9076_not
g62470 not n7447 ; n7447_not
g62471 not n9733 ; n9733_not
g62472 not n6961 ; n6961_not
g62473 not n9760 ; n9760_not
g62474 not n8590 ; n8590_not
g62475 not n9256 ; n9256_not
g62476 not n8563 ; n8563_not
g62477 not n8572 ; n8572_not
g62478 not n9445 ; n9445_not
g62479 not n9175 ; n9175_not
g62480 not n2659 ; n2659_not
g62481 not n2695 ; n2695_not
g62482 not n1489 ; n1489_not
g62483 not n7546 ; n7546_not
g62484 not n8707 ; n8707_not
g62485 not n8554 ; n8554_not
g62486 not n8851 ; n8851_not
g62487 not n1858 ; n1858_not
g62488 not n1786 ; n1786_not
g62489 not n9166 ; n9166_not
g62490 not n9751 ; n9751_not
g62491 not n1498 ; n1498_not
g62492 not n9265 ; n9265_not
g62493 not n9247 ; n9247_not
g62494 not n6952 ; n6952_not
g62495 not n1894 ; n1894_not
g62496 not n8608 ; n8608_not
g62497 not n8743 ; n8743_not
g62498 not n8536 ; n8536_not
g62499 not n6925 ; n6925_not
g62500 not n9841 ; n9841_not
g62501 not n8914 ; n8914_not
g62502 not n2497 ; n2497_not
g62503 not n8680 ; n8680_not
g62504 not n1669 ; n1669_not
g62505 not n2893 ; n2893_not
g62506 not n7087 ; n7087_not
g62507 not n1597 ; n1597_not
g62508 not n8950 ; n8950_not
g62509 not n9148 ; n9148_not
g62510 not n7483 ; n7483_not
g62511 not n6916 ; n6916_not
g62512 not n1588 ; n1588_not
g62513 not n2398 ; n2398_not
g62514 not n1876 ; n1876_not
g62515 not n8545 ; n8545_not
g62516 not n8905 ; n8905_not
g62517 not n2866 ; n2866_not
g62518 not n9157 ; n9157_not
g62519 not n9724 ; n9724_not
g62520 not n6934 ; n6934_not
g62521 not n9715 ; n9715_not
g62522 not n1885 ; n1885_not
g62523 not n2875 ; n2875_not
g62524 not n9706 ; n9706_not
g62525 not n6745 ; n6745_not
g62526 not n9328 ; n9328_not
g62527 not n7168 ; n7168_not
g62528 not n9526 ; n9526_not
g62529 not n5395 ; n5395_not
g62530 not n7753 ; n7753_not
g62531 not n5386 ; n5386_not
g62532 not n4099 ; n4099_not
g62533 not n8464 ; n8464_not
g62534 not n9553 ; n9553_not
g62535 not n8455 ; n8455_not
g62536 not n8059 ; n8059_not
g62537 not n7744 ; n7744_not
g62538 not n9364 ; n9364_not
g62539 not n3838 ; n3838_not
g62540 not n7960 ; n7960_not
g62541 not n6079 ; n6079_not
g62542 not n8248 ; n8248_not
g62543 not n7735 ; n7735_not
g62544 not n8446 ; n8446_not
g62545 not n7834 ; n7834_not
g62546 not n6088 ; n6088_not
g62547 not n5449 ; n5449_not
g62548 not n5458 ; n5458_not
g62549 not n4198 ; n4198_not
g62550 not n9535 ; n9535_not
g62551 not n4765 ; n4765_not
g62552 not n8257 ; n8257_not
g62553 not n7852 ; n7852_not
g62554 not n8491 ; n8491_not
g62555 not n4396 ; n4396_not
g62556 not n4567 ; n4567_not
g62557 not n4279 ; n4279_not
g62558 not n6277 ; n6277_not
g62559 not n4288 ; n4288_not
g62560 not n7933 ; n7933_not
g62561 not n7843 ; n7843_not
g62562 not n4378 ; n4378_not
g62563 not n4297 ; n4297_not
g62564 not n4693 ; n4693_not
g62565 not n4369 ; n4369_not
g62566 not n5098 ; n5098_not
g62567 not n6196 ; n6196_not
g62568 not n5656 ; n5656_not
g62569 not n5539 ; n5539_not
g62570 not n3784 ; n3784_not
g62571 not n5584 ; n5584_not
g62572 not n7807 ; n7807_not
g62573 not n6187 ; n6187_not
g62574 not n3793 ; n3793_not
g62575 not n6565 ; n6565_not
g62576 not n6574 ; n6574_not
g62577 not n5773 ; n5773_not
g62578 not n6583 ; n6583_not
g62579 not n9544 ; n9544_not
g62580 not n9562 ; n9562_not
g62581 not n4576 ; n4576_not
g62582 not n6097 ; n6097_not
g62583 not n4756 ; n4756_not
g62584 not n5476 ; n5476_not
g62585 not n7825 ; n7825_not
g62586 not n8239 ; n8239_not
g62587 not n7726 ; n7726_not
g62588 not n8068 ; n8068_not
g62589 not n7474 ; n7474_not
g62590 not n8419 ; n8419_not
g62591 not n5593 ; n5593_not
g62592 not n5494 ; n5494_not
g62593 not n3739 ; n3739_not
g62594 not n3748 ; n3748_not
g62595 not n7816 ; n7816_not
g62596 not n5782 ; n5782_not
g62597 not n3757 ; n3757_not
g62598 not n4738 ; n4738_not
g62599 not n4684 ; n4684_not
g62600 not n8509 ; n8509_not
g62601 not n6259 ; n6259_not
g62602 not n8275 ; n8275_not
g62603 not n4675 ; n4675_not
g62604 not n4666 ; n4666_not
g62605 not n7924 ; n7924_not
g62606 not n4657 ; n4657_not
g62607 not n4648 ; n4648_not
g62608 not n5638 ; n5638_not
g62609 not n4639 ; n4639_not
g62610 not n6286 ; n6286_not
g62611 not n7915 ; n7915_not
g62612 not n4774 ; n4774_not
g62613 not n4549 ; n4549_not
g62614 not n6178 ; n6178_not
g62615 not n5872 ; n5872_not
g62616 not n7618 ; n7618_not
g62617 not n5647 ; n5647_not
g62618 not n8473 ; n8473_not
g62619 not n4828 ; n4828_not
g62620 not n4819 ; n4819_not
g62621 not n4495 ; n4495_not
g62622 not n7780 ; n7780_not
g62623 not n7942 ; n7942_not
g62624 not n5089 ; n5089_not
g62625 not n4783 ; n4783_not
g62626 not n7762 ; n7762_not
g62627 not n4558 ; n4558_not
g62628 not n8266 ; n8266_not
g62629 not n5962 ; n5962_not
g62630 not n8284 ; n8284_not
g62631 not n4189 ; n4189_not
g62632 not n5971 ; n5971_not
g62633 not n5980 ; n5980_not
g62634 not n5629 ; n5629_not
g62635 not n4459 ; n4459_not
g62636 not n7870 ; n7870_not
g62637 not n6295 ; n6295_not
g62638 not n7861 ; n7861_not
g62639 not n4387 ; n4387_not
g62640 not n5953 ; n5953_not
g62641 not n4594 ; n4594_not
g62642 not n5944 ; n5944_not
g62643 not n7771 ; n7771_not
g62644 not n4585 ; n4585_not
g62645 not n5935 ; n5935_not
g62646 not n9409 ; n9409_not
g62647 not n2983 ; n2983_not
g62648 not n2992 ; n2992_not
g62649 not n6781 ; n6781_not
g62650 not n5719 ; n5719_not
g62651 not n5692 ; n5692_not
g62652 not n7690 ; n7690_not
g62653 not n5881 ; n5881_not
g62654 not n5665 ; n5665_not
g62655 not n7681 ; n7681_not
g62656 not n6790 ; n6790_not
g62657 not n7636 ; n7636_not
g62658 not n7672 ; n7672_not
g62659 not n6691 ; n6691_not
g62660 not n8923 ; n8923_not
g62661 not n8365 ; n8365_not
g62662 not n8176 ; n8176_not
g62663 not n9490 ; n9490_not
g62664 not n5863 ; n5863_not
g62665 not n7627 ; n7627_not
g62666 not n5728 ; n5728_not
g62667 not n5467 ; n5467_not
g62668 not n6754 ; n6754_not
g62669 not n3298 ; n3298_not
g62670 not n8194 ; n8194_not
g62671 not n5674 ; n5674_not
g62672 not n7708 ; n7708_not
g62673 not n3289 ; n3289_not
g62674 not n6763 ; n6763_not
g62675 not n8383 ; n8383_not
g62676 not n5683 ; n5683_not
g62677 not n8185 ; n8185_not
g62678 not n6772 ; n6772_not
g62679 not n8338 ; n8338_not
g62680 not n5764 ; n5764_not
g62681 not n5854 ; n5854_not
g62682 not n6844 ; n6844_not
g62683 not n8158 ; n8158_not
g62684 not n8329 ; n8329_not
g62685 not n8149 ; n8149_not
g62686 not n2929 ; n2929_not
g62687 not n6853 ; n6853_not
g62688 not n7654 ; n7654_not
g62689 not n5836 ; n5836_not
g62690 not n7645 ; n7645_not
g62691 not n5809 ; n5809_not
g62692 not n6862 ; n6862_not
g62693 not n5818 ; n5818_not
g62694 not n8356 ; n8356_not
g62695 not n7663 ; n7663_not
g62696 not n6808 ; n6808_not
g62697 not n7564 ; n7564_not
g62698 not n2884 ; n2884_not
g62699 not n6682 ; n6682_not
g62700 not n6817 ; n6817_not
g62701 not n5737 ; n5737_not
g62702 not n5746 ; n5746_not
g62703 not n6826 ; n6826_not
g62704 not n8347 ; n8347_not
g62705 not n5755 ; n5755_not
g62706 not n8167 ; n8167_not
g62707 not n6835 ; n6835_not
g62708 not n3694 ; n3694_not
g62709 not n8428 ; n8428_not
g62710 not n3685 ; n3685_not
g62711 not n3676 ; n3676_not
g62712 not n3667 ; n3667_not
g62713 not n3658 ; n3658_not
g62714 not n3649 ; n3649_not
g62715 not n5575 ; n5575_not
g62716 not n6664 ; n6664_not
g62717 not n3469 ; n3469_not
g62718 not n4729 ; n4729_not
g62719 not n3595 ; n3595_not
g62720 not n7519 ; n7519_not
g62721 not n5908 ; n5908_not
g62722 not n7717 ; n7717_not
g62723 not n3829 ; n3829_not
g62724 not n8374 ; n8374_not
g62725 not n8077 ; n8077_not
g62726 not n3766 ; n3766_not
g62727 not n6619 ; n6619_not
g62728 not n9454 ; n9454_not
g62729 not n5566 ; n5566_not
g62730 not n6709 ; n6709_not
g62731 not n3496 ; n3496_not
g62732 not n3478 ; n3478_not
g62733 not n6727 ; n6727_not
g62734 not n3388 ; n3388_not
g62735 not n5827 ; n5827_not
g62736 not n3379 ; n3379_not
g62737 not n8095 ; n8095_not
g62738 not n3586 ; n3586_not
g62739 not n5917 ; n5917_not
g62740 not n8293 ; n8293_not
g62741 not n3577 ; n3577_not
g62742 not n9922 ; n9922_not
g62743 not n8086 ; n8086_not
g62744 not n3559 ; n3559_not
g62745 not n3568 ; n3568_not
g62746 not n7835 ; n7835_not
g62747 not n8861 ; n8861_not
g62748 not n8780 ; n8780_not
g62749 not n8285 ; n8285_not
g62750 not n7826 ; n7826_not
g62751 not n8294 ; n8294_not
g62752 not n7844 ; n7844_not
g62753 not n9086 ; n9086_not
g62754 not n7853 ; n7853_not
g62755 not n7646 ; n7646_not
g62756 not n9185 ; n9185_not
g62757 not n7718 ; n7718_not
g62758 not n9194 ; n9194_not
g62759 not n9383 ; n9383_not
g62760 not n7970 ; n7970_not
g62761 not n8186 ; n8186_not
g62762 not n7727 ; n7727_not
g62763 not n8195 ; n8195_not
g62764 not n7637 ; n7637_not
g62765 not n9365 ; n9365_not
g62766 not n7736 ; n7736_not
g62767 not n8096 ; n8096_not
g62768 not n9239 ; n9239_not
g62769 not n9356 ; n9356_not
g62770 not n9248 ; n9248_not
g62771 not n7745 ; n7745_not
g62772 not n7673 ; n7673_not
g62773 not n9428 ; n9428_not
g62774 not n7682 ; n7682_not
g62775 not n7358 ; n7358_not
g62776 not n9095 ; n9095_not
g62777 not n7691 ; n7691_not
g62778 not n7448 ; n7448_not
g62779 not n8159 ; n8159_not
g62780 not n7664 ; n7664_not
g62781 not n9149 ; n9149_not
g62782 not n9158 ; n9158_not
g62783 not n8168 ; n8168_not
g62784 not n7709 ; n7709_not
g62785 not n9167 ; n9167_not
g62786 not n7655 ; n7655_not
g62787 not n9176 ; n9176_not
g62788 not n8177 ; n8177_not
g62789 not n8069 ; n8069_not
g62790 not n7943 ; n7943_not
g62791 not n7781 ; n7781_not
g62792 not n7385 ; n7385_not
g62793 not n8834 ; n8834_not
g62794 not n7934 ; n7934_not
g62795 not n8249 ; n8249_not
g62796 not n7790 ; n7790_not
g62797 not n7394 ; n7394_not
g62798 not n8258 ; n8258_not
g62799 not n7178 ; n7178_not
g62800 not n7925 ; n7925_not
g62801 not n8267 ; n8267_not
g62802 not n8807 ; n8807_not
g62803 not n7808 ; n7808_not
g62804 not n8276 ; n8276_not
g62805 not n7817 ; n7817_not
g62806 not n7628 ; n7628_not
g62807 not n8087 ; n8087_not
g62808 not n9257 ; n9257_not
g62809 not n7367 ; n7367_not
g62810 not n7754 ; n7754_not
g62811 not n9266 ; n9266_not
g62812 not n9275 ; n9275_not
g62813 not n7763 ; n7763_not
g62814 not n9338 ; n9338_not
g62815 not n7619 ; n7619_not
g62816 not n8078 ; n8078_not
g62817 not n9284 ; n9284_not
g62818 not n7376 ; n7376_not
g62819 not n9293 ; n9293_not
g62820 not n7772 ; n7772_not
g62821 not n8744 ; n8744_not
g62822 not n8735 ; n8735_not
g62823 not n8726 ; n8726_not
g62824 not n8555 ; n8555_not
g62825 not n7556 ; n7556_not
g62826 not n8717 ; n8717_not
g62827 not n8708 ; n8708_not
g62828 not n8546 ; n8546_not
g62829 not n8537 ; n8537_not
g62830 not n8528 ; n8528_not
g62831 not n8690 ; n8690_not
g62832 not n8906 ; n8906_not
g62833 not n7565 ; n7565_not
g62834 not n8681 ; n8681_not
g62835 not n8915 ; n8915_not
g62836 not n8843 ; n8843_not
g62837 not n7277 ; n7277_not
g62838 not n7538 ; n7538_not
g62839 not n7268 ; n7268_not
g62840 not n7259 ; n7259_not
g62841 not n8573 ; n8573_not
g62842 not n8771 ; n8771_not
g62843 not n8564 ; n8564_not
g62844 not n8762 ; n8762_not
g62845 not n8870 ; n8870_not
g62846 not n7529 ; n7529_not
g62847 not n8753 ; n8753_not
g62848 not n9491 ; n9491_not
g62849 not n8627 ; n8627_not
g62850 not n8618 ; n8618_not
g62851 not n7574 ; n7574_not
g62852 not n8609 ; n8609_not
g62853 not n8951 ; n8951_not
g62854 not n8960 ; n8960_not
g62855 not n8591 ; n8591_not
g62856 not n8582 ; n8582_not
g62857 not n8672 ; n8672_not
g62858 not n9446 ; n9446_not
g62859 not n8663 ; n8663_not
g62860 not n8654 ; n8654_not
g62861 not n8645 ; n8645_not
g62862 not n7196 ; n7196_not
g62863 not n8933 ; n8933_not
g62864 not n7583 ; n7583_not
g62865 not n7187 ; n7187_not
g62866 not n8636 ; n8636_not
g62867 not n8465 ; n8465_not
g62868 not n8483 ; n8483_not
g62869 not n9068 ; n9068_not
g62870 not n9455 ; n9455_not
g62871 not n9059 ; n9059_not
g62872 not n7907 ; n7907_not
g62873 not n7871 ; n7871_not
g62874 not n7862 ; n7862_not
g62875 not n8924 ; n8924_not
g62876 not n9077 ; n9077_not
g62877 not n8348 ; n8348_not
g62878 not n8366 ; n8366_not
g62879 not n8375 ; n8375_not
g62880 not n9464 ; n9464_not
g62881 not n8393 ; n8393_not
g62882 not n8438 ; n8438_not
g62883 not n7952 ; n7952_not
g62884 not n8456 ; n8456_not
g62885 not n7493 ; n7493_not
g62886 not n7349 ; n7349_not
g62887 not n7475 ; n7475_not
g62888 not n7484 ; n7484_not
g62889 not n8384 ; n8384_not
g62890 not n9473 ; n9473_not
g62891 not n7295 ; n7295_not
g62892 not n7286 ; n7286_not
g62893 not n7466 ; n7466_not
g62894 not n8474 ; n8474_not
g62895 not n9509 ; n9509_not
g62896 not n9518 ; n9518_not
g62897 not n8429 ; n8429_not
g62898 not n5279 ; n5279_not
g62899 not n6791 ; n6791_not
g62900 not n5099 ; n5099_not
g62901 not n5288 ; n5288_not
g62902 not n5297 ; n5297_not
g62903 not n6782 ; n6782_not
g62904 not n5369 ; n5369_not
g62905 not n5378 ; n5378_not
g62906 not n9824 ; n9824_not
g62907 not n5387 ; n5387_not
g62908 not n1949 ; n1949_not
g62909 not n1958 ; n1958_not
g62910 not n6773 ; n6773_not
g62911 not n5459 ; n5459_not
g62912 not n6827 ; n6827_not
g62913 not n4928 ; n4928_not
g62914 not n4919 ; n4919_not
g62915 not n4892 ; n4892_not
g62916 not n4883 ; n4883_not
g62917 not n4874 ; n4874_not
g62918 not n2498 ; n2498_not
g62919 not n4865 ; n4865_not
g62920 not n4856 ; n4856_not
g62921 not n6818 ; n6818_not
g62922 not n4847 ; n4847_not
g62923 not n4838 ; n4838_not
g62924 not n5189 ; n5189_not
g62925 not n6809 ; n6809_not
g62926 not n5198 ; n5198_not
g62927 not n2489 ; n2489_not
g62928 not n2399 ; n2399_not
g62929 not n9815 ; n9815_not
g62930 not n6692 ; n6692_not
g62931 not n5477 ; n5477_not
g62932 not n6377 ; n6377_not
g62933 not n5468 ; n5468_not
g62934 not n6386 ; n6386_not
g62935 not n6395 ; n6395_not
g62936 not n1985 ; n1985_not
g62937 not n6674 ; n6674_not
g62938 not n6656 ; n6656_not
g62939 not n6449 ; n6449_not
g62940 not n6647 ; n6647_not
g62941 not n1994 ; n1994_not
g62942 not n6458 ; n6458_not
g62943 not n5783 ; n5783_not
g62944 not n6467 ; n6467_not
g62945 not n5792 ; n5792_not
g62946 not n5774 ; n5774_not
g62947 not n6764 ; n6764_not
g62948 not n5486 ; n5486_not
g62949 not n4829 ; n4829_not
g62950 not n6755 ; n6755_not
g62951 not n5549 ; n5549_not
g62952 not n5558 ; n5558_not
g62953 not n6728 ; n6728_not
g62954 not n6719 ; n6719_not
g62955 not n6359 ; n6359_not
g62956 not n6368 ; n6368_not
g62957 not n9923 ; n9923_not
g62958 not n2786 ; n2786_not
g62959 not n4559 ; n4559_not
g62960 not n4568 ; n4568_not
g62961 not n4766 ; n4766_not
g62962 not n2777 ; n2777_not
g62963 not n2768 ; n2768_not
g62964 not n4577 ; n4577_not
g62965 not n2759 ; n2759_not
g62966 not n2669 ; n2669_not
g62967 not n6881 ; n6881_not
g62968 not n4586 ; n4586_not
g62969 not n4595 ; n4595_not
g62970 not n4937 ; n4937_not
g62971 not n6917 ; n6917_not
g62972 not n4775 ; n4775_not
g62973 not n6908 ; n6908_not
g62974 not n4793 ; n4793_not
g62975 not n4496 ; n4496_not
g62976 not n2795 ; n2795_not
g62977 not n4784 ; n4784_not
g62978 not n6890 ; n6890_not
g62979 not n2579 ; n2579_not
g62980 not n2588 ; n2588_not
g62981 not n4694 ; n4694_not
g62982 not n6845 ; n6845_not
g62983 not n4991 ; n4991_not
g62984 not n4982 ; n4982_not
g62985 not n6836 ; n6836_not
g62986 not n4973 ; n4973_not
g62987 not n4964 ; n4964_not
g62988 not n4955 ; n4955_not
g62989 not n4946 ; n4946_not
g62990 not n4739 ; n4739_not
g62991 not n6872 ; n6872_not
g62992 not n4649 ; n4649_not
g62993 not n4658 ; n4658_not
g62994 not n6863 ; n6863_not
g62995 not n4667 ; n4667_not
g62996 not n2696 ; n2696_not
g62997 not n6854 ; n6854_not
g62998 not n2678 ; n2678_not
g62999 not n6665 ; n6665_not
g63000 not n4676 ; n4676_not
g63001 not n5864 ; n5864_not
g63002 not n5675 ; n5675_not
g63003 not n5684 ; n5684_not
g63004 not n1697 ; n1697_not
g63005 not n5693 ; n5693_not
g63006 not n1598 ; n1598_not
g63007 not n1679 ; n1679_not
g63008 not n6287 ; n6287_not
g63009 not n1589 ; n1589_not
g63010 not n5837 ; n5837_not
g63011 not n5729 ; n5729_not
g63012 not n1688 ; n1688_not
g63013 not n1778 ; n1778_not
g63014 not n5972 ; n5972_not
g63015 not n5981 ; n5981_not
g63016 not n6485 ; n6485_not
g63017 not n9914 ; n9914_not
g63018 not n6476 ; n6476_not
g63019 not n5990 ; n5990_not
g63020 not n5639 ; n5639_not
g63021 not n6584 ; n6584_not
g63022 not n5882 ; n5882_not
g63023 not n5648 ; n5648_not
g63024 not n5873 ; n5873_not
g63025 not n5657 ; n5657_not
g63026 not n5666 ; n5666_not
g63027 not n5945 ; n5945_not
g63028 not n5954 ; n5954_not
g63029 not n9833 ; n9833_not
g63030 not n5963 ; n5963_not
g63031 not n6296 ; n6296_not
g63032 not n9419 ; n9419_not
g63033 not n6179 ; n6179_not
g63034 not n1787 ; n1787_not
g63035 not n6197 ; n6197_not
g63036 not n6098 ; n6098_not
g63037 not n6089 ; n6089_not
g63038 not n6269 ; n6269_not
g63039 not n5828 ; n5828_not
g63040 not n5738 ; n5738_not
g63041 not n5747 ; n5747_not
g63042 not n5819 ; n5819_not
g63043 not n5756 ; n5756_not
g63044 not n5765 ; n5765_not
g63045 not n5936 ; n5936_not
g63046 not n1796 ; n1796_not
g63047 not n6548 ; n6548_not
g63048 not n6557 ; n6557_not
g63049 not n5846 ; n5846_not
g63050 not n6629 ; n6629_not
g63051 not n6494 ; n6494_not
g63052 not n6539 ; n6539_not
g63053 not n5576 ; n5576_not
g63054 not n5567 ; n5567_not
g63055 not n5918 ; n5918_not
g63056 not n9932 ; n9932_not
g63057 not n1499 ; n1499_not
g63058 not n5585 ; n5585_not
g63059 not n5909 ; n5909_not
g63060 not n5594 ; n5594_not
g63061 not n1967 ; n1967_not
g63062 not n5891 ; n5891_not
g63063 not n6566 ; n6566_not
g63064 not n9851 ; n9851_not
g63065 not n9842 ; n9842_not
g63066 not n2993 ; n2993_not
g63067 not n4298 ; n4298_not
g63068 not n4289 ; n4289_not
g63069 not n3866 ; n3866_not
g63070 not n7088 ; n7088_not
g63071 not n2948 ; n2948_not
g63072 not n3794 ; n3794_not
g63073 not n3659 ; n3659_not
g63074 not n3668 ; n3668_not
g63075 not n3992 ; n3992_not
g63076 not n3983 ; n3983_not
g63077 not n3857 ; n3857_not
g63078 not n3677 ; n3677_not
g63079 not n4478 ; n4478_not
g63080 not n6980 ; n6980_not
g63081 not n4469 ; n4469_not
g63082 not n2876 ; n2876_not
g63083 not n2885 ; n2885_not
g63084 not n3839 ; n3839_not
g63085 not n3875 ; n3875_not
g63086 not n4199 ; n4199_not
g63087 not n4388 ; n4388_not
g63088 not n4379 ; n4379_not
g63089 not n2939 ; n2939_not
g63090 not n3587 ; n3587_not
g63091 not n3479 ; n3479_not
g63092 not n3596 ; n3596_not
g63093 not n3749 ; n3749_not
g63094 not n3758 ; n3758_not
g63095 not n3929 ; n3929_not
g63096 not n3893 ; n3893_not
g63097 not n2984 ; n2984_not
g63098 not n3884 ; n3884_not
g63099 not n3776 ; n3776_not
g63100 not n3578 ; n3578_not
g63101 not n3569 ; n3569_not
g63102 not n3848 ; n3848_not
g63103 not n7097 ; n7097_not
g63104 not n3974 ; n3974_not
g63105 not n3686 ; n3686_not
g63106 not n3965 ; n3965_not
g63107 not n3695 ; n3695_not
g63108 not n3956 ; n3956_not
g63109 not n3947 ; n3947_not
g63110 not n2975 ; n2975_not
g63111 not n3938 ; n3938_not
g63112 not n6944 ; n6944_not
g63113 not n6953 ; n6953_not
g63114 not n9941 ; n9941_not
g63115 not n2894 ; n2894_not
g63116 not n9329 ; n9329_not
g63117 not n4685 ; n4685_not
g63118 not n6962 ; n6962_not
g63119 not n9374 ; n9374_not
g63120 not n3398 ; n3398_not
g63121 not n6926 ; n6926_not
g63122 not n6935 ; n6935_not
g63123 not n3767 ; n3767_not
g63124 not n4748 ; n4748_not
g63125 not n3488 ; n3488_not
g63126 not n4397 ; n4397_not
g63127 not n2858 ; n2858_not
g63128 not n2867 ; n2867_not
g63129 not n6971 ; n6971_not
g63130 not n7079 ; n7079_not
g63131 not n4487 ; n4487_not
g63132 not n2849 ; n2849_not
g63133 not n1887 ; n1887_not
g63134 not n7656 ; n7656_not
g63135 not n1959 ; n1959_not
g63136 not n1878 ; n1878_not
g63137 not n5919 ; n5919_not
g63138 not n8394 ; n8394_not
g63139 not n8619 ; n8619_not
g63140 not n2868 ; n2868_not
g63141 not n8088 ; n8088_not
g63142 not n5883 ; n5883_not
g63143 not n3894 ; n3894_not
g63144 not n8376 ; n8376_not
g63145 not n3858 ; n3858_not
g63146 not n8925 ; n8925_not
g63147 not n7665 ; n7665_not
g63148 not n7629 ; n7629_not
g63149 not n8385 ; n8385_not
g63150 not n8727 ; n8727_not
g63151 not n8763 ; n8763_not
g63152 not n8745 ; n8745_not
g63153 not n1977 ; n1977_not
g63154 not n3876 ; n3876_not
g63155 not n7683 ; n7683_not
g63156 not n5874 ; n5874_not
g63157 not n8628 ; n8628_not
g63158 not n3867 ; n3867_not
g63159 not n2886 ; n2886_not
g63160 not n1896 ; n1896_not
g63161 not n8637 ; n8637_not
g63162 not n7674 ; n7674_not
g63163 not n3849 ; n3849_not
g63164 not n5928 ; n5928_not
g63165 not n7638 ; n7638_not
g63166 not n3768 ; n3768_not
g63167 not n7647 ; n7647_not
g63168 not n8736 ; n8736_not
g63169 not n1869 ; n1869_not
g63170 not n8097 ; n8097_not
g63171 not n9771 ; n9771_not
g63172 not n9573 ; n9573_not
g63173 not n8916 ; n8916_not
g63174 not n9339 ; n9339_not
g63175 not n8754 ; n8754_not
g63176 not n3777 ; n3777_not
g63177 not n8079 ; n8079_not
g63178 not n8718 ; n8718_not
g63179 not n9744 ; n9744_not
g63180 not n8646 ; n8646_not
g63181 not n5856 ; n5856_not
g63182 not n8709 ; n8709_not
g63183 not n3885 ; n3885_not
g63184 not n7764 ; n7764_not
g63185 not n9168 ; n9168_not
g63186 not n7755 ; n7755_not
g63187 not n9492 ; n9492_not
g63188 not n8781 ; n8781_not
g63189 not n7746 ; n7746_not
g63190 not n7962 ; n7962_not
g63191 not n5793 ; n5793_not
g63192 not n9636 ; n9636_not
g63193 not n7737 ; n7737_not
g63194 not n1788 ; n1788_not
g63195 not n8790 ; n8790_not
g63196 not n7728 ; n7728_not
g63197 not n7719 ; n7719_not
g63198 not n1689 ; n1689_not
g63199 not n9762 ; n9762_not
g63200 not n7980 ; n7980_not
g63201 not n8808 ; n8808_not
g63202 not n8871 ; n8871_not
g63203 not n3399 ; n3399_not
g63204 not n7809 ; n7809_not
g63205 not n6189 ; n6189_not
g63206 not n3498 ; n3498_not
g63207 not n8880 ; n8880_not
g63208 not n7791 ; n7791_not
g63209 not n7935 ; n7935_not
g63210 not n1797 ; n1797_not
g63211 not n7782 ; n7782_not
g63212 not n8772 ; n8772_not
g63213 not n7944 ; n7944_not
g63214 not n7773 ; n7773_not
g63215 not n3489 ; n3489_not
g63216 not n8853 ; n8853_not
g63217 not n8673 ; n8673_not
g63218 not n2967 ; n2967_not
g63219 not n8664 ; n8664_not
g63220 not n9564 ; n9564_not
g63221 not n9456 ; n9456_not
g63222 not n3759 ; n3759_not
g63223 not n9654 ; n9654_not
g63224 not n5892 ; n5892_not
g63225 not n3786 ; n3786_not
g63226 not n8655 ; n8655_not
g63227 not n9546 ; n9546_not
g63228 not n8835 ; n8835_not
g63229 not n8691 ; n8691_not
g63230 not n1698 ; n1698_not
g63231 not n9159 ; n9159_not
g63232 not n5829 ; n5829_not
g63233 not n7692 ; n7692_not
g63234 not n9591 ; n9591_not
g63235 not n9753 ; n9753_not
g63236 not n9645 ; n9645_not
g63237 not n5838 ; n5838_not
g63238 not n8682 ; n8682_not
g63239 not n5847 ; n5847_not
g63240 not n8349 ; n8349_not
g63241 not n4848 ; n4848_not
g63242 not n3966 ; n3966_not
g63243 not n4839 ; n4839_not
g63244 not n3975 ; n3975_not
g63245 not n8583 ; n8583_not
g63246 not n7890 ; n7890_not
g63247 not n2958 ; n2958_not
g63248 not n8475 ; n8475_not
g63249 not n3984 ; n3984_not
g63250 not n9807 ; n9807_not
g63251 not n3993 ; n3993_not
g63252 not n8574 ; n8574_not
g63253 not n8484 ; n8484_not
g63254 not n9528 ; n9528_not
g63255 not n9366 ; n9366_not
g63256 not n8961 ; n8961_not
g63257 not n9483 ; n9483_not
g63258 not n8358 ; n8358_not
g63259 not n8529 ; n8529_not
g63260 not n8565 ; n8565_not
g63261 not n2895 ; n2895_not
g63262 not n9852 ; n9852_not
g63263 not n4389 ; n4389_not
g63264 not n9384 ; n9384_not
g63265 not n7845 ; n7845_not
g63266 not n8547 ; n8547_not
g63267 not n4938 ; n4938_not
g63268 not n3939 ; n3939_not
g63269 not n8295 ; n8295_not
g63270 not n9465 ; n9465_not
g63271 not n4929 ; n4929_not
g63272 not n7854 ; n7854_not
g63273 not n7908 ; n7908_not
g63274 not n9816 ; n9816_not
g63275 not n9078 ; n9078_not
g63276 not n9726 ; n9726_not
g63277 not n8466 ; n8466_not
g63278 not n3948 ; n3948_not
g63279 not n4893 ; n4893_not
g63280 not n9069 ; n9069_not
g63281 not n4884 ; n4884_not
g63282 not n7863 ; n7863_not
g63283 not n8592 ; n8592_not
g63284 not n4875 ; n4875_not
g63285 not n4866 ; n4866_not
g63286 not n4857 ; n4857_not
g63287 not n5199 ; n5199_not
g63288 not n8538 ; n8538_not
g63289 not n9474 ; n9474_not
g63290 not n9690 ; n9690_not
g63291 not n3957 ; n3957_not
g63292 not n4749 ; n4749_not
g63293 not n4686 ; n4686_not
g63294 not n2769 ; n2769_not
g63295 not n4695 ; n4695_not
g63296 not n2778 ; n2778_not
g63297 not n8448 ; n8448_not
g63298 not n4776 ; n4776_not
g63299 not n2787 ; n2787_not
g63300 not n4785 ; n4785_not
g63301 not n9708 ; n9708_not
g63302 not n4794 ; n4794_not
g63303 not n2796 ; n2796_not
g63304 not n4758 ; n4758_not
g63305 not n8493 ; n8493_not
g63306 not n8556 ; n8556_not
g63307 not n4398 ; n4398_not
g63308 not n4479 ; n4479_not
g63309 not n4992 ; n4992_not
g63310 not n2688 ; n2688_not
g63311 not n2697 ; n2697_not
g63312 not n4488 ; n4488_not
g63313 not n4983 ; n4983_not
g63314 not n8970 ; n8970_not
g63315 not n9717 ; n9717_not
g63316 not n4974 ; n4974_not
g63317 not n4965 ; n4965_not
g63318 not n9375 ; n9375_not
g63319 not n4956 ; n4956_not
g63320 not n4947 ; n4947_not
g63321 not n2679 ; n2679_not
g63322 not n5388 ; n5388_not
g63323 not n9663 ; n9663_not
g63324 not n8169 ; n8169_not
g63325 not n8178 ; n8178_not
g63326 not n5298 ; n5298_not
g63327 not n8187 ; n8187_not
g63328 not n8934 ; n8934_not
g63329 not n5289 ; n5289_not
g63330 not n8196 ; n8196_not
g63331 not n5469 ; n5469_not
g63332 not n5478 ; n5478_not
g63333 not n5487 ; n5487_not
g63334 not n8439 ; n8439_not
g63335 not n1968 ; n1968_not
g63336 not n8943 ; n8943_not
g63337 not n9735 ; n9735_not
g63338 not n1995 ; n1995_not
g63339 not n9843 ; n9843_not
g63340 not n9780 ; n9780_not
g63341 not n5784 ; n5784_not
g63342 not n5379 ; n5379_not
g63343 not n9096 ; n9096_not
g63344 not n8259 ; n8259_not
g63345 not n9924 ; n9924_not
g63346 not n7818 ; n7818_not
g63347 not n9087 ; n9087_not
g63348 not n8268 ; n8268_not
g63349 not n7827 ; n7827_not
g63350 not n8277 ; n8277_not
g63351 not n9681 ; n9681_not
g63352 not n2949 ; n2949_not
g63353 not n7836 ; n7836_not
g63354 not n8286 ; n8286_not
g63355 not n9519 ; n9519_not
g63356 not n9672 ; n9672_not
g63357 not n7953 ; n7953_not
g63358 not n9825 ; n9825_not
g63359 not n9537 ; n9537_not
g63360 not n5559 ; n5559_not
g63361 not n5496 ; n5496_not
g63362 not n9555 ; n9555_not
g63363 not n6738 ; n6738_not
g63364 not n7575 ; n7575_not
g63365 not n6846 ; n6846_not
g63366 not n6666 ; n6666_not
g63367 not n6837 ; n6837_not
g63368 not n6675 ; n6675_not
g63369 not n9285 ; n9285_not
g63370 not n6828 ; n6828_not
g63371 not n7566 ; n7566_not
g63372 not n6819 ; n6819_not
g63373 not n6396 ; n6396_not
g63374 not n6387 ; n6387_not
g63375 not n6378 ; n6378_not
g63376 not n9582 ; n9582_not
g63377 not n6792 ; n6792_not
g63378 not n6486 ; n6486_not
g63379 not n9294 ; n9294_not
g63380 not n6477 ; n6477_not
g63381 not n6891 ; n6891_not
g63382 not n6468 ; n6468_not
g63383 not n7593 ; n7593_not
g63384 not n7179 ; n7179_not
g63385 not n6882 ; n6882_not
g63386 not n6459 ; n6459_not
g63387 not n6873 ; n6873_not
g63388 not n7188 ; n7188_not
g63389 not n9609 ; n9609_not
g63390 not n6864 ; n6864_not
g63391 not n7197 ; n7197_not
g63392 not n7584 ; n7584_not
g63393 not n6657 ; n6657_not
g63394 not n6855 ; n6855_not
g63395 not n9258 ; n9258_not
g63396 not n6639 ; n6639_not
g63397 not n9861 ; n9861_not
g63398 not n6594 ; n6594_not
g63399 not n6567 ; n6567_not
g63400 not n9249 ; n9249_not
g63401 not n7359 ; n7359_not
g63402 not n6585 ; n6585_not
g63403 not n7494 ; n7494_not
g63404 not n7368 ; n7368_not
g63405 not n7485 ; n7485_not
g63406 not n7377 ; n7377_not
g63407 not n6558 ; n6558_not
g63408 not n6549 ; n6549_not
g63409 not n7386 ; n7386_not
g63410 not n7476 ; n7476_not
g63411 not n9618 ; n9618_not
g63412 not n6369 ; n6369_not
g63413 not n9438 ; n9438_not
g63414 not n9276 ; n9276_not
g63415 not n6783 ; n6783_not
g63416 not n7269 ; n7269_not
g63417 not n8844 ; n8844_not
g63418 not n6774 ; n6774_not
g63419 not n7278 ; n7278_not
g63420 not n9267 ; n9267_not
g63421 not n7539 ; n7539_not
g63422 not n6765 ; n6765_not
g63423 not n7287 ; n7287_not
g63424 not n6729 ; n6729_not
g63425 not n6747 ; n6747_not
g63426 not n7296 ; n7296_not
g63427 not n9429 ; n9429_not
g63428 not n6684 ; n6684_not
g63429 not n9177 ; n9177_not
g63430 not n9186 ; n9186_not
g63431 not n9195 ; n9195_not
g63432 not n7449 ; n7449_not
g63433 not n7098 ; n7098_not
g63434 not n7458 ; n7458_not
g63435 not n7089 ; n7089_not
g63436 not n9951 ; n9951_not
g63437 not n9942 ; n9942_not
g63438 not n9627 ; n9627_not
g63439 not n9933 ; n9933_not
g63440 not n7395 ; n7395_not
g63441 not n9393 ; n9393_not
g63442 not n6981 ; n6981_not
g63443 not n6972 ; n6972_not
g63444 not n6963 ; n6963_not
g63445 not n7548 ; n7548_not
g63446 not n6954 ; n6954_not
g63447 not n6945 ; n6945_not
g63448 not n6936 ; n6936_not
g63449 not n6927 ; n6927_not
g63450 not n6918 ; n6918_not
g63451 not n6495 ; n6495_not
g63452 not n6909 ; n6909_not
g63453 not n9834 ; n9834_not
g63454 not n9348 ; n9348_not
g63455 not n6990 ; n6990_not
g63456 not n9906 ; n9906_not
g63457 not n7881 ; n7881_not
g63458 not n6297 ; n6297_not
g63459 not n1599 ; n1599_not
g63460 not n7917 ; n7917_not
g63461 not n6279 ; n6279_not
g63462 not n9943 ; n9943_not
g63463 not n7198 ; n7198_not
g63464 not n2788 ; n2788_not
g63465 not n6487 ; n6487_not
g63466 not n8881 ; n8881_not
g63467 not n9709 ; n9709_not
g63468 not n6739 ; n6739_not
g63469 not n4795 ; n4795_not
g63470 not n5839 ; n5839_not
g63471 not n8476 ; n8476_not
g63472 not n7576 ; n7576_not
g63473 not n6496 ; n6496_not
g63474 not n2797 ; n2797_not
g63475 not n8485 ; n8485_not
g63476 not n7189 ; n7189_not
g63477 not n7648 ; n7648_not
g63478 not n8188 ; n8188_not
g63479 not n9727 ; n9727_not
g63480 not n7846 ; n7846_not
g63481 not n8179 ; n8179_not
g63482 not n2779 ; n2779_not
g63483 not n9547 ; n9547_not
g63484 not n6478 ; n6478_not
g63485 not n9349 ; n9349_not
g63486 not n7657 ; n7657_not
g63487 not n8458 ; n8458_not
g63488 not n9763 ; n9763_not
g63489 not n8980 ; n8980_not
g63490 not n9646 ; n9646_not
g63491 not n4786 ; n4786_not
g63492 not n7585 ; n7585_not
g63493 not n7684 ; n7684_not
g63494 not n4687 ; n4687_not
g63495 not n9628 ; n9628_not
g63496 not n4678 ; n4678_not
g63497 not n4669 ; n4669_not
g63498 not n4597 ; n4597_not
g63499 not n6559 ; n6559_not
g63500 not n9790 ; n9790_not
g63501 not n4588 ; n4588_not
g63502 not n4399 ; n4399_not
g63503 not n7279 ; n7279_not
g63504 not n7864 ; n7864_not
g63505 not n4579 ; n4579_not
g63506 not n2869 ; n2869_not
g63507 not n9574 ; n9574_not
g63508 not n9493 ; n9493_not
g63509 not n7666 ; n7666_not
g63510 not n8098 ; n8098_not
g63511 not n7927 ; n7927_not
g63512 not n9961 ; n9961_not
g63513 not n4768 ; n4768_not
g63514 not n8089 ; n8089_not
g63515 not n9853 ; n9853_not
g63516 not n7855 ; n7855_not
g63517 not n7675 ; n7675_not
g63518 not n9556 ; n9556_not
g63519 not n7558 ; n7558_not
g63520 not n7990 ; n7990_not
g63521 not n4696 ; n4696_not
g63522 not n4885 ; n4885_not
g63523 not n4894 ; n4894_not
g63524 not n6676 ; n6676_not
g63525 not n4939 ; n4939_not
g63526 not n9817 ; n9817_not
g63527 not n9826 ; n9826_not
g63528 not n4948 ; n4948_not
g63529 not n4957 ; n4957_not
g63530 not n4966 ; n4966_not
g63531 not n7639 ; n7639_not
g63532 not n4975 ; n4975_not
g63533 not n4984 ; n4984_not
g63534 not n4858 ; n4858_not
g63535 not n9466 ; n9466_not
g63536 not n9691 ; n9691_not
g63537 not n4849 ; n4849_not
g63538 not n6685 ; n6685_not
g63539 not n9529 ; n9529_not
g63540 not n4867 ; n4867_not
g63541 not n4876 ; n4876_not
g63542 not n9808 ; n9808_not
g63543 not n7882 ; n7882_not
g63544 not n2698 ; n2698_not
g63545 not n5857 ; n5857_not
g63546 not n2689 ; n2689_not
g63547 not n8863 ; n8863_not
g63548 not n9376 ; n9376_not
g63549 not n7459 ; n7459_not
g63550 not n3499 ; n3499_not
g63551 not n5848 ; n5848_not
g63552 not n6469 ; n6469_not
g63553 not n4759 ; n4759_not
g63554 not n7594 ; n7594_not
g63555 not n9475 ; n9475_not
g63556 not n8197 ; n8197_not
g63557 not n8368 ; n8368_not
g63558 not n4993 ; n4993_not
g63559 not n6667 ; n6667_not
g63560 not n8296 ; n8296_not
g63561 not n7837 ; n7837_not
g63562 not n9664 ; n9664_not
g63563 not n8287 ; n8287_not
g63564 not n8386 ; n8386_not
g63565 not n8278 ; n8278_not
g63566 not n8395 ; n8395_not
g63567 not n8269 ; n8269_not
g63568 not n8971 ; n8971_not
g63569 not n9754 ; n9754_not
g63570 not n8827 ; n8827_not
g63571 not n7747 ; n7747_not
g63572 not n7099 ; n7099_not
g63573 not n2896 ; n2896_not
g63574 not n5794 ; n5794_not
g63575 not n7954 ; n7954_not
g63576 not n3769 ; n3769_not
g63577 not n7756 ; n7756_not
g63578 not n9772 ; n9772_not
g63579 not n1798 ; n1798_not
g63580 not n3778 ; n3778_not
g63581 not n9673 ; n9673_not
g63582 not n9619 ; n9619_not
g63583 not n3985 ; n3985_not
g63584 not n8890 ; n8890_not
g63585 not n7396 ; n7396_not
g63586 not n3994 ; n3994_not
g63587 not n9358 ; n9358_not
g63588 not n7792 ; n7792_not
g63589 not n7468 ; n7468_not
g63590 not n9781 ; n9781_not
g63591 not n8953 ; n8953_not
g63592 not n9655 ; n9655_not
g63593 not n7738 ; n7738_not
g63594 not n9916 ; n9916_not
g63595 not n1699 ; n1699_not
g63596 not n9736 ; n9736_not
g63597 not n7819 ; n7819_not
g63598 not n7774 ; n7774_not
g63599 not n3589 ; n3589_not
g63600 not n3688 ; n3688_not
g63601 not n9484 ; n9484_not
g63602 not n6289 ; n6289_not
g63603 not n3598 ; n3598_not
g63604 not n7909 ; n7909_not
g63605 not n7828 ; n7828_not
g63606 not n3697 ; n3697_not
g63607 not n3679 ; n3679_not
g63608 not n7783 ; n7783_not
g63609 not n8908 ; n8908_not
g63610 not n8359 ; n8359_not
g63611 not n7945 ; n7945_not
g63612 not n3787 ; n3787_not
g63613 not n9565 ; n9565_not
g63614 not n6757 ; n6757_not
g63615 not n9745 ; n9745_not
g63616 not n6748 ; n6748_not
g63617 not n8935 ; n8935_not
g63618 not n7765 ; n7765_not
g63619 not n9385 ; n9385_not
g63620 not n9934 ; n9934_not
g63621 not n9439 ; n9439_not
g63622 not n8926 ; n8926_not
g63623 not n9583 ; n9583_not
g63624 not n3796 ; n3796_not
g63625 not n9592 ; n9592_not
g63626 not n3976 ; n3976_not
g63627 not n2959 ; n2959_not
g63628 not n3967 ; n3967_not
g63629 not n2977 ; n2977_not
g63630 not n9637 ; n9637_not
g63631 not n3958 ; n3958_not
g63632 not n3949 ; n3949_not
g63633 not n7972 ; n7972_not
g63634 not n4498 ; n4498_not
g63635 not n4489 ; n4489_not
g63636 not n2878 ; n2878_not
g63637 not n7288 ; n7288_not
g63638 not n7693 ; n7693_not
g63639 not n6595 ; n6595_not
g63640 not n7297 ; n7297_not
g63641 not n9718 ; n9718_not
g63642 not n8494 ; n8494_not
g63643 not n8845 ; n8845_not
g63644 not n6586 ; n6586_not
g63645 not n3886 ; n3886_not
g63646 not n7378 ; n7378_not
g63647 not n3895 ; n3895_not
g63648 not n6199 ; n6199_not
g63649 not n8449 ; n8449_not
g63650 not n2995 ; n2995_not
g63651 not n7729 ; n7729_not
g63652 not n7387 ; n7387_not
g63653 not n9862 ; n9862_not
g63654 not n2986 ; n2986_not
g63655 not n7495 ; n7495_not
g63656 not n3877 ; n3877_not
g63657 not n3868 ; n3868_not
g63658 not n3859 ; n3859_not
g63659 not n7369 ; n7369_not
g63660 not n7486 ; n7486_not
g63661 not n8836 ; n8836_not
g63662 not n9952 ; n9952_not
g63663 not n5596 ; n5596_not
g63664 not n5758 ; n5758_not
g63665 not n9538 ; n9538_not
g63666 not n5767 ; n5767_not
g63667 not n5893 ; n5893_not
g63668 not n5776 ; n5776_not
g63669 not n9682 ; n9682_not
g63670 not n1969 ; n1969_not
g63671 not n5965 ; n5965_not
g63672 not n9907 ; n9907_not
g63673 not n5497 ; n5497_not
g63674 not n1888 ; n1888_not
g63675 not n5866 ; n5866_not
g63676 not n9844 ; n9844_not
g63677 not n7549 ; n7549_not
g63678 not n5749 ; n5749_not
g63679 not n5884 ; n5884_not
g63680 not n5299 ; n5299_not
g63681 not n1897 ; n1897_not
g63682 not n8854 ; n8854_not
g63683 not n5479 ; n5479_not
g63684 not n5488 ; n5488_not
g63685 not n5974 ; n5974_not
g63686 not n5587 ; n5587_not
g63687 not n8944 ; n8944_not
g63688 not n6649 ; n6649_not
g63689 not n5578 ; n5578_not
g63690 not n9394 ; n9394_not
g63691 not n5569 ; n5569_not
g63692 not n1987 ; n1987_not
g63693 not n5983 ; n5983_not
g63694 not n5785 ; n5785_not
g63695 not n5992 ; n5992_not
g63696 not n9448 ; n9448_not
g63697 not n1879 ; n1879_not
g63698 not n1978 ; n1978_not
g63699 not n5668 ; n5668_not
g63700 not n6388 ; n6388_not
g63701 not n5659 ; n5659_not
g63702 not n5956 ; n5956_not
g63703 not n6397 ; n6397_not
g63704 not n5686 ; n5686_not
g63705 not n5677 ; n5677_not
g63706 not n5695 ; n5695_not
g63707 not n6379 ; n6379_not
g63708 not n6694 ; n6694_not
g63709 not n5947 ; n5947_not
g63710 not n9871 ; n9871_not
g63711 not n7918 ; n7918_not
g63712 not n7963 ; n7963_not
g63713 not n5938 ; n5938_not
g63714 not n5678 ; n5678_not
g63715 not n9944 ; n9944_not
g63716 not n3995 ; n3995_not
g63717 not n9674 ; n9674_not
g63718 not n3977 ; n3977_not
g63719 not n8585 ; n8585_not
g63720 not n9683 ; n9683_not
g63721 not n5786 ; n5786_not
g63722 not n6686 ; n6686_not
g63723 not n7883 ; n7883_not
g63724 not n7388 ; n7388_not
g63725 not n8990 ; n8990_not
g63726 not n8594 ; n8594_not
g63727 not n3986 ; n3986_not
g63728 not n6893 ; n6893_not
g63729 not n8675 ; n8675_not
g63730 not n9836 ; n9836_not
g63731 not n2969 ; n2969_not
g63732 not n6884 ; n6884_not
g63733 not n8963 ; n8963_not
g63734 not n9827 ; n9827_not
g63735 not n8666 ; n8666_not
g63736 not n9809 ; n9809_not
g63737 not n6992 ; n6992_not
g63738 not n7892 ; n7892_not
g63739 not n5759 ; n5759_not
g63740 not n6929 ; n6929_not
g63741 not n8891 ; n8891_not
g63742 not n6938 ; n6938_not
g63743 not n3896 ; n3896_not
g63744 not n8639 ; n8639_not
g63745 not n9647 ; n9647_not
g63746 not n6965 ; n6965_not
g63747 not n1979 ; n1979_not
g63748 not n3887 ; n3887_not
g63749 not n3878 ; n3878_not
g63750 not n3869 ; n3869_not
g63751 not n9395 ; n9395_not
g63752 not n9575 ; n9575_not
g63753 not n6398 ; n6398_not
g63754 not n6947 ; n6947_not
g63755 not n9188 ; n9188_not
g63756 not n5696 ; n5696_not
g63757 not n2987 ; n2987_not
g63758 not n6677 ; n6677_not
g63759 not n1988 ; n1988_not
g63760 not n6956 ; n6956_not
g63761 not n8459 ; n8459_not
g63762 not n2978 ; n2978_not
g63763 not n8981 ; n8981_not
g63764 not n2996 ; n2996_not
g63765 not n8657 ; n8657_not
g63766 not n6983 ; n6983_not
g63767 not n7964 ; n7964_not
g63768 not n9548 ; n9548_not
g63769 not n7379 ; n7379_not
g63770 not n3968 ; n3968_not
g63771 not n9908 ; n9908_not
g63772 not n6974 ; n6974_not
g63773 not n7478 ; n7478_not
g63774 not n3959 ; n3959_not
g63775 not n7973 ; n7973_not
g63776 not n5687 ; n5687_not
g63777 not n8648 ; n8648_not
g63778 not n6389 ; n6389_not
g63779 not n5975 ; n5975_not
g63780 not n9485 ; n9485_not
g63781 not n5768 ; n5768_not
g63782 not n7496 ; n7496_not
g63783 not n6659 ; n6659_not
g63784 not n9557 ; n9557_not
g63785 not n7937 ; n7937_not
g63786 not n1889 ; n1889_not
g63787 not n9773 ; n9773_not
g63788 not n8792 ; n8792_not
g63789 not n9638 ; n9638_not
g63790 not n9854 ; n9854_not
g63791 not n3698 ; n3698_not
g63792 not n9179 ; n9179_not
g63793 not n9494 ; n9494_not
g63794 not n3689 ; n3689_not
g63795 not n1898 ; n1898_not
g63796 not n5894 ; n5894_not
g63797 not n8756 ; n8756_not
g63798 not n8855 ; n8855_not
g63799 not n2879 ; n2879_not
g63800 not n8765 ; n8765_not
g63801 not n9386 ; n9386_not
g63802 not n7199 ; n7199_not
g63803 not n3788 ; n3788_not
g63804 not n8774 ; n8774_not
g63805 not n5966 ; n5966_not
g63806 not n3779 ; n3779_not
g63807 not n7397 ; n7397_not
g63808 not n5876 ; n5876_not
g63809 not n8369 ; n8369_not
g63810 not n8783 ; n8783_not
g63811 not n8918 ; n8918_not
g63812 not n9719 ; n9719_not
g63813 not n9791 ; n9791_not
g63814 not n9746 ; n9746_not
g63815 not n8846 ; n8846_not
g63816 not n7919 ; n7919_not
g63817 not n7298 ; n7298_not
g63818 not n9665 ; n9665_not
g63819 not n5939 ; n5939_not
g63820 not n9782 ; n9782_not
g63821 not n9917 ; n9917_not
g63822 not n6497 ; n6497_not
g63823 not n8873 ; n8873_not
g63824 not n5948 ; n5948_not
g63825 not n8864 ; n8864_not
g63826 not n9629 ; n9629_not
g63827 not n8828 ; n8828_not
g63828 not n6578 ; n6578_not
g63829 not n9953 ; n9953_not
g63830 not n3599 ; n3599_not
g63831 not n5957 ; n5957_not
g63832 not n9584 ; n9584_not
g63833 not n7289 ; n7289_not
g63834 not n6857 ; n6857_not
g63835 not n7955 ; n7955_not
g63836 not n9764 ; n9764_not
g63837 not n6848 ; n6848_not
g63838 not n9359 ; n9359_not
g63839 not n6479 ; n6479_not
g63840 not n6839 ; n6839_not
g63841 not n9368 ; n9368_not
g63842 not n6488 ; n6488_not
g63843 not n6794 ; n6794_not
g63844 not n9656 ; n9656_not
g63845 not n6875 ; n6875_not
g63846 not n8684 ; n8684_not
g63847 not n9863 ; n9863_not
g63848 not n6866 ; n6866_not
g63849 not n1997 ; n1997_not
g63850 not n8693 ; n8693_not
g63851 not n8945 ; n8945_not
g63852 not n9566 ; n9566_not
g63853 not n9971 ; n9971_not
g63854 not n8738 ; n8738_not
g63855 not n9926 ; n9926_not
g63856 not n3797 ; n3797_not
g63857 not n5849 ; n5849_not
g63858 not n8747 ; n8747_not
g63859 not n6758 ; n6758_not
g63860 not n6587 ; n6587_not
g63861 not n5858 ; n5858_not
g63862 not n6299 ; n6299_not
g63863 not n6785 ; n6785_not
g63864 not n8936 ; n8936_not
g63865 not n6776 ; n6776_not
g63866 not n6596 ; n6596_not
g63867 not n8396 ; n8396_not
g63868 not n8729 ; n8729_not
g63869 not n6767 ; n6767_not
g63870 not n9755 ; n9755_not
g63871 not n4868 ; n4868_not
g63872 not n7595 ; n7595_not
g63873 not n4877 ; n4877_not
g63874 not n9539 ; n9539_not
g63875 not n4769 ; n4769_not
g63876 not n4886 ; n4886_not
g63877 not n9098 ; n9098_not
g63878 not n9692 ; n9692_not
g63879 not n4895 ; n4895_not
g63880 not n9728 ; n9728_not
g63881 not n9881 ; n9881_not
g63882 not n7928 ; n7928_not
g63883 not n2699 ; n2699_not
g63884 not n9278 ; n9278_not
g63885 not n7586 ; n7586_not
g63886 not n4949 ; n4949_not
g63887 not n9962 ; n9962_not
g63888 not n4958 ; n4958_not
g63889 not n7568 ; n7568_not
g63890 not n8495 ; n8495_not
g63891 not n4778 ; n4778_not
g63892 not n5498 ; n5498_not
g63893 not n8486 ; n8486_not
g63894 not n2798 ; n2798_not
g63895 not n5489 ; n5489_not
g63896 not n4796 ; n4796_not
g63897 not n2789 ; n2789_not
g63898 not n8468 ; n8468_not
g63899 not n5993 ; n5993_not
g63900 not n9593 ; n9593_not
g63901 not n4859 ; n4859_not
g63902 not n4976 ; n4976_not
g63903 not n4967 ; n4967_not
g63904 not n9737 ; n9737_not
g63905 not n9818 ; n9818_not
g63906 not n9872 ; n9872_not
g63907 not n6695 ; n6695_not
g63908 not n8954 ; n8954_not
g63909 not n9287 ; n9287_not
g63910 not n7559 ; n7559_not
g63911 not n9458 ; n9458_not
g63912 not n9449 ; n9449_not
g63913 not n9296 ; n9296_not
g63914 not n9089 ; n9089_not
g63915 not n8909 ; n8909_not
g63916 not n4985 ; n4985_not
g63917 not n4994 ; n4994_not
g63918 not n4688 ; n4688_not
g63919 not n8378 ; n8378_not
g63920 not n5867 ; n5867_not
g63921 not n7469 ; n7469_not
g63922 not n4589 ; n4589_not
g63923 not n8567 ; n8567_not
g63924 not n4598 ; n4598_not
g63925 not n9476 ; n9476_not
g63926 not n9197 ; n9197_not
g63927 not n5588 ; n5588_not
g63928 not n8576 ; n8576_not
g63929 not n8549 ; n8549_not
g63930 not n8558 ; n8558_not
g63931 not n4499 ; n4499_not
g63932 not n7982 ; n7982_not
g63933 not n9269 ; n9269_not
g63934 not n5597 ; n5597_not
g63935 not n2888 ; n2888_not
g63936 not n5984 ; n5984_not
g63937 not n5669 ; n5669_not
g63938 not n5579 ; n5579_not
g63939 not n8865 ; n8865_not
g63940 not n6579 ; n6579_not
g63941 not n8298 ; n8298_not
g63942 not n8784 ; n8784_not
g63943 not n6696 ; n6696_not
g63944 not n7659 ; n7659_not
g63945 not n9189 ; n9189_not
g63946 not n8289 ; n8289_not
g63947 not n5949 ; n5949_not
g63948 not n6849 ; n6849_not
g63949 not n6984 ; n6984_not
g63950 not n4689 ; n4689_not
g63951 not n9396 ; n9396_not
g63952 not n8919 ; n8919_not
g63953 not n8793 ; n8793_not
g63954 not n8199 ; n8199_not
g63955 not n7479 ; n7479_not
g63956 not n5688 ; n5688_not
g63957 not n9459 ; n9459_not
g63958 not n7965 ; n7965_not
g63959 not n5886 ; n5886_not
g63960 not n5877 ; n5877_not
g63961 not n3798 ; n3798_not
g63962 not n6786 ; n6786_not
g63963 not n8379 ; n8379_not
g63964 not n8766 ; n8766_not
g63965 not n8955 ; n8955_not
g63966 not n9918 ; n9918_not
g63967 not n8874 ; n8874_not
g63968 not n5859 ; n5859_not
g63969 not n6795 ; n6795_not
g63970 not n3789 ; n3789_not
g63971 not n5967 ; n5967_not
g63972 not n9828 ; n9828_not
g63973 not n5697 ; n5697_not
g63974 not n6975 ; n6975_not
g63975 not n6993 ; n6993_not
g63976 not n9954 ; n9954_not
g63977 not n8775 ; n8775_not
g63978 not n6939 ; n6939_not
g63979 not n5868 ; n5868_not
g63980 not n6687 ; n6687_not
g63981 not n6948 ; n6948_not
g63982 not n7785 ; n7785_not
g63983 not n8559 ; n8559_not
g63984 not n8388 ; n8388_not
g63985 not n6867 ; n6867_not
g63986 not n5958 ; n5958_not
g63987 not n5679 ; n5679_not
g63988 not n7569 ; n7569_not
g63989 not n8829 ; n8829_not
g63990 not n9936 ; n9936_not
g63991 not n6966 ; n6966_not
g63992 not n8595 ; n8595_not
g63993 not n8964 ; n8964_not
g63994 not n7668 ; n7668_not
g63995 not n9369 ; n9369_not
g63996 not n9288 ; n9288_not
g63997 not n7974 ; n7974_not
g63998 not n9963 ; n9963_not
g63999 not n7929 ; n7929_not
g64000 not n6876 ; n6876_not
g64001 not n8838 ; n8838_not
g64002 not n9873 ; n9873_not
g64003 not n8577 ; n8577_not
g64004 not n8991 ; n8991_not
g64005 not n8856 ; n8856_not
g64006 not n9468 ; n9468_not
g64007 not n6894 ; n6894_not
g64008 not n3699 ; n3699_not
g64009 not n6858 ; n6858_not
g64010 not n1899 ; n1899_not
g64011 not n8586 ; n8586_not
g64012 not n8883 ; n8883_not
g64013 not a[0] ; a[0]_not
g64014 not n8469 ; n8469_not
g64015 not n7893 ; n7893_not
g64016 not n9486 ; n9486_not
g64017 not n9819 ; n9819_not
g64018 not n8568 ; n8568_not
g64019 not n9198 ; n9198_not
g64020 not n7677 ; n7677_not
g64021 not n2979 ; n2979_not
g64022 not n6885 ; n6885_not
g64023 not n7839 ; n7839_not
g64024 not n2898 ; n2898_not
g64025 not n9882 ; n9882_not
g64026 not n7794 ; n7794_not
g64027 not n6957 ; n6957_not
g64028 not n9981 ; n9981_not
g64029 not n8694 ; n8694_not
g64030 not n6768 ; n6768_not
g64031 not n7938 ; n7938_not
g64032 not n5769 ; n5769_not
g64033 not n7866 ; n7866_not
g64034 not n7758 ; n7758_not
g64035 not n5994 ; n5994_not
g64036 not n5589 ; n5589_not
g64037 not n1989 ; n1989_not
g64038 not n5976 ; n5976_not
g64039 not n4779 ; n4779_not
g64040 not n7695 ; n7695_not
g64041 not n4599 ; n4599_not
g64042 not n9837 ; n9837_not
g64043 not n9846 ; n9846_not
g64044 not n6597 ; n6597_not
g64045 not n6777 ; n6777_not
g64046 not n7596 ; n7596_not
g64047 not n9972 ; n9972_not
g64048 not n1998 ; n1998_not
g64049 not n7767 ; n7767_not
g64050 not n7983 ; n7983_not
g64051 not n9891 ; n9891_not
g64052 not n5985 ; n5985_not
g64053 not n2997 ; n2997_not
g64054 not n8667 ; n8667_not
g64055 not n8496 ; n8496_not
g64056 not n7992 ; n7992_not
g64057 not n5787 ; n5787_not
g64058 not n8658 ; n8658_not
g64059 not n9864 ; n9864_not
g64060 not n7857 ; n7857_not
g64061 not n5499 ; n5499_not
g64062 not n8676 ; n8676_not
g64063 not n4698 ; n4698_not
g64064 not n4788 ; n4788_not
g64065 not n7749 ; n7749_not
g64066 not n7578 ; n7578_not
g64067 not n8685 ; n8685_not
g64068 not n8478 ; n8478_not
g64069 not n5778 ; n5778_not
g64070 not n8946 ; n8946_not
g64071 not n5796 ; n5796_not
g64072 not n8649 ; n8649_not
g64073 not n8739 ; n8739_not
g64074 not n9279 ; n9279_not
g64075 not n6759 ; n6759_not
g64076 not n7776 ; n7776_not
g64077 not n7686 ; n7686_not
g64078 not n8757 ; n8757_not
g64079 not n8748 ; n8748_not
g64080 not n2889 ; n2889_not
g64081 not n9909 ; n9909_not
g64082 not n2988 ; n2988_not
g64083 not n8973 ; n8973_not
g64084 not n5598 ; n5598_not
g64085 not n8928 ; n8928_not
g64086 not n7848 ; n7848_not
g64087 not n7947 ; n7947_not
g64088 not n9378 ; n9378_not
g64089 not n9927 ; n9927_not
g64090 not n9099 ; n9099_not
g64091 not n7488 ; n7488_not
g64092 not n6669 ; n6669_not
g64093 not n1999 ; n1999_not
g64094 not n9928 ; n9928_not
g64095 not n8839 ; n8839_not
g64096 not n9838 ; n9838_not
g64097 not n8965 ; n8965_not
g64098 not n8875 ; n8875_not
g64099 not n9388 ; n9388_not
g64100 not n9757 ; n9757_not
g64101 not n8956 ; n8956_not
g64102 not n9784 ; n9784_not
g64103 not n8974 ; n8974_not
g64104 not n9946 ; n9946_not
g64105 not n9766 ; n9766_not
g64106 not n9883 ; n9883_not
g64107 not n9919 ; n9919_not
g64108 not n9856 ; n9856_not
g64109 not n9847 ; n9847_not
g64110 not n8938 ; n8938_not
g64111 not n8983 ; n8983_not
g64112 not n2899 ; n2899_not
g64113 not n9874 ; n9874_not
g64114 not n9289 ; n9289_not
g64115 not n9829 ; n9829_not
g64116 not n9199 ; n9199_not
g64117 not n9964 ; n9964_not
g64118 not n9478 ; n9478_not
g64119 not n9775 ; n9775_not
g64120 not n8884 ; n8884_not
g64121 not n8893 ; n8893_not
g64122 not n9937 ; n9937_not
g64123 not n8929 ; n8929_not
g64124 not n8866 ; n8866_not
g64125 not n9793 ; n9793_not
g64126 not n8677 ; n8677_not
g64127 not n6994 ; n6994_not
g64128 not n3997 ; n3997_not
g64129 not n5887 ; n5887_not
g64130 not n5878 ; n5878_not
g64131 not n5869 ; n5869_not
g64132 not n9649 ; n9649_not
g64133 not n8668 ; n8668_not
g64134 not n8659 ; n8659_not
g64135 not n7984 ; n7984_not
g64136 not n7975 ; n7975_not
g64137 not a[1] ; a[1]_not
g64138 not n9973 ; n9973_not
g64139 not n8299 ; n8299_not
g64140 not n7957 ; n7957_not
g64141 not n7588 ; n7588_not
g64142 not n5797 ; n5797_not
g64143 not n9685 ; n9685_not
g64144 not n7939 ; n7939_not
g64145 not n7579 ; n7579_not
g64146 not n8596 ; n8596_not
g64147 not n3889 ; n3889_not
g64148 not n3898 ; n3898_not
g64149 not n6886 ; n6886_not
g64150 not n6895 ; n6895_not
g64151 not n9496 ; n9496_not
g64152 not n6949 ; n6949_not
g64153 not n9739 ; n9739_not
g64154 not n6958 ; n6958_not
g64155 not n8695 ; n8695_not
g64156 not n6967 ; n6967_not
g64157 not n6976 ; n6976_not
g64158 not n7498 ; n7498_not
g64159 not n3979 ; n3979_not
g64160 not n8686 ; n8686_not
g64161 not n6985 ; n6985_not
g64162 not n3988 ; n3988_not
g64163 not n8488 ; n8488_not
g64164 not n4798 ; n4798_not
g64165 not n9694 ; n9694_not
g64166 not n6589 ; n6589_not
g64167 not n7786 ; n7786_not
g64168 not n4789 ; n4789_not
g64169 not n4699 ; n4699_not
g64170 not n7489 ; n7489_not
g64171 not n4879 ; n4879_not
g64172 not n7795 ; n7795_not
g64173 not n4888 ; n4888_not
g64174 not n7849 ; n7849_not
g64175 not n4897 ; n4897_not
g64176 not n4996 ; n4996_not
g64177 not n9892 ; n9892_not
g64178 not n8398 ; n8398_not
g64179 not n9559 ; n9559_not
g64180 not n4987 ; n4987_not
g64181 not n9379 ; n9379_not
g64182 not n4969 ; n4969_not
g64183 not n4978 ; n4978_not
g64184 not n6499 ; n6499_not
g64185 not n9982 ; n9982_not
g64186 not n9577 ; n9577_not
g64187 not n7894 ; n7894_not
g64188 not n7669 ; n7669_not
g64189 not n7678 ; n7678_not
g64190 not n8587 ; n8587_not
g64191 not n8479 ; n8479_not
g64192 not n6697 ; n6697_not
g64193 not n8578 ; n8578_not
g64194 not n7687 ; n7687_not
g64195 not n7696 ; n7696_not
g64196 not n8569 ; n8569_not
g64197 not n7885 ; n7885_not
g64198 not n6679 ; n6679_not
g64199 not n9568 ; n9568_not
g64200 not n7876 ; n7876_not
g64201 not n7759 ; n7759_not
g64202 not n7768 ; n7768_not
g64203 not n7858 ; n7858_not
g64204 not n7777 ; n7777_not
g64205 not n9487 ; n9487_not
g64206 not n6859 ; n6859_not
g64207 not n5698 ; n5698_not
g64208 not n5599 ; n5599_not
g64209 not n5689 ; n5689_not
g64210 not n7399 ; n7399_not
g64211 not n7948 ; n7948_not
g64212 not n6796 ; n6796_not
g64213 not n6787 ; n6787_not
g64214 not n9595 ; n9595_not
g64215 not n6778 ; n6778_not
g64216 not n5896 ; n5896_not
g64217 not n6769 ; n6769_not
g64218 not n9658 ; n9658_not
g64219 not n9469 ; n9469_not
g64220 not n9991 ; n9991_not
g64221 not n9586 ; n9586_not
g64222 not n9667 ; n9667_not
g64223 not n6877 ; n6877_not
g64224 not n8848 ; n8848_not
g64225 not n7993 ; n7993_not
g64226 not n6868 ; n6868_not
g64227 not n8794 ; n8794_not
g64228 not n8758 ; n8758_not
g64229 not n9748 ; n9748_not
g64230 not n8785 ; n8785_not
g64231 not n8767 ; n8767_not
g64232 not n3799 ; n3799_not
g64233 not n8776 ; n8776_not
g64234 not n8389 ; n8389_not
g64235 not n8749 ; n8749_not
g64236 not n9676 ; n9676_not
g64237 not b[1] ; b[1]_not
g64238 not n5789 ; n5789_not
g64239 not n7859 ; n7859_not
g64240 not n5798 ; n5798_not
g64241 not n7877 ; n7877_not
g64242 not n5888 ; n5888_not
g64243 not n5978 ; n5978_not
g64244 not n7985 ; n7985_not
g64245 not n8876 ; n8876_not
g64246 not n9839 ; n9839_not
g64247 not n5897 ; n5897_not
g64248 not n5879 ; n5879_not
g64249 not n7895 ; n7895_not
g64250 not n5969 ; n5969_not
g64251 not n5987 ; n5987_not
g64252 not n5996 ; n5996_not
g64253 not n7949 ; n7949_not
g64254 not n7994 ; n7994_not
g64255 not n7967 ; n7967_not
g64256 not n9659 ; n9659_not
g64257 not n8885 ; n8885_not
g64258 not n7886 ; n7886_not
g64259 not n9893 ; n9893_not
g64260 not n8894 ; n8894_not
g64261 not n9884 ; n9884_not
g64262 not n9947 ; n9947_not
g64263 not n9299 ; n9299_not
g64264 not n9938 ; n9938_not
g64265 not n9587 ; n9587_not
g64266 not n9929 ; n9929_not
g64267 not n9398 ; n9398_not
g64268 not n9596 ; n9596_not
g64269 not n6689 ; n6689_not
g64270 not n6599 ; n6599_not
g64271 not n7769 ; n7769_not
g64272 not n7499 ; n7499_not
g64273 not n7778 ; n7778_not
g64274 not n7787 ; n7787_not
g64275 not n7796 ; n7796_not
g64276 not n9983 ; n9983_not
g64277 not n9848 ; n9848_not
g64278 not n7598 ; n7598_not
g64279 not n7589 ; n7589_not
g64280 not n9578 ; n9578_not
g64281 not n7679 ; n7679_not
g64282 not n7688 ; n7688_not
g64283 not n7697 ; n7697_not
g64284 not n9866 ; n9866_not
g64285 not n8849 ; n8849_not
g64286 not n9569 ; n9569_not
g64287 not n8966 ; n8966_not
g64288 not n9695 ; n9695_not
g64289 not n9749 ; n9749_not
g64290 not n4997 ; n4997_not
g64291 not n8399 ; n8399_not
g64292 not n3899 ; n3899_not
g64293 not n9776 ; n9776_not
g64294 not n4988 ; n4988_not
g64295 not n8948 ; n8948_not
g64296 not n4979 ; n4979_not
g64297 not n3989 ; n3989_not
g64298 not n3998 ; n3998_not
g64299 not n8975 ; n8975_not
g64300 not n9956 ; n9956_not
g64301 not n9767 ; n9767_not
g64302 not n2999 ; n2999_not
g64303 not n8489 ; n8489_not
g64304 not n9479 ; n9479_not
g64305 not n8993 ; n8993_not
g64306 not n4898 ; n4898_not
g64307 not n4889 ; n4889_not
g64308 not n9794 ; n9794_not
g64309 not n8984 ; n8984_not
g64310 not n4799 ; n4799_not
g64311 not n8498 ; n8498_not
g64312 not n9785 ; n9785_not
g64313 not n8939 ; n8939_not
g64314 not n7958 ; n7958_not
g64315 not a[2] ; a[2]_not
g64316 not n9974 ; n9974_not
g64317 not n9389 ; n9389_not
g64318 not n8858 ; n8858_not
g64319 not n9677 ; n9677_not
g64320 not n9758 ; n9758_not
g64321 not n9992 ; n9992_not
g64322 not n9686 ; n9686_not
g64323 not n9857 ; n9857_not
g64324 not n9668 ; n9668_not
g64325 not b[2] ; b[2]_not
g64326 not n6969 ; n6969_not
g64327 not n6978 ; n6978_not
g64328 not n9894 ; n9894_not
g64329 not n8769 ; n8769_not
g64330 not n6987 ; n6987_not
g64331 not n8598 ; n8598_not
g64332 not n8985 ; n8985_not
g64333 not n9876 ; n9876_not
g64334 not n9948 ; n9948_not
g64335 not n9579 ; n9579_not
g64336 not n6879 ; n6879_not
g64337 not n9786 ; n9786_not
g64338 not n8976 ; n8976_not
g64339 not n8868 ; n8868_not
g64340 not n6888 ; n6888_not
g64341 not n9939 ; n9939_not
g64342 not n9993 ; n9993_not
g64343 not n6897 ; n6897_not
g64344 not n9588 ; n9588_not
g64345 not n8895 ; n8895_not
g64346 not n9489 ; n9489_not
g64347 not n8778 ; n8778_not
g64348 not n8787 ; n8787_not
g64349 not n8796 ; n8796_not
g64350 not n9768 ; n9768_not
g64351 not n8697 ; n8697_not
g64352 not n8679 ; n8679_not
g64353 not n8688 ; n8688_not
g64354 not n6996 ; n6996_not
g64355 not n8589 ; n8589_not
g64356 not n3999 ; n3999_not
g64357 not n8958 ; n8958_not
g64358 not n9597 ; n9597_not
g64359 not n9759 ; n9759_not
g64360 not n8886 ; n8886_not
g64361 not n9777 ; n9777_not
g64362 not n7887 ; n7887_not
g64363 not n4998 ; n4998_not
g64364 not n5997 ; n5997_not
g64365 not n9678 ; n9678_not
g64366 not n9696 ; n9696_not
g64367 not n5988 ; n5988_not
g64368 not n4899 ; n4899_not
g64369 not n9867 ; n9867_not
g64370 not n5898 ; n5898_not
g64371 not n5979 ; n5979_not
g64372 not n4989 ; n4989_not
g64373 not n5889 ; n5889_not
g64374 not n7599 ; n7599_not
g64375 not n9984 ; n9984_not
g64376 not n9687 ; n9687_not
g64377 not n7977 ; n7977_not
g64378 not n5799 ; n5799_not
g64379 not n9957 ; n9957_not
g64380 not n7959 ; n7959_not
g64381 not n7869 ; n7869_not
g64382 not n9849 ; n9849_not
g64383 not n7995 ; n7995_not
g64384 not n8949 ; n8949_not
g64385 not n9669 ; n9669_not
g64386 not n8994 ; n8994_not
g64387 not n6798 ; n6798_not
g64388 not n6699 ; n6699_not
g64389 not n9399 ; n9399_not
g64390 not n8499 ; n8499_not
g64391 not n7968 ; n7968_not
g64392 not n9858 ; n9858_not
g64393 not n6789 ; n6789_not
g64394 not a[3] ; a[3]_not
g64395 not n9795 ; n9795_not
g64396 not n9966 ; n9966_not
g64397 not n8859 ; n8859_not
g64398 not n9949 ; n9949_not
g64399 not n9499 ; n9499_not
g64400 not n9679 ; n9679_not
g64401 not n9598 ; n9598_not
g64402 not b[3] ; b[3]_not
g64403 not n9778 ; n9778_not
g64404 not n9769 ; n9769_not
g64405 not n9688 ; n9688_not
g64406 not n9859 ; n9859_not
g64407 not n9697 ; n9697_not
g64408 not n9886 ; n9886_not
g64409 not n9868 ; n9868_not
g64410 not n9787 ; n9787_not
g64411 not n8995 ; n8995_not
g64412 not n9589 ; n9589_not
g64413 not n9796 ; n9796_not
g64414 not n5899 ; n5899_not
g64415 not n5998 ; n5998_not
g64416 not n5989 ; n5989_not
g64417 not n9994 ; n9994_not
g64418 not n9877 ; n9877_not
g64419 not n7699 ; n7699_not
g64420 not n7789 ; n7789_not
g64421 not n7798 ; n7798_not
g64422 not n7888 ; n7888_not
g64423 not n7897 ; n7897_not
g64424 not n7969 ; n7969_not
g64425 not n7987 ; n7987_not
g64426 not n7978 ; n7978_not
g64427 not n6799 ; n6799_not
g64428 not n6889 ; n6889_not
g64429 not n6898 ; n6898_not
g64430 not n6979 ; n6979_not
g64431 not n6988 ; n6988_not
g64432 not a[4] ; a[4]_not
g64433 not n9958 ; n9958_not
g64434 not n9967 ; n9967_not
g64435 not n8797 ; n8797_not
g64436 not n9976 ; n9976_not
g64437 not n8986 ; n8986_not
g64438 not n8896 ; n8896_not
g64439 not n8968 ; n8968_not
g64440 not n8779 ; n8779_not
g64441 not n8959 ; n8959_not
g64442 not n8599 ; n8599_not
g64443 not n8689 ; n8689_not
g64444 not n8788 ; n8788_not
g64445 not n8698 ; n8698_not
g64446 not n8869 ; n8869_not
g64447 not n8878 ; n8878_not
g64448 not b[4] ; b[4]_not
g64449 not n5999 ; n5999_not
g64450 not n9878 ; n9878_not
g64451 not n9977 ; n9977_not
g64452 not n8879 ; n8879_not
g64453 not n9887 ; n9887_not
g64454 not n9896 ; n9896_not
g64455 not n8996 ; n8996_not
g64456 not n8798 ; n8798_not
g64457 not n9869 ; n9869_not
g64458 not n8789 ; n8789_not
g64459 not n8888 ; n8888_not
g64460 not n8699 ; n8699_not
g64461 not n9959 ; n9959_not
g64462 not n8978 ; n8978_not
g64463 not a[5] ; a[5]_not
g64464 not n7799 ; n7799_not
g64465 not n9968 ; n9968_not
g64466 not n9986 ; n9986_not
g64467 not n7979 ; n7979_not
g64468 not n7988 ; n7988_not
g64469 not n8969 ; n8969_not
g64470 not n7997 ; n7997_not
g64471 not n7898 ; n7898_not
g64472 not n7889 ; n7889_not
g64473 not n6989 ; n6989_not
g64474 not n6998 ; n6998_not
g64475 not n6899 ; n6899_not
g64476 not b[5] ; b[5]_not
g64477 not n9798 ; n9798_not
g64478 not n8979 ; n8979_not
g64479 not n8988 ; n8988_not
g64480 not n9789 ; n9789_not
g64481 not n9969 ; n9969_not
g64482 not n9978 ; n9978_not
g64483 not n9888 ; n9888_not
g64484 not n8889 ; n8889_not
g64485 not n9699 ; n9699_not
g64486 not n7989 ; n7989_not
g64487 not n7998 ; n7998_not
g64488 not n7899 ; n7899_not
g64489 not n9897 ; n9897_not
g64490 not a[6] ; a[6]_not
g64491 not n9996 ; n9996_not
g64492 not n8799 ; n8799_not
g64493 not n9987 ; n9987_not
g64494 not n8898 ; n8898_not
g64495 not n9879 ; n9879_not
g64496 not b[6] ; b[6]_not
g64497 not n9898 ; n9898_not
g64498 not n9799 ; n9799_not
g64499 not n9889 ; n9889_not
g64500 not n8899 ; n8899_not
g64501 not n7999 ; n7999_not
g64502 not n9979 ; n9979_not
g64503 not a[7] ; a[7]_not
g64504 not n8998 ; n8998_not
g64505 not n9988 ; n9988_not
g64506 not n9997 ; n9997_not
g64507 not n8989 ; n8989_not
g64508 not b[7] ; b[7]_not
g64509 not n9899 ; n9899_not
g64510 not n9998 ; n9998_not
g64511 not n9989 ; n9989_not
g64512 not a[8] ; a[8]_not
g64513 not n8999 ; n8999_not
g64514 not b[8] ; b[8]_not
g64515 not n9999 ; n9999_not
g64516 not a[9] ; a[9]_not
g64517 not b[9] ; b[9]_not
g64518 not n11000 ; n11000_not
g64519 not n20000 ; n20000_not
g64520 not n10010 ; n10010_not
g64521 not n10001 ; n10001_not
g64522 not n12000 ; n12000_not
g64523 not n10110 ; n10110_not
g64524 not n20100 ; n20100_not
g64525 not n20010 ; n20010_not
g64526 not n10101 ; n10101_not
g64527 not n10020 ; n10020_not
g64528 not n21000 ; n21000_not
g64529 not n11010 ; n11010_not
g64530 not n10002 ; n10002_not
g64531 not n10200 ; n10200_not
g64532 not n30000 ; n30000_not
g64533 not n11100 ; n11100_not
g64534 not n20200 ; n20200_not
g64535 not n10120 ; n10120_not
g64536 not n10210 ; n10210_not
g64537 not n10201 ; n10201_not
g64538 not n10300 ; n10300_not
g64539 not n12100 ; n12100_not
g64540 not n11020 ; n11020_not
g64541 not n11110 ; n11110_not
g64542 not n10030 ; n10030_not
g64543 not n11101 ; n11101_not
g64544 not n20110 ; n20110_not
g64545 not n13000 ; n13000_not
g64546 not n20002 ; n20002_not
g64547 not n11200 ; n11200_not
g64548 not n30100 ; n30100_not
g64549 not n21001 ; n21001_not
g64550 not n10111 ; n10111_not
g64551 not n11002 ; n11002_not
g64552 not n10012 ; n10012_not
g64553 not n12001 ; n12001_not
g64554 not n21010 ; n21010_not
g64555 not n10102 ; n10102_not
g64556 not n10003 ; n10003_not
g64557 not n12010 ; n12010_not
g64558 not n22000 ; n22000_not
g64559 not n20020 ; n20020_not
g64560 not n21100 ; n21100_not
g64561 not n20101 ; n20101_not
g64562 not n10021 ; n10021_not
g64563 not n20021 ; n20021_not
g64564 not n21110 ; n21110_not
g64565 not n13001 ; n13001_not
g64566 not n10202 ; n10202_not
g64567 not n20201 ; n20201_not
g64568 not n10220 ; n10220_not
g64569 not n30200 ; n30200_not
g64570 not n10400 ; n10400_not
g64571 not n21101 ; n21101_not
g64572 not n11300 ; n11300_not
g64573 not n10004 ; n10004_not
g64574 not n20030 ; n20030_not
g64575 not n10301 ; n10301_not
g64576 not n10310 ; n10310_not
g64577 not n12101 ; n12101_not
g64578 not n11201 ; n11201_not
g64579 not n30110 ; n30110_not
g64580 not n10211 ; n10211_not
g64581 not n11210 ; n11210_not
g64582 not n21020 ; n21020_not
g64583 not n20120 ; n20120_not
g64584 not n40100 ; n40100_not
g64585 not n12110 ; n12110_not
g64586 not n32000 ; n32000_not
g64587 not n11003 ; n11003_not
g64588 not n13100 ; n13100_not
g64589 not n12020 ; n12020_not
g64590 not n41000 ; n41000_not
g64591 not n30002 ; n30002_not
g64592 not n12002 ; n12002_not
g64593 not n30011 ; n30011_not
g64594 not n30020 ; n30020_not
g64595 not n20003 ; n20003_not
g64596 not n21011 ; n21011_not
g64597 not n21002 ; n21002_not
g64598 not n11012 ; n11012_not
g64599 not n31100 ; n31100_not
g64600 not n30101 ; n30101_not
g64601 not n11030 ; n11030_not
g64602 not n20300 ; n20300_not
g64603 not n10022 ; n10022_not
g64604 not n13010 ; n13010_not
g64605 not n40001 ; n40001_not
g64606 not n10112 ; n10112_not
g64607 not n10040 ; n10040_not
g64608 not n10121 ; n10121_not
g64609 not n11120 ; n11120_not
g64610 not n10013 ; n10013_not
g64611 not n10103 ; n10103_not
g64612 not n20111 ; n20111_not
g64613 not n40010 ; n40010_not
g64614 not n20102 ; n20102_not
g64615 not n10031 ; n10031_not
g64616 not n21200 ; n21200_not
g64617 not n11102 ; n11102_not
g64618 not n10130 ; n10130_not
g64619 not n12011 ; n12011_not
g64620 not n20012 ; n20012_not
g64621 not n11111 ; n11111_not
g64622 not n20210 ; n20210_not
g64623 not n22001 ; n22001_not
g64624 not n22100 ; n22100_not
g64625 not n10311 ; n10311_not
g64626 not n31101 ; n31101_not
g64627 not n30111 ; n30111_not
g64628 not n31002 ; n31002_not
g64629 not n22002 ; n22002_not
g64630 not n21300 ; n21300_not
g64631 not n40002 ; n40002_not
g64632 not n20400 ; n20400_not
g64633 not n22101 ; n22101_not
g64634 not n50100 ; n50100_not
g64635 not n10320 ; n10320_not
g64636 not n30012 ; n30012_not
g64637 not n31011 ; n31011_not
g64638 not n14100 ; n14100_not
g64639 not n31110 ; n31110_not
g64640 not n30021 ; n30021_not
g64641 not n40020 ; n40020_not
g64642 not n30003 ; n30003_not
g64643 not n40011 ; n40011_not
g64644 not n14010 ; n14010_not
g64645 not n30030 ; n30030_not
g64646 not n40110 ; n40110_not
g64647 not n14001 ; n14001_not
g64648 not n12003 ; n12003_not
g64649 not n10140 ; n10140_not
g64650 not n21003 ; n21003_not
g64651 not n13101 ; n13101_not
g64652 not n41100 ; n41100_not
g64653 not n12012 ; n12012_not
g64654 not n13020 ; n13020_not
g64655 not n13110 ; n13110_not
g64656 not n12021 ; n12021_not
g64657 not n40200 ; n40200_not
g64658 not n10410 ; n10410_not
g64659 not n10401 ; n10401_not
g64660 not n22200 ; n22200_not
g64661 not n12102 ; n12102_not
g64662 not n30120 ; n30120_not
g64663 not n10203 ; n10203_not
g64664 not n13011 ; n13011_not
g64665 not n12111 ; n12111_not
g64666 not n10050 ; n10050_not
g64667 not n10041 ; n10041_not
g64668 not n20211 ; n20211_not
g64669 not n10032 ; n10032_not
g64670 not n10023 ; n10023_not
g64671 not n21120 ; n21120_not
g64672 not n10014 ; n10014_not
g64673 not n22110 ; n22110_not
g64674 not n21111 ; n21111_not
g64675 not n10104 ; n10104_not
g64676 not n21102 ; n21102_not
g64677 not n10500 ; n10500_not
g64678 not n24000 ; n24000_not
g64679 not n20220 ; n20220_not
g64680 not n10113 ; n10113_not
g64681 not n21030 ; n21030_not
g64682 not n21021 ; n21021_not
g64683 not n10122 ; n10122_not
g64684 not n10131 ; n10131_not
g64685 not n21012 ; n21012_not
g64686 not n21210 ; n21210_not
g64687 not n11040 ; n11040_not
g64688 not n20301 ; n20301_not
g64689 not n12120 ; n12120_not
g64690 not n11013 ; n11013_not
g64691 not n11004 ; n11004_not
g64692 not n12300 ; n12300_not
g64693 not n50001 ; n50001_not
g64694 not n20202 ; n20202_not
g64695 not n20310 ; n20310_not
g64696 not n12030 ; n12030_not
g64697 not n10302 ; n10302_not
g64698 not n32010 ; n32010_not
g64699 not n42000 ; n42000_not
g64700 not n10212 ; n10212_not
g64701 not n10221 ; n10221_not
g64702 not n12210 ; n12210_not
g64703 not n10230 ; n10230_not
g64704 not n32100 ; n32100_not
g64705 not n21201 ; n21201_not
g64706 not n50010 ; n50010_not
g64707 not n12201 ; n12201_not
g64708 not n11022 ; n11022_not
g64709 not n32001 ; n32001_not
g64710 not n13002 ; n13002_not
g64711 not n20130 ; n20130_not
g64712 not n15000 ; n15000_not
g64713 not n30210 ; n30210_not
g64714 not n20121 ; n20121_not
g64715 not n20112 ; n20112_not
g64716 not n41001 ; n41001_not
g64717 not n20103 ; n20103_not
g64718 not n41010 ; n41010_not
g64719 not n23001 ; n23001_not
g64720 not n30300 ; n30300_not
g64721 not n20013 ; n20013_not
g64722 not n20040 ; n20040_not
g64723 not n30201 ; n30201_not
g64724 not n20004 ; n20004_not
g64725 not n13200 ; n13200_not
g64726 not n23100 ; n23100_not
g64727 not n50002 ; n50002_not
g64728 not n32011 ; n32011_not
g64729 not n20014 ; n20014_not
g64730 not n12121 ; n12121_not
g64731 not n12112 ; n12112_not
g64732 not n12013 ; n12013_not
g64733 not n30022 ; n30022_not
g64734 not n13201 ; n13201_not
g64735 not n30220 ; n30220_not
g64736 not n12301 ; n12301_not
g64737 not n30121 ; n30121_not
g64738 not n12310 ; n12310_not
g64739 not n42010 ; n42010_not
g64740 not n12103 ; n12103_not
g64741 not n32020 ; n32020_not
g64742 not n40210 ; n40210_not
g64743 not n11014 ; n11014_not
g64744 not n12202 ; n12202_not
g64745 not n11005 ; n11005_not
g64746 not n40012 ; n40012_not
g64747 not n42100 ; n42100_not
g64748 not n20005 ; n20005_not
g64749 not n41101 ; n41101_not
g64750 not n12211 ; n12211_not
g64751 not n40003 ; n40003_not
g64752 not n12220 ; n12220_not
g64753 not n31003 ; n31003_not
g64754 not n10510 ; n10510_not
g64755 not n10501 ; n10501_not
g64756 not n30013 ; n30013_not
g64757 not n42001 ; n42001_not
g64758 not n50020 ; n50020_not
g64759 not n50011 ; n50011_not
g64760 not n30202 ; n30202_not
g64761 not n30400 ; n30400_not
g64762 not n30211 ; n30211_not
g64763 not n50101 ; n50101_not
g64764 not n10402 ; n10402_not
g64765 not n21400 ; n21400_not
g64766 not n25000 ; n25000_not
g64767 not n12400 ; n12400_not
g64768 not n10006 ; n10006_not
g64769 not n41110 ; n41110_not
g64770 not n10411 ; n10411_not
g64771 not n10420 ; n10420_not
g64772 not n30031 ; n30031_not
g64773 not n33001 ; n33001_not
g64774 not n40300 ; n40300_not
g64775 not n22210 ; n22210_not
g64776 not n22030 ; n22030_not
g64777 not n22201 ; n22201_not
g64778 not n12022 ; n12022_not
g64779 not n22111 ; n22111_not
g64780 not n51001 ; n51001_not
g64781 not n30040 ; n30040_not
g64782 not n20023 ; n20023_not
g64783 not n15100 ; n15100_not
g64784 not n22120 ; n22120_not
g64785 not n20500 ; n20500_not
g64786 not n12031 ; n12031_not
g64787 not n13300 ; n13300_not
g64788 not n30103 ; n30103_not
g64789 not n50200 ; n50200_not
g64790 not n40021 ; n40021_not
g64791 not n40120 ; n40120_not
g64792 not n34000 ; n34000_not
g64793 not n40030 ; n40030_not
g64794 not n11410 ; n11410_not
g64795 not n41011 ; n41011_not
g64796 not n11401 ; n11401_not
g64797 not n14020 ; n14020_not
g64798 not n52000 ; n52000_not
g64799 not n14011 ; n14011_not
g64800 not n41002 ; n41002_not
g64801 not n50110 ; n50110_not
g64802 not n14002 ; n14002_not
g64803 not n32101 ; n32101_not
g64804 not n30310 ; n30310_not
g64805 not n22102 ; n22102_not
g64806 not n15010 ; n15010_not
g64807 not n22012 ; n22012_not
g64808 not n14110 ; n14110_not
g64809 not n14101 ; n14101_not
g64810 not n13210 ; n13210_not
g64811 not n23101 ; n23101_not
g64812 not n14200 ; n14200_not
g64813 not n23110 ; n23110_not
g64814 not n31201 ; n31201_not
g64815 not n11500 ; n11500_not
g64816 not n23011 ; n23011_not
g64817 not n21310 ; n21310_not
g64818 not n22300 ; n22300_not
g64819 not n11140 ; n11140_not
g64820 not n11023 ; n11023_not
g64821 not n11131 ; n11131_not
g64822 not n11122 ; n11122_not
g64823 not n11113 ; n11113_not
g64824 not n12130 ; n12130_not
g64825 not n11104 ; n11104_not
g64826 not n31012 ; n31012_not
g64827 not n31021 ; n31021_not
g64828 not n11050 ; n11050_not
g64829 not n31300 ; n31300_not
g64830 not n30004 ; n30004_not
g64831 not n11032 ; n11032_not
g64832 not n30130 ; n30130_not
g64833 not n23200 ; n23200_not
g64834 not n11320 ; n11320_not
g64835 not n11311 ; n11311_not
g64836 not n11302 ; n11302_not
g64837 not n41020 ; n41020_not
g64838 not n23002 ; n23002_not
g64839 not n11230 ; n11230_not
g64840 not n11221 ; n11221_not
g64841 not n12040 ; n12040_not
g64842 not n11212 ; n11212_not
g64843 not n11203 ; n11203_not
g64844 not n41200 ; n41200_not
g64845 not n43000 ; n43000_not
g64846 not n40102 ; n40102_not
g64847 not n34100 ; n34100_not
g64848 not n41210 ; n41210_not
g64849 not n22121 ; n22121_not
g64850 not n20033 ; n20033_not
g64851 not n31004 ; n31004_not
g64852 not n12401 ; n12401_not
g64853 not n11042 ; n11042_not
g64854 not n20204 ; n20204_not
g64855 not n22310 ; n22310_not
g64856 not n41102 ; n41102_not
g64857 not n20303 ; n20303_not
g64858 not n23102 ; n23102_not
g64859 not n20213 ; n20213_not
g64860 not n21005 ; n21005_not
g64861 not n12410 ; n12410_not
g64862 not n30302 ; n30302_not
g64863 not n10610 ; n10610_not
g64864 not n41030 ; n41030_not
g64865 not n14102 ; n14102_not
g64866 not n20402 ; n20402_not
g64867 not n10601 ; n10601_not
g64868 not n11015 ; n11015_not
g64869 not n20042 ; n20042_not
g64870 not n50012 ; n50012_not
g64871 not n41111 ; n41111_not
g64872 not n11024 ; n11024_not
g64873 not n30131 ; n30131_not
g64874 not n22013 ; n22013_not
g64875 not n40022 ; n40022_not
g64876 not n13013 ; n13013_not
g64877 not n11033 ; n11033_not
g64878 not n11123 ; n11123_not
g64879 not n21410 ; n21410_not
g64880 not n12113 ; n12113_not
g64881 not n22004 ; n22004_not
g64882 not n11132 ; n11132_not
g64883 not n12302 ; n12302_not
g64884 not n22301 ; n22301_not
g64885 not n31031 ; n31031_not
g64886 not n11141 ; n11141_not
g64887 not n31130 ; n31130_not
g64888 not n10421 ; n10421_not
g64889 not n51110 ; n51110_not
g64890 not n11150 ; n11150_not
g64891 not n21221 ; n21221_not
g64892 not n14201 ; n14201_not
g64893 not n32102 ; n32102_not
g64894 not n11060 ; n11060_not
g64895 not n41300 ; n41300_not
g64896 not n30032 ; n30032_not
g64897 not n23300 ; n23300_not
g64898 not n13004 ; n13004_not
g64899 not n20114 ; n20114_not
g64900 not n16100 ; n16100_not
g64901 not n32003 ; n32003_not
g64902 not n31022 ; n31022_not
g64903 not n11600 ; n11600_not
g64904 not n12140 ; n12140_not
g64905 not n11105 ; n11105_not
g64906 not n20141 ; n20141_not
g64907 not n13202 ; n13202_not
g64908 not n11114 ; n11114_not
g64909 not n12122 ; n12122_not
g64910 not n42020 ; n42020_not
g64911 not n20231 ; n20231_not
g64912 not n42200 ; n42200_not
g64913 not n32021 ; n32021_not
g64914 not n15200 ; n15200_not
g64915 not n12203 ; n12203_not
g64916 not n10340 ; n10340_not
g64917 not n22220 ; n22220_not
g64918 not n32201 ; n32201_not
g64919 not n50030 ; n50030_not
g64920 not n31202 ; n31202_not
g64921 not n20015 ; n20015_not
g64922 not n21041 ; n21041_not
g64923 not n21212 ; n21212_not
g64924 not n42101 ; n42101_not
g64925 not n32210 ; n32210_not
g64926 not n10313 ; n10313_not
g64927 not n20240 ; n20240_not
g64928 not n30041 ; n30041_not
g64929 not n40112 ; n40112_not
g64930 not n24200 ; n24200_not
g64931 not n22202 ; n22202_not
g64932 not n10151 ; n10151_not
g64933 not n21050 ; n21050_not
g64934 not n21500 ; n21500_not
g64935 not n22211 ; n22211_not
g64936 not n41120 ; n41120_not
g64937 not n13220 ; n13220_not
g64938 not n20330 ; n20330_not
g64939 not n43001 ; n43001_not
g64940 not n52100 ; n52100_not
g64941 not n42110 ; n42110_not
g64942 not n20222 ; n20222_not
g64943 not n50021 ; n50021_not
g64944 not n20150 ; n20150_not
g64945 not n10700 ; n10700_not
g64946 not n26000 ; n26000_not
g64947 not n40220 ; n40220_not
g64948 not n13400 ; n13400_not
g64949 not n21014 ; n21014_not
g64950 not n10160 ; n10160_not
g64951 not n21032 ; n21032_not
g64952 not n22112 ; n22112_not
g64953 not n21320 ; n21320_not
g64954 not n10304 ; n10304_not
g64955 not n32120 ; n32120_not
g64956 not n22031 ; n22031_not
g64957 not n42002 ; n42002_not
g64958 not n14111 ; n14111_not
g64959 not n21023 ; n21023_not
g64960 not n30401 ; n30401_not
g64961 not n51011 ; n51011_not
g64962 not n12131 ; n12131_not
g64963 not n22400 ; n22400_not
g64964 not n43010 ; n43010_not
g64965 not n30023 ; n30023_not
g64966 not n40031 ; n40031_not
g64967 not n14012 ; n14012_not
g64968 not n32300 ; n32300_not
g64969 not n41012 ; n41012_not
g64970 not n13112 ; n13112_not
g64971 not n12221 ; n12221_not
g64972 not n31112 ; n31112_not
g64973 not n10241 ; n10241_not
g64974 not n11402 ; n11402_not
g64975 not n14021 ; n14021_not
g64976 not n20123 ; n20123_not
g64977 not n12320 ; n12320_not
g64978 not n16001 ; n16001_not
g64979 not n50210 ; n50210_not
g64980 not n13121 ; n13121_not
g64981 not n11330 ; n11330_not
g64982 not n52001 ; n52001_not
g64983 not n10232 ; n10232_not
g64984 not n50102 ; n50102_not
g64985 not n23120 ; n23120_not
g64986 not n23021 ; n23021_not
g64987 not n30113 ; n30113_not
g64988 not n31040 ; n31040_not
g64989 not n43100 ; n43100_not
g64990 not n14003 ; n14003_not
g64991 not n20105 ; n20105_not
g64992 not n34010 ; n34010_not
g64993 not n13103 ; n13103_not
g64994 not n14300 ; n14300_not
g64995 not n41021 ; n41021_not
g64996 not n23003 ; n23003_not
g64997 not n31211 ; n31211_not
g64998 not n12311 ; n12311_not
g64999 not n31103 ; n31103_not
g65000 not n16010 ; n16010_not
g65001 not n12230 ; n12230_not
g65002 not n11501 ; n11501_not
g65003 not n30005 ; n30005_not
g65004 not n40130 ; n40130_not
g65005 not n10250 ; n10250_not
g65006 not n30050 ; n30050_not
g65007 not n30014 ; n30014_not
g65008 not n30320 ; n30320_not
g65009 not n11420 ; n11420_not
g65010 not n11510 ; n11510_not
g65011 not n41003 ; n41003_not
g65012 not n13130 ; n13130_not
g65013 not n52010 ; n52010_not
g65014 not n14030 ; n14030_not
g65015 not n21230 ; n21230_not
g65016 not n50120 ; n50120_not
g65017 not n13310 ; n13310_not
g65018 not n20510 ; n20510_not
g65019 not n12050 ; n12050_not
g65020 not n14210 ; n14210_not
g65021 not n10412 ; n10412_not
g65022 not n11213 ; n11213_not
g65023 not n13040 ; n13040_not
g65024 not n11222 ; n11222_not
g65025 not n12032 ; n12032_not
g65026 not n10214 ; n10214_not
g65027 not n11231 ; n11231_not
g65028 not n51101 ; n51101_not
g65029 not n50201 ; n50201_not
g65030 not n12023 ; n12023_not
g65031 not n20411 ; n20411_not
g65032 not n11240 ; n11240_not
g65033 not n20132 ; n20132_not
g65034 not n41201 ; n41201_not
g65035 not n20420 ; n20420_not
g65036 not n13022 ; n13022_not
g65037 not n50003 ; n50003_not
g65038 not n51002 ; n51002_not
g65039 not n20312 ; n20312_not
g65040 not n13031 ; n13031_not
g65041 not n30410 ; n30410_not
g65042 not n30140 ; n30140_not
g65043 not n33200 ; n33200_not
g65044 not n20051 ; n20051_not
g65045 not n10205 ; n10205_not
g65046 not n11204 ; n11204_not
g65047 not n20321 ; n20321_not
g65048 not n10223 ; n10223_not
g65049 not n31121 ; n31121_not
g65050 not n15110 ; n15110_not
g65051 not n20060 ; n20060_not
g65052 not n11303 ; n11303_not
g65053 not n24020 ; n24020_not
g65054 not n23210 ; n23210_not
g65055 not n11312 ; n11312_not
g65056 not n24011 ; n24011_not
g65057 not n12212 ; n12212_not
g65058 not n34001 ; n34001_not
g65059 not n21203 ; n21203_not
g65060 not n11321 ; n11321_not
g65061 not n24002 ; n24002_not
g65062 not n23201 ; n23201_not
g65063 not n23111 ; n23111_not
g65064 not n21302 ; n21302_not
g65065 not n24110 ; n24110_not
g65066 not n12005 ; n12005_not
g65067 not n24101 ; n24101_not
g65068 not n40103 ; n40103_not
g65069 not n23012 ; n23012_not
g65070 not n12500 ; n12500_not
g65071 not n10511 ; n10511_not
g65072 not n33110 ; n33110_not
g65073 not n21113 ; n21113_not
g65074 not n10034 ; n10034_not
g65075 not n10133 ; n10133_not
g65076 not n30500 ; n30500_not
g65077 not n10025 ; n10025_not
g65078 not n22130 ; n22130_not
g65079 not n40004 ; n40004_not
g65080 not n10016 ; n10016_not
g65081 not n10052 ; n10052_not
g65082 not n15020 ; n15020_not
g65083 not n32030 ; n32030_not
g65084 not n10106 ; n10106_not
g65085 not n50300 ; n50300_not
g65086 not n21122 ; n21122_not
g65087 not n21104 ; n21104_not
g65088 not n22040 ; n22040_not
g65089 not n32111 ; n32111_not
g65090 not n21140 ; n21140_not
g65091 not n10043 ; n10043_not
g65092 not n40040 ; n40040_not
g65093 not n51200 ; n51200_not
g65094 not n40202 ; n40202_not
g65095 not n42011 ; n42011_not
g65096 not n33011 ; n33011_not
g65097 not n21131 ; n21131_not
g65098 not n33101 ; n33101_not
g65099 not n10124 ; n10124_not
g65100 not n40013 ; n40013_not
g65101 not n10502 ; n10502_not
g65102 not n12041 ; n12041_not
g65103 not n20024 ; n20024_not
g65104 not n30104 ; n30104_not
g65105 not n10430 ; n10430_not
g65106 not n50111 ; n50111_not
g65107 not n10115 ; n10115_not
g65108 not n13211 ; n13211_not
g65109 not n53000 ; n53000_not
g65110 not n20501 ; n20501_not
g65111 not n10061 ; n10061_not
g65112 not n44000 ; n44000_not
g65113 not n10520 ; n10520_not
g65114 not n10070 ; n10070_not
g65115 not n10142 ; n10142_not
g65116 not n15002 ; n15002_not
g65117 not n20600 ; n20600_not
g65118 not n33002 ; n33002_not
g65119 not n10322 ; n10322_not
g65120 not n13301 ; n13301_not
g65121 not n14120 ; n14120_not
g65122 not n14310 ; n14310_not
g65123 not n24003 ; n24003_not
g65124 not n40140 ; n40140_not
g65125 not n51120 ; n51120_not
g65126 not n22131 ; n22131_not
g65127 not n20700 ; n20700_not
g65128 not n15210 ; n15210_not
g65129 not n11250 ; n11250_not
g65130 not n10611 ; n10611_not
g65131 not n35010 ; n35010_not
g65132 not n23004 ; n23004_not
g65133 not n11232 ; n11232_not
g65134 not n20034 ; n20034_not
g65135 not n10701 ; n10701_not
g65136 not n12015 ; n12015_not
g65137 not n26010 ; n26010_not
g65138 not n31410 ; n31410_not
g65139 not n21060 ; n21060_not
g65140 not n14211 ; n14211_not
g65141 not n22311 ; n22311_not
g65142 not n20007 ; n20007_not
g65143 not n13140 ; n13140_not
g65144 not n14301 ; n14301_not
g65145 not n11241 ; n11241_not
g65146 not n50301 ; n50301_not
g65147 not n20133 ; n20133_not
g65148 not n10215 ; n10215_not
g65149 not n20412 ; n20412_not
g65150 not n13050 ; n13050_not
g65151 not n12006 ; n12006_not
g65152 not n10404 ; n10404_not
g65153 not n10620 ; n10620_not
g65154 not n12222 ; n12222_not
g65155 not n30501 ; n30501_not
g65156 not n20421 ; n20421_not
g65157 not n20124 ; n20124_not
g65158 not n31122 ; n31122_not
g65159 not n10080 ; n10080_not
g65160 not n21204 ; n21204_not
g65161 not n14220 ; n14220_not
g65162 not n11502 ; n11502_not
g65163 not n30123 ; n30123_not
g65164 not n15120 ; n15120_not
g65165 not n10116 ; n10116_not
g65166 not n23112 ; n23112_not
g65167 not n20205 ; n20205_not
g65168 not n16011 ; n16011_not
g65169 not n21240 ; n21240_not
g65170 not n15003 ; n15003_not
g65171 not n26100 ; n26100_not
g65172 not n22032 ; n22032_not
g65173 not n31032 ; n31032_not
g65174 not n10710 ; n10710_not
g65175 not n53001 ; n53001_not
g65176 not n13203 ; n13203_not
g65177 not n23013 ; n23013_not
g65178 not n14040 ; n14040_not
g65179 not n31500 ; n31500_not
g65180 not n13500 ; n13500_not
g65181 not n33102 ; n33102_not
g65182 not n20232 ; n20232_not
g65183 not n43101 ; n43101_not
g65184 not n42003 ; n42003_not
g65185 not n31203 ; n31203_not
g65186 not n31401 ; n31401_not
g65187 not n33201 ; n33201_not
g65188 not n21033 ; n21033_not
g65189 not n20115 ; n20115_not
g65190 not n24210 ; n24210_not
g65191 not n30141 ; n30141_not
g65192 not n12060 ; n12060_not
g65193 not n50130 ; n50130_not
g65194 not n43020 ; n43020_not
g65195 not n20313 ; n20313_not
g65196 not n31050 ; n31050_not
g65197 not n33012 ; n33012_not
g65198 not n20070 ; n20070_not
g65199 not n50202 ; n50202_not
g65200 not n21222 ; n21222_not
g65201 not n13023 ; n13023_not
g65202 not n40410 ; n40410_not
g65203 not n51003 ; n51003_not
g65204 not n32400 ; n32400_not
g65205 not n21024 ; n21024_not
g65206 not n44010 ; n44010_not
g65207 not n22320 ; n22320_not
g65208 not n23031 ; n23031_not
g65209 not n14202 ; n14202_not
g65210 not n25020 ; n25020_not
g65211 not n24012 ; n24012_not
g65212 not n50004 ; n50004_not
g65213 not n34002 ; n34002_not
g65214 not n14400 ; n14400_not
g65215 not n12042 ; n12042_not
g65216 not n16020 ; n16020_not
g65217 not n21051 ; n21051_not
g65218 not n10206 ; n10206_not
g65219 not n21150 ; n21150_not
g65220 not n32112 ; n32112_not
g65221 not n13302 ; n13302_not
g65222 not n13041 ; n13041_not
g65223 not n35100 ; n35100_not
g65224 not n11223 ; n11223_not
g65225 not n12033 ; n12033_not
g65226 not n31104 ; n31104_not
g65227 not n20403 ; n20403_not
g65228 not n22140 ; n22140_not
g65229 not n20610 ; n20610_not
g65230 not n31041 ; n31041_not
g65231 not n51210 ; n51210_not
g65232 not n21141 ; n21141_not
g65233 not n24102 ; n24102_not
g65234 not n13032 ; n13032_not
g65235 not n35001 ; n35001_not
g65236 not n32103 ; n32103_not
g65237 not n21042 ; n21042_not
g65238 not n54000 ; n54000_not
g65239 not n10251 ; n10251_not
g65240 not n11205 ; n11205_not
g65241 not n30231 ; n30231_not
g65242 not n20106 ; n20106_not
g65243 not n10521 ; n10521_not
g65244 not n20052 ; n20052_not
g65245 not n14130 ; n14130_not
g65246 not n21420 ; n21420_not
g65247 not n11214 ; n11214_not
g65248 not n43002 ; n43002_not
g65249 not n11430 ; n11430_not
g65250 not n40104 ; n40104_not
g65251 not n11412 ; n11412_not
g65252 not n50103 ; n50103_not
g65253 not n12510 ; n12510_not
g65254 not n50220 ; n50220_not
g65255 not n10044 ; n10044_not
g65256 not n13104 ; n13104_not
g65257 not n14004 ; n14004_not
g65258 not n11520 ; n11520_not
g65259 not n22014 ; n22014_not
g65260 not n12330 ; n12330_not
g65261 not n10062 ; n10062_not
g65262 not n10107 ; n10107_not
g65263 not n13410 ; n13410_not
g65264 not n10800 ; n10800_not
g65265 not n22401 ; n22401_not
g65266 not n40113 ; n40113_not
g65267 not n20340 ; n20340_not
g65268 not n30600 ; n30600_not
g65269 not n22005 ; n22005_not
g65270 not n21123 ; n21123_not
g65271 not n33300 ; n33300_not
g65272 not n20214 ; n20214_not
g65273 not n12321 ; n12321_not
g65274 not n50112 ; n50112_not
g65275 not n13320 ; n13320_not
g65276 not n25101 ; n25101_not
g65277 not n10053 ; n10053_not
g65278 not n11403 ; n11403_not
g65279 not n21303 ; n21303_not
g65280 not n10512 ; n10512_not
g65281 not n12312 ; n12312_not
g65282 not n20430 ; n20430_not
g65283 not n10242 ; n10242_not
g65284 not n30240 ; n30240_not
g65285 not n14022 ; n14022_not
g65286 not n31221 ; n31221_not
g65287 not n33021 ; n33021_not
g65288 not n21213 ; n21213_not
g65289 not n21132 ; n21132_not
g65290 not n11421 ; n11421_not
g65291 not n12213 ; n12213_not
g65292 not n24300 ; n24300_not
g65293 not n10260 ; n10260_not
g65294 not n15030 ; n15030_not
g65295 not n31113 ; n31113_not
g65296 not n20142 ; n20142_not
g65297 not n44001 ; n44001_not
g65298 not n14013 ; n14013_not
g65299 not n13122 ; n13122_not
g65300 not n25110 ; n25110_not
g65301 not n16002 ; n16002_not
g65302 not n13113 ; n13113_not
g65303 not n31023 ; n31023_not
g65304 not n30105 ; n30105_not
g65305 not n21231 ; n21231_not
g65306 not n23211 ; n23211_not
g65307 not n50040 ; n50040_not
g65308 not n23130 ; n23130_not
g65309 not n10071 ; n10071_not
g65310 not n11304 ; n11304_not
g65311 not n10017 ; n10017_not
g65312 not n27000 ; n27000_not
g65313 not n15012 ; n15012_not
g65314 not n10602 ; n10602_not
g65315 not n20331 ; n20331_not
g65316 not n24111 ; n24111_not
g65317 not n32310 ; n32310_not
g65318 not n23022 ; n23022_not
g65319 not n10224 ; n10224_not
g65320 not n11313 ; n11313_not
g65321 not n20061 ; n20061_not
g65322 not n53010 ; n53010_not
g65323 not n23220 ; n23220_not
g65324 not n25200 ; n25200_not
g65325 not n21402 ; n21402_not
g65326 not n24030 ; n24030_not
g65327 not n30330 ; n30330_not
g65328 not n10008 ; n10008_not
g65329 not n20322 ; n20322_not
g65330 not n12501 ; n12501_not
g65331 not n50031 ; n50031_not
g65332 not n12204 ; n12204_not
g65333 not n22221 ; n22221_not
g65334 not n13401 ; n13401_not
g65335 not n21114 ; n21114_not
g65336 not n11511 ; n11511_not
g65337 not n34020 ; n34020_not
g65338 not n10035 ; n10035_not
g65339 not n11340 ; n11340_not
g65340 not n22122 ; n22122_not
g65341 not n32130 ; n32130_not
g65342 not n20151 ; n20151_not
g65343 not n22212 ; n22212_not
g65344 not n10233 ; n10233_not
g65345 not n23121 ; n23121_not
g65346 not n21105 ; n21105_not
g65347 not n20223 ; n20223_not
g65348 not n20160 ; n20160_not
g65349 not n24021 ; n24021_not
g65350 not n10026 ; n10026_not
g65351 not n40122 ; n40122_not
g65352 not n11322 ; n11322_not
g65353 not n12231 ; n12231_not
g65354 not n12303 ; n12303_not
g65355 not n21330 ; n21330_not
g65356 not n22410 ; n22410_not
g65357 not n23202 ; n23202_not
g65358 not n14031 ; n14031_not
g65359 not n11331 ; n11331_not
g65360 not n14121 ; n14121_not
g65361 not n45000 ; n45000_not
g65362 not n12411 ; n12411_not
g65363 not n50013 ; n50013_not
g65364 not n12141 ; n12141_not
g65365 not n25002 ; n25002_not
g65366 not n12402 ; n12402_not
g65367 not n20520 ; n20520_not
g65368 not n12240 ; n12240_not
g65369 not n51102 ; n51102_not
g65370 not n40230 ; n40230_not
g65371 not n22500 ; n22500_not
g65372 not n11700 ; n11700_not
g65373 not n11601 ; n11601_not
g65374 not n30204 ; n30204_not
g65375 not n33111 ; n33111_not
g65376 not n32220 ; n32220_not
g65377 not n32211 ; n32211_not
g65378 not n32013 ; n32013_not
g65379 not n20025 ; n20025_not
g65380 not n13311 ; n13311_not
g65381 not n43110 ; n43110_not
g65382 not n12132 ; n12132_not
g65383 not n31140 ; n31140_not
g65384 not n20502 ; n20502_not
g65385 not n51300 ; n51300_not
g65386 not n24201 ; n24201_not
g65387 not n32202 ; n32202_not
g65388 not n26001 ; n26001_not
g65389 not n50022 ; n50022_not
g65390 not n31311 ; n31311_not
g65391 not n21600 ; n21600_not
g65392 not n34110 ; n34110_not
g65393 not n21510 ; n21510_not
g65394 not n21006 ; n21006_not
g65395 not n33003 ; n33003_not
g65396 not n34011 ; n34011_not
g65397 not n30510 ; n30510_not
g65398 not n13230 ; n13230_not
g65399 not n20250 ; n20250_not
g65400 not n31320 ; n31320_not
g65401 not n14103 ; n14103_not
g65402 not n21015 ; n21015_not
g65403 not n32121 ; n32121_not
g65404 not n22023 ; n22023_not
g65405 not n12051 ; n12051_not
g65406 not n42030 ; n42030_not
g65407 not n10170 ; n10170_not
g65408 not n22104 ; n22104_not
g65409 not n50211 ; n50211_not
g65410 not n40500 ; n40500_not
g65411 not n20043 ; n20043_not
g65412 not n43011 ; n43011_not
g65413 not n10305 ; n10305_not
g65414 not n42012 ; n42012_not
g65415 not n40320 ; n40320_not
g65416 not n44100 ; n44100_not
g65417 not n40302 ; n40302_not
g65418 not n16200 ; n16200_not
g65419 not n10350 ; n10350_not
g65420 not n31131 ; n31131_not
g65421 not n50121 ; n50121_not
g65422 not n34101 ; n34101_not
g65423 not n40311 ; n40311_not
g65424 not n32040 ; n32040_not
g65425 not n53100 ; n53100_not
g65426 not n12420 ; n12420_not
g65427 not n10152 ; n10152_not
g65428 not n10134 ; n10134_not
g65429 not n41220 ; n41220_not
g65430 not n13212 ; n13212_not
g65431 not n12123 ; n12123_not
g65432 not n23400 ; n23400_not
g65433 not n31212 ; n31212_not
g65434 not n14112 ; n14112_not
g65435 not n10161 ; n10161_not
g65436 not n22230 ; n22230_not
g65437 not n32031 ; n32031_not
g65438 not n10314 ; n10314_not
g65439 not n22050 ; n22050_not
g65440 not n10440 ; n10440_not
g65441 not n11034 ; n11034_not
g65442 not n11115 ; n11115_not
g65443 not n21312 ; n21312_not
g65444 not n51201 ; n51201_not
g65445 not n30150 ; n30150_not
g65446 not n22041 ; n22041_not
g65447 not n11124 ; n11124_not
g65448 not n13014 ; n13014_not
g65449 not n40203 ; n40203_not
g65450 not n51021 ; n51021_not
g65451 not n51111 ; n51111_not
g65452 not n31302 ; n31302_not
g65453 not n17001 ; n17001_not
g65454 not n11043 ; n11043_not
g65455 not n20304 ; n20304_not
g65456 not n11106 ; n11106_not
g65457 not n41301 ; n41301_not
g65458 not n30312 ; n30312_not
g65459 not n11151 ; n11151_not
g65460 not n41310 ; n41310_not
g65461 not n11160 ; n11160_not
g65462 not n22302 ; n22302_not
g65463 not n10125 ; n10125_not
g65464 not n30222 ; n30222_not
g65465 not n11025 ; n11025_not
g65466 not n10143 ; n10143_not
g65467 not n15102 ; n15102_not
g65468 not n11133 ; n11133_not
g65469 not n10422 ; n10422_not
g65470 not n30303 ; n30303_not
g65471 not n24120 ; n24120_not
g65472 not n11142 ; n11142_not
g65473 not n51012 ; n51012_not
g65474 not n12105 ; n12105_not
g65475 not n23310 ; n23310_not
g65476 not n13221 ; n13221_not
g65477 not n20241 ; n20241_not
g65478 not n18000 ; n18000_not
g65479 not n16110 ; n16110_not
g65480 not n32004 ; n32004_not
g65481 not n40401 ; n40401_not
g65482 not n11052 ; n11052_not
g65483 not n11007 ; n11007_not
g65484 not n34200 ; n34200_not
g65485 not n33210 ; n33210_not
g65486 not n50400 ; n50400_not
g65487 not n42021 ; n42021_not
g65488 not n33120 ; n33120_not
g65489 not n50310 ; n50310_not
g65490 not n43200 ; n43200_not
g65491 not n10431 ; n10431_not
g65492 not n30114 ; n30114_not
g65493 not n16101 ; n16101_not
g65494 not n13005 ; n13005_not
g65495 not n12150 ; n12150_not
g65496 not n11610 ; n11610_not
g65497 not n30213 ; n30213_not
g65498 not n41400 ; n41400_not
g65499 not n11061 ; n11061_not
g65500 not n40212 ; n40212_not
g65501 not n23301 ; n23301_not
g65502 not n25011 ; n25011_not
g65503 not n40501 ; n40501_not
g65504 not n50410 ; n50410_not
g65505 not n28000 ; n28000_not
g65506 not n23131 ; n23131_not
g65507 not n22330 ; n22330_not
g65508 not n32410 ; n32410_not
g65509 not n35002 ; n35002_not
g65510 not n22321 ; n22321_not
g65511 not n32122 ; n32122_not
g65512 not n22411 ; n22411_not
g65513 not n40510 ; n40510_not
g65514 not n11701 ; n11701_not
g65515 not n24013 ; n24013_not
g65516 not n23320 ; n23320_not
g65517 not n24103 ; n24103_not
g65518 not n11521 ; n11521_not
g65519 not n35020 ; n35020_not
g65520 not n51121 ; n51121_not
g65521 not n22141 ; n22141_not
g65522 not n35011 ; n35011_not
g65523 not n22402 ; n22402_not
g65524 not n24040 ; n24040_not
g65525 not n41005 ; n41005_not
g65526 not n24022 ; n24022_not
g65527 not n32140 ; n32140_not
g65528 not n23104 ; n23104_not
g65529 not n11710 ; n11710_not
g65530 not n22132 ; n22132_not
g65531 not n30052 ; n30052_not
g65532 not n30034 ; n30034_not
g65533 not n24031 ; n24031_not
g65534 not n23014 ; n23014_not
g65535 not n22114 ; n22114_not
g65536 not n32401 ; n32401_not
g65537 not n22420 ; n22420_not
g65538 not n13222 ; n13222_not
g65539 not n23122 ; n23122_not
g65540 not n23302 ; n23302_not
g65541 not n22060 ; n22060_not
g65542 not n40150 ; n40150_not
g65543 not n32131 ; n32131_not
g65544 not n11503 ; n11503_not
g65545 not n54100 ; n54100_not
g65546 not n30025 ; n30025_not
g65547 not n30340 ; n30340_not
g65548 not n30043 ; n30043_not
g65549 not n24004 ; n24004_not
g65550 not n23311 ; n23311_not
g65551 not n11800 ; n11800_not
g65552 not n13213 ; n13213_not
g65553 not n11512 ; n11512_not
g65554 not n23041 ; n23041_not
g65555 not n30403 ; n30403_not
g65556 not n13240 ; n13240_not
g65557 not n50140 ; n50140_not
g65558 not n23023 ; n23023_not
g65559 not n32500 ; n32500_not
g65560 not n22240 ; n22240_not
g65561 not n43021 ; n43021_not
g65562 not n13321 ; n13321_not
g65563 not n32320 ; n32320_not
g65564 not n50122 ; n50122_not
g65565 not n32221 ; n32221_not
g65566 not n50131 ; n50131_not
g65567 not n51013 ; n51013_not
g65568 not n41122 ; n41122_not
g65569 not n12133 ; n12133_not
g65570 not n13510 ; n13510_not
g65571 not n53101 ; n53101_not
g65572 not n13501 ; n13501_not
g65573 not n34120 ; n34120_not
g65574 not n16120 ; n16120_not
g65575 not n23401 ; n23401_not
g65576 not n16201 ; n16201_not
g65577 not n51130 ; n51130_not
g65578 not n21700 ; n21700_not
g65579 not n22600 ; n22600_not
g65580 not n13600 ; n13600_not
g65581 not n12106 ; n12106_not
g65582 not n13411 ; n13411_not
g65583 not n22222 ; n22222_not
g65584 not n51103 ; n51103_not
g65585 not n13312 ; n13312_not
g65586 not n51004 ; n51004_not
g65587 not n32230 ; n32230_not
g65588 not n45100 ; n45100_not
g65589 not n13402 ; n13402_not
g65590 not n22231 ; n22231_not
g65591 not n13420 ; n13420_not
g65592 not n23410 ; n23410_not
g65593 not n32203 ; n32203_not
g65594 not n50050 ; n50050_not
g65595 not n34210 ; n34210_not
g65596 not n43030 ; n43030_not
g65597 not n16102 ; n16102_not
g65598 not n12160 ; n12160_not
g65599 not n13006 ; n13006_not
g65600 not n50500 ; n50500_not
g65601 not n53110 ; n53110_not
g65602 not n12142 ; n12142_not
g65603 not n31006 ; n31006_not
g65604 not n12151 ; n12151_not
g65605 not n32212 ; n32212_not
g65606 not n41032 ; n41032_not
g65607 not n21610 ; n21610_not
g65608 not n21601 ; n21601_not
g65609 not n30502 ; n30502_not
g65610 not n34201 ; n34201_not
g65611 not n34102 ; n34102_not
g65612 not n31015 ; n31015_not
g65613 not n30520 ; n30520_not
g65614 not n16111 ; n16111_not
g65615 not n22024 ; n22024_not
g65616 not n12007 ; n12007_not
g65617 not n41302 ; n41302_not
g65618 not n12016 ; n12016_not
g65619 not n22042 ; n22042_not
g65620 not n20017 ; n20017_not
g65621 not n41104 ; n41104_not
g65622 not n22150 ; n22150_not
g65623 not n43300 ; n43300_not
g65624 not n53200 ; n53200_not
g65625 not n34021 ; n34021_not
g65626 not n30421 ; n30421_not
g65627 not n23500 ; n23500_not
g65628 not n53002 ; n53002_not
g65629 not n34300 ; n34300_not
g65630 not n30610 ; n30610_not
g65631 not n43111 ; n43111_not
g65632 not n30412 ; n30412_not
g65633 not n30601 ; n30601_not
g65634 not n30511 ; n30511_not
g65635 not n41311 ; n41311_not
g65636 not n53011 ; n53011_not
g65637 not n30430 ; n30430_not
g65638 not n50401 ; n50401_not
g65639 not n43012 ; n43012_not
g65640 not n41113 ; n41113_not
g65641 not n20026 ; n20026_not
g65642 not n13303 ; n13303_not
g65643 not n34111 ; n34111_not
g65644 not n41041 ; n41041_not
g65645 not n12043 ; n12043_not
g65646 not n50113 ; n50113_not
g65647 not n13141 ; n13141_not
g65648 not n43102 ; n43102_not
g65649 not n12601 ; n12601_not
g65650 not n12052 ; n12052_not
g65651 not n43003 ; n43003_not
g65652 not n53020 ; n53020_not
g65653 not n22105 ; n22105_not
g65654 not n12061 ; n12061_not
g65655 not n22006 ; n22006_not
g65656 not n41050 ; n41050_not
g65657 not n34012 ; n34012_not
g65658 not n23203 ; n23203_not
g65659 not n22510 ; n22510_not
g65660 not n13231 ; n13231_not
g65661 not n40105 ; n40105_not
g65662 not n13330 ; n13330_not
g65663 not n23032 ; n23032_not
g65664 not n22501 ; n22501_not
g65665 not n41500 ; n41500_not
g65666 not n34030 ; n34030_not
g65667 not n23212 ; n23212_not
g65668 not n11431 ; n11431_not
g65669 not n40123 ; n40123_not
g65670 not n13132 ; n13132_not
g65671 not n30700 ; n30700_not
g65672 not n30007 ; n30007_not
g65673 not n37000 ; n37000_not
g65674 not n23230 ; n23230_not
g65675 not n23140 ; n23140_not
g65676 not n16300 ; n16300_not
g65677 not n30016 ; n30016_not
g65678 not n13150 ; n13150_not
g65679 not n41401 ; n41401_not
g65680 not n41014 ; n41014_not
g65681 not n13105 ; n13105_not
g65682 not n22051 ; n22051_not
g65683 not n34003 ; n34003_not
g65684 not n13114 ; n13114_not
g65685 not n40114 ; n40114_not
g65686 not n13123 ; n13123_not
g65687 not n23221 ; n23221_not
g65688 not n22204 ; n22204_not
g65689 not n24301 ; n24301_not
g65690 not n41221 ; n41221_not
g65691 not n40600 ; n40600_not
g65692 not n13024 ; n13024_not
g65693 not n12070 ; n12070_not
g65694 not n24220 ; n24220_not
g65695 not n24211 ; n24211_not
g65696 not n51022 ; n51022_not
g65697 not n22303 ; n22303_not
g65698 not n41131 ; n41131_not
g65699 not n12115 ; n12115_not
g65700 not n13015 ; n13015_not
g65701 not n24310 ; n24310_not
g65702 not n20800 ; n20800_not
g65703 not n24130 ; n24130_not
g65704 not n32104 ; n32104_not
g65705 not n16210 ; n16210_not
g65706 not n24121 ; n24121_not
g65707 not n24112 ; n24112_not
g65708 not n13060 ; n13060_not
g65709 not n13033 ; n13033_not
g65710 not n24202 ; n24202_not
g65711 not n41023 ; n41023_not
g65712 not n13042 ; n13042_not
g65713 not n20008 ; n20008_not
g65714 not n51031 ; n51031_not
g65715 not n12025 ; n12025_not
g65716 not n13051 ; n13051_not
g65717 not n20404 ; n20404_not
g65718 not n11071 ; n11071_not
g65719 not n20413 ; n20413_not
g65720 not n20305 ; n20305_not
g65721 not n11062 ; n11062_not
g65722 not n31303 ; n31303_not
g65723 not n20422 ; n20422_not
g65724 not n10540 ; n10540_not
g65725 not n11080 ; n11080_not
g65726 not n40051 ; n40051_not
g65727 not n11053 ; n11053_not
g65728 not n15400 ; n15400_not
g65729 not n40060 ; n40060_not
g65730 not n20431 ; n20431_not
g65731 not n21430 ; n21430_not
g65732 not n10522 ; n10522_not
g65733 not n40402 ; n40402_not
g65734 not n20314 ; n20314_not
g65735 not n41140 ; n41140_not
g65736 not n33112 ; n33112_not
g65737 not n15130 ; n15130_not
g65738 not n32041 ; n32041_not
g65739 not n21016 ; n21016_not
g65740 not n11125 ; n11125_not
g65741 not n33004 ; n33004_not
g65742 not n40006 ; n40006_not
g65743 not n11116 ; n11116_not
g65744 not n21007 ; n21007_not
g65745 not n30151 ; n30151_not
g65746 not n11035 ; n11035_not
g65747 not n32050 ; n32050_not
g65748 not n40015 ; n40015_not
g65749 not n11107 ; n11107_not
g65750 not n15112 ; n15112_not
g65751 not n40024 ; n40024_not
g65752 not n20620 ; n20620_not
g65753 not n11044 ; n11044_not
g65754 not n40033 ; n40033_not
g65755 not n33103 ; n33103_not
g65756 not n31501 ; n31501_not
g65757 not n40042 ; n40042_not
g65758 not n10630 ; n10630_not
g65759 not n20602 ; n20602_not
g65760 not n20530 ; n20530_not
g65761 not n41212 ; n41212_not
g65762 not n10081 ; n10081_not
g65763 not n15022 ; n15022_not
g65764 not n33310 ; n33310_not
g65765 not n20323 ; n20323_not
g65766 not n10090 ; n10090_not
g65767 not n17002 ; n17002_not
g65768 not n31222 ; n31222_not
g65769 not n33022 ; n33022_not
g65770 not n35101 ; n35101_not
g65771 not n31312 ; n31312_not
g65772 not n20332 ; n20332_not
g65773 not n30160 ; n30160_not
g65774 not n10108 ; n10108_not
g65775 not n10117 ; n10117_not
g65776 not n31510 ; n31510_not
g65777 not n10126 ; n10126_not
g65778 not n10135 ; n10135_not
g65779 not n15004 ; n15004_not
g65780 not n10009 ; n10009_not
g65781 not n10018 ; n10018_not
g65782 not n40204 ; n40204_not
g65783 not n10027 ; n10027_not
g65784 not n20440 ; n20440_not
g65785 not n35110 ; n35110_not
g65786 not n10036 ; n10036_not
g65787 not n15040 ; n15040_not
g65788 not n10045 ; n10045_not
g65789 not n40213 ; n40213_not
g65790 not n33013 ; n33013_not
g65791 not n10603 ; n10603_not
g65792 not n11017 ; n11017_not
g65793 not n10612 ; n10612_not
g65794 not n10054 ; n10054_not
g65795 not n10063 ; n10063_not
g65796 not n10621 ; n10621_not
g65797 not n10072 ; n10072_not
g65798 not n11251 ; n11251_not
g65799 not n31042 ; n31042_not
g65800 not n10711 ; n10711_not
g65801 not n11242 ; n11242_not
g65802 not n33130 ; n33130_not
g65803 not n10702 ; n10702_not
g65804 not n21070 ; n21070_not
g65805 not n11233 ; n11233_not
g65806 not n30133 ; n30133_not
g65807 not n11224 ; n11224_not
g65808 not n15220 ; n15220_not
g65809 not n21061 ; n21061_not
g65810 not n40420 ; n40420_not
g65811 not n31051 ; n31051_not
g65812 not n11215 ; n11215_not
g65813 not n20233 ; n20233_not
g65814 not n20206 ; n20206_not
g65815 not n26200 ; n26200_not
g65816 not n20215 ; n20215_not
g65817 not n30304 ; n30304_not
g65818 not n52300 ; n52300_not
g65819 not n31033 ; n31033_not
g65820 not n21106 ; n21106_not
g65821 not n20260 ; n20260_not
g65822 not n25201 ; n25201_not
g65823 not n32005 ; n32005_not
g65824 not n25210 ; n25210_not
g65825 not n20224 ; n20224_not
g65826 not n31024 ; n31024_not
g65827 not n11260 ; n11260_not
g65828 not n42220 ; n42220_not
g65829 not n10720 ; n10720_not
g65830 not n11170 ; n11170_not
g65831 not n20251 ; n20251_not
g65832 not n20341 ; n20341_not
g65833 not n11008 ; n11008_not
g65834 not n42202 ; n42202_not
g65835 not n11161 ; n11161_not
g65836 not n41203 ; n41203_not
g65837 not n11152 ; n11152_not
g65838 not n20350 ; n20350_not
g65839 not n11143 ; n11143_not
g65840 not n21025 ; n21025_not
g65841 not n11134 ; n11134_not
g65842 not n11206 ; n11206_not
g65843 not n21052 ; n21052_not
g65844 not n15202 ; n15202_not
g65845 not n32023 ; n32023_not
g65846 not n31060 ; n31060_not
g65847 not n21043 ; n21043_not
g65848 not n35200 ; n35200_not
g65849 not n20242 ; n20242_not
g65850 not n14401 ; n14401_not
g65851 not n25300 ; n25300_not
g65852 not n42211 ; n42211_not
g65853 not n50311 ; n50311_not
g65854 not n21403 ; n21403_not
g65855 not n40411 ; n40411_not
g65856 not n21034 ; n21034_not
g65857 not n33121 ; n33121_not
g65858 not n17200 ; n17200_not
g65859 not n21340 ; n21340_not
g65860 not n42013 ; n42013_not
g65861 not n20503 ; n20503_not
g65862 not n21133 ; n21133_not
g65863 not n10504 ; n10504_not
g65864 not n42103 ; n42103_not
g65865 not n21124 ; n21124_not
g65866 not n45010 ; n45010_not
g65867 not n21502 ; n21502_not
g65868 not n40240 ; n40240_not
g65869 not n30106 ; n30106_not
g65870 not n21115 ; n21115_not
g65871 not n10405 ; n10405_not
g65872 not n50221 ; n50221_not
g65873 not n30205 ; n30205_not
g65874 not n50302 ; n50302_not
g65875 not n40132 ; n40132_not
g65876 not n20512 ; n20512_not
g65877 not n42121 ; n42121_not
g65878 not n21520 ; n21520_not
g65879 not n42031 ; n42031_not
g65880 not n14410 ; n14410_not
g65881 not n21322 ; n21322_not
g65882 not n31132 ; n31132_not
g65883 not n21160 ; n21160_not
g65884 not n21151 ; n21151_not
g65885 not n42040 ; n42040_not
g65886 not n42112 ; n42112_not
g65887 not n21142 ; n21142_not
g65888 not n31141 ; n31141_not
g65889 not n50212 ; n50212_not
g65890 not n31420 ; n31420_not
g65891 not n30223 ; n30223_not
g65892 not n10441 ; n10441_not
g65893 not n10450 ; n10450_not
g65894 not n21412 ; n21412_not
g65895 not n31402 ; n31402_not
g65896 not n30232 ; n30232_not
g65897 not n30241 ; n30241_not
g65898 not n33031 ; n33031_not
g65899 not n31150 ; n31150_not
g65900 not n40222 ; n40222_not
g65901 not n55000 ; n55000_not
g65902 not n14500 ; n14500_not
g65903 not n30214 ; n30214_not
g65904 not n10432 ; n10432_not
g65905 not n50320 ; n50320_not
g65906 not n10243 ; n10243_not
g65907 not n10252 ; n10252_not
g65908 not n10261 ; n10261_not
g65909 not n41410 ; n41410_not
g65910 not n10270 ; n10270_not
g65911 not n10306 ; n10306_not
g65912 not n10315 ; n10315_not
g65913 not n31330 ; n31330_not
g65914 not n10333 ; n10333_not
g65915 not n32014 ; n32014_not
g65916 not n10801 ; n10801_not
g65917 not n10342 ; n10342_not
g65918 not n33400 ; n33400_not
g65919 not n10810 ; n10810_not
g65920 not n10900 ; n10900_not
g65921 not n10351 ; n10351_not
g65922 not n10144 ; n10144_not
g65923 not n31213 ; n31213_not
g65924 not n10153 ; n10153_not
g65925 not n10162 ; n10162_not
g65926 not n10171 ; n10171_not
g65927 not n10180 ; n10180_not
g65928 not n26101 ; n26101_not
g65929 not n10207 ; n10207_not
g65930 not n43120 ; n43120_not
g65931 not n10216 ; n10216_not
g65932 not n31321 ; n31321_not
g65933 not n10225 ; n10225_not
g65934 not n10234 ; n10234_not
g65935 not n21205 ; n21205_not
g65936 not n21304 ; n21304_not
g65937 not n10414 ; n10414_not
g65938 not n40312 ; n40312_not
g65939 not n42022 ; n42022_not
g65940 not n30115 ; n30115_not
g65941 not n40303 ; n40303_not
g65942 not n42130 ; n42130_not
g65943 not n31123 ; n31123_not
g65944 not n26002 ; n26002_not
g65945 not n41230 ; n41230_not
g65946 not n10360 ; n10360_not
g65947 not n31105 ; n31105_not
g65948 not n31204 ; n31204_not
g65949 not n15310 ; n15310_not
g65950 not n21250 ; n21250_not
g65951 not n21241 ; n21241_not
g65952 not n21232 ; n21232_not
g65953 not n15301 ; n15301_not
g65954 not n21223 ; n21223_not
g65955 not n30124 ; n30124_not
g65956 not n26020 ; n26020_not
g65957 not n40330 ; n40330_not
g65958 not n21214 ; n21214_not
g65959 not n31114 ; n31114_not
g65960 not n40321 ; n40321_not
g65961 not n26011 ; n26011_not
g65962 not n20107 ; n20107_not
g65963 not n20071 ; n20071_not
g65964 not n52021 ; n52021_not
g65965 not n20170 ; n20170_not
g65966 not n17101 ; n17101_not
g65967 not n20062 ; n20062_not
g65968 not n30331 ; n30331_not
g65969 not n27010 ; n27010_not
g65970 not n27001 ; n27001_not
g65971 not n11611 ; n11611_not
g65972 not n20125 ; n20125_not
g65973 not n11440 ; n11440_not
g65974 not n36001 ; n36001_not
g65975 not n25012 ; n25012_not
g65976 not n42301 ; n42301_not
g65977 not n11341 ; n11341_not
g65978 not n20116 ; n20116_not
g65979 not n11350 ; n11350_not
g65980 not n15103 ; n15103_not
g65981 not n11602 ; n11602_not
g65982 not n52210 ; n52210_not
g65983 not n20080 ; n20080_not
g65984 not n11404 ; n11404_not
g65985 not n20053 ; n20053_not
g65986 not n30322 ; n30322_not
g65987 not n20143 ; n20143_not
g65988 not n25102 ; n25102_not
g65989 not n25003 ; n25003_not
g65990 not n20710 ; n20710_not
g65991 not n52030 ; n52030_not
g65992 not n27100 ; n27100_not
g65993 not n20134 ; n20134_not
g65994 not n17011 ; n17011_not
g65995 not n16003 ; n16003_not
g65996 not n52201 ; n52201_not
g65997 not n50203 ; n50203_not
g65998 not n33202 ; n33202_not
g65999 not n42310 ; n42310_not
g66000 not n25030 ; n25030_not
g66001 not n11530 ; n11530_not
g66002 not n52120 ; n52120_not
g66003 not n43201 ; n43201_not
g66004 not n52003 ; n52003_not
g66005 not n20152 ; n20152_not
g66006 not n52111 ; n52111_not
g66007 not n52012 ; n52012_not
g66008 not n36010 ; n36010_not
g66009 not n43210 ; n43210_not
g66010 not n52102 ; n52102_not
g66011 not n11305 ; n11305_not
g66012 not n11314 ; n11314_not
g66013 not n21313 ; n21313_not
g66014 not n20161 ; n20161_not
g66015 not n19000 ; n19000_not
g66016 not n11323 ; n11323_not
g66017 not n16012 ; n16012_not
g66018 not n11332 ; n11332_not
g66019 not n25021 ; n25021_not
g66020 not n16021 ; n16021_not
g66021 not n16030 ; n16030_not
g66022 not n15013 ; n15013_not
g66023 not n32113 ; n32113_not
g66024 not n33211 ; n33211_not
g66025 not n31231 ; n31231_not
g66026 not n33220 ; n33220_not
g66027 not n30313 ; n30313_not
g66028 not n20044 ; n20044_not
g66029 not n30070 ; n30070_not
g66030 not n42400 ; n42400_not
g66031 not n25120 ; n25120_not
g66032 not n30061 ; n30061_not
g66033 not n41320 ; n41320_not
g66034 not n32302 ; n32302_not
g66035 not n50230 ; n50230_not
g66036 not n25111 ; n25111_not
g66037 not n26110 ; n26110_not
g66038 not n20027 ; n20027_not
g66039 not n26030 ; n26030_not
g66040 not n33050 ; n33050_not
g66041 not n15014 ; n15014_not
g66042 not n10424 ; n10424_not
g66043 not n27101 ; n27101_not
g66044 not n13106 ; n13106_not
g66045 not n34400 ; n34400_not
g66046 not n24023 ; n24023_not
g66047 not n51122 ; n51122_not
g66048 not n21305 ; n21305_not
g66049 not n30710 ; n30710_not
g66050 not n12503 ; n12503_not
g66051 not n13250 ; n13250_not
g66052 not n32051 ; n32051_not
g66053 not n41042 ; n41042_not
g66054 not n12512 ; n12512_not
g66055 not n10460 ; n10460_not
g66056 not n36101 ; n36101_not
g66057 not n42023 ; n42023_not
g66058 not n43121 ; n43121_not
g66059 not n42140 ; n42140_not
g66060 not n10361 ; n10361_not
g66061 not n23051 ; n23051_not
g66062 not n45011 ; n45011_not
g66063 not n30620 ; n30620_not
g66064 not n50042 ; n50042_not
g66065 not n41303 ; n41303_not
g66066 not n37100 ; n37100_not
g66067 not n23006 ; n23006_not
g66068 not n24050 ; n24050_not
g66069 not n27200 ; n27200_not
g66070 not n30413 ; n30413_not
g66071 not n42320 ; n42320_not
g66072 not n22304 ; n22304_not
g66073 not n26012 ; n26012_not
g66074 not n52013 ; n52013_not
g66075 not n30323 ; n30323_not
g66076 not n32141 ; n32141_not
g66077 not n41033 ; n41033_not
g66078 not n10613 ; n10613_not
g66079 not n45020 ; n45020_not
g66080 not n15023 ; n15023_not
g66081 not n10631 ; n10631_not
g66082 not n12008 ; n12008_not
g66083 not n24032 ; n24032_not
g66084 not n13124 ; n13124_not
g66085 not n55010 ; n55010_not
g66086 not n41024 ; n41024_not
g66087 not n24041 ; n24041_not
g66088 not n50321 ; n50321_not
g66089 not n13223 ; n13223_not
g66090 not n13160 ; n13160_not
g66091 not n41600 ; n41600_not
g66092 not n52103 ; n52103_not
g66093 not n13115 ; n13115_not
g66094 not n10622 ; n10622_not
g66095 not n16211 ; n16211_not
g66096 not n21422 ; n21422_not
g66097 not n30512 ; n30512_not
g66098 not n32600 ; n32600_not
g66099 not n10604 ; n10604_not
g66100 not n13232 ; n13232_not
g66101 not n42131 ; n42131_not
g66102 not n16112 ; n16112_not
g66103 not n21404 ; n21404_not
g66104 not n30233 ; n30233_not
g66105 not n42401 ; n42401_not
g66106 not n26021 ; n26021_not
g66107 not n10406 ; n10406_not
g66108 not n13052 ; n13052_not
g66109 not n32060 ; n32060_not
g66110 not n10505 ; n10505_not
g66111 not n41006 ; n41006_not
g66112 not n42104 ; n42104_not
g66113 not n30800 ; n30800_not
g66114 not n41060 ; n41060_not
g66115 not n16130 ; n16130_not
g66116 not n40142 ; n40142_not
g66117 not n53012 ; n53012_not
g66118 not n15005 ; n15005_not
g66119 not n41510 ; n41510_not
g66120 not n13016 ; n13016_not
g66121 not n40115 ; n40115_not
g66122 not n33023 ; n33023_not
g66123 not n13061 ; n13061_not
g66124 not n52031 ; n52031_not
g66125 not n33041 ; n33041_not
g66126 not n31430 ; n31430_not
g66127 not n14420 ; n14420_not
g66128 not n32114 ; n32114_not
g66129 not n15050 ; n15050_not
g66130 not n30611 ; n30611_not
g66131 not n25301 ; n25301_not
g66132 not n13070 ; n13070_not
g66133 not n35030 ; n35030_not
g66134 not n23024 ; n23024_not
g66135 not n41321 ; n41321_not
g66136 not n41501 ; n41501_not
g66137 not n10541 ; n10541_not
g66138 not n32123 ; n32123_not
g66139 not n27110 ; n27110_not
g66140 not n21350 ; n21350_not
g66141 not n13205 ; n13205_not
g66142 not n10532 ; n10532_not
g66143 not n13034 ; n13034_not
g66144 not n40124 ; n40124_not
g66145 not n23033 ; n23033_not
g66146 not n13025 ; n13025_not
g66147 not n22106 ; n22106_not
g66148 not n18002 ; n18002_not
g66149 not n50330 ; n50330_not
g66150 not n10550 ; n10550_not
g66151 not n20540 ; n20540_not
g66152 not n15500 ; n15500_not
g66153 not n53003 ; n53003_not
g66154 not n13043 ; n13043_not
g66155 not n10019 ; n10019_not
g66156 not n22115 ; n22115_not
g66157 not n10514 ; n10514_not
g66158 not n30242 ; n30242_not
g66159 not n30602 ; n30602_not
g66160 not n18011 ; n18011_not
g66161 not n50303 ; n50303_not
g66162 not n50060 ; n50060_not
g66163 not n42122 ; n42122_not
g66164 not n24005 ; n24005_not
g66165 not n52040 ; n52040_not
g66166 not n10442 ; n10442_not
g66167 not n53030 ; n53030_not
g66168 not n50051 ; n50051_not
g66169 not n31511 ; n31511_not
g66170 not n30080 ; n30080_not
g66171 not n43112 ; n43112_not
g66172 not n12521 ; n12521_not
g66173 not n35021 ; n35021_not
g66174 not n23114 ; n23114_not
g66175 not n36200 ; n36200_not
g66176 not n37010 ; n37010_not
g66177 not n44300 ; n44300_not
g66178 not n25310 ; n25310_not
g66179 not n24014 ; n24014_not
g66180 not n40160 ; n40160_not
g66181 not n14402 ; n14402_not
g66182 not n50213 ; n50213_not
g66183 not n20720 ; n20720_not
g66184 not n21314 ; n21314_not
g66185 not n26003 ; n26003_not
g66186 not n18020 ; n18020_not
g66187 not n42113 ; n42113_not
g66188 not n21332 ; n21332_not
g66189 not n14411 ; n14411_not
g66190 not n41051 ; n41051_not
g66191 not n53021 ; n53021_not
g66192 not n32105 ; n32105_not
g66193 not n12611 ; n12611_not
g66194 not n16121 ; n16121_not
g66195 not n23105 ; n23105_not
g66196 not n41312 ; n41312_not
g66197 not n30332 ; n30332_not
g66198 not n52022 ; n52022_not
g66199 not n32132 ; n32132_not
g66200 not n33014 ; n33014_not
g66201 not n54200 ; n54200_not
g66202 not n43202 ; n43202_not
g66203 not n13007 ; n13007_not
g66204 not n30314 ; n30314_not
g66205 not n10451 ; n10451_not
g66206 not n12530 ; n12530_not
g66207 not n16202 ; n16202_not
g66208 not n43211 ; n43211_not
g66209 not n28001 ; n28001_not
g66210 not n30530 ; n30530_not
g66211 not n28010 ; n28010_not
g66212 not n44021 ; n44021_not
g66213 not n26120 ; n26120_not
g66214 not n20603 ; n20603_not
g66215 not n32033 ; n32033_not
g66216 not n36002 ; n36002_not
g66217 not n12602 ; n12602_not
g66218 not n26111 ; n26111_not
g66219 not n42500 ; n42500_not
g66220 not n42203 ; n42203_not
g66221 not n51410 ; n51410_not
g66222 not n16013 ; n16013_not
g66223 not n36011 ; n36011_not
g66224 not n44030 ; n44030_not
g66225 not n43400 ; n43400_not
g66226 not n16004 ; n16004_not
g66227 not n54110 ; n54110_not
g66228 not n41402 ; n41402_not
g66229 not n20702 ; n20702_not
g66230 not n18200 ; n18200_not
g66231 not n50015 ; n50015_not
g66232 not n40007 ; n40007_not
g66233 not n44120 ; n44120_not
g66234 not n15122 ; n15122_not
g66235 not n52211 ; n52211_not
g66236 not n35201 ; n35201_not
g66237 not n45110 ; n45110_not
g66238 not n40016 ; n40016_not
g66239 not n52202 ; n52202_not
g66240 not n40025 ; n40025_not
g66241 not n44111 ; n44111_not
g66242 not n34013 ; n34013_not
g66243 not n20630 ; n20630_not
g66244 not n44102 ; n44102_not
g66245 not n54101 ; n54101_not
g66246 not n52220 ; n52220_not
g66247 not n26102 ; n26102_not
g66248 not n15140 ; n15140_not
g66249 not n53120 ; n53120_not
g66250 not n52400 ; n52400_not
g66251 not n16040 ; n16040_not
g66252 not n53102 ; n53102_not
g66253 not n16031 ; n16031_not
g66254 not n51302 ; n51302_not
g66255 not n31610 ; n31610_not
g66256 not n32006 ; n32006_not
g66257 not n51311 ; n51311_not
g66258 not n42221 ; n42221_not
g66259 not n15302 ; n15302_not
g66260 not n51212 ; n51212_not
g66261 not n51320 ; n51320_not
g66262 not n33401 ; n33401_not
g66263 not n51203 ; n51203_not
g66264 not n51113 ; n51113_not
g66265 not n51014 ; n51014_not
g66266 not n13331 ; n13331_not
g66267 not n51230 ; n51230_not
g66268 not n26201 ; n26201_not
g66269 not n20009 ; n20009_not
g66270 not n52301 ; n52301_not
g66271 not n56000 ; n56000_not
g66272 not n43220 ; n43220_not
g66273 not n13322 ; n13322_not
g66274 not n26210 ; n26210_not
g66275 not n46100 ; n46100_not
g66276 not n42230 ; n42230_not
g66277 not n51104 ; n51104_not
g66278 not n51221 ; n51221_not
g66279 not n52310 ; n52310_not
g66280 not n30305 ; n30305_not
g66281 not n20018 ; n20018_not
g66282 not n16400 ; n16400_not
g66283 not n15221 ; n15221_not
g66284 not n34130 ; n34130_not
g66285 not n36020 ; n36020_not
g66286 not n53111 ; n53111_not
g66287 not n15320 ; n15320_not
g66288 not n42212 ; n42212_not
g66289 not n44012 ; n44012_not
g66290 not n15203 ; n15203_not
g66291 not n26300 ; n26300_not
g66292 not n51140 ; n51140_not
g66293 not n51401 ; n51401_not
g66294 not n14600 ; n14600_not
g66295 not n31601 ; n31601_not
g66296 not n32015 ; n32015_not
g66297 not n46010 ; n46010_not
g66298 not n15230 ; n15230_not
g66299 not n16022 ; n16022_not
g66300 not n50024 ; n50024_not
g66301 not n15311 ; n15311_not
g66302 not n44003 ; n44003_not
g66303 not n13313 ; n13313_not
g66304 not n33410 ; n33410_not
g66305 not n46001 ; n46001_not
g66306 not n51023 ; n51023_not
g66307 not n17003 ; n17003_not
g66308 not n30503 ; n30503_not
g66309 not n30404 ; n30404_not
g66310 not n45101 ; n45101_not
g66311 not n30431 ; n30431_not
g66312 not n52121 ; n52121_not
g66313 not n22052 ; n22052_not
g66314 not n52004 ; n52004_not
g66315 not n27002 ; n27002_not
g66316 not n38000 ; n38000_not
g66317 not n27011 ; n27011_not
g66318 not n30422 ; n30422_not
g66319 not n18101 ; n18101_not
g66320 not n23042 ; n23042_not
g66321 not n35102 ; n35102_not
g66322 not n50033 ; n50033_not
g66323 not n43130 ; n43130_not
g66324 not n22061 ; n22061_not
g66325 not n10325 ; n10325_not
g66326 not n12701 ; n12701_not
g66327 not n42311 ; n42311_not
g66328 not n10334 ; n10334_not
g66329 not n21260 ; n21260_not
g66330 not n10343 ; n10343_not
g66331 not n52112 ; n52112_not
g66332 not n13241 ; n13241_not
g66333 not n41015 ; n41015_not
g66334 not n22070 ; n22070_not
g66335 not n10352 ; n10352_not
g66336 not n16103 ; n16103_not
g66337 not n37001 ; n37001_not
g66338 not n51041 ; n51041_not
g66339 not n17012 ; n17012_not
g66340 not n20513 ; n20513_not
g66341 not n30440 ; n30440_not
g66342 not n33032 ; n33032_not
g66343 not n20504 ; n20504_not
g66344 not n16220 ; n16220_not
g66345 not n23600 ; n23600_not
g66346 not n18110 ; n18110_not
g66347 not n20612 ; n20612_not
g66348 not n40052 ; n40052_not
g66349 not n33320 ; n33320_not
g66350 not n22025 ; n22025_not
g66351 not n16310 ; n16310_not
g66352 not n40061 ; n40061_not
g66353 not n15104 ; n15104_not
g66354 not n33500 ; n33500_not
g66355 not n40034 ; n40034_not
g66356 not n44201 ; n44201_not
g66357 not n40043 ; n40043_not
g66358 not n50006 ; n50006_not
g66359 not n13340 ; n13340_not
g66360 not n41330 ; n41330_not
g66361 not n44210 ; n44210_not
g66362 not n15113 ; n15113_not
g66363 not n15401 ; n15401_not
g66364 not n15032 ; n15032_not
g66365 not n42302 ; n42302_not
g66366 not n35111 ; n35111_not
g66367 not n33302 ; n33302_not
g66368 not n34031 ; n34031_not
g66369 not n52130 ; n52130_not
g66370 not n15410 ; n15410_not
g66371 not n50312 ; n50312_not
g66372 not n51500 ; n51500_not
g66373 not n27020 ; n27020_not
g66374 not n12800 ; n12800_not
g66375 not n31520 ; n31520_not
g66376 not n41411 ; n41411_not
g66377 not n35120 ; n35120_not
g66378 not n34022 ; n34022_not
g66379 not n30521 ; n30521_not
g66380 not n55100 ; n55100_not
g66381 not n21710 ; n21710_not
g66382 not n40205 ; n40205_not
g66383 not n11045 ; n11045_not
g66384 not n11450 ; n11450_not
g66385 not n21701 ; n21701_not
g66386 not n11054 ; n11054_not
g66387 not n40403 ; n40403_not
g66388 not n11621 ; n11621_not
g66389 not n32312 ; n32312_not
g66390 not n14033 ; n14033_not
g66391 not n40610 ; n40610_not
g66392 not n12170 ; n12170_not
g66393 not n14105 ; n14105_not
g66394 not n11063 ; n11063_not
g66395 not n30008 ; n30008_not
g66396 not n11009 ; n11009_not
g66397 not n32204 ; n32204_not
g66398 not n41204 ; n41204_not
g66399 not n50141 ; n50141_not
g66400 not n14060 ; n14060_not
g66401 not n25400 ; n25400_not
g66402 not n11027 ; n11027_not
g66403 not n31016 ; n31016_not
g66404 not n14501 ; n14501_not
g66405 not n32213 ; n32213_not
g66406 not n21440 ; n21440_not
g66407 not n32330 ; n32330_not
g66408 not n29000 ; n29000_not
g66409 not n41213 ; n41213_not
g66410 not n12143 ; n12143_not
g66411 not n17111 ; n17111_not
g66412 not n14141 ; n14141_not
g66413 not n11081 ; n11081_not
g66414 not n11414 ; n11414_not
g66415 not n53300 ; n53300_not
g66416 not n41222 ; n41222_not
g66417 not n11423 ; n11423_not
g66418 not n11072 ; n11072_not
g66419 not n14150 ; n14150_not
g66420 not n32222 ; n32222_not
g66421 not n14114 ; n14114_not
g66422 not n32231 ; n32231_not
g66423 not n31214 ; n31214_not
g66424 not n31304 ; n31304_not
g66425 not n11432 ; n11432_not
g66426 not n14123 ; n14123_not
g66427 not n14132 ; n14132_not
g66428 not n12152 ; n12152_not
g66429 not n11090 ; n11090_not
g66430 not n10712 ; n10712_not
g66431 not n50132 ; n50132_not
g66432 not n24500 ; n24500_not
g66433 not n12251 ; n12251_not
g66434 not n14006 ; n14006_not
g66435 not n24302 ; n24302_not
g66436 not n30017 ; n30017_not
g66437 not n10703 ; n10703_not
g66438 not n12242 ; n12242_not
g66439 not n14015 ; n14015_not
g66440 not n40223 ; n40223_not
g66441 not n43310 ; n43310_not
g66442 not n14240 ; n14240_not
g66443 not n30170 ; n30170_not
g66444 not n35012 ; n35012_not
g66445 not n10730 ; n10730_not
g66446 not n22250 ; n22250_not
g66447 not n12260 ; n12260_not
g66448 not n30125 ; n30125_not
g66449 not n31322 ; n31322_not
g66450 not n41123 ; n41123_not
g66451 not n54011 ; n54011_not
g66452 not n10721 ; n10721_not
g66453 not n19010 ; n19010_not
g66454 not n54020 ; n54020_not
g66455 not n50123 ; n50123_not
g66456 not n31313 ; n31313_not
g66457 not n10640 ; n10640_not
g66458 not n12215 ; n12215_not
g66459 not n14042 ; n14042_not
g66460 not n12161 ; n12161_not
g66461 not n14051 ; n14051_not
g66462 not n21323 ; n21323_not
g66463 not n30134 ; n30134_not
g66464 not n12206 ; n12206_not
g66465 not n34103 ; n34103_not
g66466 not n31007 ; n31007_not
g66467 not n14024 ; n14024_not
g66468 not n24311 ; n24311_not
g66469 not n30161 ; n30161_not
g66470 not n40133 ; n40133_not
g66471 not n12233 ; n12233_not
g66472 not n19001 ; n19001_not
g66473 not n40214 ; n40214_not
g66474 not n24320 ; n24320_not
g66475 not n34112 ; n34112_not
g66476 not n12224 ; n12224_not
g66477 not n50222 ; n50222_not
g66478 not n24140 ; n24140_not
g66479 not n34040 ; n34040_not
g66480 not n21620 ; n21620_not
g66481 not n24131 ; n24131_not
g66482 not n25220 ; n25220_not
g66483 not n31241 ; n31241_not
g66484 not n14303 ; n14303_not
g66485 not n14312 ; n14312_not
g66486 not n24122 ; n24122_not
g66487 not n12017 ; n12017_not
g66488 not n21800 ; n21800_not
g66489 not n24113 ; n24113_not
g66490 not n53201 ; n53201_not
g66491 not n41231 ; n41231_not
g66492 not n22214 ; n22214_not
g66493 not n21602 ; n21602_not
g66494 not n21611 ; n21611_not
g66495 not n12035 ; n12035_not
g66496 not n50105 ; n50105_not
g66497 not n11441 ; n11441_not
g66498 not n40421 ; n40421_not
g66499 not n30116 ; n30116_not
g66500 not n14330 ; n14330_not
g66501 not n14321 ; n14321_not
g66502 not n10910 ; n10910_not
g66503 not n50240 ; n50240_not
g66504 not n24104 ; n24104_not
g66505 not n22241 ; n22241_not
g66506 not n25211 ; n25211_not
g66507 not n25202 ; n25202_not
g66508 not n22232 ; n22232_not
g66509 not n40430 ; n40430_not
g66510 not n12107 ; n12107_not
g66511 not n25103 ; n25103_not
g66512 not n31223 ; n31223_not
g66513 not n11018 ; n11018_not
g66514 not n21530 ; n21530_not
g66515 not n14204 ; n14204_not
g66516 not n14213 ; n14213_not
g66517 not n41132 ; n41132_not
g66518 not n30152 ; n30152_not
g66519 not n12125 ; n12125_not
g66520 not n53210 ; n53210_not
g66521 not n21413 ; n21413_not
g66522 not n35210 ; n35210_not
g66523 not n24230 ; n24230_not
g66524 not n24221 ; n24221_not
g66525 not n24212 ; n24212_not
g66526 not n12062 ; n12062_not
g66527 not n30143 ; n30143_not
g66528 not n25130 ; n25130_not
g66529 not n31232 ; n31232_not
g66530 not n24203 ; n24203_not
g66531 not n32240 ; n32240_not
g66532 not n12053 ; n12053_not
g66533 not n41420 ; n41420_not
g66534 not n14222 ; n14222_not
g66535 not n40601 ; n40601_not
g66536 not n25112 ; n25112_not
g66537 not n12080 ; n12080_not
g66538 not n40412 ; n40412_not
g66539 not n14231 ; n14231_not
g66540 not n25121 ; n25121_not
g66541 not n43301 ; n43301_not
g66542 not n30215 ; n30215_not
g66543 not n11603 ; n11603_not
g66544 not n40700 ; n40700_not
g66545 not n47000 ; n47000_not
g66546 not n35003 ; n35003_not
g66547 not n12071 ; n12071_not
g66548 not n41141 ; n41141_not
g66549 not n21512 ; n21512_not
g66550 not n12440 ; n12440_not
g66551 not n22007 ; n22007_not
g66552 not n22151 ; n22151_not
g66553 not n22124 ; n22124_not
g66554 not n11612 ; n11612_not
g66555 not n42041 ; n42041_not
g66556 not n22205 ; n22205_not
g66557 not n20522 ; n20522_not
g66558 not n10811 ; n10811_not
g66559 not n41150 ; n41150_not
g66560 not n10820 ; n10820_not
g66561 not n11531 ; n11531_not
g66562 not n12341 ; n12341_not
g66563 not n41105 ; n41105_not
g66564 not n30035 ; n30035_not
g66565 not n30053 ; n30053_not
g66566 not n17102 ; n17102_not
g66567 not n25013 ; n25013_not
g66568 not n41114 ; n41114_not
g66569 not n17021 ; n17021_not
g66570 not n10370 ; n10370_not
g66571 not n10802 ; n10802_not
g66572 not n40511 ; n40511_not
g66573 not n12350 ; n12350_not
g66574 not n54002 ; n54002_not
g66575 not n41240 ; n41240_not
g66576 not n22034 ; n22034_not
g66577 not n19100 ; n19100_not
g66578 not n22160 ; n22160_not
g66579 not n40232 ; n40232_not
g66580 not n12404 ; n12404_not
g66581 not n14510 ; n14510_not
g66582 not n30701 ; n30701_not
g66583 not n31160 ; n31160_not
g66584 not n13151 ; n13151_not
g66585 not n12422 ; n12422_not
g66586 not n40502 ; n40502_not
g66587 not n12413 ; n12413_not
g66588 not n10415 ; n10415_not
g66589 not n45002 ; n45002_not
g66590 not n30044 ; n30044_not
g66591 not n25004 ; n25004_not
g66592 not n40250 ; n40250_not
g66593 not n50150 ; n50150_not
g66594 not n30206 ; n30206_not
g66595 not n51032 ; n51032_not
g66596 not n42050 ; n42050_not
g66597 not n12431 ; n12431_not
g66598 not n32303 ; n32303_not
g66599 not n12116 ; n12116_not
g66600 not n45200 ; n45200_not
g66601 not n32150 ; n32150_not
g66602 not n42005 ; n42005_not
g66603 not n40340 ; n40340_not
g66604 not n40520 ; n40520_not
g66605 not n25040 ; n25040_not
g66606 not n31340 ; n31340_not
g66607 not n12305 ; n12305_not
g66608 not n31331 ; n31331_not
g66609 not n34121 ; n34121_not
g66610 not n30026 ; n30026_not
g66611 not n30062 ; n30062_not
g66612 not n22142 ; n22142_not
g66613 not n35300 ; n35300_not
g66614 not n11540 ; n11540_not
g66615 not n11513 ; n11513_not
g66616 not n12026 ; n12026_not
g66617 not n50231 ; n50231_not
g66618 not n25022 ; n25022_not
g66619 not n40313 ; n40313_not
g66620 not n12323 ; n12323_not
g66621 not n11522 ; n11522_not
g66622 not n32024 ; n32024_not
g66623 not n21503 ; n21503_not
g66624 not n12332 ; n12332_not
g66625 not n40304 ; n40304_not
g66626 not n25031 ; n25031_not
g66627 not n40331 ; n40331_not
g66628 not n31403 ; n31403_not
g66629 not n40322 ; n40322_not
g66630 not n30224 ; n30224_not
g66631 not n12314 ; n12314_not
g66632 not n41106 ; n41106_not
g66633 not n41313 ; n41313_not
g66634 not n20028 ; n20028_not
g66635 not n22107 ; n22107_not
g66636 not n43032 ; n43032_not
g66637 not n20802 ; n20802_not
g66638 not n20361 ; n20361_not
g66639 not n23034 ; n23034_not
g66640 not n33213 ; n33213_not
g66641 not n14142 ; n14142_not
g66642 not n53400 ; n53400_not
g66643 not n45102 ; n45102_not
g66644 not n15015 ; n15015_not
g66645 not n13341 ; n13341_not
g66646 not n22044 ; n22044_not
g66647 not n20019 ; n20019_not
g66648 not n33231 ; n33231_not
g66649 not n30315 ; n30315_not
g66650 not n30540 ; n30540_not
g66651 not n50430 ; n50430_not
g66652 not n14700 ; n14700_not
g66653 not n32700 ; n32700_not
g66654 not n33150 ; n33150_not
g66655 not n50223 ; n50223_not
g66656 not n20109 ; n20109_not
g66657 not n15411 ; n15411_not
g66658 not n43401 ; n43401_not
g66659 not n15150 ; n15150_not
g66660 not n33222 ; n33222_not
g66661 not n15024 ; n15024_not
g66662 not n14133 ; n14133_not
g66663 not n50160 ; n50160_not
g66664 not n13260 ; n13260_not
g66665 not n22062 ; n22062_not
g66666 not n14151 ; n14151_not
g66667 not n20325 ; n20325_not
g66668 not n30054 ; n30054_not
g66669 not n23061 ; n23061_not
g66670 not n20136 ; n20136_not
g66671 not n43212 ; n43212_not
g66672 not n14304 ; n14304_not
g66673 not n30063 ; n30063_not
g66674 not n14322 ; n14322_not
g66675 not n51024 ; n51024_not
g66676 not n22224 ; n22224_not
g66677 not n14124 ; n14124_not
g66678 not n23043 ; n23043_not
g66679 not n15033 ; n15033_not
g66680 not n13332 ; n13332_not
g66681 not n34023 ; n34023_not
g66682 not n22071 ; n22071_not
g66683 not n51051 ; n51051_not
g66684 not n30360 ; n30360_not
g66685 not n33105 ; n33105_not
g66686 not n14160 ; n14160_not
g66687 not n14313 ; n14313_not
g66688 not n15420 ; n15420_not
g66689 not n41025 ; n41025_not
g66690 not n20334 ; n20334_not
g66691 not n30009 ; n30009_not
g66692 not n13305 ; n13305_not
g66693 not n14043 ; n14043_not
g66694 not n20343 ; n20343_not
g66695 not n14214 ; n14214_not
g66696 not n33240 ; n33240_not
g66697 not n20901 ; n20901_not
g66698 not n41016 ; n41016_not
g66699 not n20730 ; n20730_not
g66700 not n21324 ; n21324_not
g66701 not n44202 ; n44202_not
g66702 not n33312 ; n33312_not
g66703 not n50142 ; n50142_not
g66704 not n14205 ; n14205_not
g66705 not n21270 ; n21270_not
g66706 not n22134 ; n22134_not
g66707 not n41052 ; n41052_not
g66708 not n15105 ; n15105_not
g66709 not n41430 ; n41430_not
g66710 not n14034 ; n14034_not
g66711 not n16320 ; n16320_not
g66712 not n43041 ; n43041_not
g66713 not n23016 ; n23016_not
g66714 not n20910 ; n20910_not
g66715 not n21333 ; n21333_not
g66716 not n32610 ; n32610_not
g66717 not n14241 ; n14241_not
g66718 not n20703 ; n20703_not
g66719 not n44310 ; n44310_not
g66720 not n22161 ; n22161_not
g66721 not n37101 ; n37101_not
g66722 not n50133 ; n50133_not
g66723 not n30090 ; n30090_not
g66724 not n14061 ; n14061_not
g66725 not n30333 ; n30333_not
g66726 not n14232 ; n14232_not
g66727 not n41034 ; n41034_not
g66728 not n41340 ; n41340_not
g66729 not n14070 ; n14070_not
g66730 not n41043 ; n41043_not
g66731 not n22152 ; n22152_not
g66732 not n30018 ; n30018_not
g66733 not n33204 ; n33204_not
g66734 not n13323 ; n13323_not
g66735 not n13800 ; n13800_not
g66736 not n30027 ; n30027_not
g66737 not n14052 ; n14052_not
g66738 not n14250 ; n14250_not
g66739 not n21315 ; n21315_not
g66740 not n14223 ; n14223_not
g66741 not n33132 ; n33132_not
g66742 not n41061 ; n41061_not
g66743 not n16302 ; n16302_not
g66744 not n50115 ; n50115_not
g66745 not n22206 ; n22206_not
g66746 not n20118 ; n20118_not
g66747 not n22116 ; n22116_not
g66748 not n30324 ; n30324_not
g66749 not n14016 ; n14016_not
g66750 not n30045 ; n30045_not
g66751 not n41322 ; n41322_not
g66752 not n20352 ; n20352_not
g66753 not n20820 ; n20820_not
g66754 not n34005 ; n34005_not
g66755 not n41070 ; n41070_not
g66756 not n55200 ; n55200_not
g66757 not n43500 ; n43500_not
g66758 not n33123 ; n33123_not
g66759 not n30351 ; n30351_not
g66760 not n20811 ; n20811_not
g66761 not n14115 ; n14115_not
g66762 not n20370 ; n20370_not
g66763 not n14007 ; n14007_not
g66764 not n33114 ; n33114_not
g66765 not n43410 ; n43410_not
g66766 not n30036 ; n30036_not
g66767 not n30261 ; n30261_not
g66768 not n30342 ; n30342_not
g66769 not n20127 ; n20127_not
g66770 not n20712 ; n20712_not
g66771 not n30144 ; n30144_not
g66772 not n30108 ; n30108_not
g66773 not n41007 ; n41007_not
g66774 not n15060 ; n15060_not
g66775 not n15114 ; n15114_not
g66776 not n33330 ; n33330_not
g66777 not n55110 ; n55110_not
g66778 not n50205 ; n50205_not
g66779 not n51033 ; n51033_not
g66780 not n44040 ; n44040_not
g66781 not n13350 ; n13350_not
g66782 not n14025 ; n14025_not
g66783 not n15123 ; n15123_not
g66784 not n15402 ; n15402_not
g66785 not n33141 ; n33141_not
g66786 not n15600 ; n15600_not
g66787 not n14106 ; n14106_not
g66788 not n21513 ; n21513_not
g66789 not n21504 ; n21504_not
g66790 not n15510 ; n15510_not
g66791 not n50412 ; n50412_not
g66792 not n37011 ; n37011_not
g66793 not n50070 ; n50070_not
g66794 not n22215 ; n22215_not
g66795 not n20208 ; n20208_not
g66796 not n37020 ; n37020_not
g66797 not n34113 ; n34113_not
g66798 not n30252 ; n30252_not
g66799 not n30414 ; n30414_not
g66800 not n41421 ; n41421_not
g66801 not n30450 ; n30450_not
g66802 not n20271 ; n20271_not
g66803 not n33060 ; n33060_not
g66804 not n22440 ; n22440_not
g66805 not n15501 ; n15501_not
g66806 not n15303 ; n15303_not
g66807 not n21342 ; n21342_not
g66808 not n30441 ; n30441_not
g66809 not n20253 ; n20253_not
g66810 not n13602 ; n13602_not
g66811 not n22512 ; n22512_not
g66812 not n21522 ; n21522_not
g66813 not n22503 ; n22503_not
g66814 not n14412 ; n14412_not
g66815 not n43104 ; n43104_not
g66816 not n40710 ; n40710_not
g66817 not n20550 ; n20550_not
g66818 not n33033 ; n33033_not
g66819 not n41232 ; n41232_not
g66820 not n20262 ; n20262_not
g66821 not n21261 ; n21261_not
g66822 not n20280 ; n20280_not
g66823 not n22413 ; n22413_not
g66824 not n21252 ; n21252_not
g66825 not n20451 ; n20451_not
g66826 not n15330 ; n15330_not
g66827 not n30270 ; n30270_not
g66828 not n34041 ; n34041_not
g66829 not n22404 ; n22404_not
g66830 not n30405 ; n30405_not
g66831 not n21243 ; n21243_not
g66832 not n13242 ; n13242_not
g66833 not n20505 ; n20505_not
g66834 not n22242 ; n22242_not
g66835 not n14340 ; n14340_not
g66836 not n14331 ; n14331_not
g66837 not n41223 ; n41223_not
g66838 not n41403 ; n41403_not
g66839 not n22080 ; n22080_not
g66840 not n22701 ; n22701_not
g66841 not n33042 ; n33042_not
g66842 not n22710 ; n22710_not
g66843 not n13233 ; n13233_not
g66844 not n34140 ; n34140_not
g66845 not n22431 ; n22431_not
g66846 not n15312 ; n15312_not
g66847 not n50340 ; n50340_not
g66848 not n34122 ; n34122_not
g66849 not n20460 ; n20460_not
g66850 not n15321 ; n15321_not
g66851 not n22422 ; n22422_not
g66852 not n50052 ; n50052_not
g66853 not n50322 ; n50322_not
g66854 not n15231 ; n15231_not
g66855 not n22602 ; n22602_not
g66856 not n20226 ; n20226_not
g66857 not n20235 ; n20235_not
g66858 not n15222 ; n15222_not
g66859 not n34203 ; n34203_not
g66860 not n21450 ; n21450_not
g66861 not n30423 ; n30423_not
g66862 not n22611 ; n22611_not
g66863 not n34230 ; n34230_not
g66864 not n45021 ; n45021_not
g66865 not n13161 ; n13161_not
g66866 not n41205 ; n41205_not
g66867 not n15240 ; n15240_not
g66868 not n50313 ; n50313_not
g66869 not n22125 ; n22125_not
g66870 not n13152 ; n13152_not
g66871 not n41250 ; n41250_not
g66872 not n21432 ; n21432_not
g66873 not n15204 ; n15204_not
g66874 not n20532 ; n20532_not
g66875 not n41412 ; n41412_not
g66876 not n14601 ; n14601_not
g66877 not n34212 ; n34212_not
g66878 not n21414 ; n21414_not
g66879 not n33006 ; n33006_not
g66880 not n21405 ; n21405_not
g66881 not n40701 ; n40701_not
g66882 not n43311 ; n43311_not
g66883 not n34221 ; n34221_not
g66884 not n43050 ; n43050_not
g66885 not n43320 ; n43320_not
g66886 not n43122 ; n43122_not
g66887 not n13143 ; n13143_not
g66888 not n55020 ; n55020_not
g66889 not n41214 ; n41214_not
g66890 not n43131 ; n43131_not
g66891 not n22170 ; n22170_not
g66892 not n14430 ; n14430_not
g66893 not n14511 ; n14511_not
g66894 not n13611 ; n13611_not
g66895 not n22530 ; n22530_not
g66896 not n13206 ; n13206_not
g66897 not n30432 ; n30432_not
g66898 not n14421 ; n14421_not
g66899 not n14520 ; n14520_not
g66900 not n50403 ; n50403_not
g66901 not n22521 ; n22521_not
g66902 not n13701 ; n13701_not
g66903 not n22620 ; n22620_not
g66904 not n43302 ; n43302_not
g66905 not n20514 ; n20514_not
g66906 not n20244 ; n20244_not
g66907 not n20217 ; n20217_not
g66908 not n50331 ; n50331_not
g66909 not n13710 ; n13710_not
g66910 not n14502 ; n14502_not
g66911 not n33024 ; n33024_not
g66912 not n13620 ; n13620_not
g66913 not n21360 ; n21360_not
g66914 not n20163 ; n20163_not
g66915 not n20640 ; n20640_not
g66916 not n44211 ; n44211_not
g66917 not n41133 ; n41133_not
g66918 not n21063 ; n21063_not
g66919 not n20604 ; n20604_not
g66920 not n13431 ; n13431_not
g66921 not n44022 ; n44022_not
g66922 not n21054 ; n21054_not
g66923 not n14610 ; n14610_not
g66924 not n20613 ; n20613_not
g66925 not n43221 ; n43221_not
g66926 not n43014 ; n43014_not
g66927 not n13422 ; n13422_not
g66928 not n50250 ; n50250_not
g66929 not n34050 ; n34050_not
g66930 not n44013 ; n44013_not
g66931 not n50421 ; n50421_not
g66932 not n20424 ; n20424_not
g66933 not n41151 ; n41151_not
g66934 not n43005 ; n43005_not
g66935 not n15132 ; n15132_not
g66936 not n20172 ; n20172_not
g66937 not n21108 ; n21108_not
g66938 not n30135 ; n30135_not
g66939 not n41142 ; n41142_not
g66940 not n43230 ; n43230_not
g66941 not n21090 ; n21090_not
g66942 not n13440 ; n13440_not
g66943 not n21081 ; n21081_not
g66944 not n21072 ; n21072_not
g66945 not n41124 ; n41124_not
g66946 not n21018 ; n21018_not
g66947 not n21009 ; n21009_not
g66948 not n20406 ; n20406_not
g66949 not n44031 ; n44031_not
g66950 not n34032 ; n34032_not
g66951 not n50232 ; n50232_not
g66952 not n41115 ; n41115_not
g66953 not n20145 ; n20145_not
g66954 not n44301 ; n44301_not
g66955 not n20415 ; n20415_not
g66956 not n20316 ; n20316_not
g66957 not n21045 ; n21045_not
g66958 not n22251 ; n22251_not
g66959 not n51006 ; n51006_not
g66960 not n45111 ; n45111_not
g66961 not n38100 ; n38100_not
g66962 not n30126 ; n30126_not
g66963 not n13413 ; n13413_not
g66964 not n21036 ; n21036_not
g66965 not n50061 ; n50061_not
g66966 not n20154 ; n20154_not
g66967 not n43023 ; n43023_not
g66968 not n13404 ; n13404_not
g66969 not n21027 ; n21027_not
g66970 not n21207 ; n21207_not
g66971 not n53310 ; n53310_not
g66972 not n22260 ; n22260_not
g66973 not n13503 ; n13503_not
g66974 not n44220 ; n44220_not
g66975 not n34302 ; n34302_not
g66976 not n20181 ; n20181_not
g66977 not n21180 ; n21180_not
g66978 not n44004 ; n44004_not
g66979 not n15042 ; n15042_not
g66980 not n22350 ; n22350_not
g66981 not n21234 ; n21234_not
g66982 not n13530 ; n13530_not
g66983 not n13251 ; n13251_not
g66984 not n21225 ; n21225_not
g66985 not n30513 ; n30513_not
g66986 not n13521 ; n13521_not
g66987 not n33303 ; n33303_not
g66988 not n20190 ; n20190_not
g66989 not n13512 ; n13512_not
g66990 not n20442 ; n20442_not
g66991 not n21216 ; n21216_not
g66992 not n20523 ; n20523_not
g66993 not n21144 ; n21144_not
g66994 not n41160 ; n41160_not
g66995 not n21135 ; n21135_not
g66996 not n22800 ; n22800_not
g66997 not n20307 ; n20307_not
g66998 not n20622 ; n20622_not
g66999 not n22314 ; n22314_not
g67000 not n43140 ; n43140_not
g67001 not n21126 ; n21126_not
g67002 not n21423 ; n21423_not
g67003 not n22305 ; n22305_not
g67004 not n34320 ; n34320_not
g67005 not n21117 ; n21117_not
g67006 not n22341 ; n22341_not
g67007 not n22035 ; n22035_not
g67008 not n34311 ; n34311_not
g67009 not n53301 ; n53301_not
g67010 not n21171 ; n21171_not
g67011 not n22332 ; n22332_not
g67012 not n30522 ; n30522_not
g67013 not n20433 ; n20433_not
g67014 not n21162 ; n21162_not
g67015 not n22323 ; n22323_not
g67016 not n21153 ; n21153_not
g67017 not n23601 ; n23601_not
g67018 not n36030 ; n36030_not
g67019 not n31017 ; n31017_not
g67020 not n12171 ; n12171_not
g67021 not n12162 ; n12162_not
g67022 not n25320 ; n25320_not
g67023 not n12207 ; n12207_not
g67024 not n41502 ; n41502_not
g67025 not n54021 ; n54021_not
g67026 not n36021 ; n36021_not
g67027 not n31422 ; n31422_not
g67028 not n12216 ; n12216_not
g67029 not n12153 ; n12153_not
g67030 not n12225 ; n12225_not
g67031 not n24420 ; n24420_not
g67032 not n29010 ; n29010_not
g67033 not n42510 ; n42510_not
g67034 not n24411 ; n24411_not
g67035 not n54030 ; n54030_not
g67036 not n42231 ; n42231_not
g67037 not n51231 ; n51231_not
g67038 not n10461 ; n10461_not
g67039 not n56001 ; n56001_not
g67040 not n31413 ; n31413_not
g67041 not n12180 ; n12180_not
g67042 not n10470 ; n10470_not
g67043 not n40170 ; n40170_not
g67044 not n12261 ; n12261_not
g67045 not n54003 ; n54003_not
g67046 not n12270 ; n12270_not
g67047 not n37110 ; n37110_not
g67048 not n32502 ; n32502_not
g67049 not n12126 ; n12126_not
g67050 not n36012 ; n36012_not
g67051 not n36003 ; n36003_not
g67052 not n31431 ; n31431_not
g67053 not n12117 ; n12117_not
g67054 not n52014 ; n52014_not
g67055 not n41511 ; n41511_not
g67056 not n31440 ; n31440_not
g67057 not n40134 ; n40134_not
g67058 not n10506 ; n10506_not
g67059 not n52104 ; n52104_not
g67060 not n40125 ; n40125_not
g67061 not n42312 ; n42312_not
g67062 not n25311 ; n25311_not
g67063 not n31008 ; n31008_not
g67064 not n51510 ; n51510_not
g67065 not n12234 ; n12234_not
g67066 not n12243 ; n12243_not
g67067 not n17400 ; n17400_not
g67068 not n55002 ; n55002_not
g67069 not n42501 ; n42501_not
g67070 not n51330 ; n51330_not
g67071 not n12252 ; n12252_not
g67072 not n40152 ; n40152_not
g67073 not n54012 ; n54012_not
g67074 not n31071 ; n31071_not
g67075 not n11910 ; n11910_not
g67076 not n10425 ; n10425_not
g67077 not n23115 ; n23115_not
g67078 not n11451 ; n11451_not
g67079 not n35400 ; n35400_not
g67080 not n31062 ; n31062_not
g67081 not n11442 ; n11442_not
g67082 not n45030 ; n45030_not
g67083 not n50520 ; n50520_not
g67084 not n45201 ; n45201_not
g67085 not n35301 ; n35301_not
g67086 not n11433 ; n11433_not
g67087 not n31053 ; n31053_not
g67088 not n11415 ; n11415_not
g67089 not n18012 ; n18012_not
g67090 not n18102 ; n18102_not
g67091 not n27012 ; n27012_not
g67092 not n10407 ; n10407_not
g67093 not n51402 ; n51402_not
g67094 not n52122 ; n52122_not
g67095 not n31080 ; n31080_not
g67096 not n17103 ; n17103_not
g67097 not n27021 ; n27021_not
g67098 not n40224 ; n40224_not
g67099 not n18003 ; n18003_not
g67100 not n11901 ; n11901_not
g67101 not n10416 ; n10416_not
g67102 not n52005 ; n52005_not
g67103 not n40215 ; n40215_not
g67104 not n12063 ; n12063_not
g67105 not n24510 ; n24510_not
g67106 not n42006 ; n42006_not
g67107 not n24501 ; n24501_not
g67108 not n10452 ; n10452_not
g67109 not n12072 ; n12072_not
g67110 not n17301 ; n17301_not
g67111 not n51312 ; n51312_not
g67112 not n51303 ; n51303_not
g67113 not n12090 ; n12090_not
g67114 not n31035 ; n31035_not
g67115 not n12108 ; n12108_not
g67116 not n41241 ; n41241_not
g67117 not n52113 ; n52113_not
g67118 not n29001 ; n29001_not
g67119 not n12135 ; n12135_not
g67120 not n31026 ; n31026_not
g67121 not n17310 ; n17310_not
g67122 not n24600 ; n24600_not
g67123 not n32340 ; n32340_not
g67124 not n42060 ; n42060_not
g67125 not n12018 ; n12018_not
g67126 not n12027 ; n12027_not
g67127 not n31044 ; n31044_not
g67128 not n12045 ; n12045_not
g67129 not n51321 ; n51321_not
g67130 not n52500 ; n52500_not
g67131 not n51501 ; n51501_not
g67132 not n29100 ; n29100_not
g67133 not n10254 ; n10254_not
g67134 not n12432 ; n12432_not
g67135 not n26220 ; n26220_not
g67136 not n42141 ; n42141_not
g67137 not n32304 ; n32304_not
g67138 not n10263 ; n10263_not
g67139 not n12036 ; n12036_not
g67140 not n54210 ; n54210_not
g67141 not n12441 ; n12441_not
g67142 not n10272 ; n10272_not
g67143 not n10281 ; n10281_not
g67144 not n30702 ; n30702_not
g67145 not n12450 ; n12450_not
g67146 not n10371 ; n10371_not
g67147 not n10191 ; n10191_not
g67148 not n12405 ; n12405_not
g67149 not n10209 ; n10209_not
g67150 not n10218 ; n10218_not
g67151 not n42132 ; n42132_not
g67152 not n52311 ; n52311_not
g67153 not n52023 ; n52023_not
g67154 not n10227 ; n10227_not
g67155 not n42033 ; n42033_not
g67156 not n10236 ; n10236_not
g67157 not n12414 ; n12414_not
g67158 not n40107 ; n40107_not
g67159 not n10245 ; n10245_not
g67160 not n12423 ; n12423_not
g67161 not n27201 ; n27201_not
g67162 not n10317 ; n10317_not
g67163 not n12504 ; n12504_not
g67164 not n10308 ; n10308_not
g67165 not n36300 ; n36300_not
g67166 not n17013 ; n17013_not
g67167 not n19101 ; n19101_not
g67168 not n34401 ; n34401_not
g67169 not n12513 ; n12513_not
g67170 not n10290 ; n10290_not
g67171 not n12522 ; n12522_not
g67172 not n30810 ; n30810_not
g67173 not n31503 ; n31503_not
g67174 not n12540 ; n12540_not
g67175 not n31611 ; n31611_not
g67176 not n30711 ; n30711_not
g67177 not n10362 ; n10362_not
g67178 not n45210 ; n45210_not
g67179 not n52032 ; n52032_not
g67180 not n17022 ; n17022_not
g67181 not n17220 ; n17220_not
g67182 not n42150 ; n42150_not
g67183 not n10344 ; n10344_not
g67184 not n10326 ; n10326_not
g67185 not n39000 ; n39000_not
g67186 not n10047 ; n10047_not
g67187 not n12333 ; n12333_not
g67188 not n10056 ; n10056_not
g67189 not n46110 ; n46110_not
g67190 not n42105 ; n42105_not
g67191 not n10065 ; n10065_not
g67192 not n42330 ; n42330_not
g67193 not n26202 ; n26202_not
g67194 not n12342 ; n12342_not
g67195 not n10074 ; n10074_not
g67196 not n10083 ; n10083_not
g67197 not n12351 ; n12351_not
g67198 not n42321 ; n42321_not
g67199 not n12306 ; n12306_not
g67200 not n10515 ; n10515_not
g67201 not n27102 ; n27102_not
g67202 not n12315 ; n12315_not
g67203 not n27111 ; n27111_not
g67204 not n41520 ; n41520_not
g67205 not n10524 ; n10524_not
g67206 not n32511 ; n32511_not
g67207 not n10029 ; n10029_not
g67208 not n12324 ; n12324_not
g67209 not n10038 ; n10038_not
g67210 not n50700 ; n50700_not
g67211 not n32061 ; n32061_not
g67212 not n42411 ; n42411_not
g67213 not n10137 ; n10137_not
g67214 not n10146 ; n10146_not
g67215 not n42123 ; n42123_not
g67216 not n10155 ; n10155_not
g67217 not n32070 ; n32070_not
g67218 not n10164 ; n10164_not
g67219 not n10434 ; n10434_not
g67220 not n10173 ; n10173_not
g67221 not n32313 ; n32313_not
g67222 not n32520 ; n32520_not
g67223 not n10182 ; n10182_not
g67224 not n26211 ; n26211_not
g67225 not n18021 ; n18021_not
g67226 not n10092 ; n10092_not
g67227 not n42114 ; n42114_not
g67228 not n36111 ; n36111_not
g67229 not n10119 ; n10119_not
g67230 not n12081 ; n12081_not
g67231 not n16410 ; n16410_not
g67232 not n12360 ; n12360_not
g67233 not n52302 ; n52302_not
g67234 not n18030 ; n18030_not
g67235 not n10128 ; n10128_not
g67236 not n51240 ; n51240_not
g67237 not n46101 ; n46101_not
g67238 not n50610 ; n50610_not
g67239 not n11037 ; n11037_not
g67240 not n26112 ; n26112_not
g67241 not n17121 ; n17121_not
g67242 not n25104 ; n25104_not
g67243 not n11406 ; n11406_not
g67244 not n51141 ; n51141_not
g67245 not n52203 ; n52203_not
g67246 not n11424 ; n11424_not
g67247 not n25401 ; n25401_not
g67248 not n11019 ; n11019_not
g67249 not n11325 ; n11325_not
g67250 not n41610 ; n41610_not
g67251 not n11334 ; n11334_not
g67252 not n35220 ; n35220_not
g67253 not n11343 ; n11343_not
g67254 not n11055 ; n11055_not
g67255 not n11352 ; n11352_not
g67256 not n25140 ; n25140_not
g67257 not n31233 ; n31233_not
g67258 not n11361 ; n11361_not
g67259 not n25131 ; n25131_not
g67260 not n11370 ; n11370_not
g67261 not n25122 ; n25122_not
g67262 not n31224 ; n31224_not
g67263 not n25113 ; n25113_not
g67264 not n31206 ; n31206_not
g67265 not n18120 ; n18120_not
g67266 not n19002 ; n19002_not
g67267 not n51420 ; n51420_not
g67268 not n11316 ; n11316_not
g67269 not n11307 ; n11307_not
g67270 not n42600 ; n42600_not
g67271 not n18300 ; n18300_not
g67272 not n51600 ; n51600_not
g67273 not n11280 ; n11280_not
g67274 not n25050 ; n25050_not
g67275 not n19011 ; n19011_not
g67276 not n11505 ; n11505_not
g67277 not n36102 ; n36102_not
g67278 not n54201 ; n54201_not
g67279 not n25410 ; n25410_not
g67280 not n52230 ; n52230_not
g67281 not n11460 ; n11460_not
g67282 not n32322 ; n32322_not
g67283 not n50511 ; n50511_not
g67284 not n11145 ; n11145_not
g67285 not n11208 ; n11208_not
g67286 not n11217 ; n11217_not
g67287 not n11136 ; n11136_not
g67288 not n11226 ; n11226_not
g67289 not n25203 ; n25203_not
g67290 not n25212 ; n25212_not
g67291 not n11235 ; n11235_not
g67292 not n51150 ; n51150_not
g67293 not n11028 ; n11028_not
g67294 not n31242 ; n31242_not
g67295 not n11127 ; n11127_not
g67296 not n18210 ; n18210_not
g67297 not n54300 ; n54300_not
g67298 not n11181 ; n11181_not
g67299 not n11172 ; n11172_not
g67300 not n35202 ; n35202_not
g67301 not n11163 ; n11163_not
g67302 not n17202 ; n17202_not
g67303 not n11190 ; n11190_not
g67304 not n11154 ; n11154_not
g67305 not n38010 ; n38010_not
g67306 not n11091 ; n11091_not
g67307 not n25014 ; n25014_not
g67308 not n31260 ; n31260_not
g67309 not n25005 ; n25005_not
g67310 not n31251 ; n31251_not
g67311 not n52212 ; n52212_not
g67312 not n41601 ; n41601_not
g67313 not n10920 ; n10920_not
g67314 not n11244 ; n11244_not
g67315 not n52221 ; n52221_not
g67316 not n11118 ; n11118_not
g67317 not n25041 ; n25041_not
g67318 not n11253 ; n11253_not
g67319 not n11109 ; n11109_not
g67320 not n11262 ; n11262_not
g67321 not n18201 ; n18201_not
g67322 not n25032 ; n25032_not
g67323 not n25023 ; n25023_not
g67324 not n11271 ; n11271_not
g67325 not n17211 ; n17211_not
g67326 not n54120 ; n54120_not
g67327 not n28011 ; n28011_not
g67328 not n32412 ; n32412_not
g67329 not n54111 ; n54111_not
g67330 not n27030 ; n27030_not
g67331 not n38001 ; n38001_not
g67332 not n11541 ; n11541_not
g67333 not n31134 ; n31134_not
g67334 not n10380 ; n10380_not
g67335 not n11532 ; n11532_not
g67336 not n32025 ; n32025_not
g67337 not n32016 ; n32016_not
g67338 not n42015 ; n42015_not
g67339 not n51213 ; n51213_not
g67340 not n46200 ; n46200_not
g67341 not n50502 ; n50502_not
g67342 not n11703 ; n11703_not
g67343 not n40260 ; n40260_not
g67344 not n31143 ; n31143_not
g67345 not n11712 ; n11712_not
g67346 not n42240 ; n42240_not
g67347 not n42024 ; n42024_not
g67348 not n11721 ; n11721_not
g67349 not n32403 ; n32403_not
g67350 not n11730 ; n11730_not
g67351 not n51411 ; n51411_not
g67352 not n42303 ; n42303_not
g67353 not n32034 ; n32034_not
g67354 not n19200 ; n19200_not
g67355 not n31107 ; n31107_not
g67356 not n32430 ; n32430_not
g67357 not n17112 ; n17112_not
g67358 not n50151 ; n50151_not
g67359 not n40242 ; n40242_not
g67360 not n52131 ; n52131_not
g67361 not n31620 ; n31620_not
g67362 not n47010 ; n47010_not
g67363 not n42051 ; n42051_not
g67364 not n32421 ; n32421_not
g67365 not n51222 ; n51222_not
g67366 not n28020 ; n28020_not
g67367 not n11523 ; n11523_not
g67368 not n42042 ; n42042_not
g67369 not n18111 ; n18111_not
g67370 not n31125 ; n31125_not
g67371 not n40143 ; n40143_not
g67372 not n11802 ; n11802_not
g67373 not n11811 ; n11811_not
g67374 not n52140 ; n52140_not
g67375 not n31116 ; n31116_not
g67376 not n11820 ; n11820_not
g67377 not n11550 ; n11550_not
g67378 not n26121 ; n26121_not
g67379 not n17031 ; n17031_not
g67380 not n19020 ; n19020_not
g67381 not n25500 ; n25500_not
g67382 not n11631 ; n11631_not
g67383 not n41700 ; n41700_not
g67384 not n35310 ; n35310_not
g67385 not n31161 ; n31161_not
g67386 not n10902 ; n10902_not
g67387 not n11640 ; n11640_not
g67388 not n28200 ; n28200_not
g67389 not n17004 ; n17004_not
g67390 not n51204 ; n51204_not
g67391 not n31152 ; n31152_not
g67392 not n31701 ; n31701_not
g67393 not n19110 ; n19110_not
g67394 not n47001 ; n47001_not
g67395 not n40233 ; n40233_not
g67396 not n26130 ; n26130_not
g67397 not n11613 ; n11613_not
g67398 not n50007 ; n50007_not
g67399 not n51114 ; n51114_not
g67400 not n23322 ; n23322_not
g67401 not n23160 ; n23160_not
g67402 not n23052 ; n23052_not
g67403 not n23250 ; n23250_not
g67404 not n23241 ; n23241_not
g67405 not n23232 ; n23232_not
g67406 not n23223 ; n23223_not
g67407 not n42420 ; n42420_not
g67408 not n23331 ; n23331_not
g67409 not n44121 ; n44121_not
g67410 not n23610 ; n23610_not
g67411 not n23313 ; n23313_not
g67412 not n12711 ; n12711_not
g67413 not n44112 ; n44112_not
g67414 not n16500 ; n16500_not
g67415 not n23304 ; n23304_not
g67416 not n20073 ; n20073_not
g67417 not n30720 ; n30720_not
g67418 not n23142 ; n23142_not
g67419 not n23151 ; n23151_not
g67420 not n13134 ; n13134_not
g67421 not n30621 ; n30621_not
g67422 not n40800 ; n40800_not
g67423 not n23340 ; n23340_not
g67424 not n42222 ; n42222_not
g67425 not n31602 ; n31602_not
g67426 not n23214 ; n23214_not
g67427 not n23205 ; n23205_not
g67428 not n51042 ; n51042_not
g67429 not n12702 ; n12702_not
g67430 not n30630 ; n30630_not
g67431 not n27300 ; n27300_not
g67432 not n20055 ; n20055_not
g67433 not n30612 ; n30612_not
g67434 not n31521 ; n31521_not
g67435 not n23430 ; n23430_not
g67436 not n20046 ; n20046_not
g67437 not n26301 ; n26301_not
g67438 not n23421 ; n23421_not
g67439 not n23412 ; n23412_not
g67440 not n44103 ; n44103_not
g67441 not n12603 ; n12603_not
g67442 not n23520 ; n23520_not
g67443 not n23511 ; n23511_not
g67444 not n23502 ; n23502_not
g67445 not n30603 ; n30603_not
g67446 not n27210 ; n27210_not
g67447 not n32043 ; n32043_not
g67448 not n12612 ; n12612_not
g67449 not n37200 ; n37200_not
g67450 not n26400 ; n26400_not
g67451 not n56010 ; n56010_not
g67452 not n20064 ; n20064_not
g67453 not n40053 ; n40053_not
g67454 not n40008 ; n40008_not
g67455 not n52401 ; n52401_not
g67456 not n23007 ; n23007_not
g67457 not n23403 ; n23403_not
g67458 not n44130 ; n44130_not
g67459 not n40062 ; n40062_not
g67460 not n30531 ; n30531_not
g67461 not n50601 ; n50601_not
g67462 not n42204 ; n42204_not
g67463 not n52320 ; n52320_not
g67464 not n20037 ; n20037_not
g67465 not n27120 ; n27120_not
g67466 not n34410 ; n34410_not
g67467 not n34500 ; n34500_not
g67468 not n50106 ; n50106_not
g67469 not n45120 ; n45120_not
g67470 not n47100 ; n47100_not
g67471 not n41331 ; n41331_not
g67472 not n35211 ; n35211_not
g67473 not n40026 ; n40026_not
g67474 not n30801 ; n30801_not
g67475 not n50034 ; n50034_not
g67476 not n40035 ; n40035_not
g67477 not n46011 ; n46011_not
g67478 not n31530 ; n31530_not
g67479 not n20091 ; n20091_not
g67480 not n46020 ; n46020_not
g67481 not n42213 ; n42213_not
g67482 not n13215 ; n13215_not
g67483 not n42402 ; n42402_not
g67484 not n52410 ; n52410_not
g67485 not n46002 ; n46002_not
g67486 not n40044 ; n40044_not
g67487 not n52050 ; n52050_not
g67488 not n12621 ; n12621_not
g67489 not n52041 ; n52041_not
g67490 not n50241 ; n50241_not
g67491 not n50016 ; n50016_not
g67492 not n23133 ; n23133_not
g67493 not n40017 ; n40017_not
g67494 not n23124 ; n23124_not
g67495 not n50025 ; n50025_not
g67496 not n20082 ; n20082_not
g67497 not n26310 ; n26310_not
g67498 not n13170 ; n13170_not
g67499 not n41224 ; n41224_not
g67500 not n44140 ; n44140_not
g67501 not n31333 ; n31333_not
g67502 not n44131 ; n44131_not
g67503 not n18112 ; n18112_not
g67504 not n25510 ; n25510_not
g67505 not n15511 ; n15511_not
g67506 not n31621 ; n31621_not
g67507 not n10345 ; n10345_not
g67508 not n18211 ; n18211_not
g67509 not n37021 ; n37021_not
g67510 not n41440 ; n41440_not
g67511 not n50413 ; n50413_not
g67512 not n21505 ; n21505_not
g67513 not n35203 ; n35203_not
g67514 not n10840 ; n10840_not
g67515 not n40306 ; n40306_not
g67516 not n21541 ; n21541_not
g67517 not n21109 ; n21109_not
g67518 not n40351 ; n40351_not
g67519 not n52600 ; n52600_not
g67520 not n32026 ; n32026_not
g67521 not n21631 ; n21631_not
g67522 not n37210 ; n37210_not
g67523 not n10912 ; n10912_not
g67524 not n40270 ; n40270_not
g67525 not n31531 ; n31531_not
g67526 not n35212 ; n35212_not
g67527 not n26140 ; n26140_not
g67528 not n32215 ; n32215_not
g67529 not n14026 ; n14026_not
g67530 not n10327 ; n10327_not
g67531 not n18400 ; n18400_not
g67532 not n53122 ; n53122_not
g67533 not n26131 ; n26131_not
g67534 not n28111 ; n28111_not
g67535 not n10381 ; n10381_not
g67536 not n45004 ; n45004_not
g67537 not n28102 ; n28102_not
g67538 not n44122 ; n44122_not
g67539 not n31360 ; n31360_not
g67540 not n42151 ; n42151_not
g67541 not n10318 ; n10318_not
g67542 not n15142 ; n15142_not
g67543 not n10264 ; n10264_not
g67544 not n14035 ; n14035_not
g67545 not n42124 ; n42124_not
g67546 not n18220 ; n18220_not
g67547 not n21640 ; n21640_not
g67548 not n43150 ; n43150_not
g67549 not n31630 ; n31630_not
g67550 not n51142 ; n51142_not
g67551 not n10273 ; n10273_not
g67552 not n17311 ; n17311_not
g67553 not n21532 ; n21532_not
g67554 not n25420 ; n25420_not
g67555 not n20452 ; n20452_not
g67556 not n30172 ; n30172_not
g67557 not n30217 ; n30217_not
g67558 not n35302 ; n35302_not
g67559 not n41233 ; n41233_not
g67560 not n26302 ; n26302_not
g67561 not n10831 ; n10831_not
g67562 not n17122 ; n17122_not
g67563 not n26311 ; n26311_not
g67564 not n25600 ; n25600_not
g67565 not n42241 ; n42241_not
g67566 not n21514 ; n21514_not
g67567 not n18202 ; n18202_not
g67568 not n31342 ; n31342_not
g67569 not n40333 ; n40333_not
g67570 not n42223 ; n42223_not
g67571 not n10309 ; n10309_not
g67572 not n42007 ; n42007_not
g67573 not n30163 ; n30163_not
g67574 not n21613 ; n21613_not
g67575 not n42700 ; n42700_not
g67576 not n10804 ; n10804_not
g67577 not n30280 ; n30280_not
g67578 not n10291 ; n10291_not
g67579 not n40243 ; n40243_not
g67580 not n17302 ; n17302_not
g67581 not n15322 ; n15322_not
g67582 not n32053 ; n32053_not
g67583 not n35320 ; n35320_not
g67584 not n20470 ; n20470_not
g67585 not n30190 ; n30190_not
g67586 not n53104 ; n53104_not
g67587 not n30181 ; n30181_not
g67588 not n10813 ; n10813_not
g67589 not n32206 ; n32206_not
g67590 not n21118 ; n21118_not
g67591 not n33106 ; n33106_not
g67592 not n42610 ; n42610_not
g67593 not n47101 ; n47101_not
g67594 not n51151 ; n51151_not
g67595 not n40324 ; n40324_not
g67596 not n51160 ; n51160_not
g67597 not n21604 ; n21604_not
g67598 not n46201 ; n46201_not
g67599 not n33142 ; n33142_not
g67600 not n50206 ; n50206_not
g67601 not n33160 ; n33160_not
g67602 not n14008 ; n14008_not
g67603 not n42133 ; n42133_not
g67604 not n33403 ; n33403_not
g67605 not n10372 ; n10372_not
g67606 not n51322 ; n51322_not
g67607 not n33007 ; n33007_not
g67608 not n53113 ; n53113_not
g67609 not n21127 ; n21127_not
g67610 not n10282 ; n10282_not
g67611 not n33070 ; n33070_not
g67612 not n53320 ; n53320_not
g67613 not n53032 ; n53032_not
g67614 not n33133 ; n33133_not
g67615 not n31540 ; n31540_not
g67616 not n25501 ; n25501_not
g67617 not n15313 ; n15313_not
g67618 not n42142 ; n42142_not
g67619 not n37201 ; n37201_not
g67620 not n20461 ; n20461_not
g67621 not n21550 ; n21550_not
g67622 not n10822 ; n10822_not
g67623 not n40342 ; n40342_not
g67624 not n18103 ; n18103_not
g67625 not n15115 ; n15115_not
g67626 not n31207 ; n31207_not
g67627 not n21622 ; n21622_not
g67628 not n40234 ; n40234_not
g67629 not n21523 ; n21523_not
g67630 not n15430 ; n15430_not
g67631 not n40315 ; n40315_not
g67632 not n33340 ; n33340_not
g67633 not n31351 ; n31351_not
g67634 not n14017 ; n14017_not
g67635 not n53410 ; n53410_not
g67636 not n15124 ; n15124_not
g67637 not n33421 ; n33421_not
g67638 not n51430 ; n51430_not
g67639 not n44041 ; n44041_not
g67640 not n17212 ; n17212_not
g67641 not n21721 ; n21721_not
g67642 not n14143 ; n14143_not
g67643 not n51421 ; n51421_not
g67644 not n51601 ; n51601_not
g67645 not n15133 ; n15133_not
g67646 not n14152 ; n14152_not
g67647 not n44032 ; n44032_not
g67648 not n35500 ; n35500_not
g67649 not n41512 ; n41512_not
g67650 not n42250 ; n42250_not
g67651 not n14161 ; n14161_not
g67652 not n21730 ; n21730_not
g67653 not n54310 ; n54310_not
g67654 not n43222 ; n43222_not
g67655 not n15205 ; n15205_not
g67656 not n30154 ; n30154_not
g67657 not n20434 ; n20434_not
g67658 not n31900 ; n31900_not
g67659 not n14107 ; n14107_not
g67660 not n11056 ; n11056_not
g67661 not n11065 ; n11065_not
g67662 not n14116 ; n14116_not
g67663 not n44050 ; n44050_not
g67664 not n32710 ; n32710_not
g67665 not n31441 ; n31441_not
g67666 not n15232 ; n15232_not
g67667 not n26320 ; n26320_not
g67668 not n21055 ; n21055_not
g67669 not n14125 ; n14125_not
g67670 not n40630 ; n40630_not
g67671 not n39100 ; n39100_not
g67672 not n21424 ; n21424_not
g67673 not n14134 ; n14134_not
g67674 not n50260 ; n50260_not
g67675 not n41413 ; n41413_not
g67676 not n42205 ; n42205_not
g67677 not n11137 ; n11137_not
g67678 not n20614 ; n20614_not
g67679 not n44005 ; n44005_not
g67680 not n14431 ; n14431_not
g67681 not n14206 ; n14206_not
g67682 not n46012 ; n46012_not
g67683 not n44014 ; n44014_not
g67684 not n46003 ; n46003_not
g67685 not n53005 ; n53005_not
g67686 not n11146 ; n11146_not
g67687 not n25321 ; n25321_not
g67688 not n14215 ; n14215_not
g67689 not n14422 ; n14422_not
g67690 not n42214 ; n42214_not
g67691 not n11155 ; n11155_not
g67692 not n54301 ; n54301_not
g67693 not n14224 ; n14224_not
g67694 not n15223 ; n15223_not
g67695 not n11164 ; n11164_not
g67696 not n21037 ; n21037_not
g67697 not n20623 ; n20623_not
g67698 not n14233 ; n14233_not
g67699 not n11173 ; n11173_not
g67700 not n33412 ; n33412_not
g67701 not n14170 ; n14170_not
g67702 not n11038 ; n11038_not
g67703 not n51412 ; n51412_not
g67704 not n44023 ; n44023_not
g67705 not n51403 ; n51403_not
g67706 not n21415 ; n21415_not
g67707 not n50512 ; n50512_not
g67708 not n20425 ; n20425_not
g67709 not n11119 ; n11119_not
g67710 not n11029 ; n11029_not
g67711 not n41521 ; n41521_not
g67712 not n43141 ; n43141_not
g67713 not n30136 ; n30136_not
g67714 not n51340 ; n51340_not
g67715 not n54040 ; n54040_not
g67716 not n11128 ; n11128_not
g67717 not n21046 ; n21046_not
g67718 not n26500 ; n26500_not
g67719 not n15214 ; n15214_not
g67720 not n50422 ; n50422_not
g67721 not n17203 ; n17203_not
g67722 not n15340 ; n15340_not
g67723 not n25330 ; n25330_not
g67724 not n21091 ; n21091_not
g67725 not n32224 ; n32224_not
g67726 not n30208 ; n30208_not
g67727 not n40225 ; n40225_not
g67728 not n44104 ; n44104_not
g67729 not n51331 ; n51331_not
g67730 not n20650 ; n20650_not
g67731 not n33115 ; n33115_not
g67732 not n20443 ; n20443_not
g67733 not n45310 ; n45310_not
g67734 not n42601 ; n42601_not
g67735 not n15160 ; n15160_not
g67736 not n21082 ; n21082_not
g67737 not n32035 ; n32035_not
g67738 not n53131 ; n53131_not
g67739 not n50161 ; n50161_not
g67740 not n37030 ; n37030_not
g67741 not n18121 ; n18121_not
g67742 not n15241 ; n15241_not
g67743 not n40360 ; n40360_not
g67744 not n26122 ; n26122_not
g67745 not n21460 ; n21460_not
g67746 not n10930 ; n10930_not
g67747 not n31324 ; n31324_not
g67748 not n53311 ; n53311_not
g67749 not n46030 ; n46030_not
g67750 not n44113 ; n44113_not
g67751 not n38101 ; n38101_not
g67752 not n18130 ; n18130_not
g67753 not n33124 ; n33124_not
g67754 not n20632 ; n20632_not
g67755 not n53023 ; n53023_not
g67756 not n42160 ; n42160_not
g67757 not n14071 ; n14071_not
g67758 not n18301 ; n18301_not
g67759 not n51610 ; n51610_not
g67760 not n17221 ; n17221_not
g67761 not n53014 ; n53014_not
g67762 not n18310 ; n18310_not
g67763 not n14080 ; n14080_not
g67764 not n33430 ; n33430_not
g67765 not n41503 ; n41503_not
g67766 not n21064 ; n21064_not
g67767 not n53140 ; n53140_not
g67768 not n11047 ; n11047_not
g67769 not n32233 ; n32233_not
g67770 not n20605 ; n20605_not
g67771 not n21703 ; n21703_not
g67772 not n46021 ; n46021_not
g67773 not n57010 ; n57010_not
g67774 not n31306 ; n31306_not
g67775 not n10525 ; n10525_not
g67776 not n40405 ; n40405_not
g67777 not n21433 ; n21433_not
g67778 not n28003 ; n28003_not
g67779 not n21712 ; n21712_not
g67780 not n28030 ; n28030_not
g67781 not n26401 ; n26401_not
g67782 not n46210 ; n46210_not
g67783 not n14521 ; n14521_not
g67784 not n14044 ; n14044_not
g67785 not n31315 ; n31315_not
g67786 not n21028 ; n21028_not
g67787 not n28021 ; n28021_not
g67788 not n26410 ; n26410_not
g67789 not n14053 ; n14053_not
g67790 not n14512 ; n14512_not
g67791 not n17230 ; n17230_not
g67792 not n25411 ; n25411_not
g67793 not n15502 ; n15502_not
g67794 not n14062 ; n14062_not
g67795 not n21073 ; n21073_not
g67796 not n15331 ; n15331_not
g67797 not n35230 ; n35230_not
g67798 not n33601 ; n33601_not
g67799 not n10129 ; n10129_not
g67800 not n20524 ; n20524_not
g67801 not n21334 ; n21334_not
g67802 not n32116 ; n32116_not
g67803 not n32080 ; n32080_not
g67804 not n40117 ; n40117_not
g67805 not n42106 ; n42106_not
g67806 not n35401 ; n35401_not
g67807 not n43015 ; n43015_not
g67808 not n31513 ; n31513_not
g67809 not n40072 ; n40072_not
g67810 not n33610 ; n33610_not
g67811 not n10093 ; n10093_not
g67812 not n10507 ; n10507_not
g67813 not n10516 ; n10516_not
g67814 not n32125 ; n32125_not
g67815 not n45202 ; n45202_not
g67816 not n31450 ; n31450_not
g67817 not n10534 ; n10534_not
g67818 not n26212 ; n26212_not
g67819 not n10156 ; n10156_not
g67820 not n14260 ; n14260_not
g67821 not n43006 ; n43006_not
g67822 not n33034 ; n33034_not
g67823 not n32071 ; n32071_not
g67824 not n10444 ; n10444_not
g67825 not n10147 ; n10147_not
g67826 not n30082 ; n30082_not
g67827 not n32107 ; n32107_not
g67828 not n14251 ; n14251_not
g67829 not n51313 ; n51313_not
g67830 not n21208 ; n21208_not
g67831 not n42115 ; n42115_not
g67832 not n46102 ; n46102_not
g67833 not n10138 ; n10138_not
g67834 not n52420 ; n52420_not
g67835 not n21325 ; n21325_not
g67836 not n33043 ; n33043_not
g67837 not n33304 ; n33304_not
g67838 not n37300 ; n37300_not
g67839 not n10462 ; n10462_not
g67840 not n10471 ; n10471_not
g67841 not n14242 ; n14242_not
g67842 not n15007 ; n15007_not
g67843 not n50152 ; n50152_not
g67844 not n50323 ; n50323_not
g67845 not n40135 ; n40135_not
g67846 not n21370 ; n21370_not
g67847 not n51520 ; n51520_not
g67848 not n10075 ; n10075_not
g67849 not n17410 ; n17410_not
g67850 not n31405 ; n31405_not
g67851 not n10057 ; n10057_not
g67852 not n51700 ; n51700_not
g67853 not n32134 ; n32134_not
g67854 not n42511 ; n42511_not
g67855 not n40144 ; n40144_not
g67856 not n15025 ; n15025_not
g67857 not n10570 ; n10570_not
g67858 not n43024 ; n43024_not
g67859 not n21190 ; n21190_not
g67860 not n46120 ; n46120_not
g67861 not n10066 ; n10066_not
g67862 not n42232 ; n42232_not
g67863 not n44302 ; n44302_not
g67864 not n17401 ; n17401_not
g67865 not n46111 ; n46111_not
g67866 not n21352 ; n21352_not
g67867 not n33520 ; n33520_not
g67868 not n10543 ; n10543_not
g67869 not n15250 ; n15250_not
g67870 not n33313 ; n33313_not
g67871 not n40081 ; n40081_not
g67872 not n10039 ; n10039_not
g67873 not n10084 ; n10084_not
g67874 not n10552 ; n10552_not
g67875 not n50530 ; n50530_not
g67876 not n30244 ; n30244_not
g67877 not n10048 ; n10048_not
g67878 not n14440 ; n14440_not
g67879 not n20533 ; n20533_not
g67880 not n31801 ; n31801_not
g67881 not n20542 ; n20542_not
g67882 not n33052 ; n33052_not
g67883 not n10561 ; n10561_not
g67884 not n10246 ; n10246_not
g67885 not n14323 ; n14323_not
g67886 not n48001 ; n48001_not
g67887 not n42070 ; n42070_not
g67888 not n18022 ; n18022_not
g67889 not n17500 ; n17500_not
g67890 not n18004 ; n18004_not
g67891 not n26041 ; n26041_not
g67892 not n21262 ; n21262_not
g67893 not n51304 ; n51304_not
g67894 not n14314 ; n14314_not
g67895 not n10237 ; n10237_not
g67896 not n10354 ; n10354_not
g67897 not n15520 ; n15520_not
g67898 not n26023 ; n26023_not
g67899 not n10228 ; n10228_not
g67900 not n33241 ; n33241_not
g67901 not n25240 ; n25240_not
g67902 not n43105 ; n43105_not
g67903 not n26230 ; n26230_not
g67904 not n42061 ; n42061_not
g67905 not n14305 ; n14305_not
g67906 not n45211 ; n45211_not
g67907 not n54031 ; n54031_not
g67908 not n33223 ; n33223_not
g67909 not n26050 ; n26050_not
g67910 not n18013 ; n18013_not
g67911 not n30262 ; n30262_not
g67912 not n10255 ; n10255_not
g67913 not n21244 ; n21244_not
g67914 not n14332 ; n14332_not
g67915 not n17014 ; n17014_not
g67916 not n25231 ; n25231_not
g67917 not n21235 ; n21235_not
g67918 not n41260 ; n41260_not
g67919 not n14350 ; n14350_not
g67920 not n33232 ; n33232_not
g67921 not n26032 ; n26032_not
g67922 not n42043 ; n42043_not
g67923 not n17032 ; n17032_not
g67924 not n33061 ; n33061_not
g67925 not n30253 ; n30253_not
g67926 not n20560 ; n20560_not
g67927 not n26014 ; n26014_not
g67928 not n43240 ; n43240_not
g67929 not n45031 ; n45031_not
g67930 not n26005 ; n26005_not
g67931 not n10183 ; n10183_not
g67932 not n26104 ; n26104_not
g67933 not n18040 ; n18040_not
g67934 not n10174 ; n10174_not
g67935 not n32008 ; n32008_not
g67936 not n21217 ; n21217_not
g67937 not n55030 ; n55030_not
g67938 not n10417 ; n10417_not
g67939 not n21307 ; n21307_not
g67940 not n33205 ; n33205_not
g67941 not n10426 ; n10426_not
g67942 not n10165 ; n10165_not
g67943 not n33214 ; n33214_not
g67944 not n42520 ; n42520_not
g67945 not n15304 ; n15304_not
g67946 not n10219 ; n10219_not
g67947 not n21280 ; n21280_not
g67948 not n18031 ; n18031_not
g67949 not n50341 ; n50341_not
g67950 not n21226 ; n21226_not
g67951 not n42052 ; n42052_not
g67952 not n31612 ; n31612_not
g67953 not n26221 ; n26221_not
g67954 not n20515 ; n20515_not
g67955 not n33250 ; n33250_not
g67956 not n17023 ; n17023_not
g67957 not n40090 ; n40090_not
g67958 not n10192 ; n10192_not
g67959 not n28210 ; n28210_not
g67960 not n10705 ; n10705_not
g67961 not n41242 ; n41242_not
g67962 not n55003 ; n55003_not
g67963 not n51214 ; n51214_not
g67964 not n43060 ; n43060_not
g67965 not n44212 ; n44212_not
g67966 not n21154 ; n21154_not
g67967 not n10714 ; n10714_not
g67968 not n56011 ; n56011_not
g67969 not n17104 ; n17104_not
g67970 not n50305 ; n50305_not
g67971 not n10723 ; n10723_not
g67972 not n21019 ; n21019_not
g67973 not n51205 ; n51205_not
g67974 not n15412 ; n15412_not
g67975 not n44221 ; n44221_not
g67976 not n54121 ; n54121_not
g67977 not n53401 ; n53401_not
g67978 not n30235 ; n30235_not
g67979 not n50521 ; n50521_not
g67980 not n32800 ; n32800_not
g67981 not n40207 ; n40207_not
g67982 not n10435 ; n10435_not
g67983 not n15403 ; n15403_not
g67984 not n15070 ; n15070_not
g67985 not n52510 ; n52510_not
g67986 not n53041 ; n53041_not
g67987 not n32170 ; n32170_not
g67988 not n15421 ; n15421_not
g67989 not n45013 ; n45013_not
g67990 not n40252 ; n40252_not
g67991 not n23611 ; n23611_not
g67992 not n51502 ; n51502_not
g67993 not n17113 ; n17113_not
g67994 not n33151 ; n33151_not
g67995 not n50404 ; n50404_not
g67996 not n21136 ; n21136_not
g67997 not n10390 ; n10390_not
g67998 not n30226 ; n30226_not
g67999 not n17320 ; n17320_not
g68000 not n54022 ; n54022_not
g68001 not n35221 ; n35221_not
g68002 not n31504 ; n31504_not
g68003 not n14530 ; n14530_not
g68004 not n10732 ; n10732_not
g68005 not n41305 ; n41305_not
g68006 not n39010 ; n39010_not
g68007 not n50350 ; n50350_not
g68008 not n30109 ; n30109_not
g68009 not n21145 ; n21145_not
g68010 not n10741 ; n10741_not
g68011 not n45040 ; n45040_not
g68012 not n44203 ; n44203_not
g68013 not n35311 ; n35311_not
g68014 not n10750 ; n10750_not
g68015 not n42016 ; n42016_not
g68016 not n31603 ; n31603_not
g68017 not n43231 ; n43231_not
g68018 not n35410 ; n35410_not
g68019 not n10615 ; n10615_not
g68020 not n55012 ; n55012_not
g68021 not n51511 ; n51511_not
g68022 not n31414 ; n31414_not
g68023 not n10624 ; n10624_not
g68024 not n51241 ; n51241_not
g68025 not n10633 ; n10633_not
g68026 not n31162 ; n31162_not
g68027 not n43042 ; n43042_not
g68028 not n32152 ; n32152_not
g68029 not n53050 ; n53050_not
g68030 not n33016 ; n33016_not
g68031 not n15034 ; n15034_not
g68032 not n31423 ; n31423_not
g68033 not n40162 ; n40162_not
g68034 not n51250 ; n51250_not
g68035 not n21181 ; n21181_not
g68036 not n44311 ; n44311_not
g68037 not n33511 ; n33511_not
g68038 not n43033 ; n43033_not
g68039 not n10480 ; n10480_not
g68040 not n10606 ; n10606_not
g68041 not n32143 ; n32143_not
g68042 not n33502 ; n33502_not
g68043 not n30307 ; n30307_not
g68044 not n10660 ; n10660_not
g68045 not n21442 ; n21442_not
g68046 not n51223 ; n51223_not
g68047 not n32044 ; n32044_not
g68048 not n32161 ; n32161_not
g68049 not n44320 ; n44320_not
g68050 not n21163 ; n21163_not
g68051 not n44401 ; n44401_not
g68052 not n45022 ; n45022_not
g68053 not n56002 ; n56002_not
g68054 not n43051 ; n43051_not
g68055 not n43132 ; n43132_not
g68056 not n40180 ; n40180_not
g68057 not n51232 ; n51232_not
g68058 not n15052 ; n15052_not
g68059 not n10642 ; n10642_not
g68060 not n30091 ; n30091_not
g68061 not n31522 ; n31522_not
g68062 not n21172 ; n21172_not
g68063 not n44230 ; n44230_not
g68064 not n10651 ; n10651_not
g68065 not n28300 ; n28300_not
g68066 not n20830 ; n20830_not
g68067 not n32530 ; n32530_not
g68068 not n23323 ; n23323_not
g68069 not n12442 ; n12442_not
g68070 not n24106 ; n24106_not
g68071 not n32305 ; n32305_not
g68072 not n29110 ; n29110_not
g68073 not n13153 ; n13153_not
g68074 not n12433 ; n12433_not
g68075 not n13702 ; n13702_not
g68076 not n12037 ; n12037_not
g68077 not n23332 ; n23332_not
g68078 not n42340 ; n42340_not
g68079 not n36310 ; n36310_not
g68080 not n23170 ; n23170_not
g68081 not n40441 ; n40441_not
g68082 not n30712 ; n30712_not
g68083 not n50062 ; n50062_not
g68084 not n30505 ; n30505_not
g68085 not n12460 ; n12460_not
g68086 not n23305 ; n23305_not
g68087 not n13162 ; n13162_not
g68088 not n40450 ; n40450_not
g68089 not n23314 ; n23314_not
g68090 not n12451 ; n12451_not
g68091 not n34204 ; n34204_not
g68092 not n12028 ; n12028_not
g68093 not n20236 ; n20236_not
g68094 not n30703 ; n30703_not
g68095 not n23044 ; n23044_not
g68096 not n23350 ; n23350_not
g68097 not n23161 ; n23161_not
g68098 not n38110 ; n38110_not
g68099 not n22540 ; n22540_not
g68100 not n24133 ; n24133_not
g68101 not n53203 ; n53203_not
g68102 not n24142 ; n24142_not
g68103 not n22531 ; n22531_not
g68104 not n13315 ; n13315_not
g68105 not n32521 ; n32521_not
g68106 not n16420 ; n16420_not
g68107 not n22171 ; n22171_not
g68108 not n24151 ; n24151_not
g68109 not n13126 ; n13126_not
g68110 not n24115 ; n24115_not
g68111 not n50710 ; n50710_not
g68112 not n13135 ; n13135_not
g68113 not n12424 ; n12424_not
g68114 not n12046 ; n12046_not
g68115 not n20245 ; n20245_not
g68116 not n23341 ; n23341_not
g68117 not n13711 ; n13711_not
g68118 not n20074 ; n20074_not
g68119 not n12415 ; n12415_not
g68120 not n50116 ; n50116_not
g68121 not n22162 ; n22162_not
g68122 not n56101 ; n56101_not
g68123 not n24124 ; n24124_not
g68124 not n29101 ; n29101_not
g68125 not n12406 ; n12406_not
g68126 not n30325 ; n30325_not
g68127 not n24007 ; n24007_not
g68128 not n43114 ; n43114_not
g68129 not n20740 ; n20740_not
g68130 not n22621 ; n22621_not
g68131 not n23233 ; n23233_not
g68132 not n20821 ; n20821_not
g68133 not n12523 ; n12523_not
g68134 not n24016 ; n24016_not
g68135 not n34420 ; n34420_not
g68136 not n34231 ; n34231_not
g68137 not n12820 ; n12820_not
g68138 not n12514 ; n12514_not
g68139 not n22612 ; n22612_not
g68140 not n23242 ; n23242_not
g68141 not n23206 ; n23206_not
g68142 not n13108 ; n13108_not
g68143 not n13621 ; n13621_not
g68144 not n30352 ; n30352_not
g68145 not n12550 ; n12550_not
g68146 not n34240 ; n34240_not
g68147 not n23215 ; n23215_not
g68148 not n20218 ; n20218_not
g68149 not n22630 ; n22630_not
g68150 not n27202 ; n27202_not
g68151 not n12541 ; n12541_not
g68152 not n22117 ; n22117_not
g68153 not n13630 ; n13630_not
g68154 not n23224 ; n23224_not
g68155 not n45400 ; n45400_not
g68156 not n16204 ; n16204_not
g68157 not n50107 ; n50107_not
g68158 not n40414 ; n40414_not
g68159 not n19111 ; n19111_not
g68160 not n24052 ; n24052_not
g68161 not n40423 ; n40423_not
g68162 not n54211 ; n54211_not
g68163 not n24061 ; n24061_not
g68164 not n30721 ; n30721_not
g68165 not n40432 ; n40432_not
g68166 not n24070 ; n24070_not
g68167 not n34213 ; n34213_not
g68168 not n13171 ; n13171_not
g68169 not n22126 ; n22126_not
g68170 not n24025 ; n24025_not
g68171 not n12505 ; n12505_not
g68172 not n22603 ; n22603_not
g68173 not n22135 ; n22135_not
g68174 not n20227 ; n20227_not
g68175 not n23251 ; n23251_not
g68176 not n36301 ; n36301_not
g68177 not n24034 ; n24034_not
g68178 not n34222 ; n34222_not
g68179 not n19102 ; n19102_not
g68180 not n23260 ; n23260_not
g68181 not n24043 ; n24043_not
g68182 not n13117 ; n13117_not
g68183 not n40702 ; n40702_not
g68184 not n23062 ; n23062_not
g68185 not n51043 ; n51043_not
g68186 not n24250 ; n24250_not
g68187 not n22423 ; n22423_not
g68188 not n42313 ; n42313_not
g68189 not n29020 ; n29020_not
g68190 not n23008 ; n23008_not
g68191 not n41350 ; n41350_not
g68192 not n37111 ; n37111_not
g68193 not n53212 ; n53212_not
g68194 not n15700 ; n15700_not
g68195 not n12118 ; n12118_not
g68196 not n22414 ; n22414_not
g68197 not n20281 ; n20281_not
g68198 not n34132 ; n34132_not
g68199 not n16105 ; n16105_not
g68200 not n22441 ; n22441_not
g68201 not n12316 ; n12316_not
g68202 not n22225 ; n22225_not
g68203 not n24232 ; n24232_not
g68204 not n42322 ; n42322_not
g68205 not n50611 ; n50611_not
g68206 not n16132 ; n16132_not
g68207 not n12307 ; n12307_not
g68208 not n34141 ; n34141_not
g68209 not n22432 ; n22432_not
g68210 not n34123 ; n34123_not
g68211 not n32314 ; n32314_not
g68212 not n19201 ; n19201_not
g68213 not n24241 ; n24241_not
g68214 not n13144 ; n13144_not
g68215 not n45112 ; n45112_not
g68216 not n55210 ; n55210_not
g68217 not n23521 ; n23521_not
g68218 not n36004 ; n36004_not
g68219 not n24304 ; n24304_not
g68220 not n22252 ; n22252_not
g68221 not n12253 ; n12253_not
g68222 not n47200 ; n47200_not
g68223 not n23530 ; n23530_not
g68224 not n12244 ; n12244_not
g68225 not n24313 ; n24313_not
g68226 not n12235 ; n12235_not
g68227 not n24322 ; n24322_not
g68228 not n20290 ; n20290_not
g68229 not n24331 ; n24331_not
g68230 not n41251 ; n41251_not
g68231 not n12226 ; n12226_not
g68232 not n12280 ; n12280_not
g68233 not n32503 ; n32503_not
g68234 not n40603 ; n40603_not
g68235 not n30550 ; n30550_not
g68236 not n22405 ; n22405_not
g68237 not n32323 ; n32323_not
g68238 not n16123 ; n16123_not
g68239 not n23503 ; n23503_not
g68240 not n12271 ; n12271_not
g68241 not n40612 ; n40612_not
g68242 not n12127 ; n12127_not
g68243 not n23134 ; n23134_not
g68244 not n23512 ; n23512_not
g68245 not n40621 ; n40621_not
g68246 not n12262 ; n12262_not
g68247 not n12136 ; n12136_not
g68248 not n16150 ; n16150_not
g68249 not n22504 ; n22504_not
g68250 not n30910 ; n30910_not
g68251 not n40513 ; n40513_not
g68252 not n12370 ; n12370_not
g68253 not n12073 ; n12073_not
g68254 not n23404 ; n23404_not
g68255 not n40522 ; n40522_not
g68256 not n12361 ; n12361_not
g68257 not n42430 ; n42430_not
g68258 not n23413 ; n23413_not
g68259 not n41710 ; n41710_not
g68260 not n27121 ; n27121_not
g68261 not n40531 ; n40531_not
g68262 not n22522 ; n22522_not
g68263 not n30901 ; n30901_not
g68264 not n22180 ; n22180_not
g68265 not n41701 ; n41701_not
g68266 not n23152 ; n23152_not
g68267 not n36121 ; n36121_not
g68268 not n40504 ; n40504_not
g68269 not n24160 ; n24160_not
g68270 not n22513 ; n22513_not
g68271 not n40711 ; n40711_not
g68272 not n20254 ; n20254_not
g68273 not n23053 ; n23053_not
g68274 not n50701 ; n50701_not
g68275 not n12334 ; n12334_not
g68276 not n34150 ; n34150_not
g68277 not n23440 ; n23440_not
g68278 not n30343 ; n30343_not
g68279 not n36103 ; n36103_not
g68280 not n12325 ; n12325_not
g68281 not n22450 ; n22450_not
g68282 not n24223 ; n24223_not
g68283 not n13801 ; n13801_not
g68284 not n22216 ; n22216_not
g68285 not n32512 ; n32512_not
g68286 not n40540 ; n40540_not
g68287 not n20272 ; n20272_not
g68288 not n54220 ; n54220_not
g68289 not n12352 ; n12352_not
g68290 not n12082 ; n12082_not
g68291 not n23422 ; n23422_not
g68292 not n23143 ; n23143_not
g68293 not n20263 ; n20263_not
g68294 not n24205 ; n24205_not
g68295 not n12343 ; n12343_not
g68296 not n12091 ; n12091_not
g68297 not n23431 ; n23431_not
g68298 not n22207 ; n22207_not
g68299 not n37120 ; n37120_not
g68300 not n42331 ; n42331_not
g68301 not n42403 ; n42403_not
g68302 not n24214 ; n24214_not
g68303 not n27112 ; n27112_not
g68304 not n16141 ; n16141_not
g68305 not n16006 ; n16006_not
g68306 not n13306 ; n13306_not
g68307 not n13432 ; n13432_not
g68308 not n12910 ; n12910_not
g68309 not n34501 ; n34501_not
g68310 not n50251 ; n50251_not
g68311 not n34330 ; n34330_not
g68312 not n12901 ; n12901_not
g68313 not n13441 ; n13441_not
g68314 not n13342 ; n13342_not
g68315 not n16024 ; n16024_not
g68316 not n13072 ; n13072_not
g68317 not n51115 ; n51115_not
g68318 not n20155 ; n20155_not
g68319 not n13414 ; n13414_not
g68320 not n23017 ; n23017_not
g68321 not n20038 ; n20038_not
g68322 not n51133 ; n51133_not
g68323 not n16015 ; n16015_not
g68324 not n34510 ; n34510_not
g68325 not n30532 ; n30532_not
g68326 not n13423 ; n13423_not
g68327 not n12703 ; n12703_not
g68328 not n22801 ; n22801_not
g68329 not n50008 ; n50008_not
g68330 not n12712 ; n12712_not
g68331 not n22027 ; n22027_not
g68332 not n36202 ; n36202_not
g68333 not n16312 ; n16312_not
g68334 not n51034 ; n51034_not
g68335 not n20164 ; n20164_not
g68336 not n16213 ; n16213_not
g68337 not n13081 ; n13081_not
g68338 not n13450 ; n13450_not
g68339 not n30523 ; n30523_not
g68340 not n50017 ; n50017_not
g68341 not n20173 ; n20173_not
g68342 not n34321 ; n34321_not
g68343 not n34006 ; n34006_not
g68344 not n13045 ; n13045_not
g68345 not n45121 ; n45121_not
g68346 not n13036 ; n13036_not
g68347 not n12604 ; n12604_not
g68348 not n16051 ; n16051_not
g68349 not n20137 ; n20137_not
g68350 not n16240 ; n16240_not
g68351 not n27130 ; n27130_not
g68352 not n13027 ; n13027_not
g68353 not n13333 ; n13333_not
g68354 not n16222 ; n16222_not
g68355 not n13063 ; n13063_not
g68356 not n27301 ; n27301_not
g68357 not n20056 ; n20056_not
g68358 not n13054 ; n13054_not
g68359 not n38020 ; n38020_not
g68360 not n13360 ; n13360_not
g68361 not n16231 ; n16231_not
g68362 not n16060 ; n16060_not
g68363 not n16033 ; n16033_not
g68364 not n48100 ; n48100_not
g68365 not n32701 ; n32701_not
g68366 not n47110 ; n47110_not
g68367 not n51124 ; n51124_not
g68368 not n20128 ; n20128_not
g68369 not n50026 ; n50026_not
g68370 not n13405 ; n13405_not
g68371 not n27400 ; n27400_not
g68372 not n16402 ; n16402_not
g68373 not n20047 ; n20047_not
g68374 not n13018 ; n13018_not
g68375 not n16042 ; n16042_not
g68376 not n12613 ; n12613_not
g68377 not n13009 ; n13009_not
g68378 not n12622 ; n12622_not
g68379 not n56020 ; n56020_not
g68380 not n20146 ; n20146_not
g68381 not n50602 ; n50602_not
g68382 not n27310 ; n27310_not
g68383 not n51016 ; n51016_not
g68384 not n52501 ; n52501_not
g68385 not n22081 ; n22081_not
g68386 not n41341 ; n41341_not
g68387 not n41602 ; n41602_not
g68388 not n22090 ; n22090_not
g68389 not n20209 ; n20209_not
g68390 not n30730 ; n30730_not
g68391 not n41332 ; n41332_not
g68392 not n12631 ; n12631_not
g68393 not n23116 ; n23116_not
g68394 not n20812 ; n20812_not
g68395 not n53500 ; n53500_not
g68396 not n22711 ; n22711_not
g68397 not n34042 ; n34042_not
g68398 not n22072 ; n22072_not
g68399 not n32602 ; n32602_not
g68400 not n27220 ; n27220_not
g68401 not n22702 ; n22702_not
g68402 not n34051 ; n34051_not
g68403 not n29200 ; n29200_not
g68404 not n12811 ; n12811_not
g68405 not n55300 ; n55300_not
g68406 not n41323 ; n41323_not
g68407 not n13612 ; n13612_not
g68408 not n34411 ; n34411_not
g68409 not n40801 ; n40801_not
g68410 not n16600 ; n16600_not
g68411 not n27211 ; n27211_not
g68412 not n41611 ; n41611_not
g68413 not n23125 ; n23125_not
g68414 not n13216 ; n13216_not
g68415 not n15043 ; n15043_not
g68416 not n13207 ; n13207_not
g68417 not n41620 ; n41620_not
g68418 not n13603 ; n13603_not
g68419 not n20182 ; n20182_not
g68420 not n22036 ; n22036_not
g68421 not n34303 ; n34303_not
g68422 not n41530 ; n41530_not
g68423 not n22045 ; n22045_not
g68424 not n51052 ; n51052_not
g68425 not n13504 ; n13504_not
g68426 not n23701 ; n23701_not
g68427 not n32620 ; n32620_not
g68428 not n13261 ; n13261_not
g68429 not n23602 ; n23602_not
g68430 not n34312 ; n34312_not
g68431 not n55120 ; n55120_not
g68432 not n12802 ; n12802_not
g68433 not n40810 ; n40810_not
g68434 not n13531 ; n13531_not
g68435 not n13090 ; n13090_not
g68436 not n12721 ; n12721_not
g68437 not n20803 ; n20803_not
g68438 not n20065 ; n20065_not
g68439 not n13243 ; n13243_not
g68440 not n13540 ; n13540_not
g68441 not n45130 ; n45130_not
g68442 not n22720 ; n22720_not
g68443 not n13513 ; n13513_not
g68444 not n20191 ; n20191_not
g68445 not n12181 ; n12181_not
g68446 not n40720 ; n40720_not
g68447 not n31270 ; n31270_not
g68448 not n13252 ; n13252_not
g68449 not n13522 ; n13522_not
g68450 not n34033 ; n34033_not
g68451 not n16510 ; n16510_not
g68452 not n17041 ; n17041_not
g68453 not n11560 ; n11560_not
g68454 not n32350 ; n32350_not
g68455 not n30073 ; n30073_not
g68456 not n24511 ; n24511_not
g68457 not n11542 ; n11542_not
g68458 not n20092 ; n20092_not
g68459 not n11533 ; n11533_not
g68460 not n11605 ; n11605_not
g68461 not n22009 ; n22009_not
g68462 not n33322 ; n33322_not
g68463 not n20380 ; n20380_not
g68464 not n31171 ; n31171_not
g68465 not n24520 ; n24520_not
g68466 not n57100 ; n57100_not
g68467 not n13270 ; n13270_not
g68468 not n36112 ; n36112_not
g68469 not n13810 ; n13810_not
g68470 not n45220 ; n45220_not
g68471 not n11470 ; n11470_not
g68472 not n21910 ; n21910_not
g68473 not n38011 ; n38011_not
g68474 not n35113 ; n35113_not
g68475 not n21901 ; n21901_not
g68476 not n13225 ; n13225_not
g68477 not n53221 ; n53221_not
g68478 not n55102 ; n55102_not
g68479 not n15601 ; n15601_not
g68480 not n11515 ; n11515_not
g68481 not n54013 ; n54013_not
g68482 not n20920 ; n20920_not
g68483 not n16330 ; n16330_not
g68484 not n43204 ; n43204_not
g68485 not n35104 ; n35104_not
g68486 not n36400 ; n36400_not
g68487 not n32332 ; n32332_not
g68488 not n53230 ; n53230_not
g68489 not n54130 ; n54130_not
g68490 not n50242 ; n50242_not
g68491 not n50503 ; n50503_not
g68492 not n31702 ; n31702_not
g68493 not n35050 ; n35050_not
g68494 not n50170 ; n50170_not
g68495 not n31144 ; n31144_not
g68496 not n11704 ; n11704_not
g68497 not n27022 ; n27022_not
g68498 not n35041 ; n35041_not
g68499 not n20902 ; n20902_not
g68500 not n54004 ; n54004_not
g68501 not n47002 ; n47002_not
g68502 not n20362 ; n20362_not
g68503 not n19120 ; n19120_not
g68504 not n11641 ; n11641_not
g68505 not n20371 ; n20371_not
g68506 not n11632 ; n11632_not
g68507 not n11623 ; n11623_not
g68508 not n22018 ; n22018_not
g68509 not n20911 ; n20911_not
g68510 not n11092 ; n11092_not
g68511 not n22054 ; n22054_not
g68512 not n11425 ; n11425_not
g68513 not n50620 ; n50620_not
g68514 not n11650 ; n11650_not
g68515 not n25222 ; n25222_not
g68516 not n21811 ; n21811_not
g68517 not n11254 ; n11254_not
g68518 not n11245 ; n11245_not
g68519 not n21802 ; n21802_not
g68520 not n14341 ; n14341_not
g68521 not n11272 ; n11272_not
g68522 not n20407 ; n20407_not
g68523 not n31252 ; n31252_not
g68524 not n21820 ; n21820_not
g68525 not n32260 ; n32260_not
g68526 not n11263 ; n11263_not
g68527 not n33700 ; n33700_not
g68528 not n23071 ; n23071_not
g68529 not n30145 ; n30145_not
g68530 not n32242 ; n32242_not
g68531 not n14404 ; n14404_not
g68532 not n11182 ; n11182_not
g68533 not n25303 ; n25303_not
g68534 not n11236 ; n11236_not
g68535 not n11227 ; n11227_not
g68536 not n41422 ; n41422_not
g68537 not n32251 ; n32251_not
g68538 not n11218 ; n11218_not
g68539 not n11209 ; n11209_not
g68540 not n31234 ; n31234_not
g68541 not n20416 ; n20416_not
g68542 not n42304 ; n42304_not
g68543 not n11191 ; n11191_not
g68544 not n11407 ; n11407_not
g68545 not n50215 ; n50215_not
g68546 not n21343 ; n21343_not
g68547 not n35131 ; n35131_not
g68548 not n45301 ; n45301_not
g68549 not n11380 ; n11380_not
g68550 not n11371 ; n11371_not
g68551 not n17131 ; n17131_not
g68552 not n11452 ; n11452_not
g68553 not n11443 ; n11443_not
g68554 not n31216 ; n31216_not
g68555 not n11416 ; n11416_not
g68556 not n35122 ; n35122_not
g68557 not n11317 ; n11317_not
g68558 not n30118 ; n30118_not
g68559 not n11308 ; n11308_not
g68560 not n24430 ; n24430_not
g68561 not n31243 ; n31243_not
g68562 not n11290 ; n11290_not
g68563 not n24421 ; n24421_not
g68564 not n20704 ; n20704_not
g68565 not n11281 ; n11281_not
g68566 not n50233 ; n50233_not
g68567 not n35140 ; n35140_not
g68568 not n50035 ; n50035_not
g68569 not n11362 ; n11362_not
g68570 not n10903 ; n10903_not
g68571 not n11353 ; n11353_not
g68572 not n11344 ; n11344_not
g68573 not n11335 ; n11335_not
g68574 not n50431 ; n50431_not
g68575 not n31009 ; n31009_not
g68576 not n11326 ; n11326_not
g68577 not n36040 ; n36040_not
g68578 not n22234 ; n22234_not
g68579 not n20119 ; n20119_not
g68580 not n24601 ; n24601_not
g68581 not n24610 ; n24610_not
g68582 not n50143 ; n50143_not
g68583 not n19300 ; n19300_not
g68584 not n20083 ; n20083_not
g68585 not n12055 ; n12055_not
g68586 not n22261 ; n22261_not
g68587 not n50440 ; n50440_not
g68588 not n20317 ; n20317_not
g68589 not n31045 ; n31045_not
g68590 not n31063 ; n31063_not
g68591 not n11920 ; n11920_not
g68592 not n36031 ; n36031_not
g68593 not n27031 ; n27031_not
g68594 not n20722 ; n20722_not
g68595 not n24700 ; n24700_not
g68596 not n11911 ; n11911_not
g68597 not n31072 ; n31072_not
g68598 not n50800 ; n50800_not
g68599 not n41800 ; n41800_not
g68600 not n31054 ; n31054_not
g68601 not n40108 ; n40108_not
g68602 not n20326 ; n20326_not
g68603 not n34015 ; n34015_not
g68604 not n13180 ; n13180_not
g68605 not n28120 ; n28120_not
g68606 not n38200 ; n38200_not
g68607 not n50080 ; n50080_not
g68608 not n22351 ; n22351_not
g68609 not n12190 ; n12190_not
g68610 not n12172 ; n12172_not
g68611 not n31018 ; n31018_not
g68612 not n22342 ; n22342_not
g68613 not n36022 ; n36022_not
g68614 not n22333 ; n22333_not
g68615 not n12217 ; n12217_not
g68616 not n24340 ; n24340_not
g68617 not n36013 ; n36013_not
g68618 not n12208 ; n12208_not
g68619 not n16114 ; n16114_not
g68620 not n22360 ; n22360_not
g68621 not n22270 ; n22270_not
g68622 not n12163 ; n12163_not
g68623 not n34105 ; n34105_not
g68624 not n20713 ; n20713_not
g68625 not n47020 ; n47020_not
g68626 not n31036 ; n31036_not
g68627 not n20308 ; n20308_not
g68628 not n51007 ; n51007_not
g68629 not n13351 ; n13351_not
g68630 not n34060 ; n34060_not
g68631 not n24403 ; n24403_not
g68632 not n22324 ; n22324_not
g68633 not n24412 ; n24412_not
g68634 not n12145 ; n12145_not
g68635 not n22315 ; n22315_not
g68636 not n31027 ; n31027_not
g68637 not n31711 ; n31711_not
g68638 not n30541 ; n30541_not
g68639 not n41431 ; n41431_not
g68640 not n35023 ; n35023_not
g68641 not n31135 ; n31135_not
g68642 not n49000 ; n49000_not
g68643 not n11803 ; n11803_not
g68644 not n20344 ; n20344_not
g68645 not n22144 ; n22144_not
g68646 not n51061 ; n51061_not
g68647 not n31126 ; n31126_not
g68648 not n35014 ; n35014_not
g68649 not n32422 ; n32422_not
g68650 not n40153 ; n40153_not
g68651 not n32404 ; n32404_not
g68652 not n11722 ; n11722_not
g68653 not n11713 ; n11713_not
g68654 not n32413 ; n32413_not
g68655 not n11740 ; n11740_not
g68656 not n11551 ; n11551_not
g68657 not n35032 ; n35032_not
g68658 not n20353 ; n20353_not
g68659 not n11731 ; n11731_not
g68660 not n23026 ; n23026_not
g68661 not n50071 ; n50071_not
g68662 not n37003 ; n37003_not
g68663 not n27004 ; n27004_not
g68664 not n50125 ; n50125_not
g68665 not n19210 ; n19210_not
g68666 not n13900 ; n13900_not
g68667 not n11902 ; n11902_not
g68668 not n11461 ; n11461_not
g68669 not n32440 ; n32440_not
g68670 not n31081 ; n31081_not
g68671 not n47011 ; n47011_not
g68672 not n27040 ; n27040_not
g68673 not n31090 ; n31090_not
g68674 not n11830 ; n11830_not
g68675 not n11821 ; n11821_not
g68676 not n11506 ; n11506_not
g68677 not n31117 ; n31117_not
g68678 not n11812 ; n11812_not
g68679 not n35005 ; n35005_not
g68680 not n54103 ; n54103_not
g68681 not n20335 ; n20335_not
g68682 not n32431 ; n32431_not
g68683 not n46300 ; n46300_not
g68684 not n16303 ; n16303_not
g68685 not n31108 ; n31108_not
g68686 not n33044 ; n33044_not
g68687 not n31802 ; n31802_not
g68688 not n17231 ; n17231_not
g68689 not n17240 ; n17240_not
g68690 not n45212 ; n45212_not
g68691 not n31811 ; n31811_not
g68692 not n31703 ; n31703_not
g68693 not n15620 ; n15620_not
g68694 not n54131 ; n54131_not
g68695 not n17501 ; n17501_not
g68696 not n17510 ; n17510_not
g68697 not n30308 ; n30308_not
g68698 not n17330 ; n17330_not
g68699 not n17321 ; n17321_not
g68700 not n31721 ; n31721_not
g68701 not n45221 ; n45221_not
g68702 not n17312 ; n17312_not
g68703 not n17420 ; n17420_not
g68704 not n31451 ; n31451_not
g68705 not n31712 ; n31712_not
g68706 not n17303 ; n17303_not
g68707 not n30191 ; n30191_not
g68708 not n31406 ; n31406_not
g68709 not n31415 ; n31415_not
g68710 not n45302 ; n45302_not
g68711 not n31424 ; n31424_not
g68712 not n30380 ; n30380_not
g68713 not n17411 ; n17411_not
g68714 not n20705 ; n20705_not
g68715 not n17402 ; n17402_not
g68716 not n47201 ; n47201_not
g68717 not n42503 ; n42503_not
g68718 not n50621 ; n50621_not
g68719 not n42800 ; n42800_not
g68720 not n20714 ; n20714_not
g68721 not n50162 ; n50162_not
g68722 not n30182 ; n30182_not
g68723 not n17222 ; n17222_not
g68724 not n45230 ; n45230_not
g68725 not n42521 ; n42521_not
g68726 not n17213 ; n17213_not
g68727 not n42422 ; n42422_not
g68728 not n17204 ; n17204_not
g68729 not n43421 ; n43421_not
g68730 not n54140 ; n54140_not
g68731 not n15008 ; n15008_not
g68732 not n31361 ; n31361_not
g68733 not n37400 ; n37400_not
g68734 not n31514 ; n31514_not
g68735 not n42413 ; n42413_not
g68736 not n42530 ; n42530_not
g68737 not n50603 ; n50603_not
g68738 not n32810 ; n32810_not
g68739 not n43403 ; n43403_not
g68740 not n54230 ; n54230_not
g68741 not n55130 ; n55130_not
g68742 not n20732 ; n20732_not
g68743 not n42440 ; n42440_not
g68744 not n50612 ; n50612_not
g68745 not n42431 ; n42431_not
g68746 not n54221 ; n54221_not
g68747 not n17600 ; n17600_not
g68748 not n20660 ; n20660_not
g68749 not n43205 ; n43205_not
g68750 not n43412 ; n43412_not
g68751 not n31370 ; n31370_not
g68752 not n50171 ; n50171_not
g68753 not n30173 ; n30173_not
g68754 not n20750 ; n20750_not
g68755 not n16061 ; n16061_not
g68756 not n30821 ; n30821_not
g68757 not n19202 ; n19202_not
g68758 not n50126 ; n50126_not
g68759 not n30812 ; n30812_not
g68760 not n19211 ; n19211_not
g68761 not n32504 ; n32504_not
g68762 not n16070 ; n16070_not
g68763 not n30803 ; n30803_not
g68764 not n16124 ; n16124_not
g68765 not n20282 ; n20282_not
g68766 not n41261 ; n41261_not
g68767 not n41252 ; n41252_not
g68768 not n43151 ; n43151_not
g68769 not n32801 ; n32801_not
g68770 not n32324 ; n32324_not
g68771 not n15701 ; n15701_not
g68772 not n20291 ; n20291_not
g68773 not n16115 ; n16115_not
g68774 not n16106 ; n16106_not
g68775 not n53204 ; n53204_not
g68776 not n32333 ; n32333_not
g68777 not n15710 ; n15710_not
g68778 not n55202 ; n55202_not
g68779 not n41243 ; n41243_not
g68780 not n31019 ; n31019_not
g68781 not n53213 ; n53213_not
g68782 not n50441 ; n50441_not
g68783 not n50450 ; n50450_not
g68784 not n30902 ; n30902_not
g68785 not n16151 ; n16151_not
g68786 not n20255 ; n20255_not
g68787 not n54401 ; n54401_not
g68788 not n16025 ; n16025_not
g68789 not n30911 ; n30911_not
g68790 not n53123 ; n53123_not
g68791 not n55220 ; n55220_not
g68792 not n50261 ; n50261_not
g68793 not n16700 ; n16700_not
g68794 not n16034 ; n16034_not
g68795 not n50702 ; n50702_not
g68796 not n16142 ; n16142_not
g68797 not n53132 ; n53132_not
g68798 not n20264 ; n20264_not
g68799 not n32513 ; n32513_not
g68800 not n16043 ; n16043_not
g68801 not n54410 ; n54410_not
g68802 not n50117 ; n50117_not
g68803 not n16403 ; n16403_not
g68804 not n47300 ; n47300_not
g68805 not n43142 ; n43142_not
g68806 not n16052 ; n16052_not
g68807 not n16133 ; n16133_not
g68808 not n53141 ; n53141_not
g68809 not n55310 ; n55310_not
g68810 not n32315 ; n32315_not
g68811 not n53150 ; n53150_not
g68812 not n20273 ; n20273_not
g68813 not n30830 ; n30830_not
g68814 not n19220 ; n19220_not
g68815 not n16214 ; n16214_not
g68816 not n30470 ; n30470_not
g68817 not n16304 ; n16304_not
g68818 not n32432 ; n32432_not
g68819 not n54500 ; n54500_not
g68820 not n16223 ; n16223_not
g68821 not n20336 ; n20336_not
g68822 not n32360 ; n32360_not
g68823 not n16232 ; n16232_not
g68824 not n31109 ; n31109_not
g68825 not n38021 ; n38021_not
g68826 not n16241 ; n16241_not
g68827 not n31118 ; n31118_not
g68828 not n16250 ; n16250_not
g68829 not n20345 ; n20345_not
g68830 not n32423 ; n32423_not
g68831 not n31127 ; n31127_not
g68832 not n54113 ; n54113_not
g68833 not n32414 ; n32414_not
g68834 not n31136 ; n31136_not
g68835 not n20354 ; n20354_not
g68836 not n32405 ; n32405_not
g68837 not n19130 ; n19130_not
g68838 not n53510 ; n53510_not
g68839 not n31145 ; n31145_not
g68840 not n31028 ; n31028_not
g68841 not n20309 ; n20309_not
g68842 not n31037 ; n31037_not
g68843 not n53222 ; n53222_not
g68844 not n41423 ; n41423_not
g68845 not n31046 ; n31046_not
g68846 not n20318 ; n20318_not
g68847 not n53240 ; n53240_not
g68848 not n16340 ; n16340_not
g68849 not n16160 ; n16160_not
g68850 not n53231 ; n53231_not
g68851 not n31055 ; n31055_not
g68852 not n41810 ; n41810_not
g68853 not n32450 ; n32450_not
g68854 not n31064 ; n31064_not
g68855 not n20327 ; n20327_not
g68856 not n31073 ; n31073_not
g68857 not n32441 ; n32441_not
g68858 not n31082 ; n31082_not
g68859 not n16205 ; n16205_not
g68860 not n38030 ; n38030_not
g68861 not n31091 ; n31091_not
g68862 not n16313 ; n16313_not
g68863 not n32630 ; n32630_not
g68864 not n43016 ; n43016_not
g68865 not n16430 ; n16430_not
g68866 not n20165 ; n20165_not
g68867 not n43007 ; n43007_not
g68868 not n20174 ; n20174_not
g68869 not n19301 ; n19301_not
g68870 not n30533 ; n30533_not
g68871 not n38111 ; n38111_not
g68872 not n32702 ; n32702_not
g68873 not n20183 ; n20183_not
g68874 not n30605 ; n30605_not
g68875 not n30614 ; n30614_not
g68876 not n30506 ; n30506_not
g68877 not n30623 ; n30623_not
g68878 not n16502 ; n16502_not
g68879 not n20192 ; n20192_not
g68880 not n30515 ; n30515_not
g68881 not n16511 ; n16511_not
g68882 not n30632 ; n30632_not
g68883 not n45131 ; n45131_not
g68884 not n43061 ; n43061_not
g68885 not n30542 ; n30542_not
g68886 not n20093 ; n20093_not
g68887 not n20084 ; n20084_not
g68888 not n50243 ; n50243_not
g68889 not n16322 ; n16322_not
g68890 not n43043 ; n43043_not
g68891 not n20075 ; n20075_not
g68892 not n53501 ; n53501_not
g68893 not n20066 ; n20066_not
g68894 not n43052 ; n43052_not
g68895 not n20129 ; n20129_not
g68896 not n30560 ; n30560_not
g68897 not n20057 ; n20057_not
g68898 not n20048 ; n20048_not
g68899 not n20138 ; n20138_not
g68900 not n43034 ; n43034_not
g68901 not n20147 ; n20147_not
g68902 not n16412 ; n16412_not
g68903 not n43025 ; n43025_not
g68904 not n20039 ; n20039_not
g68905 not n20156 ; n20156_not
g68906 not n45401 ; n45401_not
g68907 not n53060 ; n53060_not
g68908 not n20228 ; n20228_not
g68909 not n19103 ; n19103_not
g68910 not n30731 ; n30731_not
g68911 not n50108 ; n50108_not
g68912 not n30722 ; n30722_not
g68913 not n41306 ; n41306_not
g68914 not n19112 ; n19112_not
g68915 not n43124 ; n43124_not
g68916 not n19121 ; n19121_not
g68917 not n32540 ; n32540_not
g68918 not n30713 ; n30713_not
g68919 not n20237 ; n20237_not
g68920 not n32531 ; n32531_not
g68921 not n53330 ; n53330_not
g68922 not n50252 ; n50252_not
g68923 not n38120 ; n38120_not
g68924 not n50711 ; n50711_not
g68925 not n20246 ; n20246_not
g68926 not n53105 ; n53105_not
g68927 not n16007 ; n16007_not
g68928 not n32522 ; n32522_not
g68929 not n53321 ; n53321_not
g68930 not n53114 ; n53114_not
g68931 not n16016 ; n16016_not
g68932 not n30641 ; n30641_not
g68933 not n30650 ; n30650_not
g68934 not n32612 ; n32612_not
g68935 not n53420 ; n53420_not
g68936 not n41351 ; n41351_not
g68937 not n45410 ; n45410_not
g68938 not n45122 ; n45122_not
g68939 not n41342 ; n41342_not
g68940 not n53411 ; n53411_not
g68941 not n41333 ; n41333_not
g68942 not n30740 ; n30740_not
g68943 not n43106 ; n43106_not
g68944 not n53006 ; n53006_not
g68945 not n19040 ; n19040_not
g68946 not n53015 ; n53015_not
g68947 not n16601 ; n16601_not
g68948 not n53024 ; n53024_not
g68949 not n16610 ; n16610_not
g68950 not n20219 ; n20219_not
g68951 not n50720 ; n50720_not
g68952 not n53033 ; n53033_not
g68953 not n55301 ; n55301_not
g68954 not n53042 ; n53042_not
g68955 not n53051 ; n53051_not
g68956 not n31163 ; n31163_not
g68957 not n32045 ; n32045_not
g68958 not n32144 ; n32144_not
g68959 not n32054 ; n32054_not
g68960 not n55004 ; n55004_not
g68961 not n50216 ; n50216_not
g68962 not n30218 ; n30218_not
g68963 not n32135 ; n32135_not
g68964 not n33026 ; n33026_not
g68965 not n31433 ; n31433_not
g68966 not n32126 ; n32126_not
g68967 not n43250 ; n43250_not
g68968 not n43331 ; n43331_not
g68969 not n50531 ; n50531_not
g68970 not n32117 ; n32117_not
g68971 not n31460 ; n31460_not
g68972 not n20552 ; n20552_not
g68973 not n32108 ; n32108_not
g68974 not n54320 ; n54320_not
g68975 not n17042 ; n17042_not
g68976 not n17033 ; n17033_not
g68977 not n30416 ; n30416_not
g68978 not n32081 ; n32081_not
g68979 not n45320 ; n45320_not
g68980 not n37202 ; n37202_not
g68981 not n50405 ; n50405_not
g68982 not n17114 ; n17114_not
g68983 not n37211 ; n37211_not
g68984 not n32180 ; n32180_not
g68985 not n42701 ; n42701_not
g68986 not n20507 ; n20507_not
g68987 not n30425 ; n30425_not
g68988 not n43304 ; n43304_not
g68989 not n18500 ; n18500_not
g68990 not n32171 ; n32171_not
g68991 not n32036 ; n32036_not
g68992 not n42710 ; n42710_not
g68993 not n42008 ; n42008_not
g68994 not n43313 ; n43313_not
g68995 not n37220 ; n37220_not
g68996 not n55022 ; n55022_not
g68997 not n32162 ; n32162_not
g68998 not n42620 ; n42620_not
g68999 not n31172 ; n31172_not
g69000 not n50522 ; n50522_not
g69001 not n20525 ; n20525_not
g69002 not n43322 ; n43322_not
g69003 not n33008 ; n33008_not
g69004 not n50153 ; n50153_not
g69005 not n32153 ; n32153_not
g69006 not n20534 ; n20534_not
g69007 not n20615 ; n20615_not
g69008 not n32063 ; n32063_not
g69009 not n18410 ; n18410_not
g69010 not n50207 ; n50207_not
g69011 not n50630 ; n50630_not
g69012 not n20624 ; n20624_not
g69013 not n31307 ; n31307_not
g69014 not n54104 ; n54104_not
g69015 not n37310 ; n37310_not
g69016 not n31316 ; n31316_not
g69017 not n31325 ; n31325_not
g69018 not n45311 ; n45311_not
g69019 not n50540 ; n50540_not
g69020 not n31334 ; n31334_not
g69021 not n20642 ; n20642_not
g69022 not n31343 ; n31343_not
g69023 not n18320 ; n18320_not
g69024 not n31352 ; n31352_not
g69025 not n32018 ; n32018_not
g69026 not n17024 ; n17024_not
g69027 not n43241 ; n43241_not
g69028 not n54311 ; n54311_not
g69029 not n32090 ; n32090_not
g69030 not n20570 ; n20570_not
g69031 not n43340 ; n43340_not
g69032 not n30209 ; n30209_not
g69033 not n42611 ; n42611_not
g69034 not n33053 ; n33053_not
g69035 not n30407 ; n30407_not
g69036 not n30290 ; n30290_not
g69037 not n55400 ; n55400_not
g69038 not n31505 ; n31505_not
g69039 not n31262 ; n31262_not
g69040 not n31271 ; n31271_not
g69041 not n33017 ; n33017_not
g69042 not n43232 ; n43232_not
g69043 not n31280 ; n31280_not
g69044 not n37301 ; n37301_not
g69045 not n19022 ; n19022_not
g69046 not n32342 ; n32342_not
g69047 not n19013 ; n19013_not
g69048 not n41900 ; n41900_not
g69049 not n19004 ; n19004_not
g69050 not n20390 ; n20390_not
g69051 not n50432 ; n50432_not
g69052 not n41432 ; n41432_not
g69053 not n31208 ; n31208_not
g69054 not n54203 ; n54203_not
g69055 not n30452 ; n30452_not
g69056 not n17123 ; n17123_not
g69057 not n31226 ; n31226_not
g69058 not n43214 ; n43214_not
g69059 not n17141 ; n17141_not
g69060 not n31244 ; n31244_not
g69061 not n31253 ; n31253_not
g69062 not n50504 ; n50504_not
g69063 not n30263 ; n30263_not
g69064 not n20363 ; n20363_not
g69065 not n30461 ; n30461_not
g69066 not n31154 ; n31154_not
g69067 not n17006 ; n17006_not
g69068 not n20372 ; n20372_not
g69069 not n55112 ; n55112_not
g69070 not n19031 ; n19031_not
g69071 not n20381 ; n20381_not
g69072 not n31181 ; n31181_not
g69073 not n17051 ; n17051_not
g69074 not n30443 ; n30443_not
g69075 not n32009 ; n32009_not
g69076 not n20453 ; n20453_not
g69077 not n30254 ; n30254_not
g69078 not n32216 ; n32216_not
g69079 not n20462 ; n20462_not
g69080 not n32207 ; n32207_not
g69081 not n47102 ; n47102_not
g69082 not n41405 ; n41405_not
g69083 not n20471 ; n20471_not
g69084 not n50414 ; n50414_not
g69085 not n30236 ; n30236_not
g69086 not n42017 ; n42017_not
g69087 not n20480 ; n20480_not
g69088 not n55040 ; n55040_not
g69089 not n42026 ; n42026_not
g69090 not n30434 ; n30434_not
g69091 not n17132 ; n17132_not
g69092 not n30227 ; n30227_not
g69093 not n38003 ; n38003_not
g69094 not n20408 ; n20408_not
g69095 not n32603 ; n32603_not
g69096 not n32261 ; n32261_not
g69097 not n32252 ; n32252_not
g69098 not n20417 ; n20417_not
g69099 not n32243 ; n32243_not
g69100 not n47111 ; n47111_not
g69101 not n50423 ; n50423_not
g69102 not n20426 ; n20426_not
g69103 not n32900 ; n32900_not
g69104 not n50513 ; n50513_not
g69105 not n30245 ; n30245_not
g69106 not n32234 ; n32234_not
g69107 not n20435 ; n20435_not
g69108 not n45104 ; n45104_not
g69109 not n15800 ; n15800_not
g69110 not n31217 ; n31217_not
g69111 not n32225 ; n32225_not
g69112 not n20444 ; n20444_not
g69113 not n10049 ; n10049_not
g69114 not n23126 ; n23126_not
g69115 not n10058 ; n10058_not
g69116 not n12623 ; n12623_not
g69117 not n23117 ; n23117_not
g69118 not n23135 ; n23135_not
g69119 not n12641 ; n12641_not
g69120 not n23144 ; n23144_not
g69121 not n10067 ; n10067_not
g69122 not n34421 ; n34421_not
g69123 not n23153 ; n23153_not
g69124 not n23162 ; n23162_not
g69125 not n23171 ; n23171_not
g69126 not n29201 ; n29201_not
g69127 not n23180 ; n23180_not
g69128 not n10076 ; n10076_not
g69129 not n23207 ; n23207_not
g69130 not n23216 ; n23216_not
g69131 not n25304 ; n25304_not
g69132 not n40802 ; n40802_not
g69133 not n10571 ; n10571_not
g69134 not n40145 ; n40145_not
g69135 not n40811 ; n40811_not
g69136 not n28103 ; n28103_not
g69137 not n10562 ; n10562_not
g69138 not n10553 ; n10553_not
g69139 not n40127 ; n40127_not
g69140 not n10544 ; n10544_not
g69141 not n10535 ; n10535_not
g69142 not n10517 ; n10517_not
g69143 not n29120 ; n29120_not
g69144 not n10526 ; n10526_not
g69145 not n12614 ; n12614_not
g69146 not n23900 ; n23900_not
g69147 not n10472 ; n10472_not
g69148 not n23324 ; n23324_not
g69149 not n23333 ; n23333_not
g69150 not n23342 ; n23342_not
g69151 not n23351 ; n23351_not
g69152 not n12731 ; n12731_not
g69153 not n51044 ; n51044_not
g69154 not n23360 ; n23360_not
g69155 not n10139 ; n10139_not
g69156 not n10454 ; n10454_not
g69157 not n40307 ; n40307_not
g69158 not n10148 ; n10148_not
g69159 not n23405 ; n23405_not
g69160 not n23414 ; n23414_not
g69161 not n40820 ; n40820_not
g69162 not n10157 ; n10157_not
g69163 not n23423 ; n23423_not
g69164 not n23432 ; n23432_not
g69165 not n23711 ; n23711_not
g69166 not n23441 ; n23441_not
g69167 not n23225 ; n23225_not
g69168 not n52403 ; n52403_not
g69169 not n37130 ; n37130_not
g69170 not n23234 ; n23234_not
g69171 not n23243 ; n23243_not
g69172 not n10085 ; n10085_not
g69173 not n23252 ; n23252_not
g69174 not n23261 ; n23261_not
g69175 not n40019 ; n40019_not
g69176 not n23270 ; n23270_not
g69177 not n23801 ; n23801_not
g69178 not n34430 ; n34430_not
g69179 not n10481 ; n10481_not
g69180 not n10094 ; n10094_not
g69181 not n23306 ; n23306_not
g69182 not n12704 ; n12704_not
g69183 not n52412 ; n52412_not
g69184 not n23315 ; n23315_not
g69185 not n12713 ; n12713_not
g69186 not n40712 ; n40712_not
g69187 not n10427 ; n10427_not
g69188 not n29030 ; n29030_not
g69189 not n10193 ; n10193_not
g69190 not n24152 ; n24152_not
g69191 not n10184 ; n10184_not
g69192 not n10436 ; n10436_not
g69193 not n24143 ; n24143_not
g69194 not n40721 ; n40721_not
g69195 not n24134 ; n24134_not
g69196 not n10175 ; n10175_not
g69197 not n56003 ; n56003_not
g69198 not n12056 ; n12056_not
g69199 not n24125 ; n24125_not
g69200 not n12047 ; n12047_not
g69201 not n56102 ; n56102_not
g69202 not n10670 ; n10670_not
g69203 not n10445 ; n10445_not
g69204 not n24116 ; n24116_not
g69205 not n12038 ; n12038_not
g69206 not n10166 ; n10166_not
g69207 not n24107 ; n24107_not
g69208 not n52601 ; n52601_not
g69209 not n40190 ; n40190_not
g69210 not n56111 ; n56111_not
g69211 not n40244 ; n40244_not
g69212 not n12092 ; n12092_not
g69213 not n24215 ; n24215_not
g69214 not n52241 ; n52241_not
g69215 not n10742 ; n10742_not
g69216 not n10238 ; n10238_not
g69217 not n24206 ; n24206_not
g69218 not n12083 ; n12083_not
g69219 not n40235 ; n40235_not
g69220 not n52250 ; n52250_not
g69221 not n10733 ; n10733_not
g69222 not n10229 ; n10229_not
g69223 not n10724 ; n10724_not
g69224 not n37121 ; n37121_not
g69225 not n52520 ; n52520_not
g69226 not n45032 ; n45032_not
g69227 not n10715 ; n10715_not
g69228 not n24170 ; n24170_not
g69229 not n40217 ; n40217_not
g69230 not n10706 ; n10706_not
g69231 not n24161 ; n24161_not
g69232 not n35303 ; n35303_not
g69233 not n52331 ; n52331_not
g69234 not n24026 ; n24026_not
g69235 not n10616 ; n10616_not
g69236 not n52340 ; n52340_not
g69237 not n24017 ; n24017_not
g69238 not n10607 ; n10607_not
g69239 not n47030 ; n47030_not
g69240 not n35411 ; n35411_not
g69241 not n24008 ; n24008_not
g69242 not n12533 ; n12533_not
g69243 not n34700 ; n34700_not
g69244 not n12551 ; n12551_not
g69245 not n10490 ; n10490_not
g69246 not n35420 ; n35420_not
g69247 not n40154 ; n40154_not
g69248 not n10580 ; n10580_not
g69249 not n52502 ; n52502_not
g69250 not n28301 ; n28301_not
g69251 not n10661 ; n10661_not
g69252 not n35402 ; n35402_not
g69253 not n45005 ; n45005_not
g69254 not n10652 ; n10652_not
g69255 not n24080 ; n24080_not
g69256 not n52304 ; n52304_not
g69257 not n24071 ; n24071_not
g69258 not n25340 ; n25340_not
g69259 not n10643 ; n10643_not
g69260 not n24062 ; n24062_not
g69261 not n52313 ; n52313_not
g69262 not n10634 ; n10634_not
g69263 not n24053 ; n24053_not
g69264 not n52322 ; n52322_not
g69265 not n25331 ; n25331_not
g69266 not n10625 ; n10625_not
g69267 not n24044 ; n24044_not
g69268 not n56300 ; n56300_not
g69269 not n40172 ; n40172_not
g69270 not n24035 ; n24035_not
g69271 not n34403 ; n34403_not
g69272 not n13235 ; n13235_not
g69273 not n22307 ; n22307_not
g69274 not n28211 ; n28211_not
g69275 not n51053 ; n51053_not
g69276 not n23063 ; n23063_not
g69277 not n13253 ; n13253_not
g69278 not n23054 ; n23054_not
g69279 not n13262 ; n13262_not
g69280 not n47021 ; n47021_not
g69281 not n52430 ; n52430_not
g69282 not n24413 ; n24413_not
g69283 not n26114 ; n26114_not
g69284 not n23036 ; n23036_not
g69285 not n41009 ; n41009_not
g69286 not n39002 ; n39002_not
g69287 not n40064 ; n40064_not
g69288 not n13280 ; n13280_not
g69289 not n23018 ; n23018_not
g69290 not n23009 ; n23009_not
g69291 not n35501 ; n35501_not
g69292 not n13307 ; n13307_not
g69293 not n26132 ; n26132_not
g69294 not n40082 ; n40082_not
g69295 not n40433 ; n40433_not
g69296 not n13325 ; n13325_not
g69297 not n26141 ; n26141_not
g69298 not n25223 ; n25223_not
g69299 not n40046 ; n40046_not
g69300 not n26051 ; n26051_not
g69301 not n13109 ; n13109_not
g69302 not n13118 ; n13118_not
g69303 not n40424 ; n40424_not
g69304 not n13127 ; n13127_not
g69305 not n51071 ; n51071_not
g69306 not n13145 ; n13145_not
g69307 not n28220 ; n28220_not
g69308 not n13136 ; n13136_not
g69309 not n26060 ; n26060_not
g69310 not n13163 ; n13163_not
g69311 not n13172 ; n13172_not
g69312 not n23072 ; n23072_not
g69313 not n40055 ; n40055_not
g69314 not n23108 ; n23108_not
g69315 not n13190 ; n13190_not
g69316 not n23090 ; n23090_not
g69317 not n13208 ; n13208_not
g69318 not n13217 ; n13217_not
g69319 not n12830 ; n12830_not
g69320 not n13406 ; n13406_not
g69321 not n26204 ; n26204_not
g69322 not n34007 ; n34007_not
g69323 not n35222 ; n35222_not
g69324 not n51008 ; n51008_not
g69325 not n13316 ; n13316_not
g69326 not n13415 ; n13415_not
g69327 not n41036 ; n41036_not
g69328 not n44411 ; n44411_not
g69329 not n40460 ; n40460_not
g69330 not n13424 ; n13424_not
g69331 not n13433 ; n13433_not
g69332 not n26222 ; n26222_not
g69333 not n34331 ; n34331_not
g69334 not n40037 ; n40037_not
g69335 not n26231 ; n26231_not
g69336 not n34016 ; n34016_not
g69337 not n13442 ; n13442_not
g69338 not n41045 ; n41045_not
g69339 not n35213 ; n35213_not
g69340 not n13451 ; n13451_not
g69341 not n47003 ; n47003_not
g69342 not n40730 ; n40730_not
g69343 not n41054 ; n41054_not
g69344 not n28202 ; n28202_not
g69345 not n41018 ; n41018_not
g69346 not n50045 ; n50045_not
g69347 not n13343 ; n13343_not
g69348 not n13352 ; n13352_not
g69349 not n35510 ; n35510_not
g69350 not n40442 ; n40442_not
g69351 not n13361 ; n13361_not
g69352 not n47012 ; n47012_not
g69353 not n40073 ; n40073_not
g69354 not n13370 ; n13370_not
g69355 not n52421 ; n52421_not
g69356 not n12803 ; n12803_not
g69357 not n51026 ; n51026_not
g69358 not n41027 ; n41027_not
g69359 not n51710 ; n51710_not
g69360 not n12812 ; n12812_not
g69361 not n22901 ; n22901_not
g69362 not n35231 ; n35231_not
g69363 not n40451 ; n40451_not
g69364 not n34340 ; n34340_not
g69365 not n12821 ; n12821_not
g69366 not n26006 ; n26006_not
g69367 not n40334 ; n40334_not
g69368 not n40109 ; n40109_not
g69369 not n34601 ; n34601_not
g69370 not n10409 ; n10409_not
g69371 not n23621 ; n23621_not
g69372 not n23612 ; n23612_not
g69373 not n12722 ; n12722_not
g69374 not n10247 ; n10247_not
g69375 not n23603 ; n23603_not
g69376 not n22802 ; n22802_not
g69377 not n10391 ; n10391_not
g69378 not n29300 ; n29300_not
g69379 not n10256 ; n10256_not
g69380 not n51062 ; n51062_not
g69381 not n40343 ; n40343_not
g69382 not n23450 ; n23450_not
g69383 not n40316 ; n40316_not
g69384 not n40028 ; n40028_not
g69385 not n40901 ; n40901_not
g69386 not n40325 ; n40325_not
g69387 not n23504 ; n23504_not
g69388 not n23513 ; n23513_not
g69389 not n23522 ; n23522_not
g69390 not n34610 ; n34610_not
g69391 not n23531 ; n23531_not
g69392 not n23540 ; n23540_not
g69393 not n40910 ; n40910_not
g69394 not n26033 ; n26033_not
g69395 not n40406 ; n40406_not
g69396 not n51107 ; n51107_not
g69397 not n13019 ; n13019_not
g69398 not n40415 ; n40415_not
g69399 not n13028 ; n13028_not
g69400 not n50333 ; n50333_not
g69401 not n25241 ; n25241_not
g69402 not n13037 ; n13037_not
g69403 not n13046 ; n13046_not
g69404 not n10319 ; n10319_not
g69405 not n56012 ; n56012_not
g69406 not n13055 ; n13055_not
g69407 not n47120 ; n47120_not
g69408 not n13064 ; n13064_not
g69409 not n10346 ; n10346_not
g69410 not n13073 ; n13073_not
g69411 not n26042 ; n26042_not
g69412 not n13082 ; n13082_not
g69413 not n23027 ; n23027_not
g69414 not n13091 ; n13091_not
g69415 not n26015 ; n26015_not
g69416 not n45500 ; n45500_not
g69417 not n25250 ; n25250_not
g69418 not n40352 ; n40352_not
g69419 not n10265 ; n10265_not
g69420 not n40361 ; n40361_not
g69421 not n12902 ; n12902_not
g69422 not n10382 ; n10382_not
g69423 not n10274 ; n10274_not
g69424 not n12911 ; n12911_not
g69425 not n40370 ; n40370_not
g69426 not n12920 ; n12920_not
g69427 not n34520 ; n34520_not
g69428 not n52511 ; n52511_not
g69429 not n34511 ; n34511_not
g69430 not n10283 ; n10283_not
g69431 not n51134 ; n51134_not
g69432 not n26024 ; n26024_not
g69433 not n10292 ; n10292_not
g69434 not n51125 ; n51125_not
g69435 not n10364 ; n10364_not
g69436 not n56030 ; n56030_not
g69437 not n12632 ; n12632_not
g69438 not n11129 ; n11129_not
g69439 not n24710 ; n24710_not
g69440 not n25160 ; n25160_not
g69441 not n11660 ; n11660_not
g69442 not n40280 ; n40280_not
g69443 not n35060 ; n35060_not
g69444 not n11138 ; n11138_not
g69445 not n25151 ; n25151_not
g69446 not n25142 ; n25142_not
g69447 not n25133 ; n25133_not
g69448 not n52016 ; n52016_not
g69449 not n11147 ; n11147_not
g69450 not n25124 ; n25124_not
g69451 not n25115 ; n25115_not
g69452 not n35051 ; n35051_not
g69453 not n11156 ; n11156_not
g69454 not n40163 ; n40163_not
g69455 not n25106 ; n25106_not
g69456 not n11165 ; n11165_not
g69457 not n25016 ; n25016_not
g69458 not n11093 ; n11093_not
g69459 not n11615 ; n11615_not
g69460 not n25007 ; n25007_not
g69461 not n11624 ; n11624_not
g69462 not n11633 ; n11633_not
g69463 not n24530 ; n24530_not
g69464 not n25214 ; n25214_not
g69465 not n11606 ; n11606_not
g69466 not n11642 ; n11642_not
g69467 not n25205 ; n25205_not
g69468 not n52700 ; n52700_not
g69469 not n11651 ; n11651_not
g69470 not n11741 ; n11741_not
g69471 not n25025 ; n25025_not
g69472 not n11048 ; n11048_not
g69473 not n11219 ; n11219_not
g69474 not n11543 ; n11543_not
g69475 not n40505 ; n40505_not
g69476 not n11750 ; n11750_not
g69477 not n24611 ; n24611_not
g69478 not n11228 ; n11228_not
g69479 not n35024 ; n35024_not
g69480 not n11084 ; n11084_not
g69481 not n52025 ; n52025_not
g69482 not n11237 ; n11237_not
g69483 not n24620 ; n24620_not
g69484 not n56201 ; n56201_not
g69485 not n11246 ; n11246_not
g69486 not n11075 ; n11075_not
g69487 not n40514 ; n40514_not
g69488 not n25313 ; n25313_not
g69489 not n25070 ; n25070_not
g69490 not n35042 ; n35042_not
g69491 not n11174 ; n11174_not
g69492 not n28004 ; n28004_not
g69493 not n11705 ; n11705_not
g69494 not n56210 ; n56210_not
g69495 not n25061 ; n25061_not
g69496 not n11183 ; n11183_not
g69497 not n25052 ; n25052_not
g69498 not n11714 ; n11714_not
g69499 not n11192 ; n11192_not
g69500 not n25043 ; n25043_not
g69501 not n11561 ; n11561_not
g69502 not n11723 ; n11723_not
g69503 not n11039 ; n11039_not
g69504 not n25034 ; n25034_not
g69505 not n11552 ; n11552_not
g69506 not n11732 ; n11732_not
g69507 not n35033 ; n35033_not
g69508 not n35150 ; n35150_not
g69509 not n11390 ; n11390_not
g69510 not n11381 ; n11381_not
g69511 not n35114 ; n35114_not
g69512 not n11372 ; n11372_not
g69513 not n11453 ; n11453_not
g69514 not n24431 ; n24431_not
g69515 not n11363 ; n11363_not
g69516 not n11462 ; n11462_not
g69517 not n11354 ; n11354_not
g69518 not n11345 ; n11345_not
g69519 not n11336 ; n11336_not
g69520 not n11327 ; n11327_not
g69521 not n11480 ; n11480_not
g69522 not n10904 ; n10904_not
g69523 not n35141 ; n35141_not
g69524 not n10913 ; n10913_not
g69525 not n35132 ; n35132_not
g69526 not n24440 ; n24440_not
g69527 not n35123 ; n35123_not
g69528 not n11417 ; n11417_not
g69529 not n11426 ; n11426_not
g69530 not n11408 ; n11408_not
g69531 not n11435 ; n11435_not
g69532 not n11570 ; n11570_not
g69533 not n25232 ; n25232_not
g69534 not n24521 ; n24521_not
g69535 not n11318 ; n11318_not
g69536 not n52007 ; n52007_not
g69537 not n11309 ; n11309_not
g69538 not n35105 ; n35105_not
g69539 not n10940 ; n10940_not
g69540 not n11291 ; n11291_not
g69541 not n11282 ; n11282_not
g69542 not n11507 ; n11507_not
g69543 not n11273 ; n11273_not
g69544 not n11264 ; n11264_not
g69545 not n11255 ; n11255_not
g69546 not n11525 ; n11525_not
g69547 not n12137 ; n12137_not
g69548 not n29003 ; n29003_not
g69549 not n12155 ; n12155_not
g69550 not n24404 ; n24404_not
g69551 not n37103 ; n37103_not
g69552 not n56021 ; n56021_not
g69553 not n12173 ; n12173_not
g69554 not n40613 ; n40613_not
g69555 not n12182 ; n12182_not
g69556 not n29021 ; n29021_not
g69557 not n10841 ; n10841_not
g69558 not n40622 ; n40622_not
g69559 not n10832 ; n10832_not
g69560 not n10355 ; n10355_not
g69561 not n24350 ; n24350_not
g69562 not n24341 ; n24341_not
g69563 not n52133 ; n52133_not
g69564 not n52142 ; n52142_not
g69565 not n52151 ; n52151_not
g69566 not n12065 ; n12065_not
g69567 not n35330 ; n35330_not
g69568 not n24503 ; n24503_not
g69569 not n52160 ; n52160_not
g69570 not n40604 ; n40604_not
g69571 not n25601 ; n25601_not
g69572 not n25610 ; n25610_not
g69573 not n51017 ; n51017_not
g69574 not n40253 ; n40253_not
g69575 not n12128 ; n12128_not
g69576 not n25700 ; n25700_not
g69577 not n52223 ; n52223_not
g69578 not n35312 ; n35312_not
g69579 not n44330 ; n44330_not
g69580 not n24260 ; n24260_not
g69581 not n25421 ; n25421_not
g69582 not n24251 ; n24251_not
g69583 not n40262 ; n40262_not
g69584 not n24242 ; n24242_not
g69585 not n45041 ; n45041_not
g69586 not n10760 ; n10760_not
g69587 not n52232 ; n52232_not
g69588 not n24233 ; n24233_not
g69589 not n23702 ; n23702_not
g69590 not n24224 ; n24224_not
g69591 not n10751 ; n10751_not
g69592 not n56120 ; n56120_not
g69593 not n28400 ; n28400_not
g69594 not n24332 ; n24332_not
g69595 not n10823 ; n10823_not
g69596 not n24323 ; n24323_not
g69597 not n24314 ; n24314_not
g69598 not n10814 ; n10814_not
g69599 not n12146 ; n12146_not
g69600 not n40640 ; n40640_not
g69601 not n24305 ; n24305_not
g69602 not n10805 ; n10805_not
g69603 not n52205 ; n52205_not
g69604 not n45050 ; n45050_not
g69605 not n40631 ; n40631_not
g69606 not n25430 ; n25430_not
g69607 not n52214 ; n52214_not
g69608 not n35321 ; n35321_not
g69609 not n11840 ; n11840_not
g69610 not n40532 ; n40532_not
g69611 not n28031 ; n28031_not
g69612 not n52061 ; n52061_not
g69613 not n40541 ; n40541_not
g69614 not n52070 ; n52070_not
g69615 not n28040 ; n28040_not
g69616 not n40550 ; n40550_not
g69617 not n37013 ; n37013_not
g69618 not n52034 ; n52034_not
g69619 not n35015 ; n35015_not
g69620 not n40208 ; n40208_not
g69621 not n35006 ; n35006_not
g69622 not n52043 ; n52043_not
g69623 not n11516 ; n11516_not
g69624 not n11804 ; n11804_not
g69625 not n11813 ; n11813_not
g69626 not n52052 ; n52052_not
g69627 not n24800 ; n24800_not
g69628 not n11822 ; n11822_not
g69629 not n25403 ; n25403_not
g69630 not n40523 ; n40523_not
g69631 not n11831 ; n11831_not
g69632 not n35240 ; n35240_not
g69633 not n37031 ; n37031_not
g69634 not n52115 ; n52115_not
g69635 not n11930 ; n11930_not
g69636 not n37040 ; n37040_not
g69637 not n10922 ; n10922_not
g69638 not n28112 ; n28112_not
g69639 not n25511 ; n25511_not
g69640 not n52124 ; n52124_not
g69641 not n11471 ; n11471_not
g69642 not n52610 ; n52610_not
g69643 not n52106 ; n52106_not
g69644 not n40118 ; n40118_not
g69645 not n48002 ; n48002_not
g69646 not n11903 ; n11903_not
g69647 not n24701 ; n24701_not
g69648 not n11912 ; n11912_not
g69649 not n25520 ; n25520_not
g69650 not n11921 ; n11921_not
g69651 not n36212 ; n36212_not
g69652 not n27005 ; n27005_not
g69653 not n14702 ; n14702_not
g69654 not n21470 ; n21470_not
g69655 not n50315 ; n50315_not
g69656 not n14711 ; n14711_not
g69657 not n30146 ; n30146_not
g69658 not n57110 ; n57110_not
g69659 not n46202 ; n46202_not
g69660 not n14720 ; n14720_not
g69661 not n49010 ; n49010_not
g69662 not n44600 ; n44600_not
g69663 not n21452 ; n21452_not
g69664 not n36113 ; n36113_not
g69665 not n21434 ; n21434_not
g69666 not n46211 ; n46211_not
g69667 not n21425 ; n21425_not
g69668 not n43070 ; n43070_not
g69669 not n55013 ; n55013_not
g69670 not n21407 ; n21407_not
g69671 not n14621 ; n14621_not
g69672 not n21551 ; n21551_not
g69673 not n14540 ; n14540_not
g69674 not n14630 ; n14630_not
g69675 not n21542 ; n21542_not
g69676 not n21524 ; n21524_not
g69677 not n14531 ; n14531_not
g69678 not n36410 ; n36410_not
g69679 not n21515 ; n21515_not
g69680 not n39110 ; n39110_not
g69681 not n14522 ; n14522_not
g69682 not n36401 ; n36401_not
g69683 not n48200 ; n48200_not
g69684 not n45014 ; n45014_not
g69685 not n33701 ; n33701_not
g69686 not n36104 ; n36104_not
g69687 not n27014 ; n27014_not
g69688 not n21317 ; n21317_not
g69689 not n14405 ; n14405_not
g69690 not n27032 ; n27032_not
g69691 not n43610 ; n43610_not
g69692 not n27041 ; n27041_not
g69693 not n48011 ; n48011_not
g69694 not n36041 ; n36041_not
g69695 not n43601 ; n43601_not
g69696 not n21290 ; n21290_not
g69697 not n14900 ; n14900_not
g69698 not n33251 ; n33251_not
g69699 not n21272 ; n21272_not
g69700 not n21254 ; n21254_not
g69701 not n21263 ; n21263_not
g69702 not n33242 ; n33242_not
g69703 not n50324 ; n50324_not
g69704 not n30074 ; n30074_not
g69705 not n14450 ; n14450_not
g69706 not n21380 ; n21380_not
g69707 not n49001 ; n49001_not
g69708 not n14441 ; n14441_not
g69709 not n46220 ; n46220_not
g69710 not n14801 ; n14801_not
g69711 not n36122 ; n36122_not
g69712 not n14810 ; n14810_not
g69713 not n21362 ; n21362_not
g69714 not n14432 ; n14432_not
g69715 not n33611 ; n33611_not
g69716 not n21344 ; n21344_not
g69717 not n21335 ; n21335_not
g69718 not n46301 ; n46301_not
g69719 not n26150 ; n26150_not
g69720 not n21812 ; n21812_not
g69721 not n21803 ; n21803_not
g69722 not n30128 ; n30128_not
g69723 not n46112 ; n46112_not
g69724 not n14414 ; n14414_not
g69725 not n21740 ; n21740_not
g69726 not n41207 ; n41207_not
g69727 not n21731 ; n21731_not
g69728 not n46103 ; n46103_not
g69729 not n21911 ; n21911_not
g69730 not n51701 ; n51701_not
g69731 not n21902 ; n21902_not
g69732 not n30038 ; n30038_not
g69733 not n46121 ; n46121_not
g69734 not n41171 ; n41171_not
g69735 not n46130 ; n46130_not
g69736 not n30029 ; n30029_not
g69737 not n39200 ; n39200_not
g69738 not n21353 ; n21353_not
g69739 not n50225 ; n50225_not
g69740 not n41180 ; n41180_not
g69741 not n14342 ; n14342_not
g69742 not n21830 ; n21830_not
g69743 not n21821 ; n21821_not
g69744 not n14351 ; n14351_not
g69745 not n26105 ; n26105_not
g69746 not n21632 ; n21632_not
g69747 not n21623 ; n21623_not
g69748 not n21614 ; n21614_not
g69749 not n21605 ; n21605_not
g69750 not n33062 ; n33062_not
g69751 not n41225 ; n41225_not
g69752 not n14603 ; n14603_not
g69753 not n30119 ; n30119_not
g69754 not n14612 ; n14612_not
g69755 not n21560 ; n21560_not
g69756 not n33710 ; n33710_not
g69757 not n21722 ; n21722_not
g69758 not n57002 ; n57002_not
g69759 not n53303 ; n53303_not
g69760 not n21713 ; n21713_not
g69761 not n57011 ; n57011_not
g69762 not n21704 ; n21704_not
g69763 not n30155 ; n30155_not
g69764 not n21443 ; n21443_not
g69765 not n50270 ; n50270_not
g69766 not n14504 ; n14504_not
g69767 not n30164 ; n30164_not
g69768 not n41216 ; n41216_not
g69769 not n57020 ; n57020_not
g69770 not n49100 ; n49100_not
g69771 not n21650 ; n21650_not
g69772 not n21641 ; n21641_not
g69773 not n15125 ; n15125_not
g69774 not n33143 ; n33143_not
g69775 not n20930 ; n20930_not
g69776 not n33152 ; n33152_not
g69777 not n33332 ; n33332_not
g69778 not n20921 ; n20921_not
g69779 not n33161 ; n33161_not
g69780 not n30326 ; n30326_not
g69781 not n33170 ; n33170_not
g69782 not n20912 ; n20912_not
g69783 not n27401 ; n27401_not
g69784 not n33314 ; n33314_not
g69785 not n20903 ; n20903_not
g69786 not n33305 ; n33305_not
g69787 not n55103 ; n55103_not
g69788 not n33206 ; n33206_not
g69789 not n27122 ; n27122_not
g69790 not n33215 ; n33215_not
g69791 not n48101 ; n48101_not
g69792 not n33080 ; n33080_not
g69793 not n27230 ; n27230_not
g69794 not n46310 ; n46310_not
g69795 not n27212 ; n27212_not
g69796 not n48110 ; n48110_not
g69797 not n43160 ; n43160_not
g69798 not n33107 ; n33107_not
g69799 not n15143 ; n15143_not
g69800 not n39020 ; n39020_not
g69801 not n33116 ; n33116_not
g69802 not n33350 ; n33350_not
g69803 not n41315 ; n41315_not
g69804 not n15134 ; n15134_not
g69805 not n30317 ; n30317_not
g69806 not n36203 ; n36203_not
g69807 not n33125 ; n33125_not
g69808 not n27410 ; n27410_not
g69809 not n33134 ; n33134_not
g69810 not n41360 ; n41360_not
g69811 not n27320 ; n27320_not
g69812 not n20831 ; n20831_not
g69813 not n30335 ; n30335_not
g69814 not n15053 ; n15053_not
g69815 not n15044 ; n15044_not
g69816 not n20822 ; n20822_not
g69817 not n20813 ; n20813_not
g69818 not n30353 ; n30353_not
g69819 not n43430 ; n43430_not
g69820 not n15035 ; n15035_not
g69821 not n20804 ; n20804_not
g69822 not n27131 ; n27131_not
g69823 not n45140 ; n45140_not
g69824 not n50306 ; n50306_not
g69825 not n27140 ; n27140_not
g69826 not n30362 ; n30362_not
g69827 not n30371 ; n30371_not
g69828 not n33224 ; n33224_not
g69829 not n33233 ; n33233_not
g69830 not n15080 ; n15080_not
g69831 not n36221 ; n36221_not
g69832 not n27302 ; n27302_not
g69833 not n20723 ; n20723_not
g69834 not n27311 ; n27311_not
g69835 not n30344 ; n30344_not
g69836 not n33260 ; n33260_not
g69837 not n20840 ; n20840_not
g69838 not n46400 ; n46400_not
g69839 not n27104 ; n27104_not
g69840 not n21182 ; n21182_not
g69841 not n33512 ; n33512_not
g69842 not n20543 ; n20543_not
g69843 not n30272 ; n30272_not
g69844 not n36320 ; n36320_not
g69845 not n21173 ; n21173_not
g69846 not n33503 ; n33503_not
g69847 not n33323 ; n33323_not
g69848 not n15062 ; n15062_not
g69849 not n21164 ; n21164_not
g69850 not n41270 ; n41270_not
g69851 not n21155 ; n21155_not
g69852 not n21146 ; n21146_not
g69853 not n50351 ; n50351_not
g69854 not n21137 ; n21137_not
g69855 not n27050 ; n27050_not
g69856 not n21245 ; n21245_not
g69857 not n50342 ; n50342_not
g69858 not n14360 ; n14360_not
g69859 not n21236 ; n21236_not
g69860 not n43115 ; n43115_not
g69861 not n21227 ; n21227_not
g69862 not n37004 ; n37004_not
g69863 not n21218 ; n21218_not
g69864 not n33530 ; n33530_not
g69865 not n21209 ; n21209_not
g69866 not n33521 ; n33521_not
g69867 not n15017 ; n15017_not
g69868 not n21191 ; n21191_not
g69869 not n21056 ; n21056_not
g69870 not n33422 ; n33422_not
g69871 not n43520 ; n43520_not
g69872 not n21047 ; n21047_not
g69873 not n21038 ; n21038_not
g69874 not n33413 ; n33413_not
g69875 not n21029 ; n21029_not
g69876 not n33404 ; n33404_not
g69877 not n43511 ; n43511_not
g69878 not n20633 ; n20633_not
g69879 not n50360 ; n50360_not
g69880 not n27221 ; n27221_not
g69881 not n33071 ; n33071_not
g69882 not n15170 ; n15170_not
g69883 not n43502 ; n43502_not
g69884 not n27500 ; n27500_not
g69885 not n21128 ; n21128_not
g69886 not n15107 ; n15107_not
g69887 not n21119 ; n21119_not
g69888 not n36131 ; n36131_not
g69889 not n36311 ; n36311_not
g69890 not n15152 ; n15152_not
g69891 not n21092 ; n21092_not
g69892 not n21083 ; n21083_not
g69893 not n33440 ; n33440_not
g69894 not n21074 ; n21074_not
g69895 not n36302 ; n36302_not
g69896 not n21065 ; n21065_not
g69897 not n33431 ; n33431_not
g69898 not n22145 ; n22145_not
g69899 not n22091 ; n22091_not
g69900 not n50135 ; n50135_not
g69901 not n46004 ; n46004_not
g69902 not n50072 ; n50072_not
g69903 not n22154 ; n22154_not
g69904 not n46013 ; n46013_not
g69905 not n22406 ; n22406_not
g69906 not n34205 ; n34205_not
g69907 not n13901 ; n13901_not
g69908 not n35600 ; n35600_not
g69909 not n22136 ; n22136_not
g69910 not n34061 ; n34061_not
g69911 not n26312 ; n26312_not
g69912 not n34214 ; n34214_not
g69913 not n34250 ; n34250_not
g69914 not n22181 ; n22181_not
g69915 not n22172 ; n22172_not
g69916 not n41090 ; n41090_not
g69917 not n26330 ; n26330_not
g69918 not n34052 ; n34052_not
g69919 not n22109 ; n22109_not
g69920 not n22703 ; n22703_not
g69921 not n46022 ; n46022_not
g69922 not n34043 ; n34043_not
g69923 not n51800 ; n51800_not
g69924 not n22712 ; n22712_not
g69925 not n28130 ; n28130_not
g69926 not n22235 ; n22235_not
g69927 not n46031 ; n46031_not
g69928 not n30056 ; n30056_not
g69929 not n50054 ; n50054_not
g69930 not n34133 ; n34133_not
g69931 not n13226 ; n13226_not
g69932 not n41081 ; n41081_not
g69933 not n22127 ; n22127_not
g69934 not n22082 ; n22082_not
g69935 not n33620 ; n33620_not
g69936 not n22415 ; n22415_not
g69937 not n50081 ; n50081_not
g69938 not n30047 ; n30047_not
g69939 not n21533 ; n21533_not
g69940 not n34070 ; n34070_not
g69941 not n47210 ; n47210_not
g69942 not n22271 ; n22271_not
g69943 not n13631 ; n13631_not
g69944 not n26501 ; n26501_not
g69945 not n22604 ; n22604_not
g69946 not n22631 ; n22631_not
g69947 not n22352 ; n22352_not
g69948 not n22262 ; n22262_not
g69949 not n26321 ; n26321_not
g69950 not n22361 ; n22361_not
g69951 not n22334 ; n22334_not
g69952 not n22613 ; n22613_not
g69953 not n34232 ; n34232_not
g69954 not n44501 ; n44501_not
g69955 not n13640 ; n13640_not
g69956 not n22280 ; n22280_not
g69957 not n22325 ; n22325_not
g69958 not n22343 ; n22343_not
g69959 not n22622 ; n22622_not
g69960 not n22316 ; n22316_not
g69961 not n22370 ; n22370_not
g69962 not n22226 ; n22226_not
g69963 not n50801 ; n50801_not
g69964 not n34025 ; n34025_not
g69965 not n22217 ; n22217_not
g69966 not n50063 ; n50063_not
g69967 not n41126 ; n41126_not
g69968 not n13910 ; n13910_not
g69969 not n41135 ; n41135_not
g69970 not n34115 ; n34115_not
g69971 not n34223 ; n34223_not
g69972 not n50090 ; n50090_not
g69973 not n13181 ; n13181_not
g69974 not n34241 ; n34241_not
g69975 not n13622 ; n13622_not
g69976 not n22640 ; n22640_not
g69977 not n50810 ; n50810_not
g69978 not n13613 ; n13613_not
g69979 not n22244 ; n22244_not
g69980 not n26510 ; n26510_not
g69981 not n13604 ; n13604_not
g69982 not n22532 ; n22532_not
g69983 not n26600 ; n26600_not
g69984 not n30083 ; n30083_not
g69985 not n13802 ; n13802_not
g69986 not n22037 ; n22037_not
g69987 not n44402 ; n44402_not
g69988 not n41153 ; n41153_not
g69989 not n34151 ; n34151_not
g69990 not n41063 ; n41063_not
g69991 not n13505 ; n13505_not
g69992 not n22451 ; n22451_not
g69993 not n22019 ; n22019_not
g69994 not n41144 ; n41144_not
g69995 not n26240 ; n26240_not
g69996 not n22541 ; n22541_not
g69997 not n13820 ; n13820_not
g69998 not n34304 ; n34304_not
g69999 not n26411 ; n26411_not
g70000 not n13271 ; n13271_not
g70001 not n13811 ; n13811_not
g70002 not n34160 ; n34160_not
g70003 not n46040 ; n46040_not
g70004 not n26402 ; n26402_not
g70005 not n41117 ; n41117_not
g70006 not n21920 ; n21920_not
g70007 not n13460 ; n13460_not
g70008 not n34322 ; n34322_not
g70009 not n22505 ; n22505_not
g70010 not n22190 ; n22190_not
g70011 not n22811 ; n22811_not
g70012 not n34106 ; n34106_not
g70013 not n30065 ; n30065_not
g70014 not n22460 ; n22460_not
g70015 not n41162 ; n41162_not
g70016 not n22523 ; n22523_not
g70017 not n34313 ; n34313_not
g70018 not n21308 ; n21308_not
g70019 not n22514 ; n22514_not
g70020 not n41072 ; n41072_not
g70021 not n13523 ; n13523_not
g70022 not n22433 ; n22433_not
g70023 not n22064 ; n22064_not
g70024 not n41108 ; n41108_not
g70025 not n13703 ; n13703_not
g70026 not n22055 ; n22055_not
g70027 not n13532 ; n13532_not
g70028 not n34142 ; n34142_not
g70029 not n26420 ; n26420_not
g70030 not n22730 ; n22730_not
g70031 not n13541 ; n13541_not
g70032 not n28013 ; n28013_not
g70033 not n22721 ; n22721_not
g70034 not n22424 ; n22424_not
g70035 not n13550 ; n13550_not
g70036 not n22028 ; n22028_not
g70037 not n22550 ; n22550_not
g70038 not n13712 ; n13712_not
g70039 not n13514 ; n13514_not
g70040 not n22046 ; n22046_not
g70041 not n50180 ; n50180_not
g70042 not n22442 ; n22442_not
g70043 not n31560 ; n31560_not
g70044 not n42036 ; n42036_not
g70045 not n25611 ; n25611_not
g70046 not n31533 ; n31533_not
g70047 not n27141 ; n27141_not
g70048 not n40281 ; n40281_not
g70049 not n25323 ; n25323_not
g70050 not n40209 ; n40209_not
g70051 not n26520 ; n26520_not
g70052 not n31290 ; n31290_not
g70053 not n18033 ; n18033_not
g70054 not n18042 ; n18042_not
g70055 not n31281 ; n31281_not
g70056 not n18060 ; n18060_not
g70057 not n31335 ; n31335_not
g70058 not n31254 ; n31254_not
g70059 not n26511 ; n26511_not
g70060 not n31227 ; n31227_not
g70061 not n31551 ; n31551_not
g70062 not n25305 ; n25305_not
g70063 not n54303 ; n54303_not
g70064 not n26412 ; n26412_not
g70065 not n42333 ; n42333_not
g70066 not n26502 ; n26502_not
g70067 not n28221 ; n28221_not
g70068 not n26043 ; n26043_not
g70069 not n42342 ; n42342_not
g70070 not n25413 ; n25413_not
g70071 not n25215 ; n25215_not
g70072 not n18051 ; n18051_not
g70073 not n18420 ; n18420_not
g70074 not n27240 ; n27240_not
g70075 not n27312 ; n27312_not
g70076 not n28050 ; n28050_not
g70077 not n27501 ; n27501_not
g70078 not n27132 ; n27132_not
g70079 not n18015 ; n18015_not
g70080 not n31542 ; n31542_not
g70081 not n26070 ; n26070_not
g70082 not n42324 ; n42324_not
g70083 not n31326 ; n31326_not
g70084 not n52017 ; n52017_not
g70085 not n25350 ; n25350_not
g70086 not n25602 ; n25602_not
g70087 not n25521 ; n25521_not
g70088 not n18024 ; n18024_not
g70089 not n26430 ; n26430_not
g70090 not n26322 ; n26322_not
g70091 not n45312 ; n45312_not
g70092 not n28041 ; n28041_not
g70093 not n31218 ; n31218_not
g70094 not n26061 ; n26061_not
g70095 not n26331 ; n26331_not
g70096 not n18510 ; n18510_not
g70097 not n39003 ; n39003_not
g70098 not n27303 ; n27303_not
g70099 not n26052 ; n26052_not
g70100 not n52026 ; n52026_not
g70101 not n25341 ; n25341_not
g70102 not n27114 ; n27114_not
g70103 not n26421 ; n26421_not
g70104 not n39030 ; n39030_not
g70105 not n42360 ; n42360_not
g70106 not n28140 ; n28140_not
g70107 not n24711 ; n24711_not
g70108 not n50172 ; n50172_not
g70109 not n40047 ; n40047_not
g70110 not n25710 ; n25710_not
g70111 not n31812 ; n31812_not
g70112 not n39012 ; n39012_not
g70113 not n52062 ; n52062_not
g70114 not n50181 ; n50181_not
g70115 not n26214 ; n26214_not
g70116 not n25206 ; n25206_not
g70117 not n31506 ; n31506_not
g70118 not n52044 ; n52044_not
g70119 not n28131 ; n28131_not
g70120 not n52404 ; n52404_not
g70121 not n31524 ; n31524_not
g70122 not n40065 ; n40065_not
g70123 not n25701 ; n25701_not
g70124 not n40056 ; n40056_not
g70125 not n52413 ; n52413_not
g70126 not n18402 ; n18402_not
g70127 not n42171 ; n42171_not
g70128 not n26232 ; n26232_not
g70129 not n26241 ; n26241_not
g70130 not n27330 ; n27330_not
g70131 not n25152 ; n25152_not
g70132 not n50631 ; n50631_not
g70133 not n42180 ; n42180_not
g70134 not n31029 ; n31029_not
g70135 not n27150 ; n27150_not
g70136 not n54231 ; n54231_not
g70137 not n52053 ; n52053_not
g70138 not n24450 ; n24450_not
g70139 not n31821 ; n31821_not
g70140 not n25800 ; n25800_not
g70141 not n31830 ; n31830_not
g70142 not n25170 ; n25170_not
g70143 not n27321 ; n27321_not
g70144 not n51522 ; n51522_not
g70145 not n51720 ; n51720_not
g70146 not n24441 ; n24441_not
g70147 not n54240 ; n54240_not
g70148 not n40038 ; n40038_not
g70149 not n31308 ; n31308_not
g70150 not n25161 ; n25161_not
g70151 not n28005 ; n28005_not
g70152 not n40029 ; n40029_not
g70153 not n27222 ; n27222_not
g70154 not n26007 ; n26007_not
g70155 not n25620 ; n25620_not
g70156 not n46410 ; n46410_not
g70157 not n25260 ; n25260_not
g70158 not n26106 ; n26106_not
g70159 not n51540 ; n51540_not
g70160 not n25251 ; n25251_not
g70161 not n27420 ; n27420_not
g70162 not n50640 ; n50640_not
g70163 not n31272 ; n31272_not
g70164 not n38013 ; n38013_not
g70165 not n52035 ; n52035_not
g70166 not n26034 ; n26034_not
g70167 not n26403 ; n26403_not
g70168 not n52431 ; n52431_not
g70169 not n27204 ; n27204_not
g70170 not n26025 ; n26025_not
g70171 not n52080 ; n52080_not
g70172 not n28212 ; n28212_not
g70173 not n18006 ; n18006_not
g70174 not n27105 ; n27105_not
g70175 not n42153 ; n42153_not
g70176 not n26016 ; n26016_not
g70177 not n40092 ; n40092_not
g70178 not n31263 ; n31263_not
g70179 not n42162 ; n42162_not
g70180 not n24414 ; n24414_not
g70181 not n26142 ; n26142_not
g70182 not n52071 ; n52071_not
g70183 not n51702 ; n51702_not
g70184 not n44700 ; n44700_not
g70185 not n26151 ; n26151_not
g70186 not n27402 ; n27402_not
g70187 not n28122 ; n28122_not
g70188 not n50604 ; n50604_not
g70189 not n51531 ; n51531_not
g70190 not n40074 ; n40074_not
g70191 not n54204 ; n54204_not
g70192 not n26124 ; n26124_not
g70193 not n25224 ; n25224_not
g70194 not n40083 ; n40083_not
g70195 not n31317 ; n31317_not
g70196 not n25233 ; n25233_not
g70197 not n31515 ; n31515_not
g70198 not n27411 ; n27411_not
g70199 not n28203 ; n28203_not
g70200 not n26304 ; n26304_not
g70201 not n42351 ; n42351_not
g70202 not n52503 ; n52503_not
g70203 not n31362 ; n31362_not
g70204 not n18222 ; n18222_not
g70205 not n41901 ; n41901_not
g70206 not n31650 ; n31650_not
g70207 not n52512 ; n52512_not
g70208 not n18213 ; n18213_not
g70209 not n31182 ; n31182_not
g70210 not n52440 ; n52440_not
g70211 not n40227 ; n40227_not
g70212 not n42054 ; n42054_not
g70213 not n52341 ; n52341_not
g70214 not n42261 ; n42261_not
g70215 not n52530 ; n52530_not
g70216 not n18204 ; n18204_not
g70217 not n25008 ; n25008_not
g70218 not n26115 ; n26115_not
g70219 not n39120 ; n39120_not
g70220 not n31641 ; n31641_not
g70221 not n31605 ; n31605_not
g70222 not n18231 ; n18231_not
g70223 not n52332 ; n52332_not
g70224 not n54411 ; n54411_not
g70225 not n28311 ; n28311_not
g70226 not n42252 ; n42252_not
g70227 not n54330 ; n54330_not
g70228 not n31173 ; n31173_not
g70229 not n52224 ; n52224_not
g70230 not n31407 ; n31407_not
g70231 not n45006 ; n45006_not
g70232 not n51810 ; n51810_not
g70233 not n51630 ; n51630_not
g70234 not n42045 ; n42045_not
g70235 not n45042 ; n45042_not
g70236 not n31425 ; n31425_not
g70237 not n31353 ; n31353_not
g70238 not n24900 ; n24900_not
g70239 not n42117 ; n42117_not
g70240 not n31461 ; n31461_not
g70241 not n42270 ; n42270_not
g70242 not n42018 ; n42018_not
g70243 not n40272 ; n40272_not
g70244 not n52206 ; n52206_not
g70245 not n52350 ; n52350_not
g70246 not n54600 ; n54600_not
g70247 not n45303 ; n45303_not
g70248 not n52422 ; n52422_not
g70249 not n42216 ; n42216_not
g70250 not n54402 ; n54402_not
g70251 not n52215 ; n52215_not
g70252 not n40245 ; n40245_not
g70253 not n25404 ; n25404_not
g70254 not n31434 ; n31434_not
g70255 not n18303 ; n18303_not
g70256 not n40254 ; n40254_not
g70257 not n26700 ; n26700_not
g70258 not n31614 ; n31614_not
g70259 not n40155 ; n40155_not
g70260 not n52314 ; n52314_not
g70261 not n42234 ; n42234_not
g70262 not n25314 ; n25314_not
g70263 not n31371 ; n31371_not
g70264 not n40164 ; n40164_not
g70265 not n25080 ; n25080_not
g70266 not n26160 ; n26160_not
g70267 not n26610 ; n26610_not
g70268 not n45015 ; n45015_not
g70269 not n52260 ; n52260_not
g70270 not n25071 ; n25071_not
g70271 not n42081 ; n42081_not
g70272 not n42225 ; n42225_not
g70273 not n25134 ; n25134_not
g70274 not n31443 ; n31443_not
g70275 not n31380 ; n31380_not
g70276 not n26205 ; n26205_not
g70277 not n45330 ; n45330_not
g70278 not n25125 ; n25125_not
g70279 not n40137 ; n40137_not
g70280 not n52305 ; n52305_not
g70281 not n25116 ; n25116_not
g70282 not n42090 ; n42090_not
g70283 not n51711 ; n51711_not
g70284 not n25107 ; n25107_not
g70285 not n25143 ; n25143_not
g70286 not n52242 ; n52242_not
g70287 not n42243 ; n42243_not
g70288 not n25026 ; n25026_not
g70289 not n42108 ; n42108_not
g70290 not n31632 ; n31632_not
g70291 not n25017 ; n25017_not
g70292 not n54420 ; n54420_not
g70293 not n52233 ; n52233_not
g70294 not n42063 ; n42063_not
g70295 not n18240 ; n18240_not
g70296 not n27600 ; n27600_not
g70297 not n26250 ; n26250_not
g70298 not n25062 ; n25062_not
g70299 not n31623 ; n31623_not
g70300 not n26601 ; n26601_not
g70301 not n51900 ; n51900_not
g70302 not n31416 ; n31416_not
g70303 not n52251 ; n52251_not
g70304 not n25053 ; n25053_not
g70305 not n25044 ; n25044_not
g70306 not n40119 ; n40119_not
g70307 not n42072 ; n42072_not
g70308 not n40182 ; n40182_not
g70309 not n52323 ; n52323_not
g70310 not n25035 ; n25035_not
g70311 not n25530 ; n25530_not
g70312 not n45222 ; n45222_not
g70313 not n27042 ; n27042_not
g70314 not n51801 ; n51801_not
g70315 not n54501 ; n54501_not
g70316 not n51603 ; n51603_not
g70317 not n18330 ; n18330_not
g70318 not n52134 ; n52134_not
g70319 not n18105 ; n18105_not
g70320 not n42135 ; n42135_not
g70321 not n52602 ; n52602_not
g70322 not n24720 ; n24720_not
g70323 not n27006 ; n27006_not
g70324 not n52125 ; n52125_not
g70325 not n42306 ; n42306_not
g70326 not n45321 ; n45321_not
g70327 not n31209 ; n31209_not
g70328 not n27024 ; n27024_not
g70329 not n28023 ; n28023_not
g70330 not n25431 ; n25431_not
g70331 not n52107 ; n52107_not
g70332 not n42315 ; n42315_not
g70333 not n54321 ; n54321_not
g70334 not n31731 ; n31731_not
g70335 not n27510 ; n27510_not
g70336 not n54510 ; n54510_not
g70337 not n25503 ; n25503_not
g70338 not n42207 ; n42207_not
g70339 not n52116 ; n52116_not
g70340 not n27051 ; n27051_not
g70341 not n26340 ; n26340_not
g70342 not n42144 ; n42144_not
g70343 not n52620 ; n52620_not
g70344 not n52008 ; n52008_not
g70345 not n31470 ; n31470_not
g70346 not n31344 ; n31344_not
g70347 not n40218 ; n40218_not
g70348 not n28500 ; n28500_not
g70349 not n27060 ; n27060_not
g70350 not n25440 ; n25440_not
g70351 not n50622 ; n50622_not
g70352 not n42126 ; n42126_not
g70353 not n41433 ; n41433_not
g70354 not n28401 ; n28401_not
g70355 not n40263 ; n40263_not
g70356 not n27015 ; n27015_not
g70357 not n52170 ; n52170_not
g70358 not n50163 ; n50163_not
g70359 not n18150 ; n18150_not
g70360 not n17700 ; n17700_not
g70361 not n51621 ; n51621_not
g70362 not n18312 ; n18312_not
g70363 not n46500 ; n46500_not
g70364 not n42027 ; n42027_not
g70365 not n28320 ; n28320_not
g70366 not n52152 ; n52152_not
g70367 not n18123 ; n18123_not
g70368 not n47301 ; n47301_not
g70369 not n39102 ; n39102_not
g70370 not n52143 ; n52143_not
g70371 not n31713 ; n31713_not
g70372 not n18114 ; n18114_not
g70373 not n45060 ; n45060_not
g70374 not n18141 ; n18141_not
g70375 not n18321 ; n18321_not
g70376 not n52161 ; n52161_not
g70377 not n24810 ; n24810_not
g70378 not n50613 ; n50613_not
g70379 not n45600 ; n45600_not
g70380 not n28410 ; n28410_not
g70381 not n51612 ; n51612_not
g70382 not n24801 ; n24801_not
g70383 not n18132 ; n18132_not
g70384 not n31704 ; n31704_not
g70385 not n45051 ; n45051_not
g70386 not n20319 ; n20319_not
g70387 not n22227 ; n22227_not
g70388 not n50802 ; n50802_not
g70389 not n22236 ; n22236_not
g70390 not n50046 ; n50046_not
g70391 not n22254 ; n22254_not
g70392 not n50811 ; n50811_not
g70393 not n22272 ; n22272_not
g70394 not n22281 ; n22281_not
g70395 not n38220 ; n38220_not
g70396 not n41451 ; n41451_not
g70397 not n22317 ; n22317_not
g70398 not n22290 ; n22290_not
g70399 not n22326 ; n22326_not
g70400 not n30471 ; n30471_not
g70401 not n22119 ; n22119_not
g70402 not n30039 ; n30039_not
g70403 not n41442 ; n41442_not
g70404 not n20346 ; n20346_not
g70405 not n22137 ; n22137_not
g70406 not n22146 ; n22146_not
g70407 not n53520 ; n53520_not
g70408 not n20337 ; n20337_not
g70409 not n50073 ; n50073_not
g70410 not n38211 ; n38211_not
g70411 not n22164 ; n22164_not
g70412 not n22182 ; n22182_not
g70413 not n41136 ; n41136_not
g70414 not n22191 ; n22191_not
g70415 not n20328 ; n20328_not
g70416 not n22209 ; n22209_not
g70417 not n22416 ; n22416_not
g70418 not n20274 ; n20274_not
g70419 not n22425 ; n22425_not
g70420 not n22434 ; n22434_not
g70421 not n22443 ; n22443_not
g70422 not n41460 ; n41460_not
g70423 not n20265 ; n20265_not
g70424 not n22452 ; n22452_not
g70425 not n22461 ; n22461_not
g70426 not n41118 ; n41118_not
g70427 not n22470 ; n22470_not
g70428 not n20256 ; n20256_not
g70429 not n50730 ; n50730_not
g70430 not n40551 ; n40551_not
g70431 not n22335 ; n22335_not
g70432 not n22344 ; n22344_not
g70433 not n30480 ; n30480_not
g70434 not n20292 ; n20292_not
g70435 not n22353 ; n22353_not
g70436 not n22362 ; n22362_not
g70437 not n22371 ; n22371_not
g70438 not n41127 ; n41127_not
g70439 not n20283 ; n20283_not
g70440 not n22380 ; n22380_not
g70441 not n47202 ; n47202_not
g70442 not n40560 ; n40560_not
g70443 not n22245 ; n22245_not
g70444 not n22407 ; n22407_not
g70445 not n53205 ; n53205_not
g70446 not n21354 ; n21354_not
g70447 not n40614 ; n40614_not
g70448 not n21345 ; n21345_not
g70449 not n53214 ; n53214_not
g70450 not n41172 ; n41172_not
g70451 not n30453 ; n30453_not
g70452 not n40605 ; n40605_not
g70453 not n53223 ; n53223_not
g70454 not n20391 ; n20391_not
g70455 not n21903 ; n21903_not
g70456 not n53232 ; n53232_not
g70457 not n21912 ; n21912_not
g70458 not n21408 ; n21408_not
g70459 not n30147 ; n30147_not
g70460 not n20418 ; n20418_not
g70461 not n40650 ; n40650_not
g70462 not n50091 ; n50091_not
g70463 not n30138 ; n30138_not
g70464 not n21390 ; n21390_not
g70465 not n41190 ; n41190_not
g70466 not n40623 ; n40623_not
g70467 not n20409 ; n20409_not
g70468 not n21804 ; n21804_not
g70469 not n30264 ; n30264_not
g70470 not n21813 ; n21813_not
g70471 not n21822 ; n21822_not
g70472 not n21831 ; n21831_not
g70473 not n41181 ; n41181_not
g70474 not n21363 ; n21363_not
g70475 not n21840 ; n21840_not
g70476 not n53241 ; n53241_not
g70477 not n20373 ; n20373_not
g70478 not n22029 ; n22029_not
g70479 not n22047 ; n22047_not
g70480 not n22056 ; n22056_not
g70481 not n50082 ; n50082_not
g70482 not n20364 ; n20364_not
g70483 not n30066 ; n30066_not
g70484 not n22074 ; n22074_not
g70485 not n47220 ; n47220_not
g70486 not n38202 ; n38202_not
g70487 not n30057 ; n30057_not
g70488 not n53511 ; n53511_not
g70489 not n22092 ; n22092_not
g70490 not n20355 ; n20355_not
g70491 not n30048 ; n30048_not
g70492 not n21318 ; n21318_not
g70493 not n21921 ; n21921_not
g70494 not n21309 ; n21309_not
g70495 not n21930 ; n21930_not
g70496 not n45141 ; n45141_not
g70497 not n41163 ; n41163_not
g70498 not n52800 ; n52800_not
g70499 not n30093 ; n30093_not
g70500 not n30075 ; n30075_not
g70501 not n53250 ; n53250_not
g70502 not n41154 ; n41154_not
g70503 not n20382 ; n20382_not
g70504 not n30084 ; n30084_not
g70505 not n21273 ; n21273_not
g70506 not n41145 ; n41145_not
g70507 not n22623 ; n22623_not
g70508 not n22614 ; n22614_not
g70509 not n20139 ; n20139_not
g70510 not n22911 ; n22911_not
g70511 not n22605 ; n22605_not
g70512 not n41028 ; n41028_not
g70513 not n40461 ; n40461_not
g70514 not n22560 ; n22560_not
g70515 not n22551 ; n22551_not
g70516 not n22542 ; n22542_not
g70517 not n22533 ; n22533_not
g70518 not n41019 ; n41019_not
g70519 not n22524 ; n22524_not
g70520 not n50460 ; n50460_not
g70521 not n30345 ; n30345_not
g70522 not n22515 ; n22515_not
g70523 not n22704 ; n22704_not
g70524 not n20157 ; n20157_not
g70525 not n50514 ; n50514_not
g70526 not n41037 ; n41037_not
g70527 not n40740 ; n40740_not
g70528 not n41406 ; n41406_not
g70529 not n40470 ; n40470_not
g70530 not n50505 ; n50505_not
g70531 not n51009 ; n51009_not
g70532 not n53601 ; n53601_not
g70533 not n38031 ; n38031_not
g70534 not n20148 ; n20148_not
g70535 not n22650 ; n22650_not
g70536 not n22641 ; n22641_not
g70537 not n51018 ; n51018_not
g70538 not n22632 ; n22632_not
g70539 not n45150 ; n45150_not
g70540 not n23046 ; n23046_not
g70541 not n50433 ; n50433_not
g70542 not n23064 ; n23064_not
g70543 not n50424 ; n50424_not
g70544 not n23073 ; n23073_not
g70545 not n23082 ; n23082_not
g70546 not n30543 ; n30543_not
g70547 not n20094 ; n20094_not
g70548 not n51054 ; n51054_not
g70549 not n40443 ; n40443_not
g70550 not n51036 ; n51036_not
g70551 not n22506 ; n22506_not
g70552 not n40452 ; n40452_not
g70553 not n50451 ; n50451_not
g70554 not n50442 ; n50442_not
g70555 not n23019 ; n23019_not
g70556 not n53610 ; n53610_not
g70557 not n23028 ; n23028_not
g70558 not n20229 ; n20229_not
g70559 not n40533 ; n40533_not
g70560 not n30507 ; n30507_not
g70561 not n41091 ; n41091_not
g70562 not n40524 ; n40524_not
g70563 not n41082 ; n41082_not
g70564 not n40515 ; n40515_not
g70565 not n50721 ; n50721_not
g70566 not n50712 ; n50712_not
g70567 not n20247 ; n20247_not
g70568 not n50703 ; n50703_not
g70569 not n41109 ; n41109_not
g70570 not n20238 ; n20238_not
g70571 not n50901 ; n50901_not
g70572 not n22155 ; n22155_not
g70573 not n40542 ; n40542_not
g70574 not n20175 ; n20175_not
g70575 not n38301 ; n38301_not
g70576 not n30525 ; n30525_not
g70577 not n41055 ; n41055_not
g70578 not n22821 ; n22821_not
g70579 not n38310 ; n38310_not
g70580 not n20166 ; n20166_not
g70581 not n50550 ; n50550_not
g70582 not n41046 ; n41046_not
g70583 not n22740 ; n22740_not
g70584 not n50541 ; n50541_not
g70585 not n22731 ; n22731_not
g70586 not n22722 ; n22722_not
g70587 not n50532 ; n50532_not
g70588 not n22713 ; n22713_not
g70589 not n40731 ; n40731_not
g70590 not n50523 ; n50523_not
g70591 not n22065 ; n22065_not
g70592 not n41073 ; n41073_not
g70593 not n20193 ; n20193_not
g70594 not n40506 ; n40506_not
g70595 not n20184 ; n20184_not
g70596 not n38040 ; n38040_not
g70597 not n41064 ; n41064_not
g70598 not n40722 ; n40722_not
g70599 not n21093 ; n21093_not
g70600 not n30219 ; n30219_not
g70601 not n20625 ; n20625_not
g70602 not n53034 ; n53034_not
g70603 not n20580 ; n20580_not
g70604 not n30228 ; n30228_not
g70605 not n30282 ; n30282_not
g70606 not n21129 ; n21129_not
g70607 not n53043 ; n53043_not
g70608 not n21138 ; n21138_not
g70609 not n30237 ; n30237_not
g70610 not n20652 ; n20652_not
g70611 not n53007 ; n53007_not
g70612 not n21039 ; n21039_not
g70613 not n53016 ; n53016_not
g70614 not n21048 ; n21048_not
g70615 not n21057 ; n21057_not
g70616 not n21066 ; n21066_not
g70617 not n53025 ; n53025_not
g70618 not n21075 ; n21075_not
g70619 not n21084 ; n21084_not
g70620 not n20634 ; n20634_not
g70621 not n41280 ; n41280_not
g70622 not n53061 ; n53061_not
g70623 not n21219 ; n21219_not
g70624 not n41262 ; n41262_not
g70625 not n21228 ; n21228_not
g70626 not n21237 ; n21237_not
g70627 not n30408 ; n30408_not
g70628 not n20508 ; n20508_not
g70629 not n21246 ; n21246_not
g70630 not n21147 ; n21147_not
g70631 not n21156 ; n21156_not
g70632 not n20553 ; n20553_not
g70633 not n53052 ; n53052_not
g70634 not n21165 ; n21165_not
g70635 not n20544 ; n20544_not
g70636 not n30246 ; n30246_not
g70637 not n21174 ; n21174_not
g70638 not n20607 ; n20607_not
g70639 not n21183 ; n21183_not
g70640 not n20535 ; n20535_not
g70641 not n21192 ; n21192_not
g70642 not n20058 ; n20058_not
g70643 not n45132 ; n45132_not
g70644 not n20841 ; n20841_not
g70645 not n20742 ; n20742_not
g70646 not n20724 ; n20724_not
g70647 not n20850 ; n20850_not
g70648 not n20067 ; n20067_not
g70649 not n41352 ; n41352_not
g70650 not n20076 ; n20076_not
g70651 not n20715 ; n20715_not
g70652 not n20085 ; n20085_not
g70653 not n30165 ; n30165_not
g70654 not n30192 ; n30192_not
g70655 not n53430 ; n53430_not
g70656 not n41343 ; n41343_not
g70657 not n53421 ; n53421_not
g70658 not n30309 ; n30309_not
g70659 not n30183 ; n30183_not
g70660 not n20760 ; n20760_not
g70661 not n30372 ; n30372_not
g70662 not n30363 ; n30363_not
g70663 not n30318 ; n30318_not
g70664 not n30174 ; n30174_not
g70665 not n41370 ; n41370_not
g70666 not n30354 ; n30354_not
g70667 not n20805 ; n20805_not
g70668 not n20814 ; n20814_not
g70669 not n20823 ; n20823_not
g70670 not n20049 ; n20049_not
g70671 not n30156 ; n30156_not
g70672 not n20832 ; n20832_not
g70673 not n20733 ; n20733_not
g70674 not n41307 ; n41307_not
g70675 not n30390 ; n30390_not
g70676 not n20670 ; n20670_not
g70677 not n53403 ; n53403_not
g70678 not n20643 ; n20643_not
g70679 not n20904 ; n20904_not
g70680 not n20913 ; n20913_not
g70681 not n20922 ; n20922_not
g70682 not n20931 ; n20931_not
g70683 not n41325 ; n41325_not
g70684 not n20940 ; n20940_not
g70685 not n30381 ; n30381_not
g70686 not n41226 ; n41226_not
g70687 not n20481 ; n20481_not
g70688 not n21570 ; n21570_not
g70689 not n30435 ; n30435_not
g70690 not n53106 ; n53106_not
g70691 not n20472 ; n20472_not
g70692 not n21606 ; n21606_not
g70693 not n53115 ; n53115_not
g70694 not n20463 ; n20463_not
g70695 not n21615 ; n21615_not
g70696 not n21480 ; n21480_not
g70697 not n21624 ; n21624_not
g70698 not n53124 ; n53124_not
g70699 not n21507 ; n21507_not
g70700 not n30426 ; n30426_not
g70701 not n21525 ; n21525_not
g70702 not n41235 ; n41235_not
g70703 not n21534 ; n21534_not
g70704 not n21543 ; n21543_not
g70705 not n21552 ; n21552_not
g70706 not n53331 ; n53331_not
g70707 not n21561 ; n21561_not
g70708 not n20436 ; n20436_not
g70709 not n53142 ; n53142_not
g70710 not n21435 ; n21435_not
g70711 not n41415 ; n41415_not
g70712 not n21705 ; n21705_not
g70713 not n53151 ; n53151_not
g70714 not n21714 ; n21714_not
g70715 not n21723 ; n21723_not
g70716 not n53160 ; n53160_not
g70717 not n20427 ; n20427_not
g70718 not n21732 ; n21732_not
g70719 not n41208 ; n41208_not
g70720 not n21741 ; n21741_not
g70721 not n21750 ; n21750_not
g70722 not n40641 ; n40641_not
g70723 not n20454 ; n20454_not
g70724 not n21633 ; n21633_not
g70725 not n21642 ; n21642_not
g70726 not n21651 ; n21651_not
g70727 not n30273 ; n30273_not
g70728 not n53133 ; n53133_not
g70729 not n21660 ; n21660_not
g70730 not n20445 ; n20445_not
g70731 not n30129 ; n30129_not
g70732 not n53313 ; n53313_not
g70733 not n21453 ; n21453_not
g70734 not n21444 ; n21444_not
g70735 not n30444 ; n30444_not
g70736 not n21327 ; n21327_not
g70737 not n21372 ; n21372_not
g70738 not n41253 ; n41253_not
g70739 not n21282 ; n21282_not
g70740 not n30255 ; n30255_not
g70741 not n20562 ; n20562_not
g70742 not n30417 ; n30417_not
g70743 not n21462 ; n21462_not
g70744 not n20517 ; n20517_not
g70745 not n53340 ; n53340_not
g70746 not n53070 ; n53070_not
g70747 not n21417 ; n21417_not
g70748 not n51315 ; n51315_not
g70749 not n24513 ; n24513_not
g70750 not n31038 ; n31038_not
g70751 not n51324 ; n51324_not
g70752 not n24531 ; n24531_not
g70753 not n24540 ; n24540_not
g70754 not n51333 ; n51333_not
g70755 not n19320 ; n19320_not
g70756 not n30804 ; n30804_not
g70757 not n51342 ; n51342_not
g70758 not n24603 ; n24603_not
g70759 not n31047 ; n31047_not
g70760 not n51351 ; n51351_not
g70761 not n54033 ; n54033_not
g70762 not n29004 ; n29004_not
g70763 not n24423 ; n24423_not
g70764 not n54042 ; n54042_not
g70765 not n51306 ; n51306_not
g70766 not n30822 ; n30822_not
g70767 not n31065 ; n31065_not
g70768 not n24702 ; n24702_not
g70769 not n41811 ; n41811_not
g70770 not n30831 ; n30831_not
g70771 not n31074 ; n31074_not
g70772 not n41820 ; n41820_not
g70773 not n30840 ; n30840_not
g70774 not n31083 ; n31083_not
g70775 not n19311 ; n19311_not
g70776 not n54051 ; n54051_not
g70777 not n24621 ; n24621_not
g70778 not n41802 ; n41802_not
g70779 not n19302 ; n19302_not
g70780 not n24630 ; n24630_not
g70781 not n51360 ; n51360_not
g70782 not n30813 ; n30813_not
g70783 not n31056 ; n31056_not
g70784 not n54060 ; n54060_not
g70785 not n24252 ; n24252_not
g70786 not n29031 ; n29031_not
g70787 not n47310 ; n47310_not
g70788 not n24261 ; n24261_not
g70789 not n24270 ; n24270_not
g70790 not n19212 ; n19212_not
g70791 not n19221 ; n19221_not
g70792 not n51027 ; n51027_not
g70793 not n24225 ; n24225_not
g70794 not n24234 ; n24234_not
g70795 not n53304 ; n53304_not
g70796 not n51270 ; n51270_not
g70797 not n41271 ; n41271_not
g70798 not n41730 ; n41730_not
g70799 not n24243 ; n24243_not
g70800 not n19203 ; n19203_not
g70801 not n24333 ; n24333_not
g70802 not n40632 ; n40632_not
g70803 not n24342 ; n24342_not
g70804 not n24351 ; n24351_not
g70805 not n54024 ; n54024_not
g70806 not n24360 ; n24360_not
g70807 not n29022 ; n29022_not
g70808 not n23622 ; n23622_not
g70809 not n23613 ; n23613_not
g70810 not n29013 ; n29013_not
g70811 not n54006 ; n54006_not
g70812 not n50127 ; n50127_not
g70813 not n29040 ; n29040_not
g70814 not n50136 ; n50136_not
g70815 not n24306 ; n24306_not
g70816 not n19410 ; n19410_not
g70817 not n24315 ; n24315_not
g70818 not n54015 ; n54015_not
g70819 not n19401 ; n19401_not
g70820 not n24324 ; n24324_not
g70821 not n19041 ; n19041_not
g70822 not n19050 ; n19050_not
g70823 not n31137 ; n31137_not
g70824 not n31128 ; n31128_not
g70825 not n19032 ; n19032_not
g70826 not n31119 ; n31119_not
g70827 not n31191 ; n31191_not
g70828 not n19023 ; n19023_not
g70829 not n19014 ; n19014_not
g70830 not n54150 ; n54150_not
g70831 not n40173 ; n40173_not
g70832 not n31146 ; n31146_not
g70833 not n41910 ; n41910_not
g70834 not n54213 ; n54213_not
g70835 not n51513 ; n51513_not
g70836 not n31236 ; n31236_not
g70837 not n24504 ; n24504_not
g70838 not n19005 ; n19005_not
g70839 not n31092 ; n31092_not
g70840 not n51504 ; n51504_not
g70841 not n51414 ; n51414_not
g70842 not n52701 ; n52701_not
g70843 not n54105 ; n54105_not
g70844 not n51423 ; n51423_not
g70845 not n30903 ; n30903_not
g70846 not n19230 ; n19230_not
g70847 not n51405 ; n51405_not
g70848 not n40128 ; n40128_not
g70849 not n19122 ; n19122_not
g70850 not n51450 ; n51450_not
g70851 not n19113 ; n19113_not
g70852 not n30912 ; n30912_not
g70853 not n54141 ; n54141_not
g70854 not n52710 ; n52710_not
g70855 not n51432 ; n51432_not
g70856 not n28014 ; n28014_not
g70857 not n19140 ; n19140_not
g70858 not n51441 ; n51441_not
g70859 not n54123 ; n54123_not
g70860 not n53700 ; n53700_not
g70861 not n45420 ; n45420_not
g70862 not n23721 ; n23721_not
g70863 not n30624 ; n30624_not
g70864 not n40326 ; n40326_not
g70865 not n45105 ; n45105_not
g70866 not n29211 ; n29211_not
g70867 not n29220 ; n29220_not
g70868 not n40821 ; n40821_not
g70869 not n41550 ; n41550_not
g70870 not n19500 ; n19500_not
g70871 not n40317 ; n40317_not
g70872 not n30633 ; n30633_not
g70873 not n51234 ; n51234_not
g70874 not n45510 ; n45510_not
g70875 not n30642 ; n30642_not
g70876 not n41523 ; n41523_not
g70877 not n40911 ; n40911_not
g70878 not n51216 ; n51216_not
g70879 not n40344 ; n40344_not
g70880 not n30516 ; n30516_not
g70881 not n30606 ; n30606_not
g70882 not n41532 ; n41532_not
g70883 not n40902 ; n40902_not
g70884 not n40812 ; n40812_not
g70885 not n40335 ; n40335_not
g70886 not n30615 ; n30615_not
g70887 not n51225 ; n51225_not
g70888 not n41541 ; n41541_not
g70889 not n23703 ; n23703_not
g70890 not n40290 ; n40290_not
g70891 not n29202 ; n29202_not
g70892 not n41604 ; n41604_not
g70893 not n30723 ; n30723_not
g70894 not n30732 ; n30732_not
g70895 not n41613 ; n41613_not
g70896 not n51252 ; n51252_not
g70897 not n23901 ; n23901_not
g70898 not n23910 ; n23910_not
g70899 not n30750 ; n30750_not
g70900 not n29112 ; n29112_not
g70901 not n30651 ; n30651_not
g70902 not n30660 ; n30660_not
g70903 not n40830 ; n40830_not
g70904 not n41361 ; n41361_not
g70905 not n40308 ; n40308_not
g70906 not n38121 ; n38121_not
g70907 not n23811 ; n23811_not
g70908 not n45411 ; n45411_not
g70909 not n30705 ; n30705_not
g70910 not n51243 ; n51243_not
g70911 not n50361 ; n50361_not
g70912 not n50352 ; n50352_not
g70913 not n30561 ; n30561_not
g70914 not n50343 ; n50343_not
g70915 not n40434 ; n40434_not
g70916 not n51108 ; n51108_not
g70917 not n40425 ; n40425_not
g70918 not n47112 ; n47112_not
g70919 not n51117 ; n51117_not
g70920 not n40416 ; n40416_not
g70921 not n47103 ; n47103_not
g70922 not n51126 ; n51126_not
g70923 not n50415 ; n50415_not
g70924 not n30552 ; n30552_not
g70925 not n23109 ; n23109_not
g70926 not n51063 ; n51063_not
g70927 not n50406 ; n50406_not
g70928 not n47130 ; n47130_not
g70929 not n51081 ; n51081_not
g70930 not n23037 ; n23037_not
g70931 not n38004 ; n38004_not
g70932 not n50370 ; n50370_not
g70933 not n40362 ; n40362_not
g70934 not n51207 ; n51207_not
g70935 not n22812 ; n22812_not
g70936 not n40920 ; n40920_not
g70937 not n41505 ; n41505_not
g70938 not n23604 ; n23604_not
g70939 not n30570 ; n30570_not
g70940 not n40353 ; n40353_not
g70941 not n41514 ; n41514_not
g70942 not n45501 ; n45501_not
g70943 not n23631 ; n23631_not
g70944 not n38400 ; n38400_not
g70945 not n51135 ; n51135_not
g70946 not n40407 ; n40407_not
g70947 not n51144 ; n51144_not
g70948 not n22902 ; n22902_not
g70949 not n51153 ; n51153_not
g70950 not n51162 ; n51162_not
g70951 not n40380 ; n40380_not
g70952 not n51171 ; n51171_not
g70953 not n40371 ; n40371_not
g70954 not n52521 ; n52521_not
g70955 not n51180 ; n51180_not
g70956 not n51072 ; n51072_not
g70957 not n24108 ; n24108_not
g70958 not n24117 ; n24117_not
g70959 not n51261 ; n51261_not
g70960 not n29103 ; n29103_not
g70961 not n24126 ; n24126_not
g70962 not n24135 ; n24135_not
g70963 not n24144 ; n24144_not
g70964 not n24072 ; n24072_not
g70965 not n24081 ; n24081_not
g70966 not n19131 ; n19131_not
g70967 not n24090 ; n24090_not
g70968 not n24207 ; n24207_not
g70969 not n30921 ; n30921_not
g70970 not n23712 ; n23712_not
g70971 not n24216 ; n24216_not
g70972 not n41721 ; n41721_not
g70973 not n50118 ; n50118_not
g70974 not n41703 ; n41703_not
g70975 not n24153 ; n24153_not
g70976 not n24162 ; n24162_not
g70977 not n38103 ; n38103_not
g70978 not n52611 ; n52611_not
g70979 not n24171 ; n24171_not
g70980 not n24180 ; n24180_not
g70981 not n41712 ; n41712_not
g70982 not n40704 ; n40704_not
g70983 not n46401 ; n46401_not
g70984 not n41640 ; n41640_not
g70985 not n41622 ; n41622_not
g70986 not n38130 ; n38130_not
g70987 not n41631 ; n41631_not
g70988 not n24036 ; n24036_not
g70989 not n24045 ; n24045_not
g70990 not n23802 ; n23802_not
g70991 not n24054 ; n24054_not
g70992 not n24063 ; n24063_not
g70993 not n30741 ; n30741_not
g70994 not n24009 ; n24009_not
g70995 not n41316 ; n41316_not
g70996 not n24018 ; n24018_not
g70997 not n45402 ; n45402_not
g70998 not n24027 ; n24027_not
g70999 not n55014 ; n55014_not
g71000 not n43080 ; n43080_not
g71001 not n32109 ; n32109_not
g71002 not n17043 ; n17043_not
g71003 not n34143 ; n34143_not
g71004 not n13722 ; n13722_not
g71005 not n13353 ; n13353_not
g71006 not n14442 ; n14442_not
g71007 not n35142 ; n35142_not
g71008 not n16521 ; n16521_not
g71009 not n14802 ; n14802_not
g71010 not n13146 ; n13146_not
g71011 not n10905 ; n10905_not
g71012 not n55023 ; n55023_not
g71013 not n33621 ; n33621_not
g71014 not n14811 ; n14811_not
g71015 not n10914 ; n10914_not
g71016 not n10923 ; n10923_not
g71017 not n35151 ; n35151_not
g71018 not n11472 ; n11472_not
g71019 not n34800 ; n34800_not
g71020 not n11463 ; n11463_not
g71021 not n45024 ; n45024_not
g71022 not n35115 ; n35115_not
g71023 not n11445 ; n11445_not
g71024 not n11427 ; n11427_not
g71025 not n17430 ; n17430_not
g71026 not n11418 ; n11418_not
g71027 not n13740 ; n13740_not
g71028 not n32118 ; n32118_not
g71029 not n14460 ; n14460_not
g71030 not n17052 ; n17052_not
g71031 not n35124 ; n35124_not
g71032 not n43071 ; n43071_not
g71033 not n14451 ; n14451_not
g71034 not n35133 ; n35133_not
g71035 not n42630 ; n42630_not
g71036 not n43611 ; n43611_not
g71037 not n37014 ; n37014_not
g71038 not n43602 ; n43602_not
g71039 not n12633 ; n12633_not
g71040 not n14901 ; n14901_not
g71041 not n14910 ; n14910_not
g71042 not n50028 ; n50028_not
g71043 not n32091 ; n32091_not
g71044 not n42504 ; n42504_not
g71045 not n13173 ; n13173_not
g71046 not n42621 ; n42621_not
g71047 not n42450 ; n42450_not
g71048 not n37005 ; n37005_not
g71049 not n12624 ; n12624_not
g71050 not n56022 ; n56022_not
g71051 not n34503 ; n34503_not
g71052 not n14820 ; n14820_not
g71053 not n35160 ; n35160_not
g71054 not n17034 ; n17034_not
g71055 not n55212 ; n55212_not
g71056 not n50037 ; n50037_not
g71057 not n14415 ; n14415_not
g71058 not n10950 ; n10950_not
g71059 not n55140 ; n55140_not
g71060 not n43620 ; n43620_not
g71061 not n13128 ; n13128_not
g71062 not n14406 ; n14406_not
g71063 not n12642 ; n12642_not
g71064 not n13119 ; n13119_not
g71065 not n33270 ; n33270_not
g71066 not n14622 ; n14622_not
g71067 not n11571 ; n11571_not
g71068 not n56211 ; n56211_not
g71069 not n13821 ; n13821_not
g71070 not n35043 ; n35043_not
g71071 not n48021 ; n48021_not
g71072 not n32145 ; n32145_not
g71073 not n55005 ; n55005_not
g71074 not n44115 ; n44115_not
g71075 not n13812 ; n13812_not
g71076 not n14631 ; n14631_not
g71077 not n43701 ; n43701_not
g71078 not n14532 ; n14532_not
g71079 not n35052 ; n35052_not
g71080 not n33711 ; n33711_not
g71081 not n14640 ; n14640_not
g71082 not n50019 ; n50019_not
g71083 not n56040 ; n56040_not
g71084 not n34530 ; n34530_not
g71085 not n44250 ; n44250_not
g71086 not n44124 ; n44124_not
g71087 not n34125 ; n34125_not
g71088 not n56202 ; n56202_not
g71089 not n36510 ; n36510_not
g71090 not n32154 ; n32154_not
g71091 not n14604 ; n14604_not
g71092 not n35025 ; n35025_not
g71093 not n32046 ; n32046_not
g71094 not n16080 ; n16080_not
g71095 not n34134 ; n34134_not
g71096 not n11553 ; n11553_not
g71097 not n35034 ; n35034_not
g71098 not n14550 ; n14550_not
g71099 not n14613 ; n14613_not
g71100 not n14541 ; n14541_not
g71101 not n17016 ; n17016_not
g71102 not n11562 ; n11562_not
g71103 not n34107 ; n34107_not
g71104 not n17412 ; n17412_not
g71105 not n14712 ; n14712_not
g71106 not n43062 ; n43062_not
g71107 not n14721 ; n14721_not
g71108 not n32127 ; n32127_not
g71109 not n11535 ; n11535_not
g71110 not n11517 ; n11517_not
g71111 not n11508 ; n11508_not
g71112 not n11490 ; n11490_not
g71113 not n35106 ; n35106_not
g71114 not n14730 ; n14730_not
g71115 not n32064 ; n32064_not
g71116 not n17421 ; n17421_not
g71117 not n44106 ; n44106_not
g71118 not n34521 ; n34521_not
g71119 not n35061 ; n35061_not
g71120 not n32136 ; n32136_not
g71121 not n33702 ; n33702_not
g71122 not n56220 ; n56220_not
g71123 not n34116 ; n34116_not
g71124 not n35070 ; n35070_not
g71125 not n55122 ; n55122_not
g71126 not n17403 ; n17403_not
g71127 not n44610 ; n44610_not
g71128 not n14505 ; n14505_not
g71129 not n50307 ; n50307_not
g71130 not n11634 ; n11634_not
g71131 not n11616 ; n11616_not
g71132 not n11625 ; n11625_not
g71133 not n14703 ; n14703_not
g71134 not n11607 ; n11607_not
g71135 not n32055 ; n32055_not
g71136 not n32370 ; n32370_not
g71137 not n11580 ; n11580_not
g71138 not n34431 ; n34431_not
g71139 not n15225 ; n15225_not
g71140 not n33414 ; n33414_not
g71141 not n13029 ; n13029_not
g71142 not n44313 ; n44313_not
g71143 not n15234 ; n15234_not
g71144 not n16260 ; n16260_not
g71145 not n16512 ; n16512_not
g71146 not n33405 ; n33405_not
g71147 not n43512 ; n43512_not
g71148 not n15243 ; n15243_not
g71149 not n34053 ; n34053_not
g71150 not n15180 ; n15180_not
g71151 not n15252 ; n15252_not
g71152 not n13218 ; n13218_not
g71153 not n10932 ; n10932_not
g71154 not n33450 ; n33450_not
g71155 not n13047 ; n13047_not
g71156 not n15162 ; n15162_not
g71157 not n33441 ; n33441_not
g71158 not n34440 ; n34440_not
g71159 not n16503 ; n16503_not
g71160 not n33432 ; n33432_not
g71161 not n16116 ; n16116_not
g71162 not n33360 ; n33360_not
g71163 not n33423 ; n33423_not
g71164 not n13038 ; n13038_not
g71165 not n43521 ; n43521_not
g71166 not n15207 ; n15207_not
g71167 not n15216 ; n15216_not
g71168 not n33072 ; n33072_not
g71169 not n16251 ; n16251_not
g71170 not n33081 ; n33081_not
g71171 not n15153 ; n15153_not
g71172 not n15306 ; n15306_not
g71173 not n55401 ; n55401_not
g71174 not n12552 ; n12552_not
g71175 not n35331 ; n35331_not
g71176 not n15144 ; n15144_not
g71177 not n16125 ; n16125_not
g71178 not n33090 ; n33090_not
g71179 not n35340 ; n35340_not
g71180 not n15315 ; n15315_not
g71181 not n15324 ; n15324_not
g71182 not n42441 ; n42441_not
g71183 not n13137 ; n13137_not
g71184 not n15261 ; n15261_not
g71185 not n50055 ; n50055_not
g71186 not n15270 ; n15270_not
g71187 not n33054 ; n33054_not
g71188 not n43503 ; n43503_not
g71189 not n13227 ; n13227_not
g71190 not n12534 ; n12534_not
g71191 not n35313 ; n35313_not
g71192 not n33063 ; n33063_not
g71193 not n43152 ; n43152_not
g71194 not n50208 ; n50208_not
g71195 not n35322 ; n35322_not
g71196 not n33531 ; n33531_not
g71197 not n13182 ; n13182_not
g71198 not n15009 ; n15009_not
g71199 not n33522 ; n33522_not
g71200 not n17502 ; n17502_not
g71201 not n13083 ; n13083_not
g71202 not n13191 ; n13191_not
g71203 not n15027 ; n15027_not
g71204 not n33513 ; n33513_not
g71205 not n13074 ; n13074_not
g71206 not n17511 ; n17511_not
g71207 not n56013 ; n56013_not
g71208 not n33315 ; n33315_not
g71209 not n16107 ; n16107_not
g71210 not n15900 ; n15900_not
g71211 not n13092 ; n13092_not
g71212 not n14370 ; n14370_not
g71213 not n14361 ; n14361_not
g71214 not n43107 ; n43107_not
g71215 not n48003 ; n48003_not
g71216 not n14352 ; n14352_not
g71217 not n35205 ; n35205_not
g71218 not n56031 ; n56031_not
g71219 not n55050 ; n55050_not
g71220 not n34071 ; n34071_not
g71221 not n43116 ; n43116_not
g71222 not n33540 ; n33540_not
g71223 not n43125 ; n43125_not
g71224 not n35232 ; n35232_not
g71225 not n42603 ; n42603_not
g71226 not n33333 ; n33333_not
g71227 not n15090 ; n15090_not
g71228 not n55410 ; n55410_not
g71229 not n43530 ; n43530_not
g71230 not n44304 ; n44304_not
g71231 not n13056 ; n13056_not
g71232 not n15117 ; n15117_not
g71233 not n42540 ; n42540_not
g71234 not n16530 ; n16530_not
g71235 not n32073 ; n32073_not
g71236 not n45240 ; n45240_not
g71237 not n15135 ; n15135_not
g71238 not n35250 ; n35250_not
g71239 not n11085 ; n11085_not
g71240 not n15045 ; n15045_not
g71241 not n32604 ; n32604_not
g71242 not n15054 ; n15054_not
g71243 not n17007 ; n17007_not
g71244 not n11076 ; n11076_not
g71245 not n11049 ; n11049_not
g71246 not n17520 ; n17520_not
g71247 not n33504 ; n33504_not
g71248 not n34062 ; n34062_not
g71249 not n11058 ; n11058_not
g71250 not n50316 ; n50316_not
g71251 not n32325 ; n32325_not
g71252 not n15072 ; n15072_not
g71253 not n35223 ; n35223_not
g71254 not n13065 ; n13065_not
g71255 not n33324 ; n33324_not
g71256 not n14028 ; n14028_not
g71257 not n12183 ; n12183_not
g71258 not n32244 ; n32244_not
g71259 not n14019 ; n14019_not
g71260 not n12417 ; n12417_not
g71261 not n50226 ; n50226_not
g71262 not n12354 ; n12354_not
g71263 not n14208 ; n14208_not
g71264 not n16053 ; n16053_not
g71265 not n12345 ; n12345_not
g71266 not n12408 ; n12408_not
g71267 not n12336 ; n12336_not
g71268 not n12093 ; n12093_not
g71269 not n16404 ; n16404_not
g71270 not n14217 ; n14217_not
g71271 not n12327 ; n12327_not
g71272 not n13902 ; n13902_not
g71273 not n16017 ; n16017_not
g71274 not n12057 ; n12057_not
g71275 not n14181 ; n14181_not
g71276 not n12390 ; n12390_not
g71277 not n12066 ; n12066_not
g71278 not n12444 ; n12444_not
g71279 not n12381 ; n12381_not
g71280 not n14190 ; n14190_not
g71281 not n12606 ; n12606_not
g71282 not n12435 ; n12435_not
g71283 not n12426 ; n12426_not
g71284 not n12372 ; n12372_not
g71285 not n32307 ; n32307_not
g71286 not n12363 ; n12363_not
g71287 not n37113 ; n37113_not
g71288 not n14235 ; n14235_not
g71289 not n12651 ; n12651_not
g71290 not n17223 ; n17223_not
g71291 not n12282 ; n12282_not
g71292 not n16701 ; n16701_not
g71293 not n12273 ; n12273_not
g71294 not n14244 ; n14244_not
g71295 not n44151 ; n44151_not
g71296 not n34017 ; n34017_not
g71297 not n12264 ; n12264_not
g71298 not n33900 ; n33900_not
g71299 not n17232 ; n17232_not
g71300 not n32226 ; n32226_not
g71301 not n56130 ; n56130_not
g71302 not n45231 ; n45231_not
g71303 not n17205 ; n17205_not
g71304 not n56121 ; n56121_not
g71305 not n13911 ; n13911_not
g71306 not n12318 ; n12318_not
g71307 not n32235 ; n32235_not
g71308 not n13920 ; n13920_not
g71309 not n12309 ; n12309_not
g71310 not n17106 ; n17106_not
g71311 not n17214 ; n17214_not
g71312 not n16008 ; n16008_not
g71313 not n14226 ; n14226_not
g71314 not n34008 ; n34008_not
g71315 not n12291 ; n12291_not
g71316 not n34404 ; n34404_not
g71317 not n12516 ; n12516_not
g71318 not n12507 ; n12507_not
g71319 not n14109 ; n14109_not
g71320 not n34710 ; n34710_not
g71321 not n16044 ; n16044_not
g71322 not n14118 ; n14118_not
g71323 not n16035 ; n16035_not
g71324 not n17133 ; n17133_not
g71325 not n37140 ; n37140_not
g71326 not n14127 ; n14127_not
g71327 not n12480 ; n12480_not
g71328 not n44160 ; n44160_not
g71329 not n14136 ; n14136_not
g71330 not n16413 ; n16413_not
g71331 not n16620 ; n16620_not
g71332 not n14073 ; n14073_not
g71333 not n12525 ; n12525_not
g71334 not n16611 ; n16611_not
g71335 not n34701 ; n34701_not
g71336 not n14082 ; n14082_not
g71337 not n12561 ; n12561_not
g71338 not n14064 ; n14064_not
g71339 not n50145 ; n50145_not
g71340 not n14091 ; n14091_not
g71341 not n16602 ; n16602_not
g71342 not n17151 ; n17151_not
g71343 not n37050 ; n37050_not
g71344 not n37131 ; n37131_not
g71345 not n12471 ; n12471_not
g71346 not n55230 ; n55230_not
g71347 not n12462 ; n12462_not
g71348 not n12048 ; n12048_not
g71349 not n14037 ; n14037_not
g71350 not n13830 ; n13830_not
g71351 not n32253 ; n32253_not
g71352 not n56103 ; n56103_not
g71353 not n14172 ; n14172_not
g71354 not n12453 ; n12453_not
g71355 not n14145 ; n14145_not
g71356 not n14055 ; n14055_not
g71357 not n33630 ; n33630_not
g71358 not n14046 ; n14046_not
g71359 not n16026 ; n16026_not
g71360 not n14154 ; n14154_not
g71361 not n17124 ; n17124_not
g71362 not n32262 ; n32262_not
g71363 not n14163 ; n14163_not
g71364 not n48012 ; n48012_not
g71365 not n32181 ; n32181_not
g71366 not n44214 ; n44214_not
g71367 not n44601 ; n44601_not
g71368 not n44133 ; n44133_not
g71369 not n32352 ; n32352_not
g71370 not n17322 ; n17322_not
g71371 not n55032 ; n55032_not
g71372 not n37041 ; n37041_not
g71373 not n11436 ; n11436_not
g71374 not n33810 ; n33810_not
g71375 not n55320 ; n55320_not
g71376 not n16071 ; n16071_not
g71377 not n34611 ; n34611_not
g71378 not n34080 ; n34080_not
g71379 not n44142 ; n44142_not
g71380 not n32190 ; n32190_not
g71381 not n55104 ; n55104_not
g71382 not n50253 ; n50253_not
g71383 not n14424 ; n14424_not
g71384 not n17304 ; n17304_not
g71385 not n44205 ; n44205_not
g71386 not n55311 ; n55311_not
g71387 not n34620 ; n34620_not
g71388 not n50217 ; n50217_not
g71389 not n55302 ; n55302_not
g71390 not n17313 ; n17313_not
g71391 not n12732 ; n12732_not
g71392 not n44232 ; n44232_not
g71393 not n12723 ; n12723_not
g71394 not n50280 ; n50280_not
g71395 not n44241 ; n44241_not
g71396 not n32163 ; n32163_not
g71397 not n12714 ; n12714_not
g71398 not n35007 ; n35007_not
g71399 not n11526 ; n11526_not
g71400 not n35016 ; n35016_not
g71401 not n33801 ; n33801_not
g71402 not n17331 ; n17331_not
g71403 not n50262 ; n50262_not
g71404 not n16800 ; n16800_not
g71405 not n33720 ; n33720_not
g71406 not n32172 ; n32172_not
g71407 not n44223 ; n44223_not
g71408 not n14514 ; n14514_not
g71409 not n37023 ; n37023_not
g71410 not n17340 ; n17340_not
g71411 not n34602 ; n34602_not
g71412 not n11481 ; n11481_not
g71413 not n12219 ; n12219_not
g71414 not n32217 ; n32217_not
g71415 not n14271 ; n14271_not
g71416 not n34035 ; n34035_not
g71417 not n14280 ; n14280_not
g71418 not n12192 ; n12192_not
g71419 not n16710 ; n16710_not
g71420 not n12255 ; n12255_not
g71421 not n12138 ; n12138_not
g71422 not n17241 ; n17241_not
g71423 not n14253 ; n14253_not
g71424 not n50190 ; n50190_not
g71425 not n12246 ; n12246_not
g71426 not n12237 ; n12237_not
g71427 not n14262 ; n14262_not
g71428 not n12147 ; n12147_not
g71429 not n12228 ; n12228_not
g71430 not n12156 ; n12156_not
g71431 not n17250 ; n17250_not
g71432 not n12741 ; n12741_not
g71433 not n14334 ; n14334_not
g71434 not n50235 ; n50235_not
g71435 not n14343 ; n14343_not
g71436 not n12075 ; n12075_not
g71437 not n12750 ; n12750_not
g71438 not n17061 ; n17061_not
g71439 not n16062 ; n16062_not
g71440 not n32334 ; n32334_not
g71441 not n14307 ; n14307_not
g71442 not n12165 ; n12165_not
g71443 not n16440 ; n16440_not
g71444 not n32208 ; n32208_not
g71445 not n14316 ; n14316_not
g71446 not n32019 ; n32019_not
g71447 not n17142 ; n17142_not
g71448 not n14325 ; n14325_not
g71449 not n16134 ; n16134_not
g71450 not n44007 ; n44007_not
g71451 not n33045 ; n33045_not
g71452 not n13290 ; n13290_not
g71453 not n16143 ; n16143_not
g71454 not n16350 ; n16350_not
g71455 not n31920 ; n31920_not
g71456 not n43341 ; n43341_not
g71457 not n44052 ; n44052_not
g71458 not n43242 ; n43242_not
g71459 not n15801 ; n15801_not
g71460 not n32730 ; n32730_not
g71461 not n16152 ; n16152_not
g71462 not n12921 ; n12921_not
g71463 not n12912 ; n12912_not
g71464 not n35700 ; n35700_not
g71465 not n12903 ; n12903_not
g71466 not n33018 ; n33018_not
g71467 not n43350 ; n43350_not
g71468 not n33027 ; n33027_not
g71469 not n12831 ; n12831_not
g71470 not n31911 ; n31911_not
g71471 not n12822 ; n12822_not
g71472 not n16332 ; n16332_not
g71473 not n33009 ; n33009_not
g71474 not n36213 ; n36213_not
g71475 not n13281 ; n13281_not
g71476 not n43323 ; n43323_not
g71477 not n43251 ; n43251_not
g71478 not n37104 ; n37104_not
g71479 not n12813 ; n12813_not
g71480 not n43314 ; n43314_not
g71481 not n43260 ; n43260_not
g71482 not n32802 ; n32802_not
g71483 not n16206 ; n16206_not
g71484 not n13308 ; n13308_not
g71485 not n49200 ; n49200_not
g71486 not n12840 ; n12840_not
g71487 not n36501 ; n36501_not
g71488 not n13317 ; n13317_not
g71489 not n16161 ; n16161_not
g71490 not n43332 ; n43332_not
g71491 not n16170 ; n16170_not
g71492 not n34026 ; n34026_not
g71493 not n36042 ; n36042_not
g71494 not n33036 ; n33036_not
g71495 not n55500 ; n55500_not
g71496 not n35241 ; n35241_not
g71497 not n10059 ; n10059_not
g71498 not n13263 ; n13263_not
g71499 not n33171 ; n33171_not
g71500 not n12930 ; n12930_not
g71501 not n45204 ; n45204_not
g71502 not n33162 ; n33162_not
g71503 not n56400 ; n56400_not
g71504 not n44403 ; n44403_not
g71505 not n43215 ; n43215_not
g71506 not n10248 ; n10248_not
g71507 not n10239 ; n10239_not
g71508 not n10194 ; n10194_not
g71509 not n10185 ; n10185_not
g71510 not n33180 ; n33180_not
g71511 not n10176 ; n10176_not
g71512 not n10167 ; n10167_not
g71513 not n16422 ; n16422_not
g71514 not n10158 ; n10158_not
g71515 not n10149 ; n10149_not
g71516 not n44412 ; n44412_not
g71517 not n10095 ; n10095_not
g71518 not n43206 ; n43206_not
g71519 not n10086 ; n10086_not
g71520 not n10077 ; n10077_not
g71521 not n10068 ; n10068_not
g71522 not n13272 ; n13272_not
g71523 not n33117 ; n33117_not
g71524 not n15702 ; n15702_not
g71525 not n43053 ; n43053_not
g71526 not n15711 ; n15711_not
g71527 not n33108 ; n33108_not
g71528 not n36222 ; n36222_not
g71529 not n36231 ; n36231_not
g71530 not n44511 ; n44511_not
g71531 not n16323 ; n16323_not
g71532 not n44421 ; n44421_not
g71533 not n33153 ; n33153_not
g71534 not n33144 ; n33144_not
g71535 not n35610 ; n35610_not
g71536 not n33135 ; n33135_not
g71537 not n32820 ; n32820_not
g71538 not n33126 ; n33126_not
g71539 not n32811 ; n32811_not
g71540 not n44016 ; n44016_not
g71541 not n32613 ; n32613_not
g71542 not n32721 ; n32721_not
g71543 not n57300 ; n57300_not
g71544 not n36114 ; n36114_not
g71545 not n36123 ; n36123_not
g71546 not n13326 ; n13326_not
g71547 not n36141 ; n36141_not
g71548 not n57210 ; n57210_not
g71549 not n36051 ; n36051_not
g71550 not n43224 ; n43224_not
g71551 not n15630 ; n15630_not
g71552 not n50271 ; n50271_not
g71553 not n36132 ; n36132_not
g71554 not n32703 ; n32703_not
g71555 not n44034 ; n44034_not
g71556 not n44502 ; n44502_not
g71557 not n43134 ; n43134_not
g71558 not n44025 ; n44025_not
g71559 not n47121 ; n47121_not
g71560 not n42405 ; n42405_not
g71561 not n15720 ; n15720_not
g71562 not n43161 ; n43161_not
g71563 not n32640 ; n32640_not
g71564 not n32343 ; n32343_not
g71565 not n45114 ; n45114_not
g71566 not n36204 ; n36204_not
g71567 not n13335 ; n13335_not
g71568 not n16242 ; n16242_not
g71569 not n12804 ; n12804_not
g71570 not n44043 ; n44043_not
g71571 not n31902 ; n31902_not
g71572 not n16314 ; n16314_not
g71573 not n49110 ; n49110_not
g71574 not n16215 ; n16215_not
g71575 not n57012 ; n57012_not
g71576 not n16224 ; n16224_not
g71577 not n16305 ; n16305_not
g71578 not n49101 ; n49101_not
g71579 not n57030 ; n57030_not
g71580 not n43305 ; n43305_not
g71581 not n31722 ; n31722_not
g71582 not n16233 ; n16233_not
g71583 not n49002 ; n49002_not
g71584 not n36006 ; n36006_not
g71585 not n36015 ; n36015_not
g71586 not n36024 ; n36024_not
g71587 not n32712 ; n32712_not
g71588 not n57201 ; n57201_not
g71589 not n42414 ; n42414_not
g71590 not n36033 ; n36033_not
g71591 not n55203 ; n55203_not
g71592 not n42423 ; n42423_not
g71593 not n57102 ; n57102_not
g71594 not n49020 ; n49020_not
g71595 not n32901 ; n32901_not
g71596 not n32910 ; n32910_not
g71597 not n49011 ; n49011_not
g71598 not n15810 ; n15810_not
g71599 not n15441 ; n15441_not
g71600 not n10437 ; n10437_not
g71601 not n33234 ; n33234_not
g71602 not n10527 ; n10527_not
g71603 not n10671 ; n10671_not
g71604 not n33243 ; n33243_not
g71605 not n15450 ; n15450_not
g71606 not n10662 ; n10662_not
g71607 not n10446 ; n10446_not
g71608 not n33252 ; n33252_not
g71609 not n10653 ; n10653_not
g71610 not n10455 ; n10455_not
g71611 not n33261 ; n33261_not
g71612 not n33207 ; n33207_not
g71613 not n15423 ; n15423_not
g71614 not n10725 ; n10725_not
g71615 not n42531 ; n42531_not
g71616 not n10716 ; n10716_not
g71617 not n33216 ; n33216_not
g71618 not n15432 ; n15432_not
g71619 not n10707 ; n10707_not
g71620 not n33225 ; n33225_not
g71621 not n10680 ; n10680_not
g71622 not n43440 ; n43440_not
g71623 not n10608 ; n10608_not
g71624 not n10482 ; n10482_not
g71625 not n10590 ; n10590_not
g71626 not n43431 ; n43431_not
g71627 not n15504 ; n15504_not
g71628 not n42513 ; n42513_not
g71629 not n10644 ; n10644_not
g71630 not n55113 ; n55113_not
g71631 not n10635 ; n10635_not
g71632 not n15063 ; n15063_not
g71633 not n10626 ; n10626_not
g71634 not n56301 ; n56301_not
g71635 not n10617 ; n10617_not
g71636 not n10824 ; n10824_not
g71637 not n10356 ; n10356_not
g71638 not n33342 ; n33342_not
g71639 not n10815 ; n10815_not
g71640 not n10365 ; n10365_not
g71641 not n17601 ; n17601_not
g71642 not n15351 ; n15351_not
g71643 not n13155 ; n13155_not
g71644 not n10806 ; n10806_not
g71645 not n15360 ; n15360_not
g71646 not n54114 ; n54114_not
g71647 not n13236 ; n13236_not
g71648 not n10860 ; n10860_not
g71649 not n15333 ; n15333_not
g71650 not n32622 ; n32622_not
g71651 not n10842 ; n10842_not
g71652 not n10347 ; n10347_not
g71653 not n15342 ; n15342_not
g71654 not n10833 ; n10833_not
g71655 not n44322 ; n44322_not
g71656 not n10761 ; n10761_not
g71657 not n44331 ; n44331_not
g71658 not n10392 ; n10392_not
g71659 not n17610 ; n17610_not
g71660 not n34413 ; n34413_not
g71661 not n10752 ; n10752_not
g71662 not n15405 ; n15405_not
g71663 not n10743 ; n10743_not
g71664 not n15414 ; n15414_not
g71665 not n10734 ; n10734_not
g71666 not n32028 ; n32028_not
g71667 not n10770 ; n10770_not
g71668 not n43170 ; n43170_not
g71669 not n15108 ; n15108_not
g71670 not n15018 ; n15018_not
g71671 not n10419 ; n10419_not
g71672 not n44070 ; n44070_not
g71673 not n15531 ; n15531_not
g71674 not n10491 ; n10491_not
g71675 not n47211 ; n47211_not
g71676 not n15540 ; n15540_not
g71677 not n10464 ; n10464_not
g71678 not n10338 ; n10338_not
g71679 not n43413 ; n43413_not
g71680 not n10293 ; n10293_not
g71681 not n44061 ; n44061_not
g71682 not n10284 ; n10284_not
g71683 not n43404 ; n43404_not
g71684 not n10275 ; n10275_not
g71685 not n10266 ; n10266_not
g71686 not n15603 ; n15603_not
g71687 not n10257 ; n10257_not
g71688 not n13245 ; n13245_not
g71689 not n10374 ; n10374_not
g71690 not n43422 ; n43422_not
g71691 not n15522 ; n15522_not
g71692 not n10545 ; n10545_not
g71693 not n10554 ; n10554_not
g71694 not n10563 ; n10563_not
g71695 not n56310 ; n56310_not
g71696 not n15513 ; n15513_not
g71697 not n10572 ; n10572_not
g71698 not n10581 ; n10581_not
g71699 not n10509 ; n10509_not
g71700 not n10536 ; n10536_not
g71701 not n34108 ; n34108_not
g71702 not n50047 ; n50047_not
g71703 not n34117 ; n34117_not
g71704 not n41119 ; n41119_not
g71705 not n41083 ; n41083_not
g71706 not n44017 ; n44017_not
g71707 not n13543 ; n13543_not
g71708 not n22237 ; n22237_not
g71709 not n14047 ; n14047_not
g71710 not n13552 ; n13552_not
g71711 not n34018 ; n34018_not
g71712 not n34234 ; n34234_not
g71713 not n13651 ; n13651_not
g71714 not n13570 ; n13570_not
g71715 not n13561 ; n13561_not
g71716 not n50083 ; n50083_not
g71717 not n22174 ; n22174_not
g71718 not n13642 ; n13642_not
g71719 not n34216 ; n34216_not
g71720 not n13228 ; n13228_not
g71721 not n22255 ; n22255_not
g71722 not n13156 ; n13156_not
g71723 not n34027 ; n34027_not
g71724 not n50056 ; n50056_not
g71725 not n41056 ; n41056_not
g71726 not n13237 ; n13237_not
g71727 not n13516 ; n13516_not
g71728 not n22246 ; n22246_not
g71729 not n13660 ; n13660_not
g71730 not n22813 ; n22813_not
g71731 not n13453 ; n13453_not
g71732 not n13525 ; n13525_not
g71733 not n22192 ; n22192_not
g71734 not n34324 ; n34324_not
g71735 not n52405 ; n52405_not
g71736 not n14038 ; n14038_not
g71737 not n13534 ; n13534_not
g71738 not n34261 ; n34261_not
g71739 not n41047 ; n41047_not
g71740 not n13444 ; n13444_not
g71741 not n44008 ; n44008_not
g71742 not n22066 ; n22066_not
g71743 not n13624 ; n13624_not
g71744 not n22057 ; n22057_not
g71745 not n34144 ; n34144_not
g71746 not n13615 ; n13615_not
g71747 not n22147 ; n22147_not
g71748 not n50092 ; n50092_not
g71749 not n34207 ; n34207_not
g71750 not n22264 ; n22264_not
g71751 not n22075 ; n22075_not
g71752 not n47005 ; n47005_not
g71753 not n13804 ; n13804_not
g71754 not n14065 ; n14065_not
g71755 not n13606 ; n13606_not
g71756 not n52432 ; n52432_not
g71757 not n40732 ; n40732_not
g71758 not n22291 ; n22291_not
g71759 not n13831 ; n13831_not
g71760 not n13822 ; n13822_not
g71761 not n14056 ; n14056_not
g71762 not n13480 ; n13480_not
g71763 not n34306 ; n34306_not
g71764 not n34270 ; n34270_not
g71765 not n38212 ; n38212_not
g71766 not n34153 ; n34153_not
g71767 not n13372 ; n13372_not
g71768 not n38311 ; n38311_not
g71769 not n37060 ; n37060_not
g71770 not n34045 ; n34045_not
g71771 not n34126 ; n34126_not
g71772 not n50911 ; n50911_not
g71773 not n50128 ; n50128_not
g71774 not n22831 ; n22831_not
g71775 not n34081 ; n34081_not
g71776 not n13381 ; n13381_not
g71777 not n13633 ; n13633_not
g71778 not n34063 ; n34063_not
g71779 not n13282 ; n13282_not
g71780 not n13192 ; n13192_not
g71781 not n22282 ; n22282_not
g71782 not n13417 ; n13417_not
g71783 not n34036 ; n34036_not
g71784 not n13741 ; n13741_not
g71785 not n13507 ; n13507_not
g71786 not n13273 ; n13273_not
g71787 not n34180 ; n34180_not
g71788 not n13714 ; n13714_not
g71789 not n38302 ; n38302_not
g71790 not n52414 ; n52414_not
g71791 not n13147 ; n13147_not
g71792 not n34243 ; n34243_not
g71793 not n13705 ; n13705_not
g71794 not n22156 ; n22156_not
g71795 not n34225 ; n34225_not
g71796 not n41074 ; n41074_not
g71797 not n50038 ; n50038_not
g71798 not n22165 ; n22165_not
g71799 not n13390 ; n13390_not
g71800 not n13183 ; n13183_not
g71801 not n38230 ; n38230_not
g71802 not n13930 ; n13930_not
g71803 not n34072 ; n34072_not
g71804 not n13921 ; n13921_not
g71805 not n34090 ; n34090_not
g71806 not n13471 ; n13471_not
g71807 not n50065 ; n50065_not
g71808 not n50821 ; n50821_not
g71809 not n13363 ; n13363_not
g71810 not n13408 ; n13408_not
g71811 not n22219 ; n22219_not
g71812 not n13912 ; n13912_not
g71813 not n34315 ; n34315_not
g71814 not n14029 ; n14029_not
g71815 not n41065 ; n41065_not
g71816 not n34171 ; n34171_not
g71817 not n50029 ; n50029_not
g71818 not n37240 ; n37240_not
g71819 not n47203 ; n47203_not
g71820 not n40705 ; n40705_not
g71821 not n47212 ; n47212_not
g71822 not n37231 ; n37231_not
g71823 not n22804 ; n22804_not
g71824 not n34162 ; n34162_not
g71825 not n13291 ; n13291_not
g71826 not n34252 ; n34252_not
g71827 not n50830 ; n50830_not
g71828 not n38050 ; n38050_not
g71829 not n13426 ; n13426_not
g71830 not n37222 ; n37222_not
g71831 not n13246 ; n13246_not
g71832 not n38221 ; n38221_not
g71833 not n13435 ; n13435_not
g71834 not n13723 ; n13723_not
g71835 not n38041 ; n38041_not
g71836 not n13462 ; n13462_not
g71837 not n41092 ; n41092_not
g71838 not n52441 ; n52441_not
g71839 not n41128 ; n41128_not
g71840 not n20680 ; n20680_not
g71841 not n43162 ; n43162_not
g71842 not n15361 ; n15361_not
g71843 not n15352 ; n15352_not
g71844 not n30148 ; n30148_not
g71845 not n53413 ; n53413_not
g71846 not n15343 ; n15343_not
g71847 not n30319 ; n30319_not
g71848 not n41317 ; n41317_not
g71849 not n15334 ; n15334_not
g71850 not n33352 ; n33352_not
g71851 not n30157 ; n30157_not
g71852 not n15325 ; n15325_not
g71853 not n15316 ; n15316_not
g71854 not n41308 ; n41308_not
g71855 not n15145 ; n15145_not
g71856 not n41290 ; n41290_not
g71857 not n15262 ; n15262_not
g71858 not n30184 ; n30184_not
g71859 not n20635 ; n20635_not
g71860 not n15271 ; n15271_not
g71861 not n15280 ; n15280_not
g71862 not n43504 ; n43504_not
g71863 not n33046 ; n33046_not
g71864 not n15163 ; n15163_not
g71865 not n30175 ; n30175_not
g71866 not n20644 ; n20644_not
g71867 not n33370 ; n33370_not
g71868 not n15154 ; n15154_not
g71869 not n20653 ; n20653_not
g71870 not n15307 ; n15307_not
g71871 not n30166 ; n30166_not
g71872 not n45061 ; n45061_not
g71873 not n15073 ; n15073_not
g71874 not n15451 ; n15451_not
g71875 not n43450 ; n43450_not
g71876 not n15064 ; n15064_not
g71877 not n15460 ; n15460_not
g71878 not n33262 ; n33262_not
g71879 not n53431 ; n53431_not
g71880 not n41353 ; n41353_not
g71881 not n20725 ; n20725_not
g71882 not n15055 ; n15055_not
g71883 not n43441 ; n43441_not
g71884 not n20734 ; n20734_not
g71885 not n41362 ; n41362_not
g71886 not n20743 ; n20743_not
g71887 not n55114 ; n55114_not
g71888 not n33334 ; n33334_not
g71889 not n15118 ; n15118_not
g71890 not n15370 ; n15370_not
g71891 not n33325 ; n33325_not
g71892 not n30328 ; n30328_not
g71893 not n15109 ; n15109_not
g71894 not n43171 ; n43171_not
g71895 not n33307 ; n33307_not
g71896 not n15406 ; n15406_not
g71897 not n41335 ; n41335_not
g71898 not n43180 ; n43180_not
g71899 not n15415 ; n15415_not
g71900 not n55105 ; n55105_not
g71901 not n15424 ; n15424_not
g71902 not n15433 ; n15433_not
g71903 not n33280 ; n33280_not
g71904 not n15442 ; n15442_not
g71905 not n43117 ; n43117_not
g71906 not n55060 ; n55060_not
g71907 not n43126 ; n43126_not
g71908 not n30247 ; n30247_not
g71909 not n15019 ; n15019_not
g71910 not n41263 ; n41263_not
g71911 not n30265 ; n30265_not
g71912 not n47500 ; n47500_not
g71913 not n30238 ; n30238_not
g71914 not n15037 ; n15037_not
g71915 not n43540 ; n43540_not
g71916 not n43135 ; n43135_not
g71917 not n54700 ; n54700_not
g71918 not n30274 ; n30274_not
g71919 not n20545 ; n20545_not
g71920 not n48004 ; n48004_not
g71921 not n30256 ; n30256_not
g71922 not n21274 ; n21274_not
g71923 not n14380 ; n14380_not
g71924 not n21256 ; n21256_not
g71925 not n14920 ; n14920_not
g71926 not n21265 ; n21265_not
g71927 not n14371 ; n14371_not
g71928 not n37006 ; n37006_not
g71929 not n53350 ; n53350_not
g71930 not n14362 ; n14362_not
g71931 not n20509 ; n20509_not
g71932 not n14344 ; n14344_not
g71933 not n20518 ; n20518_not
g71934 not n45052 ; n45052_not
g71935 not n15172 ; n15172_not
g71936 not n50308 ; n50308_not
g71937 not n20608 ; n20608_not
g71938 not n15190 ; n15190_not
g71939 not n43522 ; n43522_not
g71940 not n37420 ; n37420_not
g71941 not n15217 ; n15217_not
g71942 not n30193 ; n30193_not
g71943 not n15226 ; n15226_not
g71944 not n15235 ; n15235_not
g71945 not n43513 ; n43513_not
g71946 not n15244 ; n15244_not
g71947 not n15253 ; n15253_not
g71948 not n47230 ; n47230_not
g71949 not n37402 ; n37402_not
g71950 not n30229 ; n30229_not
g71951 not n20554 ; n20554_not
g71952 not n15082 ; n15082_not
g71953 not n20563 ; n20563_not
g71954 not n43531 ; n43531_not
g71955 not n41272 ; n41272_not
g71956 not n33343 ; n33343_not
g71957 not n15127 ; n15127_not
g71958 not n37411 ; n37411_not
g71959 not n20590 ; n20590_not
g71960 not n30292 ; n30292_not
g71961 not n43207 ; n43207_not
g71962 not n30454 ; n30454_not
g71963 not n32605 ; n32605_not
g71964 not n43216 ; n43216_not
g71965 not n41425 ; n41425_not
g71966 not n54502 ; n54502_not
g71967 not n43234 ; n43234_not
g71968 not n50272 ; n50272_not
g71969 not n30445 ; n30445_not
g71970 not n54511 ; n54511_not
g71971 not n43252 ; n43252_not
g71972 not n37141 ; n37141_not
g71973 not n43261 ; n43261_not
g71974 not n54520 ; n54520_not
g71975 not n15802 ; n15802_not
g71976 not n43315 ; n43315_not
g71977 not n30283 ; n30283_not
g71978 not n43306 ; n43306_not
g71979 not n20491 ; n20491_not
g71980 not n43270 ; n43270_not
g71981 not n30427 ; n30427_not
g71982 not n50281 ; n50281_not
g71983 not n15820 ; n15820_not
g71984 not n30436 ; n30436_not
g71985 not n15811 ; n15811_not
g71986 not n41407 ; n41407_not
g71987 not n32920 ; n32920_not
g71988 not n15712 ; n15712_not
g71989 not n41452 ; n41452_not
g71990 not n30463 ; n30463_not
g71991 not n52720 ; n52720_not
g71992 not n30490 ; n30490_not
g71993 not n43144 ; n43144_not
g71994 not n32650 ; n32650_not
g71995 not n41461 ; n41461_not
g71996 not n53530 ; n53530_not
g71997 not n19510 ; n19510_not
g71998 not n47122 ; n47122_not
g71999 not n19501 ; n19501_not
g72000 not n41416 ; n41416_not
g72001 not n41470 ; n41470_not
g72002 not n30508 ; n30508_not
g72003 not n45106 ; n45106_not
g72004 not n45142 ; n45142_not
g72005 not n53503 ; n53503_not
g72006 not n32614 ; n32614_not
g72007 not n47113 ; n47113_not
g72008 not n32623 ; n32623_not
g72009 not n41443 ; n41443_not
g72010 not n15730 ; n15730_not
g72011 not n53521 ; n53521_not
g72012 not n50263 ; n50263_not
g72013 not n19600 ; n19600_not
g72014 not n15721 ; n15721_not
g72015 not n30472 ; n30472_not
g72016 not n15541 ; n15541_not
g72017 not n15550 ; n15550_not
g72018 not n41380 ; n41380_not
g72019 not n43423 ; n43423_not
g72020 not n20752 ; n20752_not
g72021 not n30373 ; n30373_not
g72022 not n43414 ; n43414_not
g72023 not n43405 ; n43405_not
g72024 not n15613 ; n15613_not
g72025 not n15622 ; n15622_not
g72026 not n37501 ; n37501_not
g72027 not n15631 ; n15631_not
g72028 not n20707 ; n20707_not
g72029 not n44800 ; n44800_not
g72030 not n54610 ; n54610_not
g72031 not n43432 ; n43432_not
g72032 not n15505 ; n15505_not
g72033 not n53440 ; n53440_not
g72034 not n15514 ; n15514_not
g72035 not n55123 ; n55123_not
g72036 not n30355 ; n30355_not
g72037 not n20770 ; n20770_not
g72038 not n15523 ; n15523_not
g72039 not n15028 ; n15028_not
g72040 not n15532 ; n15532_not
g72041 not n30364 ; n30364_not
g72042 not n54601 ; n54601_not
g72043 not n30409 ; n30409_not
g72044 not n20572 ; n20572_not
g72045 not n33037 ; n33037_not
g72046 not n43333 ; n43333_not
g72047 not n30418 ; n30418_not
g72048 not n33028 ; n33028_not
g72049 not n33019 ; n33019_not
g72050 not n55150 ; n55150_not
g72051 not n15208 ; n15208_not
g72052 not n43324 ; n43324_not
g72053 not n20527 ; n20527_not
g72054 not n30382 ; n30382_not
g72055 not n30391 ; n30391_not
g72056 not n20662 ; n20662_not
g72057 not n43225 ; n43225_not
g72058 not n20617 ; n20617_not
g72059 not n43360 ; n43360_not
g72060 not n43351 ; n43351_not
g72061 not n43342 ; n43342_not
g72062 not n14326 ; n14326_not
g72063 not n21355 ; n21355_not
g72064 not n21535 ; n21535_not
g72065 not n50227 ; n50227_not
g72066 not n14317 ; n14317_not
g72067 not n13750 ; n13750_not
g72068 not n50218 ; n50218_not
g72069 not n14308 ; n14308_not
g72070 not n41173 ; n41173_not
g72071 not n14290 ; n14290_not
g72072 not n37321 ; n37321_not
g72073 not n33901 ; n33901_not
g72074 not n30058 ; n30058_not
g72075 not n14254 ; n14254_not
g72076 not n14263 ; n14263_not
g72077 not n21319 ; n21319_not
g72078 not n30049 ; n30049_not
g72079 not n21328 ; n21328_not
g72080 not n53260 ; n53260_not
g72081 not n14272 ; n14272_not
g72082 not n14281 ; n14281_not
g72083 not n37330 ; n37330_not
g72084 not n41191 ; n41191_not
g72085 not n14407 ; n14407_not
g72086 not n14416 ; n14416_not
g72087 not n14434 ; n14434_not
g72088 not n40642 ; n40642_not
g72089 not n33820 ; n33820_not
g72090 not n21409 ; n21409_not
g72091 not n30139 ; n30139_not
g72092 not n21418 ; n21418_not
g72093 not n40660 ; n40660_not
g72094 not n41182 ; n41182_not
g72095 not n21364 ; n21364_not
g72096 not n48031 ; n48031_not
g72097 not n21373 ; n21373_not
g72098 not n50245 ; n50245_not
g72099 not n40651 ; n40651_not
g72100 not n38203 ; n38203_not
g72101 not n14146 ; n14146_not
g72102 not n13840 ; n13840_not
g72103 not n14155 ; n14155_not
g72104 not n30076 ; n30076_not
g72105 not n14164 ; n14164_not
g72106 not n33631 ; n33631_not
g72107 not n50173 ; n50173_not
g72108 not n22039 ; n22039_not
g72109 not n14173 ; n14173_not
g72110 not n33640 ; n33640_not
g72111 not n14182 ; n14182_not
g72112 not n50137 ; n50137_not
g72113 not n37051 ; n37051_not
g72114 not n14074 ; n14074_not
g72115 not n14083 ; n14083_not
g72116 not n33613 ; n33613_not
g72117 not n14092 ; n14092_not
g72118 not n22129 ; n22129_not
g72119 not n37303 ; n37303_not
g72120 not n50155 ; n50155_not
g72121 not n14119 ; n14119_not
g72122 not n33622 ; n33622_not
g72123 not n41137 ; n41137_not
g72124 not n14128 ; n14128_not
g72125 not n14137 ; n14137_not
g72126 not n22084 ; n22084_not
g72127 not n30085 ; n30085_not
g72128 not n43801 ; n43801_not
g72129 not n14227 ; n14227_not
g72130 not n41155 ; n41155_not
g72131 not n33910 ; n33910_not
g72132 not n30067 ; n30067_not
g72133 not n14236 ; n14236_not
g72134 not n14245 ; n14245_not
g72135 not n53251 ; n53251_not
g72136 not n41164 ; n41164_not
g72137 not n50182 ; n50182_not
g72138 not n14191 ; n14191_not
g72139 not n37312 ; n37312_not
g72140 not n53242 ; n53242_not
g72141 not n41146 ; n41146_not
g72142 not n14209 ; n14209_not
g72143 not n21283 ; n21283_not
g72144 not n14218 ; n14218_not
g72145 not n14722 ; n14722_not
g72146 not n21454 ; n21454_not
g72147 not n21445 ; n21445_not
g72148 not n14731 ; n14731_not
g72149 not n50326 ; n50326_not
g72150 not n37015 ; n37015_not
g72151 not n14740 ; n14740_not
g72152 not n21427 ; n21427_not
g72153 not n30094 ; n30094_not
g72154 not n14470 ; n14470_not
g72155 not n14461 ; n14461_not
g72156 not n43072 ; n43072_not
g72157 not n14452 ; n14452_not
g72158 not n55015 ; n55015_not
g72159 not n14650 ; n14650_not
g72160 not n38104 ; n38104_not
g72161 not n21517 ; n21517_not
g72162 not n14515 ; n14515_not
g72163 not n45016 ; n45016_not
g72164 not n14506 ; n14506_not
g72165 not n21490 ; n21490_not
g72166 not n14704 ; n14704_not
g72167 not n41245 ; n41245_not
g72168 not n21472 ; n21472_not
g72169 not n50317 ; n50317_not
g72170 not n53341 ; n53341_not
g72171 not n14713 ; n14713_not
g72172 not n21337 ; n21337_not
g72173 not n33604 ; n33604_not
g72174 not n43621 ; n43621_not
g72175 not n55024 ; n55024_not
g72176 not n43090 ; n43090_not
g72177 not n48013 ; n48013_not
g72178 not n55033 ; n55033_not
g72179 not n43612 ; n43612_not
g72180 not n43603 ; n43603_not
g72181 not n45034 ; n45034_not
g72182 not n21292 ; n21292_not
g72183 not n14902 ; n14902_not
g72184 not n14911 ; n14911_not
g72185 not n21382 ; n21382_not
g72186 not n14803 ; n14803_not
g72187 not n14812 ; n14812_not
g72188 not n14821 ; n14821_not
g72189 not n43630 ; n43630_not
g72190 not n14830 ; n14830_not
g72191 not n43081 ; n43081_not
g72192 not n14425 ; n14425_not
g72193 not n14524 ; n14524_not
g72194 not n47401 ; n47401_not
g72195 not n14542 ; n14542_not
g72196 not n33721 ; n33721_not
g72197 not n44332 ; n44332_not
g72198 not n21463 ; n21463_not
g72199 not n14551 ; n14551_not
g72200 not n33730 ; n33730_not
g72201 not n41218 ; n41218_not
g72202 not n33811 ; n33811_not
g72203 not n41209 ; n41209_not
g72204 not n33802 ; n33802_not
g72205 not n33712 ; n33712_not
g72206 not n53305 ; n53305_not
g72207 not n41227 ; n41227_not
g72208 not n21508 ; n21508_not
g72209 not n14614 ; n14614_not
g72210 not n14623 ; n14623_not
g72211 not n14632 ; n14632_not
g72212 not n14641 ; n14641_not
g72213 not n50290 ; n50290_not
g72214 not n45007 ; n45007_not
g72215 not n47410 ; n47410_not
g72216 not n53323 ; n53323_not
g72217 not n14560 ; n14560_not
g72218 not n43711 ; n43711_not
g72219 not n14605 ; n14605_not
g72220 not n37024 ; n37024_not
g72221 not n24802 ; n24802_not
g72222 not n10852 ; n10852_not
g72223 not n28420 ; n28420_not
g72224 not n52171 ; n52171_not
g72225 not n52162 ; n52162_not
g72226 not n35332 ; n35332_not
g72227 not n40327 ; n40327_not
g72228 not n35323 ; n35323_not
g72229 not n52153 ; n52153_not
g72230 not n40336 ; n40336_not
g72231 not n52144 ; n52144_not
g72232 not n52135 ; n52135_not
g72233 not n25504 ; n25504_not
g72234 not n40345 ; n40345_not
g72235 not n52126 ; n52126_not
g72236 not n10357 ; n10357_not
g72237 not n25450 ; n25450_not
g72238 not n28402 ; n28402_not
g72239 not n49201 ; n49201_not
g72240 not n40255 ; n40255_not
g72241 not n51613 ; n51613_not
g72242 not n10339 ; n10339_not
g72243 not n52180 ; n52180_not
g72244 not n40309 ; n40309_not
g72245 not n24820 ; n24820_not
g72246 not n10861 ; n10861_not
g72247 not n35350 ; n35350_not
g72248 not n24811 ; n24811_not
g72249 not n28411 ; n28411_not
g72250 not n10870 ; n10870_not
g72251 not n40318 ; n40318_not
g72252 not n10942 ; n10942_not
g72253 not n52603 ; n52603_not
g72254 not n52117 ; n52117_not
g72255 not n35017 ; n35017_not
g72256 not n52108 ; n52108_not
g72257 not n40228 ; n40228_not
g72258 not n52612 ; n52612_not
g72259 not n35026 ; n35026_not
g72260 not n10960 ; n10960_not
g72261 not n40363 ; n40363_not
g72262 not n35035 ; n35035_not
g72263 not n40219 ; n40219_not
g72264 not n52090 ; n52090_not
g72265 not n35044 ; n35044_not
g72266 not n35053 ; n35053_not
g72267 not n28312 ; n28312_not
g72268 not n35305 ; n35305_not
g72269 not n10915 ; n10915_not
g72270 not n49120 ; n49120_not
g72271 not n24730 ; n24730_not
g72272 not n25531 ; n25531_not
g72273 not n10924 ; n10924_not
g72274 not n40354 ; n40354_not
g72275 not n49111 ; n49111_not
g72276 not n24703 ; n24703_not
g72277 not n35008 ; n35008_not
g72278 not n24721 ; n24721_not
g72279 not n44314 ; n44314_not
g72280 not n25513 ; n25513_not
g72281 not n51604 ; n51604_not
g72282 not n52315 ; n52315_not
g72283 not n52306 ; n52306_not
g72284 not n25036 ; n25036_not
g72285 not n10447 ; n10447_not
g72286 not n28303 ; n28303_not
g72287 not n25351 ; n25351_not
g72288 not n25027 ; n25027_not
g72289 not n40192 ; n40192_not
g72290 not n45025 ; n45025_not
g72291 not n25018 ; n25018_not
g72292 not n25360 ; n25360_not
g72293 not n25009 ; n25009_not
g72294 not n35404 ; n35404_not
g72295 not n44341 ; n44341_not
g72296 not n52513 ; n52513_not
g72297 not n28330 ; n28330_not
g72298 not n52351 ; n52351_not
g72299 not n25324 ; n25324_not
g72300 not n25081 ; n25081_not
g72301 not n40165 ; n40165_not
g72302 not n52342 ; n52342_not
g72303 not n56302 ; n56302_not
g72304 not n35413 ; n35413_not
g72305 not n25072 ; n25072_not
g72306 not n52333 ; n52333_not
g72307 not n25063 ; n25063_not
g72308 not n40174 ; n40174_not
g72309 not n52324 ; n52324_not
g72310 not n10465 ; n10465_not
g72311 not n25054 ; n25054_not
g72312 not n10456 ; n10456_not
g72313 not n25045 ; n25045_not
g72314 not n24910 ; n24910_not
g72315 not n40264 ; n40264_not
g72316 not n24901 ; n24901_not
g72317 not n52225 ; n52225_not
g72318 not n38500 ; n38500_not
g72319 not n49210 ; n49210_not
g72320 not n52216 ; n52216_not
g72321 not n10375 ; n10375_not
g72322 not n52207 ; n52207_not
g72323 not n40273 ; n40273_not
g72324 not n10366 ; n10366_not
g72325 not n40282 ; n40282_not
g72326 not n25441 ; n25441_not
g72327 not n40291 ; n40291_not
g72328 not n52270 ; n52270_not
g72329 not n51640 ; n51640_not
g72330 not n52522 ; n52522_not
g72331 not n52261 ; n52261_not
g72332 not n40237 ; n40237_not
g72333 not n52252 ; n52252_not
g72334 not n51631 ; n51631_not
g72335 not n52243 ; n52243_not
g72336 not n48400 ; n48400_not
g72337 not n25405 ; n25405_not
g72338 not n52234 ; n52234_not
g72339 not n52540 ; n52540_not
g72340 not n25414 ; n25414_not
g72341 not n25171 ; n25171_not
g72342 not n25180 ; n25180_not
g72343 not n25261 ; n25261_not
g72344 not n51541 ; n51541_not
g72345 not n52018 ; n52018_not
g72346 not n43702 ; n43702_not
g72347 not n25207 ; n25207_not
g72348 not n25216 ; n25216_not
g72349 not n25243 ; n25243_not
g72350 not n11239 ; n11239_not
g72351 not n25234 ; n25234_not
g72352 not n11248 ; n11248_not
g72353 not n56032 ; n56032_not
g72354 not n25225 ; n25225_not
g72355 not n35161 ; n35161_not
g72356 not n25108 ; n25108_not
g72357 not n49102 ; n49102_not
g72358 not n11185 ; n11185_not
g72359 not n25117 ; n25117_not
g72360 not n40408 ; n40408_not
g72361 not n35170 ; n35170_not
g72362 not n25126 ; n25126_not
g72363 not n25135 ; n25135_not
g72364 not n11194 ; n11194_not
g72365 not n25144 ; n25144_not
g72366 not n25153 ; n25153_not
g72367 not n45070 ; n45070_not
g72368 not n25162 ; n25162_not
g72369 not n25270 ; n25270_not
g72370 not n35143 ; n35143_not
g72371 not n11338 ; n11338_not
g72372 not n24451 ; n24451_not
g72373 not n11347 ; n11347_not
g72374 not n52009 ; n52009_not
g72375 not n11356 ; n11356_not
g72376 not n56041 ; n56041_not
g72377 not n11365 ; n11365_not
g72378 not n24460 ; n24460_not
g72379 not n51514 ; n51514_not
g72380 not n11374 ; n11374_not
g72381 not n35134 ; n35134_not
g72382 not n11383 ; n11383_not
g72383 not n48301 ; n48301_not
g72384 not n11392 ; n11392_not
g72385 not n35125 ; n35125_not
g72386 not n40426 ; n40426_not
g72387 not n11419 ; n11419_not
g72388 not n11257 ; n11257_not
g72389 not n48310 ; n48310_not
g72390 not n51532 ; n51532_not
g72391 not n11266 ; n11266_not
g72392 not n11275 ; n11275_not
g72393 not n24415 ; n24415_not
g72394 not n11284 ; n11284_not
g72395 not n24424 ; n24424_not
g72396 not n11293 ; n11293_not
g72397 not n40417 ; n40417_not
g72398 not n28240 ; n28240_not
g72399 not n28600 ; n28600_not
g72400 not n35152 ; n35152_not
g72401 not n51523 ; n51523_not
g72402 not n10933 ; n10933_not
g72403 not n56230 ; n56230_not
g72404 not n11329 ; n11329_not
g72405 not n52063 ; n52063_not
g72406 not n44305 ; n44305_not
g72407 not n35233 ; n35233_not
g72408 not n35107 ; n35107_not
g72409 not n52054 ; n52054_not
g72410 not n35116 ; n35116_not
g72411 not n40390 ; n40390_not
g72412 not n52045 ; n52045_not
g72413 not n56023 ; n56023_not
g72414 not n52036 ; n52036_not
g72415 not n11059 ; n11059_not
g72416 not n40372 ; n40372_not
g72417 not n35260 ; n35260_not
g72418 not n35062 ; n35062_not
g72419 not n52081 ; n52081_not
g72420 not n35071 ; n35071_not
g72421 not n28501 ; n28501_not
g72422 not n40381 ; n40381_not
g72423 not n28510 ; n28510_not
g72424 not n35080 ; n35080_not
g72425 not n52072 ; n52072_not
g72426 not n52630 ; n52630_not
g72427 not n25423 ; n25423_not
g72428 not n35242 ; n35242_not
g72429 not n25333 ; n25333_not
g72430 not n11149 ; n11149_not
g72431 not n11158 ; n11158_not
g72432 not n11167 ; n11167_not
g72433 not n25315 ; n25315_not
g72434 not n25090 ; n25090_not
g72435 not n11176 ; n11176_not
g72436 not n25306 ; n25306_not
g72437 not n52027 ; n52027_not
g72438 not n51550 ; n51550_not
g72439 not n46501 ; n46501_not
g72440 not n11077 ; n11077_not
g72441 not n11086 ; n11086_not
g72442 not n11095 ; n11095_not
g72443 not n35215 ; n35215_not
g72444 not n36214 ; n36214_not
g72445 not n26071 ; n26071_not
g72446 not n46141 ; n46141_not
g72447 not n36403 ; n36403_not
g72448 not n26080 ; n26080_not
g72449 not n46240 ; n46240_not
g72450 not n36412 ; n36412_not
g72451 not n51901 ; n51901_not
g72452 not n36421 ; n36421_not
g72453 not n46132 ; n46132_not
g72454 not n46510 ; n46510_not
g72455 not n46231 ; n46231_not
g72456 not n36430 ; n36430_not
g72457 not n46222 ; n46222_not
g72458 not n46123 ; n46123_not
g72459 not n36007 ; n36007_not
g72460 not n49003 ; n49003_not
g72461 not n27025 ; n27025_not
g72462 not n46213 ; n46213_not
g72463 not n57130 ; n57130_not
g72464 not n27016 ; n27016_not
g72465 not n49012 ; n49012_not
g72466 not n46204 ; n46204_not
g72467 not n57121 ; n57121_not
g72468 not n49021 ; n49021_not
g72469 not n27007 ; n27007_not
g72470 not n39310 ; n39310_not
g72471 not n39301 ; n39301_not
g72472 not n39103 ; n39103_not
g72473 not n49030 ; n49030_not
g72474 not n46150 ; n46150_not
g72475 not n51721 ; n51721_not
g72476 not n36052 ; n36052_not
g72477 not n26161 ; n26161_not
g72478 not n51712 ; n51712_not
g72479 not n26170 ; n26170_not
g72480 not n36043 ; n36043_not
g72481 not n36502 ; n36502_not
g72482 not n39220 ; n39220_not
g72483 not n35800 ; n35800_not
g72484 not n36511 ; n36511_not
g72485 not n51703 ; n51703_not
g72486 not n39211 ; n39211_not
g72487 not n57022 ; n57022_not
g72488 not n26107 ; n26107_not
g72489 not n57004 ; n57004_not
g72490 not n35701 ; n35701_not
g72491 not n26116 ; n26116_not
g72492 not n26125 ; n26125_not
g72493 not n46114 ; n46114_not
g72494 not n51910 ; n51910_not
g72495 not n51127 ; n51127_not
g72496 not n46105 ; n46105_not
g72497 not n39130 ; n39130_not
g72498 not n26152 ; n26152_not
g72499 not n27205 ; n27205_not
g72500 not n27115 ; n27115_not
g72501 not n46312 ; n46312_not
g72502 not n27106 ; n27106_not
g72503 not n27223 ; n27223_not
g72504 not n27214 ; n27214_not
g72505 not n46303 ; n46303_not
g72506 not n36151 ; n36151_not
g72507 not n36304 ; n36304_not
g72508 not n46420 ; n46420_not
g72509 not n39013 ; n39013_not
g72510 not n36133 ; n36133_not
g72511 not n39004 ; n39004_not
g72512 not n36313 ; n36313_not
g72513 not n27151 ; n27151_not
g72514 not n36250 ; n36250_not
g72515 not n27142 ; n27142_not
g72516 not n39040 ; n39040_not
g72517 not n39400 ; n39400_not
g72518 not n27160 ; n27160_not
g72519 not n46330 ; n46330_not
g72520 not n36241 ; n36241_not
g72521 not n36232 ; n36232_not
g72522 not n44503 ; n44503_not
g72523 not n46402 ; n46402_not
g72524 not n46321 ; n46321_not
g72525 not n44512 ; n44512_not
g72526 not n36205 ; n36205_not
g72527 not n36061 ; n36061_not
g72528 not n27052 ; n27052_not
g72529 not n51802 ; n51802_not
g72530 not n27061 ; n27061_not
g72531 not n57220 ; n57220_not
g72532 not n57211 ; n57211_not
g72533 not n27034 ; n27034_not
g72534 not n35611 ; n35611_not
g72535 not n57202 ; n57202_not
g72536 not n36025 ; n36025_not
g72537 not n36124 ; n36124_not
g72538 not n36016 ; n36016_not
g72539 not n27070 ; n27070_not
g72540 not n27124 ; n27124_not
g72541 not n57310 ; n57310_not
g72542 not n36106 ; n36106_not
g72543 not n36322 ; n36322_not
g72544 not n36142 ; n36142_not
g72545 not n51811 ; n51811_not
g72546 not n36331 ; n36331_not
g72547 not n45700 ; n45700_not
g72548 not n36340 ; n36340_not
g72549 not n40066 ; n40066_not
g72550 not n35251 ; n35251_not
g72551 not n28213 ; n28213_not
g72552 not n40057 ; n40057_not
g72553 not n26062 ; n26062_not
g72554 not n56320 ; n56320_not
g72555 not n28231 ; n28231_not
g72556 not n40048 ; n40048_not
g72557 not n26206 ; n26206_not
g72558 not n56410 ; n56410_not
g72559 not n35530 ; n35530_not
g72560 not n56401 ; n56401_not
g72561 not n35521 ; n35521_not
g72562 not n40075 ; n40075_not
g72563 not n35512 ; n35512_not
g72564 not n28204 ; n28204_not
g72565 not n26134 ; n26134_not
g72566 not n40084 ; n40084_not
g72567 not n52423 ; n52423_not
g72568 not n35503 ; n35503_not
g72569 not n35440 ; n35440_not
g72570 not n10519 ; n10519_not
g72571 not n40129 ; n40129_not
g72572 not n56311 ; n56311_not
g72573 not n40147 ; n40147_not
g72574 not n35431 ; n35431_not
g72575 not n10492 ; n10492_not
g72576 not n52360 ; n52360_not
g72577 not n35422 ; n35422_not
g72578 not n40039 ; n40039_not
g72579 not n10384 ; n10384_not
g72580 not n10429 ; n10429_not
g72581 not n10474 ; n10474_not
g72582 not n52450 ; n52450_not
g72583 not n46042 ; n46042_not
g72584 not n46033 ; n46033_not
g72585 not n26251 ; n26251_not
g72586 not n46024 ; n46024_not
g72587 not n26260 ; n26260_not
g72588 not n46015 ; n46015_not
g72589 not n35710 ; n35710_not
g72590 not n44521 ; n44521_not
g72591 not n46006 ; n46006_not
g72592 not n46600 ; n46600_not
g72593 not n45250 ; n45250_not
g72594 not n46060 ; n46060_not
g72595 not n39202 ; n39202_not
g72596 not n26215 ; n26215_not
g72597 not n46051 ; n46051_not
g72598 not n51820 ; n51820_not
g72599 not n36601 ; n36601_not
g72600 not n26242 ; n26242_not
g72601 not n26332 ; n26332_not
g72602 not n35620 ; n35620_not
g72603 not n26314 ; n26314_not
g72604 not n28114 ; n28114_not
g72605 not n28123 ; n28123_not
g72606 not n35602 ; n35602_not
g72607 not n28132 ; n28132_not
g72608 not n56500 ; n56500_not
g72609 not n35206 ; n35206_not
g72610 not n44431 ; n44431_not
g72611 not n28141 ; n28141_not
g72612 not n39022 ; n39022_not
g72613 not n28015 ; n28015_not
g72614 not n28006 ; n28006_not
g72615 not n26224 ; n26224_not
g72616 not n44413 ; n44413_not
g72617 not n44404 ; n44404_not
g72618 not n44602 ; n44602_not
g72619 not n39112 ; n39112_not
g72620 not n26305 ; n26305_not
g72621 not n26341 ; n26341_not
g72622 not n26350 ; n26350_not
g72623 not n28033 ; n28033_not
g72624 not n36700 ; n36700_not
g72625 not n28051 ; n28051_not
g72626 not n28060 ; n28060_not
g72627 not n51730 ; n51730_not
g72628 not n51208 ; n51208_not
g72629 not n40921 ; n40921_not
g72630 not n22822 ; n22822_not
g72631 not n12265 ; n12265_not
g72632 not n44125 ; n44125_not
g72633 not n23560 ; n23560_not
g72634 not n23551 ; n23551_not
g72635 not n51064 ; n51064_not
g72636 not n12274 ; n12274_not
g72637 not n23542 ; n23542_not
g72638 not n51190 ; n51190_not
g72639 not n56050 ; n56050_not
g72640 not n23533 ; n23533_not
g72641 not n29401 ; n29401_not
g72642 not n40930 ; n40930_not
g72643 not n12283 ; n12283_not
g72644 not n23524 ; n23524_not
g72645 not n44116 ; n44116_not
g72646 not n12292 ; n12292_not
g72647 not n29311 ; n29311_not
g72648 not n12733 ; n12733_not
g72649 not n23641 ; n23641_not
g72650 not n29320 ; n29320_not
g72651 not n40912 ; n40912_not
g72652 not n34603 ; n34603_not
g72653 not n47050 ; n47050_not
g72654 not n23623 ; n23623_not
g72655 not n12724 ; n12724_not
g72656 not n23614 ; n23614_not
g72657 not n12229 ; n12229_not
g72658 not n48112 ; n48112_not
g72659 not n12238 ; n12238_not
g72660 not n23605 ; n23605_not
g72661 not n12247 ; n12247_not
g72662 not n12256 ; n12256_not
g72663 not n34522 ; n34522_not
g72664 not n51154 ; n51154_not
g72665 not n23434 ; n23434_not
g72666 not n12337 ; n12337_not
g72667 not n23425 ; n23425_not
g72668 not n51145 ; n51145_not
g72669 not n23416 ; n23416_not
g72670 not n29410 ; n29410_not
g72671 not n22903 ; n22903_not
g72672 not n23407 ; n23407_not
g72673 not n22912 ; n22912_not
g72674 not n34513 ; n34513_not
g72675 not n12346 ; n12346_not
g72676 not n38410 ; n38410_not
g72677 not n12355 ; n12355_not
g72678 not n23380 ; n23380_not
g72679 not n51136 ; n51136_not
g72680 not n23515 ; n23515_not
g72681 not n23506 ; n23506_not
g72682 not n51181 ; n51181_not
g72683 not n34540 ; n34540_not
g72684 not n51073 ; n51073_not
g72685 not n34531 ; n34531_not
g72686 not n34504 ; n34504_not
g72687 not n51172 ; n51172_not
g72688 not n51082 ; n51082_not
g72689 not n23470 ; n23470_not
g72690 not n12319 ; n12319_not
g72691 not n23461 ; n23461_not
g72692 not n44107 ; n44107_not
g72693 not n51163 ; n51163_not
g72694 not n23452 ; n23452_not
g72695 not n45115 ; n45115_not
g72696 not n12328 ; n12328_not
g72697 not n23443 ; n23443_not
g72698 not n29140 ; n29140_not
g72699 not n29131 ; n29131_not
g72700 not n37150 ; n37150_not
g72701 not n40822 ; n40822_not
g72702 not n40831 ; n40831_not
g72703 not n29122 ; n29122_not
g72704 not n12616 ; n12616_not
g72705 not n51253 ; n51253_not
g72706 not n40840 ; n40840_not
g72707 not n51037 ; n51037_not
g72708 not n12634 ; n12634_not
g72709 not n12643 ; n12643_not
g72710 not n12526 ; n12526_not
g72711 not n34702 ; n34702_not
g72712 not n34405 ; n34405_not
g72713 not n12553 ; n12553_not
g72714 not n12535 ; n12535_not
g72715 not n44161 ; n44161_not
g72716 not n40804 ; n40804_not
g72717 not n12571 ; n12571_not
g72718 not n34414 ; n34414_not
g72719 not n34441 ; n34441_not
g72720 not n23713 ; n23713_not
g72721 not n29203 ; n29203_not
g72722 not n23704 ; n23704_not
g72723 not n12193 ; n12193_not
g72724 not n34630 ; n34630_not
g72725 not n51226 ; n51226_not
g72726 not n29212 ; n29212_not
g72727 not n52531 ; n52531_not
g72728 not n34621 ; n34621_not
g72729 not n40903 ; n40903_not
g72730 not n29221 ; n29221_not
g72731 not n34450 ; n34450_not
g72732 not n44134 ; n44134_not
g72733 not n29302 ; n29302_not
g72734 not n12742 ; n12742_not
g72735 not n34612 ; n34612_not
g72736 not n29230 ; n29230_not
g72737 not n44422 ; n44422_not
g72738 not n51217 ; n51217_not
g72739 not n44152 ; n44152_not
g72740 not n12661 ; n12661_not
g72741 not n51244 ; n51244_not
g72742 not n23821 ; n23821_not
g72743 not n23803 ; n23803_not
g72744 not n12706 ; n12706_not
g72745 not n51235 ; n51235_not
g72746 not n47041 ; n47041_not
g72747 not n11635 ; n11635_not
g72748 not n23731 ; n23731_not
g72749 not n44143 ; n44143_not
g72750 not n23092 ; n23092_not
g72751 not n44071 ; n44071_not
g72752 not n23083 ; n23083_not
g72753 not n47023 ; n47023_not
g72754 not n34333 ; n34333_not
g72755 not n23074 ; n23074_not
g72756 not n34342 ; n34342_not
g72757 not n37204 ; n37204_not
g72758 not n13255 ; n13255_not
g72759 not n44062 ; n44062_not
g72760 not n23056 ; n23056_not
g72761 not n34351 ; n34351_not
g72762 not n23038 ; n23038_not
g72763 not n34360 ; n34360_not
g72764 not n51046 ; n51046_not
g72765 not n23029 ; n23029_not
g72766 not n47032 ; n47032_not
g72767 not n38005 ; n38005_not
g72768 not n23146 ; n23146_not
g72769 not n13138 ; n13138_not
g72770 not n23137 ; n23137_not
g72771 not n23128 ; n23128_not
g72772 not n13165 ; n13165_not
g72773 not n23119 ; n23119_not
g72774 not n38014 ; n38014_not
g72775 not n22921 ; n22921_not
g72776 not n44035 ; n44035_not
g72777 not n41029 ; n41029_not
g72778 not n51019 ; n51019_not
g72779 not n13327 ; n13327_not
g72780 not n38320 ; n38320_not
g72781 not n13318 ; n13318_not
g72782 not n44026 ; n44026_not
g72783 not n41038 ; n41038_not
g72784 not n44053 ; n44053_not
g72785 not n44044 ; n44044_not
g72786 not n40750 ; n40750_not
g72787 not n37213 ; n37213_not
g72788 not n13345 ; n13345_not
g72789 not n47014 ; n47014_not
g72790 not n56005 ; n56005_not
g72791 not n51028 ; n51028_not
g72792 not n40741 ; n40741_not
g72793 not n47140 ; n47140_not
g72794 not n13336 ; n13336_not
g72795 not n12391 ; n12391_not
g72796 not n23317 ; n23317_not
g72797 not n23308 ; n23308_not
g72798 not n12409 ; n12409_not
g72799 not n12418 ; n12418_not
g72800 not n23290 ; n23290_not
g72801 not n12427 ; n12427_not
g72802 not n51109 ; n51109_not
g72803 not n23281 ; n23281_not
g72804 not n12436 ; n12436_not
g72805 not n23272 ; n23272_not
g72806 not n12607 ; n12607_not
g72807 not n23371 ; n23371_not
g72808 not n12652 ; n12652_not
g72809 not n12364 ; n12364_not
g72810 not n38401 ; n38401_not
g72811 not n23362 ; n23362_not
g72812 not n23353 ; n23353_not
g72813 not n12373 ; n12373_not
g72814 not n23344 ; n23344_not
g72815 not n37114 ; n37114_not
g72816 not n23335 ; n23335_not
g72817 not n12382 ; n12382_not
g72818 not n48103 ; n48103_not
g72819 not n23326 ; n23326_not
g72820 not n51091 ; n51091_not
g72821 not n12490 ; n12490_not
g72822 not n23209 ; n23209_not
g72823 not n23191 ; n23191_not
g72824 not n12508 ; n12508_not
g72825 not n23182 ; n23182_not
g72826 not n12517 ; n12517_not
g72827 not n34423 ; n34423_not
g72828 not n12562 ; n12562_not
g72829 not n23173 ; n23173_not
g72830 not n23164 ; n23164_not
g72831 not n23047 ; n23047_not
g72832 not n23155 ; n23155_not
g72833 not n12445 ; n12445_not
g72834 not n23263 ; n23263_not
g72835 not n12454 ; n12454_not
g72836 not n23254 ; n23254_not
g72837 not n12463 ; n12463_not
g72838 not n23245 ; n23245_not
g72839 not n37105 ; n37105_not
g72840 not n23236 ; n23236_not
g72841 not n12472 ; n12472_not
g72842 not n23227 ; n23227_not
g72843 not n12481 ; n12481_not
g72844 not n23218 ; n23218_not
g72845 not n44080 ; n44080_not
g72846 not n11482 ; n11482_not
g72847 not n44233 ; n44233_not
g72848 not n40543 ; n40543_not
g72849 not n11860 ; n11860_not
g72850 not n51406 ; n51406_not
g72851 not n48202 ; n48202_not
g72852 not n11473 ; n11473_not
g72853 not n40552 ; n40552_not
g72854 not n44224 ; n44224_not
g72855 not n11905 ; n11905_not
g72856 not n40561 ; n40561_not
g72857 not n11914 ; n11914_not
g72858 not n37033 ; n37033_not
g72859 not n11923 ; n11923_not
g72860 not n28024 ; n28024_not
g72861 not n24631 ; n24631_not
g72862 not n11518 ; n11518_not
g72863 not n11806 ; n11806_not
g72864 not n24640 ; n24640_not
g72865 not n11815 ; n11815_not
g72866 not n44242 ; n44242_not
g72867 not n51415 ; n51415_not
g72868 not n40516 ; n40516_not
g72869 not n11824 ; n11824_not
g72870 not n11833 ; n11833_not
g72871 not n40138 ; n40138_not
g72872 not n40525 ; n40525_not
g72873 not n11842 ; n11842_not
g72874 not n48220 ; n48220_not
g72875 not n11491 ; n11491_not
g72876 not n40534 ; n40534_not
g72877 not n11851 ; n11851_not
g72878 not n48211 ; n48211_not
g72879 not n24613 ; n24613_not
g72880 not n51352 ; n51352_not
g72881 not n34900 ; n34900_not
g72882 not n44206 ; n44206_not
g72883 not n51343 ; n51343_not
g72884 not n11950 ; n11950_not
g72885 not n11941 ; n11941_not
g72886 not n11932 ; n11932_not
g72887 not n51334 ; n51334_not
g72888 not n24550 ; n24550_not
g72889 not n46411 ; n46411_not
g72890 not n24541 ; n24541_not
g72891 not n51325 ; n51325_not
g72892 not n11446 ; n11446_not
g72893 not n11437 ; n11437_not
g72894 not n51370 ; n51370_not
g72895 not n40570 ; n40570_not
g72896 not n51361 ; n51361_not
g72897 not n11428 ; n11428_not
g72898 not n44215 ; n44215_not
g72899 not n11563 ; n11563_not
g72900 not n11572 ; n11572_not
g72901 not n11590 ; n11590_not
g72902 not n11608 ; n11608_not
g72903 not n11617 ; n11617_not
g72904 not n40444 ; n40444_not
g72905 not n11644 ; n11644_not
g72906 not n56221 ; n56221_not
g72907 not n40453 ; n40453_not
g72908 not n52702 ; n52702_not
g72909 not n11653 ; n11653_not
g72910 not n51505 ; n51505_not
g72911 not n40435 ; n40435_not
g72912 not n11455 ; n11455_not
g72913 not n50902 ; n50902_not
g72914 not n24505 ; n24505_not
g72915 not n11527 ; n11527_not
g72916 not n11545 ; n11545_not
g72917 not n24514 ; n24514_not
g72918 not n34810 ; n34810_not
g72919 not n40183 ; n40183_not
g72920 not n11716 ; n11716_not
g72921 not n52711 ; n52711_not
g72922 not n51442 ; n51442_not
g72923 not n11725 ; n11725_not
g72924 not n24604 ; n24604_not
g72925 not n11734 ; n11734_not
g72926 not n11743 ; n11743_not
g72927 not n11752 ; n11752_not
g72928 not n56203 ; n56203_not
g72929 not n51433 ; n51433_not
g72930 not n11761 ; n11761_not
g72931 not n11536 ; n11536_not
g72932 not n11770 ; n11770_not
g72933 not n40507 ; n40507_not
g72934 not n44251 ; n44251_not
g72935 not n51424 ; n51424_not
g72936 not n11662 ; n11662_not
g72937 not n40462 ; n40462_not
g72938 not n11671 ; n11671_not
g72939 not n51460 ; n51460_not
g72940 not n40471 ; n40471_not
g72941 not n11680 ; n11680_not
g72942 not n11581 ; n11581_not
g72943 not n51451 ; n51451_not
g72944 not n44260 ; n44260_not
g72945 not n40480 ; n40480_not
g72946 not n56212 ; n56212_not
g72947 not n11707 ; n11707_not
g72948 not n23722 ; n23722_not
g72949 not n37123 ; n37123_not
g72950 not n12076 ; n12076_not
g72951 not n12067 ; n12067_not
g72952 not n40714 ; n40714_not
g72953 not n55240 ; n55240_not
g72954 not n12058 ; n12058_not
g72955 not n56104 ; n56104_not
g72956 not n51262 ; n51262_not
g72957 not n51271 ; n51271_not
g72958 not n56122 ; n56122_not
g72959 not n52621 ; n52621_not
g72960 not n34720 ; n34720_not
g72961 not n48121 ; n48121_not
g72962 not n23812 ; n23812_not
g72963 not n34711 ; n34711_not
g72964 not n44170 ; n44170_not
g72965 not n29104 ; n29104_not
g72966 not n54403 ; n54403_not
g72967 not n48022 ; n48022_not
g72968 not n51280 ; n51280_not
g72969 not n24433 ; n24433_not
g72970 not n29005 ; n29005_not
g72971 not n12148 ; n12148_not
g72972 not n12157 ; n12157_not
g72973 not n40093 ; n40093_not
g72974 not n29014 ; n29014_not
g72975 not n24523 ; n24523_not
g72976 not n51316 ; n51316_not
g72977 not n51307 ; n51307_not
g72978 not n12085 ; n12085_not
g72979 not n56131 ; n56131_not
g72980 not n40624 ; n40624_not
g72981 not n29041 ; n29041_not
g72982 not n40615 ; n40615_not
g72983 not n40606 ; n40606_not
g72984 not n48130 ; n48130_not
g72985 not n12175 ; n12175_not
g72986 not n29023 ; n29023_not
g72987 not n23632 ; n23632_not
g72988 not n56140 ; n56140_not
g72989 not n12166 ; n12166_not
g72990 not n40633 ; n40633_not
g72991 not n29032 ; n29032_not
g72992 not n19303 ; n19303_not
g72993 not n42037 ; n42037_not
g72994 not n43027 ; n43027_not
g72995 not n31471 ; n31471_not
g72996 not n42334 ; n42334_not
g72997 not n30517 ; n30517_not
g72998 not n16522 ; n16522_not
g72999 not n17800 ; n17800_not
g73000 not n32344 ; n32344_not
g73001 not n18601 ; n18601_not
g73002 not n42154 ; n42154_not
g73003 not n17053 ; n17053_not
g73004 not n31516 ; n31516_not
g73005 not n30526 ; n30526_not
g73006 not n32560 ; n32560_not
g73007 not n18322 ; n18322_not
g73008 not n32065 ; n32065_not
g73009 not n42514 ; n42514_not
g73010 not n54331 ; n54331_not
g73011 not n55213 ; n55213_not
g73012 not n42415 ; n42415_not
g73013 not n42109 ; n42109_not
g73014 not n16360 ; n16360_not
g73015 not n18007 ; n18007_not
g73016 not n31354 ; n31354_not
g73017 not n44710 ; n44710_not
g73018 not n41524 ; n41524_not
g73019 not n31840 ; n31840_not
g73020 not n42208 ; n42208_not
g73021 not n17071 ; n17071_not
g73022 not n17062 ; n17062_not
g73023 not n44620 ; n44620_not
g73024 not n42046 ; n42046_not
g73025 not n30571 ; n30571_not
g73026 not n31372 ; n31372_not
g73027 not n54025 ; n54025_not
g73028 not n16450 ; n16450_not
g73029 not n18700 ; n18700_not
g73030 not n32290 ; n32290_not
g73031 not n18340 ; n18340_not
g73032 not n54205 ; n54205_not
g73033 not n42262 ; n42262_not
g73034 not n31453 ; n31453_not
g73035 not n30580 ; n30580_not
g73036 not n42631 ; n42631_not
g73037 not n38131 ; n38131_not
g73038 not n41515 ; n41515_not
g73039 not n42406 ; n42406_not
g73040 not n45205 ; n45205_not
g73041 not n55204 ; n55204_not
g73042 not n31363 ; n31363_not
g73043 not n50191 ; n50191_not
g73044 not n31651 ; n31651_not
g73045 not n32335 ; n32335_not
g73046 not n41650 ; n41650_not
g73047 not n19024 ; n19024_not
g73048 not n31336 ; n31336_not
g73049 not n18016 ; n18016_not
g73050 not n32362 ; n32362_not
g73051 not n41542 ; n41542_not
g73052 not n54106 ; n54106_not
g73053 not n32515 ; n32515_not
g73054 not n30616 ; n30616_not
g73055 not n19033 ; n19033_not
g73056 not n32038 ; n32038_not
g73057 not n44701 ; n44701_not
g73058 not n42163 ; n42163_not
g73059 not n32524 ; n32524_not
g73060 not n17026 ; n17026_not
g73061 not n43009 ; n43009_not
g73062 not n42424 ; n42424_not
g73063 not n53701 ; n53701_not
g73064 not n31615 ; n31615_not
g73065 not n30805 ; n30805_not
g73066 not n42451 ; n42451_not
g73067 not n31570 ; n31570_not
g73068 not n32074 ; n32074_not
g73069 not n19006 ; n19006_not
g73070 not n42343 ; n42343_not
g73071 not n18115 ; n18115_not
g73072 not n31723 ; n31723_not
g73073 not n31831 ; n31831_not
g73074 not n31183 ; n31183_not
g73075 not n30607 ; n30607_not
g73076 not n30742 ; n30742_not
g73077 not n19042 ; n19042_not
g73078 not n50236 ; n50236_not
g73079 not n17044 ; n17044_not
g73080 not n32632 ; n32632_not
g73081 not n31345 ; n31345_not
g73082 not n19060 ; n19060_not
g73083 not n42253 ; n42253_not
g73084 not n42118 ; n42118_not
g73085 not n31174 ; n31174_not
g73086 not n43018 ; n43018_not
g73087 not n54034 ; n54034_not
g73088 not n41641 ; n41641_not
g73089 not n41533 ; n41533_not
g73090 not n19051 ; n19051_not
g73091 not n32506 ; n32506_not
g73092 not n54214 ; n54214_not
g73093 not n54430 ; n54430_not
g73094 not n42127 ; n42127_not
g73095 not n41920 ; n41920_not
g73096 not n42217 ; n42217_not
g73097 not n17134 ; n17134_not
g73098 not n32434 ; n32434_not
g73099 not n31417 ; n31417_not
g73100 not n54241 ; n54241_not
g73101 not n43054 ; n43054_not
g73102 not n42082 ; n42082_not
g73103 not n54007 ; n54007_not
g73104 not n30562 ; n30562_not
g73105 not n19231 ; n19231_not
g73106 not n47320 ; n47320_not
g73107 not n54340 ; n54340_not
g73108 not n42901 ; n42901_not
g73109 not n31525 ; n31525_not
g73110 not n18304 ; n18304_not
g73111 not n18133 ; n18133_not
g73112 not n31228 ; n31228_not
g73113 not n54223 ; n54223_not
g73114 not n19330 ; n19330_not
g73115 not n32443 ; n32443_not
g73116 not n19222 ; n19222_not
g73117 not n32281 ; n32281_not
g73118 not n54250 ; n54250_not
g73119 not n45232 ; n45232_not
g73120 not n30553 ; n30553_not
g73121 not n31408 ; n31408_not
g73122 not n42370 ; n42370_not
g73123 not n17161 ; n17161_not
g73124 not n31255 ; n31255_not
g73125 not n32416 ; n32416_not
g73126 not n42073 ; n42073_not
g73127 not n32272 ; n32272_not
g73128 not n17143 ; n17143_not
g73129 not n42361 ; n42361_not
g73130 not n32542 ; n32542_not
g73131 not n32425 ; n32425_not
g73132 not n41812 ; n41812_not
g73133 not n31246 ; n31246_not
g73134 not n31606 ; n31606_not
g73135 not n42550 ; n42550_not
g73136 not n32470 ; n32470_not
g73137 not n32056 ; n32056_not
g73138 not n18610 ; n18610_not
g73139 not n32317 ; n32317_not
g73140 not n42271 ; n42271_not
g73141 not n19402 ; n19402_not
g73142 not n41506 ; n41506_not
g73143 not n31381 ; n31381_not
g73144 not n30733 ; n30733_not
g73145 not n42145 ; n42145_not
g73146 not n31390 ; n31390_not
g73147 not n31732 ; n31732_not
g73148 not n41902 ; n41902_not
g73149 not n43036 ; n43036_not
g73150 not n18124 ; n18124_not
g73151 not n42091 ; n42091_not
g73152 not n31435 ; n31435_not
g73153 not n42505 ; n42505_not
g73154 not n17116 ; n17116_not
g73155 not n42541 ; n42541_not
g73156 not n54151 ; n54151_not
g73157 not n42325 ; n42325_not
g73158 not n31219 ; n31219_not
g73159 not n16405 ; n16405_not
g73160 not n19420 ; n19420_not
g73161 not n19321 ; n19321_not
g73162 not n32452 ; n32452_not
g73163 not n43045 ; n43045_not
g73164 not n54016 ; n54016_not
g73165 not n42352 ; n42352_not
g73166 not n31426 ; n31426_not
g73167 not n16432 ; n16432_not
g73168 not n42136 ; n42136_not
g73169 not n32551 ; n32551_not
g73170 not n19411 ; n19411_not
g73171 not n32461 ; n32461_not
g73172 not n42460 ; n42460_not
g73173 not n19312 ; n19312_not
g73174 not n16414 ; n16414_not
g73175 not n18061 ; n18061_not
g73176 not n16540 ; n16540_not
g73177 not n18412 ; n18412_not
g73178 not n31813 ; n31813_not
g73179 not n42820 ; n42820_not
g73180 not n54115 ; n54115_not
g73181 not n19150 ; n19150_not
g73182 not n54304 ; n54304_not
g73183 not n32353 ; n32353_not
g73184 not n32083 ; n32083_not
g73185 not n31642 ; n31642_not
g73186 not n42226 ; n42226_not
g73187 not n31912 ; n31912_not
g73188 not n30841 ; n30841_not
g73189 not n31543 ; n31543_not
g73190 not n31264 ; n31264_not
g73191 not n16531 ; n16531_not
g73192 not n30922 ; n30922_not
g73193 not n41623 ; n41623_not
g73194 not n54061 ; n54061_not
g73195 not n18502 ; n18502_not
g73196 not n30913 ; n30913_not
g73197 not n16504 ; n16504_not
g73198 not n42190 ; n42190_not
g73199 not n30832 ; n30832_not
g73200 not n17017 ; n17017_not
g73201 not n31273 ; n31273_not
g73202 not n19132 ; n19132_not
g73203 not n42811 ; n42811_not
g73204 not n16324 ; n16324_not
g73205 not n42181 ; n42181_not
g73206 not n45151 ; n45151_not
g73207 not n17008 ; n17008_not
g73208 not n42307 ; n42307_not
g73209 not n30760 ; n30760_not
g73210 not n32407 ; n32407_not
g73211 not n42613 ; n42613_not
g73212 not n41614 ; n41614_not
g73213 not n42316 ; n42316_not
g73214 not n31714 ; n31714_not
g73215 not n41830 ; n41830_not
g73216 not n53404 ; n53404_not
g73217 not n18430 ; n18430_not
g73218 not n38023 ; n38023_not
g73219 not n41605 ; n41605_not
g73220 not n54421 ; n54421_not
g73221 not n53800 ; n53800_not
g73222 not n19213 ; n19213_not
g73223 not n31633 ; n31633_not
g73224 not n42172 ; n42172_not
g73225 not n18070 ; n18070_not
g73226 not n30850 ; n30850_not
g73227 not n30715 ; n30715_not
g73228 not n45160 ; n45160_not
g73229 not n31741 ; n31741_not
g73230 not n19240 ; n19240_not
g73231 not n16315 ; n16315_not
g73232 not n31534 ; n31534_not
g73233 not n31921 ; n31921_not
g73234 not n47311 ; n47311_not
g73235 not n30814 ; n30814_not
g73236 not n18034 ; n18034_not
g73237 not n31165 ; n31165_not
g73238 not n54412 ; n54412_not
g73239 not n31318 ; n31318_not
g73240 not n31156 ; n31156_not
g73241 not n18106 ; n18106_not
g73242 not n50146 ; n50146_not
g73243 not n41560 ; n41560_not
g73244 not n54160 ; n54160_not
g73245 not n30643 ; n30643_not
g73246 not n32533 ; n32533_not
g73247 not n41236 ; n41236_not
g73248 not n38140 ; n38140_not
g73249 not n30751 ; n30751_not
g73250 not n53710 ; n53710_not
g73251 not n31822 ; n31822_not
g73252 not n19015 ; n19015_not
g73253 not n41551 ; n41551_not
g73254 not n54043 ; n54043_not
g73255 not n41371 ; n41371_not
g73256 not n18025 ; n18025_not
g73257 not n31903 ; n31903_not
g73258 not n30625 ; n30625_not
g73259 not n31327 ; n31327_not
g73260 not n42640 ; n42640_not
g73261 not n47302 ; n47302_not
g73262 not n31561 ; n31561_not
g73263 not n30634 ; n30634_not
g73264 not n31480 ; n31480_not
g73265 not n31291 ; n31291_not
g73266 not n18052 ; n18052_not
g73267 not n54133 ; n54133_not
g73268 not n30823 ; n30823_not
g73269 not n31552 ; n31552_not
g73270 not n42433 ; n42433_not
g73271 not n30670 ; n30670_not
g73272 not n16333 ; n16333_not
g73273 not n19123 ; n19123_not
g73274 not n42235 ; n42235_not
g73275 not n31282 ; n31282_not
g73276 not n32380 ; n32380_not
g73277 not n18520 ; n18520_not
g73278 not n31930 ; n31930_not
g73279 not n55132 ; n55132_not
g73280 not n31309 ; n31309_not
g73281 not n45214 ; n45214_not
g73282 not n18043 ; n18043_not
g73283 not n42244 ; n42244_not
g73284 not n30652 ; n30652_not
g73285 not n41326 ; n41326_not
g73286 not n30481 ; n30481_not
g73287 not n42802 ; n42802_not
g73288 not n32092 ; n32092_not
g73289 not n54052 ; n54052_not
g73290 not n41632 ; n41632_not
g73291 not n31624 ; n31624_not
g73292 not n30661 ; n30661_not
g73293 not n19105 ; n19105_not
g73294 not n18241 ; n18241_not
g73295 not n42064 ; n42064_not
g73296 not n47221 ; n47221_not
g73297 not n19141 ; n19141_not
g73298 not n45241 ; n45241_not
g73299 not n17710 ; n17710_not
g73300 not n54313 ; n54313_not
g73301 not n44611 ; n44611_not
g73302 not n18232 ; n18232_not
g73303 not n42604 ; n42604_not
g73304 not n42055 ; n42055_not
g73305 not n42280 ; n42280_not
g73306 not n41731 ; n41731_not
g73307 not n42721 ; n42721_not
g73308 not n32722 ; n32722_not
g73309 not n18160 ; n18160_not
g73310 not n31444 ; n31444_not
g73311 not n53602 ; n53602_not
g73312 not n41911 ; n41911_not
g73313 not n30535 ; n30535_not
g73314 not n31237 ; n31237_not
g73315 not n32308 ; n32308_not
g73316 not n32713 ; n32713_not
g73317 not n47131 ; n47131_not
g73318 not n16270 ; n16270_not
g73319 not n42730 ; n42730_not
g73320 not n30706 ; n30706_not
g73321 not n18151 ; n18151_not
g73322 not n42910 ; n42910_not
g73323 not n18250 ; n18250_not
g73324 not n41740 ; n41740_not
g73325 not n53314 ; n53314_not
g73326 not n30904 ; n30904_not
g73327 not n18205 ; n18205_not
g73328 not n41713 ; n41713_not
g73329 not n41281 ; n41281_not
g73330 not n55042 ; n55042_not
g73331 not n32029 ; n32029_not
g73332 not n42028 ; n42028_not
g73333 not n55222 ; n55222_not
g73334 not n45124 ; n45124_not
g73335 not n42703 ; n42703_not
g73336 not n41821 ; n41821_not
g73337 not n31660 ; n31660_not
g73338 not n31192 ; n31192_not
g73339 not n17152 ; n17152_not
g73340 not n18223 ; n18223_not
g73341 not n38113 ; n38113_not
g73342 not n17107 ; n17107_not
g73343 not n41722 ; n41722_not
g73344 not n41704 ; n41704_not
g73345 not n16423 ; n16423_not
g73346 not n18214 ; n18214_not
g73347 not n42712 ; n42712_not
g73348 not n30931 ; n30931_not
g73349 not n15640 ; n15640_not
g73350 not n54124 ; n54124_not
g73351 not n18403 ; n18403_not
g73352 not n16342 ; n16342_not
g73353 not n42523 ; n42523_not
g73354 not n53620 ; n53620_not
g73355 not n53611 ; n53611_not
g73356 not n18142 ; n18142_not
g73357 not n52406 ; n52406_not
g73358 not n13364 ; n13364_not
g73359 not n51029 ; n51029_not
g73360 not n21608 ; n21608_not
g73361 not n56114 ; n56114_not
g73362 not n38024 ; n38024_not
g73363 not n21626 ; n21626_not
g73364 not n22562 ; n22562_not
g73365 not n25802 ; n25802_not
g73366 not n40850 ; n40850_not
g73367 not n50093 ; n50093_not
g73368 not n50471 ; n50471_not
g73369 not n50336 ; n50336_not
g73370 not n44315 ; n44315_not
g73371 not n22256 ; n22256_not
g73372 not n52280 ; n52280_not
g73373 not n21617 ; n21617_not
g73374 not n25370 ; n25370_not
g73375 not n44324 ; n44324_not
g73376 not n10817 ; n10817_not
g73377 not n37214 ; n37214_not
g73378 not n22553 ; n22553_not
g73379 not n32345 ; n32345_not
g73380 not n22247 ; n22247_not
g73381 not n13346 ; n13346_not
g73382 not n52127 ; n52127_not
g73383 not n22544 ; n22544_not
g73384 not n42308 ; n42308_not
g73385 not n22526 ; n22526_not
g73386 not n35315 ; n35315_not
g73387 not n50057 ; n50057_not
g73388 not n53144 ; n53144_not
g73389 not n13328 ; n13328_not
g73390 not n34181 ; n34181_not
g73391 not n13724 ; n13724_not
g73392 not n10457 ; n10457_not
g73393 not n50651 ; n50651_not
g73394 not n50039 ; n50039_not
g73395 not n21644 ; n21644_not
g73396 not n42245 ; n42245_not
g73397 not n34037 ; n34037_not
g73398 not n52118 ; n52118_not
g73399 not n50714 ; n50714_not
g73400 not n10691 ; n10691_not
g73401 not n13373 ; n13373_not
g73402 not n22490 ; n22490_not
g73403 not n13742 ; n13742_not
g73404 not n54062 ; n54062_not
g73405 not n52415 ; n52415_not
g73406 not n50804 ; n50804_not
g73407 not n49310 ; n49310_not
g73408 not n38015 ; n38015_not
g73409 not n25505 ; n25505_not
g73410 not n22472 ; n22472_not
g73411 not n22535 ; n22535_not
g73412 not n10808 ; n10808_not
g73413 not n34352 ; n34352_not
g73414 not n40238 ; n40238_not
g73415 not n18404 ; n18404_not
g73416 not n10907 ; n10907_not
g73417 not n42254 ; n42254_not
g73418 not n50462 ; n50462_not
g73419 not n52433 ; n52433_not
g73420 not n22517 ; n22517_not
g73421 not n32453 ; n32453_not
g73422 not n37061 ; n37061_not
g73423 not n31058 ; n31058_not
g73424 not n13940 ; n13940_not
g73425 not n13337 ; n13337_not
g73426 not n47213 ; n47213_not
g73427 not n28421 ; n28421_not
g73428 not n21635 ; n21635_not
g73429 not n22508 ; n22508_not
g73430 not n16712 ; n16712_not
g73431 not n10466 ; n10466_not
g73432 not n31517 ; n31517_not
g73433 not n10790 ; n10790_not
g73434 not n41921 ; n41921_not
g73435 not n21563 ; n21563_not
g73436 not n31436 ; n31436_not
g73437 not n16343 ; n16343_not
g73438 not n35333 ; n35333_not
g73439 not n50822 ; n50822_not
g73440 not n34154 ; n34154_not
g73441 not n22652 ; n22652_not
g73442 not n42902 ; n42902_not
g73443 not n34190 ; n34190_not
g73444 not n53153 ; n53153_not
g73445 not n13391 ; n13391_not
g73446 not n22643 ; n22643_not
g73447 not n32318 ; n32318_not
g73448 not n10880 ; n10880_not
g73449 not n22463 ; n22463_not
g73450 not n21572 ; n21572_not
g73451 not n52154 ; n52154_not
g73452 not n42155 ; n42155_not
g73453 not n22634 ; n22634_not
g73454 not n42038 ; n42038_not
g73455 not n35306 ; n35306_not
g73456 not n16721 ; n16721_not
g73457 not n52163 ; n52163_not
g73458 not n28403 ; n28403_not
g73459 not n50516 ; n50516_not
g73460 not n10709 ; n10709_not
g73461 not n30860 ; n30860_not
g73462 not n30770 ; n30770_not
g73463 not n13418 ; n13418_not
g73464 not n34334 ; n34334_not
g73465 not n38222 ; n38222_not
g73466 not n35441 ; n35441_not
g73467 not n54008 ; n54008_not
g73468 not n21554 ; n21554_not
g73469 not n32390 ; n32390_not
g73470 not n44027 ; n44027_not
g73471 not n50048 ; n50048_not
g73472 not n50507 ; n50507_not
g73473 not n13409 ; n13409_not
g73474 not n22670 ; n22670_not
g73475 not n52271 ; n52271_not
g73476 not n25604 ; n25604_not
g73477 not n36413 ; n36413_not
g73478 not n45305 ; n45305_not
g73479 not n42236 ; n42236_not
g73480 not n16820 ; n16820_not
g73481 not n22661 ; n22661_not
g73482 not n22166 ; n22166_not
g73483 not n10844 ; n10844_not
g73484 not n43280 ; n43280_not
g73485 not n16334 ; n16334_not
g73486 not n50480 ; n50480_not
g73487 not n36422 ; n36422_not
g73488 not n52145 ; n52145_not
g73489 not n53306 ; n53306_not
g73490 not n34343 ; n34343_not
g73491 not n13733 ; n13733_not
g73492 not n50813 ; n50813_not
g73493 not n40742 ; n40742_not
g73494 not n42146 ; n42146_not
g73495 not n38330 ; n38330_not
g73496 not n10826 ; n10826_not
g73497 not n10655 ; n10655_not
g73498 not n10484 ; n10484_not
g73499 not n22580 ; n22580_not
g73500 not n44036 ; n44036_not
g73501 not n22931 ; n22931_not
g73502 not n54260 ; n54260_not
g73503 not n22571 ; n22571_not
g73504 not n52136 ; n52136_not
g73505 not n35450 ; n35450_not
g73506 not n22175 ; n22175_not
g73507 not n31049 ; n31049_not
g73508 not n50741 ; n50741_not
g73509 not n42524 ; n42524_not
g73510 not n38321 ; n38321_not
g73511 not n32462 ; n32462_not
g73512 not n22625 ; n22625_not
g73513 not n22274 ; n22274_not
g73514 not n10835 ; n10835_not
g73515 not n45026 ; n45026_not
g73516 not n21581 ; n21581_not
g73517 not n22904 ; n22904_not
g73518 not n25271 ; n25271_not
g73519 not n52442 ; n52442_not
g73520 not n22616 ; n22616_not
g73521 not n13382 ; n13382_not
g73522 not n32048 ; n32048_not
g73523 not n21590 ; n21590_not
g73524 not n54053 ; n54053_not
g73525 not n18215 ; n18215_not
g73526 not n41912 ; n41912_not
g73527 not n22913 ; n22913_not
g73528 not n22607 ; n22607_not
g73529 not n34055 ; n34055_not
g73530 not n41723 ; n41723_not
g73531 not n46115 ; n46115_not
g73532 not n13238 ; n13238_not
g73533 not n10727 ; n10727_not
g73534 not n51056 ; n51056_not
g73535 not n46052 ; n46052_not
g73536 not n54116 ; n54116_not
g73537 not n21734 ; n21734_not
g73538 not n42137 ; n42137_not
g73539 not n52505 ; n52505_not
g73540 not n43910 ; n43910_not
g73541 not n10718 ; n10718_not
g73542 not n10952 ; n10952_not
g73543 not n14048 ; n14048_not
g73544 not n50723 ; n50723_not
g73545 not n22184 ; n22184_not
g73546 not n23084 ; n23084_not
g73547 not n13445 ; n13445_not
g73548 not n32354 ; n32354_not
g73549 not n44072 ; n44072_not
g73550 not n21743 ; n21743_not
g73551 not n40751 ; n40751_not
g73552 not n26018 ; n26018_not
g73553 not n18422 ; n18422_not
g73554 not n10394 ; n10394_not
g73555 not n10736 ; n10736_not
g73556 not n22346 ; n22346_not
g73557 not n19250 ; n19250_not
g73558 not n36602 ; n36602_not
g73559 not n38033 ; n38033_not
g73560 not n25820 ; n25820_not
g73561 not n37205 ; n37205_not
g73562 not n22337 ; n22337_not
g73563 not n44063 ; n44063_not
g73564 not n36431 ; n36431_not
g73565 not n23066 ; n23066_not
g73566 not n50426 ; n50426_not
g73567 not n22328 ; n22328_not
g73568 not n41822 ; n41822_not
g73569 not n13247 ; n13247_not
g73570 not n21725 ; n21725_not
g73571 not n14039 ; n14039_not
g73572 not n13436 ; n13436_not
g73573 not n22319 ; n22319_not
g73574 not n46124 ; n46124_not
g73575 not n45206 ; n45206_not
g73576 not n41750 ; n41750_not
g73577 not n31841 ; n31841_not
g73578 not n50408 ; n50408_not
g73579 not n52082 ; n52082_not
g73580 not n34163 ; n34163_not
g73581 not n22481 ; n22481_not
g73582 not n10376 ; n10376_not
g73583 not n42326 ; n42326_not
g73584 not n13175 ; n13175_not
g73585 not n21770 ; n21770_not
g73586 not n35270 ; n35270_not
g73587 not n56006 ; n56006_not
g73588 not n42128 ; n42128_not
g73589 not n48041 ; n48041_not
g73590 not n10682 ; n10682_not
g73591 not n50732 ; n50732_not
g73592 not n32516 ; n32516_not
g73593 not n53207 ; n53207_not
g73594 not n31085 ; n31085_not
g73595 not n38213 ; n38213_not
g73596 not n47312 ; n47312_not
g73597 not n50417 ; n50417_not
g73598 not n31850 ; n31850_not
g73599 not n37250 ; n37250_not
g73600 not n21752 ; n21752_not
g73601 not n50561 ; n50561_not
g73602 not n38060 ; n38060_not
g73603 not n10673 ; n10673_not
g73604 not n19232 ; n19232_not
g73605 not n52091 ; n52091_not
g73606 not n47132 ; n47132_not
g73607 not n14057 ; n14057_not
g73608 not n32435 ; n32435_not
g73609 not n13193 ; n13193_not
g73610 not n21761 ; n21761_not
g73611 not n13454 ; n13454_not
g73612 not n54080 ; n54080_not
g73613 not n41714 ; n41714_not
g73614 not n19223 ; n19223_not
g73615 not n34406 ; n34406_not
g73616 not n52613 ; n52613_not
g73617 not n31094 ; n31094_not
g73618 not n35405 ; n35405_not
g73619 not n22454 ; n22454_not
g73620 not n41273 ; n41273_not
g73621 not n34361 ; n34361_not
g73622 not n53135 ; n53135_not
g73623 not n40229 ; n40229_not
g73624 not n22445 ; n22445_not
g73625 not n21680 ; n21680_not
g73626 not n49301 ; n49301_not
g73627 not n10439 ; n10439_not
g73628 not n10772 ; n10772_not
g73629 not n22436 ; n22436_not
g73630 not n25541 ; n25541_not
g73631 not n50444 ; n50444_not
g73632 not n31067 ; n31067_not
g73633 not n22427 ; n22427_not
g73634 not n13292 ; n13292_not
g73635 not n48410 ; n48410_not
g73636 not n44054 ; n44054_not
g73637 not n49400 ; n49400_not
g73638 not n22418 ; n22418_not
g73639 not n25532 ; n25532_not
g73640 not n21653 ; n21653_not
g73641 not n31490 ; n31490_not
g73642 not n34028 ; n34028_not
g73643 not n51038 ; n51038_not
g73644 not n50453 ; n50453_not
g73645 not n22229 ; n22229_not
g73646 not n21662 ; n21662_not
g73647 not n13931 ; n13931_not
g73648 not n18206 ; n18206_not
g73649 not n10781 ; n10781_not
g73650 not n46106 ; n46106_not
g73651 not n28322 ; n28322_not
g73652 not n16325 ; n16325_not
g73653 not n21671 ; n21671_not
g73654 not n30923 ; n30923_not
g73655 not n50066 ; n50066_not
g73656 not n44045 ; n44045_not
g73657 not n25550 ; n25550_not
g73658 not n31931 ; n31931_not
g73659 not n25514 ; n25514_not
g73660 not n22382 ; n22382_not
g73661 not n21707 ; n21707_not
g73662 not n52109 ; n52109_not
g73663 not n13427 ; n13427_not
g73664 not n31940 ; n31940_not
g73665 not n24704 ; n24704_not
g73666 not n30914 ; n30914_not
g73667 not n23039 ; n23039_not
g73668 not n26009 ; n26009_not
g73669 not n22373 ; n22373_not
g73670 not n31076 ; n31076_not
g73671 not n28304 ; n28304_not
g73672 not n13265 ; n13265_not
g73673 not n16703 ; n16703_not
g73674 not n50435 ; n50435_not
g73675 not n23048 ; n23048_not
g73676 not n21716 ; n21716_not
g73677 not n25361 ; n25361_not
g73678 not n22364 ; n22364_not
g73679 not n54071 ; n54071_not
g73680 not n51605 ; n51605_not
g73681 not n22355 ; n22355_not
g73682 not n34172 ; n34172_not
g73683 not n10763 ; n10763_not
g73684 not n13922 ; n13922_not
g73685 not n13283 ; n13283_not
g73686 not n13751 ; n13751_not
g73687 not n42317 ; n42317_not
g73688 not n22409 ; n22409_not
g73689 not n10925 ; n10925_not
g73690 not n34370 ; n34370_not
g73691 not n25811 ; n25811_not
g73692 not n10664 ; n10664_not
g73693 not n10754 ; n10754_not
g73694 not n32444 ; n32444_not
g73695 not n36800 ; n36800_not
g73696 not n22391 ; n22391_not
g73697 not n10934 ; n10934_not
g73698 not n10745 ; n10745_not
g73699 not n13661 ; n13661_not
g73700 not n13562 ; n13562_not
g73701 not n16730 ; n16730_not
g73702 not n42272 ; n42272_not
g73703 not n28340 ; n28340_not
g73704 not n50138 ; n50138_not
g73705 not n34271 ; n34271_not
g73706 not n22706 ; n22706_not
g73707 not n31454 ; n31454_not
g73708 not n53180 ; n53180_not
g73709 not n46034 ; n46034_not
g73710 not n34217 ; n34217_not
g73711 not n47150 ; n47150_not
g73712 not n47006 ; n47006_not
g73713 not n52208 ; n52208_not
g73714 not n42281 ; n42281_not
g73715 not n34046 ; n34046_not
g73716 not n52343 ; n52343_not
g73717 not n13553 ; n13553_not
g73718 not n44351 ; n44351_not
g73719 not n52550 ; n52550_not
g73720 not n22715 ; n22715_not
g73721 not n30815 ; n30815_not
g73722 not n25703 ; n25703_not
g73723 not n34262 ; n34262_not
g73724 not n10475 ; n10475_not
g73725 not n48401 ; n48401_not
g73726 not n31445 ; n31445_not
g73727 not n52334 ; n52334_not
g73728 not n40715 ; n40715_not
g73729 not n50633 ; n50633_not
g73730 not n41741 ; n41741_not
g73731 not n35414 ; n35414_not
g73732 not n13571 ; n13571_not
g73733 not n22085 ; n22085_not
g73734 not n52217 ; n52217_not
g73735 not n54026 ; n54026_not
g73736 not n18251 ; n18251_not
g73737 not n34127 ; n34127_not
g73738 not n50750 ; n50750_not
g73739 not n31904 ; n31904_not
g73740 not n40274 ; n40274_not
g73741 not n22076 ; n22076_not
g73742 not n46070 ; n46070_not
g73743 not n10367 ; n10367_not
g73744 not n37223 ; n37223_not
g73745 not n42209 ; n42209_not
g73746 not n56303 ; n56303_not
g73747 not n22733 ; n22733_not
g73748 not n18350 ; n18350_not
g73749 not n17630 ; n17630_not
g73750 not n42218 ; n42218_not
g73751 not n41075 ; n41075_not
g73752 not n13535 ; n13535_not
g73753 not n52523 ; n52523_not
g73754 not n42182 ; n42182_not
g73755 not n41246 ; n41246_not
g73756 not n32480 ; n32480_not
g73757 not n10592 ; n10592_not
g73758 not n22742 ; n22742_not
g73759 not n52190 ; n52190_not
g73760 not n30824 ; n30824_not
g73761 not n50615 ; n50615_not
g73762 not n10637 ; n10637_not
g73763 not n25316 ; n25316_not
g73764 not n50624 ; n50624_not
g73765 not n38240 ; n38240_not
g73766 not n22067 ; n22067_not
g73767 not n50543 ; n50543_not
g73768 not n34280 ; n34280_not
g73769 not n35360 ; n35360_not
g73770 not n25901 ; n25901_not
g73771 not n34118 ; n34118_not
g73772 not n50075 ; n50075_not
g73773 not n51623 ; n51623_not
g73774 not n22724 ; n22724_not
g73775 not n13544 ; n13544_not
g73776 not n45215 ; n45215_not
g73777 not n17612 ; n17612_not
g73778 not n52244 ; n52244_not
g73779 not n13670 ; n13670_not
g73780 not n54017 ; n54017_not
g73781 not n41093 ; n41093_not
g73782 not n13814 ; n13814_not
g73783 not n17702 ; n17702_not
g73784 not n30806 ; n30806_not
g73785 not n46043 ; n46043_not
g73786 not n50921 ; n50921_not
g73787 not n40247 ; n40247_not
g73788 not n34136 ; n34136_not
g73789 not n38051 ; n38051_not
g73790 not n44333 ; n44333_not
g73791 not n10619 ; n10619_not
g73792 not n13616 ; n13616_not
g73793 not n34226 ; n34226_not
g73794 not n51632 ; n51632_not
g73795 not n42506 ; n42506_not
g73796 not n34244 ; n34244_not
g73797 not n25730 ; n25730_not
g73798 not n40175 ; n40175_not
g73799 not n46061 ; n46061_not
g73800 not n13643 ; n13643_not
g73801 not n43901 ; n43901_not
g73802 not n31913 ; n31913_not
g73803 not n10628 ; n10628_not
g73804 not n19241 ; n19241_not
g73805 not n34235 ; n34235_not
g73806 not n13634 ; n13634_not
g73807 not n45620 ; n45620_not
g73808 not n18323 ; n18323_not
g73809 not n37232 ; n37232_not
g73810 not n52316 ; n52316_not
g73811 not n32507 ; n32507_not
g73812 not n25334 ; n25334_not
g73813 not n52226 ; n52226_not
g73814 not n31922 ; n31922_not
g73815 not n25406 ; n25406_not
g73816 not n13625 ; n13625_not
g73817 not n25415 ; n25415_not
g73818 not n40706 ; n40706_not
g73819 not n34253 ; n34253_not
g73820 not n25712 ; n25712_not
g73821 not n18314 ; n18314_not
g73822 not n25424 ; n25424_not
g73823 not n50642 ; n50642_not
g73824 not n41084 ; n41084_not
g73825 not n13841 ; n13841_not
g73826 not n10385 ; n10385_not
g73827 not n47330 ; n47330_not
g73828 not n13580 ; n13580_not
g73829 not n40265 ; n40265_not
g73830 not n47420 ; n47420_not
g73831 not n42191 ; n42191_not
g73832 not n45611 ; n45611_not
g73833 not n34073 ; n34073_not
g73834 not n55205 ; n55205_not
g73835 not n13607 ; n13607_not
g73836 not n18260 ; n18260_not
g73837 not n52325 ; n52325_not
g73838 not n50660 ; n50660_not
g73839 not n52235 ; n52235_not
g73840 not n16370 ; n16370_not
g73841 not n42290 ; n42290_not
g73842 not n53270 ; n53270_not
g73843 not n13832 ; n13832_not
g73844 not n13652 ; n13652_not
g73845 not n18332 ; n18332_not
g73846 not n25325 ; n25325_not
g73847 not n52532 ; n52532_not
g73848 not n25721 ; n25721_not
g73849 not n42551 ; n42551_not
g73850 not n34091 ; n34091_not
g73851 not n42533 ; n42533_not
g73852 not n22823 ; n22823_not
g73853 not n16811 ; n16811_not
g73854 not n41048 ; n41048_not
g73855 not n35351 ; n35351_not
g73856 not n47303 ; n47303_not
g73857 not n50552 ; n50552_not
g73858 not n54044 ; n54044_not
g73859 not n22760 ; n22760_not
g73860 not n42173 ; n42173_not
g73861 not n52460 ; n52460_not
g73862 not n42515 ; n42515_not
g73863 not n30941 ; n30941_not
g73864 not n42227 ; n42227_not
g73865 not n34082 ; n34082_not
g73866 not n38312 ; n38312_not
g73867 not n45710 ; n45710_not
g73868 not n30851 ; n30851_not
g73869 not n22751 ; n22751_not
g73870 not n25640 ; n25640_not
g73871 not n25460 ; n25460_not
g73872 not n40139 ; n40139_not
g73873 not n52172 ; n52172_not
g73874 not n52262 ; n52262_not
g73875 not n18233 ; n18233_not
g73876 not n45035 ; n45035_not
g73877 not n13148 ; n13148_not
g73878 not n46016 ; n46016_not
g73879 not n22814 ; n22814_not
g73880 not n25631 ; n25631_not
g73881 not n10556 ; n10556_not
g73882 not n50570 ; n50570_not
g73883 not n31481 ; n31481_not
g73884 not n10853 ; n10853_not
g73885 not n38231 ; n38231_not
g73886 not n34325 ; n34325_not
g73887 not n42263 ; n42263_not
g73888 not n17720 ; n17720_not
g73889 not n50525 ; n50525_not
g73890 not n25613 ; n25613_not
g73891 not n53162 ; n53162_not
g73892 not n41129 ; n41129_not
g73893 not n56312 ; n56312_not
g73894 not n37241 ; n37241_not
g73895 not n42164 ; n42164_not
g73896 not n25280 ; n25280_not
g73897 not n10538 ; n10538_not
g73898 not n47411 ; n47411_not
g73899 not n18224 ; n18224_not
g73900 not n22292 ; n22292_not
g73901 not n35342 ; n35342_not
g73902 not n50831 ; n50831_not
g73903 not n10646 ; n10646_not
g73904 not n51650 ; n51650_not
g73905 not n21545 ; n21545_not
g73906 not n41039 ; n41039_not
g73907 not n25622 ; n25622_not
g73908 not n44018 ; n44018_not
g73909 not n22841 ; n22841_not
g73910 not n50705 ; n50705_not
g73911 not n52370 ; n52370_not
g73912 not n13715 ; n13715_not
g73913 not n28250 ; n28250_not
g73914 not n50534 ; n50534_not
g73915 not n32471 ; n32471_not
g73916 not n10871 ; n10871_not
g73917 not n10547 ; n10547_not
g73918 not n50606 ; n50606_not
g73919 not n40157 ; n40157_not
g73920 not n55214 ; n55214_not
g73921 not n45017 ; n45017_not
g73922 not n41903 ; n41903_not
g73923 not n10583 ; n10583_not
g73924 not n30833 ; n30833_not
g73925 not n41066 ; n41066_not
g73926 not n18242 ; n18242_not
g73927 not n53216 ; n53216_not
g73928 not n51614 ; n51614_not
g73929 not n52307 ; n52307_not
g73930 not n52181 ; n52181_not
g73931 not n54035 ; n54035_not
g73932 not n13490 ; n13490_not
g73933 not n27800 ; n27800_not
g73934 not n13526 ; n13526_not
g73935 not n34208 ; n34208_not
g73936 not n13256 ; n13256_not
g73937 not n42911 ; n42911_not
g73938 not n13517 ; n13517_not
g73939 not n25910 ; n25910_not
g73940 not n22265 ; n22265_not
g73941 not n35423 ; n35423_not
g73942 not n46025 ; n46025_not
g73943 not n17603 ; n17603_not
g73944 not n13166 ; n13166_not
g73945 not n42560 ; n42560_not
g73946 not n36404 ; n36404_not
g73947 not n52253 ; n52253_not
g73948 not n52451 ; n52451_not
g73949 not n13508 ; n13508_not
g73950 not n37070 ; n37070_not
g73951 not n34316 ; n34316_not
g73952 not n28331 ; n28331_not
g73953 not n45602 ; n45602_not
g73954 not n40184 ; n40184_not
g73955 not n53171 ; n53171_not
g73956 not n41057 ; n41057_not
g73957 not n38303 ; n38303_not
g73958 not n13463 ; n13463_not
g73959 not n10565 ; n10565_not
g73960 not n13706 ; n13706_not
g73961 not n30842 ; n30842_not
g73962 not n52361 ; n52361_not
g73963 not n53261 ; n53261_not
g73964 not n22805 ; n22805_not
g73965 not n41732 ; n41732_not
g73966 not n45701 ; n45701_not
g73967 not n22157 ; n22157_not
g73968 not n34307 ; n34307_not
g73969 not n25451 ; n25451_not
g73970 not n41237 ; n41237_not
g73971 not n50903 ; n50903_not
g73972 not n13157 ; n13157_not
g73973 not n13481 ; n13481_not
g73974 not n38510 ; n38510_not
g73975 not n52352 ; n52352_not
g73976 not n18305 ; n18305_not
g73977 not n10574 ; n10574_not
g73978 not n16802 ; n16802_not
g73979 not n47600 ; n47600_not
g73980 not n44009 ; n44009_not
g73981 not n13472 ; n13472_not
g73982 not n13904 ; n13904_not
g73983 not n35432 ; n35432_not
g73984 not n11744 ; n11744_not
g73985 not n24074 ; n24074_not
g73986 not n24605 ; n24605_not
g73987 not n11618 ; n11618_not
g73988 not n52703 ; n52703_not
g73989 not n56204 ; n56204_not
g73990 not n31247 ; n31247_not
g73991 not n24065 ; n24065_not
g73992 not n32273 ; n32273_not
g73993 not n11924 ; n11924_not
g73994 not n11735 ; n11735_not
g73995 not n29123 ; n29123_not
g73996 not n45242 ; n45242_not
g73997 not n46412 ; n46412_not
g73998 not n11537 ; n11537_not
g73999 not n29114 ; n29114_not
g74000 not n11753 ; n11753_not
g74001 not n24092 ; n24092_not
g74002 not n44180 ; n44180_not
g74003 not n42740 ; n42740_not
g74004 not n51434 ; n51434_not
g74005 not n17171 ; n17171_not
g74006 not n11906 ; n11906_not
g74007 not n32264 ; n32264_not
g74008 not n24614 ; n24614_not
g74009 not n24083 ; n24083_not
g74010 not n47402 ; n47402_not
g74011 not n31256 ; n31256_not
g74012 not n11546 ; n11546_not
g74013 not n11915 ; n11915_not
g74014 not n44171 ; n44171_not
g74015 not n11951 ; n11951_not
g74016 not n24029 ; n24029_not
g74017 not n17153 ; n17153_not
g74018 not n32282 ; n32282_not
g74019 not n11960 ; n11960_not
g74020 not n48032 ; n48032_not
g74021 not n23813 ; n23813_not
g74022 not n29132 ; n29132_not
g74023 not n44423 ; n44423_not
g74024 not n32147 ; n32147_not
g74025 not n52721 ; n52721_not
g74026 not n56051 ; n56051_not
g74027 not n11708 ; n11708_not
g74028 not n23822 ; n23822_not
g74029 not n16604 ; n16604_not
g74030 not n24056 ; n24056_not
g74031 not n11933 ; n11933_not
g74032 not n48122 ; n48122_not
g74033 not n11726 ; n11726_not
g74034 not n18530 ; n18530_not
g74035 not n24047 ; n24047_not
g74036 not n11942 ; n11942_not
g74037 not n23804 ; n23804_not
g74038 not n54251 ; n54251_not
g74039 not n52730 ; n52730_not
g74040 not n46322 ; n46322_not
g74041 not n45080 ; n45080_not
g74042 not n24038 ; n24038_not
g74043 not n11717 ; n11717_not
g74044 not n51443 ; n51443_not
g74045 not n36710 ; n36710_not
g74046 not n47510 ; n47510_not
g74047 not n56105 ; n56105_not
g74048 not n24155 ; n24155_not
g74049 not n29006 ; n29006_not
g74050 not n11834 ; n11834_not
g74051 not n18413 ; n18413_not
g74052 not n24146 ; n24146_not
g74053 not n42074 ; n42074_not
g74054 not n45350 ; n45350_not
g74055 not n11843 ; n11843_not
g74056 not n51263 ; n51263_not
g74057 not n11780 ; n11780_not
g74058 not n11816 ; n11816_not
g74059 not n17360 ; n17360_not
g74060 not n31229 ; n31229_not
g74061 not n23732 ; n23732_not
g74062 not n24641 ; n24641_not
g74063 not n11807 ; n11807_not
g74064 not n24173 ; n24173_not
g74065 not n46403 ; n46403_not
g74066 not n32246 ; n32246_not
g74067 not n11825 ; n11825_not
g74068 not n51416 ; n51416_not
g74069 not n44243 ; n44243_not
g74070 not n29042 ; n29042_not
g74071 not n12068 ; n12068_not
g74072 not n24164 ; n24164_not
g74073 not n52910 ; n52910_not
g74074 not n24119 ; n24119_not
g74075 not n44252 ; n44252_not
g74076 not n16550 ; n16550_not
g74077 not n37133 ; n37133_not
g74078 not n55241 ; n55241_not
g74079 not n31238 ; n31238_not
g74080 not n54350 ; n54350_not
g74081 not n11762 ; n11762_not
g74082 not n36701 ; n36701_not
g74083 not n40148 ; n40148_not
g74084 not n40724 ; n40724_not
g74085 not n24137 ; n24137_not
g74086 not n55070 ; n55070_not
g74087 not n36512 ; n36512_not
g74088 not n51425 ; n51425_not
g74089 not n11852 ; n11852_not
g74090 not n28160 ; n28160_not
g74091 not n24128 ; n24128_not
g74092 not n11528 ; n11528_not
g74093 not n32156 ; n32156_not
g74094 not n11861 ; n11861_not
g74095 not n11771 ; n11771_not
g74096 not n32255 ; n32255_not
g74097 not n11870 ; n11870_not
g74098 not n23912 ; n23912_not
g74099 not n12437 ; n12437_not
g74100 not n45260 ; n45260_not
g74101 not n54206 ; n54206_not
g74102 not n12428 ; n12428_not
g74103 not n23903 ; n23903_not
g74104 not n53027 ; n53027_not
g74105 not n45071 ; n45071_not
g74106 not n11654 ; n11654_not
g74107 not n12419 ; n12419_not
g74108 not n40841 ; n40841_not
g74109 not n54215 ; n54215_not
g74110 not n51254 ; n51254_not
g74111 not n53018 ; n53018_not
g74112 not n36503 ; n36503_not
g74113 not n12455 ; n12455_not
g74114 not n11663 ; n11663_not
g74115 not n23921 ; n23921_not
g74116 not n54341 ; n54341_not
g74117 not n24551 ; n24551_not
g74118 not n40832 ; n40832_not
g74119 not n12446 ; n12446_not
g74120 not n12608 ; n12608_not
g74121 not n51920 ; n51920_not
g74122 not n11645 ; n11645_not
g74123 not n12374 ; n12374_not
g74124 not n12644 ; n12644_not
g74125 not n51470 ; n51470_not
g74126 not n12365 ; n12365_not
g74127 not n12653 ; n12653_not
g74128 not n46250 ; n46250_not
g74129 not n44270 ; n44270_not
g74130 not n12356 ; n12356_not
g74131 not n17072 ; n17072_not
g74132 not n12626 ; n12626_not
g74133 not n37151 ; n37151_not
g74134 not n32309 ; n32309_not
g74135 not n32228 ; n32228_not
g74136 not n17108 ; n17108_not
g74137 not n12392 ; n12392_not
g74138 not n17405 ; n17405_not
g74139 not n32219 ; n32219_not
g74140 not n12383 ; n12383_not
g74141 not n46331 ; n46331_not
g74142 not n52541 ; n52541_not
g74143 not n34424 ; n34424_not
g74144 not n53036 ; n53036_not
g74145 not n45521 ; n45521_not
g74146 not n16622 ; n16622_not
g74147 not n11690 ; n11690_not
g74148 not n56213 ; n56213_not
g74149 not n51452 ; n51452_not
g74150 not n55007 ; n55007_not
g74151 not n12554 ; n12554_not
g74152 not n44261 ; n44261_not
g74153 not n12527 ; n12527_not
g74154 not n12563 ; n12563_not
g74155 not n16631 ; n16631_not
g74156 not n12518 ; n12518_not
g74157 not n11681 ; n11681_not
g74158 not n41930 ; n41930_not
g74159 not n17144 ; n17144_not
g74160 not n44162 ; n44162_not
g74161 not n42065 ; n42065_not
g74162 not n31418 ; n31418_not
g74163 not n16613 ; n16613_not
g74164 not n12545 ; n12545_not
g74165 not n29141 ; n29141_not
g74166 not n47033 ; n47033_not
g74167 not n54233 ; n54233_not
g74168 not n11573 ; n11573_not
g74169 not n53009 ; n53009_not
g74170 not n12482 ; n12482_not
g74171 not n17126 ; n17126_not
g74172 not n24560 ; n24560_not
g74173 not n32138 ; n32138_not
g74174 not n12473 ; n12473_not
g74175 not n51461 ; n51461_not
g74176 not n12464 ; n12464_not
g74177 not n32237 ; n32237_not
g74178 not n11591 ; n11591_not
g74179 not n34415 ; n34415_not
g74180 not n52712 ; n52712_not
g74181 not n44153 ; n44153_not
g74182 not n23930 ; n23930_not
g74183 not n12509 ; n12509_not
g74184 not n45332 ; n45332_not
g74185 not n29150 ; n29150_not
g74186 not n46421 ; n46421_not
g74187 not n12491 ; n12491_not
g74188 not n12581 ; n12581_not
g74189 not n16640 ; n16640_not
g74190 not n40814 ; n40814_not
g74191 not n11582 ; n11582_not
g74192 not n11672 ; n11672_not
g74193 not n56042 ; n56042_not
g74194 not n24416 ; n24416_not
g74195 not n17117 ; n17117_not
g74196 not n17324 ; n17324_not
g74197 not n12158 ; n12158_not
g74198 not n17270 ; n17270_not
g74199 not n52820 ; n52820_not
g74200 not n24407 ; n24407_not
g74201 not n50156 ; n50156_not
g74202 not n12167 ; n12167_not
g74203 not n31184 ; n31184_not
g74204 not n42605 ; n42605_not
g74205 not n51362 ; n51362_not
g74206 not n24353 ; n24353_not
g74207 not n51281 ; n51281_not
g74208 not n24362 ; n24362_not
g74209 not n51353 ; n51353_not
g74210 not n24371 ; n24371_not
g74211 not n24623 ; n24623_not
g74212 not n56141 ; n56141_not
g74213 not n24380 ; n24380_not
g74214 not n24425 ; n24425_not
g74215 not n32183 ; n32183_not
g74216 not n55034 ; n55034_not
g74217 not n34802 ; n34802_not
g74218 not n42713 ; n42713_not
g74219 not n17333 ; n17333_not
g74220 not n29015 ; n29015_not
g74221 not n29024 ; n29024_not
g74222 not n11438 ; n11438_not
g74223 not n23624 ; n23624_not
g74224 not n51371 ; n51371_not
g74225 not n17261 ; n17261_not
g74226 not n11627 ; n11627_not
g74227 not n44216 ; n44216_not
g74228 not n23606 ; n23606_not
g74229 not n24650 ; n24650_not
g74230 not n37043 ; n37043_not
g74231 not n11636 ; n11636_not
g74232 not n52811 ; n52811_not
g74233 not n12176 ; n12176_not
g74234 not n40085 ; n40085_not
g74235 not n28070 ; n28070_not
g74236 not n24218 ; n24218_not
g74237 not n24515 ; n24515_not
g74238 not n56150 ; n56150_not
g74239 not n42614 ; n42614_not
g74240 not n24227 ; n24227_not
g74241 not n24506 ; n24506_not
g74242 not n51317 ; n51317_not
g74243 not n24236 ; n24236_not
g74244 not n17306 ; n17306_not
g74245 not n42704 ; n42704_not
g74246 not n24245 ; n24245_not
g74247 not n51326 ; n51326_not
g74248 not n40094 ; n40094_not
g74249 not n42029 ; n42029_not
g74250 not n24182 ; n24182_not
g74251 not n24533 ; n24533_not
g74252 not n42092 ; n42092_not
g74253 not n24191 ; n24191_not
g74254 not n48014 ; n48014_not
g74255 not n32192 ; n32192_not
g74256 not n24209 ; n24209_not
g74257 not n51335 ; n51335_not
g74258 not n24308 ; n24308_not
g74259 not n24461 ; n24461_not
g74260 not n24317 ; n24317_not
g74261 not n44207 ; n44207_not
g74262 not n24326 ; n24326_not
g74263 not n34514 ; n34514_not
g74264 not n51290 ; n51290_not
g74265 not n24335 ; n24335_not
g74266 not n34910 ; n34910_not
g74267 not n34820 ; n34820_not
g74268 not n24344 ; n24344_not
g74269 not n24443 ; n24443_not
g74270 not n17315 ; n17315_not
g74271 not n12077 ; n12077_not
g74272 not n24254 ; n24254_not
g74273 not n51308 ; n51308_not
g74274 not n24263 ; n24263_not
g74275 not n31193 ; n31193_not
g74276 not n24272 ; n24272_not
g74277 not n24281 ; n24281_not
g74278 not n12095 ; n12095_not
g74279 not n24290 ; n24290_not
g74280 not n38600 ; n38600_not
g74281 not n48140 ; n48140_not
g74282 not n24470 ; n24470_not
g74283 not n51344 ; n51344_not
g74284 not n52622 ; n52622_not
g74285 not n37115 ; n37115_not
g74286 not n51407 ; n51407_not
g74287 not n17216 ; n17216_not
g74288 not n11483 ; n11483_not
g74289 not n48023 ; n48023_not
g74290 not n32165 ; n32165_not
g74291 not n48212 ; n48212_not
g74292 not n45251 ; n45251_not
g74293 not n40661 ; n40661_not
g74294 not n54323 ; n54323_not
g74295 not n29051 ; n29051_not
g74296 not n52631 ; n52631_not
g74297 not n17351 ; n17351_not
g74298 not n17225 ; n17225_not
g74299 not n48203 ; n48203_not
g74300 not n56123 ; n56123_not
g74301 not n45530 ; n45530_not
g74302 not n12086 ; n12086_not
g74303 not n42731 ; n42731_not
g74304 not n38006 ; n38006_not
g74305 not n47024 ; n47024_not
g74306 not n31157 ; n31157_not
g74307 not n48230 ; n48230_not
g74308 not n23723 ; n23723_not
g74309 not n29060 ; n29060_not
g74310 not n44234 ; n44234_not
g74311 not n17207 ; n17207_not
g74312 not n42119 ; n42119_not
g74313 not n28034 ; n28034_not
g74314 not n48221 ; n48221_not
g74315 not n47501 ; n47501_not
g74316 not n23714 ; n23714_not
g74317 not n54305 ; n54305_not
g74318 not n52901 ; n52901_not
g74319 not n11492 ; n11492_not
g74320 not n18503 ; n18503_not
g74321 not n42083 ; n42083_not
g74322 not n17252 ; n17252_not
g74323 not n40634 ; n40634_not
g74324 not n11447 ; n11447_not
g74325 not n11456 ; n11456_not
g74326 not n55025 ; n55025_not
g74327 not n51272 ; n51272_not
g74328 not n51380 ; n51380_not
g74329 not n28061 ; n28061_not
g74330 not n23633 ; n23633_not
g74331 not n46313 ; n46313_not
g74332 not n32174 ; n32174_not
g74333 not n23642 ; n23642_not
g74334 not n47015 ; n47015_not
g74335 not n52802 ; n52802_not
g74336 not n44225 ; n44225_not
g74337 not n48131 ; n48131_not
g74338 not n37016 ; n37016_not
g74339 not n17234 ; n17234_not
g74340 not n46304 ; n46304_not
g74341 not n44432 ; n44432_not
g74342 not n32039 ; n32039_not
g74343 not n42722 ; n42722_not
g74344 not n40652 ; n40652_not
g74345 not n17342 ; n17342_not
g74346 not n55052 ; n55052_not
g74347 not n56132 ; n56132_not
g74348 not n37025 ; n37025_not
g74349 not n17243 ; n17243_not
g74350 not n17162 ; n17162_not
g74351 not n45341 ; n45341_not
g74352 not n37106 ; n37106_not
g74353 not n18440 ; n18440_not
g74354 not n32075 ; n32075_not
g74355 not n11168 ; n11168_not
g74356 not n51551 ; n51551_not
g74357 not n18512 ; n18512_not
g74358 not n23345 ; n23345_not
g74359 not n50228 ; n50228_not
g74360 not n47105 ; n47105_not
g74361 not n45116 ; n45116_not
g74362 not n31823 ; n31823_not
g74363 not n11159 ; n11159_not
g74364 not n23336 ; n23336_not
g74365 not n35207 ; n35207_not
g74366 not n31148 ; n31148_not
g74367 not n34505 ; n34505_not
g74368 not n23372 ; n23372_not
g74369 not n38402 ; n38402_not
g74370 not n12950 ; n12950_not
g74371 not n11186 ; n11186_not
g74372 not n17018 ; n17018_not
g74373 not n23363 ; n23363_not
g74374 not n55142 ; n55142_not
g74375 not n23354 ; n23354_not
g74376 not n11177 ; n11177_not
g74377 not n11096 ; n11096_not
g74378 not n17009 ; n17009_not
g74379 not n46160 ; n46160_not
g74380 not n17513 ; n17513_not
g74381 not n23291 ; n23291_not
g74382 not n12617 ; n12617_not
g74383 not n11087 ; n11087_not
g74384 not n31139 ; n31139_not
g74385 not n34460 ; n34460_not
g74386 not n23282 ; n23282_not
g74387 not n11078 ; n11078_not
g74388 not n42812 ; n42812_not
g74389 not n54125 ; n54125_not
g74390 not n23327 ; n23327_not
g74391 not n17504 ; n17504_not
g74392 not n19133 ; n19133_not
g74393 not n23318 ; n23318_not
g74394 not n44090 ; n44090_not
g74395 not n25343 ; n25343_not
g74396 not n23309 ; n23309_not
g74397 not n19142 ; n19142_not
g74398 not n53108 ; n53108_not
g74399 not n32408 ; n32408_not
g74400 not n42056 ; n42056_not
g74401 not n23435 ; n23435_not
g74402 not n31814 ; n31814_not
g74403 not n25253 ; n25253_not
g74404 not n12923 ; n12923_not
g74405 not n29501 ; n29501_not
g74406 not n46214 ; n46214_not
g74407 not n23426 ; n23426_not
g74408 not n48320 ; n48320_not
g74409 not n53090 ; n53090_not
g74410 not n51146 ; n51146_not
g74411 not n51542 ; n51542_not
g74412 not n23417 ; n23417_not
g74413 not n16901 ; n16901_not
g74414 not n51164 ; n51164_not
g74415 not n25235 ; n25235_not
g74416 not n56033 ; n56033_not
g74417 not n12914 ; n12914_not
g74418 not n55124 ; n55124_not
g74419 not n47321 ; n47321_not
g74420 not n23453 ; n23453_not
g74421 not n51083 ; n51083_not
g74422 not n42047 ; n42047_not
g74423 not n35180 ; n35180_not
g74424 not n10970 ; n10970_not
g74425 not n23444 ; n23444_not
g74426 not n51155 ; n51155_not
g74427 not n54143 ; n54143_not
g74428 not n51092 ; n51092_not
g74429 not n38420 ; n38420_not
g74430 not n12347 ; n12347_not
g74431 not n38411 ; n38411_not
g74432 not n42803 ; n42803_not
g74433 not n19115 ; n19115_not
g74434 not n36440 ; n36440_not
g74435 not n46205 ; n46205_not
g74436 not n23390 ; n23390_not
g74437 not n51137 ; n51137_not
g74438 not n22922 ; n22922_not
g74439 not n12941 ; n12941_not
g74440 not n42623 ; n42623_not
g74441 not n11195 ; n11195_not
g74442 not n46700 ; n46700_not
g74443 not n23381 ; n23381_not
g74444 not n34145 ; n34145_not
g74445 not n12662 ; n12662_not
g74446 not n12932 ; n12932_not
g74447 not n23408 ; n23408_not
g74448 not n16910 ; n16910_not
g74449 not n17027 ; n17027_not
g74450 not n56240 ; n56240_not
g74451 not n54314 ; n54314_not
g74452 not n23183 ; n23183_not
g74453 not n35243 ; n35243_not
g74454 not n25433 ; n25433_not
g74455 not n52064 ; n52064_not
g74456 not n46502 ; n46502_not
g74457 not n31832 ; n31832_not
g74458 not n23174 ; n23174_not
g74459 not n32426 ; n32426_not
g74460 not n30932 ; n30932_not
g74461 not n47123 ; n47123_not
g74462 not n50381 ; n50381_not
g74463 not n32066 ; n32066_not
g74464 not n13085 ; n13085_not
g74465 not n50363 ; n50363_not
g74466 not n17540 ; n17540_not
g74467 not n34433 ; n34433_not
g74468 not n12572 ; n12572_not
g74469 not n13094 ; n13094_not
g74470 not n45062 ; n45062_not
g74471 not n52055 ; n52055_not
g74472 not n44306 ; n44306_not
g74473 not n23192 ; n23192_not
g74474 not n55160 ; n55160_not
g74475 not n50372 ; n50372_not
g74476 not n32363 ; n32363_not
g74477 not n13139 ; n13139_not
g74478 not n46511 ; n46511_not
g74479 not n23138 ; n23138_not
g74480 not n41840 ; n41840_not
g74481 not n19205 ; n19205_not
g74482 not n23129 ; n23129_not
g74483 not n23165 ; n23165_not
g74484 not n35252 ; n35252_not
g74485 not n51074 ; n51074_not
g74486 not n23156 ; n23156_not
g74487 not n52073 ; n52073_not
g74488 not n46133 ; n46133_not
g74489 not n50390 ; n50390_not
g74490 not n45314 ; n45314_not
g74491 not n23147 ; n23147_not
g74492 not n23057 ; n23057_not
g74493 not n34451 ; n34451_not
g74494 not n31508 ; n31508_not
g74495 not n19160 ; n19160_not
g74496 not n52028 ; n52028_not
g74497 not n23255 ; n23255_not
g74498 not n50345 ; n50345_not
g74499 not n40760 ; n40760_not
g74500 not n13049 ; n13049_not
g74501 not n23246 ; n23246_not
g74502 not n32417 ; n32417_not
g74503 not n35225 ; n35225_not
g74504 not n51560 ; n51560_not
g74505 not n46151 ; n46151_not
g74506 not n52019 ; n52019_not
g74507 not n17522 ; n17522_not
g74508 not n23273 ; n23273_not
g74509 not n42821 ; n42821_not
g74510 not n45125 ; n45125_not
g74511 not n23264 ; n23264_not
g74512 not n56015 ; n56015_not
g74513 not n53117 ; n53117_not
g74514 not n16280 ; n16280_not
g74515 not n23219 ; n23219_not
g74516 not n28511 ; n28511_not
g74517 not n13076 ; n13076_not
g74518 not n53126 ; n53126_not
g74519 not n50147 ; n50147_not
g74520 not n42830 ; n42830_not
g74521 not n13058 ; n13058_not
g74522 not n52037 ; n52037_not
g74523 not n23237 ; n23237_not
g74524 not n17531 ; n17531_not
g74525 not n46142 ; n46142_not
g74526 not n52640 ; n52640_not
g74527 not n52046 ; n52046_not
g74528 not n23228 ; n23228_not
g74529 not n44081 ; n44081_not
g74530 not n13067 ; n13067_not
g74531 not n50354 ; n50354_not
g74532 not n12194 ; n12194_not
g74533 not n44144 ; n44144_not
g74534 not n45224 ; n45224_not
g74535 not n11465 ; n11465_not
g74536 not n29204 ; n29204_not
g74537 not n12752 ; n12752_not
g74538 not n17054 ; n17054_not
g74539 not n18602 ; n18602_not
g74540 not n43712 ; n43712_not
g74541 not n12743 ; n12743_not
g74542 not n17423 ; n17423_not
g74543 not n29231 ; n29231_not
g74544 not n12734 ; n12734_not
g74545 not n29222 ; n29222_not
g74546 not n17063 ; n17063_not
g74547 not n23741 ; n23741_not
g74548 not n29213 ; n29213_not
g74549 not n44135 ; n44135_not
g74550 not n17441 ; n17441_not
g74551 not n51218 ; n51218_not
g74552 not n11393 ; n11393_not
g74553 not n40904 ; n40904_not
g74554 not n29303 ; n29303_not
g74555 not n19043 ; n19043_not
g74556 not n11384 ; n11384_not
g74557 not n51227 ; n51227_not
g74558 not n47042 ; n47042_not
g74559 not n12770 ; n12770_not
g74560 not n51506 ; n51506_not
g74561 not n46241 ; n46241_not
g74562 not n17432 ; n17432_not
g74563 not n45503 ; n45503_not
g74564 not n53054 ; n53054_not
g74565 not n23831 ; n23831_not
g74566 not n12329 ; n12329_not
g74567 not n12671 ; n12671_not
g74568 not n17414 ; n17414_not
g74569 not n32327 ; n32327_not
g74570 not n17081 ; n17081_not
g74571 not n24524 ; n24524_not
g74572 not n12293 ; n12293_not
g74573 not n51245 ; n51245_not
g74574 not n50912 ; n50912_not
g74575 not n56222 ; n56222_not
g74576 not n12338 ; n12338_not
g74577 not n12266 ; n12266_not
g74578 not n45512 ; n45512_not
g74579 not n12257 ; n12257_not
g74580 not n12248 ; n12248_not
g74581 not n12716 ; n12716_not
g74582 not n12239 ; n12239_not
g74583 not n51047 ; n51047_not
g74584 not n37160 ; n37160_not
g74585 not n12284 ; n12284_not
g74586 not n12275 ; n12275_not
g74587 not n11555 ; n11555_not
g74588 not n32129 ; n32129_not
g74589 not n29240 ; n29240_not
g74590 not n51236 ; n51236_not
g74591 not n53045 ; n53045_not
g74592 not n29402 ; n29402_not
g74593 not n11294 ; n11294_not
g74594 not n54170 ; n54170_not
g74595 not n23525 ; n23525_not
g74596 not n44117 ; n44117_not
g74597 not n56231 ; n56231_not
g74598 not n23516 ; n23516_not
g74599 not n11285 ; n11285_not
g74600 not n10943 ; n10943_not
g74601 not n40931 ; n40931_not
g74602 not n51182 ; n51182_not
g74603 not n47060 ; n47060_not
g74604 not n12860 ; n12860_not
g74605 not n23552 ; n23552_not
g74606 not n22832 ; n22832_not
g74607 not n42641 ; n42641_not
g74608 not n46223 ; n46223_not
g74609 not n45323 ; n45323_not
g74610 not n23543 ; n23543_not
g74611 not n45107 ; n45107_not
g74612 not n24434 ; n24434_not
g74613 not n51191 ; n51191_not
g74614 not n51524 ; n51524_not
g74615 not n23534 ; n23534_not
g74616 not n40940 ; n40940_not
g74617 not n11258 ; n11258_not
g74618 not n12905 ; n12905_not
g74619 not n25226 ; n25226_not
g74620 not n23471 ; n23471_not
g74621 not n53081 ; n53081_not
g74622 not n51533 ; n51533_not
g74623 not n44108 ; n44108_not
g74624 not n11249 ; n11249_not
g74625 not n48311 ; n48311_not
g74626 not n23462 ; n23462_not
g74627 not n23507 ; n23507_not
g74628 not n31166 ; n31166_not
g74629 not n11276 ; n11276_not
g74630 not n43802 ; n43802_not
g74631 not n54161 ; n54161_not
g74632 not n53072 ; n53072_not
g74633 not n44414 ; n44414_not
g74634 not n55115 ; n55115_not
g74635 not n11267 ; n11267_not
g74636 not n48104 ; n48104_not
g74637 not n32372 ; n32372_not
g74638 not n51173 ; n51173_not
g74639 not n32084 ; n32084_not
g74640 not n23480 ; n23480_not
g74641 not n17036 ; n17036_not
g74642 not n12806 ; n12806_not
g74643 not n51515 ; n51515_not
g74644 not n11366 ; n11366_not
g74645 not n40193 ; n40193_not
g74646 not n12815 ; n12815_not
g74647 not n48113 ; n48113_not
g74648 not n12824 ; n12824_not
g74649 not n46232 ; n46232_not
g74650 not n23651 ; n23651_not
g74651 not n29312 ; n29312_not
g74652 not n56060 ; n56060_not
g74653 not n31463 ; n31463_not
g74654 not n11375 ; n11375_not
g74655 not n29321 ; n29321_not
g74656 not n48302 ; n48302_not
g74657 not n19052 ; n19052_not
g74658 not n46340 ; n46340_not
g74659 not n40913 ; n40913_not
g74660 not n28232 ; n28232_not
g74661 not n53063 ; n53063_not
g74662 not n44126 ; n44126_not
g74663 not n12707 ; n12707_not
g74664 not n23570 ; n23570_not
g74665 not n12851 ; n12851_not
g74666 not n28601 ; n28601_not
g74667 not n40922 ; n40922_not
g74668 not n19070 ; n19070_not
g74669 not n23561 ; n23561_not
g74670 not n11357 ; n11357_not
g74671 not n17450 ; n17450_not
g74672 not n43703 ; n43703_not
g74673 not n12833 ; n12833_not
g74674 not n11348 ; n11348_not
g74675 not n40805 ; n40805_not
g74676 not n37124 ; n37124_not
g74677 not n47051 ; n47051_not
g74678 not n11339 ; n11339_not
g74679 not n12842 ; n12842_not
g74680 not n51209 ; n51209_not
g74681 not n15245 ; n15245_not
g74682 not n57041 ; n57041_not
g74683 not n53441 ; n53441_not
g74684 not n15254 ; n15254_not
g74685 not n55511 ; n55511_not
g74686 not n51902 ; n51902_not
g74687 not n37430 ; n37430_not
g74688 not n45152 ; n45152_not
g74689 not n27233 ; n27233_not
g74690 not n15263 ; n15263_not
g74691 not n16514 ; n16514_not
g74692 not n33380 ; n33380_not
g74693 not n16505 ; n16505_not
g74694 not n30491 ; n30491_not
g74695 not n15218 ; n15218_not
g74696 not n20618 ; n20618_not
g74697 not n31562 ; n31562_not
g74698 not n37421 ; n37421_not
g74699 not n33416 ; n33416_not
g74700 not n41561 ; n41561_not
g74701 not n15227 ; n15227_not
g74702 not n18035 ; n18035_not
g74703 not n15236 ; n15236_not
g74704 not n33407 ; n33407_not
g74705 not n53720 ; n53720_not
g74706 not n35900 ; n35900_not
g74707 not n41363 ; n41363_not
g74708 not n53711 ; n53711_not
g74709 not n19511 ; n19511_not
g74710 not n15155 ; n15155_not
g74711 not n32615 ; n32615_not
g74712 not n31544 ; n31544_not
g74713 not n18026 ; n18026_not
g74714 not n19502 ; n19502_not
g74715 not n55502 ; n55502_not
g74716 not n26081 ; n26081_not
g74717 not n53405 ; n53405_not
g74718 not n41552 ; n41552_not
g74719 not n15308 ; n15308_not
g74720 not n33362 ; n33362_not
g74721 not n20654 ; n20654_not
g74722 not n31553 ; n31553_not
g74723 not n57050 ; n57050_not
g74724 not n15173 ; n15173_not
g74725 not n15272 ; n15272_not
g74726 not n31634 ; n31634_not
g74727 not n15164 ; n15164_not
g74728 not n19520 ; n19520_not
g74729 not n15281 ; n15281_not
g74730 not n26090 ; n26090_not
g74731 not n15290 ; n15290_not
g74732 not n20645 ; n20645_not
g74733 not n26126 ; n26126_not
g74734 not n37412 ; n37412_not
g74735 not n41138 ; n41138_not
g74736 not n14705 ; n14705_not
g74737 not n33344 ; n33344_not
g74738 not n43136 ; n43136_not
g74739 not n21095 ; n21095_not
g74740 not n26801 ; n26801_not
g74741 not n31751 ; n31751_not
g74742 not n33452 ; n33452_not
g74743 not n31571 ; n31571_not
g74744 not n54224 ; n54224_not
g74745 not n33353 ; n33353_not
g74746 not n21086 ; n21086_not
g74747 not n19601 ; n19601_not
g74748 not n15119 ; n15119_not
g74749 not n26135 ; n26135_not
g74750 not n14741 ; n14741_not
g74751 not n35711 ; n35711_not
g74752 not n36062 ; n36062_not
g74753 not n30284 ; n30284_not
g74754 not n14732 ; n14732_not
g74755 not n47222 ; n47222_not
g74756 not n35702 ; n35702_not
g74757 not n14723 ; n14723_not
g74758 not n33461 ; n33461_not
g74759 not n27701 ; n27701_not
g74760 not n14714 ; n14714_not
g74761 not n15137 ; n15137_not
g74762 not n14633 ; n14633_not
g74763 not n15182 ; n15182_not
g74764 not n14624 ; n14624_not
g74765 not n18044 ; n18044_not
g74766 not n42407 ; n42407_not
g74767 not n14615 ; n14615_not
g74768 not n21059 ; n21059_not
g74769 not n33425 ; n33425_not
g74770 not n30482 ; n30482_not
g74771 not n14606 ; n14606_not
g74772 not n20609 ; n20609_not
g74773 not n55520 ; n55520_not
g74774 not n51911 ; n51911_not
g74775 not n43145 ; n43145_not
g74776 not n57014 ; n57014_not
g74777 not n15209 ; n15209_not
g74778 not n41570 ; n41570_not
g74779 not n33443 ; n33443_not
g74780 not n14660 ; n14660_not
g74781 not n41282 ; n41282_not
g74782 not n26810 ; n26810_not
g74783 not n21077 ; n21077_not
g74784 not n14651 ; n14651_not
g74785 not n26117 ; n26117_not
g74786 not n14642 ; n14642_not
g74787 not n33434 ; n33434_not
g74788 not n21068 ; n21068_not
g74789 not n15443 ; n15443_not
g74790 not n20870 ; n20870_not
g74791 not n19403 ; n19403_not
g74792 not n27602 ; n27602_not
g74793 not n42434 ; n42434_not
g74794 not n15452 ; n15452_not
g74795 not n16460 ; n16460_not
g74796 not n33272 ; n33272_not
g74797 not n20861 ; n20861_not
g74798 not n30518 ; n30518_not
g74799 not n57113 ; n57113_not
g74800 not n33263 ; n33263_not
g74801 not n15065 ; n15065_not
g74802 not n15461 ; n15461_not
g74803 not n43181 ; n43181_not
g74804 not n31535 ; n31535_not
g74805 not n26900 ; n26900_not
g74806 not n27611 ; n27611_not
g74807 not n33290 ; n33290_not
g74808 not n19412 ; n19412_not
g74809 not n15425 ; n15425_not
g74810 not n20708 ; n20708_not
g74811 not n15083 ; n15083_not
g74812 not n15434 ; n15434_not
g74813 not n30338 ; n30338_not
g74814 not n39311 ; n39311_not
g74815 not n41345 ; n41345_not
g74816 not n15074 ; n15074_not
g74817 not n18008 ; n18008_not
g74818 not n41525 ; n41525_not
g74819 not n31625 ; n31625_not
g74820 not n20834 ; n20834_not
g74821 not n39320 ; n39320_not
g74822 not n43190 ; n43190_not
g74823 not n33245 ; n33245_not
g74824 not n20735 ; n20735_not
g74825 not n32642 ; n32642_not
g74826 not n20825 ; n20825_not
g74827 not n30527 ; n30527_not
g74828 not n31526 ; n31526_not
g74829 not n20816 ; n20816_not
g74830 not n20852 ; n20852_not
g74831 not n43028 ; n43028_not
g74832 not n57122 ; n57122_not
g74833 not n45422 ; n45422_not
g74834 not n15470 ; n15470_not
g74835 not n20843 ; n20843_not
g74836 not n27017 ; n27017_not
g74837 not n16541 ; n16541_not
g74838 not n33254 ; n33254_not
g74839 not n47231 ; n47231_not
g74840 not n41516 ; n41516_not
g74841 not n30347 ; n30347_not
g74842 not n57131 ; n57131_not
g74843 not n18017 ; n18017_not
g74844 not n26072 ; n26072_not
g74845 not n41318 ; n41318_not
g74846 not n53450 ; n53450_not
g74847 not n32624 ; n32624_not
g74848 not n15344 ; n15344_not
g74849 not n41543 ; n41543_not
g74850 not n20942 ; n20942_not
g74851 not n15128 ; n15128_not
g74852 not n15353 ; n15353_not
g74853 not n33335 ; n33335_not
g74854 not n20933 ; n20933_not
g74855 not n15317 ; n15317_not
g74856 not n20663 ; n20663_not
g74857 not n42425 ; n42425_not
g74858 not n20960 ; n20960_not
g74859 not n15326 ; n15326_not
g74860 not n53702 ; n53702_not
g74861 not n39113 ; n39113_not
g74862 not n15335 ; n15335_not
g74863 not n20951 ; n20951_not
g74864 not n20690 ; n20690_not
g74865 not n33317 ; n33317_not
g74866 not n20906 ; n20906_not
g74867 not n19430 ; n19430_not
g74868 not n27620 ; n27620_not
g74869 not n43172 ; n43172_not
g74870 not n43019 ; n43019_not
g74871 not n39302 ; n39302_not
g74872 not n53423 ; n53423_not
g74873 not n15407 ; n15407_not
g74874 not n19421 ; n19421_not
g74875 not n15416 ; n15416_not
g74876 not n41372 ; n41372_not
g74877 not n15362 ; n15362_not
g74878 not n41327 ; n41327_not
g74879 not n39104 ; n39104_not
g74880 not n31724 ; n31724_not
g74881 not n20924 ; n20924_not
g74882 not n36107 ; n36107_not
g74883 not n15371 ; n15371_not
g74884 not n30329 ; n30329_not
g74885 not n41534 ; n41534_not
g74886 not n20915 ; n20915_not
g74887 not n15380 ; n15380_not
g74888 not n41381 ; n41381_not
g74889 not n31616 ; n31616_not
g74890 not n14822 ; n14822_not
g74891 not n33614 ; n33614_not
g74892 not n53810 ; n53810_not
g74893 not n14426 ; n14426_not
g74894 not n41615 ; n41615_not
g74895 not n26225 ; n26225_not
g74896 not n43082 ; n43082_not
g74897 not n21347 ; n21347_not
g74898 not n50237 ; n50237_not
g74899 not n14831 ; n14831_not
g74900 not n41336 ; n41336_not
g74901 not n51830 ; n51830_not
g74902 not n14840 ; n14840_not
g74903 not n33605 ; n33605_not
g74904 not n14417 ; n14417_not
g74905 not n26630 ; n26630_not
g74906 not n42380 ; n42380_not
g74907 not n21374 ; n21374_not
g74908 not n30086 ; n30086_not
g74909 not n26612 ; n26612_not
g74910 not n14804 ; n14804_not
g74911 not n21365 ; n21365_not
g74912 not n14813 ; n14813_not
g74913 not n14435 ; n14435_not
g74914 not n42371 ; n42371_not
g74915 not n26621 ; n26621_not
g74916 not n55223 ; n55223_not
g74917 not n21194 ; n21194_not
g74918 not n31607 ; n31607_not
g74919 not n26207 ; n26207_not
g74920 not n50318 ; n50318_not
g74921 not n43091 ; n43091_not
g74922 not n56420 ; n56420_not
g74923 not n56411 ; n56411_not
g74924 not n14390 ; n14390_not
g74925 not n41606 ; n41606_not
g74926 not n30725 ; n30725_not
g74927 not n27710 ; n27710_not
g74928 not n14903 ; n14903_not
g74929 not n56402 ; n56402_not
g74930 not n26216 ; n26216_not
g74931 not n55610 ; n55610_not
g74932 not n21149 ; n21149_not
g74933 not n21329 ; n21329_not
g74934 not n21158 ; n21158_not
g74935 not n53801 ; n53801_not
g74936 not n21167 ; n21167_not
g74937 not n47141 ; n47141_not
g74938 not n21176 ; n21176_not
g74939 not n18080 ; n18080_not
g74940 not n42443 ; n42443_not
g74941 not n39203 ; n39203_not
g74942 not n55601 ; n55601_not
g74943 not n21185 ; n21185_not
g74944 not n36611 ; n36611_not
g74945 not n33515 ; n33515_not
g74946 not n14480 ; n14480_not
g74947 not n51803 ; n51803_not
g74948 not n21437 ; n21437_not
g74949 not n56600 ; n56600_not
g74950 not n26252 ; n26252_not
g74951 not n41192 ; n41192_not
g74952 not n14471 ; n14471_not
g74953 not n35720 ; n35720_not
g74954 not n33524 ; n33524_not
g74955 not n41624 ; n41624_not
g74956 not n26261 ; n26261_not
g74957 not n21464 ; n21464_not
g74958 not n30563 ; n30563_not
g74959 not n21455 ; n21455_not
g74960 not n30095 ; n30095_not
g74961 not n33506 ; n33506_not
g74962 not n17810 ; n17810_not
g74963 not n33560 ; n33560_not
g74964 not n41183 ; n41183_not
g74965 not n33641 ; n33641_not
g74966 not n42461 ; n42461_not
g74967 not n21392 ; n21392_not
g74968 not n33632 ; n33632_not
g74969 not n41255 ; n41255_not
g74970 not n56510 ; n56510_not
g74971 not n56501 ; n56501_not
g74972 not n26603 ; n26603_not
g74973 not n31652 ; n31652_not
g74974 not n30743 ; n30743_not
g74975 not n50327 ; n50327_not
g74976 not n14750 ; n14750_not
g74977 not n33533 ; n33533_not
g74978 not n21419 ; n21419_not
g74979 not n42362 ; n42362_not
g74980 not n44531 ; n44531_not
g74981 not n33542 ; n33542_not
g74982 not n14462 ; n14462_not
g74983 not n51812 ; n51812_not
g74984 not n33551 ; n33551_not
g74985 not n30752 ; n30752_not
g74986 not n30680 ; n30680_not
g74987 not n31580 ; n31580_not
g74988 not n15047 ; n15047_not
g74989 not n41156 ; n41156_not
g74990 not n14921 ; n14921_not
g74991 not n14912 ; n14912_not
g74992 not n26162 ; n26162_not
g74993 not n45134 ; n45134_not
g74994 not n39140 ; n39140_not
g74995 not n15029 ; n15029_not
g74996 not n39230 ; n39230_not
g74997 not n18053 ; n18053_not
g74998 not n20564 ; n20564_not
g74999 not n46520 ; n46520_not
g75000 not n20573 ; n20573_not
g75001 not n41147 ; n41147_not
g75002 not n51731 ; n51731_not
g75003 not n33470 ; n33470_not
g75004 not n53360 ; n53360_not
g75005 not n37403 ; n37403_not
g75006 not n20555 ; n20555_not
g75007 not n36053 ; n36053_not
g75008 not n19610 ; n19610_not
g75009 not n51722 ; n51722_not
g75010 not n30275 ; n30275_not
g75011 not n45413 ; n45413_not
g75012 not n15092 ; n15092_not
g75013 not n14372 ; n14372_not
g75014 not n30257 ; n30257_not
g75015 not n21257 ; n21257_not
g75016 not n14930 ; n14930_not
g75017 not n41174 ; n41174_not
g75018 not n18071 ; n18071_not
g75019 not n35801 ; n35801_not
g75020 not n21248 ; n21248_not
g75021 not n45044 ; n45044_not
g75022 not n20492 ; n20492_not
g75023 not n14381 ; n14381_not
g75024 not n21284 ; n21284_not
g75025 not n36521 ; n36521_not
g75026 not n19700 ; n19700_not
g75027 not n21239 ; n21239_not
g75028 not n31733 ; n31733_not
g75029 not n21275 ; n21275_not
g75030 not n39212 ; n39212_not
g75031 not n55043 ; n55043_not
g75032 not n21266 ; n21266_not
g75033 not n31643 ; n31643_not
g75034 not n26171 ; n26171_not
g75035 not n39221 ; n39221_not
g75036 not n30707 ; n30707_not
g75037 not n20519 ; n20519_not
g75038 not n43127 ; n43127_not
g75039 not n41165 ; n41165_not
g75040 not n53351 ; n53351_not
g75041 not n26720 ; n26720_not
g75042 not n33308 ; n33308_not
g75043 not n20528 ; n20528_not
g75044 not n51713 ; n51713_not
g75045 not n18062 ; n18062_not
g75046 not n56330 ; n56330_not
g75047 not n35810 ; n35810_not
g75048 not n56321 ; n56321_not
g75049 not n26702 ; n26702_not
g75050 not n26180 ; n26180_not
g75051 not n14345 ; n14345_not
g75052 not n45800 ; n45800_not
g75053 not n53414 ; n53414_not
g75054 not n26711 ; n26711_not
g75055 not n32705 ; n32705_not
g75056 not n20168 ; n20168_not
g75057 not n27242 ; n27242_not
g75058 not n39023 ; n39023_not
g75059 not n27206 ; n27206_not
g75060 not n20393 ; n20393_not
g75061 not n55322 ; n55322_not
g75062 not n32543 ; n32543_not
g75063 not n57410 ; n57410_not
g75064 not n30455 ; n30455_not
g75065 not n16244 ; n16244_not
g75066 not n16019 ; n16019_not
g75067 not n30374 ; n30374_not
g75068 not n27224 ; n27224_not
g75069 not n27107 ; n27107_not
g75070 not n44513 ; n44513_not
g75071 not n32561 ; n32561_not
g75072 not n43226 ; n43226_not
g75073 not n57401 ; n57401_not
g75074 not n27215 ; n27215_not
g75075 not n27422 ; n27422_not
g75076 not n55331 ; n55331_not
g75077 not n16253 ; n16253_not
g75078 not n32552 ; n32552_not
g75079 not n43217 ; n43217_not
g75080 not n27413 ; n27413_not
g75081 not n27260 ; n27260_not
g75082 not n20366 ; n20366_not
g75083 not n16046 ; n16046_not
g75084 not n53513 ; n53513_not
g75085 not n39050 ; n39050_not
g75086 not n20357 ; n20357_not
g75087 not n15740 ; n15740_not
g75088 not n16055 ; n16055_not
g75089 not n36206 ; n36206_not
g75090 not n27251 ; n27251_not
g75091 not n20384 ; n20384_not
g75092 not n32534 ; n32534_not
g75093 not n16028 ; n16028_not
g75094 not n15632 ; n15632_not
g75095 not n20177 ; n20177_not
g75096 not n41435 ; n41435_not
g75097 not n31742 ; n31742_not
g75098 not n20375 ; n20375_not
g75099 not n16037 ; n16037_not
g75100 not n30383 ; n30383_not
g75101 not n32525 ; n32525_not
g75102 not n36305 ; n36305_not
g75103 not n26423 ; n26423_not
g75104 not n30437 ; n30437_not
g75105 not n15812 ; n15812_not
g75106 not n20465 ; n20465_not
g75107 not n15920 ; n15920_not
g75108 not n26414 ; n26414_not
g75109 not n51821 ; n51821_not
g75110 not n26405 ; n26405_not
g75111 not n20456 ; n20456_not
g75112 not n36152 ; n36152_not
g75113 not n15821 ; n15821_not
g75114 not n15902 ; n15902_not
g75115 not n26441 ; n26441_not
g75116 not n20483 ; n20483_not
g75117 not n37601 ; n37601_not
g75118 not n53603 ; n53603_not
g75119 not n43271 ; n43271_not
g75120 not n26432 ; n26432_not
g75121 not n36143 ; n36143_not
g75122 not n15911 ; n15911_not
g75123 not n20474 ; n20474_not
g75124 not n20159 ; n20159_not
g75125 not n16262 ; n16262_not
g75126 not n41831 ; n41831_not
g75127 not n32903 ; n32903_not
g75128 not n20429 ; n20429_not
g75129 not n50273 ; n50273_not
g75130 not n41417 ; n41417_not
g75131 not n32714 ; n32714_not
g75132 not n43244 ; n43244_not
g75133 not n32570 ; n32570_not
g75134 not n27431 ; n27431_not
g75135 not n30446 ; n30446_not
g75136 not n55340 ; n55340_not
g75137 not n27440 ; n27440_not
g75138 not n30365 ; n30365_not
g75139 not n32921 ; n32921_not
g75140 not n41408 ; n41408_not
g75141 not n20447 ; n20447_not
g75142 not n16271 ; n16271_not
g75143 not n44522 ; n44522_not
g75144 not n43262 ; n43262_not
g75145 not n36161 ; n36161_not
g75146 not n32912 ; n32912_not
g75147 not n39014 ; n39014_not
g75148 not n45440 ; n45440_not
g75149 not n20438 ; n20438_not
g75150 not n41462 ; n41462_not
g75151 not n20258 ; n20258_not
g75152 not n16145 ; n16145_not
g75153 not n16154 ; n16154_not
g75154 not n36242 ; n36242_not
g75155 not n30428 ; n30428_not
g75156 not n27332 ; n27332_not
g75157 not n20249 ; n20249_not
g75158 not n32660 ; n32660_not
g75159 not n55304 ; n55304_not
g75160 not n45431 ; n45431_not
g75161 not n27314 ; n27314_not
g75162 not n20276 ; n20276_not
g75163 not n36260 ; n36260_not
g75164 not n44504 ; n44504_not
g75165 not n16136 ; n16136_not
g75166 not n27170 ; n27170_not
g75167 not n20267 ; n20267_not
g75168 not n27323 ; n27323_not
g75169 not n15641 ; n15641_not
g75170 not n27161 ; n27161_not
g75171 not n53531 ; n53531_not
g75172 not n16181 ; n16181_not
g75173 not n50183 ; n50183_not
g75174 not n27350 ; n27350_not
g75175 not n32750 ; n32750_not
g75176 not n41471 ; n41471_not
g75177 not n16190 ; n16190_not
g75178 not n36251 ; n36251_not
g75179 not n57500 ; n57500_not
g75180 not n43109 ; n43109_not
g75181 not n32741 ; n32741_not
g75182 not n16208 ; n16208_not
g75183 not n16163 ; n16163_not
g75184 not n30419 ; n30419_not
g75185 not n16217 ; n16217_not
g75186 not n27341 ; n27341_not
g75187 not n16172 ; n16172_not
g75188 not n15650 ; n15650_not
g75189 not n27152 ; n27152_not
g75190 not n39401 ; n39401_not
g75191 not n39410 ; n39410_not
g75192 not n16235 ; n16235_not
g75193 not n27125 ; n27125_not
g75194 not n15722 ; n15722_not
g75195 not n32822 ; n32822_not
g75196 not n16082 ; n16082_not
g75197 not n38105 ; n38105_not
g75198 not n20186 ; n20186_not
g75199 not n16091 ; n16091_not
g75200 not n27116 ; n27116_not
g75201 not n32840 ; n32840_not
g75202 not n20348 ; n20348_not
g75203 not n15731 ; n15731_not
g75204 not n32723 ; n32723_not
g75205 not n16064 ; n16064_not
g75206 not n27404 ; n27404_not
g75207 not n41444 ; n41444_not
g75208 not n41480 ; n41480_not
g75209 not n20339 ; n20339_not
g75210 not n32831 ; n32831_not
g75211 not n32633 ; n32633_not
g75212 not n16073 ; n16073_not
g75213 not n20294 ; n20294_not
g75214 not n43154 ; n43154_not
g75215 not n32732 ; n32732_not
g75216 not n55313 ; n55313_not
g75217 not n53540 ; n53540_not
g75218 not n20285 ; n20285_not
g75219 not n16118 ; n16118_not
g75220 not n16226 ; n16226_not
g75221 not n16127 ; n16127_not
g75222 not n20195 ; n20195_not
g75223 not n47240 ; n47240_not
g75224 not n41426 ; n41426_not
g75225 not n32813 ; n32813_not
g75226 not n30392 ; n30392_not
g75227 not n32804 ; n32804_not
g75228 not n41453 ; n41453_not
g75229 not n16109 ; n16109_not
g75230 not n27305 ; n27305_not
g75231 not n15623 ; n15623_not
g75232 not n33182 ; n33182_not
g75233 not n57212 ; n57212_not
g75234 not n39500 ; n39500_not
g75235 not n27044 ; n27044_not
g75236 not n19331 ; n19331_not
g75237 not n33173 ; n33173_not
g75238 not n33164 ; n33164_not
g75239 not n55421 ; n55421_not
g75240 not n20078 ; n20078_not
g75241 not n55133 ; n55133_not
g75242 not n20087 ; n20087_not
g75243 not n36350 ; n36350_not
g75244 not n20096 ; n20096_not
g75245 not n16424 ; n16424_not
g75246 not n19322 ; n19322_not
g75247 not n15614 ; n15614_not
g75248 not n16415 ; n16415_not
g75249 not n20717 ; n20717_not
g75250 not n33146 ; n33146_not
g75251 not n27530 ; n27530_not
g75252 not n27071 ; n27071_not
g75253 not n33137 ; n33137_not
g75254 not n27521 ; n27521_not
g75255 not n33128 ; n33128_not
g75256 not n55412 ; n55412_not
g75257 not n37511 ; n37511_not
g75258 not n57230 ; n57230_not
g75259 not n33155 ; n33155_not
g75260 not n19340 ; n19340_not
g75261 not n27062 ; n27062_not
g75262 not n20672 ; n20672_not
g75263 not n27035 ; n27035_not
g75264 not n20771 ; n20771_not
g75265 not n15524 ; n15524_not
g75266 not n33227 ; n33227_not
g75267 not n15533 ; n15533_not
g75268 not n43037 ; n43037_not
g75269 not n36008 ; n36008_not
g75270 not n57140 ; n57140_not
g75271 not n15506 ; n15506_not
g75272 not n27026 ; n27026_not
g75273 not n20744 ; n20744_not
g75274 not n33236 ; n33236_not
g75275 not n38114 ; n38114_not
g75276 not n20807 ; n20807_not
g75277 not n30536 ; n30536_not
g75278 not n15038 ; n15038_not
g75279 not n41507 ; n41507_not
g75280 not n15515 ; n15515_not
g75281 not n20753 ; n20753_not
g75282 not n42416 ; n42416_not
g75283 not n36026 ; n36026_not
g75284 not n37502 ; n37502_not
g75285 not n55430 ; n55430_not
g75286 not n57203 ; n57203_not
g75287 not n33191 ; n33191_not
g75288 not n20069 ; n20069_not
g75289 not n35612 ; n35612_not
g75290 not n36017 ; n36017_not
g75291 not n15542 ; n15542_not
g75292 not n33218 ; n33218_not
g75293 not n16442 ; n16442_not
g75294 not n19313 ; n19313_not
g75295 not n15551 ; n15551_not
g75296 not n35621 ; n35621_not
g75297 not n33209 ; n33209_not
g75298 not n15560 ; n15560_not
g75299 not n17900 ; n17900_not
g75300 not n26504 ; n26504_not
g75301 not n36314 ; n36314_not
g75302 not n33038 ; n33038_not
g75303 not n33029 ; n33029_not
g75304 not n27080 ; n27080_not
g75305 not n20537 ; n20537_not
g75306 not n43064 ; n43064_not
g75307 not n53612 ; n53612_not
g75308 not n43055 ; n43055_not
g75309 not n27134 ; n27134_not
g75310 not n33056 ; n33056_not
g75311 not n26522 ; n26522_not
g75312 not n53621 ; n53621_not
g75313 not n30545 ; n30545_not
g75314 not n26513 ; n26513_not
g75315 not n16307 ; n16307_not
g75316 not n46430 ; n46430_not
g75317 not n15830 ; n15830_not
g75318 not n26450 ; n26450_not
g75319 not n39005 ; n39005_not
g75320 not n53504 ; n53504_not
g75321 not n36134 ; n36134_not
g75322 not n50282 ; n50282_not
g75323 not n20627 ; n20627_not
g75324 not n36332 ; n36332_not
g75325 not n36071 ; n36071_not
g75326 not n50246 ; n50246_not
g75327 not n36341 ; n36341_not
g75328 not n55403 ; n55403_not
g75329 not n33119 ; n33119_not
g75330 not n15704 ; n15704_not
g75331 not n27512 ; n27512_not
g75332 not n27503 ; n27503_not
g75333 not n41390 ; n41390_not
g75334 not n50291 ; n50291_not
g75335 not n33065 ; n33065_not
g75336 not n30293 ; n30293_not
g75337 not n20582 ; n20582_not
g75338 not n36116 ; n36116_not
g75339 not n26540 ; n26540_not
g75340 not n16352 ; n16352_not
g75341 not n26531 ; n26531_not
g75342 not n43235 ; n43235_not
g75343 not n33092 ; n33092_not
g75344 not n31805 ; n31805_not
g75345 not n53630 ; n53630_not
g75346 not n36323 ; n36323_not
g75347 not n33083 ; n33083_not
g75348 not n57302 ; n57302_not
g75349 not n30554 ; n30554_not
g75350 not n33074 ; n33074_not
g75351 not n19151 ; n19151_not
g75352 not n14264 ; n14264_not
g75353 not n10187 ; n10187_not
g75354 not n50255 ; n50255_not
g75355 not n45170 ; n45170_not
g75356 not n14183 ; n14183_not
g75357 not n10178 ; n10178_not
g75358 not n26306 ; n26306_not
g75359 not n41291 ; n41291_not
g75360 not n37340 ; n37340_not
g75361 not n28115 ; n28115_not
g75362 not n30716 ; n30716_not
g75363 not n19106 ; n19106_not
g75364 not n10196 ; n10196_not
g75365 not n14174 ; n14174_not
g75366 not n40049 ; n40049_not
g75367 not n33830 ; n33830_not
g75368 not n21905 ; n21905_not
g75369 not n51740 ; n51740_not
g75370 not n40058 ; n40058_not
g75371 not n33920 ; n33920_not
g75372 not n28016 ; n28016_not
g75373 not n41642 ; n41642_not
g75374 not n41660 ; n41660_not
g75375 not n14552 ; n14552_not
g75376 not n18161 ; n18161_not
g75377 not n10169 ; n10169_not
g75378 not n31670 ; n31670_not
g75379 not n50192 ; n50192_not
g75380 not n36233 ; n36233_not
g75381 not n21473 ; n21473_not
g75382 not n21914 ; n21914_not
g75383 not n14192 ; n14192_not
g75384 not n14561 ; n14561_not
g75385 not n52424 ; n52424_not
g75386 not n37034 ; n37034_not
g75387 not n26315 ; n26315_not
g75388 not n53324 ; n53324_not
g75389 not n42335 ; n42335_not
g75390 not n10259 ; n10259_not
g75391 not n33740 ; n33740_not
g75392 not n14156 ; n14156_not
g75393 not n30068 ; n30068_not
g75394 not n39032 ; n39032_not
g75395 not n21941 ; n21941_not
g75396 not n33731 ; n33731_not
g75397 not n10268 ; n10268_not
g75398 not n21950 ; n21950_not
g75399 not n22049 ; n22049_not
g75400 not n30077 ; n30077_not
g75401 not n14165 ; n14165_not
g75402 not n44342 ; n44342_not
g75403 not n43721 ; n43721_not
g75404 not n35531 ; n35531_not
g75405 not n28124 ; n28124_not
g75406 not n31706 ; n31706_not
g75407 not n46601 ; n46601_not
g75408 not n18170 ; n18170_not
g75409 not n43811 ; n43811_not
g75410 not n14273 ; n14273_not
g75411 not n37331 ; n37331_not
g75412 not n53234 ; n53234_not
g75413 not n18143 ; n18143_not
g75414 not n18125 ; n18125_not
g75415 not n33812 ; n33812_not
g75416 not n40067 ; n40067_not
g75417 not n40076 ; n40076_not
g75418 not n26144 ; n26144_not
g75419 not n41651 ; n41651_not
g75420 not n10079 ; n10079_not
g75421 not n42344 ; n42344_not
g75422 not n16433 ; n16433_not
g75423 not n14246 ; n14246_not
g75424 not n26360 ; n26360_not
g75425 not n14219 ; n14219_not
g75426 not n35630 ; n35630_not
g75427 not n10088 ; n10088_not
g75428 not n38123 ; n38123_not
g75429 not n26342 ; n26342_not
g75430 not n18152 ; n18152_not
g75431 not n26351 ; n26351_not
g75432 not n35513 ; n35513_not
g75433 not n30059 ; n30059_not
g75434 not n14237 ; n14237_not
g75435 not n21428 ; n21428_not
g75436 not n40670 ; n40670_not
g75437 not n21293 ; n21293_not
g75438 not n14228 ; n14228_not
g75439 not n33911 ; n33911_not
g75440 not n42470 ; n42470_not
g75441 not n33803 ; n33803_not
g75442 not n37313 ; n37313_not
g75443 not n21923 ; n21923_not
g75444 not n53243 ; n53243_not
g75445 not n28025 ; n28025_not
g75446 not n28106 ; n28106_not
g75447 not n33722 ; n33722_not
g75448 not n35504 ; n35504_not
g75449 not n14255 ; n14255_not
g75450 not n18116 ; n18116_not
g75451 not n53315 ; n53315_not
g75452 not n33650 ; n33650_not
g75453 not n33902 ; n33902_not
g75454 not n10097 ; n10097_not
g75455 not n14516 ; n14516_not
g75456 not n28043 ; n28043_not
g75457 not n14507 ; n14507_not
g75458 not n13805 ; n13805_not
g75459 not n21932 ; n21932_not
g75460 not n45404 ; n45404_not
g75461 not n14444 ; n14444_not
g75462 not n35522 ; n35522_not
g75463 not n28205 ; n28205_not
g75464 not n26324 ; n26324_not
g75465 not n33821 ; n33821_not
g75466 not n14534 ; n14534_not
g75467 not n42353 ; n42353_not
g75468 not n21815 ; n21815_not
g75469 not n26054 ; n26054_not
g75470 not n21860 ; n21860_not
g75471 not n46610 ; n46610_not
g75472 not n28223 ; n28223_not
g75473 not n42920 ; n42920_not
g75474 not n37304 ; n37304_not
g75475 not n18134 ; n18134_not
g75476 not n10295 ; n10295_not
g75477 not n14354 ; n14354_not
g75478 not n14084 ; n14084_not
g75479 not n35261 ; n35261_not
g75480 not n31661 ; n31661_not
g75481 not n21806 ; n21806_not
g75482 not n37322 ; n37322_not
g75483 not n21842 ; n21842_not
g75484 not n14327 ; n14327_not
g75485 not n14309 ; n14309_not
g75486 not n26036 ; n26036_not
g75487 not n26063 ; n26063_not
g75488 not n25244 ; n25244_not
g75489 not n19061 ; n19061_not
g75490 not n21509 ; n21509_not
g75491 not n14093 ; n14093_not
g75492 not n53900 ; n53900_not
g75493 not n21824 ; n21824_not
g75494 not n33704 ; n33704_not
g75495 not n45008 ; n45008_not
g75496 not n14525 ; n14525_not
g75497 not n21833 ; n21833_not
g75498 not n30905 ; n30905_not
g75499 not n22139 ; n22139_not
g75500 not n10349 ; n10349_not
g75501 not n41633 ; n41633_not
g75502 not n30761 ; n30761_not
g75503 not n21851 ; n21851_not
g75504 not n28151 ; n28151_not
g75505 not n14336 ; n14336_not
g75506 not n13760 ; n13760_not
g75507 not n54134 ; n54134_not
g75508 not n45161 ; n45161_not
g75509 not n21527 ; n21527_not
g75510 not n26045 ; n26045_not
g75511 not n21383 ; n21383_not
g75512 not n38150 ; n38150_not
g75513 not n14138 ; n14138_not
g75514 not n44441 ; n44441_not
g75515 not n53225 ; n53225_not
g75516 not n26270 ; n26270_not
g75517 not n13850 ; n13850_not
g75518 not n21338 ; n21338_not
g75519 not n14282 ; n14282_not
g75520 not n48500 ; n48500_not
g75521 not n14318 ; n14318_not
g75522 not n50165 ; n50165_not
g75523 not n38204 ; n38204_not
g75524 not n55250 ; n55250_not
g75525 not n51641 ; n51641_not
g75526 not n46007 ; n46007_not
g75527 not n10277 ; n10277_not
g75528 not n28133 ; n28133_not
g75529 not n39122 ; n39122_not
g75530 not n21518 ; n21518_not
g75531 not n10286 ; n10286_not
g75532 not n14129 ; n14129_not
g75533 not n35216 ; n35216_not
g75534 not n14147 ; n14147_not
g75535 not n14066 ; n14066_not
g75536 not n38141 ; n38141_not
g75537 not n41705 ; n41705_not
g75538 not n55700 ; n55700_not
g75539 not n21482 ; n21482_not
g75540 not n53333 ; n53333_not
g75541 not n14075 ; n14075_not
g75542 not n26234 ; n26234_not
g75543 not n22094 ; n22094_not
g75544 not n26027 ; n26027_not
g75545 not n35540 ; n35540_not
g75546 not n18107 ; n18107_not
g75547 not n14291 ; n14291_not
g75548 not n55017 ; n55017_not
g75549 not n48501 ; n48501_not
g75550 not n11556 ; n11556_not
g75551 not n34920 ; n34920_not
g75552 not n41832 ; n41832_not
g75553 not n24615 ; n24615_not
g75554 not n50337 ; n50337_not
g75555 not n27036 ; n27036_not
g75556 not n17640 ; n17640_not
g75557 not n26631 ; n26631_not
g75558 not n17406 ; n17406_not
g75559 not n50607 ; n50607_not
g75560 not n24039 ; n24039_not
g75561 not n35550 ; n35550_not
g75562 not n46260 ; n46260_not
g75563 not n27441 ; n27441_not
g75564 not n27045 ; n27045_not
g75565 not n31167 ; n31167_not
g75566 not n45261 ; n45261_not
g75567 not n54351 ; n54351_not
g75568 not n44235 ; n44235_not
g75569 not n27126 ; n27126_not
g75570 not n11538 ; n11538_not
g75571 not n32049 ; n32049_not
g75572 not n46233 ; n46233_not
g75573 not n18252 ; n18252_not
g75574 not n51435 ; n51435_not
g75575 not n26640 ; n26640_not
g75576 not n44343 ; n44343_not
g75577 not n44244 ; n44244_not
g75578 not n46053 ; n46053_not
g75579 not n25812 ; n25812_not
g75580 not n51660 ; n51660_not
g75581 not n27144 ; n27144_not
g75582 not n44253 ; n44253_not
g75583 not n24606 ; n24606_not
g75584 not n56115 ; n56115_not
g75585 not n36144 ; n36144_not
g75586 not n27072 ; n27072_not
g75587 not n27027 ; n27027_not
g75588 not n52740 ; n52740_not
g75589 not n24174 ; n24174_not
g75590 not n31662 ; n31662_not
g75591 not n10683 ; n10683_not
g75592 not n50544 ; n50544_not
g75593 not n50643 ; n50643_not
g75594 not n35028 ; n35028_not
g75595 not n36126 ; n36126_not
g75596 not n24048 ; n24048_not
g75597 not n54432 ; n54432_not
g75598 not n24165 ; n24165_not
g75599 not n27234 ; n27234_not
g75600 not n57204 ; n57204_not
g75601 not n27720 ; n27720_not
g75602 not n54711 ; n54711_not
g75603 not n46413 ; n46413_not
g75604 not n54450 ; n54450_not
g75605 not n38151 ; n38151_not
g75606 not n35064 ; n35064_not
g75607 not n45252 ; n45252_not
g75608 not n46071 ; n46071_not
g75609 not n51705 ; n51705_not
g75610 not n51507 ; n51507_not
g75611 not n10476 ; n10476_not
g75612 not n45072 ; n45072_not
g75613 not n31428 ; n31428_not
g75614 not n25326 ; n25326_not
g75615 not n39501 ; n39501_not
g75616 not n57321 ; n57321_not
g75617 not n47700 ; n47700_not
g75618 not n31446 ; n31446_not
g75619 not n46440 ; n46440_not
g75620 not n11547 ; n11547_not
g75621 not n24057 ; n24057_not
g75622 not n36522 ; n36522_not
g75623 not n40194 ; n40194_not
g75624 not n45630 ; n45630_not
g75625 not n10665 ; n10665_not
g75626 not n24138 ; n24138_not
g75627 not n35532 ; n35532_not
g75628 not n40482 ; n40482_not
g75629 not n35055 ; n35055_not
g75630 not n35226 ; n35226_not
g75631 not n31419 ; n31419_not
g75632 not n51912 ; n51912_not
g75633 not n40185 ; n40185_not
g75634 not n24561 ; n24561_not
g75635 not n10647 ; n10647_not
g75636 not n24921 ; n24921_not
g75637 not n46422 ; n46422_not
g75638 not n41913 ; n41913_not
g75639 not n17820 ; n17820_not
g75640 not n28170 ; n28170_not
g75641 not n46251 ; n46251_not
g75642 not n27054 ; n27054_not
g75643 not n10638 ; n10638_not
g75644 not n34830 ; n34830_not
g75645 not n36036 ; n36036_not
g75646 not n42525 ; n42525_not
g75647 not n25344 ; n25344_not
g75648 not n50670 ; n50670_not
g75649 not n36081 ; n36081_not
g75650 not n24912 ; n24912_not
g75651 not n18270 ; n18270_not
g75652 not n43722 ; n43722_not
g75653 not n46062 ; n46062_not
g75654 not n36513 ; n36513_not
g75655 not n16740 ; n16740_not
g75656 not n27513 ; n27513_not
g75657 not n27522 ; n27522_not
g75658 not n24570 ; n24570_not
g75659 not n50661 ; n50661_not
g75660 not n50922 ; n50922_not
g75661 not n44208 ; n44208_not
g75662 not n31653 ; n31653_not
g75663 not n54720 ; n54720_not
g75664 not n51480 ; n51480_not
g75665 not n44406 ; n44406_not
g75666 not n24930 ; n24930_not
g75667 not n46305 ; n46305_not
g75668 not n10656 ; n10656_not
g75669 not n11583 ; n11583_not
g75670 not n44631 ; n44631_not
g75671 not n32139 ; n32139_not
g75672 not n51453 ; n51453_not
g75673 not n18540 ; n18540_not
g75674 not n27531 ; n27531_not
g75675 not n35046 ; n35046_not
g75676 not n27423 ; n27423_not
g75677 not n35406 ; n35406_not
g75678 not n40473 ; n40473_not
g75679 not n27405 ; n27405_not
g75680 not n46242 ; n46242_not
g75681 not n17073 ; n17073_not
g75682 not n36054 ; n36054_not
g75683 not n42516 ; n42516_not
g75684 not n27081 ; n27081_not
g75685 not n31734 ; n31734_not
g75686 not n44262 ; n44262_not
g75687 not n36063 ; n36063_not
g75688 not n45333 ; n45333_not
g75689 not n24129 ; n24129_not
g75690 not n48411 ; n48411_not
g75691 not n51606 ; n51606_not
g75692 not n31608 ; n31608_not
g75693 not n36108 ; n36108_not
g75694 not n26172 ; n26172_not
g75695 not n32148 ; n32148_not
g75696 not n43713 ; n43713_not
g75697 not n24156 ; n24156_not
g75698 not n24075 ; n24075_not
g75699 not n40464 ; n40464_not
g75700 not n35523 ; n35523_not
g75701 not n27540 ; n27540_not
g75702 not n10629 ; n10629_not
g75703 not n35037 ; n35037_not
g75704 not n44532 ; n44532_not
g75705 not n10674 ; n10674_not
g75706 not n36315 ; n36315_not
g75707 not n41814 ; n41814_not
g75708 not n44190 ; n44190_not
g75709 not n51462 ; n51462_not
g75710 not n27504 ; n27504_not
g75711 not n50652 ; n50652_not
g75712 not n50526 ; n50526_not
g75713 not n10467 ; n10467_not
g75714 not n24066 ; n24066_not
g75715 not n26226 ; n26226_not
g75716 not n27432 ; n27432_not
g75717 not n28314 ; n28314_not
g75718 not n35217 ; n35217_not
g75719 not n40149 ; n40149_not
g75720 not n31617 ; n31617_not
g75721 not n11592 ; n11592_not
g75722 not n28701 ; n28701_not
g75723 not n46314 ; n46314_not
g75724 not n50913 ; n50913_not
g75725 not n27117 ; n27117_not
g75726 not n18261 ; n18261_not
g75727 not n52731 ; n52731_not
g75728 not n25821 ; n25821_not
g75729 not n44316 ; n44316_not
g75730 not n18144 ; n18144_not
g75731 not n41841 ; n41841_not
g75732 not n54441 ; n54441_not
g75733 not n36045 ; n36045_not
g75734 not n45720 ; n45720_not
g75735 not n56043 ; n56043_not
g75736 not n44721 ; n44721_not
g75737 not n31455 ; n31455_not
g75738 not n51444 ; n51444_not
g75739 not n25335 ; n25335_not
g75740 not n27702 ; n27702_not
g75741 not n27414 ; n27414_not
g75742 not n24147 ; n24147_not
g75743 not n24903 ; n24903_not
g75744 not n25830 ; n25830_not
g75745 not n17082 ; n17082_not
g75746 not n46431 ; n46431_not
g75747 not n44640 ; n44640_not
g75748 not n24093 ; n24093_not
g75749 not n44217 ; n44217_not
g75750 not n47232 ; n47232_not
g75751 not n40491 ; n40491_not
g75752 not n44226 ; n44226_not
g75753 not n57222 ; n57222_not
g75754 not n45711 ; n45711_not
g75755 not n35541 ; n35541_not
g75756 not n40158 ; n40158_not
g75757 not n26217 ; n26217_not
g75758 not n16731 ; n16731_not
g75759 not n36324 ; n36324_not
g75760 not n24084 ; n24084_not
g75761 not n44307 ; n44307_not
g75762 not n31806 ; n31806_not
g75763 not n26181 ; n26181_not
g75764 not n50616 ; n50616_not
g75765 not n52713 ; n52713_not
g75766 not n44622 ; n44622_not
g75767 not n24651 ; n24651_not
g75768 not n27180 ; n27180_not
g75769 not n26064 ; n26064_not
g75770 not n52812 ; n52812_not
g75771 not n36207 ; n36207_not
g75772 not n49302 ; n49302_not
g75773 not n18171 ; n18171_not
g75774 not n36801 ; n36801_not
g75775 not n24660 ; n24660_not
g75776 not n27261 ; n27261_not
g75777 not n26442 ; n26442_not
g75778 not n51363 ; n51363_not
g75779 not n39033 ; n39033_not
g75780 not n28071 ; n28071_not
g75781 not n46323 ; n46323_not
g75782 not n26541 ; n26541_not
g75783 not n17109 ; n17109_not
g75784 not n10278 ; n10278_not
g75785 not n51831 ; n51831_not
g75786 not n46008 ; n46008_not
g75787 not n10872 ; n10872_not
g75788 not n17334 ; n17334_not
g75789 not n50193 ; n50193_not
g75790 not n26460 ; n26460_not
g75791 not n24633 ; n24633_not
g75792 not n39420 ; n39420_not
g75793 not n27171 ; n27171_not
g75794 not n46332 ; n46332_not
g75795 not n51354 ; n51354_not
g75796 not n17325 ; n17325_not
g75797 not n27306 ; n27306_not
g75798 not n52821 ; n52821_not
g75799 not n10449 ; n10449_not
g75800 not n17730 ; n17730_not
g75801 not n42471 ; n42471_not
g75802 not n18207 ; n18207_not
g75803 not n54171 ; n54171_not
g75804 not n31374 ; n31374_not
g75805 not n10287 ; n10287_not
g75806 not n26451 ; n26451_not
g75807 not n50571 ; n50571_not
g75808 not n36225 ; n36225_not
g75809 not n40581 ; n40581_not
g75810 not n36216 ; n36216_not
g75811 not n11448 ; n11448_not
g75812 not n27270 ; n27270_not
g75813 not n54405 ; n54405_not
g75814 not n18216 ; n18216_not
g75815 not n37026 ; n37026_not
g75816 not n31644 ; n31644_not
g75817 not n36603 ; n36603_not
g75818 not n26415 ; n26415_not
g75819 not n52443 ; n52443_not
g75820 not n36351 ; n36351_not
g75821 not n44703 ; n44703_not
g75822 not n26082 ; n26082_not
g75823 not n57420 ; n57420_not
g75824 not n21267 ; n21267_not
g75825 not n51390 ; n51390_not
g75826 not n10494 ; n10494_not
g75827 not n31383 ; n31383_not
g75828 not n11457 ; n11457_not
g75829 not n35442 ; n35442_not
g75830 not n26406 ; n26406_not
g75831 not n46026 ; n46026_not
g75832 not n50580 ; n50580_not
g75833 not n26433 ; n26433_not
g75834 not n51372 ; n51372_not
g75835 not n28215 ; n28215_not
g75836 not n26550 ; n26550_not
g75837 not n38610 ; n38610_not
g75838 not n40572 ; n40572_not
g75839 not n44820 ; n44820_not
g75840 not n35451 ; n35451_not
g75841 not n32175 ; n32175_not
g75842 not n39024 ; n39024_not
g75843 not n37035 ; n37035_not
g75844 not n54261 ; n54261_not
g75845 not n31671 ; n31671_not
g75846 not n26424 ; n26424_not
g75847 not n51381 ; n51381_not
g75848 not n10269 ; n10269_not
g75849 not n41823 ; n41823_not
g75850 not n52803 ; n52803_not
g75851 not n42615 ; n42615_not
g75852 not n28242 ; n28242_not
g75853 not n18720 ; n18720_not
g75854 not n54612 ; n54612_not
g75855 not n27342 ; n27342_not
g75856 not n25254 ; n25254_not
g75857 not n11907 ; n11907_not
g75858 not n26037 ; n26037_not
g75859 not n50562 ; n50562_not
g75860 not n11916 ; n11916_not
g75861 not n34551 ; n34551_not
g75862 not n17307 ; n17307_not
g75863 not n11925 ; n11925_not
g75864 not n45090 ; n45090_not
g75865 not n39411 ; n39411_not
g75866 not n46350 ; n46350_not
g75867 not n11934 ; n11934_not
g75868 not n34542 ; n34542_not
g75869 not n31743 ; n31743_not
g75870 not n10386 ; n10386_not
g75871 not n11943 ; n11943_not
g75872 not n51336 ; n51336_not
g75873 not n11952 ; n11952_not
g75874 not n26523 ; n26523_not
g75875 not n50535 ; n50535_not
g75876 not n46341 ; n46341_not
g75877 not n24543 ; n24543_not
g75878 not n25245 ; n25245_not
g75879 not n26505 ; n26505_not
g75880 not n48150 ; n48150_not
g75881 not n51327 ; n51327_not
g75882 not n27360 ; n27360_not
g75883 not n26028 ; n26028_not
g75884 not n36810 ; n36810_not
g75885 not n47241 ; n47241_not
g75886 not n27351 ; n27351_not
g75887 not n17127 ; n17127_not
g75888 not n39402 ; n39402_not
g75889 not n34560 ; n34560_not
g75890 not n26514 ; n26514_not
g75891 not n17703 ; n17703_not
g75892 not n36360 ; n36360_not
g75893 not n10377 ; n10377_not
g75894 not n42480 ; n42480_not
g75895 not n10359 ; n10359_not
g75896 not n26019 ; n26019_not
g75897 not n37800 ; n37800_not
g75898 not n27324 ; n27324_not
g75899 not n54126 ; n54126_not
g75900 not n35262 ; n35262_not
g75901 not n34911 ; n34911_not
g75902 not n27135 ; n27135_not
g75903 not n31752 ; n31752_not
g75904 not n28080 ; n28080_not
g75905 not n46017 ; n46017_not
g75906 not n26532 ; n26532_not
g75907 not n17316 ; n17316_not
g75908 not n27315 ; n27315_not
g75909 not n51534 ; n51534_not
g75910 not n37053 ; n37053_not
g75911 not n10296 ; n10296_not
g75912 not n40095 ; n40095_not
g75913 not n40590 ; n40590_not
g75914 not n31365 ; n31365_not
g75915 not n34533 ; n34533_not
g75916 not n27333 ; n27333_not
g75917 not n44361 ; n44361_not
g75918 not n18180 ; n18180_not
g75919 not n11961 ; n11961_not
g75920 not n55035 ; n55035_not
g75921 not n35460 ; n35460_not
g75922 not n25236 ; n25236_not
g75923 not n50553 ; n50553_not
g75924 not n35271 ; n35271_not
g75925 not n34524 ; n34524_not
g75926 not n34902 ; n34902_not
g75927 not n17910 ; n17910_not
g75928 not n51345 ; n51345_not
g75929 not n17118 ; n17118_not
g75930 not n32184 ; n32184_not
g75931 not n34146 ; n34146_not
g75932 not n27162 ; n27162_not
g75933 not n27243 ; n27243_not
g75934 not n26046 ; n26046_not
g75935 not n54603 ; n54603_not
g75936 not n48420 ; n48420_not
g75937 not n10098 ; n10098_not
g75938 not n42624 ; n42624_not
g75939 not n26136 ; n26136_not
g75940 not n27450 ; n27450_not
g75941 not n25920 ; n25920_not
g75942 not n24804 ; n24804_not
g75943 not n10089 ; n10089_not
g75944 not n50625 ; n50625_not
g75945 not n16713 ; n16713_not
g75946 not n35424 ; n35424_not
g75947 not n56061 ; n56061_not
g75948 not n26604 ; n26604_not
g75949 not n52470 ; n52470_not
g75950 not n40518 ; n40518_not
g75951 not n44712 ; n44712_not
g75952 not n48231 ; n48231_not
g75953 not n10584 ; n10584_not
g75954 not n51417 ; n51417_not
g75955 not n51570 ; n51570_not
g75956 not n24813 ; n24813_not
g75957 not n51408 ; n51408_not
g75958 not n51561 ; n51561_not
g75959 not n36153 ; n36153_not
g75960 not n40527 ; n40527_not
g75961 not n16704 ; n16704_not
g75962 not n47520 ; n47520_not
g75963 not n35505 ; n35505_not
g75964 not n45081 ; n45081_not
g75965 not n28152 ; n28152_not
g75966 not n47331 ; n47331_not
g75967 not n26127 ; n26127_not
g75968 not n10575 ; n10575_not
g75969 not n44523 ; n44523_not
g75970 not n31680 ; n31680_not
g75971 not n36333 ; n36333_not
g75972 not n17361 ; n17361_not
g75973 not n27612 ; n27612_not
g75974 not n10593 ; n10593_not
g75975 not n50634 ; n50634_not
g75976 not n54180 ; n54180_not
g75977 not n27630 ; n27630_not
g75978 not n25902 ; n25902_not
g75979 not n18153 ; n18153_not
g75980 not n35019 ; n35019_not
g75981 not n40077 ; n40077_not
g75982 not n48240 ; n48240_not
g75983 not n24624 ; n24624_not
g75984 not n17712 ; n17712_not
g75985 not n54270 ; n54270_not
g75986 not n24840 ; n24840_not
g75987 not n10485 ; n10485_not
g75988 not n51426 ; n51426_not
g75989 not n51813 ; n51813_not
g75990 not n26622 ; n26622_not
g75991 not n35514 ; n35514_not
g75992 not n26154 ; n26154_not
g75993 not n35415 ; n35415_not
g75994 not n40167 ; n40167_not
g75995 not n16722 ; n16722_not
g75996 not n40509 ; n40509_not
g75997 not n57330 ; n57330_not
g75998 not n54423 ; n54423_not
g75999 not n25911 ; n25911_not
g76000 not n18243 ; n18243_not
g76001 not n49320 ; n49320_not
g76002 not n17901 ; n17901_not
g76003 not n24822 ; n24822_not
g76004 not n27090 ; n27090_not
g76005 not n51516 ; n51516_not
g76006 not n39060 ; n39060_not
g76007 not n56052 ; n56052_not
g76008 not n26613 ; n26613_not
g76009 not n32157 ; n32157_not
g76010 not n46800 ; n46800_not
g76011 not n31626 ; n31626_not
g76012 not n50166 ; n50166_not
g76013 not n17370 ; n17370_not
g76014 not n46044 ; n46044_not
g76015 not n24831 ; n24831_not
g76016 not n24732 ; n24732_not
g76017 not n49500 ; n49500_not
g76018 not n10539 ; n10539_not
g76019 not n23922 ; n23922_not
g76020 not n44271 ; n44271_not
g76021 not n37008 ; n37008_not
g76022 not n40554 ; n40554_not
g76023 not n36612 ; n36612_not
g76024 not n31149 ; n31149_not
g76025 not n10188 ; n10188_not
g76026 not n24741 ; n24741_not
g76027 not n28044 ; n28044_not
g76028 not n23931 ; n23931_not
g76029 not n57402 ; n57402_not
g76030 not n36342 ; n36342_not
g76031 not n10179 ; n10179_not
g76032 not n17352 ; n17352_not
g76033 not n28251 ; n28251_not
g76034 not n31158 ; n31158_not
g76035 not n24750 ; n24750_not
g76036 not n40563 ; n40563_not
g76037 not n44280 ; n44280_not
g76038 not n17343 ; n17343_not
g76039 not n24714 ; n24714_not
g76040 not n51543 ; n51543_not
g76041 not n23904 ; n23904_not
g76042 not n18711 ; n18711_not
g76043 not n26091 ; n26091_not
g76044 not n11466 ; n11466_not
g76045 not n27252 ; n27252_not
g76046 not n35253 ; n35253_not
g76047 not n44433 ; n44433_not
g76048 not n51822 ; n51822_not
g76049 not n24723 ; n24723_not
g76050 not n45306 ; n45306_not
g76051 not n52452 ; n52452_not
g76052 not n23913 ; n23913_not
g76053 not n57411 ; n57411_not
g76054 not n18504 ; n18504_not
g76055 not n36900 ; n36900_not
g76056 not n18225 ; n18225_not
g76057 not n10197 ; n10197_not
g76058 not n25281 ; n25281_not
g76059 not n27207 ; n27207_not
g76060 not n46035 ; n46035_not
g76061 not n31635 ; n31635_not
g76062 not n48213 ; n48213_not
g76063 not n54360 ; n54360_not
g76064 not n26361 ; n26361_not
g76065 not n36171 ; n36171_not
g76066 not n28260 ; n28260_not
g76067 not n27216 ; n27216_not
g76068 not n40536 ; n40536_not
g76069 not n47511 ; n47511_not
g76070 not n31392 ; n31392_not
g76071 not n54414 ; n54414_not
g76072 not n45540 ; n45540_not
g76073 not n10566 ; n10566_not
g76074 not n48222 ; n48222_not
g76075 not n35433 ; n35433_not
g76076 not n11493 ; n11493_not
g76077 not n18234 ; n18234_not
g76078 not n39015 ; n39015_not
g76079 not n44514 ; n44514_not
g76080 not n10548 ; n10548_not
g76081 not n32166 ; n32166_not
g76082 not n23940 ; n23940_not
g76083 not n48204 ; n48204_not
g76084 not n18702 ; n18702_not
g76085 not n26109 ; n26109_not
g76086 not n18162 ; n18162_not
g76087 not n18513 ; n18513_not
g76088 not n51525 ; n51525_not
g76089 not n40545 ; n40545_not
g76090 not n52425 ; n52425_not
g76091 not n10557 ; n10557_not
g76092 not n45216 ; n45216_not
g76093 not n54621 ; n54621_not
g76094 not n25290 ; n25290_not
g76095 not n47502 ; n47502_not
g76096 not n51552 ; n51552_not
g76097 not n36162 ; n36162_not
g76098 not n26325 ; n26325_not
g76099 not n26730 ; n26730_not
g76100 not n44046 ; n44046_not
g76101 not n36252 ; n36252_not
g76102 not n42435 ; n42435_not
g76103 not n18045 ; n18045_not
g76104 not n10845 ; n10845_not
g76105 not n39222 ; n39222_not
g76106 not n52650 ; n52650_not
g76107 not n42561 ; n42561_not
g76108 not n25371 ; n25371_not
g76109 not n25641 ; n25641_not
g76110 not n27810 ; n27810_not
g76111 not n26721 ; n26721_not
g76112 not n25461 ; n25461_not
g76113 not n32076 ; n32076_not
g76114 not n31563 ; n31563_not
g76115 not n25380 ; n25380_not
g76116 not n26316 ; n26316_not
g76117 not n31572 ; n31572_not
g76118 not n35127 ; n35127_not
g76119 not n35136 ; n35136_not
g76120 not n17514 ; n17514_not
g76121 not n25353 ; n25353_not
g76122 not n25650 ; n25650_not
g76123 not n36234 ; n36234_not
g76124 not n44055 ; n44055_not
g76125 not n36243 ; n36243_not
g76126 not n11088 ; n11088_not
g76127 not n26910 ; n26910_not
g76128 not n26901 ; n26901_not
g76129 not n36414 ; n36414_not
g76130 not n18027 ; n18027_not
g76131 not n46530 ; n46530_not
g76132 not n46170 ; n46170_not
g76133 not n51183 ; n51183_not
g76134 not n54540 ; n54540_not
g76135 not n42606 ; n42606_not
g76136 not n45603 ; n45603_not
g76137 not n39231 ; n39231_not
g76138 not n54522 ; n54522_not
g76139 not n18036 ; n18036_not
g76140 not n51192 ; n51192_not
g76141 not n17523 ; n17523_not
g76142 not n46080 ; n46080_not
g76143 not n45450 ; n45450_not
g76144 not n35235 ; n35235_not
g76145 not n36270 ; n36270_not
g76146 not n51228 ; n51228_not
g76147 not n28521 ; n28521_not
g76148 not n26307 ; n26307_not
g76149 not n51237 ; n51237_not
g76150 not n18072 ; n18072_not
g76151 not n44028 ; n44028_not
g76152 not n26190 ; n26190_not
g76153 not n45810 ; n45810_not
g76154 not n25623 ; n25623_not
g76155 not n48600 ; n48600_not
g76156 not n45315 ; n45315_not
g76157 not n49104 ; n49104_not
g76158 not n17541 ; n17541_not
g76159 not n31509 ; n31509_not
g76160 not n25416 ; n25416_not
g76161 not n18081 ; n18081_not
g76162 not n45441 ; n45441_not
g76163 not n25470 ; n25470_not
g76164 not n35352 ; n35352_not
g76165 not n18063 ; n18063_not
g76166 not n44037 ; n44037_not
g76167 not n45801 ; n45801_not
g76168 not n26712 ; n26712_not
g76169 not n18054 ; n18054_not
g76170 not n46107 ; n46107_not
g76171 not n51750 ; n51750_not
g76172 not n25632 ; n25632_not
g76173 not n35118 ; n35118_not
g76174 not n27603 ; n27603_not
g76175 not n46161 ; n46161_not
g76176 not n36261 ; n36261_not
g76177 not n17532 ; n17532_not
g76178 not n51219 ; n51219_not
g76179 not n36504 ; n36504_not
g76180 not n26703 ; n26703_not
g76181 not n18108 ; n18108_not
g76182 not n54225 ; n54225_not
g76183 not n45900 ; n45900_not
g76184 not n40392 ; n40392_not
g76185 not n31581 ; n31581_not
g76186 not n35109 ; n35109_not
g76187 not n17604 ; n17604_not
g76188 not n35172 ; n35172_not
g76189 not n45207 ; n45207_not
g76190 not n49131 ; n49131_not
g76191 not n11187 ; n11187_not
g76192 not n51903 ; n51903_not
g76193 not n52560 ; n52560_not
g76194 not n46116 ; n46116_not
g76195 not n40293 ; n40293_not
g76196 not n18522 ; n18522_not
g76197 not n31491 ; n31491_not
g76198 not n35163 ; n35163_not
g76199 not n11178 ; n11178_not
g76200 not n47313 ; n47313_not
g76201 not n10818 ; n10818_not
g76202 not n54306 ; n54306_not
g76203 not n25308 ; n25308_not
g76204 not n45513 ; n45513_not
g76205 not n46215 ; n46215_not
g76206 not n17019 ; n17019_not
g76207 not n54513 ; n54513_not
g76208 not n11169 ; n11169_not
g76209 not n27711 ; n27711_not
g76210 not n35640 ; n35640_not
g76211 not n26802 ; n26802_not
g76212 not n36450 ; n36450_not
g76213 not n51732 ; n51732_not
g76214 not n46224 ; n46224_not
g76215 not n37512 ; n37512_not
g76216 not n49122 ; n49122_not
g76217 not n44073 ; n44073_not
g76218 not n10809 ; n10809_not
g76219 not n35703 ; n35703_not
g76220 not n54504 ; n54504_not
g76221 not n51129 ; n51129_not
g76222 not n50832 ; n50832_not
g76223 not n11196 ; n11196_not
g76224 not n45522 ; n45522_not
g76225 not n27801 ; n27801_not
g76226 not n48321 ; n48321_not
g76227 not n27900 ; n27900_not
g76228 not n46710 ; n46710_not
g76229 not n51156 ; n51156_not
g76230 not n18360 ; n18360_not
g76231 not n10827 ; n10827_not
g76232 not n35145 ; n35145_not
g76233 not n18009 ; n18009_not
g76234 not n32085 ; n32085_not
g76235 not n51165 ; n51165_not
g76236 not n49203 ; n49203_not
g76237 not n46206 ; n46206_not
g76238 not n35721 ; n35721_not
g76239 not n11097 ; n11097_not
g76240 not n10836 ; n10836_not
g76241 not n54135 ; n54135_not
g76242 not n31707 ; n31707_not
g76243 not n39240 ; n39240_not
g76244 not n51174 ; n51174_not
g76245 not n18018 ; n18018_not
g76246 not n51615 ; n51615_not
g76247 not n51147 ; n51147_not
g76248 not n50760 ; n50760_not
g76249 not n45504 ; n45504_not
g76250 not n41931 ; n41931_not
g76251 not n44064 ; n44064_not
g76252 not n26145 ; n26145_not
g76253 not n35712 ; n35712_not
g76254 not n45225 ; n45225_not
g76255 not n51723 ; n51723_not
g76256 not n35154 ; n35154_not
g76257 not n49140 ; n49140_not
g76258 not n17505 ; n17505_not
g76259 not n35208 ; n35208_not
g76260 not n28008 ; n28008_not
g76261 not n50814 ; n50814_not
g76262 not n26280 ; n26280_not
g76263 not n48330 ; n48330_not
g76264 not n40239 ; n40239_not
g76265 not n36432 ; n36432_not
g76266 not n51309 ; n51309_not
g76267 not n25524 ; n25524_not
g76268 not n40338 ; n40338_not
g76269 not n39150 ; n39150_not
g76270 not n49221 ; n49221_not
g76271 not n45360 ; n45360_not
g76272 not n35730 ; n35730_not
g76273 not n31536 ; n31536_not
g76274 not n18090 ; n18090_not
g76275 not n49113 ; n49113_not
g76276 not n51291 ; n51291_not
g76277 not n16911 ; n16911_not
g76278 not n36441 ; n36441_not
g76279 not n45270 ; n45270_not
g76280 not n46602 ; n46602_not
g76281 not n49212 ; n49212_not
g76282 not n54234 ; n54234_not
g76283 not n10944 ; n10944_not
g76284 not n25506 ; n25506_not
g76285 not n52605 ; n52605_not
g76286 not n26235 ; n26235_not
g76287 not n36405 ; n36405_not
g76288 not n35325 ; n35325_not
g76289 not n25515 ; n25515_not
g76290 not n10935 ; n10935_not
g76291 not n32058 ; n32058_not
g76292 not n18405 ; n18405_not
g76293 not n35307 ; n35307_not
g76294 not n45342 ; n45342_not
g76295 not n17802 ; n17802_not
g76296 not n38520 ; n38520_not
g76297 not n25560 ; n25560_not
g76298 not n26262 ; n26262_not
g76299 not n28431 ; n28431_not
g76300 not n40347 ; n40347_not
g76301 not n26271 ; n26271_not
g76302 not n18414 ; n18414_not
g76303 not n31545 ; n31545_not
g76304 not n10890 ; n10890_not
g76305 not n54900 ; n54900_not
g76306 not n45351 ; n45351_not
g76307 not n46521 ; n46521_not
g76308 not n46125 ; n46125_not
g76309 not n25542 ; n25542_not
g76310 not n51318 ; n51318_not
g76311 not n40356 ; n40356_not
g76312 not n56700 ; n56700_not
g76313 not n10917 ; n10917_not
g76314 not n45324 ; n45324_not
g76315 not n47223 ; n47223_not
g76316 not n54090 ; n54090_not
g76317 not n16920 ; n16920_not
g76318 not n25551 ; n25551_not
g76319 not n36621 ; n36621_not
g76320 not n51255 ; n51255_not
g76321 not n25443 ; n25443_not
g76322 not n52623 ; n52623_not
g76323 not n10980 ; n10980_not
g76324 not n35073 ; n35073_not
g76325 not n36531 ; n36531_not
g76326 not n40383 ; n40383_not
g76327 not n35343 ; n35343_not
g76328 not n49230 ; n49230_not
g76329 not n45423 ; n45423_not
g76330 not n39114 ; n39114_not
g76331 not n17550 ; n17550_not
g76332 not n45414 ; n45414_not
g76333 not n39204 ; n39204_not
g76334 not n51840 ; n51840_not
g76335 not n42570 ; n42570_not
g76336 not n39132 ; n39132_not
g76337 not n10854 ; n10854_not
g76338 not n35091 ; n35091_not
g76339 not n51246 ; n51246_not
g76340 not n52632 ; n52632_not
g76341 not n39213 ; n39213_not
g76342 not n25425 ; n25425_not
g76343 not n31554 ; n31554_not
g76344 not n27621 ; n27621_not
g76345 not n46503 ; n46503_not
g76346 not n31590 ; n31590_not
g76347 not n28413 ; n28413_not
g76348 not n31518 ; n31518_not
g76349 not n35082 ; n35082_not
g76350 not n42453 ; n42453_not
g76351 not n39105 ; n39105_not
g76352 not n44019 ; n44019_not
g76353 not n46152 ; n46152_not
g76354 not n31716 ; n31716_not
g76355 not n45432 ; n45432_not
g76356 not n18450 ; n18450_not
g76357 not n25614 ; n25614_not
g76358 not n28503 ; n28503_not
g76359 not n18126 ; n18126_not
g76360 not n51282 ; n51282_not
g76361 not n36306 ; n36306_not
g76362 not n40248 ; n40248_not
g76363 not n50805 ; n50805_not
g76364 not n40329 ; n40329_not
g76365 not n10962 ; n10962_not
g76366 not n36423 ; n36423_not
g76367 not n46512 ; n46512_not
g76368 not n46134 ; n46134_not
g76369 not n40365 ; n40365_not
g76370 not n44541 ; n44541_not
g76371 not n18432 ; n18432_not
g76372 not n44802 ; n44802_not
g76373 not n18135 ; n18135_not
g76374 not n50823 ; n50823_not
g76375 not n35280 ; n35280_not
g76376 not n31527 ; n31527_not
g76377 not n51264 ; n51264_not
g76378 not n45405 ; n45405_not
g76379 not n25605 ; n25605_not
g76380 not n51273 ; n51273_not
g76381 not n40374 ; n40374_not
g76382 not n18117 ; n18117_not
g76383 not n16902 ; n16902_not
g76384 not n54531 ; n54531_not
g76385 not n46143 ; n46143_not
g76386 not n42543 ; n42543_not
g76387 not n24264 ; n24264_not
g76388 not n49032 ; n49032_not
g76389 not n10737 ; n10737_not
g76390 not n40437 ; n40437_not
g76391 not n44730 ; n44730_not
g76392 not n44136 ; n44136_not
g76393 not n25083 ; n25083_not
g76394 not n39312 ; n39312_not
g76395 not n28125 ; n28125_not
g76396 not n24273 ; n24273_not
g76397 not n50715 ; n50715_not
g76398 not n49023 ; n49023_not
g76399 not n24480 ; n24480_not
g76400 not n17433 ; n17433_not
g76401 not n57105 ; n57105_not
g76402 not n25092 ; n25092_not
g76403 not n24282 ; n24282_not
g76404 not n35181 ; n35181_not
g76405 not n56007 ; n56007_not
g76406 not n10728 ; n10728_not
g76407 not n42417 ; n42417_not
g76408 not n36117 ; n36117_not
g76409 not n11475 ; n11475_not
g76410 not n57123 ; n57123_not
g76411 not n25065 ; n25065_not
g76412 not n50706 ; n50706_not
g76413 not n24255 ; n24255_not
g76414 not n34803 ; n34803_not
g76415 not n18603 ; n18603_not
g76416 not n54144 ; n54144_not
g76417 not n49014 ; n49014_not
g76418 not n25074 ; n25074_not
g76419 not n57114 ; n57114_not
g76420 not n36720 ; n36720_not
g76421 not n52533 ; n52533_not
g76422 not n51471 ; n51471_not
g76423 not n45621 ; n45621_not
g76424 not n10755 ; n10755_not
g76425 not n25119 ; n25119_not
g76426 not n11376 ; n11376_not
g76427 not n24309 ; n24309_not
g76428 not n40428 ; n40428_not
g76429 not n10395 ; n10395_not
g76430 not n44118 ; n44118_not
g76431 not n11367 ; n11367_not
g76432 not n25128 ; n25128_not
g76433 not n36711 ; n36711_not
g76434 not n54810 ; n54810_not
g76435 not n10746 ; n10746_not
g76436 not n44127 ; n44127_not
g76437 not n49041 ; n49041_not
g76438 not n44451 ; n44451_not
g76439 not n45036 ; n45036_not
g76440 not n24291 ; n24291_not
g76441 not n11394 ; n11394_not
g76442 not n28341 ; n28341_not
g76443 not n17442 ; n17442_not
g76444 not n39303 ; n39303_not
g76445 not n54630 ; n54630_not
g76446 not n24471 ; n24471_not
g76447 not n11385 ; n11385_not
g76448 not n28116 ; n28116_not
g76449 not n54702 ; n54702_not
g76450 not n35622 ; n35622_not
g76451 not n44424 ; n44424_not
g76452 not n24525 ; n24525_not
g76453 not n52515 ; n52515_not
g76454 not n39510 ; n39510_not
g76455 not n35631 ; n35631_not
g76456 not n47322 ; n47322_not
g76457 not n39330 ; n39330_not
g76458 not n51642 ; n51642_not
g76459 not n17415 ; n17415_not
g76460 not n48510 ; n48510_not
g76461 not n40446 ; n40446_not
g76462 not n45027 ; n45027_not
g76463 not n44181 ; n44181_not
g76464 not n40455 ; n40455_not
g76465 not n44613 ; n44613_not
g76466 not n28323 ; n28323_not
g76467 not n25803 ; n25803_not
g76468 not n24183 ; n24183_not
g76469 not n11628 ; n11628_not
g76470 not n27009 ; n27009_not
g76471 not n10692 ; n10692_not
g76472 not n54801 ; n54801_not
g76473 not n17064 ; n17064_not
g76474 not n18630 ; n18630_not
g76475 not n24534 ; n24534_not
g76476 not n26244 ; n26244_not
g76477 not n44172 ; n44172_not
g76478 not n24192 ; n24192_not
g76479 not n28332 ; n28332_not
g76480 not n44154 ; n44154_not
g76481 not n49005 ; n49005_not
g76482 not n31464 ; n31464_not
g76483 not n50904 ; n50904_not
g76484 not n25047 ; n25047_not
g76485 not n57132 ; n57132_not
g76486 not n38700 ; n38700_not
g76487 not n24237 ; n24237_not
g76488 not n46701 ; n46701_not
g76489 not n18612 ; n18612_not
g76490 not n39321 ; n39321_not
g76491 not n28035 ; n28035_not
g76492 not n25056 ; n25056_not
g76493 not n24246 ; n24246_not
g76494 not n17424 ; n17424_not
g76495 not n18306 ; n18306_not
g76496 not n44145 ; n44145_not
g76497 not n11565 ; n11565_not
g76498 not n57150 ; n57150_not
g76499 not n37503 ; n37503_not
g76500 not n28026 ; n28026_not
g76501 not n24516 ; n24516_not
g76502 not n25029 ; n25029_not
g76503 not n18621 ; n18621_not
g76504 not n24219 ; n24219_not
g76505 not n44163 ; n44163_not
g76506 not n44604 ; n44604_not
g76507 not n45612 ; n45612_not
g76508 not n25038 ; n25038_not
g76509 not n28143 ; n28143_not
g76510 not n24228 ; n24228_not
g76511 not n10719 ; n10719_not
g76512 not n48402 ; n48402_not
g76513 not n11268 ; n11268_not
g76514 not n17037 ; n17037_not
g76515 not n10953 ; n10953_not
g76516 not n25218 ; n25218_not
g76517 not n24408 ; n24408_not
g76518 not n44091 ; n44091_not
g76519 not n57033 ; n57033_not
g76520 not n41922 ; n41922_not
g76521 not n11259 ; n11259_not
g76522 not n42426 ; n42426_not
g76523 not n25227 ; n25227_not
g76524 not n18342 ; n18342_not
g76525 not n11286 ; n11286_not
g76526 not n16812 ; n16812_not
g76527 not n26811 ; n26811_not
g76528 not n26352 ; n26352_not
g76529 not n35370 ; n35370_not
g76530 not n24390 ; n24390_not
g76531 not n11277 ; n11277_not
g76532 not n10782 ; n10782_not
g76533 not n31473 ; n31473_not
g76534 not n25704 ; n25704_not
g76535 not n54216 ; n54216_not
g76536 not n54315 ; n54315_not
g76537 not n57042 ; n57042_not
g76538 not n26820 ; n26820_not
g76539 not n25209 ; n25209_not
g76540 not n44811 ; n44811_not
g76541 not n47601 ; n47601_not
g76542 not n47610 ; n47610_not
g76543 not n40419 ; n40419_not
g76544 not n44082 ; n44082_not
g76545 not n35190 ; n35190_not
g76546 not n25263 ; n25263_not
g76547 not n32094 ; n32094_not
g76548 not n16830 ; n16830_not
g76549 not n50751 ; n50751_not
g76550 not n40284 ; n40284_not
g76551 not n25434 ; n25434_not
g76552 not n16821 ; n16821_not
g76553 not n28053 ; n28053_not
g76554 not n42633 ; n42633_not
g76555 not n44442 ; n44442_not
g76556 not n17028 ; n17028_not
g76557 not n10791 ; n10791_not
g76558 not n39123 ; n39123_not
g76559 not n48312 ; n48312_not
g76560 not n36072 ; n36072_not
g76561 not n45531 ; n45531_not
g76562 not n49410 ; n49410_not
g76563 not n40275 ; n40275_not
g76564 not n57006 ; n57006_not
g76565 not n51741 ; n51741_not
g76566 not n50742 ; n50742_not
g76567 not n35361 ; n35361_not
g76568 not n51651 ; n51651_not
g76569 not n10908 ; n10908_not
g76570 not n25146 ; n25146_not
g76571 not n10764 ; n10764_not
g76572 not n24336 ; n24336_not
g76573 not n49050 ; n49050_not
g76574 not n43704 ; n43704_not
g76575 not n25731 ; n25731_not
g76576 not n25155 ; n25155_not
g76577 not n56016 ; n56016_not
g76578 not n24345 ; n24345_not
g76579 not n26334 ; n26334_not
g76580 not n42642 ; n42642_not
g76581 not n16803 ; n16803_not
g76582 not n35316 ; n35316_not
g76583 not n45045 ; n45045_not
g76584 not n25740 ; n25740_not
g76585 not n24318 ; n24318_not
g76586 not n28224 ; n28224_not
g76587 not n28107 ; n28107_not
g76588 not n11358 ; n11358_not
g76589 not n25137 ; n25137_not
g76590 not n50724 ; n50724_not
g76591 not n24327 ; n24327_not
g76592 not n44109 ; n44109_not
g76593 not n17631 ; n17631_not
g76594 not n17451 ; n17451_not
g76595 not n11349 ; n11349_not
g76596 not n40257 ; n40257_not
g76597 not n52542 ; n52542_not
g76598 not n17622 ; n17622_not
g76599 not n28350 ; n28350_not
g76600 not n25182 ; n25182_not
g76601 not n10773 ; n10773_not
g76602 not n24372 ; n24372_not
g76603 not n25713 ; n25713_not
g76604 not n11295 ; n11295_not
g76605 not n50733 ; n50733_not
g76606 not n24426 ; n24426_not
g76607 not n25191 ; n25191_not
g76608 not n24381 ; n24381_not
g76609 not n57051 ; n57051_not
g76610 not n50157 ; n50157_not
g76611 not n31761 ; n31761_not
g76612 not n39042 ; n39042_not
g76613 not n57060 ; n57060_not
g76614 not n46611 ; n46611_not
g76615 not n54324 ; n54324_not
g76616 not n24444 ; n24444_not
g76617 not n25164 ; n25164_not
g76618 not n28611 ; n28611_not
g76619 not n24354 ; n24354_not
g76620 not n25722 ; n25722_not
g76621 not n48303 ; n48303_not
g76622 not n36702 ; n36702_not
g76623 not n24435 ; n24435_not
g76624 not n25173 ; n25173_not
g76625 not n24363 ; n24363_not
g76626 not n17460 ; n17460_not
g76627 not n33651 ; n33651_not
g76628 not n14238 ; n14238_not
g76629 not n44352 ; n44352_not
g76630 not n13653 ; n13653_not
g76631 not n21942 ; n21942_not
g76632 not n53253 ; n53253_not
g76633 not n41292 ; n41292_not
g76634 not n33903 ; n33903_not
g76635 not n33750 ; n33750_not
g76636 not n21195 ; n21195_not
g76637 not n21933 ; n21933_not
g76638 not n14247 ; n14247_not
g76639 not n33534 ; n33534_not
g76640 not n40851 ; n40851_not
g76641 not n13662 ; n13662_not
g76642 not n30096 ; n30096_not
g76643 not n21186 ; n21186_not
g76644 not n21924 ; n21924_not
g76645 not n33660 ; n33660_not
g76646 not n30708 ; n30708_not
g76647 not n32247 ; n32247_not
g76648 not n14256 ; n14256_not
g76649 not n16434 ; n16434_not
g76650 not n55233 ; n55233_not
g76651 not n21258 ; n21258_not
g76652 not n21249 ; n21249_not
g76653 not n33912 ; n33912_not
g76654 not n43470 ; n43470_not
g76655 not n13626 ; n13626_not
g76656 not n45135 ; n45135_not
g76657 not n40671 ; n40671_not
g76658 not n21285 ; n21285_not
g76659 not n43803 ; n43803_not
g76660 not n13635 ; n13635_not
g76661 not n53244 ; n53244_not
g76662 not n33543 ; n33543_not
g76663 not n53334 ; n53334_not
g76664 not n21960 ; n21960_not
g76665 not n14229 ; n14229_not
g76666 not n13644 ; n13644_not
g76667 not n53910 ; n53910_not
g76668 not n37314 ; n37314_not
g76669 not n21294 ; n21294_not
g76670 not n21951 ; n21951_not
g76671 not n13761 ; n13761_not
g76672 not n19611 ; n19611_not
g76673 not n33507 ; n33507_not
g76674 not n14292 ; n14292_not
g76675 not n37323 ; n37323_not
g76676 not n21339 ; n21339_not
g76677 not n13707 ; n13707_not
g76678 not n43506 ; n43506_not
g76679 not n21870 ; n21870_not
g76680 not n21348 ; n21348_not
g76681 not n13716 ; n13716_not
g76682 not n13752 ; n13752_not
g76683 not n21861 ; n21861_not
g76684 not n16443 ; n16443_not
g76685 not n30717 ; n30717_not
g76686 not n21852 ; n21852_not
g76687 not n19620 ; n19620_not
g76688 not n14319 ; n14319_not
g76689 not n53271 ; n53271_not
g76690 not n45162 ; n45162_not
g76691 not n21177 ; n21177_not
g76692 not n21915 ; n21915_not
g76693 not n13671 ; n13671_not
g76694 not n33525 ; n33525_not
g76695 not n32391 ; n32391_not
g76696 not n19602 ; n19602_not
g76697 not n21168 ; n21168_not
g76698 not n21906 ; n21906_not
g76699 not n48033 ; n48033_not
g76700 not n14265 ; n14265_not
g76701 not n13680 ; n13680_not
g76702 not n21159 ; n21159_not
g76703 not n16650 ; n16650_not
g76704 not n53901 ; n53901_not
g76705 not n33516 ; n33516_not
g76706 not n14274 ; n14274_not
g76707 not n37044 ; n37044_not
g76708 not n13770 ; n13770_not
g76709 not n40662 ; n40662_not
g76710 not n14283 ; n14283_not
g76711 not n14094 ; n14094_not
g76712 not n13509 ; n13509_not
g76713 not n43434 ; n43434_not
g76714 not n33615 ; n33615_not
g76715 not n50148 ; n50148_not
g76716 not n43821 ; n43821_not
g76717 not n13518 ; n13518_not
g76718 not n13527 ; n13527_not
g76719 not n53226 ; n53226_not
g76720 not n43443 ; n43443_not
g76721 not n13860 ; n13860_not
g76722 not n13536 ; n13536_not
g76723 not n13851 ; n13851_not
g76724 not n33606 ; n33606_not
g76725 not n13545 ; n13545_not
g76726 not n43452 ; n43452_not
g76727 not n19161 ; n19161_not
g76728 not n22086 ; n22086_not
g76729 not n14139 ; n14139_not
g76730 not n55800 ; n55800_not
g76731 not n22176 ; n22176_not
g76732 not n13464 ; n13464_not
g76733 not n19521 ; n19521_not
g76734 not n22167 ; n22167_not
g76735 not n14058 ; n14058_not
g76736 not n13473 ; n13473_not
g76737 not n55224 ; n55224_not
g76738 not n50076 ; n50076_not
g76739 not n14067 ; n14067_not
g76740 not n13482 ; n13482_not
g76741 not n19530 ; n19530_not
g76742 not n43425 ; n43425_not
g76743 not n30906 ; n30906_not
g76744 not n32229 ; n32229_not
g76745 not n22149 ; n22149_not
g76746 not n14076 ; n14076_not
g76747 not n13491 ; n13491_not
g76748 not n53316 ; n53316_not
g76749 not n14085 ; n14085_not
g76750 not n13590 ; n13590_not
g76751 not n30681 ; n30681_not
g76752 not n33930 ; n33930_not
g76753 not n14184 ; n14184_not
g76754 not n33561 ; n33561_not
g76755 not n43461 ; n43461_not
g76756 not n38115 ; n38115_not
g76757 not n32238 ; n32238_not
g76758 not n33642 ; n33642_not
g76759 not n33921 ; n33921_not
g76760 not n53325 ; n53325_not
g76761 not n14193 ; n14193_not
g76762 not n33552 ; n33552_not
g76763 not n13608 ; n13608_not
g76764 not n19143 ; n19143_not
g76765 not n13815 ; n13815_not
g76766 not n42930 ; n42930_not
g76767 not n30078 ; n30078_not
g76768 not n13617 ; n13617_not
g76769 not n13806 ; n13806_not
g76770 not n13554 ; n13554_not
g76771 not n22077 ; n22077_not
g76772 not n13842 ; n13842_not
g76773 not n42921 ; n42921_not
g76774 not n37305 ; n37305_not
g76775 not n14148 ; n14148_not
g76776 not n41283 ; n41283_not
g76777 not n13563 ; n13563_not
g76778 not n19152 ; n19152_not
g76779 not n38106 ; n38106_not
g76780 not n22059 ; n22059_not
g76781 not n14157 ; n14157_not
g76782 not n13572 ; n13572_not
g76783 not n50175 ; n50175_not
g76784 not n14166 ; n14166_not
g76785 not n13581 ; n13581_not
g76786 not n40680 ; n40680_not
g76787 not n33570 ; n33570_not
g76788 not n16425 ; n16425_not
g76789 not n14175 ; n14175_not
g76790 not n14526 ; n14526_not
g76791 not n33417 ; n33417_not
g76792 not n20934 ; n20934_not
g76793 not n21672 ; n21672_not
g76794 not n14544 ; n14544_not
g76795 not n40635 ; n40635_not
g76796 not n20925 ; n20925_not
g76797 not n21663 ; n21663_not
g76798 not n30168 ; n30168_not
g76799 not n20916 ; n20916_not
g76800 not n21654 ; n21654_not
g76801 not n16605 ; n16605_not
g76802 not n33408 ; n33408_not
g76803 not n21465 ; n21465_not
g76804 not n20907 ; n20907_not
g76805 not n21645 ; n21645_not
g76806 not n50283 ; n50283_not
g76807 not n13365 ; n13365_not
g76808 not n47412 ; n47412_not
g76809 not n21429 ; n21429_not
g76810 not n20970 ; n20970_not
g76811 not n21708 ; n21708_not
g76812 not n21438 ; n21438_not
g76813 not n50265 ; n50265_not
g76814 not n20961 ; n20961_not
g76815 not n33426 ; n33426_not
g76816 not n47403 ; n47403_not
g76817 not n53361 ; n53361_not
g76818 not n20952 ; n20952_not
g76819 not n21690 ; n21690_not
g76820 not n14049 ; n14049_not
g76821 not n30159 ; n30159_not
g76822 not n16614 ; n16614_not
g76823 not n14517 ; n14517_not
g76824 not n20943 ; n20943_not
g76825 not n21681 ; n21681_not
g76826 not n30177 ; n30177_not
g76827 not n43623 ; n43623_not
g76828 not n20871 ; n20871_not
g76829 not n21609 ; n21609_not
g76830 not n37350 ; n37350_not
g76831 not n14580 ; n14580_not
g76832 not n33741 ; n33741_not
g76833 not n20862 ; n20862_not
g76834 not n47421 ; n47421_not
g76835 not n43632 ; n43632_not
g76836 not n14562 ; n14562_not
g76837 not n33732 ; n33732_not
g76838 not n55710 ; n55710_not
g76839 not n20853 ; n20853_not
g76840 not n21591 ; n21591_not
g76841 not n43641 ; n43641_not
g76842 not n20844 ; n20844_not
g76843 not n21582 ; n21582_not
g76844 not n30186 ; n30186_not
g76845 not n43731 ; n43731_not
g76846 not n21636 ; n21636_not
g76847 not n43605 ; n43605_not
g76848 not n53370 ; n53370_not
g76849 not n37341 ; n37341_not
g76850 not n48024 ; n48024_not
g76851 not n21474 ; n21474_not
g76852 not n43614 ; n43614_not
g76853 not n21627 ; n21627_not
g76854 not n14571 ; n14571_not
g76855 not n50292 ; n50292_not
g76856 not n21483 ; n21483_not
g76857 not n20880 ; n20880_not
g76858 not n21618 ; n21618_not
g76859 not n32283 ; n32283_not
g76860 not n14364 ; n14364_not
g76861 not n21069 ; n21069_not
g76862 not n21807 ; n21807_not
g76863 not n53280 ; n53280_not
g76864 not n43515 ; n43515_not
g76865 not n16632 ; n16632_not
g76866 not n33840 ; n33840_not
g76867 not n33471 ; n33471_not
g76868 not n21384 ; n21384_not
g76869 not n50247 ; n50247_not
g76870 not n14382 ; n14382_not
g76871 not n43524 ; n43524_not
g76872 not n21393 ; n21393_not
g76873 not n37332 ; n37332_not
g76874 not n21780 ; n21780_not
g76875 not n33831 ; n33831_not
g76876 not n14391 ; n14391_not
g76877 not n21843 ; n21843_not
g76878 not n16641 ; n16641_not
g76879 not n19116 ; n19116_not
g76880 not n14328 ; n14328_not
g76881 not n13734 ; n13734_not
g76882 not n21096 ; n21096_not
g76883 not n21834 ; n21834_not
g76884 not n30726 ; n30726_not
g76885 not n21087 ; n21087_not
g76886 not n21825 ; n21825_not
g76887 not n32256 ; n32256_not
g76888 not n19107 ; n19107_not
g76889 not n21078 ; n21078_not
g76890 not n21816 ; n21816_not
g76891 not n33480 ; n33480_not
g76892 not n50238 ; n50238_not
g76893 not n21375 ; n21375_not
g76894 not n33705 ; n33705_not
g76895 not n21744 ; n21744_not
g76896 not n37701 ; n37701_not
g76897 not n16623 ; n16623_not
g76898 not n33813 ; n33813_not
g76899 not n33444 ; n33444_not
g76900 not n21735 ; n21735_not
g76901 not n14454 ; n14454_not
g76902 not n43551 ; n43551_not
g76903 not n21726 ; n21726_not
g76904 not n38133 ; n38133_not
g76905 not n33804 ; n33804_not
g76906 not n14472 ; n14472_not
g76907 not n21717 ; n21717_not
g76908 not n14481 ; n14481_not
g76909 not n33435 ; n33435_not
g76910 not n43560 ; n43560_not
g76911 not n43533 ; n43533_not
g76912 not n33462 ; n33462_not
g76913 not n21771 ; n21771_not
g76914 not n14409 ; n14409_not
g76915 not n21762 ; n21762_not
g76916 not n32265 ; n32265_not
g76917 not n33822 ; n33822_not
g76918 not n14427 ; n14427_not
g76919 not n21753 ; n21753_not
g76920 not n43542 ; n43542_not
g76921 not n14436 ; n14436_not
g76922 not n33453 ; n33453_not
g76923 not n32274 ; n32274_not
g76924 not n34128 ; n34128_not
g76925 not n13167 ; n13167_not
g76926 not n22581 ; n22581_not
g76927 not n41256 ; n41256_not
g76928 not n22572 ; n22572_not
g76929 not n34083 ; n34083_not
g76930 not n13158 ; n13158_not
g76931 not n19422 ; n19422_not
g76932 not n54009 ; n54009_not
g76933 not n22563 ; n22563_not
g76934 not n43902 ; n43902_not
g76935 not n30762 ; n30762_not
g76936 not n30564 ; n30564_not
g76937 not n22554 ; n22554_not
g76938 not n32328 ; n32328_not
g76939 not n22626 ; n22626_not
g76940 not n47016 ; n47016_not
g76941 not n22617 ; n22617_not
g76942 not n45126 ; n45126_not
g76943 not n19404 ; n19404_not
g76944 not n37233 ; n37233_not
g76945 not n22608 ; n22608_not
g76946 not n50058 ; n50058_not
g76947 not n47142 ; n47142_not
g76948 not n19233 ; n19233_not
g76949 not n19413 ; n19413_not
g76950 not n13176 ; n13176_not
g76951 not n22590 ; n22590_not
g76952 not n16380 ; n16380_not
g76953 not n37080 ; n37080_not
g76954 not n50067 ; n50067_not
g76955 not n19440 ; n19440_not
g76956 not n22491 ; n22491_not
g76957 not n38061 ; n38061_not
g76958 not n22482 ; n22482_not
g76959 not n37251 ; n37251_not
g76960 not n22473 ; n22473_not
g76961 not n22545 ; n22545_not
g76962 not n19431 ; n19431_not
g76963 not n37242 ; n37242_not
g76964 not n22536 ; n22536_not
g76965 not n22527 ; n22527_not
g76966 not n34092 ; n34092_not
g76967 not n42903 ; n42903_not
g76968 not n22518 ; n22518_not
g76969 not n22185 ; n22185_not
g76970 not n22509 ; n22509_not
g76971 not n41238 ; n41238_not
g76972 not n19350 ; n19350_not
g76973 not n37710 ; n37710_not
g76974 not n22770 ; n22770_not
g76975 not n13266 ; n13266_not
g76976 not n22761 ; n22761_not
g76977 not n40716 ; n40716_not
g76978 not n50049 ; n50049_not
g76979 not n13257 ; n13257_not
g76980 not n22752 ; n22752_not
g76981 not n22743 ; n22743_not
g76982 not n13248 ; n13248_not
g76983 not n22734 ; n22734_not
g76984 not n44901 ; n44901_not
g76985 not n47007 ; n47007_not
g76986 not n32193 ; n32193_not
g76987 not n19323 ; n19323_not
g76988 not n16344 ; n16344_not
g76989 not n22833 ; n22833_not
g76990 not n22824 ; n22824_not
g76991 not n13293 ; n13293_not
g76992 not n19332 ; n19332_not
g76993 not n22806 ; n22806_not
g76994 not n16353 ; n16353_not
g76995 not n19341 ; n19341_not
g76996 not n53172 ; n53172_not
g76997 not n54036 ; n54036_not
g76998 not n40725 ; n40725_not
g76999 not n38043 ; n38043_not
g77000 not n22095 ; n22095_not
g77001 not n34056 ; n34056_not
g77002 not n22671 ; n22671_not
g77003 not n19251 ; n19251_not
g77004 not n50931 ; n50931_not
g77005 not n22662 ; n22662_not
g77006 not n40707 ; n40707_not
g77007 not n45171 ; n45171_not
g77008 not n50490 ; n50490_not
g77009 not n22653 ; n22653_not
g77010 not n53190 ; n53190_not
g77011 not n54018 ; n54018_not
g77012 not n19242 ; n19242_not
g77013 not n22644 ; n22644_not
g77014 not n47160 ; n47160_not
g77015 not n22635 ; n22635_not
g77016 not n41247 ; n41247_not
g77017 not n34038 ; n34038_not
g77018 not n22725 ; n22725_not
g77019 not n37224 ; n37224_not
g77020 not n54027 ; n54027_not
g77021 not n22716 ; n22716_not
g77022 not n52461 ; n52461_not
g77023 not n47151 ; n47151_not
g77024 not n22707 ; n22707_not
g77025 not n53181 ; n53181_not
g77026 not n34047 ; n34047_not
g77027 not n44910 ; n44910_not
g77028 not n22680 ; n22680_not
g77029 not n21546 ; n21546_not
g77030 not n13392 ; n13392_not
g77031 not n48060 ; n48060_not
g77032 not n13383 ; n13383_not
g77033 not n13932 ; n13932_not
g77034 not n13374 ; n13374_not
g77035 not n43353 ; n43353_not
g77036 not n13941 ; n13941_not
g77037 not n30933 ; n30933_not
g77038 not n22275 ; n22275_not
g77039 not n13446 ; n13446_not
g77040 not n22347 ; n22347_not
g77041 not n53217 ; n53217_not
g77042 not n13437 ; n13437_not
g77043 not n21573 ; n21573_not
g77044 not n13428 ; n13428_not
g77045 not n50841 ; n50841_not
g77046 not n22338 ; n22338_not
g77047 not n43344 ; n43344_not
g77048 not n21564 ; n21564_not
g77049 not n13419 ; n13419_not
g77050 not n13914 ; n13914_not
g77051 not n55215 ; n55215_not
g77052 not n22329 ; n22329_not
g77053 not n42912 ; n42912_not
g77054 not n37071 ; n37071_not
g77055 not n21555 ; n21555_not
g77056 not n22239 ; n22239_not
g77057 not n19503 ; n19503_not
g77058 not n48051 ; n48051_not
g77059 not n43407 ; n43407_not
g77060 not n19512 ; n19512_not
g77061 not n13905 ; n13905_not
g77062 not n22194 ; n22194_not
g77063 not n13455 ; n13455_not
g77064 not n43416 ; n43416_not
g77065 not n22284 ; n22284_not
g77066 not n34065 ; n34065_not
g77067 not n13347 ; n13347_not
g77068 not n13950 ; n13950_not
g77069 not n50085 ; n50085_not
g77070 not n43362 ; n43362_not
g77071 not n22266 ; n22266_not
g77072 not n43371 ; n43371_not
g77073 not n22257 ; n22257_not
g77074 not n43380 ; n43380_not
g77075 not n30924 ; n30924_not
g77076 not n22437 ; n22437_not
g77077 not n43290 ; n43290_not
g77078 not n22428 ; n22428_not
g77079 not n13824 ; n13824_not
g77080 not n22419 ; n22419_not
g77081 not n53208 ; n53208_not
g77082 not n22464 ; n22464_not
g77083 not n38070 ; n38070_not
g77084 not n22455 ; n22455_not
g77085 not n34137 ; n34137_not
g77086 not n22446 ; n22446_not
g77087 not n32319 ; n32319_not
g77088 not n47205 ; n47205_not
g77089 not n22374 ; n22374_not
g77090 not n37260 ; n37260_not
g77091 not n43326 ; n43326_not
g77092 not n22365 ; n22365_not
g77093 not n30951 ; n30951_not
g77094 not n22356 ; n22356_not
g77095 not n43335 ; n43335_not
g77096 not n22392 ; n22392_not
g77097 not n19206 ; n19206_not
g77098 not n43308 ; n43308_not
g77099 not n22383 ; n22383_not
g77100 not n43317 ; n43317_not
g77101 not n32454 ; n32454_not
g77102 not n33147 ; n33147_not
g77103 not n30339 ; n30339_not
g77104 not n20664 ; n20664_not
g77105 not n50382 ; n50382_not
g77106 not n55134 ; n55134_not
g77107 not n33138 ; n33138_not
g77108 not n20655 ; n20655_not
g77109 not n32445 ; n32445_not
g77110 not n43047 ; n43047_not
g77111 not n33129 ; n33129_not
g77112 not n47133 ; n47133_not
g77113 not n37521 ; n37521_not
g77114 not n55404 ; n55404_not
g77115 not n20637 ; n20637_not
g77116 not n32436 ; n32436_not
g77117 not n15606 ; n15606_not
g77118 not n32463 ; n32463_not
g77119 not n33183 ; n33183_not
g77120 not n15624 ; n15624_not
g77121 not n50373 ; n50373_not
g77122 not n20709 ; n20709_not
g77123 not n33174 ; n33174_not
g77124 not n55413 ; n55413_not
g77125 not n53451 ; n53451_not
g77126 not n16407 ; n16407_not
g77127 not n41382 ; n41382_not
g77128 not n15642 ; n15642_not
g77129 not n33165 ; n33165_not
g77130 not n15651 ; n15651_not
g77131 not n33156 ; n33156_not
g77132 not n20682 ; n20682_not
g77133 not n20088 ; n20088_not
g77134 not n33066 ; n33066_not
g77135 not n30537 ; n30537_not
g77136 not n53622 ; n53622_not
g77137 not n30348 ; n30348_not
g77138 not n20574 ; n20574_not
g77139 not n43245 ; n43245_not
g77140 not n33057 ; n33057_not
g77141 not n33039 ; n33039_not
g77142 not n20565 ; n20565_not
g77143 not n30285 ; n30285_not
g77144 not n20097 ; n20097_not
g77145 not n15804 ; n15804_not
g77146 not n33048 ; n33048_not
g77147 not n32418 ; n32418_not
g77148 not n30357 ; n30357_not
g77149 not n53613 ; n53613_not
g77150 not n20547 ; n20547_not
g77151 not n16335 ; n16335_not
g77152 not n30294 ; n30294_not
g77153 not n43227 ; n43227_not
g77154 not n30546 ; n30546_not
g77155 not n15714 ; n15714_not
g77156 not n32670 ; n32670_not
g77157 not n53631 ; n53631_not
g77158 not n20619 ; n20619_not
g77159 not n15732 ; n15732_not
g77160 not n50391 ; n50391_not
g77161 not n55143 ; n55143_not
g77162 not n15741 ; n15741_not
g77163 not n43056 ; n43056_not
g77164 not n33093 ; n33093_not
g77165 not n20079 ; n20079_not
g77166 not n33084 ; n33084_not
g77167 not n32427 ; n32427_not
g77168 not n33075 ; n33075_not
g77169 not n16362 ; n16362_not
g77170 not n20592 ; n20592_not
g77171 not n43236 ; n43236_not
g77172 not n53433 ; n53433_not
g77173 not n30591 ; n30591_not
g77174 not n41355 ; n41355_not
g77175 not n32490 ; n32490_not
g77176 not n30582 ; n30582_not
g77177 not n43029 ; n43029_not
g77178 not n20835 ; n20835_not
g77179 not n32922 ; n32922_not
g77180 not n41391 ; n41391_not
g77181 not n33246 ; n33246_not
g77182 not n20826 ; n20826_not
g77183 not n30528 ; n30528_not
g77184 not n15048 ; n15048_not
g77185 not n30573 ; n30573_not
g77186 not n32508 ; n32508_not
g77187 not n50364 ; n50364_not
g77188 not n41337 ; n41337_not
g77189 not n15093 ; n15093_not
g77190 not n32634 ; n32634_not
g77191 not n16470 ; n16470_not
g77192 not n15084 ; n15084_not
g77193 not n33282 ; n33282_not
g77194 not n15075 ; n15075_not
g77195 not n20718 ; n20718_not
g77196 not n33264 ; n33264_not
g77197 not n43182 ; n43182_not
g77198 not n47034 ; n47034_not
g77199 not n43038 ; n43038_not
g77200 not n33219 ; n33219_not
g77201 not n20763 ; n20763_not
g77202 not n19305 ; n19305_not
g77203 not n32472 ; n32472_not
g77204 not n53640 ; n53640_not
g77205 not n20754 ; n20754_not
g77206 not n55431 ; n55431_not
g77207 not n32652 ; n32652_not
g77208 not n20745 ; n20745_not
g77209 not n55125 ; n55125_not
g77210 not n33192 ; n33192_not
g77211 not n55422 ; n55422_not
g77212 not n20727 ; n20727_not
g77213 not n20817 ; n20817_not
g77214 not n33237 ; n33237_not
g77215 not n15039 ; n15039_not
g77216 not n20808 ; n20808_not
g77217 not n16452 ; n16452_not
g77218 not n55440 ; n55440_not
g77219 not n33228 ; n33228_not
g77220 not n32481 ; n32481_not
g77221 not n43191 ; n43191_not
g77222 not n41373 ; n41373_not
g77223 not n19314 ; n19314_not
g77224 not n32517 ; n32517_not
g77225 not n47070 ; n47070_not
g77226 not n32823 ; n32823_not
g77227 not n16083 ; n16083_not
g77228 not n30474 ; n30474_not
g77229 not n43164 ; n43164_not
g77230 not n20187 ; n20187_not
g77231 not n50463 ; n50463_not
g77232 not n16092 ; n16092_not
g77233 not n32814 ; n32814_not
g77234 not n32643 ; n32643_not
g77235 not n55314 ; n55314_not
g77236 not n32805 ; n32805_not
g77237 not n47061 ; n47061_not
g77238 not n30465 ; n30465_not
g77239 not n20295 ; n20295_not
g77240 not n16227 ; n16227_not
g77241 not n53541 ; n53541_not
g77242 not n32850 ; n32850_not
g77243 not n40860 ; n40860_not
g77244 not n16047 ; n16047_not
g77245 not n20178 ; n20178_not
g77246 not n20358 ; n20358_not
g77247 not n32535 ; n32535_not
g77248 not n50436 ; n50436_not
g77249 not n41427 ; n41427_not
g77250 not n16056 ; n16056_not
g77251 not n32841 ; n32841_not
g77252 not n20349 ; n20349_not
g77253 not n32625 ; n32625_not
g77254 not n16065 ; n16065_not
g77255 not n32526 ; n32526_not
g77256 not n32724 ; n32724_not
g77257 not n32832 ; n32832_not
g77258 not n53523 ; n53523_not
g77259 not n16074 ; n16074_not
g77260 not n16236 ; n16236_not
g77261 not n43092 ; n43092_not
g77262 not n55305 ; n55305_not
g77263 not n16164 ; n16164_not
g77264 not n50454 ; n50454_not
g77265 not n16218 ; n16218_not
g77266 not n16173 ; n16173_not
g77267 not n50256 ; n50256_not
g77268 not n32760 ; n32760_not
g77269 not n43119 ; n43119_not
g77270 not n16182 ; n16182_not
g77271 not n32751 ; n32751_not
g77272 not n47052 ; n47052_not
g77273 not n16191 ; n16191_not
g77274 not n16209 ; n16209_not
g77275 not n45117 ; n45117_not
g77276 not n15660 ; n15660_not
g77277 not n32742 ; n32742_not
g77278 not n30483 ; n30483_not
g77279 not n20286 ; n20286_not
g77280 not n15705 ; n15705_not
g77281 not n16119 ; n16119_not
g77282 not n20277 ; n20277_not
g77283 not n16128 ; n16128_not
g77284 not n32733 ; n32733_not
g77285 not n43146 ; n43146_not
g77286 not n20196 ; n20196_not
g77287 not n41418 ; n41418_not
g77288 not n16137 ; n16137_not
g77289 not n50445 ; n50445_not
g77290 not n20268 ; n20268_not
g77291 not n30492 ; n30492_not
g77292 not n43137 ; n43137_not
g77293 not n20259 ; n20259_not
g77294 not n16146 ; n16146_not
g77295 not n16155 ; n16155_not
g77296 not n16290 ; n16290_not
g77297 not n15822 ; n15822_not
g77298 not n15903 ; n15903_not
g77299 not n20484 ; n20484_not
g77300 not n50409 ; n50409_not
g77301 not n47106 ; n47106_not
g77302 not n43272 ; n43272_not
g77303 not n53460 ; n53460_not
g77304 not n37602 ; n37602_not
g77305 not n43074 ; n43074_not
g77306 not n20475 ; n20475_not
g77307 not n15912 ; n15912_not
g77308 not n37611 ; n37611_not
g77309 not n43281 ; n43281_not
g77310 not n20466 ; n20466_not
g77311 not n15921 ; n15921_not
g77312 not n16272 ; n16272_not
g77313 not n32409 ; n32409_not
g77314 not n32931 ; n32931_not
g77315 not n20457 ; n20457_not
g77316 not n32715 ; n32715_not
g77317 not n15831 ; n15831_not
g77318 not n50472 ; n50472_not
g77319 not n20529 ; n20529_not
g77320 not n15840 ; n15840_not
g77321 not n16317 ; n16317_not
g77322 not n47043 ; n47043_not
g77323 not n20493 ; n20493_not
g77324 not n53604 ; n53604_not
g77325 not n50427 ; n50427_not
g77326 not n16254 ; n16254_not
g77327 not n55332 ; n55332_not
g77328 not n32571 ; n32571_not
g77329 not n53514 ; n53514_not
g77330 not n20169 ; n20169_not
g77331 not n55323 ; n55323_not
g77332 not n32562 ; n32562_not
g77333 not n43209 ; n43209_not
g77334 not n20394 ; n20394_not
g77335 not n16245 ; n16245_not
g77336 not n20385 ; n20385_not
g77337 not n32553 ; n32553_not
g77338 not n16029 ; n16029_not
g77339 not n32544 ; n32544_not
g77340 not n20376 ; n20376_not
g77341 not n53505 ; n53505_not
g77342 not n15750 ; n15750_not
g77343 not n16038 ; n16038_not
g77344 not n30258 ; n30258_not
g77345 not n20367 ; n20367_not
g77346 not n15930 ; n15930_not
g77347 not n20448 ; n20448_not
g77348 not n20439 ; n20439_not
g77349 not n50418 ; n50418_not
g77350 not n43254 ; n43254_not
g77351 not n55350 ; n55350_not
g77352 not n55170 ; n55170_not
g77353 not n32904 ; n32904_not
g77354 not n19800 ; n19800_not
g77355 not n55341 ; n55341_not
g77356 not n37620 ; n37620_not
g77357 not n30249 ; n30249_not
g77358 not n33273 ; n33273_not
g77359 not n55602 ; n55602_not
g77360 not n19710 ; n19710_not
g77361 not n16560 ; n16560_not
g77362 not n30618 ; n30618_not
g77363 not n33390 ; n33390_not
g77364 not n19701 ; n19701_not
g77365 not n53811 ; n53811_not
g77366 not n21357 ; n21357_not
g77367 not n45144 ; n45144_not
g77368 not n30735 ; n30735_not
g77369 not n55611 ; n55611_not
g77370 not n53802 ; n53802_not
g77371 not n30609 ; n30609_not
g77372 not n50481 ; n50481_not
g77373 not n55044 ; n55044_not
g77374 not n14355 ; n14355_not
g77375 not n41346 ; n41346_not
g77376 not n55053 ; n55053_not
g77377 not n30654 ; n30654_not
g77378 not n30627 ; n30627_not
g77379 not n53406 ; n53406_not
g77380 not n55260 ; n55260_not
g77381 not n16551 ; n16551_not
g77382 not n30636 ; n30636_not
g77383 not n48006 ; n48006_not
g77384 not n30645 ; n30645_not
g77385 not n30195 ; n30195_not
g77386 not n45009 ; n45009_not
g77387 not n21519 ; n21519_not
g77388 not n21492 ; n21492_not
g77389 not n55251 ; n55251_not
g77390 not n53343 ; n53343_not
g77391 not n41229 ; n41229_not
g77392 not n43650 ; n43650_not
g77393 not n55701 ; n55701_not
g77394 not n19071 ; n19071_not
g77395 not n30753 ; n30753_not
g77396 not n38142 ; n38142_not
g77397 not n19062 ; n19062_not
g77398 not n21528 ; n21528_not
g77399 not n33714 ; n33714_not
g77400 not n14535 ; n14535_not
g77401 not n50328 ; n50328_not
g77402 not n47430 ; n47430_not
g77403 not n41328 ; n41328_not
g77404 not n53820 ; n53820_not
g77405 not n33624 ; n33624_not
g77406 not n14445 ; n14445_not
g77407 not n55620 ; n55620_not
g77408 not n47025 ; n47025_not
g77409 not n19053 ; n19053_not
g77410 not n43065 ; n43065_not
g77411 not n14490 ; n14490_not
g77412 not n55008 ; n55008_not
g77413 not n21447 ; n21447_not
g77414 not n32580 ; n32580_not
g77415 not n15183 ; n15183_not
g77416 not n55512 ; n55512_not
g77417 not n15174 ; n15174_not
g77418 not n37431 ; n37431_not
g77419 not n53712 ; n53712_not
g77420 not n55080 ; n55080_not
g77421 not n16515 ; n16515_not
g77422 not n15165 ; n15165_not
g77423 not n43155 ; n43155_not
g77424 not n33372 ; n33372_not
g77425 not n33363 ; n33363_not
g77426 not n53730 ; n53730_not
g77427 not n15192 ; n15192_not
g77428 not n55521 ; n55521_not
g77429 not n37422 ; n37422_not
g77430 not n53721 ; n53721_not
g77431 not n20628 ; n20628_not
g77432 not n53415 ; n53415_not
g77433 not n33327 ; n33327_not
g77434 not n33309 ; n33309_not
g77435 not n55503 ; n55503_not
g77436 not n53703 ; n53703_not
g77437 not n42444 ; n42444_not
g77438 not n33354 ; n33354_not
g77439 not n15138 ; n15138_not
g77440 not n33345 ; n33345_not
g77441 not n15129 ; n15129_not
g77442 not n20673 ; n20673_not
g77443 not n30690 ; n30690_not
g77444 not n53424 ; n53424_not
g77445 not n15057 ; n15057_not
g77446 not n32607 ; n32607_not
g77447 not n37404 ; n37404_not
g77448 not n38124 ; n38124_not
g77449 not n45054 ; n45054_not
g77450 not n30663 ; n30663_not
g77451 not n30672 ; n30672_not
g77452 not n41265 ; n41265_not
g77453 not n30267 ; n30267_not
g77454 not n20538 ; n20538_not
g77455 not n50346 ; n50346_not
g77456 not n33318 ; n33318_not
g77457 not n15147 ; n15147_not
g77458 not n50355 ; n50355_not
g77459 not n37413 ; n37413_not
g77460 not n55530 ; n55530_not
g77461 not n47250 ; n47250_not
g77462 not n20583 ; n20583_not
g77463 not n51093 ; n51093_not
g77464 not n29520 ; n29520_not
g77465 not n22914 ; n22914_not
g77466 not n17226 ; n17226_not
g77467 not n23814 ; n23814_not
g77468 not n12654 ; n12654_not
g77469 not n42750 ; n42750_not
g77470 not n23391 ; n23391_not
g77471 not n54243 ; n54243_not
g77472 not n12942 ; n12942_not
g77473 not n34506 ; n34506_not
g77474 not n23409 ; n23409_not
g77475 not n12195 ; n12195_not
g77476 not n17172 ; n17172_not
g77477 not n45234 ; n45234_not
g77478 not n12933 ; n12933_not
g77479 not n23751 ; n23751_not
g77480 not n17154 ; n17154_not
g77481 not n31248 ; n31248_not
g77482 not n11745 ; n11745_not
g77483 not n34704 ; n34704_not
g77484 not n23373 ; n23373_not
g77485 not n42804 ; n42804_not
g77486 not n22932 ; n22932_not
g77487 not n12951 ; n12951_not
g77488 not n34155 ; n34155_not
g77489 not n12267 ; n12267_not
g77490 not n12519 ; n12519_not
g77491 not n23364 ; n23364_not
g77492 not n29250 ; n29250_not
g77493 not n12726 ; n12726_not
g77494 not n34164 ; n34164_not
g77495 not n12276 ; n12276_not
g77496 not n34344 ; n34344_not
g77497 not n34650 ; n34650_not
g77498 not n29223 ; n29223_not
g77499 not n23382 ; n23382_not
g77500 not n42723 ; n42723_not
g77501 not n29052 ; n29052_not
g77502 not n22923 ; n22923_not
g77503 not n29502 ; n29502_not
g77504 not n11736 ; n11736_not
g77505 not n11763 ; n11763_not
g77506 not n34713 ; n34713_not
g77507 not n29205 ; n29205_not
g77508 not n23445 ; n23445_not
g77509 not n12186 ; n12186_not
g77510 not n23436 ; n23436_not
g77511 not n12663 ; n12663_not
g77512 not n23463 ; n23463_not
g77513 not n11772 ; n11772_not
g77514 not n12744 ; n12744_not
g77515 not n17217 ; n17217_not
g77516 not n54153 ; n54153_not
g77517 not n12672 ; n12672_not
g77518 not n12915 ; n12915_not
g77519 not n23454 ; n23454_not
g77520 not n51084 ; n51084_not
g77521 not n29070 ; n29070_not
g77522 not n34515 ; n34515_not
g77523 not n31194 ; n31194_not
g77524 not n23418 ; n23418_not
g77525 not n37161 ; n37161_not
g77526 not n32382 ; n32382_not
g77527 not n29511 ; n29511_not
g77528 not n29106 ; n29106_not
g77529 not n19017 ; n19017_not
g77530 not n12285 ; n12285_not
g77531 not n29061 ; n29061_not
g77532 not n12294 ; n12294_not
g77533 not n31068 ; n31068_not
g77534 not n11754 ; n11754_not
g77535 not n12924 ; n12924_not
g77536 not n23427 ; n23427_not
g77537 not n55062 ; n55062_not
g77538 not n12492 ; n12492_not
g77539 not n53091 ; n53091_not
g77540 not n29214 ; n29214_not
g77541 not n34461 ; n34461_not
g77542 not n34227 ; n34227_not
g77543 not n12546 ; n12546_not
g77544 not n29034 ; n29034_not
g77545 not n23832 ; n23832_not
g77546 not n23292 ; n23292_not
g77547 not n40761 ; n40761_not
g77548 not n47115 ; n47115_not
g77549 not n56025 ; n56025_not
g77550 not n34470 ; n34470_not
g77551 not n34218 ; n34218_not
g77552 not n12627 ; n12627_not
g77553 not n34731 ; n34731_not
g77554 not n12708 ; n12708_not
g77555 not n12618 ; n12618_not
g77556 not n54333 ; n54333_not
g77557 not n53109 ; n53109_not
g77558 not n42822 ; n42822_not
g77559 not n23265 ; n23265_not
g77560 not n23652 ; n23652_not
g77561 not n53118 ; n53118_not
g77562 not n34335 ; n34335_not
g77563 not n29241 ; n29241_not
g77564 not n11691 ; n11691_not
g77565 not n12258 ; n12258_not
g77566 not n23256 ; n23256_not
g77567 not n23283 ; n23283_not
g77568 not n12609 ; n12609_not
g77569 not n31086 ; n31086_not
g77570 not n34236 ; n34236_not
g77571 not n23274 ; n23274_not
g77572 not n53046 ; n53046_not
g77573 not n32373 ; n32373_not
g77574 not n34245 ; n34245_not
g77575 not n34173 ; n34173_not
g77576 not n31239 ; n31239_not
g77577 not n23346 ; n23346_not
g77578 not n29043 ; n29043_not
g77579 not n34182 ; n34182_not
g77580 not n32337 ; n32337_not
g77581 not n31077 ; n31077_not
g77582 not n43812 ; n43812_not
g77583 not n17163 ; n17163_not
g77584 not n23355 ; n23355_not
g77585 not n37143 ; n37143_not
g77586 not n52506 ; n52506_not
g77587 not n29232 ; n29232_not
g77588 not n19125 ; n19125_not
g77589 not n12960 ; n12960_not
g77590 not n34740 ; n34740_not
g77591 not n11727 ; n11727_not
g77592 not n42813 ; n42813_not
g77593 not n34191 ; n34191_not
g77594 not n11718 ; n11718_not
g77595 not n52641 ; n52641_not
g77596 not n12249 ; n12249_not
g77597 not n23319 ; n23319_not
g77598 not n17244 ; n17244_not
g77599 not n55152 ; n55152_not
g77600 not n34209 ; n34209_not
g77601 not n11709 ; n11709_not
g77602 not n23337 ; n23337_not
g77603 not n40770 ; n40770_not
g77604 not n23823 ; n23823_not
g77605 not n17235 ; n17235_not
g77606 not n12528 ; n12528_not
g77607 not n34290 ; n34290_not
g77608 not n40644 ; n40644_not
g77609 not n23328 ; n23328_not
g77610 not n48042 ; n48042_not
g77611 not n12717 ; n12717_not
g77612 not n16542 ; n16542_not
g77613 not n12834 ; n12834_not
g77614 not n12384 ; n12384_not
g77615 not n38502 ; n38502_not
g77616 not n34380 ; n34380_not
g77617 not n55107 ; n55107_not
g77618 not n23616 ; n23616_not
g77619 not n12456 ; n12456_not
g77620 not n12825 ; n12825_not
g77621 not n34623 ; n34623_not
g77622 not n48123 ; n48123_not
g77623 not n31284 ; n31284_not
g77624 not n23607 ; n23607_not
g77625 not n11853 ; n11853_not
g77626 not n51048 ; n51048_not
g77627 not n11835 ; n11835_not
g77628 not n23571 ; n23571_not
g77629 not n23733 ; n23733_not
g77630 not n12852 ; n12852_not
g77631 not n37125 ; n37125_not
g77632 not n32364 ; n32364_not
g77633 not n11844 ; n11844_not
g77634 not n12843 ; n12843_not
g77635 not n52911 ; n52911_not
g77636 not n12375 ; n12375_not
g77637 not n34263 ; n34263_not
g77638 not n23742 ; n23742_not
g77639 not n23580 ; n23580_not
g77640 not n53064 ; n53064_not
g77641 not n29313 ; n29313_not
g77642 not n40806 ; n40806_not
g77643 not n12438 ; n12438_not
g77644 not n34254 ; n34254_not
g77645 not n51057 ; n51057_not
g77646 not n23643 ; n23643_not
g77647 not n37170 ; n37170_not
g77648 not n34605 ; n34605_not
g77649 not n17046 ; n17046_not
g77650 not n34614 ; n34614_not
g77651 not n12447 ; n12447_not
g77652 not n29304 ; n29304_not
g77653 not n31266 ; n31266_not
g77654 not n23661 ; n23661_not
g77655 not n19044 ; n19044_not
g77656 not n48114 ; n48114_not
g77657 not n40734 ; n40734_not
g77658 not n52920 ; n52920_not
g77659 not n11871 ; n11871_not
g77660 not n53055 ; n53055_not
g77661 not n40815 ; n40815_not
g77662 not n32355 ; n32355_not
g77663 not n11862 ; n11862_not
g77664 not n50508 ; n50508_not
g77665 not n42741 ; n42741_not
g77666 not n12393 ; n12393_not
g77667 not n12816 ; n12816_not
g77668 not n12429 ; n12429_not
g77669 not n18900 ; n18900_not
g77670 not n19035 ; n19035_not
g77671 not n23634 ; n23634_not
g77672 not n29322 ; n29322_not
g77673 not n11880 ; n11880_not
g77674 not n17181 ; n17181_not
g77675 not n31275 ; n31275_not
g77676 not n12807 ; n12807_not
g77677 not n31176 ; n31176_not
g77678 not n12780 ; n12780_not
g77679 not n12087 ; n12087_not
g77680 not n29421 ; n29421_not
g77681 not n34641 ; n34641_not
g77682 not n12483 ; n12483_not
g77683 not n29430 ; n29430_not
g77684 not n53073 ; n53073_not
g77685 not n12753 ; n12753_not
g77686 not n23724 ; n23724_not
g77687 not n12096 ; n12096_not
g77688 not n23490 ; n23490_not
g77689 not n12474 ; n12474_not
g77690 not n23517 ; n23517_not
g77691 not n29412 ; n29412_not
g77692 not n31059 ; n31059_not
g77693 not n12339 ; n12339_not
g77694 not n41940 ; n41940_not
g77695 not n18423 ; n18423_not
g77696 not n23508 ; n23508_not
g77697 not n34353 ; n34353_not
g77698 not n12177 ; n12177_not
g77699 not n12906 ; n12906_not
g77700 not n11637 ; n11637_not
g77701 not n23472 ; n23472_not
g77702 not n34281 ; n34281_not
g77703 not n53082 ; n53082_not
g77704 not n11790 ; n11790_not
g77705 not n17208 ; n17208_not
g77706 not n37116 ; n37116_not
g77707 not n11781 ; n11781_not
g77708 not n23481 ; n23481_not
g77709 not n29115 ; n29115_not
g77710 not n34632 ; n34632_not
g77711 not n23706 ; n23706_not
g77712 not n31293 ; n31293_not
g77713 not n23544 ; n23544_not
g77714 not n12357 ; n12357_not
g77715 not n12078 ; n12078_not
g77716 not n34272 ; n34272_not
g77717 not n23562 ; n23562_not
g77718 not n12771 ; n12771_not
g77719 not n34362 ; n34362_not
g77720 not n12366 ; n12366_not
g77721 not n23553 ; n23553_not
g77722 not n12465 ; n12465_not
g77723 not n12861 ; n12861_not
g77724 not n11826 ; n11826_not
g77725 not n29403 ; n29403_not
g77726 not n34722 ; n34722_not
g77727 not n52902 ; n52902_not
g77728 not n11808 ; n11808_not
g77729 not n23526 ; n23526_not
g77730 not n19080 ; n19080_not
g77731 not n40752 ; n40752_not
g77732 not n48105 ; n48105_not
g77733 not n11817 ; n11817_not
g77734 not n42732 ; n42732_not
g77735 not n23535 ; n23535_not
g77736 not n19026 ; n19026_not
g77737 not n18333 ; n18333_not
g77738 not n22842 ; n22842_not
g77739 not n12870 ; n12870_not
g77740 not n12348 ; n12348_not
g77741 not n53136 ; n53136_not
g77742 not n29700 ; n29700_not
g77743 not n29133 ; n29133_not
g77744 not n17091 ; n17091_not
g77745 not n54063 ; n54063_not
g77746 not n51039 ; n51039_not
g77747 not n34371 ; n34371_not
g77748 not n17280 ; n17280_not
g77749 not n42705 ; n42705_not
g77750 not n53145 ; n53145_not
g77751 not n29142 ; n29142_not
g77752 not n23841 ; n23841_not
g77753 not n24453 ; n24453_not
g77754 not n38016 ; n38016_not
g77755 not n12591 ; n12591_not
g77756 not n29610 ; n29610_not
g77757 not n23058 ; n23058_not
g77758 not n11682 ; n11682_not
g77759 not n11673 ; n11673_not
g77760 not n17271 ; n17271_not
g77761 not n23085 ; n23085_not
g77762 not n11655 ; n11655_not
g77763 not n11664 ; n11664_not
g77764 not n34812 ; n34812_not
g77765 not n29160 ; n29160_not
g77766 not n34326 ; n34326_not
g77767 not n23076 ; n23076_not
g77768 not n34425 ; n34425_not
g77769 not n13275 ; n13275_not
g77770 not n19260 ; n19260_not
g77771 not n41805 ; n41805_not
g77772 not n23049 ; n23049_not
g77773 not n37206 ; n37206_not
g77774 not n42534 ; n42534_not
g77775 not n12681 ; n12681_not
g77776 not n31347 ; n31347_not
g77777 not n31356 ; n31356_not
g77778 not n38034 ; n38034_not
g77779 not n53154 ; n53154_not
g77780 not n22851 ; n22851_not
g77781 not n53163 ; n53163_not
g77782 not n29124 ; n29124_not
g77783 not n53028 ; n53028_not
g77784 not n45180 ; n45180_not
g77785 not n54045 ; n54045_not
g77786 not n41436 ; n41436_not
g77787 not n50517 ; n50517_not
g77788 not n40842 ; n40842_not
g77789 not n22941 ; n22941_not
g77790 not n53037 ; n53037_not
g77791 not n37215 ; n37215_not
g77792 not n48141 ; n48141_not
g77793 not n40824 ; n40824_not
g77794 not n34416 ; n34416_not
g77795 not n13338 ; n13338_not
g77796 not n34308 ; n34308_not
g77797 not n29601 ; n29601_not
g77798 not n52830 ; n52830_not
g77799 not n12636 ; n12636_not
g77800 not n38025 ; n38025_not
g77801 not n34317 ; n34317_not
g77802 not n54054 ; n54054_not
g77803 not n52551 ; n52551_not
g77804 not n53019 ; n53019_not
g77805 not n37152 ; n37152_not
g77806 not n29025 ; n29025_not
g77807 not n41850 ; n41850_not
g77808 not n42831 ; n42831_not
g77809 not n17136 ; n17136_not
g77810 not n12564 ; n12564_not
g77811 not n23184 ; n23184_not
g77812 not n12168 ; n12168_not
g77813 not n29151 ; n29151_not
g77814 not n13086 ; n13086_not
g77815 not n40626 ; n40626_not
g77816 not n31095 ; n31095_not
g77817 not n32292 ; n32292_not
g77818 not n13095 ; n13095_not
g77819 not n23193 ; n23193_not
g77820 not n31338 ; n31338_not
g77821 not n23157 ; n23157_not
g77822 not n40617 ; n40617_not
g77823 not n18801 ; n18801_not
g77824 not n23175 ; n23175_not
g77825 not n17262 ; n17262_not
g77826 not n23166 ; n23166_not
g77827 not n34434 ; n34434_not
g77828 not n19170 ; n19170_not
g77829 not n13059 ; n13059_not
g77830 not n23238 ; n23238_not
g77831 not n18810 ; n18810_not
g77832 not n23247 ; n23247_not
g77833 not n17253 ; n17253_not
g77834 not n31329 ; n31329_not
g77835 not n42714 ; n42714_not
g77836 not n12582 ; n12582_not
g77837 not n13077 ; n13077_not
g77838 not n19008 ; n19008_not
g77839 not n12573 ; n12573_not
g77840 not n53127 ; n53127_not
g77841 not n34443 ; n34443_not
g77842 not n23229 ; n23229_not
g77843 not n54108 ; n54108_not
g77844 not n13068 ; n13068_not
g77845 not n48132 ; n48132_not
g77846 not n13185 ; n13185_not
g77847 not n30942 ; n30942_not
g77848 not n47340 ; n47340_not
g77849 not n19215 ; n19215_not
g77850 not n51066 ; n51066_not
g77851 not n56070 ; n56070_not
g77852 not n16308 ; n16308_not
g77853 not n23067 ; n23067_not
g77854 not n40608 ; n40608_not
g77855 not n11646 ; n11646_not
g77856 not n42840 ; n42840_not
g77857 not n37134 ; n37134_not
g77858 not n23148 ; n23148_not
g77859 not n23139 ; n23139_not
g77860 not n33391 ; n33391_not
g77861 not n35803 ; n35803_not
g77862 not n32266 ; n32266_not
g77863 not n46432 ; n46432_not
g77864 not n36037 ; n36037_not
g77865 not n28720 ; n28720_not
g77866 not n34705 ; n34705_not
g77867 not n39250 ; n39250_not
g77868 not n30493 ; n30493_not
g77869 not n34642 ; n34642_not
g77870 not n36505 ; n36505_not
g77871 not n50482 ; n50482_not
g77872 not n32248 ; n32248_not
g77873 not n34516 ; n34516_not
g77874 not n26830 ; n26830_not
g77875 not n51850 ; n51850_not
g77876 not n36082 ; n36082_not
g77877 not n39115 ; n39115_not
g77878 not n28702 ; n28702_not
g77879 not n29107 ; n29107_not
g77880 not n49105 ; n49105_not
g77881 not n35722 ; n35722_not
g77882 not n46540 ; n46540_not
g77883 not n38305 ; n38305_not
g77884 not n36514 ; n36514_not
g77885 not n50680 ; n50680_not
g77886 not n29116 ; n29116_not
g77887 not n29125 ; n29125_not
g77888 not n47530 ; n47530_not
g77889 not n30259 ; n30259_not
g77890 not n39214 ; n39214_not
g77891 not n47440 ; n47440_not
g77892 not n30664 ; n30664_not
g77893 not n49141 ; n49141_not
g77894 not n51139 ; n51139_not
g77895 not n31753 ; n31753_not
g77896 not n48250 ; n48250_not
g77897 not n48700 ; n48700_not
g77898 not n35038 ; n35038_not
g77899 not n39223 ; n39223_not
g77900 not n48601 ; n48601_not
g77901 not n34633 ; n34633_not
g77902 not n31906 ; n31906_not
g77903 not n30277 ; n30277_not
g77904 not n31249 ; n31249_not
g77905 not n34651 ; n34651_not
g77906 not n29161 ; n29161_not
g77907 not n26920 ; n26920_not
g77908 not n32086 ; n32086_not
g77909 not n36064 ; n36064_not
g77910 not n29071 ; n29071_not
g77911 not n32239 ; n32239_not
g77912 not n37009 ; n37009_not
g77913 not n33328 ; n33328_not
g77914 not n35911 ; n35911_not
g77915 not n35713 ; n35713_not
g77916 not n30682 ; n30682_not
g77917 not n27415 ; n27415_not
g77918 not n46522 ; n46522_not
g77919 not n37135 ; n37135_not
g77920 not n32257 ; n32257_not
g77921 not n47512 ; n47512_not
g77922 not n48223 ; n48223_not
g77923 not n50338 ; n50338_not
g77924 not n30466 ; n30466_not
g77925 not n30655 ; n30655_not
g77926 not n38161 ; n38161_not
g77927 not n31069 ; n31069_not
g77928 not n51931 ; n51931_not
g77929 not n34723 ; n34723_not
g77930 not n29152 ; n29152_not
g77931 not n35056 ; n35056_not
g77932 not n32275 ; n32275_not
g77933 not n51913 ; n51913_not
g77934 not n46423 ; n46423_not
g77935 not n32545 ; n32545_not
g77936 not n30691 ; n30691_not
g77937 not n51922 ; n51922_not
g77938 not n29170 ; n29170_not
g77939 not n33319 ; n33319_not
g77940 not n35731 ; n35731_not
g77941 not n49132 ; n49132_not
g77942 not n50932 ; n50932_not
g77943 not n50671 ; n50671_not
g77944 not n35812 ; n35812_not
g77945 not n39133 ; n39133_not
g77946 not n48232 ; n48232_not
g77947 not n30646 ; n30646_not
g77948 not n35047 ; n35047_not
g77949 not n49114 ; n49114_not
g77950 not n35821 ; n35821_not
g77951 not n48241 ; n48241_not
g77952 not n31258 ; n31258_not
g77953 not n34624 ; n34624_not
g77954 not n38314 ; n38314_not
g77955 not n26902 ; n26902_not
g77956 not n39232 ; n39232_not
g77957 not n39241 ; n39241_not
g77958 not n46513 ; n46513_not
g77959 not n33373 ; n33373_not
g77960 not n27433 ; n27433_not
g77961 not n28711 ; n28711_not
g77962 not n31744 ; n31744_not
g77963 not n49123 ; n49123_not
g77964 not n35902 ; n35902_not
g77965 not n47503 ; n47503_not
g77966 not n35830 ; n35830_not
g77967 not n38116 ; n38116_not
g77968 not n32554 ; n32554_not
g77969 not n39124 ; n39124_not
g77970 not n49204 ; n49204_not
g77971 not n32284 ; n32284_not
g77972 not n34714 ; n34714_not
g77973 not n47521 ; n47521_not
g77974 not n30673 ; n30673_not
g77975 not n50662 ; n50662_not
g77976 not n32536 ; n32536_not
g77977 not n35029 ; n35029_not
g77978 not n36073 ; n36073_not
g77979 not n49150 ; n49150_not
g77980 not n33355 ; n33355_not
g77981 not n33364 ; n33364_not
g77982 not n34840 ; n34840_not
g77983 not n30295 ; n30295_not
g77984 not n34390 ; n34390_not
g77985 not n50923 ; n50923_not
g77986 not n32914 ; n32914_not
g77987 not n31870 ; n31870_not
g77988 not n34912 ; n34912_not
g77989 not n30367 ; n30367_not
g77990 not n32923 ; n32923_not
g77991 not n36154 ; n36154_not
g77992 not n48115 ; n48115_not
g77993 not n31825 ; n31825_not
g77994 not n26605 ; n26605_not
g77995 not n48160 ; n48160_not
g77996 not n30439 ; n30439_not
g77997 not n31375 ; n31375_not
g77998 not n32941 ; n32941_not
g77999 not n31339 ; n31339_not
g78000 not n49006 ; n49006_not
g78001 not n26614 ; n26614_not
g78002 not n27091 ; n27091_not
g78003 not n37603 ; n37603_not
g78004 not n34804 ; n34804_not
g78005 not n29017 ; n29017_not
g78006 not n27271 ; n27271_not
g78007 not n32608 ; n32608_not
g78008 not n30268 ; n30268_not
g78009 not n30376 ; n30376_not
g78010 not n47350 ; n47350_not
g78011 not n34525 ; n34525_not
g78012 not n47107 ; n47107_not
g78013 not n30448 ; n30448_not
g78014 not n49015 ; n49015_not
g78015 not n31834 ; n31834_not
g78016 not n31762 ; n31762_not
g78017 not n36181 ; n36181_not
g78018 not n32590 ; n32590_not
g78019 not n37045 ; n37045_not
g78020 not n32905 ; n32905_not
g78021 not n37144 ; n37144_not
g78022 not n36163 ; n36163_not
g78023 not n50581 ; n50581_not
g78024 not n48106 ; n48106_not
g78025 not n26650 ; n26650_not
g78026 not n32680 ; n32680_not
g78027 not n29008 ; n29008_not
g78028 not n33049 ; n33049_not
g78029 not n37108 ; n37108_not
g78030 not n30547 ; n30547_not
g78031 not n33058 ; n33058_not
g78032 not n39070 ; n39070_not
g78033 not n36118 ; n36118_not
g78034 not n37900 ; n37900_not
g78035 not n30538 ; n30538_not
g78036 not n35920 ; n35920_not
g78037 not n36109 ; n36109_not
g78038 not n33067 ; n33067_not
g78039 not n29026 ; n29026_not
g78040 not n31096 ; n31096_not
g78041 not n33076 ; n33076_not
g78042 not n31807 ; n31807_not
g78043 not n26623 ; n26623_not
g78044 not n47800 ; n47800_not
g78045 not n48124 ; n48124_not
g78046 not n50590 ; n50590_not
g78047 not n38206 ; n38206_not
g78048 not n37036 ; n37036_not
g78049 not n26632 ; n26632_not
g78050 not n47332 ; n47332_not
g78051 not n27082 ; n27082_not
g78052 not n36136 ; n36136_not
g78053 not n32392 ; n32392_not
g78054 not n26641 ; n26641_not
g78055 not n48007 ; n48007_not
g78056 not n34534 ; n34534_not
g78057 not n31816 ; n31816_not
g78058 not n32725 ; n32725_not
g78059 not n50608 ; n50608_not
g78060 not n26542 ; n26542_not
g78061 not n32734 ; n32734_not
g78062 not n50257 ; n50257_not
g78063 not n31357 ; n31357_not
g78064 not n32653 ; n32653_not
g78065 not n50536 ; n50536_not
g78066 not n31852 ; n31852_not
g78067 not n37063 ; n37063_not
g78068 not n48142 ; n48142_not
g78069 not n37081 ; n37081_not
g78070 not n49042 ; n49042_not
g78071 not n30457 ; n30457_not
g78072 not n50527 ; n50527_not
g78073 not n38224 ; n38224_not
g78074 not n51841 ; n51841_not
g78075 not n38602 ; n38602_not
g78076 not n32644 ; n32644_not
g78077 not n48151 ; n48151_not
g78078 not n32806 ; n32806_not
g78079 not n31366 ; n31366_not
g78080 not n30394 ; n30394_not
g78081 not n32743 ; n32743_not
g78082 not n26524 ; n26524_not
g78083 not n38233 ; n38233_not
g78084 not n27145 ; n27145_not
g78085 not n50545 ; n50545_not
g78086 not n32752 ; n32752_not
g78087 not n50554 ; n50554_not
g78088 not n49060 ; n49060_not
g78089 not n31861 ; n31861_not
g78090 not n32761 ; n32761_not
g78091 not n26533 ; n26533_not
g78092 not n32770 ; n32770_not
g78093 not n37612 ; n37612_not
g78094 not n27136 ; n27136_not
g78095 not n49051 ; n49051_not
g78096 not n47242 ; n47242_not
g78097 not n52048 ; n52048_not
g78098 not n32842 ; n32842_not
g78099 not n49033 ; n49033_not
g78100 not n30385 ; n30385_not
g78101 not n50509 ; n50509_not
g78102 not n28081 ; n28081_not
g78103 not n32851 ; n32851_not
g78104 not n47116 ; n47116_not
g78105 not n36172 ; n36172_not
g78106 not n27253 ; n27253_not
g78107 not n32860 ; n32860_not
g78108 not n38242 ; n38242_not
g78109 not n49024 ; n49024_not
g78110 not n50248 ; n50248_not
g78111 not n34822 ; n34822_not
g78112 not n31348 ; n31348_not
g78113 not n52039 ; n52039_not
g78114 not n48133 ; n48133_not
g78115 not n34903 ; n34903_not
g78116 not n26551 ; n26551_not
g78117 not n30475 ; n30475_not
g78118 not n27127 ; n27127_not
g78119 not n36226 ; n36226_not
g78120 not n50563 ; n50563_not
g78121 not n32815 ; n32815_not
g78122 not n46405 ; n46405_not
g78123 not n32635 ; n32635_not
g78124 not n49420 ; n49420_not
g78125 not n26560 ; n26560_not
g78126 not n47251 ; n47251_not
g78127 not n27244 ; n27244_not
g78128 not n32824 ; n32824_not
g78129 not n50266 ; n50266_not
g78130 not n38215 ; n38215_not
g78131 not n28900 ; n28900_not
g78132 not n36217 ; n36217_not
g78133 not n37090 ; n37090_not
g78134 not n31843 ; n31843_not
g78135 not n32833 ; n32833_not
g78136 not n50572 ; n50572_not
g78137 not n50518 ; n50518_not
g78138 not n29062 ; n29062_not
g78139 not n29080 ; n29080_not
g78140 not n50635 ; n50635_not
g78141 not n30583 ; n30583_not
g78142 not n31294 ; n31294_not
g78143 not n32482 ; n32482_not
g78144 not n38170 ; n38170_not
g78145 not n39313 ; n39313_not
g78146 not n30592 ; n30592_not
g78147 not n34750 ; n34750_not
g78148 not n31771 ; n31771_not
g78149 not n33274 ; n33274_not
g78150 not n37441 ; n37441_not
g78151 not n50491 ; n50491_not
g78152 not n47710 ; n47710_not
g78153 not n47341 ; n47341_not
g78154 not n32491 ; n32491_not
g78155 not n33229 ; n33229_not
g78156 not n38260 ; n38260_not
g78157 not n50167 ; n50167_not
g78158 not n35632 ; n35632_not
g78159 not n47611 ; n47611_not
g78160 not n26731 ; n26731_not
g78161 not n27343 ; n27343_not
g78162 not n32473 ; n32473_not
g78163 not n31393 ; n31393_not
g78164 not n33238 ; n33238_not
g78165 not n28801 ; n28801_not
g78166 not n38008 ; n38008_not
g78167 not n26740 ; n26740_not
g78168 not n35641 ; n35641_not
g78169 not n30574 ; n30574_not
g78170 not n39322 ; n39322_not
g78171 not n32932 ; n32932_not
g78172 not n33247 ; n33247_not
g78173 not n31276 ; n31276_not
g78174 not n32518 ; n32518_not
g78175 not n48205 ; n48205_not
g78176 not n26812 ; n26812_not
g78177 not n30628 ; n30628_not
g78178 not n51940 ; n51940_not
g78179 not n48214 ; n48214_not
g78180 not n50653 ; n50653_not
g78181 not n32617 ; n32617_not
g78182 not n34732 ; n34732_not
g78183 not n26821 ; n26821_not
g78184 not n33382 ; n33382_not
g78185 not n31267 ; n31267_not
g78186 not n32527 ; n32527_not
g78187 not n30637 ; n30637_not
g78188 not n34615 ; n34615_not
g78189 not n33292 ; n33292_not
g78190 not n37126 ; n37126_not
g78191 not n47602 ; n47602_not
g78192 not n39304 ; n39304_not
g78193 not n34381 ; n34381_not
g78194 not n37450 ; n37450_not
g78195 not n31168 ; n31168_not
g78196 not n50644 ; n50644_not
g78197 not n34741 ; n34741_not
g78198 not n31285 ; n31285_not
g78199 not n32509 ; n32509_not
g78200 not n27361 ; n27361_not
g78201 not n34606 ; n34606_not
g78202 not n33337 ; n33337_not
g78203 not n26803 ; n26803_not
g78204 not n30619 ; n30619_not
g78205 not n32437 ; n32437_not
g78206 not n50293 ; n50293_not
g78207 not n50176 ; n50176_not
g78208 not n27055 ; n27055_not
g78209 not n33139 ; n33139_not
g78210 not n34552 ; n34552_not
g78211 not n39340 ; n39340_not
g78212 not n38251 ; n38251_not
g78213 not n36019 ; n36019_not
g78214 not n32662 ; n32662_not
g78215 not n33148 ; n33148_not
g78216 not n50626 ; n50626_not
g78217 not n36028 ; n36028_not
g78218 not n37513 ; n37513_not
g78219 not n27046 ; n27046_not
g78220 not n32446 ; n32446_not
g78221 not n34561 ; n34561_not
g78222 not n33157 ; n33157_not
g78223 not n46450 ; n46450_not
g78224 not n32419 ; n32419_not
g78225 not n30556 ; n30556_not
g78226 not n50617 ; n50617_not
g78227 not n33085 ; n33085_not
g78228 not n37531 ; n37531_not
g78229 not n33094 ; n33094_not
g78230 not n30358 ; n30358_not
g78231 not n36091 ; n36091_not
g78232 not n38620 ; n38620_not
g78233 not n28054 ; n28054_not
g78234 not n34543 ; n34543_not
g78235 not n31384 ; n31384_not
g78236 not n47233 ; n47233_not
g78237 not n32428 ; n32428_not
g78238 not n31087 ; n31087_not
g78239 not n27307 ; n27307_not
g78240 not n37018 ; n37018_not
g78241 not n31780 ; n31780_not
g78242 not n27037 ; n27037_not
g78243 not n47701 ; n47701_not
g78244 not n34570 ; n34570_not
g78245 not n47620 ; n47620_not
g78246 not n32464 ; n32464_not
g78247 not n36127 ; n36127_not
g78248 not n39331 ; n39331_not
g78249 not n31177 ; n31177_not
g78250 not n35623 ; n35623_not
g78251 not n26722 ; n26722_not
g78252 not n37504 ; n37504_not
g78253 not n36046 ; n36046_not
g78254 not n33166 ; n33166_not
g78255 not n33175 ; n33175_not
g78256 not n49510 ; n49510_not
g78257 not n26704 ; n26704_not
g78258 not n27325 ; n27325_not
g78259 not n33184 ; n33184_not
g78260 not n32455 ; n32455_not
g78261 not n31078 ; n31078_not
g78262 not n28144 ; n28144_not
g78263 not n28810 ; n28810_not
g78264 not n35614 ; n35614_not
g78265 not n33193 ; n33193_not
g78266 not n26713 ; n26713_not
g78267 not n50347 ; n50347_not
g78268 not n35218 ; n35218_not
g78269 not n34237 ; n34237_not
g78270 not n47206 ; n47206_not
g78271 not n35281 ; n35281_not
g78272 not n50833 ; n50833_not
g78273 not n29602 ; n29602_not
g78274 not n30934 ; n30934_not
g78275 not n34075 ; n34075_not
g78276 not n35227 ; n35227_not
g78277 not n50356 ; n50356_not
g78278 not n51094 ; n51094_not
g78279 not n38080 ; n38080_not
g78280 not n47305 ; n47305_not
g78281 not n28252 ; n28252_not
g78282 not n38800 ; n38800_not
g78283 not n32365 ; n32365_not
g78284 not n27613 ; n27613_not
g78285 not n28531 ; n28531_not
g78286 not n34246 ; n34246_not
g78287 not n30943 ; n30943_not
g78288 not n27604 ; n27604_not
g78289 not n28522 ; n28522_not
g78290 not n50815 ; n50815_not
g78291 not n34255 ; n34255_not
g78292 not n50365 ; n50365_not
g78293 not n48043 ; n48043_not
g78294 not n50068 ; n50068_not
g78295 not n30916 ; n30916_not
g78296 not n49312 ; n49312_not
g78297 not n47431 ; n47431_not
g78298 not n34219 ; n34219_not
g78299 not n34228 ; n34228_not
g78300 not n50095 ; n50095_not
g78301 not n34048 ; n34048_not
g78302 not n35272 ; n35272_not
g78303 not n34057 ; n34057_not
g78304 not n47215 ; n47215_not
g78305 not n28540 ; n28540_not
g78306 not n28243 ; n28243_not
g78307 not n34453 ; n34453_not
g78308 not n48430 ; n48430_not
g78309 not n50824 ; n50824_not
g78310 not n47125 ; n47125_not
g78311 not n50770 ; n50770_not
g78312 not n28504 ; n28504_not
g78313 not n50383 ; n50383_not
g78314 not n50761 ; n50761_not
g78315 not n33760 ; n33760_not
g78316 not n32068 ; n32068_not
g78317 not n34129 ; n34129_not
g78318 not n47422 ; n47422_not
g78319 not n50392 ; n50392_not
g78320 not n30961 ; n30961_not
g78321 not n51076 ; n51076_not
g78322 not n32149 ; n32149_not
g78323 not n37720 ; n37720_not
g78324 not n50806 ; n50806_not
g78325 not n38071 ; n38071_not
g78326 not n34138 ; n34138_not
g78327 not n51652 ; n51652_not
g78328 not n35263 ; n35263_not
g78329 not n50752 ; n50752_not
g78330 not n48322 ; n48322_not
g78331 not n34147 ; n34147_not
g78332 not n48421 ; n48421_not
g78333 not n28261 ; n28261_not
g78334 not n27622 ; n27622_not
g78335 not n51670 ; n51670_not
g78336 not n34093 ; n34093_not
g78337 not n34264 ; n34264_not
g78338 not n34435 ; n34435_not
g78339 not n50374 ; n50374_not
g78340 not n27640 ; n27640_not
g78341 not n34273 ; n34273_not
g78342 not n50077 ; n50077_not
g78343 not n29620 ; n29620_not
g78344 not n34426 ; n34426_not
g78345 not n35245 ; n35245_not
g78346 not n34282 ; n34282_not
g78347 not n50851 ; n50851_not
g78348 not n27631 ; n27631_not
g78349 not n28513 ; n28513_not
g78350 not n49303 ; n49303_not
g78351 not n34291 ; n34291_not
g78352 not n50185 ; n50185_not
g78353 not n31681 ; n31681_not
g78354 not n36613 ; n36613_not
g78355 not n28207 ; n28207_not
g78356 not n33562 ; n33562_not
g78357 not n47161 ; n47161_not
g78358 not n38413 ; n38413_not
g78359 not n48034 ; n48034_not
g78360 not n35191 ; n35191_not
g78361 not n29503 ; n29503_not
g78362 not n33751 ; n33751_not
g78363 not n35092 ; n35092_not
g78364 not n30880 ; n30880_not
g78365 not n29512 ; n29512_not
g78366 not n33571 ; n33571_not
g78367 not n29530 ; n29530_not
g78368 not n31951 ; n31951_not
g78369 not n35182 ; n35182_not
g78370 not n33544 ; n33544_not
g78371 not n36622 ; n36622_not
g78372 not n48313 ; n48313_not
g78373 not n30862 ; n30862_not
g78374 not n32374 ; n32374_not
g78375 not n35236 ; n35236_not
g78376 not n27460 ; n27460_not
g78377 not n38422 ; n38422_not
g78378 not n30907 ; n30907_not
g78379 not n33553 ; n33553_not
g78380 not n37522 ; n37522_not
g78381 not n33652 ; n33652_not
g78382 not n27910 ; n27910_not
g78383 not n30088 ; n30088_not
g78384 not n31483 ; n31483_not
g78385 not n30871 ; n30871_not
g78386 not n30079 ; n30079_not
g78387 not n27532 ; n27532_not
g78388 not n34165 ; n34165_not
g78389 not n36604 ; n36604_not
g78390 not n33616 ; n33616_not
g78391 not n35065 ; n35065_not
g78392 not n34174 ; n34174_not
g78393 not n31429 ; n31429_not
g78394 not n27550 ; n27550_not
g78395 not n37054 ; n37054_not
g78396 not n31960 ; n31960_not
g78397 not n34183 ; n34183_not
g78398 not n34480 ; n34480_not
g78399 not n28234 ; n28234_not
g78400 not n37801 ; n37801_not
g78401 not n34192 ; n34192_not
g78402 not n34471 ; n34471_not
g78403 not n33580 ; n33580_not
g78404 not n27901 ; n27901_not
g78405 not n35083 ; n35083_not
g78406 not n32095 ; n32095_not
g78407 not n35074 ; n35074_not
g78408 not n38404 ; n38404_not
g78409 not n32383 ; n32383_not
g78410 not n50086 ; n50086_not
g78411 not n47152 ; n47152_not
g78412 not n27514 ; n27514_not
g78413 not n37810 ; n37810_not
g78414 not n50158 ; n50158_not
g78415 not n34156 ; n34156_not
g78416 not n33625 ; n33625_not
g78417 not n35317 ; n35317_not
g78418 not n32329 ; n32329_not
g78419 not n38332 ; n38332_not
g78420 not n31474 ; n31474_not
g78421 not n51625 ; n51625_not
g78422 not n35326 ; n35326_not
g78423 not n27820 ; n27820_not
g78424 not n27721 ; n27721_not
g78425 not n29800 ; n29800_not
g78426 not n38026 ; n38026_not
g78427 not n38323 ; n38323_not
g78428 not n48340 ; n48340_not
g78429 not n50464 ; n50464_not
g78430 not n38341 ; n38341_not
g78431 not n28360 ; n28360_not
g78432 not n47404 ; n47404_not
g78433 not n50473 ; n50473_not
g78434 not n32176 ; n32176_not
g78435 not n35308 ; n35308_not
g78436 not n34345 ; n34345_not
g78437 not n38503 ; n38503_not
g78438 not n50941 ; n50941_not
g78439 not n28405 ; n28405_not
g78440 not n35353 ; n35353_not
g78441 not n27811 ; n27811_not
g78442 not n34318 ; n34318_not
g78443 not n38035 ; n38035_not
g78444 not n46531 ; n46531_not
g78445 not n35344 ; n35344_not
g78446 not n34327 ; n34327_not
g78447 not n28423 ; n28423_not
g78448 not n34336 ; n34336_not
g78449 not n47143 ; n47143_not
g78450 not n47413 ; n47413_not
g78451 not n35335 ; n35335_not
g78452 not n32185 ; n32185_not
g78453 not n37711 ; n37711_not
g78454 not n32338 ; n32338_not
g78455 not n38044 ; n38044_not
g78456 not n34309 ; n34309_not
g78457 not n28414 ; n28414_not
g78458 not n32194 ; n32194_not
g78459 not n50725 ; n50725_not
g78460 not n28315 ; n28315_not
g78461 not n50842 ; n50842_not
g78462 not n50428 ; n50428_not
g78463 not n38530 ; n38530_not
g78464 not n30952 ; n30952_not
g78465 not n50437 ; n50437_not
g78466 not n28324 ; n28324_not
g78467 not n51049 ; n51049_not
g78468 not n49330 ; n49330_not
g78469 not n50716 ; n50716_not
g78470 not n48403 ; n48403_not
g78471 not n48412 ; n48412_not
g78472 not n50419 ; n50419_not
g78473 not n50743 ; n50743_not
g78474 not n34408 ; n34408_not
g78475 not n27712 ; n27712_not
g78476 not n28306 ; n28306_not
g78477 not n31456 ; n31456_not
g78478 not n50734 ; n50734_not
g78479 not n51058 ; n51058_not
g78480 not n27730 ; n27730_not
g78481 not n32158 ; n32158_not
g78482 not n51643 ; n51643_not
g78483 not n50455 ; n50455_not
g78484 not n38053 ; n38053_not
g78485 not n29701 ; n29701_not
g78486 not n50914 ; n50914_not
g78487 not n47323 ; n47323_not
g78488 not n32167 ; n32167_not
g78489 not n34354 ; n34354_not
g78490 not n34066 ; n34066_not
g78491 not n48331 ; n48331_not
g78492 not n51634 ; n51634_not
g78493 not n29710 ; n29710_not
g78494 not n28432 ; n28432_not
g78495 not n31465 ; n31465_not
g78496 not n28450 ; n28450_not
g78497 not n50446 ; n50446_not
g78498 not n50707 ; n50707_not
g78499 not n38350 ; n38350_not
g78500 not n30763 ; n30763_not
g78501 not n35290 ; n35290_not
g78502 not n34363 ; n34363_not
g78503 not n48052 ; n48052_not
g78504 not n34372 ; n34372_not
g78505 not n28333 ; n28333_not
g78506 not n49402 ; n49402_not
g78507 not n47170 ; n47170_not
g78508 not n27703 ; n27703_not
g78509 not n28441 ; n28441_not
g78510 not n33463 ; n33463_not
g78511 not n38701 ; n38701_not
g78512 not n33454 ; n33454_not
g78513 not n27541 ; n27541_not
g78514 not n33706 ; n33706_not
g78515 not n33445 ; n33445_not
g78516 not n46603 ; n46603_not
g78517 not n30196 ; n30196_not
g78518 not n27523 ; n27523_not
g78519 not n30772 ; n30772_not
g78520 not n49240 ; n49240_not
g78521 not n33436 ; n33436_not
g78522 not n33517 ; n33517_not
g78523 not n33508 ; n33508_not
g78524 not n34813 ; n34813_not
g78525 not n29242 ; n29242_not
g78526 not n30565 ; n30565_not
g78527 not n33490 ; n33490_not
g78528 not n38134 ; n38134_not
g78529 not n38152 ; n38152_not
g78530 not n39160 ; n39160_not
g78531 not n33481 ; n33481_not
g78532 not n32572 ; n32572_not
g78533 not n33472 ; n33472_not
g78534 not n49222 ; n49222_not
g78535 not n45262 ; n45262_not
g78536 not n27442 ; n27442_not
g78537 not n38125 ; n38125_not
g78538 not n34444 ; n34444_not
g78539 not n33409 ; n33409_not
g78540 not n32563 ; n32563_not
g78541 not n27424 ; n27424_not
g78542 not n38710 ; n38710_not
g78543 not n32347 ; n32347_not
g78544 not n30790 ; n30790_not
g78545 not n33742 ; n33742_not
g78546 not n30178 ; n30178_not
g78547 not n39142 ; n39142_not
g78548 not n48610 ; n48610_not
g78549 not n27505 ; n27505_not
g78550 not n46612 ; n46612_not
g78551 not n29260 ; n29260_not
g78552 not n33427 ; n33427_not
g78553 not n36631 ; n36631_not
g78554 not n30781 ; n30781_not
g78555 not n49231 ; n49231_not
g78556 not n33418 ; n33418_not
g78557 not n51760 ; n51760_not
g78558 not n33724 ; n33724_not
g78559 not n30187 ; n30187_not
g78560 not n27451 ; n27451_not
g78561 not n30727 ; n30727_not
g78562 not n31915 ; n31915_not
g78563 not n34660 ; n34660_not
g78564 not n32059 ; n32059_not
g78565 not n51832 ; n51832_not
g78566 not n33607 ; n33607_not
g78567 not n51823 ; n51823_not
g78568 not n30718 ; n30718_not
g78569 not n33283 ; n33283_not
g78570 not n36523 ; n36523_not
g78571 not n49213 ; n49213_not
g78572 not n39205 ; n39205_not
g78573 not n48304 ; n48304_not
g78574 not n36541 ; n36541_not
g78575 not n46441 ; n46441_not
g78576 not n31717 ; n31717_not
g78577 not n31708 ; n31708_not
g78578 not n31924 ; n31924_not
g78579 not n36532 ; n36532_not
g78580 not n48016 ; n48016_not
g78581 not n33535 ; n33535_not
g78582 not n33661 ; n33661_not
g78583 not n33526 ; n33526_not
g78584 not n51805 ; n51805_not
g78585 not n31726 ; n31726_not
g78586 not n31438 ; n31438_not
g78587 not n30745 ; n30745_not
g78588 not n32581 ; n32581_not
g78589 not n50329 ; n50329_not
g78590 not n33634 ; n33634_not
g78591 not n35740 ; n35740_not
g78592 not n28045 ; n28045_not
g78593 not n30826 ; n30826_not
g78594 not n28603 ; n28603_not
g78595 not n48520 ; n48520_not
g78596 not n28135 ; n28135_not
g78597 not n27334 ; n27334_not
g78598 not n28036 ; n28036_not
g78599 not n35173 ; n35173_not
g78600 not n39025 ; n39025_not
g78601 not n48511 ; n48511_not
g78602 not n35155 ; n35155_not
g78603 not n35164 ; n35164_not
g78604 not n37702 ; n37702_not
g78605 not n27352 ; n27352_not
g78606 not n28621 ; n28621_not
g78607 not n39034 ; n39034_not
g78608 not n35605 ; n35605_not
g78609 not n28108 ; n28108_not
g78610 not n28612 ; n28612_not
g78611 not n38431 ; n38431_not
g78612 not n27280 ; n27280_not
g78613 not n28117 ; n28117_not
g78614 not n35146 ; n35146_not
g78615 not n38440 ; n38440_not
g78616 not n51067 ; n51067_not
g78617 not n27316 ; n27316_not
g78618 not n29350 ; n29350_not
g78619 not n31942 ; n31942_not
g78620 not n29440 ; n29440_not
g78621 not n27406 ; n27406_not
g78622 not n33670 ; n33670_not
g78623 not n35128 ; n35128_not
g78624 not n29341 ; n29341_not
g78625 not n28171 ; n28171_not
g78626 not n31159 ; n31159_not
g78627 not n51715 ; n51715_not
g78628 not n30853 ; n30853_not
g78629 not n28180 ; n28180_not
g78630 not n35119 ; n35119_not
g78631 not n39007 ; n39007_not
g78632 not n29404 ; n29404_not
g78633 not n30835 ; n30835_not
g78634 not n27370 ; n27370_not
g78635 not n29413 ; n29413_not
g78636 not n48502 ; n48502_not
g78637 not n30844 ; n30844_not
g78638 not n28009 ; n28009_not
g78639 not n28162 ; n28162_not
g78640 not n29422 ; n29422_not
g78641 not n47260 ; n47260_not
g78642 not n35137 ; n35137_not
g78643 not n29431 ; n29431_not
g78644 not n28018 ; n28018_not
g78645 not n35650 ; n35650_not
g78646 not n30169 ; n30169_not
g78647 not n31933 ; n31933_not
g78648 not n38512 ; n38512_not
g78649 not n50275 ; n50275_not
g78650 not n28216 ; n28216_not
g78651 not n51742 ; n51742_not
g78652 not n46621 ; n46621_not
g78653 not n31186 ; n31186_not
g78654 not n27262 ; n27262_not
g78655 not n28630 ; n28630_not
g78656 not n39052 ; n39052_not
g78657 not n27217 ; n27217_not
g78658 not n29332 ; n29332_not
g78659 not n28090 ; n28090_not
g78660 not n30736 ; n30736_not
g78661 not n30817 ; n30817_not
g78662 not n30808 ; n30808_not
g78663 not n51733 ; n51733_not
g78664 not n28063 ; n28063_not
g78665 not n33715 ; n33715_not
g78666 not n32293 ; n32293_not
g78667 not n53065 ; n53065_not
g78668 not n13771 ; n13771_not
g78669 not n13672 ; n13672_not
g78670 not n23563 ; n23563_not
g78671 not n23095 ; n23095_not
g78672 not n54631 ; n54631_not
g78673 not n22780 ; n22780_not
g78674 not n40924 ; n40924_not
g78675 not n23554 ; n23554_not
g78676 not n54244 ; n54244_not
g78677 not n13762 ; n13762_not
g78678 not n42292 ; n42292_not
g78679 not n10963 ; n10963_not
g78680 not n22771 ; n22771_not
g78681 not n10954 ; n10954_not
g78682 not n13681 ; n13681_not
g78683 not n23545 ; n23545_not
g78684 not n45253 ; n45253_not
g78685 not n10729 ; n10729_not
g78686 not n43903 ; n43903_not
g78687 not n22834 ; n22834_not
g78688 not n22762 ; n22762_not
g78689 not n23536 ; n23536_not
g78690 not n43651 ; n43651_not
g78691 not n13690 ; n13690_not
g78692 not n40852 ; n40852_not
g78693 not n22753 ; n22753_not
g78694 not n10657 ; n10657_not
g78695 not n23590 ; n23590_not
g78696 not n13627 ; n13627_not
g78697 not n56242 ; n56242_not
g78698 not n10990 ; n10990_not
g78699 not n22807 ; n22807_not
g78700 not n11197 ; n11197_not
g78701 not n13636 ; n13636_not
g78702 not n10666 ; n10666_not
g78703 not n13645 ; n13645_not
g78704 not n43660 ; n43660_not
g78705 not n10675 ; n10675_not
g78706 not n43912 ; n43912_not
g78707 not n13654 ; n13654_not
g78708 not n54640 ; n54640_not
g78709 not n10684 ; n10684_not
g78710 not n23581 ; n23581_not
g78711 not n54235 ; n54235_not
g78712 not n17740 ; n17740_not
g78713 not n56116 ; n56116_not
g78714 not n23572 ; n23572_not
g78715 not n10693 ; n10693_not
g78716 not n13663 ; n13663_not
g78717 not n42274 ; n42274_not
g78718 not n45217 ; n45217_not
g78719 not n44812 ; n44812_not
g78720 not n10765 ; n10765_not
g78721 not n23491 ; n23491_not
g78722 not n54613 ; n54613_not
g78723 not n53074 ; n53074_not
g78724 not n10774 ; n10774_not
g78725 not n10783 ; n10783_not
g78726 not n13735 ; n13735_not
g78727 not n54604 ; n54604_not
g78728 not n42265 ; n42265_not
g78729 not n10792 ; n10792_not
g78730 not n22708 ; n22708_not
g78731 not n10918 ; n10918_not
g78732 not n13717 ; n13717_not
g78733 not n23482 ; n23482_not
g78734 not n55900 ; n55900_not
g78735 not n10909 ; n10909_not
g78736 not n40942 ; n40942_not
g78737 not n52516 ; n52516_not
g78738 not n10819 ; n10819_not
g78739 not n11359 ; n11359_not
g78740 not n10828 ; n10828_not
g78741 not n23473 ; n23473_not
g78742 not n13708 ; n13708_not
g78743 not n11269 ; n11269_not
g78744 not n23527 ; n23527_not
g78745 not n54622 ; n54622_not
g78746 not n22843 ; n22843_not
g78747 not n22744 ; n22744_not
g78748 not n23518 ; n23518_not
g78749 not n22852 ; n22852_not
g78750 not n22735 ; n22735_not
g78751 not n10738 ; n10738_not
g78752 not n43291 ; n43291_not
g78753 not n23509 ; n23509_not
g78754 not n42283 ; n42283_not
g78755 not n10945 ; n10945_not
g78756 not n11278 ; n11278_not
g78757 not n40933 ; n40933_not
g78758 not n56233 ; n56233_not
g78759 not n10747 ; n10747_not
g78760 not n11287 ; n11287_not
g78761 not n22726 ; n22726_not
g78762 not n17713 ; n17713_not
g78763 not n13744 ; n13744_not
g78764 not n10756 ; n10756_not
g78765 not n11296 ; n11296_not
g78766 not n17704 ; n17704_not
g78767 not n22717 ; n22717_not
g78768 not n40825 ; n40825_not
g78769 not n13519 ; n13519_not
g78770 not n23365 ; n23365_not
g78771 not n10648 ; n10648_not
g78772 not n23743 ; n23743_not
g78773 not n23374 ; n23374_not
g78774 not n10639 ; n10639_not
g78775 not n13528 ; n13528_not
g78776 not n23734 ; n23734_not
g78777 not n23383 ; n23383_not
g78778 not n56026 ; n56026_not
g78779 not n40816 ; n40816_not
g78780 not n23392 ; n23392_not
g78781 not n42346 ; n42346_not
g78782 not n10594 ; n10594_not
g78783 not n41851 ; n41851_not
g78784 not n23716 ; n23716_not
g78785 not n23419 ; n23419_not
g78786 not n17803 ; n17803_not
g78787 not n23428 ; n23428_not
g78788 not n10585 ; n10585_not
g78789 not n23437 ; n23437_not
g78790 not n13537 ; n13537_not
g78791 not n23446 ; n23446_not
g78792 not n23806 ; n23806_not
g78793 not n13474 ; n13474_not
g78794 not n23257 ; n23257_not
g78795 not n23266 ; n23266_not
g78796 not n54190 ; n54190_not
g78797 not n23275 ; n23275_not
g78798 not n40870 ; n40870_not
g78799 not n23284 ; n23284_not
g78800 not n13483 ; n13483_not
g78801 not n13492 ; n13492_not
g78802 not n23293 ; n23293_not
g78803 not n42355 ; n42355_not
g78804 not n53047 ; n53047_not
g78805 not n41842 ; n41842_not
g78806 not n23329 ; n23329_not
g78807 not n54712 ; n54712_not
g78808 not n13861 ; n13861_not
g78809 not n13852 ; n13852_not
g78810 not n23761 ; n23761_not
g78811 not n23338 ; n23338_not
g78812 not n23347 ; n23347_not
g78813 not n23356 ; n23356_not
g78814 not n54703 ; n54703_not
g78815 not n10567 ; n10567_not
g78816 not n10576 ; n10576_not
g78817 not n40807 ; n40807_not
g78818 not n23644 ; n23644_not
g78819 not n13573 ; n13573_not
g78820 not n42328 ; n42328_not
g78821 not n13582 ; n13582_not
g78822 not n13816 ; n13816_not
g78823 not n13591 ; n13591_not
g78824 not n40915 ; n40915_not
g78825 not n11179 ; n11179_not
g78826 not n13807 ; n13807_not
g78827 not n13609 ; n13609_not
g78828 not n23626 ; n23626_not
g78829 not n11188 ; n11188_not
g78830 not n54226 ; n54226_not
g78831 not n42319 ; n42319_not
g78832 not n13618 ; n13618_not
g78833 not n13546 ; n13546_not
g78834 not n23455 ; n23455_not
g78835 not n23464 ; n23464_not
g78836 not n42337 ; n42337_not
g78837 not n10558 ; n10558_not
g78838 not n10549 ; n10549_not
g78839 not n13834 ; n13834_not
g78840 not n53056 ; n53056_not
g78841 not n23671 ; n23671_not
g78842 not n13555 ; n13555_not
g78843 not n40906 ; n40906_not
g78844 not n13564 ; n13564_not
g78845 not n11098 ; n11098_not
g78846 not n56251 ; n56251_not
g78847 not n23653 ; n23653_not
g78848 not n22429 ; n22429_not
g78849 not n11557 ; n11557_not
g78850 not n23194 ; n23194_not
g78851 not n54532 ; n54532_not
g78852 not n42184 ; n42184_not
g78853 not n53128 ; n53128_not
g78854 not n41941 ; n41941_not
g78855 not n23185 ; n23185_not
g78856 not n44920 ; n44920_not
g78857 not n23176 ; n23176_not
g78858 not n11575 ; n11575_not
g78859 not n22393 ; n22393_not
g78860 not n23167 ; n23167_not
g78861 not n18415 ; n18415_not
g78862 not n43327 ; n43327_not
g78863 not n18424 ; n18424_not
g78864 not n22384 ; n22384_not
g78865 not n23158 ; n23158_not
g78866 not n42175 ; n42175_not
g78867 not n22375 ; n22375_not
g78868 not n22492 ; n22492_not
g78869 not n42193 ; n42193_not
g78870 not n22483 ; n22483_not
g78871 not n41932 ; n41932_not
g78872 not n53119 ; n53119_not
g78873 not n22474 ; n22474_not
g78874 not n23248 ; n23248_not
g78875 not n22465 ; n22465_not
g78876 not n23239 ; n23239_not
g78877 not n22456 ; n22456_not
g78878 not n22447 ; n22447_not
g78879 not n11548 ; n11548_not
g78880 not n22438 ; n22438_not
g78881 not n44911 ; n44911_not
g78882 not n22339 ; n22339_not
g78883 not n22348 ; n22348_not
g78884 not n23059 ; n23059_not
g78885 not n22357 ; n22357_not
g78886 not n22366 ; n22366_not
g78887 not n42157 ; n42157_not
g78888 not n43336 ; n43336_not
g78889 not n53137 ; n53137_not
g78890 not n11647 ; n11647_not
g78891 not n23149 ; n23149_not
g78892 not n11593 ; n11593_not
g78893 not n18442 ; n18442_not
g78894 not n42166 ; n42166_not
g78895 not n43633 ; n43633_not
g78896 not n23068 ; n23068_not
g78897 not n18460 ; n18460_not
g78898 not n56224 ; n56224_not
g78899 not n23077 ; n23077_not
g78900 not n11629 ; n11629_not
g78901 not n23086 ; n23086_not
g78902 not n11638 ; n11638_not
g78903 not n21547 ; n21547_not
g78904 not n52507 ; n52507_not
g78905 not n22654 ; n22654_not
g78906 not n13168 ; n13168_not
g78907 not n17650 ; n17650_not
g78908 not n22645 ; n22645_not
g78909 not n42229 ; n42229_not
g78910 not n43309 ; n43309_not
g78911 not n22636 ; n22636_not
g78912 not n54280 ; n54280_not
g78913 not n10873 ; n10873_not
g78914 not n22627 ; n22627_not
g78915 not n53092 ; n53092_not
g78916 not n43642 ; n43642_not
g78917 not n40960 ; n40960_not
g78918 not n54550 ; n54550_not
g78919 not n22618 ; n22618_not
g78920 not n40780 ; n40780_not
g78921 not n13177 ; n13177_not
g78922 not n11368 ; n11368_not
g78923 not n42256 ; n42256_not
g78924 not n22690 ; n22690_not
g78925 not n10837 ; n10837_not
g78926 not n53083 ; n53083_not
g78927 not n22681 ; n22681_not
g78928 not n11377 ; n11377_not
g78929 not n42247 ; n42247_not
g78930 not n10846 ; n10846_not
g78931 not n40951 ; n40951_not
g78932 not n22672 ; n22672_not
g78933 not n11386 ; n11386_not
g78934 not n54271 ; n54271_not
g78935 not n42238 ; n42238_not
g78936 not n22663 ; n22663_not
g78937 not n11395 ; n11395_not
g78938 not n13186 ; n13186_not
g78939 not n22564 ; n22564_not
g78940 not n43318 ; n43318_not
g78941 not n22555 ; n22555_not
g78942 not n18352 ; n18352_not
g78943 not n22546 ; n22546_not
g78944 not n54541 ; n54541_not
g78945 not n11485 ; n11485_not
g78946 not n22537 ; n22537_not
g78947 not n22528 ; n22528_not
g78948 not n22519 ; n22519_not
g78949 not n40762 ; n40762_not
g78950 not n18370 ; n18370_not
g78951 not n18316 ; n18316_not
g78952 not n22609 ; n22609_not
g78953 not n18325 ; n18325_not
g78954 not n22924 ; n22924_not
g78955 not n40771 ; n40771_not
g78956 not n22591 ; n22591_not
g78957 not n18334 ; n18334_not
g78958 not n11458 ; n11458_not
g78959 not n22933 ; n22933_not
g78960 not n22582 ; n22582_not
g78961 not n11467 ; n11467_not
g78962 not n41923 ; n41923_not
g78963 not n22942 ; n22942_not
g78964 not n22573 ; n22573_not
g78965 not n24751 ; n24751_not
g78966 not n17434 ; n17434_not
g78967 not n13780 ; n13780_not
g78968 not n24670 ; n24670_not
g78969 not n23950 ; n23950_not
g78970 not n42652 ; n42652_not
g78971 not n17443 ; n17443_not
g78972 not n24742 ; n24742_not
g78973 not n23941 ; n23941_not
g78974 not n40555 ; n40555_not
g78975 not n42643 ; n42643_not
g78976 not n24733 ; n24733_not
g78977 not n16804 ; n16804_not
g78978 not n17047 ; n17047_not
g78979 not n10495 ; n10495_not
g78980 not n23932 ; n23932_not
g78981 not n17452 ; n17452_not
g78982 not n16813 ; n16813_not
g78983 not n17038 ; n17038_not
g78984 not n56305 ; n56305_not
g78985 not n10486 ; n10486_not
g78986 not n24724 ; n24724_not
g78987 not n23923 ; n23923_not
g78988 not n17461 ; n17461_not
g78989 not n16822 ; n16822_not
g78990 not n24715 ; n24715_not
g78991 not n17470 ; n17470_not
g78992 not n23914 ; n23914_not
g78993 not n17380 ; n17380_not
g78994 not n24823 ; n24823_not
g78995 not n24634 ; n24634_not
g78996 not n44344 ; n44344_not
g78997 not n16741 ; n16741_not
g78998 not n42625 ; n42625_not
g78999 not n24814 ; n24814_not
g79000 not n55009 ; n55009_not
g79001 not n40519 ; n40519_not
g79002 not n16750 ; n16750_not
g79003 not n24805 ; n24805_not
g79004 not n17074 ; n17074_not
g79005 not n52750 ; n52750_not
g79006 not n45082 ; n45082_not
g79007 not n40528 ; n40528_not
g79008 not n17407 ; n17407_not
g79009 not n40537 ; n40537_not
g79010 not n17416 ; n17416_not
g79011 not n42661 ; n42661_not
g79012 not n24661 ; n24661_not
g79013 not n56314 ; n56314_not
g79014 not n24760 ; n24760_not
g79015 not n40546 ; n40546_not
g79016 not n17425 ; n17425_not
g79017 not n42634 ; n42634_not
g79018 not n17533 ; n17533_not
g79019 not n54082 ; n54082_not
g79020 not n17542 ; n17542_not
g79021 not n52813 ; n52813_not
g79022 not n40582 ; n40582_not
g79023 not n16903 ; n16903_not
g79024 not n54910 ; n54910_not
g79025 not n17551 ; n17551_not
g79026 not n24643 ; n24643_not
g79027 not n16912 ; n16912_not
g79028 not n44326 ; n44326_not
g79029 not n24625 ; n24625_not
g79030 not n24616 ; n24616_not
g79031 not n17560 ; n17560_not
g79032 not n24049 ; n24049_not
g79033 not n16921 ; n16921_not
g79034 not n24058 ; n24058_not
g79035 not n24067 ; n24067_not
g79036 not n24076 ; n24076_not
g79037 not n54901 ; n54901_not
g79038 not n52822 ; n52822_not
g79039 not n54091 ; n54091_not
g79040 not n24085 ; n24085_not
g79041 not n43804 ; n43804_not
g79042 not n16930 ; n16930_not
g79043 not n24706 ; n24706_not
g79044 not n40564 ; n40564_not
g79045 not n16831 ; n16831_not
g79046 not n17029 ; n17029_not
g79047 not n44353 ; n44353_not
g79048 not n23905 ; n23905_not
g79049 not n10477 ; n10477_not
g79050 not n52804 ; n52804_not
g79051 not n16840 ; n16840_not
g79052 not n42616 ; n42616_not
g79053 not n17506 ; n17506_not
g79054 not n40573 ; n40573_not
g79055 not n17515 ; n17515_not
g79056 not n17524 ; n17524_not
g79057 not n24544 ; n24544_not
g79058 not n24184 ; n24184_not
g79059 not n10189 ; n10189_not
g79060 not n17263 ; n17263_not
g79061 not n52705 ; n52705_not
g79062 not n24175 ; n24175_not
g79063 not n16624 ; n16624_not
g79064 not n10198 ; n10198_not
g79065 not n17272 ; n17272_not
g79066 not n40465 ; n40465_not
g79067 not n45244 ; n45244_not
g79068 not n24166 ; n24166_not
g79069 not n55045 ; n55045_not
g79070 not n56332 ; n56332_not
g79071 not n16633 ; n16633_not
g79072 not n24157 ; n24157_not
g79073 not n17281 ; n17281_not
g79074 not n42706 ; n42706_not
g79075 not n24148 ; n24148_not
g79076 not n40168 ; n40168_not
g79077 not n24940 ; n24940_not
g79078 not n56323 ; n56323_not
g79079 not n10279 ; n10279_not
g79080 not n10288 ; n10288_not
g79081 not n40474 ; n40474_not
g79082 not n56350 ; n56350_not
g79083 not n17227 ; n17227_not
g79084 not n14356 ; n14356_not
g79085 not n14338 ; n14338_not
g79086 not n25057 ; n25057_not
g79087 not n24256 ; n24256_not
g79088 not n17164 ; n17164_not
g79089 not n17236 ; n17236_not
g79090 not n25048 ; n25048_not
g79091 not n55054 ; n55054_not
g79092 not n17245 ; n17245_not
g79093 not n24247 ; n24247_not
g79094 not n25039 ; n25039_not
g79095 not n24238 ; n24238_not
g79096 not n14347 ; n14347_not
g79097 not n42715 ; n42715_not
g79098 not n24229 ; n24229_not
g79099 not n40447 ; n40447_not
g79100 not n24526 ; n24526_not
g79101 not n56341 ; n56341_not
g79102 not n44371 ; n44371_not
g79103 not n16606 ; n16606_not
g79104 not n17254 ; n17254_not
g79105 not n24535 ; n24535_not
g79106 not n24193 ; n24193_not
g79107 not n16615 ; n16615_not
g79108 not n40456 ; n40456_not
g79109 not n24094 ; n24094_not
g79110 not n40492 ; n40492_not
g79111 not n16705 ; n16705_not
g79112 not n10387 ; n10387_not
g79113 not n10396 ; n10396_not
g79114 not n52732 ; n52732_not
g79115 not n17353 ; n17353_not
g79116 not n16714 ; n16714_not
g79117 not n17362 ; n17362_not
g79118 not n10459 ; n10459_not
g79119 not n52741 ; n52741_not
g79120 not n16723 ; n16723_not
g79121 not n24850 ; n24850_not
g79122 not n17092 ; n17092_not
g79123 not n17371 ; n17371_not
g79124 not n24841 ; n24841_not
g79125 not n16732 ; n16732_not
g79126 not n17083 ; n17083_not
g79127 not n24832 ; n24832_not
g79128 not n16642 ; n16642_not
g79129 not n17137 ; n17137_not
g79130 not n17290 ; n17290_not
g79131 not n10297 ; n10297_not
g79132 not n16651 ; n16651_not
g79133 not n24139 ; n24139_not
g79134 not n17128 ; n17128_not
g79135 not n24931 ; n24931_not
g79136 not n24571 ; n24571_not
g79137 not n16660 ; n16660_not
g79138 not n40159 ; n40159_not
g79139 not n17308 ; n17308_not
g79140 not n24922 ; n24922_not
g79141 not n52714 ; n52714_not
g79142 not n40483 ; n40483_not
g79143 not n17119 ; n17119_not
g79144 not n17317 ; n17317_not
g79145 not n17326 ; n17326_not
g79146 not n24913 ; n24913_not
g79147 not n24580 ; n24580_not
g79148 not n10369 ; n10369_not
g79149 not n17335 ; n17335_not
g79150 not n24904 ; n24904_not
g79151 not n17344 ; n17344_not
g79152 not n55027 ; n55027_not
g79153 not n52723 ; n52723_not
g79154 not n13942 ; n13942_not
g79155 not n42409 ; n42409_not
g79156 not n45091 ; n45091_not
g79157 not n56260 ; n56260_not
g79158 not n41806 ; n41806_not
g79159 not n13951 ; n13951_not
g79160 not n13348 ; n13348_not
g79161 not n23824 ; n23824_not
g79162 not n23833 ; n23833_not
g79163 not n13357 ; n13357_not
g79164 not n13366 ; n13366_not
g79165 not n42391 ; n42391_not
g79166 not n23842 ; n23842_not
g79167 not n52561 ; n52561_not
g79168 not n13375 ; n13375_not
g79169 not n23707 ; n23707_not
g79170 not n17812 ; n17812_not
g79171 not n42445 ; n42445_not
g79172 not n52903 ; n52903_not
g79173 not n42436 ; n42436_not
g79174 not n54136 ; n54136_not
g79175 not n17830 ; n17830_not
g79176 not n10882 ; n10882_not
g79177 not n52912 ; n52912_not
g79178 not n54811 ; n54811_not
g79179 not n40717 ; n40717_not
g79180 not n23752 ; n23752_not
g79181 not n42418 ; n42418_not
g79182 not n16543 ; n16543_not
g79183 not n40726 ; n40726_not
g79184 not n52606 ; n52606_not
g79185 not n52921 ; n52921_not
g79186 not n54802 ; n54802_not
g79187 not n52930 ; n52930_not
g79188 not n54145 ; n54145_not
g79189 not n40744 ; n40744_not
g79190 not n54154 ; n54154_not
g79191 not n54181 ; n54181_not
g79192 not n23851 ; n23851_not
g79193 not n42373 ; n42373_not
g79194 not n41833 ; n41833_not
g79195 not n13438 ; n13438_not
g79196 not n54730 ; n54730_not
g79197 not n10972 ; n10972_not
g79198 not n44362 ; n44362_not
g79199 not n13447 ; n13447_not
g79200 not n42364 ; n42364_not
g79201 not n13456 ; n13456_not
g79202 not n13465 ; n13465_not
g79203 not n54721 ; n54721_not
g79204 not n10927 ; n10927_not
g79205 not n13384 ; n13384_not
g79206 not n52552 ; n52552_not
g79207 not n13924 ; n13924_not
g79208 not n42382 ; n42382_not
g79209 not n13393 ; n13393_not
g79210 not n45226 ; n45226_not
g79211 not n40834 ; n40834_not
g79212 not n52543 ; n52543_not
g79213 not n53029 ; n53029_not
g79214 not n40843 ; n40843_not
g79215 not n44803 ; n44803_not
g79216 not n13906 ; n13906_not
g79217 not n53038 ; n53038_not
g79218 not n13429 ; n13429_not
g79219 not n24508 ; n24508_not
g79220 not n42535 ; n42535_not
g79221 not n24265 ; n24265_not
g79222 not n42526 ; n42526_not
g79223 not n24490 ; n24490_not
g79224 not n24274 ; n24274_not
g79225 not n24283 ; n24283_not
g79226 not n24481 ; n24481_not
g79227 not n24292 ; n24292_not
g79228 not n24319 ; n24319_not
g79229 not n24463 ; n24463_not
g79230 not n42580 ; n42580_not
g79231 not n42571 ; n42571_not
g79232 not n13825 ; n13825_not
g79233 not n40591 ; n40591_not
g79234 not n54109 ; n54109_not
g79235 not n17605 ; n17605_not
g79236 not n56008 ; n56008_not
g79237 not n44335 ; n44335_not
g79238 not n24553 ; n24553_not
g79239 not n17623 ; n17623_not
g79240 not n42553 ; n42553_not
g79241 not n17632 ; n17632_not
g79242 not n42490 ; n42490_not
g79243 not n52651 ; n52651_not
g79244 not n13870 ; n13870_not
g79245 not n23617 ; n23617_not
g79246 not n52840 ; n52840_not
g79247 not n42481 ; n42481_not
g79248 not n40618 ; n40618_not
g79249 not n40078 ; n40078_not
g79250 not n45235 ; n45235_not
g79251 not n52642 ; n52642_not
g79252 not n40636 ; n40636_not
g79253 not n23662 ; n23662_not
g79254 not n43831 ; n43831_not
g79255 not n52633 ; n52633_not
g79256 not n40654 ; n40654_not
g79257 not n44443 ; n44443_not
g79258 not n42463 ; n42463_not
g79259 not n13915 ; n13915_not
g79260 not n40672 ; n40672_not
g79261 not n55810 ; n55810_not
g79262 not n40681 ; n40681_not
g79263 not n56017 ; n56017_not
g79264 not n54820 ; n54820_not
g79265 not n24328 ; n24328_not
g79266 not n43813 ; n43813_not
g79267 not n24337 ; n24337_not
g79268 not n42508 ; n42508_not
g79269 not n24346 ; n24346_not
g79270 not n24445 ; n24445_not
g79271 not n24355 ; n24355_not
g79272 not n24364 ; n24364_not
g79273 not n24436 ; n24436_not
g79274 not n24373 ; n24373_not
g79275 not n24382 ; n24382_not
g79276 not n24391 ; n24391_not
g79277 not n17722 ; n17722_not
g79278 not n52831 ; n52831_not
g79279 not n24418 ; n24418_not
g79280 not n24409 ; n24409_not
g79281 not n40609 ; n40609_not
g79282 not n20269 ; n20269_not
g79283 not n45181 ; n45181_not
g79284 not n19090 ; n19090_not
g79285 not n41707 ; n41707_not
g79286 not n11953 ; n11953_not
g79287 not n41293 ; n41293_not
g79288 not n41095 ; n41095_not
g79289 not n41086 ; n41086_not
g79290 not n11944 ; n11944_not
g79291 not n19108 ; n19108_not
g79292 not n41077 ; n41077_not
g79293 not n11935 ; n11935_not
g79294 not n19117 ; n19117_not
g79295 not n41716 ; n41716_not
g79296 not n20665 ; n20665_not
g79297 not n41068 ; n41068_not
g79298 not n11926 ; n11926_not
g79299 not n41059 ; n41059_not
g79300 not n20674 ; n20674_not
g79301 not n20197 ; n20197_not
g79302 not n20683 ; n20683_not
g79303 not n20188 ; n20188_not
g79304 not n11917 ; n11917_not
g79305 not n20179 ; n20179_not
g79306 not n19135 ; n19135_not
g79307 not n53416 ; n53416_not
g79308 not n11908 ; n11908_not
g79309 not n20539 ; n20539_not
g79310 not n41158 ; n41158_not
g79311 not n20548 ; n20548_not
g79312 not n12583 ; n12583_not
g79313 not n19063 ; n19063_not
g79314 not n19072 ; n19072_not
g79315 not n11962 ; n11962_not
g79316 not n20395 ; n20395_not
g79317 not n41149 ; n41149_not
g79318 not n20386 ; n20386_not
g79319 not n41275 ; n41275_not
g79320 not n20575 ; n20575_not
g79321 not n20377 ; n20377_not
g79322 not n20368 ; n20368_not
g79323 not n20584 ; n20584_not
g79324 not n20359 ; n20359_not
g79325 not n20593 ; n20593_not
g79326 not n43570 ; n43570_not
g79327 not n12592 ; n12592_not
g79328 not n53371 ; n53371_not
g79329 not n53380 ; n53380_not
g79330 not n43444 ; n43444_not
g79331 not n20296 ; n20296_not
g79332 not n20287 ; n20287_not
g79333 not n54163 ; n54163_not
g79334 not n20629 ; n20629_not
g79335 not n20278 ; n20278_not
g79336 not n20638 ; n20638_not
g79337 not n20755 ; n20755_not
g79338 not n11872 ; n11872_not
g79339 not n20773 ; n20773_not
g79340 not n45136 ; n45136_not
g79341 not n11863 ; n11863_not
g79342 not n20764 ; n20764_not
g79343 not n12637 ; n12637_not
g79344 not n20737 ; n20737_not
g79345 not n20089 ; n20089_not
g79346 not n11854 ; n11854_not
g79347 not n41761 ; n41761_not
g79348 not n20098 ; n20098_not
g79349 not n20719 ; n20719_not
g79350 not n11845 ; n11845_not
g79351 not n20692 ; n20692_not
g79352 not n11836 ; n11836_not
g79353 not n19207 ; n19207_not
g79354 not n54073 ; n54073_not
g79355 not n41383 ; n41383_not
g79356 not n56152 ; n56152_not
g79357 not n53425 ; n53425_not
g79358 not n54118 ; n54118_not
g79359 not n41338 ; n41338_not
g79360 not n41725 ; n41725_not
g79361 not n11890 ; n11890_not
g79362 not n41347 ; n41347_not
g79363 not n12619 ; n12619_not
g79364 not n19153 ; n19153_not
g79365 not n41860 ; n41860_not
g79366 not n20728 ; n20728_not
g79367 not n19162 ; n19162_not
g79368 not n41734 ; n41734_not
g79369 not n53443 ; n53443_not
g79370 not n41365 ; n41365_not
g79371 not n11881 ; n11881_not
g79372 not n12628 ; n12628_not
g79373 not n41743 ; n41743_not
g79374 not n19180 ; n19180_not
g79375 not n20791 ; n20791_not
g79376 not n43453 ; n43453_not
g79377 not n20782 ; n20782_not
g79378 not n41752 ; n41752_not
g79379 not n20818 ; n20818_not
g79380 not n20827 ; n20827_not
g79381 not n20836 ; n20836_not
g79382 not n20845 ; n20845_not
g79383 not n20854 ; n20854_not
g79384 not n20863 ; n20863_not
g79385 not n20872 ; n20872_not
g79386 not n21484 ; n21484_not
g79387 not n20881 ; n20881_not
g79388 not n20890 ; n20890_not
g79389 not n21475 ; n21475_not
g79390 not n41662 ; n41662_not
g79391 not n19018 ; n19018_not
g79392 not n20908 ; n20908_not
g79393 not n20917 ; n20917_not
g79394 not n20926 ; n20926_not
g79395 not n21457 ; n21457_not
g79396 not n54208 ; n54208_not
g79397 not n21493 ; n21493_not
g79398 not n41644 ; n41644_not
g79399 not n41905 ; n41905_not
g79400 not n53326 ; n53326_not
g79401 not n41653 ; n41653_not
g79402 not n13096 ; n13096_not
g79403 not n53335 ; n53335_not
g79404 not n18343 ; n18343_not
g79405 not n20809 ; n20809_not
g79406 not n19009 ; n19009_not
g79407 not n21529 ; n21529_not
g79408 not n41671 ; n41671_not
g79409 not n21349 ; n21349_not
g79410 not n21169 ; n21169_not
g79411 not n21178 ; n21178_not
g79412 not n21187 ; n21187_not
g79413 not n21196 ; n21196_not
g79414 not n56161 ; n56161_not
g79415 not n21295 ; n21295_not
g79416 not n41257 ; n41257_not
g79417 not n19045 ; n19045_not
g79418 not n21277 ; n21277_not
g79419 not n21268 ; n21268_not
g79420 not n21259 ; n21259_not
g79421 not n41176 ; n41176_not
g79422 not n11980 ; n11980_not
g79423 not n13078 ; n13078_not
g79424 not n20485 ; n20485_not
g79425 not n41167 ; n41167_not
g79426 not n53353 ; n53353_not
g79427 not n20476 ; n20476_not
g79428 not n20467 ; n20467_not
g79429 not n20458 ; n20458_not
g79430 not n13069 ; n13069_not
g79431 not n20449 ; n20449_not
g79432 not n41680 ; n41680_not
g79433 not n20935 ; n20935_not
g79434 not n20944 ; n20944_not
g79435 not n20953 ; n20953_not
g79436 not n21439 ; n21439_not
g79437 not n20962 ; n20962_not
g79438 not n41194 ; n41194_not
g79439 not n20971 ; n20971_not
g79440 not n45190 ; n45190_not
g79441 not n20980 ; n20980_not
g79442 not n13087 ; n13087_not
g79443 not n41248 ; n41248_not
g79444 not n19027 ; n19027_not
g79445 not n43822 ; n43822_not
g79446 not n41185 ; n41185_not
g79447 not n21394 ; n21394_not
g79448 not n21385 ; n21385_not
g79449 not n12574 ; n12574_not
g79450 not n21079 ; n21079_not
g79451 not n21088 ; n21088_not
g79452 not n21367 ; n21367_not
g79453 not n21097 ; n21097_not
g79454 not n12097 ; n12097_not
g79455 not n53290 ; n53290_not
g79456 not n53470 ; n53470_not
g79457 not n44830 ; n44830_not
g79458 not n12088 ; n12088_not
g79459 not n12835 ; n12835_not
g79460 not n56053 ; n56053_not
g79461 not n56107 ; n56107_not
g79462 not n41527 ; n41527_not
g79463 not n12826 ; n12826_not
g79464 not n12718 ; n12718_not
g79465 not n53461 ; n53461_not
g79466 not n41536 ; n41536_not
g79467 not n12817 ; n12817_not
g79468 not n12727 ; n12727_not
g79469 not n41545 ; n41545_not
g79470 not n19171 ; n19171_not
g79471 not n12808 ; n12808_not
g79472 not n55243 ; n55243_not
g79473 not n43543 ; n43543_not
g79474 not n41554 ; n41554_not
g79475 not n19900 ; n19900_not
g79476 not n19252 ; n19252_not
g79477 not n41770 ; n41770_not
g79478 not n12880 ; n12880_not
g79479 not n53506 ; n53506_not
g79480 not n56134 ; n56134_not
g79481 not n45172 ; n45172_not
g79482 not n19243 ; n19243_not
g79483 not n41491 ; n41491_not
g79484 not n43480 ; n43480_not
g79485 not n12871 ; n12871_not
g79486 not n12862 ; n12862_not
g79487 not n53281 ; n53281_not
g79488 not n41392 ; n41392_not
g79489 not n56125 ; n56125_not
g79490 not n19216 ; n19216_not
g79491 not n12853 ; n12853_not
g79492 not n41509 ; n41509_not
g79493 not n41266 ; n41266_not
g79494 not n12844 ; n12844_not
g79495 not n12709 ; n12709_not
g79496 not n43552 ; n43552_not
g79497 not n41518 ; n41518_not
g79498 not n41590 ; n41590_not
g79499 not n12556 ; n12556_not
g79500 not n12178 ; n12178_not
g79501 not n43507 ; n43507_not
g79502 not n12736 ; n12736_not
g79503 not n19810 ; n19810_not
g79504 not n41608 ; n41608_not
g79505 not n12691 ; n12691_not
g79506 not n19081 ; n19081_not
g79507 not n41617 ; n41617_not
g79508 not n43516 ; n43516_not
g79509 not n12673 ; n12673_not
g79510 not n12664 ; n12664_not
g79511 not n41635 ; n41635_not
g79512 not n41626 ; n41626_not
g79513 not n12646 ; n12646_not
g79514 not n12790 ; n12790_not
g79515 not n56062 ; n56062_not
g79516 not n12781 ; n12781_not
g79517 not n41563 ; n41563_not
g79518 not n53434 ; n53434_not
g79519 not n41572 ; n41572_not
g79520 not n43534 ; n43534_not
g79521 not n19126 ; n19126_not
g79522 not n41356 ; n41356_not
g79523 not n53344 ; n53344_not
g79524 not n56080 ; n56080_not
g79525 not n41581 ; n41581_not
g79526 not n43525 ; n43525_not
g79527 not n12547 ; n12547_not
g79528 not n12754 ; n12754_not
g79529 not n12961 ; n12961_not
g79530 not n20557 ; n20557_not
g79531 not n19225 ; n19225_not
g79532 not n12952 ; n12952_not
g79533 not n43462 ; n43462_not
g79534 not n11782 ; n11782_not
g79535 not n20494 ; n20494_not
g79536 not n56035 ; n56035_not
g79537 not n11773 ; n11773_not
g79538 not n11827 ; n11827_not
g79539 not n11818 ; n11818_not
g79540 not n12970 ; n12970_not
g79541 not n20647 ; n20647_not
g79542 not n11809 ; n11809_not
g79543 not n11791 ; n11791_not
g79544 not n56143 ; n56143_not
g79545 not n53533 ; n53533_not
g79546 not n11692 ; n11692_not
g79547 not n12916 ; n12916_not
g79548 not n11683 ; n11683_not
g79549 not n12907 ; n12907_not
g79550 not n41455 ; n41455_not
g79551 not n53542 ; n53542_not
g79552 not n43471 ; n43471_not
g79553 not n11674 ; n11674_not
g79554 not n11665 ; n11665_not
g79555 not n11656 ; n11656_not
g79556 not n41464 ; n41464_not
g79557 not n12682 ; n12682_not
g79558 not n41473 ; n41473_not
g79559 not n53524 ; n53524_not
g79560 not n43561 ; n43561_not
g79561 not n53515 ; n53515_not
g79562 not n19261 ; n19261_not
g79563 not n41482 ; n41482_not
g79564 not n11764 ; n11764_not
g79565 not n12943 ; n12943_not
g79566 not n11755 ; n11755_not
g79567 not n53245 ; n53245_not
g79568 not n41815 ; n41815_not
g79569 not n11746 ; n11746_not
g79570 not n12934 ; n12934_not
g79571 not n45145 ; n45145_not
g79572 not n11737 ; n11737_not
g79573 not n41428 ; n41428_not
g79574 not n11728 ; n11728_not
g79575 not n19270 ; n19270_not
g79576 not n41437 ; n41437_not
g79577 not n12925 ; n12925_not
g79578 not n11719 ; n11719_not
g79579 not n53254 ; n53254_not
g79580 not n41446 ; n41446_not
g79581 not n21925 ; n21925_not
g79582 not n54451 ; n54451_not
g79583 not n21916 ; n21916_not
g79584 not n45127 ; n45127_not
g79585 not n18640 ; n18640_not
g79586 not n42085 ; n42085_not
g79587 not n22096 ; n22096_not
g79588 not n21907 ; n21907_not
g79589 not n43723 ; n43723_not
g79590 not n13276 ; n13276_not
g79591 not n52453 ; n52453_not
g79592 not n53191 ; n53191_not
g79593 not n21880 ; n21880_not
g79594 not n21871 ; n21871_not
g79595 not n54442 ; n54442_not
g79596 not n43372 ; n43372_not
g79597 not n21862 ; n21862_not
g79598 not n42076 ; n42076_not
g79599 not n21853 ; n21853_not
g79600 not n53173 ; n53173_not
g79601 not n56206 ; n56206_not
g79602 not n43354 ; n43354_not
g79603 not n13258 ; n13258_not
g79604 not n18622 ; n18622_not
g79605 not n43363 ; n43363_not
g79606 not n42094 ; n42094_not
g79607 not n18550 ; n18550_not
g79608 not n21970 ; n21970_not
g79609 not n18631 ; n18631_not
g79610 not n21961 ; n21961_not
g79611 not n21952 ; n21952_not
g79612 not n21943 ; n21943_not
g79613 not n53182 ; n53182_not
g79614 not n43615 ; n43615_not
g79615 not n21934 ; n21934_not
g79616 not n13267 ; n13267_not
g79617 not n22087 ; n22087_not
g79618 not n22186 ; n22186_not
g79619 not n21745 ; n21745_not
g79620 not n18703 ; n18703_not
g79621 not n22195 ; n22195_not
g79622 not n21736 ; n21736_not
g79623 not n18505 ; n18505_not
g79624 not n18712 ; n18712_not
g79625 not n21727 ; n21727_not
g79626 not n43381 ; n43381_not
g79627 not n54406 ; n54406_not
g79628 not n18721 ; n18721_not
g79629 not n21718 ; n21718_not
g79630 not n42049 ; n42049_not
g79631 not n21709 ; n21709_not
g79632 not n53209 ; n53209_not
g79633 not n18730 ; n18730_not
g79634 not n21691 ; n21691_not
g79635 not n54370 ; n54370_not
g79636 not n21682 ; n21682_not
g79637 not n21673 ; n21673_not
g79638 not n21664 ; n21664_not
g79639 not n21655 ; n21655_not
g79640 not n21646 ; n21646_not
g79641 not n21844 ; n21844_not
g79642 not n54433 ; n54433_not
g79643 not n21835 ; n21835_not
g79644 not n43606 ; n43606_not
g79645 not n21826 ; n21826_not
g79646 not n21817 ; n21817_not
g79647 not n43732 ; n43732_not
g79648 not n42067 ; n42067_not
g79649 not n21808 ; n21808_not
g79650 not n18523 ; n18523_not
g79651 not n54424 ; n54424_not
g79652 not n18514 ; n18514_not
g79653 not n21790 ; n21790_not
g79654 not n21781 ; n21781_not
g79655 not n21772 ; n21772_not
g79656 not n22177 ; n22177_not
g79657 not n21763 ; n21763_not
g79658 not n21754 ; n21754_not
g79659 not n54415 ; n54415_not
g79660 not n54361 ; n54361_not
g79661 not n42058 ; n42058_not
g79662 not n54505 ; n54505_not
g79663 not n18532 ; n18532_not
g79664 not n42139 ; n42139_not
g79665 not n56215 ; n56215_not
g79666 not n43345 ; n43345_not
g79667 not n43624 ; n43624_not
g79668 not n22906 ; n22906_not
g79669 not n54523 ; n54523_not
g79670 not n43714 ; n43714_not
g79671 not n53146 ; n53146_not
g79672 not n54514 ; n54514_not
g79673 not n42148 ; n42148_not
g79674 not n22951 ; n22951_not
g79675 not n54325 ; n54325_not
g79676 not n11566 ; n11566_not
g79677 not n53164 ; n53164_not
g79678 not n22816 ; n22816_not
g79679 not n54334 ; n54334_not
g79680 not n18604 ; n18604_not
g79681 not n54460 ; n54460_not
g79682 not n52462 ; n52462_not
g79683 not n18613 ; n18613_not
g79684 not n54316 ; n54316_not
g79685 not n53155 ; n53155_not
g79686 not n52471 ; n52471_not
g79687 not n22861 ; n22861_not
g79688 not n44902 ; n44902_not
g79689 not n40735 ; n40735_not
g79690 not n44434 ; n44434_not
g79691 not n52426 ; n52426_not
g79692 not n53236 ; n53236_not
g79693 not n44821 ; n44821_not
g79694 not n18901 ; n18901_not
g79695 not n43417 ; n43417_not
g79696 not n53227 ; n53227_not
g79697 not n13285 ; n13285_not
g79698 not n22069 ; n22069_not
g79699 not n40645 ; n40645_not
g79700 not n53308 ; n53308_not
g79701 not n21448 ; n21448_not
g79702 not n43426 ; n43426_not
g79703 not n53263 ; n53263_not
g79704 not n41950 ; n41950_not
g79705 not n18910 ; n18910_not
g79706 not n21358 ; n21358_not
g79707 not n43435 ; n43435_not
g79708 not n54253 ; n54253_not
g79709 not n13195 ; n13195_not
g79710 not n21556 ; n21556_not
g79711 not n21565 ; n21565_not
g79712 not n21574 ; n21574_not
g79713 not n54343 ; n54343_not
g79714 not n22276 ; n22276_not
g79715 not n21583 ; n21583_not
g79716 not n56071 ; n56071_not
g79717 not n18802 ; n18802_not
g79718 not n21592 ; n21592_not
g79719 not n22267 ; n22267_not
g79720 not n21619 ; n21619_not
g79721 not n21628 ; n21628_not
g79722 not n22249 ; n22249_not
g79723 not n44407 ; n44407_not
g79724 not n21637 ; n21637_not
g79725 not n40690 ; n40690_not
g79726 not n11476 ; n11476_not
g79727 not n43390 ; n43390_not
g79728 not n22285 ; n22285_not
g79729 not n53218 ; n53218_not
g79730 not n22294 ; n22294_not
g79731 not n22159 ; n22159_not
g79732 not n18433 ; n18433_not
g79733 not n18811 ; n18811_not
g79734 not n43408 ; n43408_not
g79735 not n18820 ; n18820_not
g79736 not n56170 ; n56170_not
g79737 not n56431 ; n56431_not
g79738 not n16525 ; n16525_not
g79739 not n45631 ; n45631_not
g79740 not n15247 ; n15247_not
g79741 not n55135 ; n55135_not
g79742 not n55513 ; n55513_not
g79743 not n45721 ; n45721_not
g79744 not n26146 ; n26146_not
g79745 not n44713 ; n44713_not
g79746 not n15535 ; n15535_not
g79747 not n26137 ; n26137_not
g79748 not n14761 ; n14761_not
g79749 not n16516 ; n16516_not
g79750 not n40087 ; n40087_not
g79751 not n16534 ; n16534_not
g79752 not n26119 ; n26119_not
g79753 not n52165 ; n52165_not
g79754 not n57313 ; n57313_not
g79755 not n26182 ; n26182_not
g79756 not n15517 ; n15517_not
g79757 not n45622 ; n45622_not
g79758 not n43075 ; n43075_not
g79759 not n55270 ; n55270_not
g79760 not n52417 ; n52417_not
g79761 not n43282 ; n43282_not
g79762 not n40069 ; n40069_not
g79763 not n56422 ; n56422_not
g79764 not n15184 ; n15184_not
g79765 not n26164 ; n26164_not
g79766 not n15526 ; n15526_not
g79767 not n52156 ; n52156_not
g79768 not n52138 ; n52138_not
g79769 not n25228 ; n25228_not
g79770 not n43066 ; n43066_not
g79771 not n39511 ; n39511_not
g79772 not n15553 ; n15553_not
g79773 not n16480 ; n16480_not
g79774 not n26047 ; n26047_not
g79775 not n26038 ; n26038_not
g79776 not n14743 ; n14743_not
g79777 not n52129 ; n52129_not
g79778 not n26029 ; n26029_not
g79779 not n25246 ; n25246_not
g79780 not n57331 ; n57331_not
g79781 not n15652 ; n15652_not
g79782 not n25255 ; n25255_not
g79783 not n25264 ; n25264_not
g79784 not n52435 ; n52435_not
g79785 not n15175 ; n15175_not
g79786 not n43147 ; n43147_not
g79787 not n55252 ; n55252_not
g79788 not n26092 ; n26092_not
g79789 not n55261 ; n55261_not
g79790 not n52147 ; n52147_not
g79791 not n57322 ; n57322_not
g79792 not n26074 ; n26074_not
g79793 not n26056 ; n26056_not
g79794 not n56440 ; n56440_not
g79795 not n42454 ; n42454_not
g79796 not n15544 ; n15544_not
g79797 not n14752 ; n14752_not
g79798 not n26065 ; n26065_not
g79799 not n15661 ; n15661_not
g79800 not n15256 ; n15256_not
g79801 not n45550 ; n45550_not
g79802 not n26272 ; n26272_not
g79803 not n14626 ; n14626_not
g79804 not n15418 ; n15418_not
g79805 not n44551 ; n44551_not
g79806 not n16390 ; n16390_not
g79807 not n15427 ; n15427_not
g79808 not n55018 ; n55018_not
g79809 not n16417 ; n16417_not
g79810 not n15724 ; n15724_not
g79811 not n44641 ; n44641_not
g79812 not n14455 ; n14455_not
g79813 not n14617 ; n14617_not
g79814 not n15436 ; n15436_not
g79815 not n16435 ; n16435_not
g79816 not n43039 ; n43039_not
g79817 not n26254 ; n26254_not
g79818 not n45604 ; n45604_not
g79819 not n14608 ; n14608_not
g79820 not n14644 ; n14644_not
g79821 not n52192 ; n52192_not
g79822 not n16372 ; n16372_not
g79823 not n45532 ; n45532_not
g79824 not n15382 ; n15382_not
g79825 not n15751 ; n15751_not
g79826 not n14635 ; n14635_not
g79827 not n15391 ; n15391_not
g79828 not n15742 ; n15742_not
g79829 not n45541 ; n45541_not
g79830 not n26911 ; n26911_not
g79831 not n14446 ; n14446_not
g79832 not n15409 ; n15409_not
g79833 not n26281 ; n26281_not
g79834 not n44533 ; n44533_not
g79835 not n15229 ; n15229_not
g79836 not n15481 ; n15481_not
g79837 not n26209 ; n26209_not
g79838 not n52174 ; n52174_not
g79839 not n55405 ; n55405_not
g79840 not n15490 ; n15490_not
g79841 not n14770 ; n14770_not
g79842 not n45613 ; n45613_not
g79843 not n56413 ; n56413_not
g79844 not n15193 ; n15193_not
g79845 not n44650 ; n44650_not
g79846 not n15508 ; n15508_not
g79847 not n26191 ; n26191_not
g79848 not n15238 ; n15238_not
g79849 not n16444 ; n16444_not
g79850 not n15445 ; n15445_not
g79851 not n52183 ; n52183_not
g79852 not n45730 ; n45730_not
g79853 not n15454 ; n15454_not
g79854 not n15463 ; n15463_not
g79855 not n56404 ; n56404_not
g79856 not n26236 ; n26236_not
g79857 not n15706 ; n15706_not
g79858 not n26227 ; n26227_not
g79859 not n52408 ; n52408_not
g79860 not n16462 ; n16462_not
g79861 not n55630 ; n55630_not
g79862 not n39502 ; n39502_not
g79863 not n15472 ; n15472_not
g79864 not n15292 ; n15292_not
g79865 not n42913 ; n42913_not
g79866 not n55423 ; n55423_not
g79867 not n25381 ; n25381_not
g79868 not n52525 ; n52525_not
g79869 not n27109 ; n27109_not
g79870 not n56611 ; n56611_not
g79871 not n14545 ; n14545_not
g79872 not n25390 ; n25390_not
g79873 not n55702 ; n55702_not
g79874 not n42904 ; n42904_not
g79875 not n45037 ; n45037_not
g79876 not n40195 ; n40195_not
g79877 not n44524 ; n44524_not
g79878 not n55414 ; n55414_not
g79879 not n42922 ; n42922_not
g79880 not n15607 ; n15607_not
g79881 not n25822 ; n25822_not
g79882 not n55225 ; n55225_not
g79883 not n25813 ; n25813_not
g79884 not n56602 ; n56602_not
g79885 not n16408 ; n16408_not
g79886 not n25804 ; n25804_not
g79887 not n14536 ; n14536_not
g79888 not n55432 ; n55432_not
g79889 not n40267 ; n40267_not
g79890 not n26515 ; n26515_not
g79891 not n56710 ; n56710_not
g79892 not n25714 ; n25714_not
g79893 not n14572 ; n14572_not
g79894 not n26506 ; n26506_not
g79895 not n56701 ; n56701_not
g79896 not n15562 ; n15562_not
g79897 not n16363 ; n16363_not
g79898 not n25705 ; n25705_not
g79899 not n25426 ; n25426_not
g79900 not n16354 ; n16354_not
g79901 not n15580 ; n15580_not
g79902 not n40249 ; n40249_not
g79903 not n56620 ; n56620_not
g79904 not n25750 ; n25750_not
g79905 not n25741 ; n25741_not
g79906 not n55504 ; n55504_not
g79907 not n25732 ; n25732_not
g79908 not n55207 ; n55207_not
g79909 not n25723 ; n25723_not
g79910 not n15571 ; n15571_not
g79911 not n25291 ; n25291_not
g79912 not n45640 ; n45640_not
g79913 not n14491 ; n14491_not
g79914 not n45703 ; n45703_not
g79915 not n57340 ; n57340_not
g79916 not n14707 ; n14707_not
g79917 not n25930 ; n25930_not
g79918 not n25921 ; n25921_not
g79919 not n16453 ; n16453_not
g79920 not n25309 ; n25309_not
g79921 not n45019 ; n45019_not
g79922 not n27019 ; n27019_not
g79923 not n56800 ; n56800_not
g79924 not n14734 ; n14734_not
g79925 not n56503 ; n56503_not
g79926 not n14482 ; n14482_not
g79927 not n14725 ; n14725_not
g79928 not n45154 ; n45154_not
g79929 not n15265 ; n15265_not
g79930 not n14716 ; n14716_not
g79931 not n40177 ; n40177_not
g79932 not n15283 ; n15283_not
g79933 not n25336 ; n25336_not
g79934 not n14662 ; n14662_not
g79935 not n42931 ; n42931_not
g79936 not n25345 ; n25345_not
g79937 not n14653 ; n14653_not
g79938 not n25840 ; n25840_not
g79939 not n25354 ; n25354_not
g79940 not n55234 ; n55234_not
g79941 not n25831 ; n25831_not
g79942 not n14527 ; n14527_not
g79943 not n15625 ; n15625_not
g79944 not n15274 ; n15274_not
g79945 not n25912 ; n25912_not
g79946 not n25903 ; n25903_not
g79947 not n56512 ; n56512_not
g79948 not n56521 ; n56521_not
g79949 not n27064 ; n27064_not
g79950 not n42940 ; n42940_not
g79951 not n52480 ; n52480_not
g79952 not n14680 ; n14680_not
g79953 not n15634 ; n15634_not
g79954 not n56530 ; n56530_not
g79955 not n14671 ; n14671_not
g79956 not n45334 ; n45334_not
g79957 not n45325 ; n45325_not
g79958 not n55315 ; n55315_not
g79959 not n44605 ; n44605_not
g79960 not n14806 ; n14806_not
g79961 not n26155 ; n26155_not
g79962 not n45316 ; n45316_not
g79963 not n45307 ; n45307_not
g79964 not n16093 ; n16093_not
g79965 not n45901 ; n45901_not
g79966 not n14932 ; n14932_not
g79967 not n15085 ; n15085_not
g79968 not n45910 ; n45910_not
g79969 not n45280 ; n45280_not
g79970 not n52264 ; n52264_not
g79971 not n55360 ; n55360_not
g79972 not n57034 ; n57034_not
g79973 not n14950 ; n14950_not
g79974 not n43174 ; n43174_not
g79975 not n45361 ; n45361_not
g79976 not n14833 ; n14833_not
g79977 not n16075 ; n16075_not
g79978 not n14824 ; n14824_not
g79979 not n42850 ; n42850_not
g79980 not n57142 ; n57142_not
g79981 not n45352 ; n45352_not
g79982 not n14365 ; n14365_not
g79983 not n57025 ; n57025_not
g79984 not n45343 ; n45343_not
g79985 not n14941 ; n14941_not
g79986 not n15904 ; n15904_not
g79987 not n52345 ; n52345_not
g79988 not n16084 ; n16084_not
g79989 not n14815 ; n14815_not
g79990 not n16147 ; n16147_not
g79991 not n52363 ; n52363_not
g79992 not n52255 ; n52255_not
g79993 not n45514 ; n45514_not
g79994 not n14905 ; n14905_not
g79995 not n45271 ; n45271_not
g79996 not n45523 ; n45523_not
g79997 not n55306 ; n55306_not
g79998 not n16156 ; n16156_not
g79999 not n15841 ; n15841_not
g80000 not n26290 ; n26290_not
g80001 not n52354 ; n52354_not
g80002 not n15715 ; n15715_not
g80003 not n45505 ; n45505_not
g80004 not n43156 ; n43156_not
g80005 not n14923 ; n14923_not
g80006 not n55531 ; n55531_not
g80007 not n15832 ; n15832_not
g80008 not n16129 ; n16129_not
g80009 not n16138 ; n16138_not
g80010 not n14914 ; n14914_not
g80011 not n15094 ; n15094_not
g80012 not n55180 ; n55180_not
g80013 not n45460 ; n45460_not
g80014 not n55063 ; n55063_not
g80015 not n45811 ; n45811_not
g80016 not n43219 ; n43219_not
g80017 not n55351 ; n55351_not
g80018 not n55324 ; n55324_not
g80019 not n45424 ; n45424_not
g80020 not n52309 ; n52309_not
g80021 not n52282 ; n52282_not
g80022 not n43264 ; n43264_not
g80023 not n44731 ; n44731_not
g80024 not n15940 ; n15940_not
g80025 not n15760 ; n15760_not
g80026 not n15805 ; n15805_not
g80027 not n45415 ; n45415_not
g80028 not n55540 ; n55540_not
g80029 not n52291 ; n52291_not
g80030 not n42724 ; n42724_not
g80031 not n51706 ; n51706_not
g80032 not n55342 ; n55342_not
g80033 not n43237 ; n43237_not
g80034 not n45451 ; n45451_not
g80035 not n43246 ; n43246_not
g80036 not n42733 ; n42733_not
g80037 not n42742 ; n42742_not
g80038 not n45820 ; n45820_not
g80039 not n44740 ; n44740_not
g80040 not n45442 ; n45442_not
g80041 not n42751 ; n42751_not
g80042 not n57070 ; n57070_not
g80043 not n55333 ; n55333_not
g80044 not n45433 ; n45433_not
g80045 not n42760 ; n42760_not
g80046 not n16048 ; n16048_not
g80047 not n14851 ; n14851_not
g80048 not n57124 ; n57124_not
g80049 not n26245 ; n26245_not
g80050 not n42832 ; n42832_not
g80051 not n52327 ; n52327_not
g80052 not n14842 ; n14842_not
g80053 not n16057 ; n16057_not
g80054 not n57043 ; n57043_not
g80055 not n15913 ; n15913_not
g80056 not n45046 ; n45046_not
g80057 not n16066 ; n16066_not
g80058 not n15067 ; n15067_not
g80059 not n45370 ; n45370_not
g80060 not n42841 ; n42841_not
g80061 not n52336 ; n52336_not
g80062 not n57106 ; n57106_not
g80063 not n15931 ; n15931_not
g80064 not n45109 ; n45109_not
g80065 not n15049 ; n15049_not
g80066 not n45406 ; n45406_not
g80067 not n57115 ; n57115_not
g80068 not n42805 ; n42805_not
g80069 not n14860 ; n14860_not
g80070 not n52273 ; n52273_not
g80071 not n57052 ; n57052_not
g80072 not n43192 ; n43192_not
g80073 not n52318 ; n52318_not
g80074 not n42814 ; n42814_not
g80075 not n16039 ; n16039_not
g80076 not n42823 ; n42823_not
g80077 not n15922 ; n15922_not
g80078 not n43084 ; n43084_not
g80079 not n16264 ; n16264_not
g80080 not n16273 ; n16273_not
g80081 not n16282 ; n16282_not
g80082 not n26344 ; n26344_not
g80083 not n39601 ; n39601_not
g80084 not n39403 ; n39403_not
g80085 not n14437 ; n14437_not
g80086 not n52219 ; n52219_not
g80087 not n16255 ; n16255_not
g80088 not n25534 ; n25534_not
g80089 not n44623 ; n44623_not
g80090 not n15814 ; n15814_not
g80091 not n15139 ; n15139_not
g80092 not n15157 ; n15157_not
g80093 not n26317 ; n26317_not
g80094 not n39430 ; n39430_not
g80095 not n57250 ; n57250_not
g80096 not n15346 ; n15346_not
g80097 not n55522 ; n55522_not
g80098 not n15355 ; n15355_not
g80099 not n15364 ; n15364_not
g80100 not n16345 ; n16345_not
g80101 not n15373 ; n15373_not
g80102 not n39412 ; n39412_not
g80103 not n15319 ; n15319_not
g80104 not n55144 ; n55144_not
g80105 not n51751 ; n51751_not
g80106 not n16309 ; n16309_not
g80107 not n44542 ; n44542_not
g80108 not n57241 ; n57241_not
g80109 not n15328 ; n15328_not
g80110 not n39421 ; n39421_not
g80111 not n15337 ; n15337_not
g80112 not n16327 ; n16327_not
g80113 not n44632 ; n44632_not
g80114 not n55621 ; n55621_not
g80115 not n26326 ; n26326_not
g80116 not n55603 ; n55603_not
g80117 not n15670 ; n15670_not
g80118 not n16183 ; n16183_not
g80119 not n15850 ; n15850_not
g80120 not n26335 ; n26335_not
g80121 not n52381 ; n52381_not
g80122 not n16192 ; n16192_not
g80123 not n44614 ; n44614_not
g80124 not n16165 ; n16165_not
g80125 not n43129 ; n43129_not
g80126 not n51661 ; n51661_not
g80127 not n52372 ; n52372_not
g80128 not n14392 ; n14392_not
g80129 not n43255 ; n43255_not
g80130 not n16174 ; n16174_not
g80131 not n52246 ; n52246_not
g80132 not n16228 ; n16228_not
g80133 not n26362 ; n26362_not
g80134 not n52228 ; n52228_not
g80135 not n16237 ; n16237_not
g80136 not n26371 ; n26371_not
g80137 not n57214 ; n57214_not
g80138 not n44722 ; n44722_not
g80139 not n16246 ; n16246_not
g80140 not n52237 ; n52237_not
g80141 not n16219 ; n16219_not
g80142 not n55612 ; n55612_not
g80143 not n55153 ; n55153_not
g80144 not n52390 ; n52390_not
g80145 not n25165 ; n25165_not
g80146 not n43741 ; n43741_not
g80147 not n45064 ; n45064_not
g80148 not n26461 ; n26461_not
g80149 not n25516 ; n25516_not
g80150 not n25174 ; n25174_not
g80151 not n40357 ; n40357_not
g80152 not n52057 ; n52057_not
g80153 not n25543 ; n25543_not
g80154 not n25552 ; n25552_not
g80155 not n40348 ; n40348_not
g80156 not n26443 ; n26443_not
g80157 not n14464 ; n14464_not
g80158 not n43165 ; n43165_not
g80159 not n16570 ; n16570_not
g80160 not n25570 ; n25570_not
g80161 not n17173 ; n17173_not
g80162 not n17056 ; n17056_not
g80163 not n26416 ; n26416_not
g80164 not n52084 ; n52084_not
g80165 not n26425 ; n26425_not
g80166 not n16561 ; n16561_not
g80167 not n25408 ; n25408_not
g80168 not n25147 ; n25147_not
g80169 not n40339 ; n40339_not
g80170 not n25561 ; n25561_not
g80171 not n25156 ; n25156_not
g80172 not n55162 ; n55162_not
g80173 not n42544 ; n42544_not
g80174 not n25435 ; n25435_not
g80175 not n55720 ; n55720_not
g80176 not n26407 ; n26407_not
g80177 not n14554 ; n14554_not
g80178 not n14419 ; n14419_not
g80179 not n57412 ; n57412_not
g80180 not n44416 ; n44416_not
g80181 not n40375 ; n40375_not
g80182 not n26470 ; n26470_not
g80183 not n17146 ; n17146_not
g80184 not n14509 ; n14509_not
g80185 not n25480 ; n25480_not
g80186 not n25471 ; n25471_not
g80187 not n52660 ; n52660_not
g80188 not n52615 ; n52615_not
g80189 not n27172 ; n27172_not
g80190 not n40366 ; n40366_not
g80191 not n25273 ; n25273_not
g80192 not n55117 ; n55117_not
g80193 not n27226 ; n27226_not
g80194 not n25453 ; n25453_not
g80195 not n44704 ; n44704_not
g80196 not n55090 ; n55090_not
g80197 not n15058 ; n15058_not
g80198 not n25183 ; n25183_not
g80199 not n44461 ; n44461_not
g80200 not n40384 ; n40384_not
g80201 not n52075 ; n52075_not
g80202 not n57430 ; n57430_not
g80203 not n55108 ; n55108_not
g80204 not n25192 ; n25192_not
g80205 not n25525 ; n25525_not
g80206 not n26434 ; n26434_not
g80207 not n57403 ; n57403_not
g80208 not n14374 ; n14374_not
g80209 not n40294 ; n40294_not
g80210 not n26452 ; n26452_not
g80211 not n52066 ; n52066_not
g80212 not n40258 ; n40258_not
g80213 not n25651 ; n25651_not
g80214 not n17191 ; n17191_not
g80215 not n55072 ; n55072_not
g80216 not n25093 ; n25093_not
g80217 not n25660 ; n25660_not
g80218 not n16552 ; n16552_not
g80219 not n27181 ; n27181_not
g80220 not n15148 ; n15148_not
g80221 not n25075 ; n25075_not
g80222 not n17218 ; n17218_not
g80223 not n52093 ; n52093_not
g80224 not n40285 ; n40285_not
g80225 not n27154 ; n27154_not
g80226 not n55711 ; n55711_not
g80227 not n25066 ; n25066_not
g80228 not n44452 ; n44452_not
g80229 not n25363 ; n25363_not
g80230 not n57502 ; n57502_not
g80231 not n17182 ; n17182_not
g80232 not n25084 ; n25084_not
g80233 not n17209 ; n17209_not
g80234 not n25444 ; n25444_not
g80235 not n40438 ; n40438_not
g80236 not n55801 ; n55801_not
g80237 not n10099 ; n10099_not
g80238 not n25318 ; n25318_not
g80239 not n25129 ; n25129_not
g80240 not n44506 ; n44506_not
g80241 not n25606 ; n25606_not
g80242 not n16318 ; n16318_not
g80243 not n25615 ; n25615_not
g80244 not n40429 ; n40429_not
g80245 not n24454 ; n24454_not
g80246 not n55450 ; n55450_not
g80247 not n27190 ; n27190_not
g80248 not n25138 ; n25138_not
g80249 not n40393 ; n40393_not
g80250 not n39043 ; n39043_not
g80251 not n55441 ; n55441_not
g80252 not n25633 ; n25633_not
g80253 not n52570 ; n52570_not
g80254 not n25624 ; n25624_not
g80255 not n45055 ; n45055_not
g80256 not n25642 ; n25642_not
g80257 not n43283 ; n43283_not
g80258 not n12980 ; n12980_not
g80259 not n12755 ; n12755_not
g80260 not n14816 ; n14816_not
g80261 not n15851 ; n15851_not
g80262 not n54245 ; n54245_not
g80263 not n30836 ; n30836_not
g80264 not n34517 ; n34517_not
g80265 not n37226 ; n37226_not
g80266 not n32780 ; n32780_not
g80267 not n43823 ; n43823_not
g80268 not n12773 ; n12773_not
g80269 not n34391 ; n34391_not
g80270 not n18380 ; n18380_not
g80271 not n53804 ; n53804_not
g80272 not n43922 ; n43922_not
g80273 not n14825 ; n14825_not
g80274 not n12764 ; n12764_not
g80275 not n12944 ; n12944_not
g80276 not n30854 ; n30854_not
g80277 not n53903 ; n53903_not
g80278 not n32762 ; n32762_not
g80279 not n37262 ; n37262_not
g80280 not n41672 ; n41672_not
g80281 not n53552 ; n53552_not
g80282 not n14753 ; n14753_not
g80283 not n30863 ; n30863_not
g80284 not n15095 ; n15095_not
g80285 not n55406 ; n55406_not
g80286 not n41438 ; n41438_not
g80287 not n41933 ; n41933_not
g80288 not n13097 ; n13097_not
g80289 not n32753 ; n32753_not
g80290 not n31259 ; n31259_not
g80291 not n15437 ; n15437_not
g80292 not n32735 ; n32735_not
g80293 not n18911 ; n18911_not
g80294 not n30647 ; n30647_not
g80295 not n19136 ; n19136_not
g80296 not n53750 ; n53750_not
g80297 not n15842 ; n15842_not
g80298 not n33284 ; n33284_not
g80299 not n34445 ; n34445_not
g80300 not n37235 ; n37235_not
g80301 not n33329 ; n33329_not
g80302 not n13187 ; n13187_not
g80303 not n18920 ; n18920_not
g80304 not n56063 ; n56063_not
g80305 not n30665 ; n30665_not
g80306 not n19622 ; n19622_not
g80307 not n12962 ; n12962_not
g80308 not n12971 ; n12971_not
g80309 not n41681 ; n41681_not
g80310 not n44066 ; n44066_not
g80311 not n19118 ; n19118_not
g80312 not n19127 ; n19127_not
g80313 not n37244 ; n37244_not
g80314 not n32771 ; n32771_not
g80315 not n13079 ; n13079_not
g80316 not n31268 ; n31268_not
g80317 not n44138 ; n44138_not
g80318 not n12953 ; n12953_not
g80319 not n41942 ; n41942_not
g80320 not n13178 ; n13178_not
g80321 not n54263 ; n54263_not
g80322 not n13088 ; n13088_not
g80323 not n38126 ; n38126_not
g80324 not n33464 ; n33464_not
g80325 not n30845 ; n30845_not
g80326 not n43445 ; n43445_not
g80327 not n37253 ; n37253_not
g80328 not n30656 ; n30656_not
g80329 not n19613 ; n19613_not
g80330 not n43517 ; n43517_not
g80331 not n19604 ; n19604_not
g80332 not n54236 ; n54236_not
g80333 not n53813 ; n53813_not
g80334 not n19631 ; n19631_not
g80335 not n53336 ; n53336_not
g80336 not n44408 ; n44408_not
g80337 not n33338 ; n33338_not
g80338 not n32744 ; n32744_not
g80339 not n15383 ; n15383_not
g80340 not n18434 ; n18434_not
g80341 not n12674 ; n12674_not
g80342 not n14771 ; n14771_not
g80343 not n15815 ; n15815_not
g80344 not n53642 ; n53642_not
g80345 not n30593 ; n30593_not
g80346 not n19073 ; n19073_not
g80347 not n15275 ; n15275_not
g80348 not n15059 ; n15059_not
g80349 not n12854 ; n12854_not
g80350 not n42671 ; n42671_not
g80351 not n32906 ; n32906_not
g80352 not n19703 ; n19703_not
g80353 not n44048 ; n44048_not
g80354 not n37613 ; n37613_not
g80355 not n32933 ; n32933_not
g80356 not n37154 ; n37154_not
g80357 not n18830 ; n18830_not
g80358 not n15923 ; n15923_not
g80359 not n55532 ; n55532_not
g80360 not n43274 ; n43274_not
g80361 not n43526 ; n43526_not
g80362 not n30782 ; n30782_not
g80363 not n30746 ; n30746_not
g80364 not n12872 ; n12872_not
g80365 not n43175 ; n43175_not
g80366 not n32870 ; n32870_not
g80367 not n13295 ; n13295_not
g80368 not n33491 ; n33491_not
g80369 not n37172 ; n37172_not
g80370 not n32951 ; n32951_not
g80371 not n12863 ; n12863_not
g80372 not n44147 ; n44147_not
g80373 not n53840 ; n53840_not
g80374 not n49340 ; n49340_not
g80375 not n37604 ; n37604_not
g80376 not n45191 ; n45191_not
g80377 not n37163 ; n37163_not
g80378 not n49241 ; n49241_not
g80379 not n30791 ; n30791_not
g80380 not n15266 ; n15266_not
g80381 not n42662 ; n42662_not
g80382 not n53651 ; n53651_not
g80383 not n43427 ; n43427_not
g80384 not n12683 ; n12683_not
g80385 not n15914 ; n15914_not
g80386 not n38144 ; n38144_not
g80387 not n12809 ; n12809_not
g80388 not n37622 ; n37622_not
g80389 not n54335 ; n54335_not
g80390 not n18812 ; n18812_not
g80391 not n43256 ; n43256_not
g80392 not n32708 ; n32708_not
g80393 not n44840 ; n44840_not
g80394 not n53624 ; n53624_not
g80395 not n12791 ; n12791_not
g80396 not n30773 ; n30773_not
g80397 not n19721 ; n19721_not
g80398 not n15950 ; n15950_not
g80399 not n43247 ; n43247_not
g80400 not n18803 ; n18803_not
g80401 not n19730 ; n19730_not
g80402 not n30575 ; n30575_not
g80403 not n55343 ; n55343_not
g80404 not n50276 ; n50276_not
g80405 not n43418 ; n43418_not
g80406 not n12656 ; n12656_not
g80407 not n30557 ; n30557_not
g80408 not n54326 ; n54326_not
g80409 not n18443 ; n18443_not
g80410 not n14780 ; n14780_not
g80411 not n41069 ; n41069_not
g80412 not n15806 ; n15806_not
g80413 not n15392 ; n15392_not
g80414 not n12845 ; n12845_not
g80415 not n53633 ; n53633_not
g80416 not n15284 ; n15284_not
g80417 not n18821 ; n18821_not
g80418 not n55064 ; n55064_not
g80419 not n15932 ; n15932_not
g80420 not n19712 ; n19712_not
g80421 not n30584 ; n30584_not
g80422 not n41636 ; n41636_not
g80423 not n45335 ; n45335_not
g80424 not n15293 ; n15293_not
g80425 not n55541 ; n55541_not
g80426 not n12836 ; n12836_not
g80427 not n43166 ; n43166_not
g80428 not n49232 ; n49232_not
g80429 not n33509 ; n33509_not
g80430 not n12827 ; n12827_not
g80431 not n15941 ; n15941_not
g80432 not n12818 ; n12818_not
g80433 not n55352 ; n55352_not
g80434 not n12917 ; n12917_not
g80435 not n14762 ; n14762_not
g80436 not n53723 ; n53723_not
g80437 not n55370 ; n55370_not
g80438 not n13268 ; n13268_not
g80439 not n14807 ; n14807_not
g80440 not n43265 ; n43265_not
g80441 not n12908 ; n12908_not
g80442 not n32807 ; n32807_not
g80443 not n30629 ; n30629_not
g80444 not n15419 ; n15419_not
g80445 not n54281 ; n54281_not
g80446 not n37217 ; n37217_not
g80447 not n41960 ; n41960_not
g80448 not n53354 ; n53354_not
g80449 not n15239 ; n15239_not
g80450 not n13277 ; n13277_not
g80451 not n31286 ; n31286_not
g80452 not n12746 ; n12746_not
g80453 not n53714 ; n53714_not
g80454 not n34436 ; n34436_not
g80455 not n37208 ; n37208_not
g80456 not n15428 ; n15428_not
g80457 not n12935 ; n12935_not
g80458 not n30638 ; n30638_not
g80459 not n19640 ; n19640_not
g80460 not n53741 ; n53741_not
g80461 not n41096 ; n41096_not
g80462 not n33473 ; n33473_not
g80463 not n41663 ; n41663_not
g80464 not n43832 ; n43832_not
g80465 not n53345 ; n53345_not
g80466 not n18902 ; n18902_not
g80467 not n47801 ; n47801_not
g80468 not n30827 ; n30827_not
g80469 not n12926 ; n12926_not
g80470 not n31277 ; n31277_not
g80471 not n53732 ; n53732_not
g80472 not n55154 ; n55154_not
g80473 not n55073 ; n55073_not
g80474 not n15374 ; n15374_not
g80475 not n43436 ; n43436_not
g80476 not n49250 ; n49250_not
g80477 not n30728 ; n30728_not
g80478 not n32843 ; n32843_not
g80479 not n55361 ; n55361_not
g80480 not n54308 ; n54308_not
g80481 not n30737 ; n30737_not
g80482 not n12881 ; n12881_not
g80483 not n41078 ; n41078_not
g80484 not n41645 ; n41645_not
g80485 not n32852 ; n32852_not
g80486 not n19082 ; n19082_not
g80487 not n34373 ; n34373_not
g80488 not n37190 ; n37190_not
g80489 not n15077 ; n15077_not
g80490 not n15257 ; n15257_not
g80491 not n37451 ; n37451_not
g80492 not n18425 ; n18425_not
g80493 not n38135 ; n38135_not
g80494 not n32861 ; n32861_not
g80495 not n37181 ; n37181_not
g80496 not n53660 ; n53660_not
g80497 not n15905 ; n15905_not
g80498 not n32816 ; n32816_not
g80499 not n54290 ; n54290_not
g80500 not n55163 ; n55163_not
g80501 not n30818 ; n30818_not
g80502 not n53705 ; n53705_not
g80503 not n45092 ; n45092_not
g80504 not n37406 ; n37406_not
g80505 not n41087 ; n41087_not
g80506 not n41654 ; n41654_not
g80507 not n32825 ; n32825_not
g80508 not n12890 ; n12890_not
g80509 not n45344 ; n45344_not
g80510 not n44057 ; n44057_not
g80511 not n32834 ; n32834_not
g80512 not n33482 ; n33482_not
g80513 not n31295 ; n31295_not
g80514 not n12728 ; n12728_not
g80515 not n15248 ; n15248_not
g80516 not n19091 ; n19091_not
g80517 not n30809 ; n30809_not
g80518 not n12719 ; n12719_not
g80519 not n41852 ; n41852_not
g80520 not n54038 ; n54038_not
g80521 not n19271 ; n19271_not
g80522 not n19352 ; n19352_not
g80523 not n12629 ; n12629_not
g80524 not n14654 ; n14654_not
g80525 not n37343 ; n37343_not
g80526 not n56045 ; n56045_not
g80527 not n19262 ; n19262_not
g80528 not n56027 ; n56027_not
g80529 not n19172 ; n19172_not
g80530 not n19361 ; n19361_not
g80531 not n43814 ; n43814_not
g80532 not n38045 ; n38045_not
g80533 not n41780 ; n41780_not
g80534 not n43463 ; n43463_not
g80535 not n19163 ; n19163_not
g80536 not n44084 ; n44084_not
g80537 not n19370 ; n19370_not
g80538 not n38036 ; n38036_not
g80539 not n19334 ; n19334_not
g80540 not n14663 ; n14663_not
g80541 not n37352 ; n37352_not
g80542 not n33059 ; n33059_not
g80543 not n54056 ; n54056_not
g80544 not n41843 ; n41843_not
g80545 not n53264 ; n53264_not
g80546 not n19190 ; n19190_not
g80547 not n15329 ; n15329_not
g80548 not n55118 ; n55118_not
g80549 not n47342 ; n47342_not
g80550 not n37433 ; n37433_not
g80551 not n43490 ; n43490_not
g80552 not n15491 ; n15491_not
g80553 not n19343 ; n19343_not
g80554 not n45056 ; n45056_not
g80555 not n45371 ; n45371_not
g80556 not n15644 ; n15644_not
g80557 not n54047 ; n54047_not
g80558 not n37334 ; n37334_not
g80559 not n30917 ; n30917_not
g80560 not n14645 ; n14645_not
g80561 not n41762 ; n41762_not
g80562 not n55451 ; n55451_not
g80563 not n54128 ; n54128_not
g80564 not n19415 ; n19415_not
g80565 not n14636 ; n14636_not
g80566 not n19424 ; n19424_not
g80567 not n30566 ; n30566_not
g80568 not n19226 ; n19226_not
g80569 not n19433 ; n19433_not
g80570 not n30908 ; n30908_not
g80571 not n41186 ; n41186_not
g80572 not n54029 ; n54029_not
g80573 not n14717 ; n14717_not
g80574 not n56018 ; n56018_not
g80575 not n19253 ; n19253_not
g80576 not n38018 ; n38018_not
g80577 not n34490 ; n34490_not
g80578 not n33383 ; n33383_not
g80579 not n41771 ; n41771_not
g80580 not n37424 ; n37424_not
g80581 not n34463 ; n34463_not
g80582 not n14870 ; n14870_not
g80583 not n19145 ; n19145_not
g80584 not n33392 ; n33392_not
g80585 not n15482 ; n15482_not
g80586 not n12692 ; n12692_not
g80587 not n41195 ; n41195_not
g80588 not n19406 ; n19406_not
g80589 not n15338 ; n15338_not
g80590 not n55334 ; n55334_not
g80591 not n41816 ; n41816_not
g80592 not n14924 ; n14924_not
g80593 not n15572 ; n15572_not
g80594 not n14960 ; n14960_not
g80595 not n15536 ; n15536_not
g80596 not n33365 ; n33365_not
g80597 not n15158 ; n15158_not
g80598 not n14681 ; n14681_not
g80599 not n30953 ; n30953_not
g80600 not n14708 ; n14708_not
g80601 not n43157 ; n43157_not
g80602 not n14915 ; n14915_not
g80603 not n44417 ; n44417_not
g80604 not n54065 ; n54065_not
g80605 not n33374 ; n33374_not
g80606 not n43481 ; n43481_not
g80607 not n54083 ; n54083_not
g80608 not n43472 ; n43472_not
g80609 not n15581 ; n15581_not
g80610 not n14942 ; n14942_not
g80611 not n15554 ; n15554_not
g80612 not n55433 ; n55433_not
g80613 not n41825 ; n41825_not
g80614 not n15149 ; n15149_not
g80615 not n14690 ; n14690_not
g80616 not n45362 ; n45362_not
g80617 not n19235 ; n19235_not
g80618 not n15563 ; n15563_not
g80619 not n41807 ; n41807_not
g80620 not n54074 ; n54074_not
g80621 not n30944 ; n30944_not
g80622 not n34508 ; n34508_not
g80623 not n49313 ; n49313_not
g80624 not n14951 ; n14951_not
g80625 not n14933 ; n14933_not
g80626 not n15545 ; n15545_not
g80627 not n12647 ; n12647_not
g80628 not n53255 ; n53255_not
g80629 not n37415 ; n37415_not
g80630 not n15626 ; n15626_not
g80631 not n55505 ; n55505_not
g80632 not n19316 ; n19316_not
g80633 not n37361 ; n37361_not
g80634 not n15608 ; n15608_not
g80635 not n14672 ; n14672_not
g80636 not n15509 ; n15509_not
g80637 not n19325 ; n19325_not
g80638 not n55442 ; n55442_not
g80639 not n34481 ; n34481_not
g80640 not n19217 ; n19217_not
g80641 not n19280 ; n19280_not
g80642 not n30962 ; n30962_not
g80643 not n55424 ; n55424_not
g80644 not n15590 ; n15590_not
g80645 not n32942 ; n32942_not
g80646 not n15527 ; n15527_not
g80647 not n14906 ; n14906_not
g80648 not n15518 ; n15518_not
g80649 not n45074 ; n45074_not
g80650 not n37442 ; n37442_not
g80651 not n12638 ; n12638_not
g80652 not n44093 ; n44093_not
g80653 not n18605 ; n18605_not
g80654 not n19208 ; n19208_not
g80655 not n47333 ; n47333_not
g80656 not n37370 ; n37370_not
g80657 not n55415 ; n55415_not
g80658 not n19307 ; n19307_not
g80659 not n37541 ; n37541_not
g80660 not n19019 ; n19019_not
g80661 not n15167 ; n15167_not
g80662 not n33437 ; n33437_not
g80663 not n19532 ; n19532_not
g80664 not n18335 ; n18335_not
g80665 not n15356 ; n15356_not
g80666 not n14744 ; n14744_not
g80667 not n19541 ; n19541_not
g80668 not n41708 ; n41708_not
g80669 not n37280 ; n37280_not
g80670 not n43508 ; n43508_not
g80671 not n33446 ; n33446_not
g80672 not n33275 ; n33275_not
g80673 not n43454 ; n43454_not
g80674 not n55145 ; n55145_not
g80675 not n49304 ; n49304_not
g80676 not n53912 ; n53912_not
g80677 not n30926 ; n30926_not
g80678 not n44129 ; n44129_not
g80679 not n18317 ; n18317_not
g80680 not n37307 ; n37307_not
g80681 not n19028 ; n19028_not
g80682 not n33257 ; n33257_not
g80683 not n15734 ; n15734_not
g80684 not n41276 ; n41276_not
g80685 not n15455 ; n15455_not
g80686 not n19181 ; n19181_not
g80687 not n19514 ; n19514_not
g80688 not n41717 ; n41717_not
g80689 not n45380 ; n45380_not
g80690 not n33428 ; n33428_not
g80691 not n31196 ; n31196_not
g80692 not n15752 ; n15752_not
g80693 not n19523 ; n19523_not
g80694 not n15761 ; n15761_not
g80695 not n55307 ; n55307_not
g80696 not n53921 ; n53921_not
g80697 not n37109 ; n37109_not
g80698 not n44075 ; n44075_not
g80699 not n33455 ; n33455_not
g80700 not n41690 ; n41690_not
g80701 not n12557 ; n12557_not
g80702 not n34454 ; n34454_not
g80703 not n34418 ; n34418_not
g80704 not n15824 ; n15824_not
g80705 not n54218 ; n54218_not
g80706 not n53831 ; n53831_not
g80707 not n41915 ; n41915_not
g80708 not n30872 ; n30872_not
g80709 not n15365 ; n15365_not
g80710 not n32717 ; n32717_not
g80711 not n53822 ; n53822_not
g80712 not n30674 ; n30674_not
g80713 not n19550 ; n19550_not
g80714 not n14834 ; n14834_not
g80715 not n15446 ; n15446_not
g80716 not n18344 ; n18344_not
g80717 not n38108 ; n38108_not
g80718 not n55316 ; n55316_not
g80719 not n12737 ; n12737_not
g80720 not n30890 ; n30890_not
g80721 not n53930 ; n53930_not
g80722 not n55523 ; n55523_not
g80723 not n37271 ; n37271_not
g80724 not n30692 ; n30692_not
g80725 not n18353 ; n18353_not
g80726 not n54191 ; n54191_not
g80727 not n55460 ; n55460_not
g80728 not n47270 ; n47270_not
g80729 not n30881 ; n30881_not
g80730 not n15671 ; n15671_not
g80731 not n15473 ; n15473_not
g80732 not n15185 ; n15185_not
g80733 not n14627 ; n14627_not
g80734 not n19460 ; n19460_not
g80735 not n41177 ; n41177_not
g80736 not n41744 ; n41744_not
g80737 not n55109 ; n55109_not
g80738 not n45353 ; n45353_not
g80739 not n41168 ; n41168_not
g80740 not n33347 ; n33347_not
g80741 not n41870 ; n41870_not
g80742 not n41753 ; n41753_not
g80743 not n38063 ; n38063_not
g80744 not n15662 ; n15662_not
g80745 not n45182 ; n45182_not
g80746 not n54146 ; n54146_not
g80747 not n14726 ; n14726_not
g80748 not n54155 ; n54155_not
g80749 not n19442 ; n19442_not
g80750 not n47315 ; n47315_not
g80751 not n12593 ; n12593_not
g80752 not n55325 ; n55325_not
g80753 not n37514 ; n37514_not
g80754 not n41258 ; n41258_not
g80755 not n37325 ; n37325_not
g80756 not n19451 ; n19451_not
g80757 not n30971 ; n30971_not
g80758 not n14861 ; n14861_not
g80759 not n37316 ; n37316_not
g80760 not n15707 ; n15707_not
g80761 not n15068 ; n15068_not
g80762 not n14609 ; n14609_not
g80763 not n19037 ; n19037_not
g80764 not n41159 ; n41159_not
g80765 not n41726 ; n41726_not
g80766 not n15716 ; n15716_not
g80767 not n33266 ; n33266_not
g80768 not n15194 ; n15194_not
g80769 not n33419 ; n33419_not
g80770 not n38090 ; n38090_not
g80771 not n14735 ; n14735_not
g80772 not n53309 ; n53309_not
g80773 not n14843 ; n14843_not
g80774 not n19505 ; n19505_not
g80775 not n53291 ; n53291_not
g80776 not n31169 ; n31169_not
g80777 not n15347 ; n15347_not
g80778 not n41735 ; n41735_not
g80779 not n12584 ; n12584_not
g80780 not n14618 ; n14618_not
g80781 not n37523 ; n37523_not
g80782 not n19055 ; n19055_not
g80783 not n55514 ; n55514_not
g80784 not n31178 ; n31178_not
g80785 not n14852 ; n14852_not
g80786 not n54173 ; n54173_not
g80787 not n15464 ; n15464_not
g80788 not n41267 ; n41267_not
g80789 not n38081 ; n38081_not
g80790 not n19046 ; n19046_not
g80791 not n17192 ; n17192_not
g80792 not n43607 ; n43607_not
g80793 not n44354 ; n44354_not
g80794 not n42419 ; n42419_not
g80795 not n43391 ; n43391_not
g80796 not n13970 ; n13970_not
g80797 not n54803 ; n54803_not
g80798 not n33905 ; n33905_not
g80799 not n13961 ; n13961_not
g80800 not n43382 ; n43382_not
g80801 not n43616 ; n43616_not
g80802 not n31880 ; n31880_not
g80803 not n43724 ; n43724_not
g80804 not n16319 ; n16319_not
g80805 not n33752 ; n33752_not
g80806 not n48053 ; n48053_not
g80807 not n55172 ; n55172_not
g80808 not n31907 ; n31907_not
g80809 not n33932 ; n33932_not
g80810 not n42428 ; n42428_not
g80811 not n31718 ; n31718_not
g80812 not n17840 ; n17840_not
g80813 not n33923 ; n33923_not
g80814 not n42536 ; n42536_not
g80815 not n31727 ; n31727_not
g80816 not n54812 ; n54812_not
g80817 not n43733 ; n43733_not
g80818 not n37064 ; n37064_not
g80819 not n42653 ; n42653_not
g80820 not n55730 ; n55730_not
g80821 not n33914 ; n33914_not
g80822 not n31862 ; n31862_not
g80823 not n16328 ; n16328_not
g80824 not n43364 ; n43364_not
g80825 not n48026 ; n48026_not
g80826 not n47243 ; n47243_not
g80827 not n45272 ; n45272_not
g80828 not n34067 ; n34067_not
g80829 not n33860 ; n33860_not
g80830 not n17921 ; n17921_not
g80831 not n48062 ; n48062_not
g80832 not n31853 ; n31853_not
g80833 not n33851 ; n33851_not
g80834 not n55712 ; n55712_not
g80835 not n43355 ; n43355_not
g80836 not n42392 ; n42392_not
g80837 not n43373 ; n43373_not
g80838 not n54164 ; n54164_not
g80839 not n17903 ; n17903_not
g80840 not n50087 ; n50087_not
g80841 not n31871 ; n31871_not
g80842 not n47153 ; n47153_not
g80843 not n55721 ; n55721_not
g80844 not n17912 ; n17912_not
g80845 not n50186 ; n50186_not
g80846 not n13952 ; n13952_not
g80847 not n34058 ; n34058_not
g80848 not n42473 ; n42473_not
g80849 not n16283 ; n16283_not
g80850 not n37811 ; n37811_not
g80851 not n31952 ; n31952_not
g80852 not n14069 ; n14069_not
g80853 not n31943 ; n31943_not
g80854 not n54830 ; n54830_not
g80855 not n37820 ; n37820_not
g80856 not n14096 ; n14096_not
g80857 not n31682 ; n31682_not
g80858 not n37532 ; n37532_not
g80859 not n33725 ; n33725_not
g80860 not n13871 ; n13871_not
g80861 not n37802 ; n37802_not
g80862 not n14087 ; n14087_not
g80863 not n31961 ; n31961_not
g80864 not n13880 ; n13880_not
g80865 not n17750 ; n17750_not
g80866 not n14078 ; n14078_not
g80867 not n14546 ; n14546_not
g80868 not n31925 ; n31925_not
g80869 not n50285 ; n50285_not
g80870 not n31709 ; n31709_not
g80871 not n48044 ; n48044_not
g80872 not n43409 ; n43409_not
g80873 not n43841 ; n43841_not
g80874 not n33950 ; n33950_not
g80875 not n31916 ; n31916_not
g80876 not n37055 ; n37055_not
g80877 not n17822 ; n17822_not
g80878 not n55820 ; n55820_not
g80879 not n33941 ; n33941_not
g80880 not n33770 ; n33770_not
g80881 not n55802 ; n55802_not
g80882 not n45209 ; n45209_not
g80883 not n13907 ; n13907_not
g80884 not n31934 ; n31934_not
g80885 not n42455 ; n42455_not
g80886 not n37721 ; n37721_not
g80887 not n54821 ; n54821_not
g80888 not n17804 ; n17804_not
g80889 not n13916 ; n13916_not
g80890 not n42446 ; n42446_not
g80891 not n13925 ; n13925_not
g80892 not n17813 ; n17813_not
g80893 not n54704 ; n54704_not
g80894 not n55217 ; n55217_not
g80895 not n43661 ; n43661_not
g80896 not n33716 ; n33716_not
g80897 not n14537 ; n14537_not
g80898 not n16409 ; n16409_not
g80899 not n42347 ; n42347_not
g80900 not n42491 ; n42491_not
g80901 not n54209 ; n54209_not
g80902 not n16418 ; n16418_not
g80903 not n50168 ; n50168_not
g80904 not n55703 ; n55703_not
g80905 not n14555 ; n14555_not
g80906 not n43706 ; n43706_not
g80907 not n43328 ; n43328_not
g80908 not n43652 ; n43652_not
g80909 not n37910 ; n37910_not
g80910 not n43319 ; n43319_not
g80911 not n42356 ; n42356_not
g80912 not n54713 ; n54713_not
g80913 not n13862 ; n13862_not
g80914 not n18038 ; n18038_not
g80915 not n31754 ; n31754_not
g80916 not n13826 ; n13826_not
g80917 not n42329 ; n42329_not
g80918 not n45164 ; n45164_not
g80919 not n18047 ; n18047_not
g80920 not n13817 ; n13817_not
g80921 not n41861 ; n41861_not
g80922 not n13844 ; n13844_not
g80923 not n44363 ; n44363_not
g80924 not n33707 ; n33707_not
g80925 not n42338 ; n42338_not
g80926 not n43670 ; n43670_not
g80927 not n31763 ; n31763_not
g80928 not n18029 ; n18029_not
g80929 not n55235 ; n55235_not
g80930 not n31835 ; n31835_not
g80931 not n42383 ; n42383_not
g80932 not n33824 ; n33824_not
g80933 not n33743 ; n33743_not
g80934 not n50177 ; n50177_not
g80935 not n37712 ; n37712_not
g80936 not n47261 ; n47261_not
g80937 not n45227 ; n45227_not
g80938 not n55190 ; n55190_not
g80939 not n31826 ; n31826_not
g80940 not n13934 ; n13934_not
g80941 not n33842 ; n33842_not
g80942 not n43625 ; n43625_not
g80943 not n31844 ; n31844_not
g80944 not n17930 ; n17930_not
g80945 not n32348 ; n32348_not
g80946 not n14573 ; n14573_not
g80947 not n33833 ; n33833_not
g80948 not n43634 ; n43634_not
g80949 not n32339 ; n32339_not
g80950 not n47252 ; n47252_not
g80951 not n34085 ; n34085_not
g80952 not n50078 ; n50078_not
g80953 not n16364 ; n16364_not
g80954 not n37901 ; n37901_not
g80955 not n43346 ; n43346_not
g80956 not n31808 ; n31808_not
g80957 not n43337 ; n43337_not
g80958 not n42365 ; n42365_not
g80959 not n43643 ; n43643_not
g80960 not n33734 ; n33734_not
g80961 not n16373 ; n16373_not
g80962 not n54722 ; n54722_not
g80963 not n42509 ; n42509_not
g80964 not n33815 ; n33815_not
g80965 not n54740 ; n54740_not
g80966 not n16355 ; n16355_not
g80967 not n33806 ; n33806_not
g80968 not n31817 ; n31817_not
g80969 not n42374 ; n42374_not
g80970 not n31772 ; n31772_not
g80971 not n54731 ; n54731_not
g80972 not n45245 ; n45245_not
g80973 not n14258 ; n14258_not
g80974 not n32285 ; n32285_not
g80975 not n42626 ; n42626_not
g80976 not n43544 ; n43544_not
g80977 not n32258 ; n32258_not
g80978 not n32087 ; n32087_not
g80979 not n14276 ; n14276_not
g80980 not n17138 ; n17138_not
g80981 not n45254 ; n45254_not
g80982 not n13772 ; n13772_not
g80983 not n32294 ; n32294_not
g80984 not n32159 ; n32159_not
g80985 not n32276 ; n32276_not
g80986 not n17093 ; n17093_not
g80987 not n17156 ; n17156_not
g80988 not n55082 ; n55082_not
g80989 not n55019 ; n55019_not
g80990 not n44327 ; n44327_not
g80991 not n14285 ; n14285_not
g80992 not n47162 ; n47162_not
g80993 not n17084 ; n17084_not
g80994 not n32267 ; n32267_not
g80995 not n14429 ; n14429_not
g80996 not n42581 ; n42581_not
g80997 not n14195 ; n14195_not
g80998 not n14186 ; n14186_not
g80999 not n43553 ; n43553_not
g81000 not n17039 ; n17039_not
g81001 not n32096 ; n32096_not
g81002 not n42635 ; n42635_not
g81003 not n50195 ; n50195_not
g81004 not n32249 ; n32249_not
g81005 not n14267 ; n14267_not
g81006 not n17129 ; n17129_not
g81007 not n14249 ; n14249_not
g81008 not n33662 ; n33662_not
g81009 not n17057 ; n17057_not
g81010 not n45236 ; n45236_not
g81011 not n32069 ; n32069_not
g81012 not n17048 ; n17048_not
g81013 not n17147 ; n17147_not
g81014 not n14294 ; n14294_not
g81015 not n17183 ; n17183_not
g81016 not n32195 ; n32195_not
g81017 not n13745 ; n13745_not
g81018 not n42590 ; n42590_not
g81019 not n55055 ; n55055_not
g81020 not n14348 ; n14348_not
g81021 not n17174 ; n17174_not
g81022 not n14357 ; n14357_not
g81023 not n14339 ; n14339_not
g81024 not n14366 ; n14366_not
g81025 not n33671 ; n33671_not
g81026 not n43535 ; n43535_not
g81027 not n32168 ; n32168_not
g81028 not n33680 ; n33680_not
g81029 not n32186 ; n32186_not
g81030 not n14384 ; n14384_not
g81031 not n55037 ; n55037_not
g81032 not n47171 ; n47171_not
g81033 not n32177 ; n32177_not
g81034 not n33635 ; n33635_not
g81035 not n17660 ; n17660_not
g81036 not n43571 ; n43571_not
g81037 not n32384 ; n32384_not
g81038 not n13835 ; n13835_not
g81039 not n14492 ; n14492_not
g81040 not n54119 ; n54119_not
g81041 not n14159 ; n14159_not
g81042 not n42518 ; n42518_not
g81043 not n50267 ; n50267_not
g81044 not n17615 ; n17615_not
g81045 not n55127 ; n55127_not
g81046 not n42545 ; n42545_not
g81047 not n17642 ; n17642_not
g81048 not n14168 ; n14168_not
g81049 not n43751 ; n43751_not
g81050 not n32375 ; n32375_not
g81051 not n37730 ; n37730_not
g81052 not n50258 ; n50258_not
g81053 not n17732 ; n17732_not
g81054 not n43580 ; n43580_not
g81055 not n33617 ; n33617_not
g81056 not n47207 ; n47207_not
g81057 not n47216 ; n47216_not
g81058 not n33626 ; n33626_not
g81059 not n17705 ; n17705_not
g81060 not n17714 ; n17714_not
g81061 not n42554 ; n42554_not
g81062 not n14519 ; n14519_not
g81063 not n42608 ; n42608_not
g81064 not n54920 ; n54920_not
g81065 not n32078 ; n32078_not
g81066 not n54911 ; n54911_not
g81067 not n17066 ; n17066_not
g81068 not n37046 ; n37046_not
g81069 not n14447 ; n14447_not
g81070 not n13781 ; n13781_not
g81071 not n14177 ; n14177_not
g81072 not n13790 ; n13790_not
g81073 not n45263 ; n45263_not
g81074 not n32357 ; n32357_not
g81075 not n43562 ; n43562_not
g81076 not n42563 ; n42563_not
g81077 not n14474 ; n14474_not
g81078 not n17633 ; n17633_not
g81079 not n54902 ; n54902_not
g81080 not n14456 ; n14456_not
g81081 not n15680 ; n15680_not
g81082 not n31475 ; n31475_not
g81083 not n16157 ; n16157_not
g81084 not n32663 ; n32663_not
g81085 not n41537 ; n41537_not
g81086 not n18560 ; n18560_not
g81087 not n45317 ; n45317_not
g81088 not n31493 ; n31493_not
g81089 not n16175 ; n16175_not
g81090 not n18524 ; n18524_not
g81091 not n54506 ; n54506_not
g81092 not n47126 ; n47126_not
g81093 not n33581 ; n33581_not
g81094 not n41546 ; n41546_not
g81095 not n18542 ; n18542_not
g81096 not n16166 ; n16166_not
g81097 not n41519 ; n41519_not
g81098 not n32645 ; n32645_not
g81099 not n54470 ; n54470_not
g81100 not n54461 ; n54461_not
g81101 not n14375 ; n14375_not
g81102 not n18614 ; n18614_not
g81103 not n47117 ; n47117_not
g81104 not n31466 ; n31466_not
g81105 not n16148 ; n16148_not
g81106 not n32654 ; n32654_not
g81107 not n33572 ; n33572_not
g81108 not n41528 ; n41528_not
g81109 not n48008 ; n48008_not
g81110 not n44903 ; n44903_not
g81111 not n43139 ; n43139_not
g81112 not n16139 ; n16139_not
g81113 not n41573 ; n41573_not
g81114 not n42167 ; n42167_not
g81115 not n33608 ; n33608_not
g81116 not n18083 ; n18083_not
g81117 not n55613 ; n55613_not
g81118 not n41951 ; n41951_not
g81119 not n37091 ; n37091_not
g81120 not n18074 ; n18074_not
g81121 not n16229 ; n16229_not
g81122 not n18065 ; n18065_not
g81123 not n18470 ; n18470_not
g81124 not n41564 ; n41564_not
g81125 not n42176 ; n42176_not
g81126 not n18137 ; n18137_not
g81127 not n31529 ; n31529_not
g81128 not n18128 ; n18128_not
g81129 not n43085 ; n43085_not
g81130 not n16247 ; n16247_not
g81131 not n18119 ; n18119_not
g81132 not n15635 ; n15635_not
g81133 not n18452 ; n18452_not
g81134 not n16238 ; n16238_not
g81135 not n18092 ; n18092_not
g81136 not n16193 ; n16193_not
g81137 not n33590 ; n33590_not
g81138 not n16184 ; n16184_not
g81139 not n55604 ; n55604_not
g81140 not n41555 ; n41555_not
g81141 not n54515 ; n54515_not
g81142 not n42149 ; n42149_not
g81143 not n18515 ; n18515_not
g81144 not n44912 ; n44912_not
g81145 not n18056 ; n18056_not
g81146 not n43094 ; n43094_not
g81147 not n42158 ; n42158_not
g81148 not n55028 ; n55028_not
g81149 not n54524 ; n54524_not
g81150 not n45119 ; n45119_not
g81151 not n31376 ; n31376_not
g81152 not n18731 ; n18731_not
g81153 not n31187 ; n31187_not
g81154 not n54371 ; n54371_not
g81155 not n32609 ; n32609_not
g81156 not n18740 ; n18740_not
g81157 not n41447 ; n41447_not
g81158 not n42059 ; n42059_not
g81159 not n18704 ; n18704_not
g81160 not n45047 ; n45047_not
g81161 not n31385 ; n31385_not
g81162 not n18713 ; n18713_not
g81163 not n54407 ; n54407_not
g81164 not n32618 ; n32618_not
g81165 not n18722 ; n18722_not
g81166 not n33536 ; n33536_not
g81167 not n41456 ; n41456_not
g81168 not n53570 ; n53570_not
g81169 not n43229 ; n43229_not
g81170 not n31349 ; n31349_not
g81171 not n47108 ; n47108_not
g81172 not n54353 ; n54353_not
g81173 not n33518 ; n33518_not
g81174 not n53606 ; n53606_not
g81175 not n44039 ; n44039_not
g81176 not n53615 ; n53615_not
g81177 not n31367 ; n31367_not
g81178 not n15770 ; n15770_not
g81179 not n54380 ; n54380_not
g81180 not n55550 ; n55550_not
g81181 not n53561 ; n53561_not
g81182 not n33527 ; n33527_not
g81183 not n31358 ; n31358_not
g81184 not n16085 ; n16085_not
g81185 not n54452 ; n54452_not
g81186 not n41492 ; n41492_not
g81187 not n15725 ; n15725_not
g81188 not n16076 ; n16076_not
g81189 not n18641 ; n18641_not
g81190 not n54344 ; n54344_not
g81191 not n42086 ; n42086_not
g81192 not n45326 ; n45326_not
g81193 not n18650 ; n18650_not
g81194 not n33554 ; n33554_not
g81195 not n33563 ; n33563_not
g81196 not n31448 ; n31448_not
g81197 not n18623 ; n18623_not
g81198 not n16094 ; n16094_not
g81199 not n42095 ; n42095_not
g81200 not n18632 ; n18632_not
g81201 not n42068 ; n42068_not
g81202 not n33545 ; n33545_not
g81203 not n54425 ; n54425_not
g81204 not n43184 ; n43184_not
g81205 not n16049 ; n16049_not
g81206 not n41465 ; n41465_not
g81207 not n54416 ; n54416_not
g81208 not n31394 ; n31394_not
g81209 not n54443 ; n54443_not
g81210 not n33293 ; n33293_not
g81211 not n41483 ; n41483_not
g81212 not n16067 ; n16067_not
g81213 not n42077 ; n42077_not
g81214 not n18533 ; n18533_not
g81215 not n54434 ; n54434_not
g81216 not n13286 ; n13286_not
g81217 not n16058 ; n16058_not
g81218 not n41474 ; n41474_not
g81219 not n31673 ; n31673_not
g81220 not n42275 ; n42275_not
g81221 not n16535 ; n16535_not
g81222 not n54614 ; n54614_not
g81223 not n18182 ; n18182_not
g81224 not n31664 ; n31664_not
g81225 not n54254 ; n54254_not
g81226 not n18191 ; n18191_not
g81227 not n54605 ; n54605_not
g81228 not n43931 ; n43931_not
g81229 not n37019 ; n37019_not
g81230 not n13754 ; n13754_not
g81231 not n42284 ; n42284_not
g81232 not n55640 ; n55640_not
g81233 not n45137 ; n45137_not
g81234 not n16490 ; n16490_not
g81235 not n18164 ; n18164_not
g81236 not n18173 ; n18173_not
g81237 not n18236 ; n18236_not
g81238 not n55271 ; n55271_not
g81239 not n55910 ; n55910_not
g81240 not n31637 ; n31637_not
g81241 not n32627 ; n32627_not
g81242 not n42248 ; n42248_not
g81243 not n43940 ; n43940_not
g81244 not n41906 ; n41906_not
g81245 not n55631 ; n55631_not
g81246 not n18245 ; n18245_not
g81247 not n31628 ; n31628_not
g81248 not n33644 ; n33644_not
g81249 not n16526 ; n16526_not
g81250 not n42266 ; n42266_not
g81251 not n31655 ; n31655_not
g81252 not n18209 ; n18209_not
g81253 not n55262 ; n55262_not
g81254 not n14465 ; n14465_not
g81255 not n18218 ; n18218_not
g81256 not n16508 ; n16508_not
g81257 not n31646 ; n31646_not
g81258 not n31439 ; n31439_not
g81259 not n42257 ; n42257_not
g81260 not n44372 ; n44372_not
g81261 not n18227 ; n18227_not
g81262 not n16454 ; n16454_not
g81263 not n54650 ; n54650_not
g81264 not n16463 ; n16463_not
g81265 not n54641 ; n54641_not
g81266 not n37703 ; n37703_not
g81267 not n16445 ; n16445_not
g81268 not n45281 ; n45281_not
g81269 not n43292 ; n43292_not
g81270 not n43904 ; n43904_not
g81271 not n31736 ; n31736_not
g81272 not n43058 ; n43058_not
g81273 not n45290 ; n45290_not
g81274 not n32582 ; n32582_not
g81275 not n18146 ; n18146_not
g81276 not n45146 ; n45146_not
g81277 not n17723 ; n17723_not
g81278 not n55253 ; n55253_not
g81279 not n43067 ; n43067_not
g81280 not n54623 ; n54623_not
g81281 not n31691 ; n31691_not
g81282 not n18155 ; n18155_not
g81283 not n43913 ; n43913_not
g81284 not n54632 ; n54632_not
g81285 not n55622 ; n55622_not
g81286 not n42293 ; n42293_not
g81287 not n42464 ; n42464_not
g81288 not n47306 ; n47306_not
g81289 not n13196 ; n13196_not
g81290 not n31565 ; n31565_not
g81291 not n31484 ; n31484_not
g81292 not n42194 ; n42194_not
g81293 not n32690 ; n32690_not
g81294 not n41609 ; n41609_not
g81295 not n18272 ; n18272_not
g81296 not n18263 ; n18263_not
g81297 not n18362 ; n18362_not
g81298 not n31574 ; n31574_not
g81299 not n18254 ; n18254_not
g81300 not n16337 ; n16337_not
g81301 not n43049 ; n43049_not
g81302 not n31547 ; n31547_not
g81303 not n16256 ; n16256_not
g81304 not n18407 ; n18407_not
g81305 not n45308 ; n45308_not
g81306 not n41582 ; n41582_not
g81307 not n31538 ; n31538_not
g81308 not n31556 ; n31556_not
g81309 not n16292 ; n16292_not
g81310 not n41591 ; n41591_not
g81311 not n44921 ; n44921_not
g81312 not n43076 ; n43076_not
g81313 not n54533 ; n54533_not
g81314 not n42185 ; n42185_not
g81315 not n18281 ; n18281_not
g81316 not n41627 ; n41627_not
g81317 not n18290 ; n18290_not
g81318 not n34076 ; n34076_not
g81319 not n54551 ; n54551_not
g81320 not n55280 ; n55280_not
g81321 not n18308 ; n18308_not
g81322 not n42239 ; n42239_not
g81323 not n16472 ; n16472_not
g81324 not n31619 ; n31619_not
g81325 not n44930 ; n44930_not
g81326 not n54560 ; n54560_not
g81327 not n16382 ; n16382_not
g81328 not n32672 ; n32672_not
g81329 not n31583 ; n31583_not
g81330 not n54542 ; n54542_not
g81331 not n41618 ; n41618_not
g81332 not n55208 ; n55208_not
g81333 not n16427 ; n16427_not
g81334 not n18326 ; n18326_not
g81335 not n31592 ; n31592_not
g81336 not n45029 ; n45029_not
g81337 not n24293 ; n24293_not
g81338 not n51266 ; n51266_not
g81339 not n35363 ; n35363_not
g81340 not n23654 ; n23654_not
g81341 not n45830 ; n45830_not
g81342 not n46550 ; n46550_not
g81343 not n52850 ; n52850_not
g81344 not n51833 ; n51833_not
g81345 not n24329 ; n24329_not
g81346 not n49214 ; n49214_not
g81347 not n56720 ; n56720_not
g81348 not n52643 ; n52643_not
g81349 not n24338 ; n24338_not
g81350 not n10784 ; n10784_not
g81351 not n35318 ; n35318_not
g81352 not n24347 ; n24347_not
g81353 not n40079 ; n40079_not
g81354 not n57062 ; n57062_not
g81355 not n29027 ; n29027_not
g81356 not n44444 ; n44444_not
g81357 not n27830 ; n27830_not
g81358 not n49205 ; n49205_not
g81359 not n29054 ; n29054_not
g81360 not n35354 ; n35354_not
g81361 not n24266 ; n24266_not
g81362 not n10838 ; n10838_not
g81363 not n10829 ; n10829_not
g81364 not n46091 ; n46091_not
g81365 not n24275 ; n24275_not
g81366 not n23672 ; n23672_not
g81367 not n29045 ; n29045_not
g81368 not n36407 ; n36407_not
g81369 not n10793 ; n10793_not
g81370 not n24284 ; n24284_not
g81371 not n23663 ; n23663_not
g81372 not n40646 ; n40646_not
g81373 not n44741 ; n44741_not
g81374 not n51275 ; n51275_not
g81375 not n35372 ; n35372_not
g81376 not n46082 ; n46082_not
g81377 not n29009 ; n29009_not
g81378 not n49223 ; n49223_not
g81379 not n24383 ; n24383_not
g81380 not n24374 ; n24374_not
g81381 not n24428 ; n24428_not
g81382 not n24365 ; n24365_not
g81383 not n24356 ; n24356_not
g81384 not n51284 ; n51284_not
g81385 not n46073 ; n46073_not
g81386 not n36092 ; n36092_not
g81387 not n24446 ; n24446_not
g81388 not n36416 ; n36416_not
g81389 not n10766 ; n10766_not
g81390 not n52841 ; n52841_not
g81391 not n23627 ; n23627_not
g81392 not n40619 ; n40619_not
g81393 not n35930 ; n35930_not
g81394 not n40088 ; n40088_not
g81395 not n23618 ; n23618_not
g81396 not n56270 ; n56270_not
g81397 not n10775 ; n10775_not
g81398 not n29018 ; n29018_not
g81399 not n56621 ; n56621_not
g81400 not n23609 ; n23609_not
g81401 not n24392 ; n24392_not
g81402 not n52832 ; n52832_not
g81403 not n29108 ; n29108_not
g81404 not n52922 ; n52922_not
g81405 not n47027 ; n47027_not
g81406 not n49160 ; n49160_not
g81407 not n46118 ; n46118_not
g81408 not n27803 ; n27803_not
g81409 not n40727 ; n40727_not
g81410 not n23762 ; n23762_not
g81411 not n23753 ; n23753_not
g81412 not n35327 ; n35327_not
g81413 not n52913 ; n52913_not
g81414 not n26192 ; n26192_not
g81415 not n46406 ; n46406_not
g81416 not n51248 ; n51248_not
g81417 not n34940 ; n34940_not
g81418 not n23744 ; n23744_not
g81419 not n29090 ; n29090_not
g81420 not n49142 ; n49142_not
g81421 not n23807 ; n23807_not
g81422 not n49151 ; n49151_not
g81423 not n40754 ; n40754_not
g81424 not n51239 ; n51239_not
g81425 not n24059 ; n24059_not
g81426 not n10892 ; n10892_not
g81427 not n52940 ; n52940_not
g81428 not n24068 ; n24068_not
g81429 not n24077 ; n24077_not
g81430 not n24086 ; n24086_not
g81431 not n52931 ; n52931_not
g81432 not n40736 ; n40736_not
g81433 not n24095 ; n24095_not
g81434 not n56261 ; n56261_not
g81435 not n10847 ; n10847_not
g81436 not n45821 ; n45821_not
g81437 not n10874 ; n10874_not
g81438 not n29072 ; n29072_not
g81439 not n40691 ; n40691_not
g81440 not n45524 ; n45524_not
g81441 not n44318 ; n44318_not
g81442 not n40682 ; n40682_not
g81443 not n24239 ; n24239_not
g81444 not n27821 ; n27821_not
g81445 not n24248 ; n24248_not
g81446 not n56612 ; n56612_not
g81447 not n35336 ; n35336_not
g81448 not n51842 ; n51842_not
g81449 not n24257 ; n24257_not
g81450 not n40664 ; n40664_not
g81451 not n24149 ; n24149_not
g81452 not n52292 ; n52292_not
g81453 not n24158 ; n24158_not
g81454 not n40709 ; n40709_not
g81455 not n52607 ; n52607_not
g81456 not n24167 ; n24167_not
g81457 not n24176 ; n24176_not
g81458 not n52904 ; n52904_not
g81459 not n24185 ; n24185_not
g81460 not n56603 ; n56603_not
g81461 not n51257 ; n51257_not
g81462 not n24194 ; n24194_not
g81463 not n46109 ; n46109_not
g81464 not n23717 ; n23717_not
g81465 not n52616 ; n52616_not
g81466 not n23708 ; n23708_not
g81467 not n57035 ; n57035_not
g81468 not n38612 ; n38612_not
g81469 not n23924 ; n23924_not
g81470 not n24680 ; n24680_not
g81471 not n23915 ; n23915_not
g81472 not n52337 ; n52337_not
g81473 not n10649 ; n10649_not
g81474 not n39170 ; n39170_not
g81475 not n28064 ; n28064_not
g81476 not n23906 ; n23906_not
g81477 not n51383 ; n51383_not
g81478 not n36074 ; n36074_not
g81479 not n44309 ; n44309_not
g81480 not n10595 ; n10595_not
g81481 not n51329 ; n51329_not
g81482 not n35417 ; n35417_not
g81483 not n40565 ; n40565_not
g81484 not n51392 ; n51392_not
g81485 not n36821 ; n36821_not
g81486 not n10586 ; n10586_not
g81487 not n40583 ; n40583_not
g81488 not n52814 ; n52814_not
g81489 not n26246 ; n26246_not
g81490 not n24653 ; n24653_not
g81491 not n23960 ; n23960_not
g81492 not n23951 ; n23951_not
g81493 not n48710 ; n48710_not
g81494 not n10667 ; n10667_not
g81495 not n51365 ; n51365_not
g81496 not n10658 ; n10658_not
g81497 not n35408 ; n35408_not
g81498 not n46037 ; n46037_not
g81499 not n23942 ; n23942_not
g81500 not n52805 ; n52805_not
g81501 not n23933 ; n23933_not
g81502 not n40574 ; n40574_not
g81503 not n24671 ; n24671_not
g81504 not n51374 ; n51374_not
g81505 not n26255 ; n26255_not
g81506 not n38630 ; n38630_not
g81507 not n24743 ; n24743_not
g81508 not n57026 ; n57026_not
g81509 not n51347 ; n51347_not
g81510 not n10568 ; n10568_not
g81511 not n10496 ; n10496_not
g81512 not n24752 ; n24752_not
g81513 not n10559 ; n10559_not
g81514 not n35435 ; n35435_not
g81515 not n52346 ; n52346_not
g81516 not n40547 ; n40547_not
g81517 not n28802 ; n28802_not
g81518 not n57017 ; n57017_not
g81519 not n24761 ; n24761_not
g81520 not n24770 ; n24770_not
g81521 not n40538 ; n40538_not
g81522 not n35039 ; n35039_not
g81523 not n46028 ; n46028_not
g81524 not n36443 ; n36443_not
g81525 not n10487 ; n10487_not
g81526 not n49322 ; n49322_not
g81527 not n24716 ; n24716_not
g81528 not n35291 ; n35291_not
g81529 not n24725 ; n24725_not
g81530 not n56306 ; n56306_not
g81531 not n10577 ; n10577_not
g81532 not n28136 ; n28136_not
g81533 not n35426 ; n35426_not
g81534 not n28820 ; n28820_not
g81535 not n46019 ; n46019_not
g81536 not n51338 ; n51338_not
g81537 not n40556 ; n40556_not
g81538 not n24734 ; n24734_not
g81539 not n35282 ; n35282_not
g81540 not n36083 ; n36083_not
g81541 not n39800 ; n39800_not
g81542 not n24536 ; n24536_not
g81543 not n24545 ; n24545_not
g81544 not n10748 ; n10748_not
g81545 not n46064 ; n46064_not
g81546 not n10397 ; n10397_not
g81547 not n47018 ; n47018_not
g81548 not n36425 ; n36425_not
g81549 not n24563 ; n24563_not
g81550 not n10739 ; n10739_not
g81551 not n24455 ; n24455_not
g81552 not n51293 ; n51293_not
g81553 not n10757 ; n10757_not
g81554 not n35921 ; n35921_not
g81555 not n24473 ; n24473_not
g81556 not n35381 ; n35381_not
g81557 not n24491 ; n24491_not
g81558 not n52652 ; n52652_not
g81559 not n24518 ; n24518_not
g81560 not n35912 ; n35912_not
g81561 not n51815 ; n51815_not
g81562 not n36830 ; n36830_not
g81563 not n24608 ; n24608_not
g81564 not n36434 ; n36434_not
g81565 not n57044 ; n57044_not
g81566 not n46046 ; n46046_not
g81567 not n24626 ; n24626_not
g81568 not n24635 ; n24635_not
g81569 not n52328 ; n52328_not
g81570 not n52661 ; n52661_not
g81571 not n51356 ; n51356_not
g81572 not n10685 ; n10685_not
g81573 not n35903 ; n35903_not
g81574 not n10676 ; n10676_not
g81575 not n40592 ; n40592_not
g81576 not n52319 ; n52319_not
g81577 not n35390 ; n35390_not
g81578 not n56630 ; n56630_not
g81579 not n26237 ; n26237_not
g81580 not n44570 ; n44570_not
g81581 not n24581 ; n24581_not
g81582 not n44336 ; n44336_not
g81583 not n56711 ; n56711_not
g81584 not n46055 ; n46055_not
g81585 not n28910 ; n28910_not
g81586 not n52823 ; n52823_not
g81587 not n24590 ; n24590_not
g81588 not n10694 ; n10694_not
g81589 not n23096 ; n23096_not
g81590 not n36902 ; n36902_not
g81591 not n51194 ; n51194_not
g81592 not n51176 ; n51176_not
g81593 not n10955 ; n10955_not
g81594 not n40925 ; n40925_not
g81595 not n47063 ; n47063_not
g81596 not n44291 ; n44291_not
g81597 not n39134 ; n39134_not
g81598 not n10964 ; n10964_not
g81599 not n49106 ; n49106_not
g81600 not n56036 ; n56036_not
g81601 not n48701 ; n48701_not
g81602 not n10973 ; n10973_not
g81603 not n29423 ; n29423_not
g81604 not n22853 ; n22853_not
g81605 not n36119 ; n36119_not
g81606 not n47072 ; n47072_not
g81607 not n29360 ; n29360_not
g81608 not n46523 ; n46523_not
g81609 not n29414 ; n29414_not
g81610 not n56234 ; n56234_not
g81611 not n51185 ; n51185_not
g81612 not n53066 ; n53066_not
g81613 not n36362 ; n36362_not
g81614 not n29405 ; n29405_not
g81615 not n46163 ; n46163_not
g81616 not n22844 ; n22844_not
g81617 not n35633 ; n35633_not
g81618 not n51068 ; n51068_not
g81619 not n26921 ; n26921_not
g81620 not n53057 ; n53057_not
g81621 not n52265 ; n52265_not
g81622 not n29342 ; n29342_not
g81623 not n56243 ; n56243_not
g81624 not n57134 ; n57134_not
g81625 not n35174 ; n35174_not
g81626 not n38504 ; n38504_not
g81627 not n40916 ; n40916_not
g81628 not n29333 ; n29333_not
g81629 not n35165 ; n35165_not
g81630 not n46532 ; n46532_not
g81631 not n26930 ; n26930_not
g81632 not n35183 ; n35183_not
g81633 not n51059 ; n51059_not
g81634 not n22817 ; n22817_not
g81635 not n52526 ; n52526_not
g81636 not n39701 ; n39701_not
g81637 not n56531 ; n56531_not
g81638 not n29306 ; n29306_not
g81639 not n22808 ; n22808_not
g81640 not n49412 ; n49412_not
g81641 not n29315 ; n29315_not
g81642 not n47054 ; n47054_not
g81643 not n35192 ; n35192_not
g81644 not n26156 ; n26156_not
g81645 not n29324 ; n29324_not
g81646 not n49052 ; n49052_not
g81647 not n53084 ; n53084_not
g81648 not n46190 ; n46190_not
g81649 not n51149 ; n51149_not
g81650 not n40781 ; n40781_not
g81651 not n40952 ; n40952_not
g81652 not n51158 ; n51158_not
g81653 not n38423 ; n38423_not
g81654 not n57170 ; n57170_not
g81655 not n44282 ; n44282_not
g81656 not n46181 ; n46181_not
g81657 not n47090 ; n47090_not
g81658 not n56504 ; n56504_not
g81659 not n40790 ; n40790_not
g81660 not n52256 ; n52256_not
g81661 not n36353 ; n36353_not
g81662 not n29513 ; n29513_not
g81663 not n38414 ; n38414_not
g81664 not n51905 ; n51905_not
g81665 not n52247 ; n52247_not
g81666 not n39125 ; n39125_not
g81667 not n29504 ; n29504_not
g81668 not n22907 ; n22907_not
g81669 not n35606 ; n35606_not
g81670 not n52508 ; n52508_not
g81671 not n10883 ; n10883_not
g81672 not n34733 ; n34733_not
g81673 not n26147 ; n26147_not
g81674 not n36911 ; n36911_not
g81675 not n36542 ; n36542_not
g81676 not n56513 ; n56513_not
g81677 not n51167 ; n51167_not
g81678 not n29441 ; n29441_not
g81679 not n10928 ; n10928_not
g81680 not n49070 ; n49070_not
g81681 not n49430 ; n49430_not
g81682 not n40934 ; n40934_not
g81683 not n29432 ; n29432_not
g81684 not n38450 ; n38450_not
g81685 not n22862 ; n22862_not
g81686 not n51077 ; n51077_not
g81687 not n44606 ; n44606_not
g81688 not n56522 ; n56522_not
g81689 not n52517 ; n52517_not
g81690 not n40943 ; n40943_not
g81691 not n34742 ; n34742_not
g81692 not n38432 ; n38432_not
g81693 not n49061 ; n49061_not
g81694 not n57161 ; n57161_not
g81695 not n46172 ; n46172_not
g81696 not n29450 ; n29450_not
g81697 not n53075 ; n53075_not
g81698 not n38441 ; n38441_not
g81699 not n10919 ; n10919_not
g81700 not n34751 ; n34751_not
g81701 not n47081 ; n47081_not
g81702 not n40844 ; n40844_not
g81703 not n29180 ; n29180_not
g81704 not n35651 ; n35651_not
g81705 not n40826 ; n40826_not
g81706 not n40817 ; n40817_not
g81707 not n29171 ; n29171_not
g81708 not n10937 ; n10937_not
g81709 not n57107 ; n57107_not
g81710 not n52553 ; n52553_not
g81711 not n49115 ; n49115_not
g81712 not n23852 ; n23852_not
g81713 not n52274 ; n52274_not
g81714 not n29207 ; n29207_not
g81715 not n35048 ; n35048_not
g81716 not n46145 ; n46145_not
g81717 not n57116 ; n57116_not
g81718 not n40835 ; n40835_not
g81719 not n23861 ; n23861_not
g81720 not n35273 ; n35273_not
g81721 not n49124 ; n49124_not
g81722 not n52283 ; n52283_not
g81723 not n29144 ; n29144_not
g81724 not n49133 ; n49133_not
g81725 not n40772 ; n40772_not
g81726 not n29135 ; n29135_not
g81727 not n29081 ; n29081_not
g81728 not n46127 ; n46127_not
g81729 not n46136 ; n46136_not
g81730 not n23843 ; n23843_not
g81731 not n47036 ; n47036_not
g81732 not n29153 ; n29153_not
g81733 not n51707 ; n51707_not
g81734 not n52562 ; n52562_not
g81735 not n51860 ; n51860_not
g81736 not n44732 ; n44732_not
g81737 not n36380 ; n36380_not
g81738 not n23834 ; n23834_not
g81739 not n45515 ; n45515_not
g81740 not n52571 ; n52571_not
g81741 not n35129 ; n35129_not
g81742 not n38522 ; n38522_not
g81743 not n29270 ; n29270_not
g81744 not n35228 ; n35228_not
g81745 not n23726 ; n23726_not
g81746 not n35237 ; n35237_not
g81747 not n26165 ; n26165_not
g81748 not n53048 ; n53048_not
g81749 not n29243 ; n29243_not
g81750 not n56540 ; n56540_not
g81751 not n23636 ; n23636_not
g81752 not n39143 ; n39143_not
g81753 not n35156 ; n35156_not
g81754 not n35147 ; n35147_not
g81755 not n47045 ; n47045_not
g81756 not n40907 ; n40907_not
g81757 not n56252 ; n56252_not
g81758 not n35138 ; n35138_not
g81759 not n23681 ; n23681_not
g81760 not n35075 ; n35075_not
g81761 not n35255 ; n35255_not
g81762 not n29225 ; n29225_not
g81763 not n23816 ; n23816_not
g81764 not n35066 ; n35066_not
g81765 not n29216 ; n29216_not
g81766 not n51716 ; n51716_not
g81767 not n38540 ; n38540_not
g81768 not n35057 ; n35057_not
g81769 not n53039 ; n53039_not
g81770 not n29252 ; n29252_not
g81771 not n40880 ; n40880_not
g81772 not n35093 ; n35093_not
g81773 not n44804 ; n44804_not
g81774 not n45506 ; n45506_not
g81775 not n23771 ; n23771_not
g81776 not n46154 ; n46154_not
g81777 not n36371 ; n36371_not
g81778 not n35084 ; n35084_not
g81779 not n10982 ; n10982_not
g81780 not n29234 ; n29234_not
g81781 not n35642 ; n35642_not
g81782 not n35471 ; n35471_not
g81783 not n44516 ; n44516_not
g81784 not n45425 ; n45425_not
g81785 not n28370 ; n28370_not
g81786 not n40286 ; n40286_not
g81787 not n25436 ; n25436_not
g81788 not n36623 ; n36623_not
g81789 not n38405 ; n38405_not
g81790 not n35462 ; n35462_not
g81791 not n40277 ; n40277_not
g81792 not n51626 ; n51626_not
g81793 not n45605 ; n45605_not
g81794 not n26354 ; n26354_not
g81795 not n25553 ; n25553_not
g81796 not n45434 ; n45434_not
g81797 not n25562 ; n25562_not
g81798 not n35453 ; n35453_not
g81799 not n25706 ; n25706_not
g81800 not n46631 ; n46631_not
g81801 not n40268 ; n40268_not
g81802 not n45416 ; n45416_not
g81803 not n38513 ; n38513_not
g81804 not n35480 ; n35480_not
g81805 not n35732 ; n35732_not
g81806 not n39062 ; n39062_not
g81807 not n48611 ; n48611_not
g81808 not n25670 ; n25670_not
g81809 not n35813 ; n35813_not
g81810 not n28073 ; n28073_not
g81811 not n46541 ; n46541_not
g81812 not n25544 ; n25544_not
g81813 not n25571 ; n25571_not
g81814 not n45443 ; n45443_not
g81815 not n36506 ; n36506_not
g81816 not n28091 ; n28091_not
g81817 not n25391 ; n25391_not
g81818 not n45623 ; n45623_not
g81819 not n27227 ; n27227_not
g81820 not n25580 ; n25580_not
g81821 not n39044 ; n39044_not
g81822 not n51617 ; n51617_not
g81823 not n28325 ; n28325_not
g81824 not n45632 ; n45632_not
g81825 not n45452 ; n45452_not
g81826 not n25805 ; n25805_not
g81827 not n35705 ; n35705_not
g81828 not n25715 ; n25715_not
g81829 not n25724 ; n25724_not
g81830 not n40259 ; n40259_not
g81831 not n35444 ; n35444_not
g81832 not n25733 ; n25733_not
g81833 not n28352 ; n28352_not
g81834 not n25409 ; n25409_not
g81835 not n36614 ; n36614_not
g81836 not n51635 ; n51635_not
g81837 not n45614 ; n45614_not
g81838 not n25742 ; n25742_not
g81839 not n35741 ; n35741_not
g81840 not n28343 ; n28343_not
g81841 not n25751 ; n25751_not
g81842 not n52535 ; n52535_not
g81843 not n25760 ; n25760_not
g81844 not n25526 ; n25526_not
g81845 not n28442 ; n28442_not
g81846 not n51608 ; n51608_not
g81847 not n35516 ; n35516_not
g81848 not n40358 ; n40358_not
g81849 not n46820 ; n46820_not
g81850 not n52391 ; n52391_not
g81851 not n36047 ; n36047_not
g81852 not n45407 ; n45407_not
g81853 not n35507 ; n35507_not
g81854 not n28424 ; n28424_not
g81855 not n40349 ; n40349_not
g81856 not n35552 ; n35552_not
g81857 not n28460 ; n28460_not
g81858 not n38351 ; n38351_not
g81859 not n39602 ; n39602_not
g81860 not n35543 ; n35543_not
g81861 not n25508 ; n25508_not
g81862 not n35534 ; n35534_not
g81863 not n35660 ; n35660_not
g81864 not n35525 ; n35525_not
g81865 not n38360 ; n38360_not
g81866 not n44462 ; n44462_not
g81867 not n28406 ; n28406_not
g81868 not n48602 ; n48602_not
g81869 not n25625 ; n25625_not
g81870 not n46802 ; n46802_not
g81871 not n28055 ; n28055_not
g81872 not n25634 ; n25634_not
g81873 not n26372 ; n26372_not
g81874 not n25643 ; n25643_not
g81875 not n36641 ; n36641_not
g81876 not n55811 ; n55811_not
g81877 not n25652 ; n25652_not
g81878 not n56900 ; n56900_not
g81879 not n25454 ; n25454_not
g81880 not n25661 ; n25661_not
g81881 not n40295 ; n40295_not
g81882 not n25445 ; n25445_not
g81883 not n51455 ; n51455_not
g81884 not n50834 ; n50834_not
g81885 not n46811 ; n46811_not
g81886 not n28046 ; n28046_not
g81887 not n35822 ; n35822_not
g81888 not n25490 ; n25490_not
g81889 not n52580 ; n52580_not
g81890 not n25481 ; n25481_not
g81891 not n25607 ; n25607_not
g81892 not n25616 ; n25616_not
g81893 not n56810 ; n56810_not
g81894 not n28226 ; n28226_not
g81895 not n51536 ; n51536_not
g81896 not n26264 ; n26264_not
g81897 not n40097 ; n40097_not
g81898 not n45560 ; n45560_not
g81899 not n46703 ; n46703_not
g81900 not n26048 ; n26048_not
g81901 not n26039 ; n26039_not
g81902 not n26084 ; n26084_not
g81903 not n51527 ; n51527_not
g81904 not n52427 ; n52427_not
g81905 not n26129 ; n26129_not
g81906 not n25940 ; n25940_not
g81907 not n51518 ; n51518_not
g81908 not n45740 ; n45740_not
g81909 not n51545 ; n51545_not
g81910 not n45533 ; n45533_not
g81911 not n28244 ; n28244_not
g81912 not n52445 ; n52445_not
g81913 not n25274 ; n25274_not
g81914 not n26282 ; n26282_not
g81915 not n46721 ; n46721_not
g81916 not n25265 ; n25265_not
g81917 not n56801 ; n56801_not
g81918 not n25256 ; n25256_not
g81919 not n45542 ; n45542_not
g81920 not n28235 ; n28235_not
g81921 not n46712 ; n46712_not
g81922 not n25229 ; n25229_not
g81923 not n45551 ; n45551_not
g81924 not n51491 ; n51491_not
g81925 not n25841 ; n25841_not
g81926 not n25832 ; n25832_not
g81927 not n28019 ; n28019_not
g81928 not n28154 ; n28154_not
g81929 not n36524 ; n36524_not
g81930 not n28172 ; n28172_not
g81931 not n25823 ; n25823_not
g81932 not n51482 ; n51482_not
g81933 not n25814 ; n25814_not
g81934 not n26219 ; n26219_not
g81935 not n52409 ; n52409_not
g81936 not n36533 ; n36533_not
g81937 not n28163 ; n28163_not
g81938 not n39017 ; n39017_not
g81939 not n25931 ; n25931_not
g81940 not n25922 ; n25922_not
g81941 not n51509 ; n51509_not
g81942 not n25913 ; n25913_not
g81943 not n25904 ; n25904_not
g81944 not n36551 ; n36551_not
g81945 not n44543 ; n44543_not
g81946 not n45731 ; n45731_not
g81947 not n39530 ; n39530_not
g81948 not n26174 ; n26174_not
g81949 not n28181 ; n28181_not
g81950 not n25850 ; n25850_not
g81951 not n25346 ; n25346_not
g81952 not n40187 ; n40187_not
g81953 not n26327 ; n26327_not
g81954 not n45461 ; n45461_not
g81955 not n52490 ; n52490_not
g81956 not n51653 ; n51653_not
g81957 not n45470 ; n45470_not
g81958 not n51590 ; n51590_not
g81959 not n28109 ; n28109_not
g81960 not n40169 ; n40169_not
g81961 not n44534 ; n44534_not
g81962 not n26309 ; n26309_not
g81963 not n51464 ; n51464_not
g81964 not n26336 ; n26336_not
g81965 not n35804 ; n35804_not
g81966 not n45641 ; n45641_not
g81967 not n28316 ; n28316_not
g81968 not n25364 ; n25364_not
g81969 not n39035 ; n39035_not
g81970 not n25355 ; n25355_not
g81971 not n35723 ; n35723_not
g81972 not n51725 ; n51725_not
g81973 not n28307 ; n28307_not
g81974 not n45803 ; n45803_not
g81975 not n45650 ; n45650_not
g81976 not n51563 ; n51563_not
g81977 not n52463 ; n52463_not
g81978 not n46730 ; n46730_not
g81979 not n51554 ; n51554_not
g81980 not n28253 ; n28253_not
g81981 not n26291 ; n26291_not
g81982 not n28127 ; n28127_not
g81983 not n35750 ; n35750_not
g81984 not n45713 ; n45713_not
g81985 not n51680 ; n51680_not
g81986 not n51662 ; n51662_not
g81987 not n51581 ; n51581_not
g81988 not n52472 ; n52472_not
g81989 not n25319 ; n25319_not
g81990 not n51572 ; n51572_not
g81991 not n51473 ; n51473_not
g81992 not n28271 ; n28271_not
g81993 not n48620 ; n48620_not
g81994 not n40457 ; n40457_not
g81995 not n40178 ; n40178_not
g81996 not n45920 ; n45920_not
g81997 not n40448 ; n40448_not
g81998 not n56342 ; n56342_not
g81999 not n24509 ; n24509_not
g82000 not n25049 ; n25049_not
g82001 not n44264 ; n44264_not
g82002 not n46442 ; n46442_not
g82003 not n25058 ; n25058_not
g82004 not n28208 ; n28208_not
g82005 not n35246 ; n35246_not
g82006 not n28712 ; n28712_not
g82007 not n24941 ; n24941_not
g82008 not n56324 ; n56324_not
g82009 not n24950 ; n24950_not
g82010 not n38180 ; n38180_not
g82011 not n46433 ; n46433_not
g82012 not n40466 ; n40466_not
g82013 not n24554 ; n24554_not
g82014 not n56333 ; n56333_not
g82015 not n51770 ; n51770_not
g82016 not n36470 ; n36470_not
g82017 not n44273 ; n44273_not
g82018 not n28640 ; n28640_not
g82019 not n25094 ; n25094_not
g82020 not n52670 ; n52670_not
g82021 not n44246 ; n44246_not
g82022 not n45911 ; n45911_not
g82023 not n46451 ; n46451_not
g82024 not n44237 ; n44237_not
g82025 not n44228 ; n44228_not
g82026 not n24464 ; n24464_not
g82027 not n38225 ; n38225_not
g82028 not n38603 ; n38603_not
g82029 not n28622 ; n28622_not
g82030 not n25139 ; n25139_not
g82031 not n36038 ; n36038_not
g82032 not n25148 ; n25148_not
g82033 not n46613 ; n46613_not
g82034 not n56351 ; n56351_not
g82035 not n38207 ; n38207_not
g82036 not n25067 ; n25067_not
g82037 not n25076 ; n25076_not
g82038 not n40439 ; n40439_not
g82039 not n44255 ; n44255_not
g82040 not n56360 ; n56360_not
g82041 not n25085 ; n25085_not
g82042 not n44381 ; n44381_not
g82043 not n38216 ; n38216_not
g82044 not n52364 ; n52364_not
g82045 not n44561 ; n44561_not
g82046 not n24824 ; n24824_not
g82047 not n50942 ; n50942_not
g82048 not n52742 ; n52742_not
g82049 not n24833 ; n24833_not
g82050 not n27920 ; n27920_not
g82051 not n24842 ; n24842_not
g82052 not n51428 ; n51428_not
g82053 not n50933 ; n50933_not
g82054 not n10469 ; n10469_not
g82055 not n24851 ; n24851_not
g82056 not n24860 ; n24860_not
g82057 not n52706 ; n52706_not
g82058 not n51437 ; n51437_not
g82059 not n47009 ; n47009_not
g82060 not n36812 ; n36812_not
g82061 not n36452 ; n36452_not
g82062 not n27911 ; n27911_not
g82063 not n52760 ; n52760_not
g82064 not n56315 ; n56315_not
g82065 not n40529 ; n40529_not
g82066 not n52751 ; n52751_not
g82067 not n24644 ; n24644_not
g82068 not n24806 ; n24806_not
g82069 not n39152 ; n39152_not
g82070 not n51419 ; n51419_not
g82071 not n24815 ; n24815_not
g82072 not n50924 ; n50924_not
g82073 not n28730 ; n28730_not
g82074 not n24914 ; n24914_not
g82075 not n40484 ; n40484_not
g82076 not n24923 ; n24923_not
g82077 not n38162 ; n38162_not
g82078 not n24932 ; n24932_not
g82079 not n40475 ; n40475_not
g82080 not n38171 ; n38171_not
g82081 not n51671 ; n51671_not
g82082 not n38153 ; n38153_not
g82083 not n52733 ; n52733_not
g82084 not n36803 ; n36803_not
g82085 not n40493 ; n40493_not
g82086 not n10379 ; n10379_not
g82087 not n24905 ; n24905_not
g82088 not n51446 ; n51446_not
g82089 not n52355 ; n52355_not
g82090 not n36461 ; n36461_not
g82091 not n25418 ; n25418_not
g82092 not n45065 ; n45065_not
g82093 not n35840 ; n35840_not
g82094 not n38315 ; n38315_not
g82095 not n44453 ; n44453_not
g82096 not n28280 ; n28280_not
g82097 not n40385 ; n40385_not
g82098 not n35615 ; n35615_not
g82099 not n25373 ; n25373_not
g82100 not n28532 ; n28532_not
g82101 not n38306 ; n38306_not
g82102 not n36722 ; n36722_not
g82103 not n40394 ; n40394_not
g82104 not n48530 ; n48530_not
g82105 not n28514 ; n28514_not
g82106 not n44750 ; n44750_not
g82107 not n50843 ; n50843_not
g82108 not n35570 ; n35570_not
g82109 not n26345 ; n26345_not
g82110 not n38342 ; n38342_not
g82111 not n35561 ; n35561_not
g82112 not n28028 ; n28028_not
g82113 not n35831 ; n35831_not
g82114 not n40367 ; n40367_not
g82115 not n36713 ; n36713_not
g82116 not n38324 ; n38324_not
g82117 not n46640 ; n46640_not
g82118 not n52625 ; n52625_not
g82119 not n52382 ; n52382_not
g82120 not n50852 ; n50852_not
g82121 not n39080 ; n39080_not
g82122 not n36704 ; n36704_not
g82123 not n38333 ; n38333_not
g82124 not n44471 ; n44471_not
g82125 not n25463 ; n25463_not
g82126 not n40376 ; n40376_not
g82127 not n25184 ; n25184_not
g82128 not n25193 ; n25193_not
g82129 not n56432 ; n56432_not
g82130 not n24419 ; n24419_not
g82131 not n25238 ; n25238_not
g82132 not n44192 ; n44192_not
g82133 not n38252 ; n38252_not
g82134 not n56441 ; n56441_not
g82135 not n44183 ; n44183_not
g82136 not n39107 ; n39107_not
g82137 not n44219 ; n44219_not
g82138 not n38234 ; n38234_not
g82139 not n56405 ; n56405_not
g82140 not n25157 ; n25157_not
g82141 not n56414 ; n56414_not
g82142 not n28604 ; n28604_not
g82143 not n38243 ; n38243_not
g82144 not n25166 ; n25166_not
g82145 not n56423 ; n56423_not
g82146 not n25175 ; n25175_not
g82147 not n28550 ; n28550_not
g82148 not n44156 ; n44156_not
g82149 not n51743 ; n51743_not
g82150 not n25328 ; n25328_not
g82151 not n36740 ; n36740_not
g82152 not n46622 ; n46622_not
g82153 not n55901 ; n55901_not
g82154 not n36029 ; n36029_not
g82155 not n46901 ; n46901_not
g82156 not n36731 ; n36731_not
g82157 not n56450 ; n56450_not
g82158 not n51752 ; n51752_not
g82159 not n44174 ; n44174_not
g82160 not n36632 ; n36632_not
g82161 not n38261 ; n38261_not
g82162 not n52373 ; n52373_not
g82163 not n25283 ; n25283_not
g82164 not n44426 ; n44426_not
g82165 not n44165 ; n44165_not
g82166 not n46910 ; n46910_not
g82167 not n38270 ; n38270_not
g82168 not n20657 ; n20657_not
g82169 not n34607 ; n34607_not
g82170 not n20675 ; n20675_not
g82171 not n45704 ; n45704_not
g82172 not n30386 ; n30386_not
g82173 not n20684 ; n20684_not
g82174 not n20729 ; n20729_not
g82175 not n30377 ; n30377_not
g82176 not n27092 ; n27092_not
g82177 not n20747 ; n20747_not
g82178 not n48017 ; n48017_not
g82179 not n20765 ; n20765_not
g82180 not n27056 ; n27056_not
g82181 not n30368 ; n30368_not
g82182 not n53453 ; n53453_not
g82183 not n37073 ; n37073_not
g82184 not n41375 ; n41375_not
g82185 not n20495 ; n20495_not
g82186 not n36164 ; n36164_not
g82187 not n41393 ; n41393_not
g82188 not n34625 ; n34625_not
g82189 not n20549 ; n20549_not
g82190 not n27119 ; n27119_not
g82191 not n20567 ; n20567_not
g82192 not n46325 ; n46325_not
g82193 not n34616 ; n34616_not
g82194 not n20585 ; n20585_not
g82195 not n27065 ; n27065_not
g82196 not n20594 ; n20594_not
g82197 not n34850 ; n34850_not
g82198 not n20639 ; n20639_not
g82199 not n30395 ; n30395_not
g82200 not n44660 ; n44660_not
g82201 not n53426 ; n53426_not
g82202 not n34562 ; n34562_not
g82203 not n20693 ; n20693_not
g82204 not n36146 ; n36146_not
g82205 not n34553 ; n34553_not
g82206 not n50096 ; n50096_not
g82207 not n51806 ; n51806_not
g82208 not n34544 ; n34544_not
g82209 not n56153 ; n56153_not
g82210 not n20783 ; n20783_not
g82211 not n20792 ; n20792_not
g82212 not n34580 ; n34580_not
g82213 not n34571 ; n34571_not
g82214 not n20738 ; n20738_not
g82215 not n46316 ; n46316_not
g82216 not n27074 ; n27074_not
g82217 not n53435 ; n53435_not
g82218 not n41357 ; n41357_not
g82219 not n41348 ; n41348_not
g82220 not n53543 ; n53543_not
g82221 not n34814 ; n34814_not
g82222 not n30485 ; n30485_not
g82223 not n30467 ; n30467_not
g82224 not n36290 ; n36290_not
g82225 not n30476 ; n30476_not
g82226 not n34670 ; n34670_not
g82227 not n36173 ; n36173_not
g82228 not n53525 ; n53525_not
g82229 not n34706 ; n34706_not
g82230 not n12188 ; n12188_not
g82231 not n19910 ; n19910_not
g82232 not n34805 ; n34805_not
g82233 not n52094 ; n52094_not
g82234 not n53534 ; n53534_not
g82235 not n12098 ; n12098_not
g82236 not n46334 ; n46334_not
g82237 not n34643 ; n34643_not
g82238 not n53480 ; n53480_not
g82239 not n53471 ; n53471_not
g82240 not n30269 ; n30269_not
g82241 not n56144 ; n56144_not
g82242 not n34634 ; n34634_not
g82243 not n30278 ; n30278_not
g82244 not n53516 ; n53516_not
g82245 not n27146 ; n27146_not
g82246 not n27137 ; n27137_not
g82247 not n34661 ; n34661_not
g82248 not n40871 ; n40871_not
g82249 not n30458 ; n30458_not
g82250 not n19820 ; n19820_not
g82251 not n34652 ; n34652_not
g82252 not n34832 ; n34832_not
g82253 not n30449 ; n30449_not
g82254 not n21719 ; n21719_not
g82255 not n21728 ; n21728_not
g82256 not n53156 ; n53156_not
g82257 not n21737 ; n21737_not
g82258 not n21746 ; n21746_not
g82259 not n34913 ; n34913_not
g82260 not n21755 ; n21755_not
g82261 not n53165 ; n53165_not
g82262 not n21764 ; n21764_not
g82263 not n21395 ; n21395_not
g82264 not n21773 ; n21773_not
g82265 not n34931 ; n34931_not
g82266 not n57323 ; n57323_not
g82267 not n53174 ; n53174_not
g82268 not n21485 ; n21485_not
g82269 not n21629 ; n21629_not
g82270 not n53318 ; n53318_not
g82271 not n36128 ; n36128_not
g82272 not n21638 ; n21638_not
g82273 not n21647 ; n21647_not
g82274 not n52139 ; n52139_not
g82275 not n34526 ; n34526_not
g82276 not n21656 ; n21656_not
g82277 not n21458 ; n21458_not
g82278 not n21665 ; n21665_not
g82279 not n53129 ; n53129_not
g82280 not n21449 ; n21449_not
g82281 not n34904 ; n34904_not
g82282 not n21674 ; n21674_not
g82283 not n21683 ; n21683_not
g82284 not n21692 ; n21692_not
g82285 not n53138 ; n53138_not
g82286 not n53147 ; n53147_not
g82287 not n21854 ; n21854_not
g82288 not n21863 ; n21863_not
g82289 not n21872 ; n21872_not
g82290 not n49016 ; n49016_not
g82291 not n21881 ; n21881_not
g82292 not n21890 ; n21890_not
g82293 not n53219 ; n53219_not
g82294 not n44651 ; n44651_not
g82295 not n21908 ; n21908_not
g82296 not n53228 ; n53228_not
g82297 not n21917 ; n21917_not
g82298 not n30098 ; n30098_not
g82299 not n21926 ; n21926_not
g82300 not n21935 ; n21935_not
g82301 not n39521 ; n39521_not
g82302 not n21944 ; n21944_not
g82303 not n21782 ; n21782_not
g82304 not n47225 ; n47225_not
g82305 not n40655 ; n40655_not
g82306 not n21791 ; n21791_not
g82307 not n46460 ; n46460_not
g82308 not n52148 ; n52148_not
g82309 not n53183 ; n53183_not
g82310 not n21809 ; n21809_not
g82311 not n21818 ; n21818_not
g82312 not n53192 ; n53192_not
g82313 not n21368 ; n21368_not
g82314 not n21827 ; n21827_not
g82315 not n21359 ; n21359_not
g82316 not n21836 ; n21836_not
g82317 not n21845 ; n21845_not
g82318 not n53273 ; n53273_not
g82319 not n30287 ; n30287_not
g82320 not n11990 ; n11990_not
g82321 not n53363 ; n53363_not
g82322 not n20558 ; n20558_not
g82323 not n11981 ; n11981_not
g82324 not n53408 ; n53408_not
g82325 not n27047 ; n27047_not
g82326 not n57350 ; n57350_not
g82327 not n34535 ; n34535_not
g82328 not n20648 ; n20648_not
g82329 not n49043 ; n49043_not
g82330 not n36308 ; n36308_not
g82331 not n46307 ; n46307_not
g82332 not n53390 ; n53390_not
g82333 not n53381 ; n53381_not
g82334 not n56081 ; n56081_not
g82335 not n41285 ; n41285_not
g82336 not n21494 ; n21494_not
g82337 not n56072 ; n56072_not
g82338 not n30197 ; n30197_not
g82339 not n21539 ; n21539_not
g82340 not n57332 ; n57332_not
g82341 not n21548 ; n21548_not
g82342 not n21557 ; n21557_not
g82343 not n21566 ; n21566_not
g82344 not n53093 ; n53093_not
g82345 not n30188 ; n30188_not
g82346 not n21575 ; n21575_not
g82347 not n21584 ; n21584_not
g82348 not n49025 ; n49025_not
g82349 not n21593 ; n21593_not
g82350 not n30179 ; n30179_not
g82351 not n21269 ; n21269_not
g82352 not n21287 ; n21287_not
g82353 not n49034 ; n49034_not
g82354 not n30089 ; n30089_not
g82355 not n21377 ; n21377_not
g82356 not n27029 ; n27029_not
g82357 not n56162 ; n56162_not
g82358 not n44822 ; n44822_not
g82359 not n34922 ; n34922_not
g82360 not n21467 ; n21467_not
g82361 not n30548 ; n30548_not
g82362 not n12494 ; n12494_not
g82363 not n27182 ; n27182_not
g82364 not n44507 ; n44507_not
g82365 not n36236 ; n36236_not
g82366 not n30683 ; n30683_not
g82367 not n56180 ; n56180_not
g82368 not n36209 ; n36209_not
g82369 not n12467 ; n12467_not
g82370 not n46370 ; n46370_not
g82371 not n56090 ; n56090_not
g82372 not n27191 ; n27191_not
g82373 not n36263 ; n36263_not
g82374 not n41366 ; n41366_not
g82375 not n53444 ; n53444_not
g82376 not n12458 ; n12458_not
g82377 not n39053 ; n39053_not
g82378 not n12485 ; n12485_not
g82379 not n56171 ; n56171_not
g82380 not n37136 ; n37136_not
g82381 not n52067 ; n52067_not
g82382 not n36227 ; n36227_not
g82383 not n12476 ; n12476_not
g82384 not n56135 ; n56135_not
g82385 not n27155 ; n27155_not
g82386 not n36245 ; n36245_not
g82387 not n36182 ; n36182_not
g82388 not n56126 ; n56126_not
g82389 not n30755 ; n30755_not
g82390 not n52058 ; n52058_not
g82391 not n37145 ; n37145_not
g82392 not n12566 ; n12566_not
g82393 not n52049 ; n52049_not
g82394 not n34409 ; n34409_not
g82395 not n36254 ; n36254_not
g82396 not n19802 ; n19802_not
g82397 not n57404 ; n57404_not
g82398 not n12278 ; n12278_not
g82399 not n12269 ; n12269_not
g82400 not n46352 ; n46352_not
g82401 not n51851 ; n51851_not
g82402 not n36281 ; n36281_not
g82403 not n46415 ; n46415_not
g82404 not n56225 ; n56225_not
g82405 not n12287 ; n12287_not
g82406 not n52085 ; n52085_not
g82407 not n34724 ; n34724_not
g82408 not n46343 ; n46343_not
g82409 not n27164 ; n27164_not
g82410 not n34715 ; n34715_not
g82411 not n12197 ; n12197_not
g82412 not n39008 ; n39008_not
g82413 not n36191 ; n36191_not
g82414 not n30359 ; n30359_not
g82415 not n49403 ; n49403_not
g82416 not n12395 ; n12395_not
g82417 not n44831 ; n44831_not
g82418 not n12386 ; n12386_not
g82419 not n40970 ; n40970_not
g82420 not n56207 ; n56207_not
g82421 not n52076 ; n52076_not
g82422 not n12377 ; n12377_not
g82423 not n40961 ; n40961_not
g82424 not n56108 ; n56108_not
g82425 not n12449 ; n12449_not
g82426 not n45155 ; n45155_not
g82427 not n36218 ; n36218_not
g82428 not n34760 ; n34760_not
g82429 not n44705 ; n44705_not
g82430 not n37118 ; n37118_not
g82431 not n27209 ; n27209_not
g82432 not n36272 ; n36272_not
g82433 not n12296 ; n12296_not
g82434 not n12368 ; n12368_not
g82435 not n12359 ; n12359_not
g82436 not n46361 ; n46361_not
g82437 not n57422 ; n57422_not
g82438 not n56216 ; n56216_not
g82439 not n22826 ; n22826_not
g82440 not n51941 ; n51941_not
g82441 not n29801 ; n29801_not
g82442 not n57251 ; n57251_not
g82443 not n11558 ; n11558_not
g82444 not n46244 ; n46244_not
g82445 not n29810 ; n29810_not
g82446 not n50951 ; n50951_not
g82447 not n36344 ; n36344_not
g82448 not n26075 ; n26075_not
g82449 not n29603 ; n29603_not
g82450 not n57233 ; n57233_not
g82451 not n22943 ; n22943_not
g82452 not n22934 ; n22934_not
g82453 not n36056 ; n36056_not
g82454 not n40745 ; n40745_not
g82455 not n46235 ; n46235_not
g82456 not n22916 ; n22916_not
g82457 not n44633 ; n44633_not
g82458 not n11567 ; n11567_not
g82459 not n22871 ; n22871_not
g82460 not n11576 ; n11576_not
g82461 not n46505 ; n46505_not
g82462 not n49520 ; n49520_not
g82463 not n57242 ; n57242_not
g82464 not n47180 ; n47180_not
g82465 not n49610 ; n49610_not
g82466 not n22187 ; n22187_not
g82467 not n36335 ; n36335_not
g82468 not n26912 ; n26912_not
g82469 not n36137 ; n36137_not
g82470 not n46262 ; n46262_not
g82471 not n22196 ; n22196_not
g82472 not n29900 ; n29900_not
g82473 not n44642 ; n44642_not
g82474 not n11486 ; n11486_not
g82475 not n11477 ; n11477_not
g82476 not n52184 ; n52184_not
g82477 not n51950 ; n51950_not
g82478 not n22097 ; n22097_not
g82479 not n52193 ; n52193_not
g82480 not n51761 ; n51761_not
g82481 not n46253 ; n46253_not
g82482 not n49601 ; n49601_not
g82483 not n50906 ; n50906_not
g82484 not n57260 ; n57260_not
g82485 not n38054 ; n38054_not
g82486 not n22952 ; n22952_not
g82487 not n57206 ; n57206_not
g82488 not n36920 ; n36920_not
g82489 not n11495 ; n11495_not
g82490 not n52229 ; n52229_not
g82491 not n29612 ; n29612_not
g82492 not n44723 ; n44723_not
g82493 not n29522 ; n29522_not
g82494 not n44813 ; n44813_not
g82495 not n44552 ; n44552_not
g82496 not n11468 ; n11468_not
g82497 not n46208 ; n46208_not
g82498 not n29540 ; n29540_not
g82499 not n44615 ; n44615_not
g82500 not n52238 ; n52238_not
g82501 not n49502 ; n49502_not
g82502 not n23069 ; n23069_not
g82503 not n29630 ; n29630_not
g82504 not n39611 ; n39611_not
g82505 not n23078 ; n23078_not
g82506 not n51932 ; n51932_not
g82507 not n22961 ; n22961_not
g82508 not n52481 ; n52481_not
g82509 not n44624 ; n44624_not
g82510 not n46226 ; n46226_not
g82511 not n47135 ; n47135_not
g82512 not n51086 ; n51086_not
g82513 not n46217 ; n46217_not
g82514 not n34823 ; n34823_not
g82515 not n38009 ; n38009_not
g82516 not n29531 ; n29531_not
g82517 not n11585 ; n11585_not
g82518 not n51923 ; n51923_not
g82519 not n49007 ; n49007_not
g82520 not n49700 ; n49700_not
g82521 not n52166 ; n52166_not
g82522 not n43742 ; n43742_not
g82523 not n44714 ; n44714_not
g82524 not n22079 ; n22079_not
g82525 not n36317 ; n36317_not
g82526 not n22277 ; n22277_not
g82527 not n46271 ; n46271_not
g82528 not n57314 ; n57314_not
g82529 not n22286 ; n22286_not
g82530 not n22295 ; n22295_not
g82531 not n46280 ; n46280_not
g82532 not n57305 ; n57305_not
g82533 not n22259 ; n22259_not
g82534 not n50825 ; n50825_not
g82535 not n52436 ; n52436_not
g82536 not n52175 ; n52175_not
g82537 not n37028 ; n37028_not
g82538 not n22169 ; n22169_not
g82539 not n21953 ; n21953_not
g82540 not n36326 ; n36326_not
g82541 not n21962 ; n21962_not
g82542 not n21971 ; n21971_not
g82543 not n21980 ; n21980_not
g82544 not n21278 ; n21278_not
g82545 not n52157 ; n52157_not
g82546 not n50861 ; n50861_not
g82547 not n57450 ; n57450_not
g82548 not n37407 ; n37407_not
g82549 not n35814 ; n35814_not
g82550 not n56622 ; n56622_not
g82551 not n36219 ; n36219_not
g82552 not n56127 ; n56127_not
g82553 not n57036 ; n57036_not
g82554 not n35508 ; n35508_not
g82555 not n56325 ; n56325_not
g82556 not n56442 ; n56442_not
g82557 not n14826 ; n14826_not
g82558 not n36084 ; n36084_not
g82559 not n56361 ; n56361_not
g82560 not n14727 ; n14727_not
g82561 not n14835 ; n14835_not
g82562 not n43626 ; n43626_not
g82563 not n56190 ; n56190_not
g82564 not n14772 ; n14772_not
g82565 not n56406 ; n56406_not
g82566 not n14196 ; n14196_not
g82567 not n56136 ; n56136_not
g82568 not n57441 ; n57441_not
g82569 not n33159 ; n33159_not
g82570 not n35382 ; n35382_not
g82571 not n33168 ; n33168_not
g82572 not n56334 ; n56334_not
g82573 not n43167 ; n43167_not
g82574 not n44580 ; n44580_not
g82575 not n35580 ; n35580_not
g82576 not n35904 ; n35904_not
g82577 not n35517 ; n35517_not
g82578 not n36507 ; n36507_not
g82579 not n36318 ; n36318_not
g82580 not n44571 ; n44571_not
g82581 not n33339 ; n33339_not
g82582 not n14736 ; n14736_not
g82583 not n36264 ; n36264_not
g82584 not n36246 ; n36246_not
g82585 not n37371 ; n37371_not
g82586 not n14745 ; n14745_not
g82587 not n14790 ; n14790_not
g82588 not n44742 ; n44742_not
g82589 not n57180 ; n57180_not
g82590 not n14187 ; n14187_not
g82591 not n56532 ; n56532_not
g82592 not n43482 ; n43482_not
g82593 not n57162 ; n57162_not
g82594 not n14655 ; n14655_not
g82595 not n15069 ; n15069_not
g82596 not n56631 ; n56631_not
g82597 not n35616 ; n35616_not
g82598 not n57054 ; n57054_not
g82599 not n33348 ; n33348_not
g82600 not n44940 ; n44940_not
g82601 not n14844 ; n14844_not
g82602 not n37146 ; n37146_not
g82603 not n14709 ; n14709_not
g82604 not n48261 ; n48261_not
g82605 not n48162 ; n48162_not
g82606 not n44607 ; n44607_not
g82607 not n44085 ; n44085_not
g82608 not n56217 ; n56217_not
g82609 not n56721 ; n56721_not
g82610 not n56901 ; n56901_not
g82611 not n14781 ; n14781_not
g82612 not n33609 ; n33609_not
g82613 not n48801 ; n48801_not
g82614 not n36048 ; n36048_not
g82615 not n35832 ; n35832_not
g82616 not n56820 ; n56820_not
g82617 not n56316 ; n56316_not
g82618 not n44922 ; n44922_not
g82619 not n44553 ; n44553_not
g82620 not n57324 ; n57324_not
g82621 not n43545 ; n43545_not
g82622 not n35373 ; n35373_not
g82623 not n44508 ; n44508_not
g82624 not n56541 ; n56541_not
g82625 not n35733 ; n35733_not
g82626 not n48126 ; n48126_not
g82627 not n56208 ; n56208_not
g82628 not n43563 ; n43563_not
g82629 not n35922 ; n35922_not
g82630 not n35805 ; n35805_not
g82631 not n14718 ; n14718_not
g82632 not n50349 ; n50349_not
g82633 not n43923 ; n43923_not
g82634 not n57225 ; n57225_not
g82635 not n36129 ; n36129_not
g82636 not n48081 ; n48081_not
g82637 not n56307 ; n56307_not
g82638 not n43941 ; n43941_not
g82639 not n36237 ; n36237_not
g82640 not n35931 ; n35931_not
g82641 not n48153 ; n48153_not
g82642 not n14808 ; n14808_not
g82643 not n56352 ; n56352_not
g82644 not n48225 ; n48225_not
g82645 not n36516 ; n36516_not
g82646 not n43635 ; n43635_not
g82647 not n14754 ; n14754_not
g82648 not n14169 ; n14169_not
g82649 not n36192 ; n36192_not
g82650 not n36183 ; n36183_not
g82651 not n14763 ; n14763_not
g82652 not n48072 ; n48072_not
g82653 not n57153 ; n57153_not
g82654 not n43950 ; n43950_not
g82655 not n56523 ; n56523_not
g82656 not n36426 ; n36426_not
g82657 not n48603 ; n48603_not
g82658 not n56163 ; n56163_not
g82659 not n56370 ; n56370_not
g82660 not n56460 ; n56460_not
g82661 not n43077 ; n43077_not
g82662 not n43527 ; n43527_not
g82663 not n56514 ; n56514_not
g82664 not n43473 ; n43473_not
g82665 not n48216 ; n48216_not
g82666 not n35913 ; n35913_not
g82667 not n37425 ; n37425_not
g82668 not n56145 ; n56145_not
g82669 not n33627 ; n33627_not
g82670 not n35742 ; n35742_not
g82671 not n33375 ; n33375_not
g82672 not n56811 ; n56811_not
g82673 not n35607 ; n35607_not
g82674 not n56640 ; n56640_not
g82675 not n56154 ; n56154_not
g82676 not n48720 ; n48720_not
g82677 not n35391 ; n35391_not
g82678 not n44616 ; n44616_not
g82679 not n36354 ; n36354_not
g82680 not n44058 ; n44058_not
g82681 not n56181 ; n56181_not
g82682 not n36228 ; n36228_not
g82683 not n14637 ; n14637_not
g82684 not n36417 ; n36417_not
g82685 not n14817 ; n14817_not
g82686 not n57315 ; n57315_not
g82687 not n36147 ; n36147_not
g82688 not n43572 ; n43572_not
g82689 not n33294 ; n33294_not
g82690 not n56343 ; n56343_not
g82691 not n36174 ; n36174_not
g82692 not n44076 ; n44076_not
g82693 not n14646 ; n14646_not
g82694 not n44544 ; n44544_not
g82695 not n36435 ; n36435_not
g82696 not n48702 ; n48702_not
g82697 not n33636 ; n33636_not
g82698 not n35823 ; n35823_not
g82699 not n14178 ; n14178_not
g82700 not n56172 ; n56172_not
g82701 not n15087 ; n15087_not
g82702 not n45066 ; n45066_not
g82703 not n56505 ; n56505_not
g82704 not n56451 ; n56451_not
g82705 not n43554 ; n43554_not
g82706 not n48711 ; n48711_not
g82707 not n57171 ; n57171_not
g82708 not n44751 ; n44751_not
g82709 not n36255 ; n36255_not
g82710 not n35751 ; n35751_not
g82711 not n36039 ; n36039_not
g82712 not n35490 ; n35490_not
g82713 not n36363 ; n36363_not
g82714 not n48270 ; n48270_not
g82715 not n14943 ; n14943_not
g82716 not n33384 ; n33384_not
g82717 not n57270 ; n57270_not
g82718 not n14907 ; n14907_not
g82719 not n44715 ; n44715_not
g82720 not n48135 ; n48135_not
g82721 not n56730 ; n56730_not
g82722 not n56226 ; n56226_not
g82723 not n56604 ; n56604_not
g82724 not n56235 ; n56235_not
g82725 not n36381 ; n36381_not
g82726 not n35535 ; n35535_not
g82727 not n35661 ; n35661_not
g82728 not n15168 ; n15168_not
g82729 not n56271 ; n56271_not
g82730 not n36336 ; n36336_not
g82731 not n14277 ; n14277_not
g82732 not n14691 ; n14691_not
g82733 not n14619 ; n14619_not
g82734 not n14673 ; n14673_not
g82735 not n44067 ; n44067_not
g82736 not n48243 ; n48243_not
g82737 not n44931 ; n44931_not
g82738 not n33078 ; n33078_not
g82739 not n14628 ; n14628_not
g82740 not n37380 ; n37380_not
g82741 not n44049 ; n44049_not
g82742 not n15177 ; n15177_not
g82743 not n55065 ; n55065_not
g82744 not n35940 ; n35940_not
g82745 not n56262 ; n56262_not
g82746 not n36291 ; n36291_not
g82747 not n33087 ; n33087_not
g82748 not n57342 ; n57342_not
g82749 not n48144 ; n48144_not
g82750 not n35436 ; n35436_not
g82751 not n55038 ; n55038_not
g82752 not n43932 ; n43932_not
g82753 not n14268 ; n14268_not
g82754 not n43536 ; n43536_not
g82755 not n45057 ; n45057_not
g82756 not n36057 ; n36057_not
g82757 not n35553 ; n35553_not
g82758 not n14925 ; n14925_not
g82759 not n44733 ; n44733_not
g82760 not n37434 ; n37434_not
g82761 not n57081 ; n57081_not
g82762 not n55074 ; n55074_not
g82763 not n35850 ; n35850_not
g82764 not n15159 ; n15159_not
g82765 not n48180 ; n48180_not
g82766 not n56910 ; n56910_not
g82767 not n15195 ; n15195_not
g82768 not n36390 ; n36390_not
g82769 not n14295 ; n14295_not
g82770 not n14934 ; n14934_not
g82771 not n44661 ; n44661_not
g82772 not n45039 ; n45039_not
g82773 not n36327 ; n36327_not
g82774 not n14376 ; n14376_not
g82775 not n48117 ; n48117_not
g82776 not n36093 ; n36093_not
g82777 not n35454 ; n35454_not
g82778 not n14682 ; n14682_not
g82779 not n36156 ; n36156_not
g82780 not n56280 ; n56280_not
g82781 not n35706 ; n35706_not
g82782 not n36462 ; n36462_not
g82783 not n33069 ; n33069_not
g82784 not n35652 ; n35652_not
g82785 not n14385 ; n14385_not
g82786 not n44643 ; n44643_not
g82787 not n35841 ; n35841_not
g82788 not n36138 ; n36138_not
g82789 not n43518 ; n43518_not
g82790 not n35463 ; n35463_not
g82791 not n14916 ; n14916_not
g82792 not n36471 ; n36471_not
g82793 not n48108 ; n48108_not
g82794 not n35544 ; n35544_not
g82795 not n57090 ; n57090_not
g82796 not n14286 ; n14286_not
g82797 not n35445 ; n35445_not
g82798 not n44706 ; n44706_not
g82799 not n43590 ; n43590_not
g82800 not n44517 ; n44517_not
g82801 not n57243 ; n57243_not
g82802 not n14853 ; n14853_not
g82803 not n48090 ; n48090_not
g82804 not n57126 ; n57126_not
g82805 not n56550 ; n56550_not
g82806 not n57027 ; n57027_not
g82807 not n14970 ; n14970_not
g82808 not n56424 ; n56424_not
g82809 not n56415 ; n56415_not
g82810 not n36282 ; n36282_not
g82811 not n44652 ; n44652_not
g82812 not n14862 ; n14862_not
g82813 not n35643 ; n35643_not
g82814 not n14961 ; n14961_not
g82815 not n48234 ; n48234_not
g82816 not n43581 ; n43581_not
g82817 not n55083 ; n55083_not
g82818 not n48207 ; n48207_not
g82819 not n57018 ; n57018_not
g82820 not n48612 ; n48612_not
g82821 not n35418 ; n35418_not
g82822 not n35571 ; n35571_not
g82823 not n57234 ; n57234_not
g82824 not n36444 ; n36444_not
g82825 not n43509 ; n43509_not
g82826 not n36408 ; n36408_not
g82827 not n57306 ; n57306_not
g82828 not n35409 ; n35409_not
g82829 not n56433 ; n56433_not
g82830 not n44724 ; n44724_not
g82831 not n48252 ; n48252_not
g82832 not n44625 ; n44625_not
g82833 not n43617 ; n43617_not
g82834 not n36273 ; n36273_not
g82835 not n57414 ; n57414_not
g82836 not n35481 ; n35481_not
g82837 not n37416 ; n37416_not
g82838 not n55029 ; n55029_not
g82839 not n14664 ; n14664_not
g82840 not n56244 ; n56244_not
g82841 not n36453 ; n36453_not
g82842 not n33258 ; n33258_not
g82843 not n14259 ; n14259_not
g82844 not n48009 ; n48009_not
g82845 not n33096 ; n33096_not
g82846 not n14871 ; n14871_not
g82847 not n57252 ; n57252_not
g82848 not n43095 ; n43095_not
g82849 not n44670 ; n44670_not
g82850 not n48171 ; n48171_not
g82851 not n50358 ; n50358_not
g82852 not n36480 ; n36480_not
g82853 not n57009 ; n57009_not
g82854 not n36309 ; n36309_not
g82855 not n14880 ; n14880_not
g82856 not n43491 ; n43491_not
g82857 not n57108 ; n57108_not
g82858 not n44634 ; n44634_not
g82859 not n48621 ; n48621_not
g82860 not n44562 ; n44562_not
g82861 not n33285 ; n33285_not
g82862 not n35562 ; n35562_not
g82863 not n33357 ; n33357_not
g82864 not n36372 ; n36372_not
g82865 not n35526 ; n35526_not
g82866 not n56253 ; n56253_not
g82867 not n36066 ; n36066_not
g82868 not n43086 ; n43086_not
g82869 not n56613 ; n56613_not
g82870 not n35427 ; n35427_not
g82871 not n43608 ; n43608_not
g82872 not n14952 ; n14952_not
g82873 not n35472 ; n35472_not
g82874 not n14367 ; n14367_not
g82875 not n36345 ; n36345_not
g82876 not n33942 ; n33942_not
g82877 not n13485 ; n13485_not
g82878 not n11784 ; n11784_not
g82879 not n13476 ; n13476_not
g82880 not n13278 ; n13278_not
g82881 not n44247 ; n44247_not
g82882 not n13467 ; n13467_not
g82883 not n33951 ; n33951_not
g82884 not n11793 ; n11793_not
g82885 not n37218 ; n37218_not
g82886 not n34860 ; n34860_not
g82887 not n11829 ; n11829_not
g82888 not n49602 ; n49602_not
g82889 not n44814 ; n44814_not
g82890 not n13458 ; n13458_not
g82891 not n13287 ; n13287_not
g82892 not n11496 ; n11496_not
g82893 not n49611 ; n49611_not
g82894 not n11838 ; n11838_not
g82895 not n44238 ; n44238_not
g82896 not n49620 ; n49620_not
g82897 not n13449 ; n13449_not
g82898 not n13296 ; n13296_not
g82899 not n33960 ; n33960_not
g82900 not n11577 ; n11577_not
g82901 not n11685 ; n11685_not
g82902 not n13548 ; n13548_not
g82903 not n33915 ; n33915_not
g82904 not n11694 ; n11694_not
g82905 not n11568 ; n11568_not
g82906 not n34284 ; n34284_not
g82907 not n13539 ; n13539_not
g82908 not n44256 ; n44256_not
g82909 not n33924 ; n33924_not
g82910 not n49530 ; n49530_not
g82911 not n44229 ; n44229_not
g82912 not n34293 ; n34293_not
g82913 not n11739 ; n11739_not
g82914 not n33933 ; n33933_not
g82915 not n11748 ; n11748_not
g82916 not n11757 ; n11757_not
g82917 not n13494 ; n13494_not
g82918 not n11766 ; n11766_not
g82919 not n11775 ; n11775_not
g82920 not n12783 ; n12783_not
g82921 not n43842 ; n43842_not
g82922 not n34356 ; n34356_not
g82923 not n49710 ; n49710_not
g82924 not n11892 ; n11892_not
g82925 not n34365 ; n34365_not
g82926 not n43833 ; n43833_not
g82927 not n34374 ; n34374_not
g82928 not n37209 ; n37209_not
g82929 not n11919 ; n11919_not
g82930 not n34383 ; n34383_not
g82931 not n11928 ; n11928_not
g82932 not n37038 ; n37038_not
g82933 not n11937 ; n11937_not
g82934 not n44409 ; n44409_not
g82935 not n11946 ; n11946_not
g82936 not n11487 ; n11487_not
g82937 not n11847 ; n11847_not
g82938 not n11856 ; n11856_not
g82939 not n34329 ; n34329_not
g82940 not n11478 ; n11478_not
g82941 not n11865 ; n11865_not
g82942 not n43734 ; n43734_not
g82943 not n11874 ; n11874_not
g82944 not n49701 ; n49701_not
g82945 not n12774 ; n12774_not
g82946 not n13359 ; n13359_not
g82947 not n34347 ; n34347_not
g82948 not n11883 ; n11883_not
g82949 not n13368 ; n13368_not
g82950 not n13377 ; n13377_not
g82951 not n13386 ; n13386_not
g82952 not n49503 ; n49503_not
g82953 not n13395 ; n13395_not
g82954 not n34338 ; n34338_not
g82955 not n11379 ; n11379_not
g82956 not n34086 ; n34086_not
g82957 not n10884 ; n10884_not
g82958 not n56037 ; n56037_not
g82959 not n13683 ; n13683_not
g82960 not n11388 ; n11388_not
g82961 not n49440 ; n49440_not
g82962 not n33843 ; n33843_not
g82963 not n34077 ; n34077_not
g82964 not n11397 ; n11397_not
g82965 not n44265 ; n44265_not
g82966 not n13674 ; n13674_not
g82967 not n13665 ; n13665_not
g82968 not n33852 ; n33852_not
g82969 not n10875 ; n10875_not
g82970 not n13656 ; n13656_not
g82971 not n55920 ; n55920_not
g82972 not n44373 ; n44373_not
g82973 not n33861 ; n33861_not
g82974 not n13647 ; n13647_not
g82975 not n49422 ; n49422_not
g82976 not n34176 ; n34176_not
g82977 not n13746 ; n13746_not
g82978 not n11289 ; n11289_not
g82979 not n48306 ; n48306_not
g82980 not n33816 ; n33816_not
g82981 not n10938 ; n10938_not
g82982 not n37245 ; n37245_not
g82983 not n11298 ; n11298_not
g82984 not n10929 ; n10929_not
g82985 not n10893 ; n10893_not
g82986 not n37236 ; n37236_not
g82987 not n13692 ; n13692_not
g82988 not n33834 ; n33834_not
g82989 not n44283 ; n44283_not
g82990 not n55902 ; n55902_not
g82991 not n34194 ; n34194_not
g82992 not n13719 ; n13719_not
g82993 not n33825 ; n33825_not
g82994 not n13728 ; n13728_not
g82995 not n44274 ; n44274_not
g82996 not n36912 ; n36912_not
g82997 not n13737 ; n13737_not
g82998 not n43707 ; n43707_not
g82999 not n34185 ; n34185_not
g83000 not n13584 ; n13584_not
g83001 not n34257 ; n34257_not
g83002 not n44148 ; n44148_not
g83003 not n34824 ; n34824_not
g83004 not n13575 ; n13575_not
g83005 not n11649 ; n11649_not
g83006 not n49512 ; n49512_not
g83007 not n11658 ; n11658_not
g83008 not n56046 ; n56046_not
g83009 not n34833 ; n34833_not
g83010 not n34266 ; n34266_not
g83011 not n11667 ; n11667_not
g83012 not n37227 ; n37227_not
g83013 not n13566 ; n13566_not
g83014 not n11586 ; n11586_not
g83015 not n33906 ; n33906_not
g83016 not n44904 ; n44904_not
g83017 not n11676 ; n11676_not
g83018 not n13557 ; n13557_not
g83019 not n34275 ; n34275_not
g83020 not n34068 ; n34068_not
g83021 not n13638 ; n13638_not
g83022 not n36534 ; n36534_not
g83023 not n13188 ; n13188_not
g83024 not n33870 ; n33870_not
g83025 not n13629 ; n13629_not
g83026 not n34239 ; n34239_not
g83027 not n36921 ; n36921_not
g83028 not n11595 ; n11595_not
g83029 not n44913 ; n44913_not
g83030 not n13593 ; n13593_not
g83031 not n34815 ; n34815_not
g83032 not n34248 ; n34248_not
g83033 not n36930 ; n36930_not
g83034 not n44382 ; n44382_not
g83035 not n11199 ; n11199_not
g83036 not n13197 ; n13197_not
g83037 not n12765 ; n12765_not
g83038 not n49323 ; n49323_not
g83039 not n34752 ; n34752_not
g83040 not n34581 ; n34581_not
g83041 not n56109 ; n56109_not
g83042 not n12369 ; n12369_not
g83043 not n34743 ; n34743_not
g83044 not n12378 ; n12378_not
g83045 not n37128 ; n37128_not
g83046 not n34590 ; n34590_not
g83047 not n37173 ; n37173_not
g83048 not n12387 ; n12387_not
g83049 not n44166 ; n44166_not
g83050 not n12396 ; n12396_not
g83051 not n34734 ; n34734_not
g83052 not n44184 ; n44184_not
g83053 not n34464 ; n34464_not
g83054 not n12729 ; n12729_not
g83055 not n34725 ; n34725_not
g83056 not n34455 ; n34455_not
g83057 not n44418 ; n44418_not
g83058 not n12459 ; n12459_not
g83059 not n37119 ; n37119_not
g83060 not n12693 ; n12693_not
g83061 not n34554 ; n34554_not
g83062 not n44850 ; n44850_not
g83063 not n12279 ; n12279_not
g83064 not n49314 ; n49314_not
g83065 not n34563 ; n34563_not
g83066 not n34770 ; n34770_not
g83067 not n48027 ; n48027_not
g83068 not n12288 ; n12288_not
g83069 not n37182 ; n37182_not
g83070 not n12297 ; n12297_not
g83071 not n34572 ; n34572_not
g83072 not n34761 ; n34761_not
g83073 not n56055 ; n56055_not
g83074 not n12756 ; n12756_not
g83075 not n34635 ; n34635_not
g83076 not n56073 ; n56073_not
g83077 not n12549 ; n12549_not
g83078 not n12558 ; n12558_not
g83079 not n44427 ; n44427_not
g83080 not n12738 ; n12738_not
g83081 not n34644 ; n34644_not
g83082 not n12576 ; n12576_not
g83083 not n44157 ; n44157_not
g83084 not n34680 ; n34680_not
g83085 not n12684 ; n12684_not
g83086 not n34653 ; n34653_not
g83087 not n34419 ; n34419_not
g83088 not n12594 ; n12594_not
g83089 not n44175 ; n44175_not
g83090 not n37155 ; n37155_not
g83091 not n34662 ; n34662_not
g83092 not n12666 ; n12666_not
g83093 not n49350 ; n49350_not
g83094 not n34671 ; n34671_not
g83095 not n12639 ; n12639_not
g83096 not n12648 ; n12648_not
g83097 not n34608 ; n34608_not
g83098 not n12468 ; n12468_not
g83099 not n44832 ; n44832_not
g83100 not n34716 ; n34716_not
g83101 not n34617 ; n34617_not
g83102 not n12477 ; n12477_not
g83103 not n44139 ; n44139_not
g83104 not n12486 ; n12486_not
g83105 not n11991 ; n11991_not
g83106 not n37164 ; n37164_not
g83107 not n56082 ; n56082_not
g83108 not n12747 ; n12747_not
g83109 not n44841 ; n44841_not
g83110 not n34626 ; n34626_not
g83111 not n34707 ; n34707_not
g83112 not n12495 ; n12495_not
g83113 not n34446 ; n34446_not
g83114 not n34518 ; n34518_not
g83115 not n37056 ; n37056_not
g83116 not n34527 ; n34527_not
g83117 not n43752 ; n43752_not
g83118 not n34536 ; n34536_not
g83119 not n34545 ; n34545_not
g83120 not n37065 ; n37065_not
g83121 not n34473 ; n34473_not
g83122 not n44823 ; n44823_not
g83123 not n49800 ; n49800_not
g83124 not n43824 ; n43824_not
g83125 not n11955 ; n11955_not
g83126 not n34932 ; n34932_not
g83127 not n34905 ; n34905_not
g83128 not n49305 ; n49305_not
g83129 not n43743 ; n43743_not
g83130 not n34923 ; n34923_not
g83131 not n11964 ; n11964_not
g83132 not n34428 ; n34428_not
g83133 not n12567 ; n12567_not
g83134 not n48018 ; n48018_not
g83135 not n49413 ; n49413_not
g83136 not n37191 ; n37191_not
g83137 not n12189 ; n12189_not
g83138 not n12198 ; n12198_not
g83139 not n49404 ; n49404_not
g83140 not n56091 ; n56091_not
g83141 not n34491 ; n34491_not
g83142 not n44193 ; n44193_not
g83143 not n56028 ; n56028_not
g83144 not n44094 ; n44094_not
g83145 not n37083 ; n37083_not
g83146 not n34509 ; n34509_not
g83147 not n12657 ; n12657_not
g83148 not n34842 ; n34842_not
g83149 not n44454 ; n44454_not
g83150 not n33807 ; n33807_not
g83151 not n36714 ; n36714_not
g83152 not n14466 ; n14466_not
g83153 not n48531 ; n48531_not
g83154 not n14457 ; n14457_not
g83155 not n47802 ; n47802_not
g83156 not n36723 ; n36723_not
g83157 not n48522 ; n48522_not
g83158 not n35193 ; n35193_not
g83159 not n36642 ; n36642_not
g83160 not n36732 ; n36732_not
g83161 not n43761 ; n43761_not
g83162 not n44436 ; n44436_not
g83163 not n48513 ; n48513_not
g83164 not n36633 ; n36633_not
g83165 not n14439 ; n14439_not
g83166 not n36741 ; n36741_not
g83167 not n33726 ; n33726_not
g83168 not n14556 ; n14556_not
g83169 not n14547 ; n14547_not
g83170 not n33780 ; n33780_not
g83171 not n35670 ; n35670_not
g83172 not n37335 ; n37335_not
g83173 not n50277 ; n50277_not
g83174 not n48441 ; n48441_not
g83175 not n14529 ; n14529_not
g83176 not n50268 ; n50268_not
g83177 not n48450 ; n48450_not
g83178 not n33717 ; n33717_not
g83179 not n48504 ; n48504_not
g83180 not n44481 ; n44481_not
g83181 not n44337 ; n44337_not
g83182 not n48540 ; n48540_not
g83183 not n36705 ; n36705_not
g83184 not n35625 ; n35625_not
g83185 not n14484 ; n14484_not
g83186 not n44463 ; n44463_not
g83187 not n35247 ; n35247_not
g83188 not n33681 ; n33681_not
g83189 not n37326 ; n37326_not
g83190 not n13962 ; n13962_not
g83191 not n35256 ; n35256_not
g83192 not n44364 ; n44364_not
g83193 not n10299 ; n10299_not
g83194 not n13755 ; n13755_not
g83195 not n55911 ; n55911_not
g83196 not n36750 ; n36750_not
g83197 not n36624 ; n36624_not
g83198 not n14394 ; n14394_not
g83199 not n14349 ; n14349_not
g83200 not n35238 ; n35238_not
g83201 not n33690 ; n33690_not
g83202 not n44391 ; n44391_not
g83203 not n35346 ; n35346_not
g83204 not n43653 ; n43653_not
g83205 not n14097 ; n14097_not
g83206 not n48342 ; n48342_not
g83207 not n33672 ; n33672_not
g83208 not n14088 ; n14088_not
g83209 not n48351 ; n48351_not
g83210 not n43662 ; n43662_not
g83211 not n48360 ; n48360_not
g83212 not n48630 ; n48630_not
g83213 not n14079 ; n14079_not
g83214 not n43671 ; n43671_not
g83215 not n37362 ; n37362_not
g83216 not n43680 ; n43680_not
g83217 not n48405 ; n48405_not
g83218 not n48315 ; n48315_not
g83219 not n36543 ; n36543_not
g83220 not n35364 ; n35364_not
g83221 not n48324 ; n48324_not
g83222 not n43644 ; n43644_not
g83223 not n35760 ; n35760_not
g83224 not n14475 ; n14475_not
g83225 not n35355 ; n35355_not
g83226 not n36561 ; n36561_not
g83227 not n44472 ; n44472_not
g83228 not n48333 ; n48333_not
g83229 not n33654 ; n33654_not
g83230 not n37353 ; n37353_not
g83231 not n43716 ; n43716_not
g83232 not n33744 ; n33744_not
g83233 not n13971 ; n13971_not
g83234 not n55803 ; n55803_not
g83235 not n48414 ; n48414_not
g83236 not n14583 ; n14583_not
g83237 not n33735 ; n33735_not
g83238 not n37029 ; n37029_not
g83239 not n50295 ; n50295_not
g83240 not n37344 ; n37344_not
g83241 not n48423 ; n48423_not
g83242 not n14565 ; n14565_not
g83243 not n55812 ; n55812_not
g83244 not n55821 ; n55821_not
g83245 not n36651 ; n36651_not
g83246 not n48432 ; n48432_not
g83247 not n44760 ; n44760_not
g83248 not n36606 ; n36606_not
g83249 not n44526 ; n44526_not
g83250 not n35715 ; n35715_not
g83251 not n56703 ; n56703_not
g83252 not n14592 ; n14592_not
g83253 not n13980 ; n13980_not
g83254 not n43374 ; n43374_not
g83255 not n55830 ; n55830_not
g83256 not n37281 ; n37281_not
g83257 not n50097 ; n50097_not
g83258 not n43365 ; n43365_not
g83259 not n50088 ; n50088_not
g83260 not n13953 ; n13953_not
g83261 not n43356 ; n43356_not
g83262 not n47343 ; n47343_not
g83263 not n13944 ; n13944_not
g83264 not n48063 ; n48063_not
g83265 not n43347 ; n43347_not
g83266 not n35292 ; n35292_not
g83267 not n13926 ; n13926_not
g83268 not n37272 ; n37272_not
g83269 not n35283 ; n35283_not
g83270 not n10947 ; n10947_not
g83271 not n44319 ; n44319_not
g83272 not n10866 ; n10866_not
g83273 not n13917 ; n13917_not
g83274 not n35328 ; n35328_not
g83275 not n35337 ; n35337_not
g83276 not n37290 ; n37290_not
g83277 not n43392 ; n43392_not
g83278 not n13935 ; n13935_not
g83279 not n43383 ; n43383_not
g83280 not n48054 ; n48054_not
g83281 not n43851 ; n43851_not
g83282 not n44805 ; n44805_not
g83283 not n43284 ; n43284_not
g83284 not n13809 ; n13809_not
g83285 not n34149 ; n34149_not
g83286 not n42672 ; n42672_not
g83287 not n13791 ; n13791_not
g83288 not n13782 ; n13782_not
g83289 not n10983 ; n10983_not
g83290 not n35184 ; n35184_not
g83291 not n34158 ; n34158_not
g83292 not n36552 ; n36552_not
g83293 not n10974 ; n10974_not
g83294 not n43914 ; n43914_not
g83295 not n44292 ; n44292_not
g83296 not n10965 ; n10965_not
g83297 not n13764 ; n13764_not
g83298 not n34167 ; n34167_not
g83299 not n36903 ; n36903_not
g83300 not n37074 ; n37074_not
g83301 not n34095 ; n34095_not
g83302 not n37263 ; n37263_not
g83303 not n43338 ; n43338_not
g83304 not n35265 ; n35265_not
g83305 not n43329 ; n43329_not
g83306 not n13881 ; n13881_not
g83307 not n13872 ; n13872_not
g83308 not n13827 ; n13827_not
g83309 not n13836 ; n13836_not
g83310 not n43293 ; n43293_not
g83311 not n37254 ; n37254_not
g83312 not n33771 ; n33771_not
g83313 not n13854 ; n13854_not
g83314 not n10992 ; n10992_not
g83315 not n50187 ; n50187_not
g83316 not n36822 ; n36822_not
g83317 not n44346 ; n44346_not
g83318 not n44328 ; n44328_not
g83319 not n43464 ; n43464_not
g83320 not n49332 ; n49332_not
g83321 not n43806 ; n43806_not
g83322 not n36831 ; n36831_not
g83323 not n10389 ; n10389_not
g83324 not n36804 ; n36804_not
g83325 not n10479 ; n10479_not
g83326 not n48036 ; n48036_not
g83327 not n10497 ; n10497_not
g83328 not n37317 ; n37317_not
g83329 not n36813 ; n36813_not
g83330 not n43437 ; n43437_not
g83331 not n43428 ; n43428_not
g83332 not n43419 ; n43419_not
g83333 not n13890 ; n13890_not
g83334 not n33645 ; n33645_not
g83335 not n50178 ; n50178_not
g83336 not n43455 ; n43455_not
g83337 not n37308 ; n37308_not
g83338 not n43446 ; n43446_not
g83339 not n13845 ; n13845_not
g83340 not n36840 ; n36840_not
g83341 not n38136 ; n38136_not
g83342 not n29802 ; n29802_not
g83343 not n22539 ; n22539_not
g83344 not n22548 ; n22548_not
g83345 not n22557 ; n22557_not
g83346 not n38055 ; n38055_not
g83347 not n22566 ; n22566_not
g83348 not n22575 ; n22575_not
g83349 not n47172 ; n47172_not
g83350 not n22584 ; n22584_not
g83351 not n47163 ; n47163_not
g83352 not n22593 ; n22593_not
g83353 not n50916 ; n50916_not
g83354 not n22629 ; n22629_not
g83355 not n22638 ; n22638_not
g83356 not n22647 ; n22647_not
g83357 not n22656 ; n22656_not
g83358 not n22665 ; n22665_not
g83359 not n38046 ; n38046_not
g83360 not n22674 ; n22674_not
g83361 not n50844 ; n50844_not
g83362 not n22368 ; n22368_not
g83363 not n50853 ; n50853_not
g83364 not n22377 ; n22377_not
g83365 not n52437 ; n52437_not
g83366 not n22386 ; n22386_not
g83367 not n22395 ; n22395_not
g83368 not n50871 ; n50871_not
g83369 not n22449 ; n22449_not
g83370 not n22458 ; n22458_not
g83371 not n47190 ; n47190_not
g83372 not n29910 ; n29910_not
g83373 not n22467 ; n22467_not
g83374 not n22476 ; n22476_not
g83375 not n40692 ; n40692_not
g83376 not n29901 ; n29901_not
g83377 not n22197 ; n22197_not
g83378 not n22485 ; n22485_not
g83379 not n52446 ; n52446_not
g83380 not n38064 ; n38064_not
g83381 not n22494 ; n22494_not
g83382 not n29730 ; n29730_not
g83383 not n22863 ; n22863_not
g83384 not n40737 ; n40737_not
g83385 not n22881 ; n22881_not
g83386 not n52473 ; n52473_not
g83387 not n29703 ; n29703_not
g83388 not n22908 ; n22908_not
g83389 not n29712 ; n29712_not
g83390 not n29721 ; n29721_not
g83391 not n22926 ; n22926_not
g83392 not n22944 ; n22944_not
g83393 not n22953 ; n22953_not
g83394 not n22971 ; n22971_not
g83395 not n29604 ; n29604_not
g83396 not n40746 ; n40746_not
g83397 not n29613 ; n29613_not
g83398 not n38019 ; n38019_not
g83399 not n40755 ; n40755_not
g83400 not n22296 ; n22296_not
g83401 not n23088 ; n23088_not
g83402 not n50934 ; n50934_not
g83403 not n22683 ; n22683_not
g83404 not n22692 ; n22692_not
g83405 not n50943 ; n50943_not
g83406 not n22719 ; n22719_not
g83407 not n22728 ; n22728_not
g83408 not n22737 ; n22737_not
g83409 not n22746 ; n22746_not
g83410 not n22755 ; n22755_not
g83411 not n29820 ; n29820_not
g83412 not n22764 ; n22764_not
g83413 not n22773 ; n22773_not
g83414 not n22782 ; n22782_not
g83415 not n22791 ; n22791_not
g83416 not n50961 ; n50961_not
g83417 not n47145 ; n47145_not
g83418 not n22809 ; n22809_not
g83419 not n22818 ; n22818_not
g83420 not n22836 ; n22836_not
g83421 not n29532 ; n29532_not
g83422 not n22854 ; n22854_not
g83423 not n20973 ; n20973_not
g83424 not n41097 ; n41097_not
g83425 not n20649 ; n20649_not
g83426 not n20982 ; n20982_not
g83427 not n20991 ; n20991_not
g83428 not n41295 ; n41295_not
g83429 not n53391 ; n53391_not
g83430 not n30297 ; n30297_not
g83431 not n53373 ; n53373_not
g83432 not n20595 ; n20595_not
g83433 not n21099 ; n21099_not
g83434 not n41277 ; n41277_not
g83435 not n20568 ; n20568_not
g83436 not n30279 ; n30279_not
g83437 not n20559 ; n20559_not
g83438 not n41268 ; n41268_not
g83439 not n41169 ; n41169_not
g83440 not n21189 ; n21189_not
g83441 not n53355 ; n53355_not
g83442 not n21198 ; n21198_not
g83443 not n41178 ; n41178_not
g83444 not n21279 ; n21279_not
g83445 not n21297 ; n21297_not
g83446 not n41187 ; n41187_not
g83447 not n53445 ; n53445_not
g83448 not n20748 ; n20748_not
g83449 not n53436 ; n53436_not
g83450 not n20739 ; n20739_not
g83451 not n41358 ; n41358_not
g83452 not n20829 ; n20829_not
g83453 not n20838 ; n20838_not
g83454 not n20847 ; n20847_not
g83455 not n20856 ; n20856_not
g83456 not n20865 ; n20865_not
g83457 not n20874 ; n20874_not
g83458 not n20883 ; n20883_not
g83459 not n20892 ; n20892_not
g83460 not n20694 ; n20694_not
g83461 not n53418 ; n53418_not
g83462 not n20685 ; n20685_not
g83463 not n20919 ; n20919_not
g83464 not n50745 ; n50745_not
g83465 not n20928 ; n20928_not
g83466 not n20937 ; n20937_not
g83467 not n20946 ; n20946_not
g83468 not n41079 ; n41079_not
g83469 not n20955 ; n20955_not
g83470 not n20964 ; n20964_not
g83471 not n41088 ; n41088_not
g83472 not n20658 ; n20658_not
g83473 not n53247 ; n53247_not
g83474 not n53238 ; n53238_not
g83475 not n50763 ; n50763_not
g83476 not n22089 ; n22089_not
g83477 not n50772 ; n50772_not
g83478 not n47217 ; n47217_not
g83479 not n38091 ; n38091_not
g83480 not n50781 ; n50781_not
g83481 not n22179 ; n22179_not
g83482 not n50790 ; n50790_not
g83483 not n50808 ; n50808_not
g83484 not n22269 ; n22269_not
g83485 not n50817 ; n50817_not
g83486 not n47208 ; n47208_not
g83487 not n50826 ; n50826_not
g83488 not n22287 ; n22287_not
g83489 not n22359 ; n22359_not
g83490 not n21369 ; n21369_not
g83491 not n21387 ; n21387_not
g83492 not n53346 ; n53346_not
g83493 not n41196 ; n41196_not
g83494 not n30099 ; n30099_not
g83495 not n21459 ; n21459_not
g83496 not n21477 ; n21477_not
g83497 not n21495 ; n21495_not
g83498 not n53328 ; n53328_not
g83499 not n21468 ; n21468_not
g83500 not n40638 ; n40638_not
g83501 not n40647 ; n40647_not
g83502 not n50754 ; n50754_not
g83503 not n53283 ; n53283_not
g83504 not n21378 ; n21378_not
g83505 not n40656 ; n40656_not
g83506 not n40665 ; n40665_not
g83507 not n53265 ; n53265_not
g83508 not n53256 ; n53256_not
g83509 not n21288 ; n21288_not
g83510 not n29343 ; n29343_not
g83511 not n23592 ; n23592_not
g83512 not n23619 ; n23619_not
g83513 not n38406 ; n38406_not
g83514 not n23583 ; n23583_not
g83515 not n29280 ; n29280_not
g83516 not n23628 ; n23628_not
g83517 not n23574 ; n23574_not
g83518 not n38505 ; n38505_not
g83519 not n29244 ; n29244_not
g83520 not n23565 ; n23565_not
g83521 not n29325 ; n29325_not
g83522 not n23556 ; n23556_not
g83523 not n29253 ; n29253_not
g83524 not n23547 ; n23547_not
g83525 not n23646 ; n23646_not
g83526 not n29316 ; n29316_not
g83527 not n38514 ; n38514_not
g83528 not n23538 ; n23538_not
g83529 not n23529 ; n23529_not
g83530 not n47046 ; n47046_not
g83531 not n29307 ; n29307_not
g83532 not n51195 ; n51195_not
g83533 not n47064 ; n47064_not
g83534 not n29370 ; n29370_not
g83535 not n38451 ; n38451_not
g83536 not n22827 ; n22827_not
g83537 not n38442 ; n38442_not
g83538 not n38433 ; n38433_not
g83539 not n38424 ; n38424_not
g83540 not n38415 ; n38415_not
g83541 not n47055 ; n47055_not
g83542 not n29352 ; n29352_not
g83543 not n29334 ; n29334_not
g83544 not n23754 ; n23754_not
g83545 not n23763 ; n23763_not
g83546 not n38352 ; n38352_not
g83547 not n38532 ; n38532_not
g83548 not n23781 ; n23781_not
g83549 not n23295 ; n23295_not
g83550 not n40827 ; n40827_not
g83551 not n52536 ; n52536_not
g83552 not n23286 ; n23286_not
g83553 not n23277 ; n23277_not
g83554 not n23268 ; n23268_not
g83555 not n38343 ; n38343_not
g83556 not n29154 ; n29154_not
g83557 not n23259 ; n23259_not
g83558 not n23808 ; n23808_not
g83559 not n29226 ; n29226_not
g83560 not n23826 ; n23826_not
g83561 not n40863 ; n40863_not
g83562 not n38334 ; n38334_not
g83563 not n29217 ; n29217_not
g83564 not n40845 ; n40845_not
g83565 not n23196 ; n23196_not
g83566 not n40836 ; n40836_not
g83567 not n23664 ; n23664_not
g83568 not n23673 ; n23673_not
g83569 not n23493 ; n23493_not
g83570 not n23484 ; n23484_not
g83571 not n23475 ; n23475_not
g83572 not n38370 ; n38370_not
g83573 not n23466 ; n23466_not
g83574 not n23691 ; n23691_not
g83575 not n23457 ; n23457_not
g83576 not n52527 ; n52527_not
g83577 not n23448 ; n23448_not
g83578 not n23439 ; n23439_not
g83579 not n23709 ; n23709_not
g83580 not n23718 ; n23718_not
g83581 not n23394 ; n23394_not
g83582 not n38361 ; n38361_not
g83583 not n23385 ; n23385_not
g83584 not n23736 ; n23736_not
g83585 not n23376 ; n23376_not
g83586 not n23367 ; n23367_not
g83587 not n29262 ; n29262_not
g83588 not n23358 ; n23358_not
g83589 not n23349 ; n23349_not
g83590 not n29514 ; n29514_not
g83591 not n22962 ; n22962_not
g83592 not n29523 ; n29523_not
g83593 not n23079 ; n23079_not
g83594 not n52482 ; n52482_not
g83595 not n29550 ; n29550_not
g83596 not n51069 ; n51069_not
g83597 not n29640 ; n29640_not
g83598 not n29541 ; n29541_not
g83599 not n47127 ; n47127_not
g83600 not n51078 ; n51078_not
g83601 not n23169 ; n23169_not
g83602 not n23178 ; n23178_not
g83603 not n23187 ; n23187_not
g83604 not n29622 ; n29622_not
g83605 not n47118 ; n47118_not
g83606 not n52491 ; n52491_not
g83607 not n51096 ; n51096_not
g83608 not n22872 ; n22872_not
g83609 not n29451 ; n29451_not
g83610 not n29442 ; n29442_not
g83611 not n40791 ; n40791_not
g83612 not n51177 ; n51177_not
g83613 not n29433 ; n29433_not
g83614 not n52518 ; n52518_not
g83615 not n47073 ; n47073_not
g83616 not n29424 ; n29424_not
g83617 not n38460 ; n38460_not
g83618 not n29415 ; n29415_not
g83619 not n51186 ; n51186_not
g83620 not n47091 ; n47091_not
g83621 not n22917 ; n22917_not
g83622 not n40782 ; n40782_not
g83623 not n51159 ; n51159_not
g83624 not n51087 ; n51087_not
g83625 not n51168 ; n51168_not
g83626 not n46371 ; n46371_not
g83627 not n30693 ; n30693_not
g83628 not n53553 ; n53553_not
g83629 not n41439 ; n41439_not
g83630 not n50709 ; n50709_not
g83631 not n30882 ; n30882_not
g83632 not n19146 ; n19146_not
g83633 not n53922 ; n53922_not
g83634 not n38118 ; n38118_not
g83635 not n19137 ; n19137_not
g83636 not n30873 ; n30873_not
g83637 not n53913 ; n53913_not
g83638 not n30864 ; n30864_not
g83639 not n19128 ; n19128_not
g83640 not n47262 ; n47262_not
g83641 not n19605 ; n19605_not
g83642 not n37641 ; n37641_not
g83643 not n30855 ; n30855_not
g83644 not n53904 ; n53904_not
g83645 not n19614 ; n19614_not
g83646 not n30846 ; n30846_not
g83647 not n19623 ; n19623_not
g83648 not n19632 ; n19632_not
g83649 not n19191 ; n19191_not
g83650 not n37713 ; n37713_not
g83651 not n19182 ; n19182_not
g83652 not n19506 ; n19506_not
g83653 not n37704 ; n37704_not
g83654 not n19515 ; n19515_not
g83655 not n30918 ; n30918_not
g83656 not n19173 ; n19173_not
g83657 not n19524 ; n19524_not
g83658 not n19533 ; n19533_not
g83659 not n53319 ; n53319_not
g83660 not n19542 ; n19542_not
g83661 not n53940 ; n53940_not
g83662 not n19551 ; n19551_not
g83663 not n47280 ; n47280_not
g83664 not n41286 ; n41286_not
g83665 not n19560 ; n19560_not
g83666 not n53931 ; n53931_not
g83667 not n30891 ; n30891_not
g83668 not n47253 ; n47253_not
g83669 not n30747 ; n30747_not
g83670 not n19704 ; n19704_not
g83671 not n50727 ; n50727_not
g83672 not n30783 ; n30783_not
g83673 not n30756 ; n30756_not
g83674 not n19713 ; n19713_not
g83675 not n30774 ; n30774_not
g83676 not n19722 ; n19722_not
g83677 not n19731 ; n19731_not
g83678 not n53832 ; n53832_not
g83679 not n30765 ; n30765_not
g83680 not n19056 ; n19056_not
g83681 not n30558 ; n30558_not
g83682 not n19740 ; n19740_not
g83683 not n30567 ; n30567_not
g83684 not n53823 ; n53823_not
g83685 not n30576 ; n30576_not
g83686 not n30585 ; n30585_not
g83687 not n45165 ; n45165_not
g83688 not n30837 ; n30837_not
g83689 not n19641 ; n19641_not
g83690 not n30828 ; n30828_not
g83691 not n19650 ; n19650_not
g83692 not n50718 ; n50718_not
g83693 not n30819 ; n30819_not
g83694 not n19092 ; n19092_not
g83695 not n53364 ; n53364_not
g83696 not n30738 ; n30738_not
g83697 not n19083 ; n19083_not
g83698 not n53850 ; n53850_not
g83699 not n53841 ; n53841_not
g83700 not n30792 ; n30792_not
g83701 not n18642 ; n18642_not
g83702 not n18633 ; n18633_not
g83703 not n37812 ; n37812_not
g83704 not n18624 ; n18624_not
g83705 not n41808 ; n41808_not
g83706 not n18615 ; n18615_not
g83707 not n19290 ; n19290_not
g83708 not n54057 ; n54057_not
g83709 not n30963 ; n30963_not
g83710 not n19308 ; n19308_not
g83711 not n54048 ; n54048_not
g83712 not n19317 ; n19317_not
g83713 not n30972 ; n30972_not
g83714 not n50655 ; n50655_not
g83715 not n19326 ; n19326_not
g83716 not n19281 ; n19281_not
g83717 not n19335 ; n19335_not
g83718 not n19272 ; n19272_not
g83719 not n19344 ; n19344_not
g83720 not n37803 ; n37803_not
g83721 not n54039 ; n54039_not
g83722 not n41781 ; n41781_not
g83723 not n31098 ; n31098_not
g83724 not n18741 ; n18741_not
g83725 not n38028 ; n38028_not
g83726 not n50646 ; n50646_not
g83727 not n19218 ; n19218_not
g83728 not n41835 ; n41835_not
g83729 not n18732 ; n18732_not
g83730 not n46641 ; n46641_not
g83731 not n19227 ; n19227_not
g83732 not n18723 ; n18723_not
g83733 not n31089 ; n31089_not
g83734 not n41790 ; n41790_not
g83735 not n18714 ; n18714_not
g83736 not n37821 ; n37821_not
g83737 not n18705 ; n18705_not
g83738 not n19245 ; n19245_not
g83739 not n41817 ; n41817_not
g83740 not n18660 ; n18660_not
g83741 not n19263 ; n19263_not
g83742 not n30954 ; n30954_not
g83743 not n54066 ; n54066_not
g83744 not n18651 ; n18651_not
g83745 not n19434 ; n19434_not
g83746 not n30981 ; n30981_not
g83747 not n50682 ; n50682_not
g83748 not n19443 ; n19443_not
g83749 not n19452 ; n19452_not
g83750 not n38073 ; n38073_not
g83751 not n19461 ; n19461_not
g83752 not n50691 ; n50691_not
g83753 not n19470 ; n19470_not
g83754 not n37740 ; n37740_not
g83755 not n47307 ; n47307_not
g83756 not n37731 ; n37731_not
g83757 not n37722 ; n37722_not
g83758 not n30936 ; n30936_not
g83759 not n19353 ; n19353_not
g83760 not n19362 ; n19362_not
g83761 not n19371 ; n19371_not
g83762 not n19380 ; n19380_not
g83763 not n50664 ; n50664_not
g83764 not n53274 ; n53274_not
g83765 not n19407 ; n19407_not
g83766 not n19236 ; n19236_not
g83767 not n19416 ; n19416_not
g83768 not n30990 ; n30990_not
g83769 not n50673 ; n50673_not
g83770 not n47325 ; n47325_not
g83771 not n19425 ; n19425_not
g83772 not n20199 ; n20199_not
g83773 not n19920 ; n19920_not
g83774 not n53571 ; n53571_not
g83775 not n40908 ; n40908_not
g83776 not n53526 ; n53526_not
g83777 not n53562 ; n53562_not
g83778 not n30495 ; n30495_not
g83779 not n30459 ; n30459_not
g83780 not n20289 ; n20289_not
g83781 not n20298 ; n20298_not
g83782 not n30477 ; n30477_not
g83783 not n53535 ; n53535_not
g83784 not n40890 ; n40890_not
g83785 not n30468 ; n30468_not
g83786 not n40881 ; n40881_not
g83787 not n53508 ; n53508_not
g83788 not n30549 ; n30549_not
g83789 not n40935 ; n40935_not
g83790 not n53490 ; n53490_not
g83791 not n53625 ; n53625_not
g83792 not n30369 ; n30369_not
g83793 not n45147 ; n45147_not
g83794 not n53616 ; n53616_not
g83795 not n53607 ; n53607_not
g83796 not n30378 ; n30378_not
g83797 not n40926 ; n40926_not
g83798 not n30387 ; n30387_not
g83799 not n30396 ; n30396_not
g83800 not n40917 ; n40917_not
g83801 not n53580 ; n53580_not
g83802 not n30288 ; n30288_not
g83803 not n20577 ; n20577_not
g83804 not n40944 ; n40944_not
g83805 not n38109 ; n38109_not
g83806 not n47235 ; n47235_not
g83807 not n20667 ; n20667_not
g83808 not n40953 ; n40953_not
g83809 not n41385 ; n41385_not
g83810 not n40962 ; n40962_not
g83811 not n20757 ; n20757_not
g83812 not n20766 ; n20766_not
g83813 not n40971 ; n40971_not
g83814 not n20784 ; n20784_not
g83815 not n20793 ; n20793_not
g83816 not n40980 ; n40980_not
g83817 not n41367 ; n41367_not
g83818 not n19830 ; n19830_not
g83819 not n20379 ; n20379_not
g83820 not n20388 ; n20388_not
g83821 not n40872 ; n40872_not
g83822 not n20397 ; n20397_not
g83823 not n53481 ; n53481_not
g83824 not n19803 ; n19803_not
g83825 not n20469 ; n20469_not
g83826 not n53463 ; n53463_not
g83827 not n20478 ; n20478_not
g83828 not n20487 ; n20487_not
g83829 not n20496 ; n20496_not
g83830 not n30684 ; n30684_not
g83831 not n53751 ; n53751_not
g83832 not n30675 ; n30675_not
g83833 not n53742 ; n53742_not
g83834 not n30666 ; n30666_not
g83835 not n30657 ; n30657_not
g83836 not n53733 ; n53733_not
g83837 not n30486 ; n30486_not
g83838 not n30648 ; n30648_not
g83839 not n53724 ; n53724_not
g83840 not n30639 ; n30639_not
g83841 not n53814 ; n53814_not
g83842 not n30594 ; n30594_not
g83843 not n53805 ; n53805_not
g83844 not n53409 ; n53409_not
g83845 not n19812 ; n19812_not
g83846 not n45156 ; n45156_not
g83847 not n53760 ; n53760_not
g83848 not n38145 ; n38145_not
g83849 not n53661 ; n53661_not
g83850 not n50736 ; n50736_not
g83851 not n53652 ; n53652_not
g83852 not n53643 ; n53643_not
g83853 not n53634 ; n53634_not
g83854 not n53715 ; n53715_not
g83855 not n19902 ; n19902_not
g83856 not n53706 ; n53706_not
g83857 not n53454 ; n53454_not
g83858 not n41376 ; n41376_not
g83859 not n53670 ; n53670_not
g83860 not n51528 ; n51528_not
g83861 not n26652 ; n26652_not
g83862 not n26661 ; n26661_not
g83863 not n39702 ; n39702_not
g83864 not n51519 ; n51519_not
g83865 not n39207 ; n39207_not
g83866 not n26670 ; n26670_not
g83867 not n27813 ; n27813_not
g83868 not n52293 ; n52293_not
g83869 not n39153 ; n39153_not
g83870 not n51843 ; n51843_not
g83871 not n39180 ; n39180_not
g83872 not n46542 ; n46542_not
g83873 not n46119 ; n46119_not
g83874 not n51852 ; n51852_not
g83875 not n52284 ; n52284_not
g83876 not n39216 ; n39216_not
g83877 not n46128 ; n46128_not
g83878 not n51708 ; n51708_not
g83879 not n39144 ; n39144_not
g83880 not n46137 ; n46137_not
g83881 not n26706 ; n26706_not
g83882 not n52275 ; n52275_not
g83883 not n26175 ; n26175_not
g83884 not n26715 ; n26715_not
g83885 not n45804 ; n45804_not
g83886 not n51870 ; n51870_not
g83887 not n26247 ; n26247_not
g83888 not n26580 ; n26580_not
g83889 not n52329 ; n52329_not
g83890 not n46047 ; n46047_not
g83891 not n39810 ; n39810_not
g83892 not n39171 ; n39171_not
g83893 not n51546 ; n51546_not
g83894 not n46056 ; n46056_not
g83895 not n26607 ; n26607_not
g83896 not n39801 ; n39801_not
g83897 not n46065 ; n46065_not
g83898 not n26616 ; n26616_not
g83899 not n51825 ; n51825_not
g83900 not n45840 ; n45840_not
g83901 not n51537 ; n51537_not
g83902 not n26625 ; n26625_not
g83903 not n46560 ; n46560_not
g83904 not n46074 ; n46074_not
g83905 not n26634 ; n26634_not
g83906 not n46083 ; n46083_not
g83907 not n27840 ; n27840_not
g83908 not n45831 ; n45831_not
g83909 not n27831 ; n27831_not
g83910 not n26643 ; n26643_not
g83911 not n46092 ; n46092_not
g83912 not n39243 ; n39243_not
g83913 not n51483 ; n51483_not
g83914 not n27732 ; n27732_not
g83915 not n26940 ; n26940_not
g83916 not n39252 ; n39252_not
g83917 not n26760 ; n26760_not
g83918 not n46173 ; n46173_not
g83919 not n39261 ; n39261_not
g83920 not n27723 ; n27723_not
g83921 not n52257 ; n52257_not
g83922 not n51726 ; n51726_not
g83923 not n39270 ; n39270_not
g83924 not n46182 ; n46182_not
g83925 not n27714 ; n27714_not
g83926 not n51474 ; n51474_not
g83927 not n46191 ; n46191_not
g83928 not n52248 ; n52248_not
g83929 not n27705 ; n27705_not
g83930 not n39306 ; n39306_not
g83931 not n39315 ; n39315_not
g83932 not n51465 ; n51465_not
g83933 not n39324 ; n39324_not
g83934 not n52239 ; n52239_not
g83935 not n39333 ; n39333_not
g83936 not n46146 ; n46146_not
g83937 not n26166 ; n26166_not
g83938 not n26724 ; n26724_not
g83939 not n51492 ; n51492_not
g83940 not n46533 ; n46533_not
g83941 not n39711 ; n39711_not
g83942 not n26733 ; n26733_not
g83943 not n39225 ; n39225_not
g83944 not n46155 ; n46155_not
g83945 not n52266 ; n52266_not
g83946 not n26922 ; n26922_not
g83947 not n26157 ; n26157_not
g83948 not n26742 ; n26742_not
g83949 not n39234 ; n39234_not
g83950 not n27750 ; n27750_not
g83951 not n39135 ; n39135_not
g83952 not n51717 ; n51717_not
g83953 not n27741 ; n27741_not
g83954 not n26931 ; n26931_not
g83955 not n26751 ; n26751_not
g83956 not n46164 ; n46164_not
g83957 not n28056 ; n28056_not
g83958 not n38820 ; n38820_not
g83959 not n51618 ; n51618_not
g83960 not n39072 ; n39072_not
g83961 not n51735 ; n51735_not
g83962 not n26373 ; n26373_not
g83963 not n38811 ; n38811_not
g83964 not n38802 ; n38802_not
g83965 not n26382 ; n26382_not
g83966 not n52392 ; n52392_not
g83967 not n28038 ; n28038_not
g83968 not n26355 ; n26355_not
g83969 not n26391 ; n26391_not
g83970 not n51609 ; n51609_not
g83971 not n26346 ; n26346_not
g83972 not n26409 ; n26409_not
g83973 not n52383 ; n52383_not
g83974 not n26337 ; n26337_not
g83975 not n26418 ; n26418_not
g83976 not n39603 ; n39603_not
g83977 not n26427 ; n26427_not
g83978 not n39090 ; n39090_not
g83979 not n26436 ; n26436_not
g83980 not n46623 ; n46623_not
g83981 not n28155 ; n28155_not
g83982 not n28146 ; n28146_not
g83983 not n28029 ; n28029_not
g83984 not n26256 ; n26256_not
g83985 not n45741 ; n45741_not
g83986 not n45750 ; n45750_not
g83987 not n38901 ; n38901_not
g83988 not n39027 ; n39027_not
g83989 not n51636 ; n51636_not
g83990 not n26274 ; n26274_not
g83991 not n26292 ; n26292_not
g83992 not n28119 ; n28119_not
g83993 not n28065 ; n28065_not
g83994 not n26319 ; n26319_not
g83995 not n28092 ; n28092_not
g83996 not n39045 ; n39045_not
g83997 not n27228 ; n27228_not
g83998 not n45813 ; n45813_not
g83999 not n28083 ; n28083_not
g84000 not n39054 ; n39054_not
g84001 not n46650 ; n46650_not
g84002 not n51627 ; n51627_not
g84003 not n26508 ; n26508_not
g84004 not n27930 ; n27930_not
g84005 not n26517 ; n26517_not
g84006 not n27921 ; n27921_not
g84007 not n46605 ; n46605_not
g84008 not n51573 ; n51573_not
g84009 not n26526 ; n26526_not
g84010 not n26535 ; n26535_not
g84011 not n52347 ; n52347_not
g84012 not n39162 ; n39162_not
g84013 not n26544 ; n26544_not
g84014 not n51672 ; n51672_not
g84015 not n27903 ; n27903_not
g84016 not n38154 ; n38154_not
g84017 not n26265 ; n26265_not
g84018 not n26553 ; n26553_not
g84019 not n51564 ; n51564_not
g84020 not n26562 ; n26562_not
g84021 not n52338 ; n52338_not
g84022 not n46029 ; n46029_not
g84023 not n51681 ; n51681_not
g84024 not n51807 ; n51807_not
g84025 not n26571 ; n26571_not
g84026 not n51555 ; n51555_not
g84027 not n46038 ; n46038_not
g84028 not n39612 ; n39612_not
g84029 not n26445 ; n26445_not
g84030 not n45921 ; n45921_not
g84031 not n26454 ; n26454_not
g84032 not n52374 ; n52374_not
g84033 not n26463 ; n26463_not
g84034 not n45903 ; n45903_not
g84035 not n51591 ; n51591_not
g84036 not n26472 ; n26472_not
g84037 not n51753 ; n51753_not
g84038 not n26481 ; n26481_not
g84039 not n39900 ; n39900_not
g84040 not n52365 ; n52365_not
g84041 not n51762 ; n51762_not
g84042 not n51663 ; n51663_not
g84043 not n26490 ; n26490_not
g84044 not n39117 ; n39117_not
g84045 not n38730 ; n38730_not
g84046 not n45246 ; n45246_not
g84047 not n51582 ; n51582_not
g84048 not n38721 ; n38721_not
g84049 not n38712 ; n38712_not
g84050 not n51780 ; n51780_not
g84051 not n38703 ; n38703_not
g84052 not n52356 ; n52356_not
g84053 not n27147 ; n27147_not
g84054 not n52095 ; n52095_not
g84055 not n39360 ; n39360_not
g84056 not n27480 ; n27480_not
g84057 not n51249 ; n51249_not
g84058 not n27156 ; n27156_not
g84059 not n51816 ; n51816_not
g84060 not n27471 ; n27471_not
g84061 not n46344 ; n46344_not
g84062 not n27174 ; n27174_not
g84063 not n39063 ; n39063_not
g84064 not n27462 ; n27462_not
g84065 not n46425 ; n46425_not
g84066 not n39009 ; n39009_not
g84067 not n27453 ; n27453_not
g84068 not n46353 ; n46353_not
g84069 not n52086 ; n52086_not
g84070 not n27444 ; n27444_not
g84071 not n27192 ; n27192_not
g84072 not n39018 ; n39018_not
g84073 not n51258 ; n51258_not
g84074 not n45714 ; n45714_not
g84075 not n51339 ; n51339_not
g84076 not n46308 ; n46308_not
g84077 not n27534 ; n27534_not
g84078 not n27057 ; n27057_not
g84079 not n27066 ; n27066_not
g84080 not n45705 ; n45705_not
g84081 not n39342 ; n39342_not
g84082 not n27525 ; n27525_not
g84083 not n51861 ; n51861_not
g84084 not n46317 ; n46317_not
g84085 not n27084 ; n27084_not
g84086 not n27516 ; n27516_not
g84087 not n46443 ; n46443_not
g84088 not n27507 ; n27507_not
g84089 not n46326 ; n46326_not
g84090 not n39351 ; n39351_not
g84091 not n27129 ; n27129_not
g84092 not n46335 ; n46335_not
g84093 not n27075 ; n27075_not
g84094 not n27291 ; n27291_not
g84095 not n27390 ; n27390_not
g84096 not n39423 ; n39423_not
g84097 not n46380 ; n46380_not
g84098 not n51285 ; n51285_not
g84099 not n27309 ; n27309_not
g84100 not n27318 ; n27318_not
g84101 not n27381 ; n27381_not
g84102 not n52059 ; n52059_not
g84103 not n27165 ; n27165_not
g84104 not n27327 ; n27327_not
g84105 not n39414 ; n39414_not
g84106 not n27372 ; n27372_not
g84107 not n27336 ; n27336_not
g84108 not n27345 ; n27345_not
g84109 not n39405 ; n39405_not
g84110 not n27363 ; n27363_not
g84111 not n27354 ; n27354_not
g84112 not n51276 ; n51276_not
g84113 not n27435 ; n27435_not
g84114 not n39450 ; n39450_not
g84115 not n52077 ; n52077_not
g84116 not n27426 ; n27426_not
g84117 not n27237 ; n27237_not
g84118 not n27246 ; n27246_not
g84119 not n46407 ; n46407_not
g84120 not n27417 ; n27417_not
g84121 not n27255 ; n27255_not
g84122 not n39441 ; n39441_not
g84123 not n51294 ; n51294_not
g84124 not n27264 ; n27264_not
g84125 not n27408 ; n27408_not
g84126 not n27273 ; n27273_not
g84127 not n52068 ; n52068_not
g84128 not n27282 ; n27282_not
g84129 not n39432 ; n39432_not
g84130 not n18327 ; n18327_not
g84131 not n51267 ; n51267_not
g84132 not n46236 ; n46236_not
g84133 not n51429 ; n51429_not
g84134 not n27651 ; n27651_not
g84135 not n26085 ; n26085_not
g84136 not n51942 ; n51942_not
g84137 not n26076 ; n26076_not
g84138 not n27642 ; n27642_not
g84139 not n46245 ; n46245_not
g84140 not n52194 ; n52194_not
g84141 not n51951 ; n51951_not
g84142 not n26067 ; n26067_not
g84143 not n27633 ; n27633_not
g84144 not n26904 ; n26904_not
g84145 not n39108 ; n39108_not
g84146 not n26805 ; n26805_not
g84147 not n51456 ; n51456_not
g84148 not n51915 ; n51915_not
g84149 not n26814 ; n26814_not
g84150 not n46209 ; n46209_not
g84151 not n26823 ; n26823_not
g84152 not n39621 ; n39621_not
g84153 not n46515 ; n46515_not
g84154 not n51447 ; n51447_not
g84155 not n26832 ; n26832_not
g84156 not n46218 ; n46218_not
g84157 not n51924 ; n51924_not
g84158 not n26841 ; n26841_not
g84159 not n26850 ; n26850_not
g84160 not n46227 ; n46227_not
g84161 not n51438 ; n51438_not
g84162 not n51906 ; n51906_not
g84163 not n51933 ; n51933_not
g84164 not n27660 ; n27660_not
g84165 not n39531 ; n39531_not
g84166 not n51384 ; n51384_not
g84167 not n52158 ; n52158_not
g84168 not n39522 ; n39522_not
g84169 not n51375 ; n51375_not
g84170 not n52149 ; n52149_not
g84171 not n46290 ; n46290_not
g84172 not n27570 ; n27570_not
g84173 not n51366 ; n51366_not
g84174 not n39513 ; n39513_not
g84175 not n27561 ; n27561_not
g84176 not n51357 ; n51357_not
g84177 not n39504 ; n39504_not
g84178 not n51348 ; n51348_not
g84179 not n27552 ; n27552_not
g84180 not n46452 ; n46452_not
g84181 not n27543 ; n27543_not
g84182 not n27039 ; n27039_not
g84183 not n26913 ; n26913_not
g84184 not n51960 ; n51960_not
g84185 not n27624 ; n27624_not
g84186 not n46254 ; n46254_not
g84187 not n46263 ; n46263_not
g84188 not n52185 ; n52185_not
g84189 not n27615 ; n27615_not
g84190 not n46470 ; n46470_not
g84191 not n27606 ; n27606_not
g84192 not n46272 ; n46272_not
g84193 not n52176 ; n52176_not
g84194 not n51771 ; n51771_not
g84195 not n51393 ; n51393_not
g84196 not n46281 ; n46281_not
g84197 not n52167 ; n52167_not
g84198 not n38622 ; n38622_not
g84199 not n38190 ; n38190_not
g84200 not n24717 ; n24717_not
g84201 not n38181 ; n38181_not
g84202 not n24726 ; n24726_not
g84203 not n24681 ; n24681_not
g84204 not n28830 ; n28830_not
g84205 not n24735 ; n24735_not
g84206 not n38172 ; n38172_not
g84207 not n24744 ; n24744_not
g84208 not n50952 ; n50952_not
g84209 not n38163 ; n38163_not
g84210 not n24753 ; n24753_not
g84211 not n28812 ; n28812_not
g84212 not n24762 ; n24762_not
g84213 not n24771 ; n24771_not
g84214 not n46416 ; n46416_not
g84215 not n24780 ; n24780_not
g84216 not n24654 ; n24654_not
g84217 not n24645 ; n24645_not
g84218 not n24807 ; n24807_not
g84219 not n24636 ; n24636_not
g84220 not n28911 ; n28911_not
g84221 not n38226 ; n38226_not
g84222 not n38604 ; n38604_not
g84223 not n24591 ; n24591_not
g84224 not n28902 ; n28902_not
g84225 not n38217 ; n38217_not
g84226 not n24618 ; n24618_not
g84227 not n52662 ; n52662_not
g84228 not n28074 ; n28074_not
g84229 not n24663 ; n24663_not
g84230 not n38208 ; n38208_not
g84231 not n28128 ; n28128_not
g84232 not n24690 ; n24690_not
g84233 not n52671 ; n52671_not
g84234 not n24942 ; n24942_not
g84235 not n24564 ; n24564_not
g84236 not n24951 ; n24951_not
g84237 not n24555 ; n24555_not
g84238 not n24960 ; n24960_not
g84239 not n28704 ; n28704_not
g84240 not n52707 ; n52707_not
g84241 not n24546 ; n24546_not
g84242 not n45075 ; n45075_not
g84243 not n24519 ; n24519_not
g84244 not n50907 ; n50907_not
g84245 not n40179 ; n40179_not
g84246 not n25059 ; n25059_not
g84247 not n52680 ; n52680_not
g84248 not n25068 ; n25068_not
g84249 not n25077 ; n25077_not
g84250 not n38613 ; n38613_not
g84251 not n24816 ; n24816_not
g84252 not n38640 ; n38640_not
g84253 not n24825 ; n24825_not
g84254 not n24834 ; n24834_not
g84255 not n24843 ; n24843_not
g84256 not n24852 ; n24852_not
g84257 not n24861 ; n24861_not
g84258 not n24609 ; n24609_not
g84259 not n24870 ; n24870_not
g84260 not n24906 ; n24906_not
g84261 not n28740 ; n28740_not
g84262 not n24915 ; n24915_not
g84263 not n24924 ; n24924_not
g84264 not n24933 ; n24933_not
g84265 not n52716 ; n52716_not
g84266 not n28722 ; n28722_not
g84267 not n23844 ; n23844_not
g84268 not n52563 ; n52563_not
g84269 not n38307 ; n38307_not
g84270 not n52572 ; n52572_not
g84271 not n29136 ; n29136_not
g84272 not n23817 ; n23817_not
g84273 not n52581 ; n52581_not
g84274 not n40764 ; n40764_not
g84275 not n29127 ; n29127_not
g84276 not n29082 ; n29082_not
g84277 not n47028 ; n47028_not
g84278 not n29118 ; n29118_not
g84279 not n23772 ; n23772_not
g84280 not n38280 ; n38280_not
g84281 not n40719 ; n40719_not
g84282 not n29028 ; n29028_not
g84283 not n29208 ; n29208_not
g84284 not n23853 ; n23853_not
g84285 not n40854 ; n40854_not
g84286 not n29181 ; n29181_not
g84287 not n23871 ; n23871_not
g84288 not n38325 ; n38325_not
g84289 not n29190 ; n29190_not
g84290 not n40278 ; n40278_not
g84291 not n23862 ; n23862_not
g84292 not n38316 ; n38316_not
g84293 not n38550 ; n38550_not
g84294 not n29163 ; n29163_not
g84295 not n40809 ; n40809_not
g84296 not n47037 ; n47037_not
g84297 not n40629 ; n40629_not
g84298 not n23637 ; n23637_not
g84299 not n29019 ; n29019_not
g84300 not n40089 ; n40089_not
g84301 not n24438 ; n24438_not
g84302 not n38244 ; n38244_not
g84303 not n24456 ; n24456_not
g84304 not n24465 ; n24465_not
g84305 not n24483 ; n24483_not
g84306 not n52653 ; n52653_not
g84307 not n40098 ; n40098_not
g84308 not n47019 ; n47019_not
g84309 not n24528 ; n24528_not
g84310 not n38235 ; n38235_not
g84311 not n28920 ; n28920_not
g84312 not n24573 ; n24573_not
g84313 not n52608 ; n52608_not
g84314 not n29046 ; n29046_not
g84315 not n38271 ; n38271_not
g84316 not n23727 ; n23727_not
g84317 not n52617 ; n52617_not
g84318 not n52626 ; n52626_not
g84319 not n38262 ; n38262_not
g84320 not n40674 ; n40674_not
g84321 not n29055 ; n29055_not
g84322 not n23682 ; n23682_not
g84323 not n38253 ; n38253_not
g84324 not n29037 ; n29037_not
g84325 not n25446 ; n25446_not
g84326 not n27804 ; n27804_not
g84327 not n28380 ; n28380_not
g84328 not n40269 ; n40269_not
g84329 not n52545 ; n52545_not
g84330 not n28344 ; n28344_not
g84331 not n38910 ; n38910_not
g84332 not n28353 ; n28353_not
g84333 not n28362 ; n28362_not
g84334 not n25419 ; n25419_not
g84335 not n28335 ; n28335_not
g84336 not n25518 ; n25518_not
g84337 not n46821 ; n46821_not
g84338 not n28452 ; n28452_not
g84339 not n25527 ; n25527_not
g84340 not n25509 ; n25509_not
g84341 not n38523 ; n38523_not
g84342 not n46812 ; n46812_not
g84343 not n28434 ; n28434_not
g84344 not n52590 ; n52590_not
g84345 not n25491 ; n25491_not
g84346 not n46803 ; n46803_not
g84347 not n28416 ; n28416_not
g84348 not n25464 ; n25464_not
g84349 not n25455 ; n25455_not
g84350 not n28236 ; n28236_not
g84351 not n46713 ; n46713_not
g84352 not n25239 ; n25239_not
g84353 not n28227 ; n28227_not
g84354 not n26058 ; n26058_not
g84355 not n46704 ; n46704_not
g84356 not n28218 ; n28218_not
g84357 not n51690 ; n51690_not
g84358 not n26094 ; n26094_not
g84359 not n26139 ; n26139_not
g84360 not n28191 ; n28191_not
g84361 not n26184 ; n26184_not
g84362 not n28173 ; n28173_not
g84363 not n45723 ; n45723_not
g84364 not n28164 ; n28164_not
g84365 not n26229 ; n26229_not
g84366 not n25374 ; n25374_not
g84367 not n46551 ; n46551_not
g84368 not n51645 ; n51645_not
g84369 not n25365 ; n25365_not
g84370 not n28317 ; n28317_not
g84371 not n25356 ; n25356_not
g84372 not n40197 ; n40197_not
g84373 not n28308 ; n28308_not
g84374 not n28290 ; n28290_not
g84375 not n25329 ; n25329_not
g84376 not n46740 ; n46740_not
g84377 not n46731 ; n46731_not
g84378 not n28263 ; n28263_not
g84379 not n46722 ; n46722_not
g84380 not n28245 ; n28245_not
g84381 not n52455 ; n52455_not
g84382 not n25284 ; n25284_not
g84383 not n25275 ; n25275_not
g84384 not n25266 ; n25266_not
g84385 not n25194 ; n25194_not
g84386 not n25248 ; n25248_not
g84387 not n25185 ; n25185_not
g84388 not n46920 ; n46920_not
g84389 not n25176 ; n25176_not
g84390 not n25167 ; n25167_not
g84391 not n25158 ; n25158_not
g84392 not n25149 ; n25149_not
g84393 not n25293 ; n25293_not
g84394 not n46911 ; n46911_not
g84395 not n25095 ; n25095_not
g84396 not n25086 ; n25086_not
g84397 not n28560 ; n28560_not
g84398 not n40188 ; n40188_not
g84399 not n28650 ; n28650_not
g84400 not n24474 ; n24474_not
g84401 not n28632 ; n28632_not
g84402 not n28614 ; n28614_not
g84403 not n46461 ; n46461_not
g84404 not n24429 ; n24429_not
g84405 not n28506 ; n28506_not
g84406 not n25473 ; n25473_not
g84407 not n46830 ; n46830_not
g84408 not n28470 ; n28470_not
g84409 not n25338 ; n25338_not
g84410 not n46902 ; n46902_not
g84411 not n28542 ; n28542_not
g84412 not n25383 ; n25383_not
g84413 not n50862 ; n50862_not
g84414 not n28272 ; n28272_not
g84415 not n46506 ; n46506_not
g84416 not n28524 ; n28524_not
g84417 not n52635 ; n52635_not
g84418 not n25428 ; n25428_not
g84419 not n42771 ; n42771_not
g84420 not n17076 ; n17076_not
g84421 not n42654 ; n42654_not
g84422 not n54633 ; n54633_not
g84423 not n17094 ; n17094_not
g84424 not n42762 ; n42762_not
g84425 not n55092 ; n55092_not
g84426 not n54642 ; n54642_not
g84427 not n54651 ; n54651_not
g84428 not n42753 ; n42753_not
g84429 not n32295 ; n32295_not
g84430 not n17139 ; n17139_not
g84431 not n17148 ; n17148_not
g84432 not n32277 ; n32277_not
g84433 not n54660 ; n54660_not
g84434 not n42744 ; n42744_not
g84435 not n17166 ; n17166_not
g84436 not n32385 ; n32385_not
g84437 not n55137 ; n55137_not
g84438 not n54561 ; n54561_not
g84439 not n42555 ; n42555_not
g84440 not n32088 ; n32088_not
g84441 not n54570 ; n54570_not
g84442 not n42564 ; n42564_not
g84443 not n55119 ; n55119_not
g84444 not n45219 ; n45219_not
g84445 not n54606 ; n54606_not
g84446 not n32367 ; n32367_not
g84447 not n37632 ; n37632_not
g84448 not n17049 ; n17049_not
g84449 not n32349 ; n32349_not
g84450 not n54615 ; n54615_not
g84451 not n42780 ; n42780_not
g84452 not n17058 ; n17058_not
g84453 not n54624 ; n54624_not
g84454 not n17265 ; n17265_not
g84455 not n42609 ; n42609_not
g84456 not n17274 ; n17274_not
g84457 not n42708 ; n42708_not
g84458 not n55047 ; n55047_not
g84459 not n17283 ; n17283_not
g84460 not n54723 ; n54723_not
g84461 not n17292 ; n17292_not
g84462 not n54732 ; n54732_not
g84463 not n17319 ; n17319_not
g84464 not n54741 ; n54741_not
g84465 not n47640 ; n47640_not
g84466 not n17328 ; n17328_not
g84467 not n54750 ; n54750_not
g84468 not n17337 ; n17337_not
g84469 not n17346 ; n17346_not
g84470 not n42690 ; n42690_not
g84471 not n17355 ; n17355_not
g84472 not n31980 ; n31980_not
g84473 not n42591 ; n42591_not
g84474 not n42735 ; n42735_not
g84475 not n17184 ; n17184_not
g84476 not n17193 ; n17193_not
g84477 not n45237 ; n45237_not
g84478 not n42726 ; n42726_not
g84479 not n17229 ; n17229_not
g84480 not n17238 ; n17238_not
g84481 not n54705 ; n54705_not
g84482 not n42717 ; n42717_not
g84483 not n17247 ; n17247_not
g84484 not n17157 ; n17157_not
g84485 not n17256 ; n17256_not
g84486 not n54714 ; n54714_not
g84487 not n32493 ; n32493_not
g84488 not n16761 ; n16761_not
g84489 not n54435 ; n54435_not
g84490 not n16770 ; n16770_not
g84491 not n32484 ; n32484_not
g84492 not n16365 ; n16365_not
g84493 not n54444 ; n54444_not
g84494 not n50493 ; n50493_not
g84495 not n54453 ; n54453_not
g84496 not n32475 ; n32475_not
g84497 not n16806 ; n16806_not
g84498 not n42519 ; n42519_not
g84499 not n16815 ; n16815_not
g84500 not n42870 ; n42870_not
g84501 not n32466 ; n32466_not
g84502 not n16824 ; n16824_not
g84503 not n45192 ; n45192_not
g84504 not n54462 ; n54462_not
g84505 not n16338 ; n16338_not
g84506 not n16833 ; n16833_not
g84507 not n16671 ; n16671_not
g84508 not n42924 ; n42924_not
g84509 not n16419 ; n16419_not
g84510 not n16680 ; n16680_not
g84511 not n55227 ; n55227_not
g84512 not n54408 ; n54408_not
g84513 not n16707 ; n16707_not
g84514 not n16716 ; n16716_not
g84515 not n42915 ; n42915_not
g84516 not n16725 ; n16725_not
g84517 not n16734 ; n16734_not
g84518 not n45174 ; n45174_not
g84519 not n54417 ; n54417_not
g84520 not n42906 ; n42906_not
g84521 not n16743 ; n16743_not
g84522 not n16383 ; n16383_not
g84523 not n16752 ; n16752_not
g84524 not n54426 ; n54426_not
g84525 not n55209 ; n55209_not
g84526 not n16374 ; n16374_not
g84527 not n16293 ; n16293_not
g84528 not n16914 ; n16914_not
g84529 not n16284 ; n16284_not
g84530 not n16923 ; n16923_not
g84531 not n42825 ; n42825_not
g84532 not n54516 ; n54516_not
g84533 not n16932 ; n16932_not
g84534 not n55155 ; n55155_not
g84535 not n16275 ; n16275_not
g84536 not n42546 ; n42546_not
g84537 not n16941 ; n16941_not
g84538 not n54525 ; n54525_not
g84539 not n42816 ; n42816_not
g84540 not n16950 ; n16950_not
g84541 not n54534 ; n54534_not
g84542 not n54543 ; n54543_not
g84543 not n42807 ; n42807_not
g84544 not n32394 ; n32394_not
g84545 not n54552 ; n54552_not
g84546 not n42861 ; n42861_not
g84547 not n32457 ; n32457_not
g84548 not n16329 ; n16329_not
g84549 not n16842 ; n16842_not
g84550 not n54471 ; n54471_not
g84551 not n42852 ; n42852_not
g84552 not n32448 ; n32448_not
g84553 not n16851 ; n16851_not
g84554 not n55182 ; n55182_not
g84555 not n16860 ; n16860_not
g84556 not n54480 ; n54480_not
g84557 not n32439 ; n32439_not
g84558 not n32358 ; n32358_not
g84559 not n42843 ; n42843_not
g84560 not n54507 ; n54507_not
g84561 not n42834 ; n42834_not
g84562 not n55164 ; n55164_not
g84563 not n16905 ; n16905_not
g84564 not n31953 ; n31953_not
g84565 not n17382 ; n17382_not
g84566 not n54831 ; n54831_not
g84567 not n17373 ; n17373_not
g84568 not n42465 ; n42465_not
g84569 not n17364 ; n17364_not
g84570 not n31944 ; n31944_not
g84571 not n42456 ; n42456_not
g84572 not n31935 ; n31935_not
g84573 not n54822 ; n54822_not
g84574 not n47226 ; n47226_not
g84575 not n31926 ; n31926_not
g84576 not n17805 ; n17805_not
g84577 not n17724 ; n17724_not
g84578 not n17454 ; n17454_not
g84579 not n50556 ; n50556_not
g84580 not n17445 ; n17445_not
g84581 not n17436 ; n17436_not
g84582 not n31971 ; n31971_not
g84583 not n42483 ; n42483_not
g84584 not n17427 ; n17427_not
g84585 not n17742 ; n17742_not
g84586 not n31683 ; n31683_not
g84587 not n17418 ; n17418_not
g84588 not n54129 ; n54129_not
g84589 not n31962 ; n31962_not
g84590 not n17409 ; n17409_not
g84591 not n31692 ; n31692_not
g84592 not n17391 ; n17391_not
g84593 not n50196 ; n50196_not
g84594 not n17760 ; n17760_not
g84595 not n37524 ; n37524_not
g84596 not n50565 ; n50565_not
g84597 not n50574 ; n50574_not
g84598 not n31728 ; n31728_not
g84599 not n47541 ; n47541_not
g84600 not n31881 ; n31881_not
g84601 not n31737 ; n31737_not
g84602 not n54156 ; n54156_not
g84603 not n31872 ; n31872_not
g84604 not n17904 ; n17904_not
g84605 not n47532 ; n47532_not
g84606 not n54165 ; n54165_not
g84607 not n17913 ; n17913_not
g84608 not n50583 ; n50583_not
g84609 not n31863 ; n31863_not
g84610 not n17850 ; n17850_not
g84611 not n47523 ; n47523_not
g84612 not n31854 ; n31854_not
g84613 not n17814 ; n17814_not
g84614 not n31917 ; n31917_not
g84615 not n37830 ; n37830_not
g84616 not n42438 ; n42438_not
g84617 not n17832 ; n17832_not
g84618 not n31908 ; n31908_not
g84619 not n31719 ; n31719_not
g84620 not n54813 ; n54813_not
g84621 not n47550 ; n47550_not
g84622 not n54804 ; n54804_not
g84623 not n31890 ; n31890_not
g84624 not n42645 ; n42645_not
g84625 not n17463 ; n17463_not
g84626 not n41448 ; n41448_not
g84627 not n17472 ; n17472_not
g84628 not n17481 ; n17481_not
g84629 not n54903 ; n54903_not
g84630 not n17490 ; n17490_not
g84631 not n32079 ; n32079_not
g84632 not n54912 ; n54912_not
g84633 not n42618 ; n42618_not
g84634 not n17508 ; n17508_not
g84635 not n17517 ; n17517_not
g84636 not n31809 ; n31809_not
g84637 not n17526 ; n17526_not
g84638 not n54084 ; n54084_not
g84639 not n17535 ; n17535_not
g84640 not n17544 ; n17544_not
g84641 not n42681 ; n42681_not
g84642 not n42636 ; n42636_not
g84643 not n17067 ; n17067_not
g84644 not n50529 ; n50529_not
g84645 not n54840 ; n54840_not
g84646 not n17580 ; n17580_not
g84647 not n17571 ; n17571_not
g84648 not n17562 ; n17562_not
g84649 not n42528 ; n42528_not
g84650 not n17553 ; n17553_not
g84651 not n17670 ; n17670_not
g84652 not n47613 ; n47613_not
g84653 not n37542 ; n37542_not
g84654 not n50547 ; n50547_not
g84655 not n47604 ; n47604_not
g84656 not n17715 ; n17715_not
g84657 not n37533 ; n37533_not
g84658 not n47181 ; n47181_not
g84659 not n47631 ; n47631_not
g84660 not n54075 ; n54075_not
g84661 not n50538 ; n50538_not
g84662 not n42573 ; n42573_not
g84663 not n47622 ; n47622_not
g84664 not n17607 ; n17607_not
g84665 not n17616 ; n17616_not
g84666 not n17634 ; n17634_not
g84667 not n17652 ; n17652_not
g84668 not n15348 ; n15348_not
g84669 not n15339 ; n15339_not
g84670 not n50394 ; n50394_not
g84671 not n15294 ; n15294_not
g84672 not n15285 ; n15285_not
g84673 not n15807 ; n15807_not
g84674 not n15276 ; n15276_not
g84675 not n32718 ; n32718_not
g84676 not n15816 ; n15816_not
g84677 not n37551 ; n37551_not
g84678 not n15267 ; n15267_not
g84679 not n32727 ; n32727_not
g84680 not n15258 ; n15258_not
g84681 not n15249 ; n15249_not
g84682 not n15834 ; n15834_not
g84683 not n47811 ; n47811_not
g84684 not n15438 ; n15438_not
g84685 not n15726 ; n15726_not
g84686 not n15429 ; n15429_not
g84687 not n15744 ; n15744_not
g84688 not n15393 ; n15393_not
g84689 not n15384 ; n15384_not
g84690 not n15375 ; n15375_not
g84691 not n15366 ; n15366_not
g84692 not n15762 ; n15762_not
g84693 not n15357 ; n15357_not
g84694 not n15771 ; n15771_not
g84695 not n32925 ; n32925_not
g84696 not n43266 ; n43266_not
g84697 not n32916 ; n32916_not
g84698 not n32709 ; n32709_not
g84699 not n32583 ; n32583_not
g84700 not n43257 ; n43257_not
g84701 not n37623 ; n37623_not
g84702 not n55173 ; n55173_not
g84703 not n43239 ; n43239_not
g84704 not n15780 ; n15780_not
g84705 not n15852 ; n15852_not
g84706 not n50286 ; n50286_not
g84707 not n15825 ; n15825_not
g84708 not n32961 ; n32961_not
g84709 not n43275 ; n43275_not
g84710 not n32943 ; n32943_not
g84711 not n32934 ; n32934_not
g84712 not n37614 ; n37614_not
g84713 not n33249 ; n33249_not
g84714 not n50367 ; n50367_not
g84715 not n32952 ; n32952_not
g84716 not n47901 ; n47901_not
g84717 not n55128 ; n55128_not
g84718 not n33177 ; n33177_not
g84719 not n33186 ; n33186_not
g84720 not n33195 ; n33195_not
g84721 not n37452 ; n37452_not
g84722 not n43176 ; n43176_not
g84723 not n15078 ; n15078_not
g84724 not n37443 ; n37443_not
g84725 not n37461 ; n37461_not
g84726 not n43185 ; n43185_not
g84727 not n33267 ; n33267_not
g84728 not n15537 ; n15537_not
g84729 not n15528 ; n15528_not
g84730 not n15672 ; n15672_not
g84731 not n15519 ; n15519_not
g84732 not n45084 ; n45084_not
g84733 not n50385 ; n50385_not
g84734 not n15681 ; n15681_not
g84735 not n15492 ; n15492_not
g84736 not n15483 ; n15483_not
g84737 not n15474 ; n15474_not
g84738 not n15465 ; n15465_not
g84739 not n15456 ; n15456_not
g84740 not n15447 ; n15447_not
g84741 not n15717 ; n15717_not
g84742 not n15618 ; n15618_not
g84743 not n15627 ; n15627_not
g84744 not n15636 ; n15636_not
g84745 not n15591 ; n15591_not
g84746 not n37506 ; n37506_not
g84747 not n15582 ; n15582_not
g84748 not n50376 ; n50376_not
g84749 not n15573 ; n15573_not
g84750 not n15564 ; n15564_not
g84751 not n15654 ; n15654_not
g84752 not n15555 ; n15555_not
g84753 not n15546 ; n15546_not
g84754 not n42429 ; n42429_not
g84755 not n16455 ; n16455_not
g84756 not n16464 ; n16464_not
g84757 not n32637 ; n32637_not
g84758 not n45129 ; n45129_not
g84759 not n16482 ; n16482_not
g84760 not n55218 ; n55218_not
g84761 not n32619 ; n32619_not
g84762 not n16509 ; n16509_not
g84763 not n16518 ; n16518_not
g84764 not n16527 ; n16527_not
g84765 not n16536 ; n16536_not
g84766 not n16545 ; n16545_not
g84767 not n47712 ; n47712_not
g84768 not n50466 ; n50466_not
g84769 not n16266 ; n16266_not
g84770 not n32682 ; n32682_not
g84771 not n16347 ; n16347_not
g84772 not n43059 ; n43059_not
g84773 not n47721 ; n47721_not
g84774 not n47136 ; n47136_not
g84775 not n32664 ; n32664_not
g84776 not n16392 ; n16392_not
g84777 not n50475 ; n50475_not
g84778 not n32655 ; n32655_not
g84779 not n16437 ; n16437_not
g84780 not n32556 ; n32556_not
g84781 not n16617 ; n16617_not
g84782 not n42474 ; n42474_not
g84783 not n42951 ; n42951_not
g84784 not n16626 ; n16626_not
g84785 not n32547 ; n32547_not
g84786 not n16635 ; n16635_not
g84787 not n42942 ; n42942_not
g84788 not n16644 ; n16644_not
g84789 not n32538 ; n32538_not
g84790 not n16653 ; n16653_not
g84791 not n42933 ; n42933_not
g84792 not n55236 ; n55236_not
g84793 not n32529 ; n32529_not
g84794 not n16662 ; n16662_not
g84795 not n16428 ; n16428_not
g84796 not n16554 ; n16554_not
g84797 not n16563 ; n16563_not
g84798 not n32592 ; n32592_not
g84799 not n50484 ; n50484_not
g84800 not n16572 ; n16572_not
g84801 not n16581 ; n16581_not
g84802 not n16473 ; n16473_not
g84803 not n32574 ; n32574_not
g84804 not n16590 ; n16590_not
g84805 not n42960 ; n42960_not
g84806 not n32565 ; n32565_not
g84807 not n47703 ; n47703_not
g84808 not n16608 ; n16608_not
g84809 not n15735 ; n15735_not
g84810 not n50439 ; n50439_not
g84811 not n43194 ; n43194_not
g84812 not n32628 ; n32628_not
g84813 not n15645 ; n15645_not
g84814 not n47730 ; n47730_not
g84815 not n43149 ; n43149_not
g84816 not n15690 ; n15690_not
g84817 not n50448 ; n50448_not
g84818 not n50457 ; n50457_not
g84819 not n32673 ; n32673_not
g84820 not n41592 ; n41592_not
g84821 not n18435 ; n18435_not
g84822 not n18444 ; n18444_not
g84823 not n42168 ; n42168_not
g84824 not n18462 ; n18462_not
g84825 not n41583 ; n41583_not
g84826 not n42159 ; n42159_not
g84827 not n31269 ; n31269_not
g84828 not n41952 ; n41952_not
g84829 not n41574 ; n41574_not
g84830 not n18480 ; n18480_not
g84831 not n18507 ; n18507_not
g84832 not n54309 ; n54309_not
g84833 not n47316 ; n47316_not
g84834 not n37920 ; n37920_not
g84835 not n41961 ; n41961_not
g84836 not n41565 ; n41565_not
g84837 not n18525 ; n18525_not
g84838 not n37911 ; n37911_not
g84839 not n18354 ; n18354_not
g84840 not n31575 ; n31575_not
g84841 not n47415 ; n47415_not
g84842 not n31476 ; n31476_not
g84843 not n41619 ; n41619_not
g84844 not n50628 ; n50628_not
g84845 not n18372 ; n18372_not
g84846 not n42195 ; n42195_not
g84847 not n31566 ; n31566_not
g84848 not n54291 ; n54291_not
g84849 not n31557 ; n31557_not
g84850 not n31485 ; n31485_not
g84851 not n18390 ; n18390_not
g84852 not n42186 ; n42186_not
g84853 not n31548 ; n31548_not
g84854 not n31494 ; n31494_not
g84855 not n18417 ; n18417_not
g84856 not n31539 ; n31539_not
g84857 not n42177 ; n42177_not
g84858 not n47406 ; n47406_not
g84859 not n41943 ; n41943_not
g84860 not n47370 ; n47370_not
g84861 not n17922 ; n17922_not
g84862 not n42087 ; n42087_not
g84863 not n17931 ; n17931_not
g84864 not n18543 ; n18543_not
g84865 not n17940 ; n17940_not
g84866 not n18534 ; n18534_not
g84867 not n42078 ; n42078_not
g84868 not n54345 ; n54345_not
g84869 not n41493 ; n41493_not
g84870 not n54354 ; n54354_not
g84871 not n41556 ; n41556_not
g84872 not n18552 ; n18552_not
g84873 not n41547 ; n41547_not
g84874 not n41538 ; n41538_not
g84875 not n18570 ; n18570_not
g84876 not n41529 ; n41529_not
g84877 not n31458 ; n31458_not
g84878 not n54336 ; n54336_not
g84879 not n37902 ; n37902_not
g84880 not n42096 ; n42096_not
g84881 not n50619 ; n50619_not
g84882 not n18156 ; n18156_not
g84883 not n54246 ; n54246_not
g84884 not n18165 ; n18165_not
g84885 not n47442 ; n47442_not
g84886 not n42276 ; n42276_not
g84887 not n18174 ; n18174_not
g84888 not n41691 ; n41691_not
g84889 not n31665 ; n31665_not
g84890 not n18183 ; n18183_not
g84891 not n18192 ; n18192_not
g84892 not n42267 ; n42267_not
g84893 not n31656 ; n31656_not
g84894 not n54255 ; n54255_not
g84895 not n41682 ; n41682_not
g84896 not n54264 ; n54264_not
g84897 not n18075 ; n18075_not
g84898 not n18084 ; n18084_not
g84899 not n18093 ; n18093_not
g84900 not n41871 ; n41871_not
g84901 not n41727 ; n41727_not
g84902 not n41718 ; n41718_not
g84903 not n42294 ; n42294_not
g84904 not n18129 ; n18129_not
g84905 not n17733 ; n17733_not
g84906 not n18138 ; n18138_not
g84907 not n41709 ; n41709_not
g84908 not n18147 ; n18147_not
g84909 not n42285 ; n42285_not
g84910 not n41916 ; n41916_not
g84911 not n41646 ; n41646_not
g84912 not n18282 ; n18282_not
g84913 not n18291 ; n18291_not
g84914 not n17643 ; n17643_not
g84915 not n41637 ; n41637_not
g84916 not n18309 ; n18309_not
g84917 not n47424 ; n47424_not
g84918 not n31593 ; n31593_not
g84919 not n18318 ; n18318_not
g84920 not n41628 ; n41628_not
g84921 not n31584 ; n31584_not
g84922 not n18345 ; n18345_not
g84923 not n42258 ; n42258_not
g84924 not n18219 ; n18219_not
g84925 not n31647 ; n31647_not
g84926 not n41673 ; n41673_not
g84927 not n18228 ; n18228_not
g84928 not n42249 ; n42249_not
g84929 not n31638 ; n31638_not
g84930 not n18237 ; n18237_not
g84931 not n47433 ; n47433_not
g84932 not n41664 ; n41664_not
g84933 not n18246 ; n18246_not
g84934 not n31629 ; n31629_not
g84935 not n31449 ; n31449_not
g84936 not n18255 ; n18255_not
g84937 not n18264 ; n18264_not
g84938 not n41907 ; n41907_not
g84939 not n41655 ; n41655_not
g84940 not n18273 ; n18273_not
g84941 not n54183 ; n54183_not
g84942 not n31188 ; n31188_not
g84943 not n19029 ; n19029_not
g84944 not n31179 ; n31179_not
g84945 not n19065 ; n19065_not
g84946 not n18930 ; n18930_not
g84947 not n41925 ; n41925_not
g84948 not n54228 ; n54228_not
g84949 not n18363 ; n18363_not
g84950 not n18840 ; n18840_not
g84951 not n41745 ; n41745_not
g84952 not n18831 ; n18831_not
g84953 not n41853 ; n41853_not
g84954 not n18822 ; n18822_not
g84955 not n30927 ; n30927_not
g84956 not n18813 ; n18813_not
g84957 not n18804 ; n18804_not
g84958 not n41754 ; n41754_not
g84959 not n41763 ; n41763_not
g84960 not n54093 ; n54093_not
g84961 not n41772 ; n41772_not
g84962 not n18750 ; n18750_not
g84963 not n41880 ; n41880_not
g84964 not n54138 ; n54138_not
g84965 not n18921 ; n18921_not
g84966 not n18912 ; n18912_not
g84967 not n18903 ; n18903_not
g84968 not n41862 ; n41862_not
g84969 not n19155 ; n19155_not
g84970 not n41736 ; n41736_not
g84971 not n18048 ; n18048_not
g84972 not n18057 ; n18057_not
g84973 not n31197 ; n31197_not
g84974 not n54363 ; n54363_not
g84975 not n18066 ; n18066_not
g84976 not n41457 ; n41457_not
g84977 not n41466 ; n41466_not
g84978 not n41475 ; n41475_not
g84979 not n50637 ; n50637_not
g84980 not n42069 ; n42069_not
g84981 not n41484 ; n41484_not
g84982 not n47361 ; n47361_not
g84983 not n18039 ; n18039_not
g84984 not n54381 ; n54381_not
g84985 not n18408 ; n18408_not
g84986 not n54273 ; n54273_not
g84987 not n18453 ; n18453_not
g84988 not n54318 ; n54318_not
g84989 not n47352 ; n47352_not
g84990 not n41970 ; n41970_not
g84991 not n42357 ; n42357_not
g84992 not n31818 ; n31818_not
g84993 not n31746 ; n31746_not
g84994 not n47271 ; n47271_not
g84995 not n50592 ; n50592_not
g84996 not n41826 ; n41826_not
g84997 not n31836 ; n31836_not
g84998 not n42393 ; n42393_not
g84999 not n42384 ; n42384_not
g85000 not n47451 ; n47451_not
g85001 not n31773 ; n31773_not
g85002 not n47460 ; n47460_not
g85003 not n42348 ; n42348_not
g85004 not n54219 ; n54219_not
g85005 not n31764 ; n31764_not
g85006 not n47505 ; n47505_not
g85007 not n42375 ; n42375_not
g85008 not n31845 ; n31845_not
g85009 not n42339 ; n42339_not
g85010 not n42366 ; n42366_not
g85011 not n31782 ; n31782_not
g85012 not n17823 ; n17823_not
g85013 not n54174 ; n54174_not
g85014 not n47514 ; n47514_not
g85015 not n31827 ; n31827_not
g85016 not n42682 ; n42682_not
g85017 not n38704 ; n38704_not
g85018 not n44581 ; n44581_not
g85019 not n42934 ; n42934_not
g85020 not n37129 ; n37129_not
g85021 not n38128 ; n38128_not
g85022 not n45841 ; n45841_not
g85023 not n37192 ; n37192_not
g85024 not n39703 ; n39703_not
g85025 not n45346 ; n45346_not
g85026 not n39262 ; n39262_not
g85027 not n36418 ; n36418_not
g85028 not n47263 ; n47263_not
g85029 not n45274 ; n45274_not
g85030 not n45472 ; n45472_not
g85031 not n37147 ; n37147_not
g85032 not n39154 ; n39154_not
g85033 not n41683 ; n41683_not
g85034 not n36409 ; n36409_not
g85035 not n48073 ; n48073_not
g85036 not n44590 ; n44590_not
g85037 not n46552 ; n46552_not
g85038 not n42376 ; n42376_not
g85039 not n43951 ; n43951_not
g85040 not n46084 ; n46084_not
g85041 not n41962 ; n41962_not
g85042 not n39172 ; n39172_not
g85043 not n44194 ; n44194_not
g85044 not n41296 ; n41296_not
g85045 not n39253 ; n39253_not
g85046 not n46075 ; n46075_not
g85047 not n41539 ; n41539_not
g85048 not n40765 ; n40765_not
g85049 not n46039 ; n46039_not
g85050 not n37633 ; n37633_not
g85051 not n46570 ; n46570_not
g85052 not n37165 ; n37165_not
g85053 not n45850 ; n45850_not
g85054 not n38380 ; n38380_not
g85055 not n39280 ; n39280_not
g85056 not n48712 ; n48712_not
g85057 not n43924 ; n43924_not
g85058 not n36436 ; n36436_not
g85059 not n46048 ; n46048_not
g85060 not n36364 ; n36364_not
g85061 not n41575 ; n41575_not
g85062 not n47092 ; n47092_not
g85063 not n42925 ; n42925_not
g85064 not n39163 ; n39163_not
g85065 not n41674 ; n41674_not
g85066 not n46066 ; n46066_not
g85067 not n47173 ; n47173_not
g85068 not n42943 ; n42943_not
g85069 not n38056 ; n38056_not
g85070 not n39271 ; n39271_not
g85071 not n46057 ; n46057_not
g85072 not n36427 ; n36427_not
g85073 not n44554 ; n44554_not
g85074 not n39235 ; n39235_not
g85075 not n41278 ; n41278_not
g85076 not n38137 ; n38137_not
g85077 not n44563 ; n44563_not
g85078 not n39217 ; n39217_not
g85079 not n43843 ; n43843_not
g85080 not n45166 ; n45166_not
g85081 not n36382 ; n36382_not
g85082 not n43267 ; n43267_not
g85083 not n45814 ; n45814_not
g85084 not n38272 ; n38272_not
g85085 not n39208 ; n39208_not
g85086 not n39712 ; n39712_not
g85087 not n43933 ; n43933_not
g85088 not n41557 ; n41557_not
g85089 not n41692 ; n41692_not
g85090 not n37174 ; n37174_not
g85091 not n37606 ; n37606_not
g85092 not n38371 ; n38371_not
g85093 not n36373 ; n36373_not
g85094 not n43276 ; n43276_not
g85095 not n39721 ; n39721_not
g85096 not n37156 ; n37156_not
g85097 not n46138 ; n46138_not
g85098 not n39730 ; n39730_not
g85099 not n42394 ; n42394_not
g85100 not n39145 ; n39145_not
g85101 not n42673 ; n42673_not
g85102 not n45805 ; n45805_not
g85103 not n46129 ; n46129_not
g85104 not n44419 ; n44419_not
g85105 not n46147 ; n46147_not
g85106 not n44086 ; n44086_not
g85107 not n40756 ; n40756_not
g85108 not n44482 ; n44482_not
g85109 not n46543 ; n46543_not
g85110 not n41548 ; n41548_not
g85111 not n46156 ; n46156_not
g85112 not n42385 ; n42385_not
g85113 not n37624 ; n37624_not
g85114 not n43942 ; n43942_not
g85115 not n46093 ; n46093_not
g85116 not n37183 ; n37183_not
g85117 not n37354 ; n37354_not
g85118 not n43249 ; n43249_not
g85119 not n48280 ; n48280_not
g85120 not n39244 ; n39244_not
g85121 not n36094 ; n36094_not
g85122 not n45391 ; n45391_not
g85123 not n36922 ; n36922_not
g85124 not n41287 ; n41287_not
g85125 not n41953 ; n41953_not
g85126 not n47272 ; n47272_not
g85127 not n36391 ; n36391_not
g85128 not n44077 ; n44077_not
g85129 not n39226 ; n39226_not
g85130 not n41566 ; n41566_not
g85131 not n48730 ; n48730_not
g85132 not n47740 ; n47740_not
g85133 not n41629 ; n41629_not
g85134 not n38407 ; n38407_not
g85135 not n39424 ; n39424_not
g85136 not n41836 ; n41836_not
g85137 not n42349 ; n42349_not
g85138 not n39064 ; n39064_not
g85139 not n45823 ; n45823_not
g85140 not n39055 ; n39055_not
g85141 not n39433 ; n39433_not
g85142 not n38416 ; n38416_not
g85143 not n38146 ; n38146_not
g85144 not n46651 ; n46651_not
g85145 not n46624 ; n46624_not
g85146 not n41458 ; n41458_not
g85147 not n39604 ; n39604_not
g85148 not n36049 ; n36049_not
g85149 not n37651 ; n37651_not
g85150 not n37642 ; n37642_not
g85151 not n36490 ; n36490_not
g85152 not n39406 ; n39406_not
g85153 not n39082 ; n39082_not
g85154 not n39415 ; n39415_not
g85155 not n43096 ; n43096_not
g85156 not n41449 ; n41449_not
g85157 not n43852 ; n43852_not
g85158 not n45490 ; n45490_not
g85159 not n47731 ; n47731_not
g85160 not n42367 ; n42367_not
g85161 not n38425 ; n38425_not
g85162 not n45733 ; n45733_not
g85163 not n36526 ; n36526_not
g85164 not n39019 ; n39019_not
g85165 not n43087 ; n43087_not
g85166 not n45337 ; n45337_not
g85167 not n39505 ; n39505_not
g85168 not n39514 ; n39514_not
g85169 not n43960 ; n43960_not
g85170 not n39523 ; n39523_not
g85171 not n47083 ; n47083_not
g85172 not n39442 ; n39442_not
g85173 not n47218 ; n47218_not
g85174 not n37336 ; n37336_not
g85175 not n46660 ; n46660_not
g85176 not n36508 ; n36508_not
g85177 not n39037 ; n39037_not
g85178 not n39451 ; n39451_not
g85179 not n48217 ; n48217_not
g85180 not n42466 ; n42466_not
g85181 not n46606 ; n46606_not
g85182 not n39460 ; n39460_not
g85183 not n45760 ; n45760_not
g85184 not n45751 ; n45751_not
g85185 not n43177 ; n43177_not
g85186 not n41656 ; n41656_not
g85187 not n45904 ; n45904_not
g85188 not n36454 ; n36454_not
g85189 not n39334 ; n39334_not
g85190 not n41494 ; n41494_not
g85191 not n43834 ; n43834_not
g85192 not n48703 ; n48703_not
g85193 not n39343 ; n39343_not
g85194 not n45940 ; n45940_not
g85195 not n41485 ; n41485_not
g85196 not n36067 ; n36067_not
g85197 not n42970 ; n42970_not
g85198 not n45931 ; n45931_not
g85199 not n47560 ; n47560_not
g85200 not n45922 ; n45922_not
g85201 not n41980 ; n41980_not
g85202 not n42952 ; n42952_not
g85203 not n41665 ; n41665_not
g85204 not n42448 ; n42448_not
g85205 not n44095 ; n44095_not
g85206 not n36445 ; n36445_not
g85207 not n39307 ; n39307_not
g85208 not n43186 ; n43186_not
g85209 not n45049 ; n45049_not
g85210 not n42961 ; n42961_not
g85211 not n39316 ; n39316_not
g85212 not n48046 ; n48046_not
g85213 not n48226 ; n48226_not
g85214 not n39325 ; n39325_not
g85215 not n43159 ; n43159_not
g85216 not n43708 ; n43708_not
g85217 not n39370 ; n39370_not
g85218 not n45913 ; n45913_not
g85219 not n39622 ; n39622_not
g85220 not n48118 ; n48118_not
g85221 not n41638 ; n41638_not
g85222 not n38263 ; n38263_not
g85223 not n42358 ; n42358_not
g85224 not n39613 ; n39613_not
g85225 not n41467 ; n41467_not
g85226 not n36481 ; n36481_not
g85227 not n39352 ; n39352_not
g85228 not n41647 ; n41647_not
g85229 not n39127 ; n39127_not
g85230 not n36463 ; n36463_not
g85231 not n47353 ; n47353_not
g85232 not n45247 ; n45247_not
g85233 not n36058 ; n36058_not
g85234 not n41476 ; n41476_not
g85235 not n44473 ; n44473_not
g85236 not n45481 ; n45481_not
g85237 not n37417 ; n37417_not
g85238 not n46615 ; n46615_not
g85239 not n39361 ; n39361_not
g85240 not n39109 ; n39109_not
g85241 not n36472 ; n36472_not
g85242 not n47182 ; n47182_not
g85243 not n37345 ; n37345_not
g85244 not n37381 ; n37381_not
g85245 not n38821 ; n38821_not
g85246 not n41863 ; n41863_not
g85247 not n36292 ; n36292_not
g85248 not n41791 ; n41791_not
g85249 not n39073 ; n39073_not
g85250 not n37372 ; n37372_not
g85251 not n37363 ; n37363_not
g85252 not n46327 ; n46327_not
g85253 not n38029 ; n38029_not
g85254 not n42790 ; n42790_not
g85255 not n45373 ; n45373_not
g85256 not n38812 ; n38812_not
g85257 not n45076 ; n45076_not
g85258 not n44518 ; n44518_not
g85259 not n47506 ; n47506_not
g85260 not n37408 ; n37408_not
g85261 not n41719 ; n41719_not
g85262 not n36283 ; n36283_not
g85263 not n46345 ; n46345_not
g85264 not n42808 ; n42808_not
g85265 not n38317 ; n38317_not
g85266 not n38830 ; n38830_not
g85267 not n46435 ; n46435_not
g85268 not n37390 ; n37390_not
g85269 not n46336 ; n46336_not
g85270 not n47533 ; n47533_not
g85271 not n48253 ; n48253_not
g85272 not n42781 ; n42781_not
g85273 not n47137 ; n47137_not
g85274 not n37516 ; n37516_not
g85275 not n48064 ; n48064_not
g85276 not n38335 ; n38335_not
g85277 not n46453 ; n46453_not
g85278 not n40747 ; n40747_not
g85279 not n45715 ; n45715_not
g85280 not n41773 ; n41773_not
g85281 not n43861 ; n43861_not
g85282 not n38038 ; n38038_not
g85283 not n46318 ; n46318_not
g85284 not n36157 ; n36157_not
g85285 not n38326 ; n38326_not
g85286 not n45706 ; n45706_not
g85287 not n44059 ; n44059_not
g85288 not n38290 ; n38290_not
g85289 not n44527 ; n44527_not
g85290 not n41782 ; n41782_not
g85291 not n41872 ; n41872_not
g85292 not n47335 ; n47335_not
g85293 not n36148 ; n36148_not
g85294 not n46309 ; n46309_not
g85295 not n38803 ; n38803_not
g85296 not n42871 ; n42871_not
g85297 not n37453 ; n37453_not
g85298 not n45067 ; n45067_not
g85299 not n46363 ; n46363_not
g85300 not n41818 ; n41818_not
g85301 not n41746 ; n41746_not
g85302 not n47524 ; n47524_not
g85303 not n37435 ; n37435_not
g85304 not n46372 ; n46372_not
g85305 not n41827 ; n41827_not
g85306 not n39028 ; n39028_not
g85307 not n41737 ; n41737_not
g85308 not n42862 ; n42862_not
g85309 not n37444 ; n37444_not
g85310 not n47515 ; n47515_not
g85311 not n48802 ; n48802_not
g85312 not n41764 ; n41764_not
g85313 not n45463 ; n45463_not
g85314 not n42853 ; n42853_not
g85315 not n46390 ; n46390_not
g85316 not n48244 ; n48244_not
g85317 not n36517 ; n36517_not
g85318 not n41755 ; n41755_not
g85319 not n36256 ; n36256_not
g85320 not n41845 ; n41845_not
g85321 not n42844 ; n42844_not
g85322 not n37426 ; n37426_not
g85323 not n43195 ; n43195_not
g85324 not n41728 ; n41728_not
g85325 not n41809 ; n41809_not
g85326 not n46354 ; n46354_not
g85327 not n36274 ; n36274_not
g85328 not n38920 ; n38920_not
g85329 not n37471 ; n37471_not
g85330 not n43807 ; n43807_not
g85331 not n42817 ; n42817_not
g85332 not n45364 ; n45364_not
g85333 not n46417 ; n46417_not
g85334 not n42835 ; n42835_not
g85335 not n47911 ; n47911_not
g85336 not n38902 ; n38902_not
g85337 not n38308 ; n38308_not
g85338 not n37066 ; n37066_not
g85339 not n44509 ; n44509_not
g85340 not n36265 ; n36265_not
g85341 not n42880 ; n42880_not
g85342 not n42826 ; n42826_not
g85343 not n46408 ; n46408_not
g85344 not n38911 ; n38911_not
g85345 not n46219 ; n46219_not
g85346 not n41917 ; n41917_not
g85347 not n38731 ; n38731_not
g85348 not n48271 ; n48271_not
g85349 not n37273 ; n37273_not
g85350 not n48037 ; n48037_not
g85351 not n38083 ; n38083_not
g85352 not n38281 ; n38281_not
g85353 not n47821 ; n47821_not
g85354 not n39631 ; n39631_not
g85355 not n38362 ; n38362_not
g85356 not n37264 ; n37264_not
g85357 not n46507 ; n46507_not
g85358 not n36346 ; n36346_not
g85359 not n42736 ; n42736_not
g85360 not n44068 ; n44068_not
g85361 not n41908 ; n41908_not
g85362 not n38740 ; n38740_not
g85363 not n47128 ; n47128_not
g85364 not n37282 ; n37282_not
g85365 not n39118 ; n39118_not
g85366 not n42916 ; n42916_not
g85367 not n42727 ; n42727_not
g85368 not n46228 ; n46228_not
g85369 not n46174 ; n46174_not
g85370 not n42709 ; n42709_not
g85371 not n37228 ; n37228_not
g85372 not n38713 ; n38713_not
g85373 not n45094 ; n45094_not
g85374 not n47290 ; n47290_not
g85375 not n42691 ; n42691_not
g85376 not n46165 ; n46165_not
g85377 not n37219 ; n37219_not
g85378 not n41584 ; n41584_not
g85379 not n46525 ; n46525_not
g85380 not n47551 ; n47551_not
g85381 not n41593 ; n41593_not
g85382 not n38722 ; n38722_not
g85383 not n41935 ; n41935_not
g85384 not n37255 ; n37255_not
g85385 not n37561 ; n37561_not
g85386 not n42718 ; n42718_not
g85387 not n46192 ; n46192_not
g85388 not n37246 ; n37246_not
g85389 not n36931 ; n36931_not
g85390 not n46183 ; n46183_not
g85391 not n37237 ; n37237_not
g85392 not n47803 ; n47803_not
g85393 not n36355 ; n36355_not
g85394 not n46282 ; n46282_not
g85395 not n43717 ; n43717_not
g85396 not n47542 ; n47542_not
g85397 not n36319 ; n36319_not
g85398 not n45175 ; n45175_not
g85399 not n42907 ; n42907_not
g85400 not n45382 ; n45382_not
g85401 not n39541 ; n39541_not
g85402 not n46273 ; n46273_not
g85403 not n42754 ; n42754_not
g85404 not n37318 ; n37318_not
g85405 not n36139 ; n36139_not
g85406 not n45355 ; n45355_not
g85407 not n38344 ; n38344_not
g85408 not n46291 ; n46291_not
g85409 not n42772 ; n42772_not
g85410 not n47236 ; n47236_not
g85411 not n37327 ; n37327_not
g85412 not n45724 ; n45724_not
g85413 not n46462 ; n46462_not
g85414 not n41890 ; n41890_not
g85415 not n42763 ; n42763_not
g85416 not n39532 ; n39532_not
g85417 not n42745 ; n42745_not
g85418 not n46246 ; n46246_not
g85419 not n36940 ; n36940_not
g85420 not n37534 ; n37534_not
g85421 not n37291 ; n37291_not
g85422 not n47308 ; n47308_not
g85423 not n47227 ; n47227_not
g85424 not n47155 ; n47155_not
g85425 not n37507 ; n37507_not
g85426 not n46237 ; n46237_not
g85427 not n37543 ; n37543_not
g85428 not n38353 ; n38353_not
g85429 not n36328 ; n36328_not
g85430 not n46264 ; n46264_not
g85431 not n48262 ; n48262_not
g85432 not n46255 ; n46255_not
g85433 not n37309 ; n37309_not
g85434 not n47317 ; n47317_not
g85435 not n46480 ; n46480_not
g85436 not n36337 ; n36337_not
g85437 not n48235 ; n48235_not
g85438 not n48109 ; n48109_not
g85439 not n38065 ; n38065_not
g85440 not n45544 ; n45544_not
g85441 not n44374 ; n44374_not
g85442 not n42556 ; n42556_not
g85443 not n45085 ; n45085_not
g85444 not n47425 ; n47425_not
g85445 not n48424 ; n48424_not
g85446 not n43753 ; n43753_not
g85447 not n47623 ; n47623_not
g85448 not n42169 ; n42169_not
g85449 not n38515 ; n38515_not
g85450 not n42565 ; n42565_not
g85451 not n36814 ; n36814_not
g85452 not n38155 ; n38155_not
g85453 not n40549 ; n40549_not
g85454 not n40486 ; n40486_not
g85455 not n45283 ; n45283_not
g85456 not n42187 ; n42187_not
g85457 not n38650 ; n38650_not
g85458 not n45553 ; n45553_not
g85459 not n40495 ; n40495_not
g85460 not n44293 ; n44293_not
g85461 not n43744 ; n43744_not
g85462 not n36805 ; n36805_not
g85463 not n48172 ; n48172_not
g85464 not n47191 ; n47191_not
g85465 not n48433 ; n48433_not
g85466 not n45436 ; n45436_not
g85467 not n42178 ; n42178_not
g85468 not n45229 ; n45229_not
g85469 not n38191 ; n38191_not
g85470 not n38614 ; n38614_not
g85471 not n36823 ; n36823_not
g85472 not n44437 ; n44437_not
g85473 not n38524 ; n38524_not
g85474 not n38182 ; n38182_not
g85475 not n40576 ; n40576_not
g85476 not n47434 ; n47434_not
g85477 not n48145 ; n48145_not
g85478 not n45454 ; n45454_not
g85479 not n45535 ; n45535_not
g85480 not n42583 ; n42583_not
g85481 not n40585 ; n40585_not
g85482 not n38605 ; n38605_not
g85483 not n48406 ; n48406_not
g85484 not n38632 ; n38632_not
g85485 not n41395 ; n41395_not
g85486 not n44356 ; n44356_not
g85487 not n38164 ; n38164_not
g85488 not n40558 ; n40558_not
g85489 not n48415 ; n48415_not
g85490 not n38173 ; n38173_not
g85491 not n42574 ; n42574_not
g85492 not n44149 ; n44149_not
g85493 not n40567 ; n40567_not
g85494 not n48181 ; n48181_not
g85495 not n44266 ; n44266_not
g85496 not n47281 ; n47281_not
g85497 not n47614 ; n47614_not
g85498 not n44275 ; n44275_not
g85499 not n42196 ; n42196_not
g85500 not n45562 ; n45562_not
g85501 not n42529 ; n42529_not
g85502 not n38218 ; n38218_not
g85503 not n44239 ; n44239_not
g85504 not n42259 ; n42259_not
g85505 not n44248 ; n44248_not
g85506 not n47461 ; n47461_not
g85507 not n44383 ; n44383_not
g85508 not n44257 ; n44257_not
g85509 not n43726 ; n43726_not
g85510 not n46426 ; n46426_not
g85511 not n36607 ; n36607_not
g85512 not n48451 ; n48451_not
g85513 not n40477 ; n40477_not
g85514 not n47047 ; n47047_not
g85515 not n48019 ; n48019_not
g85516 not n41926 ; n41926_not
g85517 not n48442 ; n48442_not
g85518 not n37093 ; n37093_not
g85519 not n38623 ; n38623_not
g85520 not n40459 ; n40459_not
g85521 not n48028 ; n48028_not
g85522 not n48460 ; n48460_not
g85523 not n48136 ; n48136_not
g85524 not n44284 ; n44284_not
g85525 not n40468 ; n40468_not
g85526 not n47416 ; n47416_not
g85527 not n42538 ; n42538_not
g85528 not n38209 ; n38209_not
g85529 not n42619 ; n42619_not
g85530 not n36562 ; n36562_not
g85531 not n47029 ; n47029_not
g85532 not n48334 ; n48334_not
g85533 not n41881 ; n41881_not
g85534 not n40396 ; n40396_not
g85535 not n38560 ; n38560_not
g85536 not n45526 ; n45526_not
g85537 not n47443 ; n47443_not
g85538 not n47452 ; n47452_not
g85539 not n48343 ; n48343_not
g85540 not n47641 ; n47641_not
g85541 not n42286 ; n42286_not
g85542 not n37084 ; n37084_not
g85543 not n40729 ; n40729_not
g85544 not n40819 ; n40819_not
g85545 not n40837 ; n40837_not
g85546 not n40297 ; n40297_not
g85547 not n38542 ; n38542_not
g85548 not n40288 ; n40288_not
g85549 not n47038 ; n47038_not
g85550 not n37048 ; n37048_not
g85551 not n36553 ; n36553_not
g85552 not n42646 ; n42646_not
g85553 not n48325 ; n48325_not
g85554 not n40855 ; n40855_not
g85555 not n40774 ; n40774_not
g85556 not n42628 ; n42628_not
g85557 not n40387 ; n40387_not
g85558 not n40378 ; n40378_not
g85559 not n40369 ; n40369_not
g85560 not n43915 ; n43915_not
g85561 not n48154 ; n48154_not
g85562 not n43906 ; n43906_not
g85563 not n44347 ; n44347_not
g85564 not n40792 ; n40792_not
g85565 not n45517 ; n45517_not
g85566 not n45256 ; n45256_not
g85567 not n42295 ; n42295_not
g85568 not n45292 ; n45292_not
g85569 not n40864 ; n40864_not
g85570 not n47632 ; n47632_not
g85571 not n38227 ; n38227_not
g85572 not n37039 ; n37039_not
g85573 not n41368 ; n41368_not
g85574 not n45508 ; n45508_not
g85575 not n45445 ; n45445_not
g85576 not n36841 ; n36841_not
g85577 not n44338 ; n44338_not
g85578 not n47650 ; n47650_not
g85579 not n38236 ; n38236_not
g85580 not n40675 ; n40675_not
g85581 not n44329 ; n44329_not
g85582 not n37075 ; n37075_not
g85583 not n36832 ; n36832_not
g85584 not n37552 ; n37552_not
g85585 not n40099 ; n40099_not
g85586 not n41377 ; n41377_not
g85587 not n48082 ; n48082_not
g85588 not n43771 ; n43771_not
g85589 not n40594 ; n40594_not
g85590 not n40657 ; n40657_not
g85591 not n42088 ; n42088_not
g85592 not n40666 ; n40666_not
g85593 not n42277 ; n42277_not
g85594 not n40684 ; n40684_not
g85595 not n42079 ; n42079_not
g85596 not n38254 ; n38254_not
g85597 not n37462 ; n37462_not
g85598 not n47902 ; n47902_not
g85599 not n48352 ; n48352_not
g85600 not n48163 ; n48163_not
g85601 not n48370 ; n48370_not
g85602 not n36850 ; n36850_not
g85603 not n42268 ; n42268_not
g85604 not n40639 ; n40639_not
g85605 not n45265 ; n45265_not
g85606 not n42097 ; n42097_not
g85607 not n38245 ; n38245_not
g85608 not n48361 ; n48361_not
g85609 not n40279 ; n40279_not
g85610 not n45607 ; n45607_not
g85611 not n47380 ; n47380_not
g85612 not n36634 ; n36634_not
g85613 not n38119 ; n38119_not
g85614 not n45328 ; n45328_not
g85615 not n48091 ; n48091_not
g85616 not n48307 ; n48307_not
g85617 not n47371 ; n47371_not
g85618 not n45625 ; n45625_not
g85619 not n36616 ; n36616_not
g85620 not n45616 ; n45616_not
g85621 not n38074 ; n38074_not
g85622 not n45139 ; n45139_not
g85623 not n38452 ; n38452_not
g85624 not n47326 ; n47326_not
g85625 not n47146 ; n47146_not
g85626 not n44491 ; n44491_not
g85627 not n46822 ; n46822_not
g85628 not n43762 ; n43762_not
g85629 not n36229 ; n36229_not
g85630 not n38533 ; n38533_not
g85631 not n45157 ; n45157_not
g85632 not n44392 ; n44392_not
g85633 not n38461 ; n38461_not
g85634 not n36643 ; n36643_not
g85635 not n46804 ; n46804_not
g85636 not n45418 ; n45418_not
g85637 not n47704 ; n47704_not
g85638 not n46813 ; n46813_not
g85639 not n36661 ; n36661_not
g85640 not n46705 ; n46705_not
g85641 not n38434 ; n38434_not
g85642 not n36913 ; n36913_not
g85643 not n46714 ; n46714_not
g85644 not n42475 ; n42475_not
g85645 not n48208 ; n48208_not
g85646 not n36571 ; n36571_not
g85647 not n46723 ; n46723_not
g85648 not n48640 ; n48640_not
g85649 not n36544 ; n36544_not
g85650 not n43069 ; n43069_not
g85651 not n47362 ; n47362_not
g85652 not n45409 ; n45409_not
g85653 not n47722 ; n47722_not
g85654 not n40189 ; n40189_not
g85655 not n45652 ; n45652_not
g85656 not n38443 ; n38443_not
g85657 not n44464 ; n44464_not
g85658 not n47713 ; n47713_not
g85659 not n42439 ; n42439_not
g85660 not n47470 ; n47470_not
g85661 not n45643 ; n45643_not
g85662 not n37138 ; n37138_not
g85663 not n45634 ; n45634_not
g85664 not n47074 ; n47074_not
g85665 not n48622 ; n48622_not
g85666 not n46732 ; n46732_not
g85667 not n38470 ; n38470_not
g85668 not n48613 ; n48613_not
g85669 not n44185 ; n44185_not
g85670 not n46741 ; n46741_not
g85671 not n45670 ; n45670_not
g85672 not n46561 ; n46561_not
g85673 not n46750 ; n46750_not
g85674 not n44536 ; n44536_not
g85675 not n45661 ; n45661_not
g85676 not n46471 ; n46471_not
g85677 not n36742 ; n36742_not
g85678 not n44428 ; n44428_not
g85679 not n44176 ; n44176_not
g85680 not n46912 ; n46912_not
g85681 not n48505 ; n48505_not
g85682 not n45571 ; n45571_not
g85683 not n48316 ; n48316_not
g85684 not n45184 ; n45184_not
g85685 not n36751 ; n36751_not
g85686 not n44158 ; n44158_not
g85687 not n47812 ; n47812_not
g85688 not n48514 ; n48514_not
g85689 not n46903 ; n46903_not
g85690 not n44167 ; n44167_not
g85691 not n47605 ; n47605_not
g85692 not n46930 ; n46930_not
g85693 not n36760 ; n36760_not
g85694 not n47407 ; n47407_not
g85695 not n46921 ; n46921_not
g85696 not n40198 ; n40198_not
g85697 not n47056 ; n47056_not
g85698 not n45427 ; n45427_not
g85699 not n36706 ; n36706_not
g85700 not n42493 ; n42493_not
g85701 not n47245 ; n47245_not
g85702 not n42484 ; n42484_not
g85703 not n46840 ; n46840_not
g85704 not n36652 ; n36652_not
g85705 not n48127 ; n48127_not
g85706 not n41386 ; n41386_not
g85707 not n41971 ; n41971_not
g85708 not n47065 ; n47065_not
g85709 not n46381 ; n46381_not
g85710 not n48550 ; n48550_not
g85711 not n46516 ; n46516_not
g85712 not n46831 ; n46831_not
g85713 not n48532 ; n48532_not
g85714 not n43681 ; n43681_not
g85715 not n48541 ; n48541_not
g85716 not n36904 ; n36904_not
g85717 not n36724 ; n36724_not
g85718 not n48523 ; n48523_not
g85719 not n43816 ; n43816_not
g85720 not n36733 ; n36733_not
g85721 not n45580 ; n45580_not
g85722 not n36715 ; n36715_not
g85723 not n45319 ; n45319_not
g85724 not n44446 ; n44446_not
g85725 not n48190 ; n48190_not
g85726 not n31792 ; n31792_not
g85727 not n23836 ; n23836_not
g85728 not n17428 ; n17428_not
g85729 not n26914 ; n26914_not
g85730 not n17194 ; n17194_not
g85731 not n17437 ; n17437_not
g85732 not n50593 ; n50593_not
g85733 not n17446 ; n17446_not
g85734 not n17455 ; n17455_not
g85735 not n23818 ; n23818_not
g85736 not n17464 ; n17464_not
g85737 not n17473 ; n17473_not
g85738 not n23809 ; n23809_not
g85739 not n17482 ; n17482_not
g85740 not n31774 ; n31774_not
g85741 not n54940 ; n54940_not
g85742 not n17491 ; n17491_not
g85743 not n54922 ; n54922_not
g85744 not n17356 ; n17356_not
g85745 not n17365 ; n17365_not
g85746 not n17374 ; n17374_not
g85747 not n31846 ; n31846_not
g85748 not n17383 ; n17383_not
g85749 not n27760 ; n27760_not
g85750 not n17392 ; n17392_not
g85751 not n17077 ; n17077_not
g85752 not n31837 ; n31837_not
g85753 not n51196 ; n51196_not
g85754 not n17068 ; n17068_not
g85755 not n31828 ; n31828_not
g85756 not n51880 ; n51880_not
g85757 not n17419 ; n17419_not
g85758 not n17059 ; n17059_not
g85759 not n31819 ; n31819_not
g85760 not n17572 ; n17572_not
g85761 not n17581 ; n17581_not
g85762 not n51259 ; n51259_not
g85763 not n54067 ; n54067_not
g85764 not n23773 ; n23773_not
g85765 not n31666 ; n31666_not
g85766 not n17590 ; n17590_not
g85767 not n54058 ; n54058_not
g85768 not n31657 ; n31657_not
g85769 not n31648 ; n31648_not
g85770 not n54049 ; n54049_not
g85771 not n31639 ; n31639_not
g85772 not n23764 ; n23764_not
g85773 not n17608 ; n17608_not
g85774 not n16951 ; n16951_not
g85775 not n52726 ; n52726_not
g85776 not n17626 ; n17626_not
g85777 not n31459 ; n31459_not
g85778 not n31594 ; n31594_not
g85779 not n54931 ; n54931_not
g85780 not n31783 ; n31783_not
g85781 not n17509 ; n17509_not
g85782 not n17518 ; n17518_not
g85783 not n23791 ; n23791_not
g85784 not n31756 ; n31756_not
g85785 not n17527 ; n17527_not
g85786 not n51862 ; n51862_not
g85787 not n17536 ; n17536_not
g85788 not n51853 ; n51853_not
g85789 not n17545 ; n17545_not
g85790 not n31738 ; n31738_not
g85791 not n31729 ; n31729_not
g85792 not n17554 ; n17554_not
g85793 not n54085 ; n54085_not
g85794 not n27805 ; n27805_not
g85795 not n17563 ; n17563_not
g85796 not n54094 ; n54094_not
g85797 not n31693 ; n31693_not
g85798 not n27724 ; n27724_not
g85799 not n23908 ; n23908_not
g85800 not n51169 ; n51169_not
g85801 not n27733 ; n27733_not
g85802 not n52546 ; n52546_not
g85803 not n31936 ; n31936_not
g85804 not n55084 ; n55084_not
g85805 not n17149 ; n17149_not
g85806 not n17158 ; n17158_not
g85807 not n31927 ; n31927_not
g85808 not n51178 ; n51178_not
g85809 not n55075 ; n55075_not
g85810 not n31918 ; n31918_not
g85811 not n26932 ; n26932_not
g85812 not n17176 ; n17176_not
g85813 not n16528 ; n16528_not
g85814 not n31909 ; n31909_not
g85815 not n27742 ; n27742_not
g85816 not n52537 ; n52537_not
g85817 not n50557 ; n50557_not
g85818 not n23935 ; n23935_not
g85819 not n23863 ; n23863_not
g85820 not n55147 ; n55147_not
g85821 not n51907 ; n51907_not
g85822 not n23926 ; n23926_not
g85823 not n31963 ; n31963_not
g85824 not n27706 ; n27706_not
g85825 not n55129 ; n55129_not
g85826 not n23872 ; n23872_not
g85827 not n23917 ; n23917_not
g85828 not n26950 ; n26950_not
g85829 not n31954 ; n31954_not
g85830 not n27715 ; n27715_not
g85831 not n50566 ; n50566_not
g85832 not n26941 ; n26941_not
g85833 not n17086 ; n17086_not
g85834 not n31945 ; n31945_not
g85835 not n17275 ; n17275_not
g85836 not n31873 ; n31873_not
g85837 not n17284 ; n17284_not
g85838 not n23854 ; n23854_not
g85839 not n17293 ; n17293_not
g85840 not n27751 ; n27751_not
g85841 not n55039 ; n55039_not
g85842 not n31864 ; n31864_not
g85843 not n17329 ; n17329_not
g85844 not n31747 ; n31747_not
g85845 not n50584 ; n50584_not
g85846 not n17338 ; n17338_not
g85847 not n31855 ; n31855_not
g85848 not n17347 ; n17347_not
g85849 not n23881 ; n23881_not
g85850 not n50188 ; n50188_not
g85851 not n55057 ; n55057_not
g85852 not n17167 ; n17167_not
g85853 not n31891 ; n31891_not
g85854 not n17239 ; n17239_not
g85855 not n51187 ; n51187_not
g85856 not n50575 ; n50575_not
g85857 not n17248 ; n17248_not
g85858 not n17257 ; n17257_not
g85859 not n31882 ; n31882_not
g85860 not n17266 ; n17266_not
g85861 not n53086 ; n53086_not
g85862 not n30919 ; n30919_not
g85863 not n53905 ; n53905_not
g85864 not n22909 ; n22909_not
g85865 not n51385 ; n51385_not
g85866 not n23395 ; n23395_not
g85867 not n17815 ; n17815_not
g85868 not n51772 ; n51772_not
g85869 not n53095 ; n53095_not
g85870 not n22918 ; n22918_not
g85871 not n53860 ; n53860_not
g85872 not n51394 ; n51394_not
g85873 not n23386 ; n23386_not
g85874 not n53851 ; n53851_not
g85875 not n22927 ; n22927_not
g85876 not n23377 ; n23377_not
g85877 not n51763 ; n51763_not
g85878 not n53842 ; n53842_not
g85879 not n23476 ; n23476_not
g85880 not n50692 ; n50692_not
g85881 not n54166 ; n54166_not
g85882 not n53941 ; n53941_not
g85883 not n27931 ; n27931_not
g85884 not n22873 ; n22873_not
g85885 not n53932 ; n53932_not
g85886 not n30946 ; n30946_not
g85887 not n23467 ; n23467_not
g85888 not n51376 ; n51376_not
g85889 not n22882 ; n22882_not
g85890 not n54175 ; n54175_not
g85891 not n53923 ; n53923_not
g85892 not n27940 ; n27940_not
g85893 not n23458 ; n23458_not
g85894 not n54184 ; n54184_not
g85895 not n23449 ; n23449_not
g85896 not n53914 ; n53914_not
g85897 not n17833 ; n17833_not
g85898 not n30928 ; n30928_not
g85899 not n17824 ; n17824_not
g85900 not n30748 ; n30748_not
g85901 not n53806 ; n53806_not
g85902 not n23287 ; n23287_not
g85903 not n17725 ; n17725_not
g85904 not n30685 ; n30685_not
g85905 not n23278 ; n23278_not
g85906 not n30478 ; n30478_not
g85907 not n52492 ; n52492_not
g85908 not n23269 ; n23269_not
g85909 not n51448 ; n51448_not
g85910 not n30487 ; n30487_not
g85911 not n30496 ; n30496_not
g85912 not n23197 ; n23197_not
g85913 not n50098 ; n50098_not
g85914 not n54256 ; n54256_not
g85915 not n23188 ; n23188_not
g85916 not n23179 ; n23179_not
g85917 not n23368 ; n23368_not
g85918 not n17770 ; n17770_not
g85919 not n54229 ; n54229_not
g85920 not n53833 ; n53833_not
g85921 not n23359 ; n23359_not
g85922 not n50719 ; n50719_not
g85923 not n53824 ; n53824_not
g85924 not n22954 ; n22954_not
g85925 not n22963 ; n22963_not
g85926 not n50728 ; n50728_not
g85927 not n53815 ; n53815_not
g85928 not n22972 ; n22972_not
g85929 not n51439 ; n51439_not
g85930 not n17743 ; n17743_not
g85931 not n23296 ; n23296_not
g85932 not n30757 ; n30757_not
g85933 not n51745 ; n51745_not
g85934 not n17734 ; n17734_not
g85935 not n31369 ; n31369_not
g85936 not n31378 ; n31378_not
g85937 not n17680 ; n17680_not
g85938 not n27841 ; n27841_not
g85939 not n51286 ; n51286_not
g85940 not n31387 ; n31387_not
g85941 not n52528 ; n52528_not
g85942 not n31396 ; n31396_not
g85943 not n17707 ; n17707_not
g85944 not n23683 ; n23683_not
g85945 not n27850 ; n27850_not
g85946 not n31189 ; n31189_not
g85947 not n31198 ; n31198_not
g85948 not n50638 ; n50638_not
g85949 not n51295 ; n51295_not
g85950 not n23674 ; n23674_not
g85951 not n31297 ; n31297_not
g85952 not n31288 ; n31288_not
g85953 not n31279 ; n31279_not
g85954 not n17617 ; n17617_not
g85955 not n31585 ; n31585_not
g85956 not n23746 ; n23746_not
g85957 not n17635 ; n17635_not
g85958 not n31576 ; n31576_not
g85959 not n17644 ; n17644_not
g85960 not n31567 ; n31567_not
g85961 not n27823 ; n27823_not
g85962 not n50629 ; n50629_not
g85963 not n31558 ; n31558_not
g85964 not n31486 ; n31486_not
g85965 not n31549 ; n31549_not
g85966 not n51268 ; n51268_not
g85967 not n31495 ; n31495_not
g85968 not n17662 ; n17662_not
g85969 not n51277 ; n51277_not
g85970 not n51835 ; n51835_not
g85971 not n23728 ; n23728_not
g85972 not n23719 ; n23719_not
g85973 not n31468 ; n31468_not
g85974 not n23557 ; n23557_not
g85975 not n54139 ; n54139_not
g85976 not n51790 ; n51790_not
g85977 not n22828 ; n22828_not
g85978 not n51358 ; n51358_not
g85979 not n23548 ; n23548_not
g85980 not n22837 ; n22837_not
g85981 not n50674 ; n50674_not
g85982 not n23539 ; n23539_not
g85983 not n27913 ; n27913_not
g85984 not n30766 ; n30766_not
g85985 not n53068 ; n53068_not
g85986 not n17842 ; n17842_not
g85987 not n51367 ; n51367_not
g85988 not n23494 ; n23494_not
g85989 not n17860 ; n17860_not
g85990 not n50683 ; n50683_not
g85991 not n22864 ; n22864_not
g85992 not n23485 ; n23485_not
g85993 not n53077 ; n53077_not
g85994 not n30973 ; n30973_not
g85995 not n53950 ; n53950_not
g85996 not n30964 ; n30964_not
g85997 not n23656 ; n23656_not
g85998 not n23638 ; n23638_not
g85999 not n17752 ; n17752_not
g86000 not n51817 ; n51817_not
g86001 not n30937 ; n30937_not
g86002 not n31099 ; n31099_not
g86003 not n51808 ; n51808_not
g86004 not n23629 ; n23629_not
g86005 not n50647 ; n50647_not
g86006 not n51349 ; n51349_not
g86007 not n50656 ; n50656_not
g86008 not n53059 ; n53059_not
g86009 not n23593 ; n23593_not
g86010 not n23584 ; n23584_not
g86011 not n23575 ; n23575_not
g86012 not n22819 ; n22819_not
g86013 not n30982 ; n30982_not
g86014 not n23566 ; n23566_not
g86015 not n50665 ; n50665_not
g86016 not n15655 ; n15655_not
g86017 not n52618 ; n52618_not
g86018 not n32746 ; n32746_not
g86019 not n15862 ; n15862_not
g86020 not n15646 ; n15646_not
g86021 not n32755 ; n32755_not
g86022 not n27508 ; n27508_not
g86023 not n32764 ; n32764_not
g86024 not n15637 ; n15637_not
g86025 not n32773 ; n32773_not
g86026 not n27517 ; n27517_not
g86027 not n32782 ; n32782_not
g86028 not n16249 ; n16249_not
g86029 not n32791 ; n32791_not
g86030 not n16258 ; n16258_not
g86031 not n24196 ; n24196_not
g86032 not n15619 ; n15619_not
g86033 not n32809 ; n32809_not
g86034 not n32818 ; n32818_not
g86035 not n33097 ; n33097_not
g86036 not n24259 ; n24259_not
g86037 not n16168 ; n16168_not
g86038 not n33088 ; n33088_not
g86039 not n50287 ; n50287_not
g86040 not n27076 ; n27076_not
g86041 not n16177 ; n16177_not
g86042 not n33079 ; n33079_not
g86043 not n27481 ; n27481_not
g86044 not n16186 ; n16186_not
g86045 not n23692 ; n23692_not
g86046 not n27490 ; n27490_not
g86047 not n50395 ; n50395_not
g86048 not n32728 ; n32728_not
g86049 not n16195 ; n16195_not
g86050 not n55246 ; n55246_not
g86051 not n32737 ; n32737_not
g86052 not n27067 ; n27067_not
g86053 not n32953 ; n32953_not
g86054 not n16375 ; n16375_not
g86055 not n55291 ; n55291_not
g86056 not n16087 ; n16087_not
g86057 not n32881 ; n32881_not
g86058 not n16384 ; n16384_not
g86059 not n32944 ; n32944_not
g86060 not n16078 ; n16078_not
g86061 not n27544 ; n27544_not
g86062 not n32890 ; n32890_not
g86063 not n16069 ; n16069_not
g86064 not n24178 ; n24178_not
g86065 not n32908 ; n32908_not
g86066 not n16429 ; n16429_not
g86067 not n55282 ; n55282_not
g86068 not n15970 ; n15970_not
g86069 not n32926 ; n32926_not
g86070 not n16447 ; n16447_not
g86071 not n15961 ; n15961_not
g86072 not n32917 ; n32917_not
g86073 not n32584 ; n32584_not
g86074 not n15952 ; n15952_not
g86075 not n32593 ; n32593_not
g86076 not n16267 ; n16267_not
g86077 not n32827 ; n32827_not
g86078 not n16276 ; n16276_not
g86079 not n27526 ; n27526_not
g86080 not n32836 ; n32836_not
g86081 not n32971 ; n32971_not
g86082 not n16285 ; n16285_not
g86083 not n16294 ; n16294_not
g86084 not n32845 ; n32845_not
g86085 not n24187 ; n24187_not
g86086 not n32854 ; n32854_not
g86087 not n16339 ; n16339_not
g86088 not n16159 ; n16159_not
g86089 not n32863 ; n32863_not
g86090 not n16357 ; n16357_not
g86091 not n27535 ; n27535_not
g86092 not n52906 ; n52906_not
g86093 not n50278 ; n50278_not
g86094 not n16096 ; n16096_not
g86095 not n32872 ; n32872_not
g86096 not n33277 ; n33277_not
g86097 not n24349 ; n24349_not
g86098 not n33259 ; n33259_not
g86099 not n27373 ; n27373_not
g86100 not n33268 ; n33268_not
g86101 not n27382 ; n27382_not
g86102 not n23647 ; n23647_not
g86103 not n27391 ; n27391_not
g86104 not n50368 ; n50368_not
g86105 not n55318 ; n55318_not
g86106 not n15745 ; n15745_not
g86107 not n15736 ; n15736_not
g86108 not n27409 ; n27409_not
g86109 not n27157 ; n27157_not
g86110 not n33394 ; n33394_not
g86111 not n55336 ; n55336_not
g86112 not n33385 ; n33385_not
g86113 not n27337 ; n27337_not
g86114 not n24376 ; n24376_not
g86115 not n27346 ; n27346_not
g86116 not n33367 ; n33367_not
g86117 not n55183 ; n55183_not
g86118 not n15772 ; n15772_not
g86119 not n33349 ; n33349_not
g86120 not n24367 ; n24367_not
g86121 not n55327 ; n55327_not
g86122 not n52843 ; n52843_not
g86123 not n27355 ; n27355_not
g86124 not n24358 ; n24358_not
g86125 not n27364 ; n27364_not
g86126 not n33295 ; n33295_not
g86127 not n52636 ; n52636_not
g86128 not n33169 ; n33169_not
g86129 not n50377 ; n50377_not
g86130 not n24277 ; n24277_not
g86131 not n27463 ; n27463_not
g86132 not n15691 ; n15691_not
g86133 not n52870 ; n52870_not
g86134 not n55309 ; n55309_not
g86135 not n50296 ; n50296_not
g86136 not n50386 ; n50386_not
g86137 not n24268 ; n24268_not
g86138 not n52627 ; n52627_not
g86139 not n15682 ; n15682_not
g86140 not n27085 ; n27085_not
g86141 not n27472 ; n27472_not
g86142 not n27418 ; n27418_not
g86143 not n27427 ; n27427_not
g86144 not n15727 ; n15727_not
g86145 not n52852 ; n52852_not
g86146 not n33196 ; n33196_not
g86147 not n32962 ; n32962_not
g86148 not n27436 ; n27436_not
g86149 not n33187 ; n33187_not
g86150 not n27445 ; n27445_not
g86151 not n24295 ; n24295_not
g86152 not n52861 ; n52861_not
g86153 not n33178 ; n33178_not
g86154 not n27454 ; n27454_not
g86155 not n24286 ; n24286_not
g86156 not n16753 ; n16753_not
g86157 not n52960 ; n52960_not
g86158 not n32377 ; n32377_not
g86159 not n32359 ; n32359_not
g86160 not n16762 ; n16762_not
g86161 not n16771 ; n16771_not
g86162 not n32287 ; n32287_not
g86163 not n32278 ; n32278_not
g86164 not n27634 ; n27634_not
g86165 not n16780 ; n16780_not
g86166 not n32269 ; n32269_not
g86167 not n23827 ; n23827_not
g86168 not n52573 ; n52573_not
g86169 not n16807 ; n16807_not
g86170 not n27643 ; n27643_not
g86171 not n55192 ; n55192_not
g86172 not n16348 ; n16348_not
g86173 not n16816 ; n16816_not
g86174 not n31990 ; n31990_not
g86175 not n32494 ; n32494_not
g86176 not n16681 ; n16681_not
g86177 not n32485 ; n32485_not
g86178 not n52591 ; n52591_not
g86179 not n32476 ; n32476_not
g86180 not n50494 ; n50494_not
g86181 not n16690 ; n16690_not
g86182 not n32467 ; n32467_not
g86183 not n32458 ; n32458_not
g86184 not n16708 ; n16708_not
g86185 not n55219 ; n55219_not
g86186 not n16717 ; n16717_not
g86187 not n32449 ; n32449_not
g86188 not n27625 ; n27625_not
g86189 not n52951 ; n52951_not
g86190 not n32368 ; n32368_not
g86191 not n16726 ; n16726_not
g86192 not n16393 ; n16393_not
g86193 not n16735 ; n16735_not
g86194 not n52582 ; n52582_not
g86195 not n32395 ; n32395_not
g86196 not n16744 ; n16744_not
g86197 not n55174 ; n55174_not
g86198 not n23962 ; n23962_not
g86199 not n55165 ; n55165_not
g86200 not n16906 ; n16906_not
g86201 not n16915 ; n16915_not
g86202 not n23953 ; n23953_not
g86203 not n50548 ; n50548_not
g86204 not n16924 ; n16924_not
g86205 not n50197 ; n50197_not
g86206 not n16933 ; n16933_not
g86207 not n23944 ; n23944_not
g86208 not n16825 ; n16825_not
g86209 not n32197 ; n32197_not
g86210 not n16834 ; n16834_not
g86211 not n27652 ; n27652_not
g86212 not n32188 ; n32188_not
g86213 not n32179 ; n32179_not
g86214 not n16843 ; n16843_not
g86215 not n32098 ; n32098_not
g86216 not n23980 ; n23980_not
g86217 not n16852 ; n16852_not
g86218 not n16861 ; n16861_not
g86219 not n27661 ; n27661_not
g86220 not n23971 ; n23971_not
g86221 not n50539 ; n50539_not
g86222 not n16870 ; n16870_not
g86223 not n27670 ; n27670_not
g86224 not n55264 ; n55264_not
g86225 not n27562 ; n27562_not
g86226 not n16537 ; n16537_not
g86227 not n50449 ; n50449_not
g86228 not n16546 ; n16546_not
g86229 not n27571 ; n27571_not
g86230 not n16555 ; n16555_not
g86231 not n32665 ; n32665_not
g86232 not n50458 ; n50458_not
g86233 not n16564 ; n16564_not
g86234 not n51871 ; n51871_not
g86235 not n27580 ; n27580_not
g86236 not n32674 ; n32674_not
g86237 not n55255 ; n55255_not
g86238 not n15943 ; n15943_not
g86239 not n15934 ; n15934_not
g86240 not n16465 ; n16465_not
g86241 not n15925 ; n15925_not
g86242 not n16474 ; n16474_not
g86243 not n15916 ; n15916_not
g86244 not n24169 ; n24169_not
g86245 not n15907 ; n15907_not
g86246 not n27553 ; n27553_not
g86247 not n23737 ; n23737_not
g86248 not n55273 ; n55273_not
g86249 not n16492 ; n16492_not
g86250 not n15880 ; n15880_not
g86251 not n15871 ; n15871_not
g86252 not n32629 ; n32629_not
g86253 not n32638 ; n32638_not
g86254 not n55237 ; n55237_not
g86255 not n16627 ; n16627_not
g86256 not n24088 ; n24088_not
g86257 not n23782 ; n23782_not
g86258 not n27607 ; n27607_not
g86259 not n16636 ; n16636_not
g86260 not n24079 ; n24079_not
g86261 not n50485 ; n50485_not
g86262 not n16645 ; n16645_not
g86263 not n32566 ; n32566_not
g86264 not n16438 ; n16438_not
g86265 not n16654 ; n16654_not
g86266 not n32557 ; n32557_not
g86267 not n16663 ; n16663_not
g86268 not n32548 ; n32548_not
g86269 not n27616 ; n27616_not
g86270 not n32539 ; n32539_not
g86271 not n52942 ; n52942_not
g86272 not n16672 ; n16672_not
g86273 not n53563 ; n53563_not
g86274 not n32683 ; n32683_not
g86275 not n16483 ; n16483_not
g86276 not n52915 ; n52915_not
g86277 not n16573 ; n16573_not
g86278 not n16582 ; n16582_not
g86279 not n50467 ; n50467_not
g86280 not n52924 ; n52924_not
g86281 not n55228 ; n55228_not
g86282 not n16591 ; n16591_not
g86283 not n32692 ; n32692_not
g86284 not n24097 ; n24097_not
g86285 not n16609 ; n16609_not
g86286 not n52933 ; n52933_not
g86287 not n16618 ; n16618_not
g86288 not n32647 ; n32647_not
g86289 not n50476 ; n50476_not
g86290 not n28831 ; n28831_not
g86291 not n19444 ; n19444_not
g86292 not n53284 ; n53284_not
g86293 not n19453 ; n19453_not
g86294 not n19462 ; n19462_not
g86295 not n28309 ; n28309_not
g86296 not n53554 ; n53554_not
g86297 not n28822 ; n28822_not
g86298 not n28813 ; n28813_not
g86299 not n21928 ; n21928_not
g86300 not n19471 ; n19471_not
g86301 not n21919 ; n21919_not
g86302 not n19480 ; n19480_not
g86303 not n28804 ; n28804_not
g86304 not n50944 ; n50944_not
g86305 not n19192 ; n19192_not
g86306 not n21892 ; n21892_not
g86307 not n19183 ; n19183_not
g86308 not n19507 ; n19507_not
g86309 not n19516 ; n19516_not
g86310 not n19525 ; n19525_not
g86311 not n19336 ; n19336_not
g86312 not n21946 ; n21946_not
g86313 not n19273 ; n19273_not
g86314 not n19345 ; n19345_not
g86315 not n28084 ; n28084_not
g86316 not n19354 ; n19354_not
g86317 not n19363 ; n19363_not
g86318 not n53266 ; n53266_not
g86319 not n19372 ; n19372_not
g86320 not n19381 ; n19381_not
g86321 not n19390 ; n19390_not
g86322 not n19246 ; n19246_not
g86323 not n50962 ; n50962_not
g86324 not n19237 ; n19237_not
g86325 not n21937 ; n21937_not
g86326 not n19408 ; n19408_not
g86327 not n51619 ; n51619_not
g86328 not n53275 ; n53275_not
g86329 not n50953 ; n50953_not
g86330 not n19417 ; n19417_not
g86331 not n19228 ; n19228_not
g86332 not n19426 ; n19426_not
g86333 not n28840 ; n28840_not
g86334 not n19435 ; n19435_not
g86335 not n19624 ; n19624_not
g86336 not n19633 ; n19633_not
g86337 not n51637 ; n51637_not
g86338 not n19642 ; n19642_not
g86339 not n19651 ; n19651_not
g86340 not n28714 ; n28714_not
g86341 not n19660 ; n19660_not
g86342 not n28705 ; n28705_not
g86343 not n19093 ; n19093_not
g86344 not n53356 ; n53356_not
g86345 not n28192 ; n28192_not
g86346 not n53365 ; n53365_not
g86347 not n53374 ; n53374_not
g86348 not n21856 ; n21856_not
g86349 not n19705 ; n19705_not
g86350 not n19714 ; n19714_not
g86351 not n19066 ; n19066_not
g86352 not n19723 ; n19723_not
g86353 not n21847 ; n21847_not
g86354 not n19534 ; n19534_not
g86355 not n28750 ; n28750_not
g86356 not n28741 ; n28741_not
g86357 not n19543 ; n19543_not
g86358 not n19552 ; n19552_not
g86359 not n19156 ; n19156_not
g86360 not n19561 ; n19561_not
g86361 not n19147 ; n19147_not
g86362 not n21883 ; n21883_not
g86363 not n19570 ; n19570_not
g86364 not n21874 ; n21874_not
g86365 not n53329 ; n53329_not
g86366 not n28732 ; n28732_not
g86367 not n28723 ; n28723_not
g86368 not n19138 ; n19138_not
g86369 not n28327 ; n28327_not
g86370 not n19606 ; n19606_not
g86371 not n19615 ; n19615_not
g86372 not n21865 ; n21865_not
g86373 not n51673 ; n51673_not
g86374 not n29254 ; n29254_not
g86375 not n19165 ; n19165_not
g86376 not n51565 ; n51565_not
g86377 not n51574 ; n51574_not
g86378 not n29155 ; n29155_not
g86379 not n22279 ; n22279_not
g86380 not n29227 ; n29227_not
g86381 not n29164 ; n29164_not
g86382 not n29218 ; n29218_not
g86383 not n29209 ; n29209_not
g86384 not n29191 ; n29191_not
g86385 not n22189 ; n22189_not
g86386 not n29173 ; n29173_not
g86387 not n22099 ; n22099_not
g86388 not n51583 ; n51583_not
g86389 not n51682 ; n51682_not
g86390 not n29281 ; n29281_not
g86391 not n51556 ; n51556_not
g86392 not n29263 ; n29263_not
g86393 not n54148 ; n54148_not
g86394 not n28255 ; n28255_not
g86395 not n22378 ; n22378_not
g86396 not n52438 ; n52438_not
g86397 not n22369 ; n22369_not
g86398 not n22297 ; n22297_not
g86399 not n29272 ; n29272_not
g86400 not n51592 ; n51592_not
g86401 not n29074 ; n29074_not
g86402 not n29065 ; n29065_not
g86403 not n29056 ; n29056_not
g86404 not n53239 ; n53239_not
g86405 not n28291 ; n28291_not
g86406 not n29047 ; n29047_not
g86407 not n19282 ; n19282_not
g86408 not n29038 ; n29038_not
g86409 not n29029 ; n29029_not
g86410 not n21964 ; n21964_not
g86411 not n21289 ; n21289_not
g86412 not n51655 ; n51655_not
g86413 not n18607 ; n18607_not
g86414 not n21955 ; n21955_not
g86415 not n19309 ; n19309_not
g86416 not n21298 ; n21298_not
g86417 not n19291 ; n19291_not
g86418 not n19318 ; n19318_not
g86419 not n28903 ; n28903_not
g86420 not n19327 ; n19327_not
g86421 not n28912 ; n28912_not
g86422 not n52429 ; n52429_not
g86423 not n29146 ; n29146_not
g86424 not n28282 ; n28282_not
g86425 not n29137 ; n29137_not
g86426 not n54076 ; n54076_not
g86427 not n21991 ; n21991_not
g86428 not n29092 ; n29092_not
g86429 not n19255 ; n19255_not
g86430 not n21982 ; n21982_not
g86431 not n29083 ; n29083_not
g86432 not n53248 ; n53248_not
g86433 not n21973 ; n21973_not
g86434 not n20497 ; n20497_not
g86435 not n21586 ; n21586_not
g86436 not n20569 ; n20569_not
g86437 not n28264 ; n28264_not
g86438 not n20587 ; n20587_not
g86439 not n28543 ; n28543_not
g86440 not n28426 ; n28426_not
g86441 not n53455 ; n53455_not
g86442 not n20659 ; n20659_not
g86443 not n21577 ; n21577_not
g86444 not n28534 ; n28534_not
g86445 not n20677 ; n20677_not
g86446 not n28525 ; n28525_not
g86447 not n20695 ; n20695_not
g86448 not n20749 ; n20749_not
g86449 not n21568 ; n21568_not
g86450 not n21559 ; n21559_not
g86451 not n20767 ; n20767_not
g86452 not n20758 ; n20758_not
g86453 not n20785 ; n20785_not
g86454 not n20794 ; n20794_not
g86455 not n28435 ; n28435_not
g86456 not n28516 ; n28516_not
g86457 not n53446 ; n53446_not
g86458 not n19840 ; n19840_not
g86459 not n52771 ; n52771_not
g86460 not n28552 ; n28552_not
g86461 not n50863 ; n50863_not
g86462 not n52780 ; n52780_not
g86463 not n21649 ; n21649_not
g86464 not n20389 ; n20389_not
g86465 not n53491 ; n53491_not
g86466 not n28417 ; n28417_not
g86467 not n20398 ; n20398_not
g86468 not n21469 ; n21469_not
g86469 not n52807 ; n52807_not
g86470 not n19813 ; n19813_not
g86471 not n21478 ; n21478_not
g86472 not n19804 ; n19804_not
g86473 not n52816 ; n52816_not
g86474 not n52825 ; n52825_not
g86475 not n52834 ; n52834_not
g86476 not n53473 ; n53473_not
g86477 not n20479 ; n20479_not
g86478 not n21595 ; n21595_not
g86479 not n20668 ; n20668_not
g86480 not n20956 ; n20956_not
g86481 not n28480 ; n28480_not
g86482 not n21397 ; n21397_not
g86483 not n20965 ; n20965_not
g86484 not n20974 ; n20974_not
g86485 not n21379 ; n21379_not
g86486 not n20983 ; n20983_not
g86487 not n20992 ; n20992_not
g86488 not n28471 ; n28471_not
g86489 not n28453 ; n28453_not
g86490 not n53383 ; n53383_not
g86491 not n21199 ; n21199_not
g86492 not n20578 ; n20578_not
g86493 not n28462 ; n28462_not
g86494 not n53338 ; n53338_not
g86495 not n28507 ; n28507_not
g86496 not n20839 ; n20839_not
g86497 not n20848 ; n20848_not
g86498 not n20857 ; n20857_not
g86499 not n50854 ; n50854_not
g86500 not n20866 ; n20866_not
g86501 not n20875 ; n20875_not
g86502 not n21487 ; n21487_not
g86503 not n53428 ; n53428_not
g86504 not n20884 ; n20884_not
g86505 not n20893 ; n20893_not
g86506 not n20929 ; n20929_not
g86507 not n20938 ; n20938_not
g86508 not n28444 ; n28444_not
g86509 not n20947 ; n20947_not
g86510 not n21388 ; n21388_not
g86511 not n28660 ; n28660_not
g86512 not n28363 ; n28363_not
g86513 not n28651 ; n28651_not
g86514 not n53176 ; n53176_not
g86515 not n19912 ; n19912_not
g86516 not n28642 ; n28642_not
g86517 not n51628 ; n51628_not
g86518 not n28372 ; n28372_not
g86519 not n21784 ; n21784_not
g86520 not n28633 ; n28633_not
g86521 not n19930 ; n19930_not
g86522 not n50827 ; n50827_not
g86523 not n21775 ; n21775_not
g86524 not n53464 ; n53464_not
g86525 not n50917 ; n50917_not
g86526 not n19057 ; n19057_not
g86527 not n19732 ; n19732_not
g86528 not n19741 ; n19741_not
g86529 not n50908 ; n50908_not
g86530 not n19048 ; n19048_not
g86531 not n21838 ; n21838_not
g86532 not n53194 ; n53194_not
g86533 not n28345 ; n28345_not
g86534 not n21829 ; n21829_not
g86535 not n53185 ; n53185_not
g86536 not n19822 ; n19822_not
g86537 not n53419 ; n53419_not
g86538 not n21793 ; n21793_not
g86539 not n21694 ; n21694_not
g86540 not n21685 ; n21685_not
g86541 not n21676 ; n21676_not
g86542 not n19903 ; n19903_not
g86543 not n27814 ; n27814_not
g86544 not n28570 ; n28570_not
g86545 not n53536 ; n53536_not
g86546 not n27904 ; n27904_not
g86547 not n50872 ; n50872_not
g86548 not n53545 ; n53545_not
g86549 not n21667 ; n21667_not
g86550 not n28561 ; n28561_not
g86551 not n20299 ; n20299_not
g86552 not n52735 ; n52735_not
g86553 not n28408 ; n28408_not
g86554 not n52744 ; n52744_not
g86555 not n21658 ; n21658_not
g86556 not n52753 ; n52753_not
g86557 not n53518 ; n53518_not
g86558 not n52762 ; n52762_not
g86559 not n28624 ; n28624_not
g86560 not n28615 ; n28615_not
g86561 not n28381 ; n28381_not
g86562 not n21766 ; n21766_not
g86563 not n53167 ; n53167_not
g86564 not n28336 ; n28336_not
g86565 not n21757 ; n21757_not
g86566 not n53293 ; n53293_not
g86567 not n28606 ; n28606_not
g86568 not n21748 ; n21748_not
g86569 not n21739 ; n21739_not
g86570 not n53509 ; n53509_not
g86571 not n28390 ; n28390_not
g86572 not n53158 ; n53158_not
g86573 not n53149 ; n53149_not
g86574 not n18490 ; n18490_not
g86575 not n29713 ; n29713_not
g86576 not n18517 ; n18517_not
g86577 not n53680 ; n53680_not
g86578 not n29704 ; n29704_not
g86579 not n17950 ; n17950_not
g86580 not n18535 ; n18535_not
g86581 not n17941 ; n17941_not
g86582 not n18544 ; n18544_not
g86583 not n17932 ; n17932_not
g86584 not n51466 ; n51466_not
g86585 not n50926 ; n50926_not
g86586 not n54319 ; n54319_not
g86587 not n17923 ; n17923_not
g86588 not n17914 ; n17914_not
g86589 not n17905 ; n17905_not
g86590 not n18562 ; n18562_not
g86591 not n29830 ; n29830_not
g86592 not n18427 ; n18427_not
g86593 not n18148 ; n18148_not
g86594 not n29911 ; n29911_not
g86595 not n18139 ; n18139_not
g86596 not n18445 ; n18445_not
g86597 not n53707 ; n53707_not
g86598 not n50881 ; n50881_not
g86599 not n18454 ; n18454_not
g86600 not n18094 ; n18094_not
g86601 not n28075 ; n28075_not
g86602 not n22846 ; n22846_not
g86603 not n18085 ; n18085_not
g86604 not n29740 ; n29740_not
g86605 not n18076 ; n18076_not
g86606 not n18067 ; n18067_not
g86607 not n18472 ; n18472_not
g86608 not n18058 ; n18058_not
g86609 not n29722 ; n29722_not
g86610 not n18049 ; n18049_not
g86611 not n29731 ; n29731_not
g86612 not n22747 ; n22747_not
g86613 not n18553 ; n18553_not
g86614 not n28039 ; n28039_not
g86615 not n53626 ; n53626_not
g86616 not n28138 ; n28138_not
g86617 not n22738 ; n22738_not
g86618 not n54346 ; n54346_not
g86619 not n53617 ; n53617_not
g86620 not n28147 ; n28147_not
g86621 not n22729 ; n22729_not
g86622 not n29650 ; n29650_not
g86623 not n53608 ; n53608_not
g86624 not n22693 ; n22693_not
g86625 not n29605 ; n29605_not
g86626 not n28156 ; n28156_not
g86627 not n53671 ; n53671_not
g86628 not n28093 ; n28093_not
g86629 not n53662 ; n53662_not
g86630 not n22783 ; n22783_not
g86631 not n51727 ; n51727_not
g86632 not n18580 ; n18580_not
g86633 not n53653 ; n53653_not
g86634 not n50971 ; n50971_not
g86635 not n22774 ; n22774_not
g86636 not n53644 ; n53644_not
g86637 not n51475 ; n51475_not
g86638 not n22765 ; n22765_not
g86639 not n28066 ; n28066_not
g86640 not n53635 ; n53635_not
g86641 not n22756 ; n22756_not
g86642 not n51457 ; n51457_not
g86643 not n22981 ; n22981_not
g86644 not n50746 ; n50746_not
g86645 not n50755 ; n50755_not
g86646 not n50764 ; n50764_not
g86647 not n53743 ; n53743_not
g86648 not n17653 ; n17653_not
g86649 not n29902 ; n29902_not
g86650 not n50773 ; n50773_not
g86651 not n22936 ; n22936_not
g86652 not n53734 ; n53734_not
g86653 not n50782 ; n50782_not
g86654 not n50791 ; n50791_not
g86655 not n50737 ; n50737_not
g86656 not n53770 ; n53770_not
g86657 not n52483 ; n52483_not
g86658 not n23089 ; n23089_not
g86659 not n54265 ; n54265_not
g86660 not n30469 ; n30469_not
g86661 not n30289 ; n30289_not
g86662 not n53761 ; n53761_not
g86663 not n28048 ; n28048_not
g86664 not n30298 ; n30298_not
g86665 not n54274 ; n54274_not
g86666 not n53752 ; n53752_not
g86667 not n30199 ; n30199_not
g86668 not n18238 ; n18238_not
g86669 not n18229 ; n18229_not
g86670 not n18382 ; n18382_not
g86671 not n53716 ; n53716_not
g86672 not n18193 ; n18193_not
g86673 not n18184 ; n18184_not
g86674 not n29920 ; n29920_not
g86675 not n18409 ; n18409_not
g86676 not n18175 ; n18175_not
g86677 not n18166 ; n18166_not
g86678 not n18157 ; n18157_not
g86679 not n53725 ; n53725_not
g86680 not n50809 ; n50809_not
g86681 not n18319 ; n18319_not
g86682 not n18328 ; n18328_not
g86683 not n22891 ; n22891_not
g86684 not n29821 ; n29821_not
g86685 not n18337 ; n18337_not
g86686 not n18292 ; n18292_not
g86687 not n18283 ; n18283_not
g86688 not n18274 ; n18274_not
g86689 not n18355 ; n18355_not
g86690 not n18265 ; n18265_not
g86691 not n50836 ; n50836_not
g86692 not n18364 ; n18364_not
g86693 not n18256 ; n18256_not
g86694 not n18247 ; n18247_not
g86695 not n22558 ; n22558_not
g86696 not n29353 ; n29353_not
g86697 not n28228 ; n28228_not
g86698 not n22549 ; n22549_not
g86699 not n22495 ; n22495_not
g86700 not n29326 ; n29326_not
g86701 not n54238 ; n54238_not
g86702 not n29317 ; n29317_not
g86703 not n51547 ; n51547_not
g86704 not n22486 ; n22486_not
g86705 not n28237 ; n28237_not
g86706 not n22576 ; n22576_not
g86707 not n51538 ; n51538_not
g86708 not n28219 ; n28219_not
g86709 not n29461 ; n29461_not
g86710 not n18418 ; n18418_not
g86711 not n29470 ; n29470_not
g86712 not n22567 ; n22567_not
g86713 not n54283 ; n54283_not
g86714 not n51079 ; n51079_not
g86715 not n29344 ; n29344_not
g86716 not n29290 ; n29290_not
g86717 not n22459 ; n22459_not
g86718 not n29308 ; n29308_not
g86719 not n29362 ; n29362_not
g86720 not n19039 ; n19039_not
g86721 not n22396 ; n22396_not
g86722 not n19075 ; n19075_not
g86723 not n29335 ; n29335_not
g86724 not n22387 ; n22387_not
g86725 not n29407 ; n29407_not
g86726 not n18373 ; n18373_not
g86727 not n22477 ; n22477_not
g86728 not n29380 ; n29380_not
g86729 not n54193 ; n54193_not
g86730 not n22468 ; n22468_not
g86731 not n52456 ; n52456_not
g86732 not n29524 ; n29524_not
g86733 not n51493 ; n51493_not
g86734 not n28183 ; n28183_not
g86735 not n54382 ; n54382_not
g86736 not n29533 ; n29533_not
g86737 not n29632 ; n29632_not
g86738 not n29542 ; n29542_not
g86739 not n29551 ; n29551_not
g86740 not n22648 ; n22648_not
g86741 not n29560 ; n29560_not
g86742 not n51088 ; n51088_not
g86743 not n29614 ; n29614_not
g86744 not n54373 ; n54373_not
g86745 not n53572 ; n53572_not
g86746 not n22639 ; n22639_not
g86747 not n54355 ; n54355_not
g86748 not n22684 ; n22684_not
g86749 not n51484 ; n51484_not
g86750 not n54364 ; n54364_not
g86751 not n53590 ; n53590_not
g86752 not n29623 ; n29623_not
g86753 not n51718 ; n51718_not
g86754 not n18508 ; n18508_not
g86755 not n22675 ; n22675_not
g86756 not n28165 ; n28165_not
g86757 not n53581 ; n53581_not
g86758 not n22666 ; n22666_not
g86759 not n22657 ; n22657_not
g86760 not n22594 ; n22594_not
g86761 not n29515 ; n29515_not
g86762 not n52447 ; n52447_not
g86763 not n54328 ; n54328_not
g86764 not n51097 ; n51097_not
g86765 not n22585 ; n22585_not
g86766 not n29506 ; n29506_not
g86767 not n51529 ; n51529_not
g86768 not n18463 ; n18463_not
g86769 not n13909 ; n13909_not
g86770 not n13927 ; n13927_not
g86771 not n49126 ; n49126_not
g86772 not n25618 ; n25618_not
g86773 not n48631 ; n48631_not
g86774 not n13936 ; n13936_not
g86775 not n55714 ; n55714_not
g86776 not n26815 ; n26815_not
g86777 not n25537 ; n25537_not
g86778 not n12784 ; n12784_not
g86779 not n35464 ; n35464_not
g86780 not n10687 ; n10687_not
g86781 not n35293 ; n35293_not
g86782 not n13954 ; n13954_not
g86783 not n55723 ; n55723_not
g86784 not n13945 ; n13945_not
g86785 not n49405 ; n49405_not
g86786 not n10678 ; n10678_not
g86787 not n10669 ; n10669_not
g86788 not n49117 ; n49117_not
g86789 not n55651 ; n55651_not
g86790 not n13819 ; n13819_not
g86791 not n10768 ; n10768_not
g86792 not n55660 ; n55660_not
g86793 not n13837 ; n13837_not
g86794 not n13846 ; n13846_not
g86795 not n35338 ; n35338_not
g86796 not n49360 ; n49360_not
g86797 not n10759 ; n10759_not
g86798 not n26806 ; n26806_not
g86799 not n25465 ; n25465_not
g86800 not n13864 ; n13864_not
g86801 not n25627 ; n25627_not
g86802 not n10696 ; n10696_not
g86803 not n13882 ; n13882_not
g86804 not n55705 ; n55705_not
g86805 not n13891 ; n13891_not
g86806 not n25960 ; n25960_not
g86807 not n35860 ; n35860_not
g86808 not n25474 ; n25474_not
g86809 not n55840 ; n55840_not
g86810 not n10588 ; n10588_not
g86811 not n25591 ; n25591_not
g86812 not n49108 ; n49108_not
g86813 not n35167 ; n35167_not
g86814 not n35482 ; n35482_not
g86815 not n26833 ; n26833_not
g86816 not n13855 ; n13855_not
g86817 not n10579 ; n10579_not
g86818 not n35158 ; n35158_not
g86819 not n49432 ; n49432_not
g86820 not n35149 ; n35149_not
g86821 not n26824 ; n26824_not
g86822 not n25609 ; n25609_not
g86823 not n35275 ; n35275_not
g86824 not n55732 ; n55732_not
g86825 not n35473 ; n35473_not
g86826 not n35257 ; n35257_not
g86827 not n35248 ; n35248_not
g86828 not n26626 ; n26626_not
g86829 not n55741 ; n55741_not
g86830 not n55822 ; n55822_not
g86831 not n55750 ; n55750_not
g86832 not n35185 ; n35185_not
g86833 not n55813 ; n55813_not
g86834 not n10597 ; n10597_not
g86835 not n25276 ; n25276_not
g86836 not n35176 ; n35176_not
g86837 not n49414 ; n49414_not
g86838 not n25294 ; n25294_not
g86839 not n55543 ; n55543_not
g86840 not n25663 ; n25663_not
g86841 not n55930 ; n55930_not
g86842 not n13198 ; n13198_not
g86843 not n55552 ; n55552_not
g86844 not n49324 ; n49324_not
g86845 not n13639 ; n13639_not
g86846 not n55561 ; n55561_not
g86847 not n13648 ; n13648_not
g86848 not n49144 ; n49144_not
g86849 not n13657 ; n13657_not
g86850 not n35842 ; n35842_not
g86851 not n13666 ; n13666_not
g86852 not n55516 ; n55516_not
g86853 not n25942 ; n25942_not
g86854 not n35833 ; n35833_not
g86855 not n13558 ; n13558_not
g86856 not n25681 ; n25681_not
g86857 not n52555 ; n52555_not
g86858 not n13567 ; n13567_not
g86859 not n10885 ; n10885_not
g86860 not n55525 ; n55525_not
g86861 not n13576 ; n13576_not
g86862 not n10867 ; n10867_not
g86863 not n25672 ; n25672_not
g86864 not n13585 ; n13585_not
g86865 not n55534 ; n55534_not
g86866 not n49315 ; n49315_not
g86867 not n35437 ; n35437_not
g86868 not n13594 ; n13594_not
g86869 not n10849 ; n10849_not
g86870 not n55606 ; n55606_not
g86871 not n49135 ; n49135_not
g86872 not n13756 ; n13756_not
g86873 not n35851 ; n35851_not
g86874 not n25645 ; n25645_not
g86875 not n55615 ; n55615_not
g86876 not n26635 ; n26635_not
g86877 not n55624 ; n55624_not
g86878 not n25636 ; n25636_not
g86879 not n13774 ; n13774_not
g86880 not n55633 ; n55633_not
g86881 not n35455 ; n35455_not
g86882 not n51736 ; n51736_not
g86883 not n35347 ; n35347_not
g86884 not n35707 ; n35707_not
g86885 not n13792 ; n13792_not
g86886 not n55642 ; n55642_not
g86887 not n25951 ; n25951_not
g86888 not n55570 ; n55570_not
g86889 not n13675 ; n13675_not
g86890 not n10795 ; n10795_not
g86891 not n25654 ; n25654_not
g86892 not n13684 ; n13684_not
g86893 not n35446 ; n35446_not
g86894 not n49342 ; n49342_not
g86895 not n55912 ; n55912_not
g86896 not n35716 ; n35716_not
g86897 not n13693 ; n13693_not
g86898 not n55903 ; n55903_not
g86899 not n25456 ; n25456_not
g86900 not n13729 ; n13729_not
g86901 not n10786 ; n10786_not
g86902 not n13738 ; n13738_not
g86903 not n25285 ; n25285_not
g86904 not n10777 ; n10777_not
g86905 not n13747 ; n13747_not
g86906 not n14566 ; n14566_not
g86907 not n49603 ; n49603_not
g86908 not n49540 ; n49540_not
g86909 not n14575 ; n14575_not
g86910 not n49612 ; n49612_not
g86911 not n13981 ; n13981_not
g86912 not n14557 ; n14557_not
g86913 not n14584 ; n14584_not
g86914 not n25933 ; n25933_not
g86915 not n49621 ; n49621_not
g86916 not n35923 ; n35923_not
g86917 not n13972 ; n13972_not
g86918 not n26068 ; n26068_not
g86919 not n14539 ; n14539_not
g86920 not n25519 ; n25519_not
g86921 not n26590 ; n26590_not
g86922 not n26077 ; n26077_not
g86923 not n26086 ; n26086_not
g86924 not n13990 ; n13990_not
g86925 not n35914 ; n35914_not
g86926 not n55921 ; n55921_not
g86927 not n49072 ; n49072_not
g86928 not n25528 ; n25528_not
g86929 not n35518 ; n35518_not
g86930 not n35932 ; n35932_not
g86931 not n26176 ; n26176_not
g86932 not n25870 ; n25870_not
g86933 not n49513 ; n49513_not
g86934 not n26059 ; n26059_not
g86935 not n49054 ; n49054_not
g86936 not n26572 ; n26572_not
g86937 not n35536 ; n35536_not
g86938 not n35662 ; n35662_not
g86939 not n49504 ; n49504_not
g86940 not n25861 ; n25861_not
g86941 not n14089 ; n14089_not
g86942 not n14098 ; n14098_not
g86943 not n25438 ; n25438_not
g86944 not n34960 ; n34960_not
g86945 not n14593 ; n14593_not
g86946 not n49630 ; n49630_not
g86947 not n34870 ; n34870_not
g86948 not n26581 ; n26581_not
g86949 not n25483 ; n25483_not
g86950 not n25924 ; n25924_not
g86951 not n49063 ; n49063_not
g86952 not n35527 ; n35527_not
g86953 not n26149 ; n26149_not
g86954 not n25915 ; n25915_not
g86955 not n35671 ; n35671_not
g86956 not n25906 ; n25906_not
g86957 not n26167 ; n26167_not
g86958 not n25564 ; n25564_not
g86959 not n26851 ; n26851_not
g86960 not n14359 ; n14359_not
g86961 not n35086 ; n35086_not
g86962 not n51691 ; n51691_not
g86963 not n14296 ; n14296_not
g86964 not n14377 ; n14377_not
g86965 not n26608 ; n26608_not
g86966 not n49090 ; n49090_not
g86967 not n14287 ; n14287_not
g86968 not n14386 ; n14386_not
g86969 not n14278 ; n14278_not
g86970 not n35077 ; n35077_not
g86971 not n26617 ; n26617_not
g86972 not n10489 ; n10489_not
g86973 not n34780 ; n34780_not
g86974 not n25582 ; n25582_not
g86975 not n10399 ; n10399_not
g86976 not n26842 ; n26842_not
g86977 not n49450 ; n49450_not
g86978 not n25573 ; n25573_not
g86979 not n35491 ; n35491_not
g86980 not n35095 ; n35095_not
g86981 not n13765 ; n13765_not
g86982 not n14449 ; n14449_not
g86983 not n26095 ; n26095_not
g86984 not n14467 ; n14467_not
g86985 not n25546 ; n25546_not
g86986 not n49522 ; n49522_not
g86987 not n14476 ; n14476_not
g86988 not n34834 ; n34834_not
g86989 not n35509 ; n35509_not
g86990 not n26860 ; n26860_not
g86991 not n34843 ; n34843_not
g86992 not n14494 ; n14494_not
g86993 not n25555 ; n25555_not
g86994 not n25249 ; n25249_not
g86995 not n14269 ; n14269_not
g86996 not n35068 ; n35068_not
g86997 not n14197 ; n14197_not
g86998 not n34825 ; n34825_not
g86999 not n35059 ; n35059_not
g87000 not n35905 ; n35905_not
g87001 not n14188 ; n14188_not
g87002 not n49081 ; n49081_not
g87003 not n14179 ; n14179_not
g87004 not n12478 ; n12478_not
g87005 not n12487 ; n12487_not
g87006 not n49234 ; n49234_not
g87007 not n12496 ; n12496_not
g87008 not n35680 ; n35680_not
g87009 not n56083 ; n56083_not
g87010 not n11992 ; n11992_not
g87011 not n11587 ; n11587_not
g87012 not n11983 ; n11983_not
g87013 not n12559 ; n12559_not
g87014 not n12568 ; n12568_not
g87015 not n26725 ; n26725_not
g87016 not n25375 ; n25375_not
g87017 not n11659 ; n11659_not
g87018 not n56092 ; n56092_not
g87019 not n12289 ; n12289_not
g87020 not n11596 ; n11596_not
g87021 not n12298 ; n12298_not
g87022 not n56119 ; n56119_not
g87023 not n12379 ; n12379_not
g87024 not n12388 ; n12388_not
g87025 not n25807 ; n25807_not
g87026 not n12397 ; n12397_not
g87027 not n12469 ; n12469_not
g87028 not n26716 ; n26716_not
g87029 not n12757 ; n12757_not
g87030 not n35545 ; n35545_not
g87031 not n12748 ; n12748_not
g87032 not n35383 ; n35383_not
g87033 not n56065 ; n56065_not
g87034 not n12739 ; n12739_not
g87035 not n12793 ; n12793_not
g87036 not n25384 ; n25384_not
g87037 not n35554 ; n35554_not
g87038 not n49243 ; n49243_not
g87039 not n26734 ; n26734_not
g87040 not n26662 ; n26662_not
g87041 not n12829 ; n12829_not
g87042 not n12838 ; n12838_not
g87043 not n25780 ; n25780_not
g87044 not n12847 ; n12847_not
g87045 not n12586 ; n12586_not
g87046 not n11578 ; n11578_not
g87047 not n12649 ; n12649_not
g87048 not n12658 ; n12658_not
g87049 not n11497 ; n11497_not
g87050 not n11488 ; n11488_not
g87051 not n12676 ; n12676_not
g87052 not n12694 ; n12694_not
g87053 not n35653 ; n35653_not
g87054 not n35761 ; n35761_not
g87055 not n49216 ; n49216_not
g87056 not n11758 ; n11758_not
g87057 not n35374 ; n35374_not
g87058 not n11848 ; n11848_not
g87059 not n35770 ; n35770_not
g87060 not n11749 ; n11749_not
g87061 not n11857 ; n11857_not
g87062 not n25852 ; n25852_not
g87063 not n11866 ; n11866_not
g87064 not n11875 ; n11875_not
g87065 not n56047 ; n56047_not
g87066 not n11884 ; n11884_not
g87067 not n11893 ; n11893_not
g87068 not n25843 ; n25843_not
g87069 not n35743 ; n35743_not
g87070 not n11776 ; n11776_not
g87071 not n56056 ; n56056_not
g87072 not n35365 ; n35365_not
g87073 not n11785 ; n11785_not
g87074 not n25339 ; n25339_not
g87075 not n26680 ; n26680_not
g87076 not n11794 ; n11794_not
g87077 not n11767 ; n11767_not
g87078 not n35356 ; n35356_not
g87079 not n49207 ; n49207_not
g87080 not n11299 ; n11299_not
g87081 not n35752 ; n35752_not
g87082 not n11839 ; n11839_not
g87083 not n35725 ; n35725_not
g87084 not n35419 ; n35419_not
g87085 not n35428 ; n35428_not
g87086 not n11677 ; n11677_not
g87087 not n26707 ; n26707_not
g87088 not n12199 ; n12199_not
g87089 not n25816 ; n25816_not
g87090 not n11668 ; n11668_not
g87091 not n25366 ; n25366_not
g87092 not n49225 ; n49225_not
g87093 not n11389 ; n11389_not
g87094 not n11929 ; n11929_not
g87095 not n11398 ; n11398_not
g87096 not n11938 ; n11938_not
g87097 not n26185 ; n26185_not
g87098 not n11947 ; n11947_not
g87099 not n35392 ; n35392_not
g87100 not n25834 ; n25834_not
g87101 not n11956 ; n11956_not
g87102 not n11974 ; n11974_not
g87103 not n11695 ; n11695_not
g87104 not n26671 ; n26671_not
g87105 not n11686 ; n11686_not
g87106 not n25825 ; n25825_not
g87107 not n35815 ; n35815_not
g87108 not n25735 ; n25735_not
g87109 not n13369 ; n13369_not
g87110 not n13378 ; n13378_not
g87111 not n55417 ; n55417_not
g87112 not n13387 ; n13387_not
g87113 not n13396 ; n13396_not
g87114 not n55426 ; n55426_not
g87115 not n10984 ; n10984_not
g87116 not n25726 ; n25726_not
g87117 not n55435 ; n55435_not
g87118 not n12973 ; n12973_not
g87119 not n12964 ; n12964_not
g87120 not n12955 ; n12955_not
g87121 not n12946 ; n12946_not
g87122 not n12937 ; n12937_not
g87123 not n12928 ; n12928_not
g87124 not n12919 ; n12919_not
g87125 not n49270 ; n49270_not
g87126 not n12892 ; n12892_not
g87127 not n12883 ; n12883_not
g87128 not n13288 ; n13288_not
g87129 not n12874 ; n12874_not
g87130 not n13297 ; n13297_not
g87131 not n12865 ; n12865_not
g87132 not n25744 ; n25744_not
g87133 not n12856 ; n12856_not
g87134 not n26770 ; n26770_not
g87135 not n55471 ; n55471_not
g87136 not n13495 ; n13495_not
g87137 not n25429 ; n25429_not
g87138 not n55480 ; n55480_not
g87139 not n35824 ; n35824_not
g87140 not n26644 ; n26644_not
g87141 not n25690 ; n25690_not
g87142 not n55507 ; n55507_not
g87143 not n10939 ; n10939_not
g87144 not n35266 ; n35266_not
g87145 not n10894 ; n10894_not
g87146 not n13549 ; n13549_not
g87147 not n26761 ; n26761_not
g87148 not n10975 ; n10975_not
g87149 not n55444 ; n55444_not
g87150 not n25717 ; n25717_not
g87151 not n55453 ; n55453_not
g87152 not n52465 ; n52465_not
g87153 not n13459 ; n13459_not
g87154 not n49153 ; n49153_not
g87155 not n13468 ; n13468_not
g87156 not n25708 ; n25708_not
g87157 not n55462 ; n55462_not
g87158 not n13477 ; n13477_not
g87159 not n10957 ; n10957_not
g87160 not n13486 ; n13486_not
g87161 not n35590 ; n35590_not
g87162 not n25771 ; n25771_not
g87163 not n55345 ; n55345_not
g87164 not n26743 ; n26743_not
g87165 not n56038 ; n56038_not
g87166 not n10948 ; n10948_not
g87167 not n55354 ; n55354_not
g87168 not n12667 ; n12667_not
g87169 not n49171 ; n49171_not
g87170 not n35563 ; n35563_not
g87171 not n35572 ; n35572_not
g87172 not n49180 ; n49180_not
g87173 not n35581 ; n35581_not
g87174 not n35635 ; n35635_not
g87175 not n12991 ; n12991_not
g87176 not n25753 ; n25753_not
g87177 not n55381 ; n55381_not
g87178 not n55390 ; n55390_not
g87179 not n35806 ; n35806_not
g87180 not n49162 ; n49162_not
g87181 not n26752 ; n26752_not
g87182 not n12577 ; n12577_not
g87183 not n49261 ; n49261_not
g87184 not n10993 ; n10993_not
g87185 not n13099 ; n13099_not
g87186 not n55408 ; n55408_not
g87187 not n12982 ; n12982_not
g87188 not n35617 ; n35617_not
g87189 not n26653 ; n26653_not
g87190 not n35608 ; n35608_not
g87191 not n25762 ; n25762_not
g87192 not n49252 ; n49252_not
g87193 not n55363 ; n55363_not
g87194 not n55372 ; n55372_not
g87195 not n33835 ; n33835_not
g87196 not n33844 ; n33844_not
g87197 not n34078 ; n34078_not
g87198 not n33853 ; n33853_not
g87199 not n33862 ; n33862_not
g87200 not n27166 ; n27166_not
g87201 not n33871 ; n33871_not
g87202 not n15475 ; n15475_not
g87203 not n33880 ; n33880_not
g87204 not n33907 ; n33907_not
g87205 not n15466 ; n15466_not
g87206 not n24664 ; n24664_not
g87207 not n33916 ; n33916_not
g87208 not n33925 ; n33925_not
g87209 not n33781 ; n33781_not
g87210 not n57226 ; n57226_not
g87211 not n33790 ; n33790_not
g87212 not n33808 ; n33808_not
g87213 not n33817 ; n33817_not
g87214 not n57235 ; n57235_not
g87215 not n33826 ; n33826_not
g87216 not n15493 ; n15493_not
g87217 not n34087 ; n34087_not
g87218 not n15484 ; n15484_not
g87219 not n15385 ; n15385_not
g87220 not n15376 ; n15376_not
g87221 not n15754 ; n15754_not
g87222 not n15367 ; n15367_not
g87223 not n15358 ; n15358_not
g87224 not n15349 ; n15349_not
g87225 not n33637 ; n33637_not
g87226 not n52681 ; n52681_not
g87227 not n15781 ; n15781_not
g87228 not n33646 ; n33646_not
g87229 not n33655 ; n33655_not
g87230 not n27184 ; n27184_not
g87231 not n36166 ; n36166_not
g87232 not n26392 ; n26392_not
g87233 not n26356 ; n26356_not
g87234 not n33934 ; n33934_not
g87235 not n15457 ; n15457_not
g87236 not n15709 ; n15709_not
g87237 not n33943 ; n33943_not
g87238 not n15448 ; n15448_not
g87239 not n33952 ; n33952_not
g87240 not n33961 ; n33961_not
g87241 not n15439 ; n15439_not
g87242 not n33970 ; n33970_not
g87243 not n56830 ; n56830_not
g87244 not n15394 ; n15394_not
g87245 not n26383 ; n26383_not
g87246 not n57244 ; n57244_not
g87247 not n57172 ; n57172_not
g87248 not n34294 ; n34294_not
g87249 not n34285 ; n34285_not
g87250 not n48910 ; n48910_not
g87251 not n57190 ; n57190_not
g87252 not n34276 ; n34276_not
g87253 not n26509 ; n26509_not
g87254 not n34267 ; n34267_not
g87255 not n15592 ; n15592_not
g87256 not n26365 ; n26365_not
g87257 not n15556 ; n15556_not
g87258 not n34393 ; n34393_not
g87259 not n57163 ; n57163_not
g87260 not n15565 ; n15565_not
g87261 not n15574 ; n15574_not
g87262 not n34375 ; n34375_not
g87263 not n24646 ; n24646_not
g87264 not n15583 ; n15583_not
g87265 not n34357 ; n34357_not
g87266 not n34348 ; n34348_not
g87267 not n34339 ; n34339_not
g87268 not n57217 ; n57217_not
g87269 not n34096 ; n34096_not
g87270 not n56821 ; n56821_not
g87271 not n34177 ; n34177_not
g87272 not n15547 ; n15547_not
g87273 not n55138 ; n55138_not
g87274 not n34168 ; n34168_not
g87275 not n34159 ; n34159_not
g87276 not n15538 ; n15538_not
g87277 not n33772 ; n33772_not
g87278 not n15664 ; n15664_not
g87279 not n24655 ; n24655_not
g87280 not n15529 ; n15529_not
g87281 not n34258 ; n34258_not
g87282 not n34249 ; n34249_not
g87283 not n27139 ; n27139_not
g87284 not n48901 ; n48901_not
g87285 not n34195 ; n34195_not
g87286 not n34186 ; n34186_not
g87287 not n33556 ; n33556_not
g87288 not n48820 ; n48820_not
g87289 not n24565 ; n24565_not
g87290 not n27292 ; n27292_not
g87291 not n33547 ; n33547_not
g87292 not n24556 ; n24556_not
g87293 not n33538 ; n33538_not
g87294 not n33529 ; n33529_not
g87295 not n24538 ; n24538_not
g87296 not n48811 ; n48811_not
g87297 not n24493 ; n24493_not
g87298 not n33592 ; n33592_not
g87299 not n27274 ; n27274_not
g87300 not n57370 ; n57370_not
g87301 not n26428 ; n26428_not
g87302 not n24628 ; n24628_not
g87303 not n33583 ; n33583_not
g87304 not n56920 ; n56920_not
g87305 not n33574 ; n33574_not
g87306 not n27283 ; n27283_not
g87307 not n26437 ; n26437_not
g87308 not n36193 ; n36193_not
g87309 not n24583 ; n24583_not
g87310 not n33565 ; n33565_not
g87311 not n26446 ; n26446_not
g87312 not n57406 ; n57406_not
g87313 not n33358 ; n33358_not
g87314 not n15790 ; n15790_not
g87315 not n26464 ; n26464_not
g87316 not n24448 ; n24448_not
g87317 not n36184 ; n36184_not
g87318 not n27319 ; n27319_not
g87319 not n50359 ; n50359_not
g87320 not n57460 ; n57460_not
g87321 not n36247 ; n36247_not
g87322 not n24394 ; n24394_not
g87323 not n27328 ; n27328_not
g87324 not n24385 ; n24385_not
g87325 not n26473 ; n26473_not
g87326 not n57433 ; n57433_not
g87327 not n33493 ; n33493_not
g87328 not n26455 ; n26455_not
g87329 not n33484 ; n33484_not
g87330 not n57442 ; n57442_not
g87331 not n33475 ; n33475_not
g87332 not n24475 ; n24475_not
g87333 not n33466 ; n33466_not
g87334 not n24466 ; n24466_not
g87335 not n36238 ; n36238_not
g87336 not n33457 ; n33457_not
g87337 not n33448 ; n33448_not
g87338 not n27175 ; n27175_not
g87339 not n57451 ; n57451_not
g87340 not n33439 ; n33439_not
g87341 not n24691 ; n24691_not
g87342 not n57307 ; n57307_not
g87343 not n33727 ; n33727_not
g87344 not n33763 ; n33763_not
g87345 not n24673 ; n24673_not
g87346 not n27238 ; n27238_not
g87347 not n33745 ; n33745_not
g87348 not n26347 ; n26347_not
g87349 not n33736 ; n33736_not
g87350 not n15295 ; n15295_not
g87351 not n15286 ; n15286_not
g87352 not n15277 ; n15277_not
g87353 not n15268 ; n15268_not
g87354 not n15259 ; n15259_not
g87355 not n15817 ; n15817_not
g87356 not n15826 ; n15826_not
g87357 not n57262 ; n57262_not
g87358 not n33682 ; n33682_not
g87359 not n15844 ; n15844_not
g87360 not n15853 ; n15853_not
g87361 not n52672 ; n52672_not
g87362 not n26491 ; n26491_not
g87363 not n33691 ; n33691_not
g87364 not n26482 ; n26482_not
g87365 not n33664 ; n33664_not
g87366 not n27265 ; n27265_not
g87367 not n33619 ; n33619_not
g87368 not n56911 ; n56911_not
g87369 not n57316 ; n57316_not
g87370 not n33754 ; n33754_not
g87371 not n15835 ; n15835_not
g87372 not n57334 ; n57334_not
g87373 not n51826 ; n51826_not
g87374 not n27247 ; n27247_not
g87375 not n52663 ; n52663_not
g87376 not n26419 ; n26419_not
g87377 not n33709 ; n33709_not
g87378 not n27256 ; n27256_not
g87379 not n57361 ; n57361_not
g87380 not n26257 ; n26257_not
g87381 not n24484 ; n24484_not
g87382 not n56740 ; n56740_not
g87383 not n14980 ; n14980_not
g87384 not n26266 ; n26266_not
g87385 not n34807 ; n34807_not
g87386 not n26536 ; n26536_not
g87387 not n51781 ; n51781_not
g87388 not n56803 ; n56803_not
g87389 not n25258 ; n25258_not
g87390 not n49018 ; n49018_not
g87391 not n34852 ; n34852_not
g87392 not n56713 ; n56713_not
g87393 not n24439 ; n24439_not
g87394 not n56731 ; n56731_not
g87395 not n55048 ; n55048_not
g87396 not n49009 ; n49009_not
g87397 not n49423 ; n49423_not
g87398 not n15079 ; n15079_not
g87399 not n35626 ; n35626_not
g87400 not n15097 ; n15097_not
g87401 not n26284 ; n26284_not
g87402 not n34384 ; n34384_not
g87403 not n52708 ; n52708_not
g87404 not n15169 ; n15169_not
g87405 not n15187 ; n15187_not
g87406 not n26527 ; n26527_not
g87407 not n26275 ; n26275_not
g87408 not n24529 ; n24529_not
g87409 not n52690 ; n52690_not
g87410 not n34762 ; n34762_not
g87411 not n49900 ; n49900_not
g87412 not n25393 ; n25393_not
g87413 not n55831 ; n55831_not
g87414 not n34942 ; n34942_not
g87415 not n52645 ; n52645_not
g87416 not n35950 ; n35950_not
g87417 not n26554 ; n26554_not
g87418 not n26239 ; n26239_not
g87419 not n34933 ; n34933_not
g87420 not n34915 ; n34915_not
g87421 not n49702 ; n49702_not
g87422 not n35941 ; n35941_not
g87423 not n14485 ; n14485_not
g87424 not n26194 ; n26194_not
g87425 not n49711 ; n49711_not
g87426 not n26563 ; n26563_not
g87427 not n34951 ; n34951_not
g87428 not n49720 ; n49720_not
g87429 not n49045 ; n49045_not
g87430 not n26545 ; n26545_not
g87431 not n14395 ; n14395_not
g87432 not n49801 ; n49801_not
g87433 not n49810 ; n49810_not
g87434 not n49036 ; n49036_not
g87435 not n34924 ; n34924_not
g87436 not n34906 ; n34906_not
g87437 not n49027 ; n49027_not
g87438 not n25348 ; n25348_not
g87439 not n27049 ; n27049_not
g87440 not n57073 ; n57073_not
g87441 not n55093 ; n55093_not
g87442 not n34429 ; n34429_not
g87443 not n27094 ; n27094_not
g87444 not n36076 ; n36076_not
g87445 not n57118 ; n57118_not
g87446 not n57082 ; n57082_not
g87447 not n26329 ; n26329_not
g87448 not n15088 ; n15088_not
g87449 not n34474 ; n34474_not
g87450 not n57091 ; n57091_not
g87451 not n34465 ; n34465_not
g87452 not n26518 ; n26518_not
g87453 not n51646 ; n51646_not
g87454 not n24619 ; n24619_not
g87455 not n34456 ; n34456_not
g87456 not n49333 ; n49333_not
g87457 not n34438 ; n34438_not
g87458 not n57019 ; n57019_not
g87459 not n57028 ; n57028_not
g87460 not n57154 ; n57154_not
g87461 not n56704 ; n56704_not
g87462 not n52717 ; n52717_not
g87463 not n15178 ; n15178_not
g87464 not n48721 ; n48721_not
g87465 not n57046 ; n57046_not
g87466 not n51916 ; n51916_not
g87467 not n57145 ; n57145_not
g87468 not n24574 ; n24574_not
g87469 not n34483 ; n34483_not
g87470 not n52727 ; n52727_not
g87471 not n26249 ; n26249_not
g87472 not n26087 ; n26087_not
g87473 not n22397 ; n22397_not
g87474 not n39506 ; n39506_not
g87475 not n40559 ; n40559_not
g87476 not n39443 ; n39443_not
g87477 not n39920 ; n39920_not
g87478 not n21677 ; n21677_not
g87479 not n25592 ; n25592_not
g87480 not n21884 ; n21884_not
g87481 not n25538 ; n25538_not
g87482 not n26096 ; n26096_not
g87483 not n25628 ; n25628_not
g87484 not n25286 ; n25286_not
g87485 not n53249 ; n53249_not
g87486 not n39533 ; n39533_not
g87487 not n26438 ; n26438_not
g87488 not n45806 ; n45806_not
g87489 not n26465 ; n26465_not
g87490 not n53348 ; n53348_not
g87491 not n26186 ; n26186_not
g87492 not n21839 ; n21839_not
g87493 not n21866 ; n21866_not
g87494 not n21875 ; n21875_not
g87495 not n25943 ; n25943_not
g87496 not n25952 ; n25952_not
g87497 not n39911 ; n39911_not
g87498 not n21299 ; n21299_not
g87499 not n45725 ; n45725_not
g87500 not n25619 ; n25619_not
g87501 not n20498 ; n20498_not
g87502 not n39515 ; n39515_not
g87503 not n26456 ; n26456_not
g87504 not n26159 ; n26159_not
g87505 not n21848 ; n21848_not
g87506 not n40595 ; n40595_not
g87507 not n45815 ; n45815_not
g87508 not n25871 ; n25871_not
g87509 not n21659 ; n21659_not
g87510 not n26177 ; n26177_not
g87511 not n26339 ; n26339_not
g87512 not n40568 ; n40568_not
g87513 not n25880 ; n25880_not
g87514 not n21389 ; n21389_not
g87515 not n26366 ; n26366_not
g87516 not n26447 ; n26447_not
g87517 not n52376 ; n52376_not
g87518 not n45716 ; n45716_not
g87519 not n21983 ; n21983_not
g87520 not n39614 ; n39614_not
g87521 not n39542 ; n39542_not
g87522 not n21992 ; n21992_not
g87523 not n21668 ; n21668_not
g87524 not n39452 ; n39452_not
g87525 not n26357 ; n26357_not
g87526 not n52367 ; n52367_not
g87527 not n21974 ; n21974_not
g87528 not n21857 ; n21857_not
g87529 not n40676 ; n40676_not
g87530 not n25916 ; n25916_not
g87531 not n26276 ; n26276_not
g87532 not n39425 ; n39425_not
g87533 not n21947 ; n21947_not
g87534 not n52358 ; n52358_not
g87535 not n26393 ; n26393_not
g87536 not n26294 ; n26294_not
g87537 not n26267 ; n26267_not
g87538 not n45770 ; n45770_not
g87539 not n21749 ; n21749_not
g87540 not n25556 ; n25556_not
g87541 not n45851 ; n45851_not
g87542 not n51638 ; n51638_not
g87543 not n40685 ; n40685_not
g87544 not n51647 ; n51647_not
g87545 not n21929 ; n21929_not
g87546 not n39470 ; n39470_not
g87547 not n25259 ; n25259_not
g87548 not n21785 ; n21785_not
g87549 not n21587 ; n21587_not
g87550 not n45833 ; n45833_not
g87551 not n21767 ; n21767_not
g87552 not n45761 ; n45761_not
g87553 not n21578 ; n21578_not
g87554 not n45455 ; n45455_not
g87555 not n22298 ; n22298_not
g87556 not n52394 ; n52394_not
g87557 not n41198 ; n41198_not
g87558 not n25925 ; n25925_not
g87559 not n21398 ; n21398_not
g87560 not n40667 ; n40667_not
g87561 not n21758 ; n21758_not
g87562 not n26384 ; n26384_not
g87563 not n22289 ; n22289_not
g87564 not n25970 ; n25970_not
g87565 not n45680 ; n45680_not
g87566 not n25547 ; n25547_not
g87567 not n21569 ; n21569_not
g87568 not n21776 ; n21776_not
g87569 not n21938 ; n21938_not
g87570 not n52448 ; n52448_not
g87571 not n21695 ; n21695_not
g87572 not n22199 ; n22199_not
g87573 not n22388 ; n22388_not
g87574 not n21893 ; n21893_not
g87575 not n25583 ; n25583_not
g87576 not n21794 ; n21794_not
g87577 not n52349 ; n52349_not
g87578 not n39434 ; n39434_not
g87579 not n21686 ; n21686_not
g87580 not n45743 ; n45743_not
g87581 not n52457 ; n52457_not
g87582 not n21479 ; n21479_not
g87583 not n26069 ; n26069_not
g87584 not n51656 ; n51656_not
g87585 not n21488 ; n21488_not
g87586 not n53276 ; n53276_not
g87587 not n21965 ; n21965_not
g87588 not n52475 ; n52475_not
g87589 not n39407 ; n39407_not
g87590 not n26429 ; n26429_not
g87591 not n40586 ; n40586_not
g87592 not n22379 ; n22379_not
g87593 not n52385 ; n52385_not
g87594 not n20795 ; n20795_not
g87595 not n53285 ; n53285_not
g87596 not n45860 ; n45860_not
g87597 not n25907 ; n25907_not
g87598 not n39416 ; n39416_not
g87599 not n21956 ; n21956_not
g87600 not n40577 ; n40577_not
g87601 not n41189 ; n41189_not
g87602 not n25934 ; n25934_not
g87603 not n25295 ; n25295_not
g87604 not n25565 ; n25565_not
g87605 not n39461 ; n39461_not
g87606 not n26375 ; n26375_not
g87607 not n25961 ; n25961_not
g87608 not n21497 ; n21497_not
g87609 not n21596 ; n21596_not
g87610 not n25574 ; n25574_not
g87611 not n53258 ; n53258_not
g87612 not n40829 ; n40829_not
g87613 not n40469 ; n40469_not
g87614 not n23927 ; n23927_not
g87615 not n52547 ; n52547_not
g87616 not n23864 ; n23864_not
g87617 not n24953 ; n24953_not
g87618 not n23936 ; n23936_not
g87619 not n24944 ; n24944_not
g87620 not n24566 ; n24566_not
g87621 not n23945 ; n23945_not
g87622 not n52556 ; n52556_not
g87623 not n40478 ; n40478_not
g87624 not n24935 ; n24935_not
g87625 not n23954 ; n23954_not
g87626 not n23189 ; n23189_not
g87627 not n52718 ; n52718_not
g87628 not n52682 ; n52682_not
g87629 not n51971 ; n51971_not
g87630 not n51962 ; n51962_not
g87631 not n51953 ; n51953_not
g87632 not n24539 ; n24539_not
g87633 not n23882 ; n23882_not
g87634 not n23909 ; n23909_not
g87635 not n39740 ; n39740_not
g87636 not n51944 ; n51944_not
g87637 not n24980 ; n24980_not
g87638 not n51935 ; n51935_not
g87639 not n23873 ; n23873_not
g87640 not n24971 ; n24971_not
g87641 not n51926 ; n51926_not
g87642 not n23918 ; n23918_not
g87643 not n24962 ; n24962_not
g87644 not n23981 ; n23981_not
g87645 not n23837 ; n23837_not
g87646 not n23990 ; n23990_not
g87647 not n40784 ; n40784_not
g87648 not n52736 ; n52736_not
g87649 not n24872 ; n24872_not
g87650 not n23828 ; n23828_not
g87651 not n24863 ; n24863_not
g87652 not n52970 ; n52970_not
g87653 not n24854 ; n24854_not
g87654 not n23819 ; n23819_not
g87655 not n24845 ; n24845_not
g87656 not n24926 ; n24926_not
g87657 not n24575 ; n24575_not
g87658 not n24917 ; n24917_not
g87659 not n24584 ; n24584_not
g87660 not n23963 ; n23963_not
g87661 not n40487 ; n40487_not
g87662 not n45554 ; n45554_not
g87663 not n23198 ; n23198_not
g87664 not n24908 ; n24908_not
g87665 not n23972 ; n23972_not
g87666 not n24890 ; n24890_not
g87667 not n45518 ; n45518_not
g87668 not n45077 ; n45077_not
g87669 not n40496 ; n40496_not
g87670 not n24881 ; n24881_not
g87671 not n40397 ; n40397_not
g87672 not n25385 ; n25385_not
g87673 not n40847 ; n40847_not
g87674 not n25376 ; n25376_not
g87675 not n23846 ; n23846_not
g87676 not n52655 ; n52655_not
g87677 not n40289 ; n40289_not
g87678 not n23288 ; n23288_not
g87679 not n23279 ; n23279_not
g87680 not n40388 ; n40388_not
g87681 not n52628 ; n52628_not
g87682 not n52637 ; n52637_not
g87683 not n40865 ; n40865_not
g87684 not n25169 ; n25169_not
g87685 not n24449 ; n24449_not
g87686 not n24476 ; n24476_not
g87687 not n52538 ; n52538_not
g87688 not n25097 ; n25097_not
g87689 not n25088 ; n25088_not
g87690 not n24485 ; n24485_not
g87691 not n52673 ; n52673_not
g87692 not n25079 ; n25079_not
g87693 not n24494 ; n24494_not
g87694 not n40838 ; n40838_not
g87695 not n51980 ; n51980_not
g87696 not n45563 ; n45563_not
g87697 not n23891 ; n23891_not
g87698 not n45572 ; n45572_not
g87699 not n40199 ; n40199_not
g87700 not n40856 ; n40856_not
g87701 not n25358 ; n25358_not
g87702 not n25268 ; n25268_not
g87703 not n25178 ; n25178_not
g87704 not n25187 ; n25187_not
g87705 not n25196 ; n25196_not
g87706 not n24665 ; n24665_not
g87707 not n23684 ; n23684_not
g87708 not n24656 ; n24656_not
g87709 not n23495 ; n23495_not
g87710 not n24269 ; n24269_not
g87711 not n52871 ; n52871_not
g87712 not n52817 ; n52817_not
g87713 not n24638 ; n24638_not
g87714 not n24278 ; n24278_not
g87715 not n24287 ; n24287_not
g87716 not n40649 ; n40649_not
g87717 not n52790 ; n52790_not
g87718 not n40694 ; n40694_not
g87719 not n23459 ; n23459_not
g87720 not n24683 ; n24683_not
g87721 not n23468 ; n23468_not
g87722 not n23693 ; n23693_not
g87723 not n23477 ; n23477_not
g87724 not n52880 ; n52880_not
g87725 not n52808 ; n52808_not
g87726 not n23486 ; n23486_not
g87727 not n23567 ; n23567_not
g87728 not n23639 ; n23639_not
g87729 not n23576 ; n23576_not
g87730 not n45086 ; n45086_not
g87731 not n52844 ; n52844_not
g87732 not n24458 ; n24458_not
g87733 not n23585 ; n23585_not
g87734 not n24359 ; n24359_not
g87735 not n23594 ; n23594_not
g87736 not n24368 ; n24368_not
g87737 not n52835 ; n52835_not
g87738 not n24386 ; n24386_not
g87739 not n24377 ; n24377_not
g87740 not n52862 ; n52862_not
g87741 not n24296 ; n24296_not
g87742 not n24593 ; n24593_not
g87743 not n23657 ; n23657_not
g87744 not n52853 ; n52853_not
g87745 not n52826 ; n52826_not
g87746 not n23549 ; n23549_not
g87747 not n23648 ; n23648_not
g87748 not n24548 ; n24548_not
g87749 not n23558 ; n23558_not
g87750 not n52646 ; n52646_not
g87751 not n52943 ; n52943_not
g87752 not n52754 ; n52754_not
g87753 not n24791 ; n24791_not
g87754 not n23792 ; n23792_not
g87755 not n23783 ; n23783_not
g87756 not n52592 ; n52592_not
g87757 not n52934 ; n52934_not
g87758 not n24089 ; n24089_not
g87759 not n40739 ; n40739_not
g87760 not n24782 ; n24782_not
g87761 not n23774 ; n23774_not
g87762 not n24098 ; n24098_not
g87763 not n52925 ; n52925_not
g87764 not n52763 ; n52763_not
g87765 not n52961 ; n52961_not
g87766 not n24836 ; n24836_not
g87767 not n40766 ; n40766_not
g87768 not n24629 ; n24629_not
g87769 not n45545 ; n45545_not
g87770 not n52583 ; n52583_not
g87771 not n24827 ; n24827_not
g87772 not n40757 ; n40757_not
g87773 not n52952 ; n52952_not
g87774 not n24818 ; n24818_not
g87775 not n52745 ; n52745_not
g87776 not n24809 ; n24809_not
g87777 not n23297 ; n23297_not
g87778 not n24179 ; n24179_not
g87779 not n24755 ; n24755_not
g87780 not n24674 ; n24674_not
g87781 not n24746 ; n24746_not
g87782 not n52781 ; n52781_not
g87783 not n24737 ; n24737_not
g87784 not n24728 ; n24728_not
g87785 not n45536 ; n45536_not
g87786 not n24188 ; n24188_not
g87787 not n45527 ; n45527_not
g87788 not n24719 ; n24719_not
g87789 not n24197 ; n24197_not
g87790 not n52916 ; n52916_not
g87791 not n52691 ; n52691_not
g87792 not n23369 ; n23369_not
g87793 not n23378 ; n23378_not
g87794 not n23747 ; n23747_not
g87795 not n24773 ; n24773_not
g87796 not n23387 ; n23387_not
g87797 not n23738 ; n23738_not
g87798 not n45095 ; n45095_not
g87799 not n23396 ; n23396_not
g87800 not n52772 ; n52772_not
g87801 not n52907 ; n52907_not
g87802 not n23729 ; n23729_not
g87803 not n24764 ; n24764_not
g87804 not n22838 ; n22838_not
g87805 not n25745 ; n25745_not
g87806 not n22856 ; n22856_not
g87807 not n25736 ; n25736_not
g87808 not n45617 ; n45617_not
g87809 not n53159 ; n53159_not
g87810 not n25727 ; n25727_not
g87811 not n25718 ; n25718_not
g87812 not n22874 ; n22874_not
g87813 not n25709 ; n25709_not
g87814 not n22883 ; n22883_not
g87815 not n25763 ; n25763_not
g87816 not n45626 ; n45626_not
g87817 not n22775 ; n22775_not
g87818 not n22784 ; n22784_not
g87819 not n45464 ; n45464_not
g87820 not n22793 ; n22793_not
g87821 not n52466 ; n52466_not
g87822 not n25754 ; n25754_not
g87823 not n53168 ; n53168_not
g87824 not n22829 ; n22829_not
g87825 not n22991 ; n22991_not
g87826 not n25664 ; n25664_not
g87827 not n40298 ; n40298_not
g87828 not n23099 ; n23099_not
g87829 not n52187 ; n52187_not
g87830 not n25655 ; n25655_not
g87831 not n52565 ; n52565_not
g87832 not n52493 ; n52493_not
g87833 not n22982 ; n22982_not
g87834 not n45473 ; n45473_not
g87835 not n45608 ; n45608_not
g87836 not n25691 ; n25691_not
g87837 not n22919 ; n22919_not
g87838 not n22928 ; n22928_not
g87839 not n25439 ; n25439_not
g87840 not n22946 ; n22946_not
g87841 not n25682 ; n25682_not
g87842 not n52196 ; n52196_not
g87843 not n22964 ; n22964_not
g87844 not n25673 ; n25673_not
g87845 not n22973 ; n22973_not
g87846 not n52295 ; n52295_not
g87847 not n45653 ; n45653_not
g87848 not n25826 ; n25826_not
g87849 not n22568 ; n22568_not
g87850 not n22577 ; n22577_not
g87851 not n25817 ; n25817_not
g87852 not n22586 ; n22586_not
g87853 not n41099 ; n41099_not
g87854 not n25808 ; n25808_not
g87855 not n45644 ; n45644_not
g87856 not n22595 ; n22595_not
g87857 not n53195 ; n53195_not
g87858 not n22469 ; n22469_not
g87859 not n45662 ; n45662_not
g87860 not n39902 ; n39902_not
g87861 not n22478 ; n22478_not
g87862 not n25862 ; n25862_not
g87863 not n22487 ; n22487_not
g87864 not n22496 ; n22496_not
g87865 not n25853 ; n25853_not
g87866 not n25349 ; n25349_not
g87867 not n25844 ; n25844_not
g87868 not n22559 ; n22559_not
g87869 not n25835 ; n25835_not
g87870 not n22685 ; n22685_not
g87871 not n22694 ; n22694_not
g87872 not n39812 ; n39812_not
g87873 not n52259 ; n52259_not
g87874 not n25772 ; n25772_not
g87875 not n22739 ; n22739_not
g87876 not n53177 ; n53177_not
g87877 not n22748 ; n22748_not
g87878 not n22757 ; n22757_not
g87879 not n39803 ; n39803_not
g87880 not n25394 ; n25394_not
g87881 not n22766 ; n22766_not
g87882 not n52286 ; n52286_not
g87883 not n52277 ; n52277_not
g87884 not n25790 ; n25790_not
g87885 not n22649 ; n22649_not
g87886 not n39830 ; n39830_not
g87887 not n45635 ; n45635_not
g87888 not n22658 ; n22658_not
g87889 not n22667 ; n22667_not
g87890 not n39821 ; n39821_not
g87891 not n53186 ; n53186_not
g87892 not n22676 ; n22676_not
g87893 not n52268 ; n52268_not
g87894 not n25781 ; n25781_not
g87895 not n40892 ; n40892_not
g87896 not n45509 ; n45509_not
g87897 not n23666 ; n23666_not
g87898 not n25475 ; n25475_not
g87899 not n25466 ; n25466_not
g87900 not n40874 ; n40874_not
g87901 not n40379 ; n40379_not
g87902 not n45581 ; n45581_not
g87903 not n52079 ; n52079_not
g87904 not n25448 ; n25448_not
g87905 not n40883 ; n40883_not
g87906 not n23756 ; n23756_not
g87907 not n25493 ; n25493_not
g87908 not n52097 ; n52097_not
g87909 not n52088 ; n52088_not
g87910 not n40775 ; n40775_not
g87911 not n53096 ; n53096_not
g87912 not n45482 ; n45482_not
g87913 not n40964 ; n40964_not
g87914 not n52169 ; n52169_not
g87915 not n53087 ; n53087_not
g87916 not n40955 ; n40955_not
g87917 not n22892 ; n22892_not
g87918 not n25646 ; n25646_not
g87919 not n40991 ; n40991_not
g87920 not n52178 ; n52178_not
g87921 not n25637 ; n25637_not
g87922 not n40982 ; n40982_not
g87923 not n22937 ; n22937_not
g87924 not n40973 ; n40973_not
g87925 not n40928 ; n40928_not
g87926 not n45590 ; n45590_not
g87927 not n40919 ; n40919_not
g87928 not n25484 ; n25484_not
g87929 not n45491 ; n45491_not
g87930 not n40946 ; n40946_not
g87931 not n53078 ; n53078_not
g87932 not n40937 ; n40937_not
g87933 not n53069 ; n53069_not
g87934 not n22847 ; n22847_not
g87935 not n43628 ; n43628_not
g87936 not n14828 ; n14828_not
g87937 not n14837 ; n14837_not
g87938 not n55247 ; n55247_not
g87939 not n14846 ; n14846_not
g87940 not n14855 ; n14855_not
g87941 not n43619 ; n43619_not
g87942 not n14864 ; n14864_not
g87943 not n55607 ; n55607_not
g87944 not n14873 ; n14873_not
g87945 not n14396 ; n14396_not
g87946 not n14882 ; n14882_not
g87947 not n14891 ; n14891_not
g87948 not n43097 ; n43097_not
g87949 not n14387 ; n14387_not
g87950 not n14909 ; n14909_not
g87951 not n43592 ; n43592_not
g87952 not n14918 ; n14918_not
g87953 not n14927 ; n14927_not
g87954 not n14936 ; n14936_not
g87955 not n44960 ; n44960_not
g87956 not n55580 ; n55580_not
g87957 not n55652 ; n55652_not
g87958 not n14495 ; n14495_not
g87959 not n43664 ; n43664_not
g87960 not n14486 ; n14486_not
g87961 not n14729 ; n14729_not
g87962 not n14477 ; n14477_not
g87963 not n14738 ; n14738_not
g87964 not n55643 ; n55643_not
g87965 not n43655 ; n43655_not
g87966 not n14747 ; n14747_not
g87967 not n14756 ; n14756_not
g87968 not n14765 ; n14765_not
g87969 not n55634 ; n55634_not
g87970 not n43646 ; n43646_not
g87971 not n14774 ; n14774_not
g87972 not n14783 ; n14783_not
g87973 not n55625 ; n55625_not
g87974 not n43637 ; n43637_not
g87975 not n14792 ; n14792_not
g87976 not n14819 ; n14819_not
g87977 not n55616 ; n55616_not
g87978 not n42944 ; n42944_not
g87979 not n55544 ; n55544_not
g87980 not n43538 ; n43538_not
g87981 not n55535 ; n55535_not
g87982 not n42935 ; n42935_not
g87983 not n15089 ; n15089_not
g87984 not n43529 ; n43529_not
g87985 not n55526 ; n55526_not
g87986 not n42926 ; n42926_not
g87987 not n15179 ; n15179_not
g87988 not n15197 ; n15197_not
g87989 not n42917 ; n42917_not
g87990 not n55517 ; n55517_not
g87991 not n15188 ; n15188_not
g87992 not n42908 ; n42908_not
g87993 not n44933 ; n44933_not
g87994 not n55508 ; n55508_not
g87995 not n45059 ; n45059_not
g87996 not n43583 ; n43583_not
g87997 not n14945 ; n14945_not
g87998 not n42980 ; n42980_not
g87999 not n14954 ; n14954_not
g88000 not n44951 ; n44951_not
g88001 not n43574 ; n43574_not
g88002 not n14963 ; n14963_not
g88003 not n42971 ; n42971_not
g88004 not n55571 ; n55571_not
g88005 not n14972 ; n14972_not
g88006 not n43565 ; n43565_not
g88007 not n55049 ; n55049_not
g88008 not n42962 ; n42962_not
g88009 not n14981 ; n14981_not
g88010 not n55562 ; n55562_not
g88011 not n43556 ; n43556_not
g88012 not n42953 ; n42953_not
g88013 not n55058 ; n55058_not
g88014 not n44942 ; n44942_not
g88015 not n55553 ; n55553_not
g88016 not n14990 ; n14990_not
g88017 not n43547 ; n43547_not
g88018 not n44582 ; n44582_not
g88019 not n43844 ; n43844_not
g88020 not n55805 ; n55805_not
g88021 not n13892 ; n13892_not
g88022 not n43826 ; n43826_not
g88023 not n44348 ; n44348_not
g88024 not n54923 ; n54923_not
g88025 not n13865 ; n13865_not
g88026 not n13856 ; n13856_not
g88027 not n13847 ; n13847_not
g88028 not n43808 ; n43808_not
g88029 not n55760 ; n55760_not
g88030 not n55751 ; n55751_not
g88031 not n54950 ; n54950_not
g88032 not n55742 ; n55742_not
g88033 not n13775 ; n13775_not
g88034 not n13766 ; n13766_not
g88035 not n43916 ; n43916_not
g88036 not n13784 ; n13784_not
g88037 not n43277 ; n43277_not
g88038 not n42674 ; n42674_not
g88039 not n13829 ; n13829_not
g88040 not n13874 ; n13874_not
g88041 not n55850 ; n55850_not
g88042 not n13919 ; n13919_not
g88043 not n43871 ; n43871_not
g88044 not n13937 ; n13937_not
g88045 not n13946 ; n13946_not
g88046 not n13955 ; n13955_not
g88047 not n55832 ; n55832_not
g88048 not n43853 ; n43853_not
g88049 not n55823 ; n55823_not
g88050 not n44357 ; n44357_not
g88051 not n43718 ; n43718_not
g88052 not n14585 ; n14585_not
g88053 not n14594 ; n14594_not
g88054 not n43709 ; n43709_not
g88055 not n55706 ; n55706_not
g88056 not n14639 ; n14639_not
g88057 not n14648 ; n14648_not
g88058 not n14657 ; n14657_not
g88059 not n43691 ; n43691_not
g88060 not n14666 ; n14666_not
g88061 not n43682 ; n43682_not
g88062 not n14675 ; n14675_not
g88063 not n55670 ; n55670_not
g88064 not n14684 ; n14684_not
g88065 not n55661 ; n55661_not
g88066 not n14693 ; n14693_not
g88067 not n43673 ; n43673_not
g88068 not n13757 ; n13757_not
g88069 not n55733 ; n55733_not
g88070 not n43781 ; n43781_not
g88071 not n14369 ; n14369_not
g88072 not n44339 ; n44339_not
g88073 not n43763 ; n43763_not
g88074 not n14459 ; n14459_not
g88075 not n43754 ; n43754_not
g88076 not n55724 ; n55724_not
g88077 not n14549 ; n14549_not
g88078 not n43736 ; n43736_not
g88079 not n55715 ; n55715_not
g88080 not n14567 ; n14567_not
g88081 not n15944 ; n15944_not
g88082 not n43259 ; n43259_not
g88083 not n15863 ; n15863_not
g88084 not n15953 ; n15953_not
g88085 not n15791 ; n15791_not
g88086 not n42719 ; n42719_not
g88087 not n55346 ; n55346_not
g88088 not n15962 ; n15962_not
g88089 not n42728 ; n42728_not
g88090 not n42737 ; n42737_not
g88091 not n15971 ; n15971_not
g88092 not n15782 ; n15782_not
g88093 not n42746 ; n42746_not
g88094 not n55175 ; n55175_not
g88095 not n55337 ; n55337_not
g88096 not n42755 ; n42755_not
g88097 not n55364 ; n55364_not
g88098 not n42692 ; n42692_not
g88099 not n44861 ; n44861_not
g88100 not n43286 ; n43286_not
g88101 not n15908 ; n15908_not
g88102 not n42683 ; n42683_not
g88103 not n15917 ; n15917_not
g88104 not n15926 ; n15926_not
g88105 not n44852 ; n44852_not
g88106 not n15935 ; n15935_not
g88107 not n55355 ; n55355_not
g88108 not n55319 ; n55319_not
g88109 not n42818 ; n42818_not
g88110 not n15746 ; n15746_not
g88111 not n42827 ; n42827_not
g88112 not n43187 ; n43187_not
g88113 not n42836 ; n42836_not
g88114 not n15737 ; n15737_not
g88115 not n42845 ; n42845_not
g88116 not n42854 ; n42854_not
g88117 not n42863 ; n42863_not
g88118 not n43169 ; n43169_not
g88119 not n16079 ; n16079_not
g88120 not n42872 ; n42872_not
g88121 not n15980 ; n15980_not
g88122 not n42764 ; n42764_not
g88123 not n42773 ; n42773_not
g88124 not n55328 ; n55328_not
g88125 not n42782 ; n42782_not
g88126 not n42791 ; n42791_not
g88127 not n44843 ; n44843_not
g88128 not n55184 ; n55184_not
g88129 not n42809 ; n42809_not
g88130 not n15755 ; n15755_not
g88131 not n43196 ; n43196_not
g88132 not n55454 ; n55454_not
g88133 not n43439 ; n43439_not
g88134 not n55445 ; n55445_not
g88135 not n55436 ; n55436_not
g88136 not n44906 ; n44906_not
g88137 not n55427 ; n55427_not
g88138 not n55418 ; n55418_not
g88139 not n15629 ; n15629_not
g88140 not n43394 ; n43394_not
g88141 not n15647 ; n15647_not
g88142 not n15656 ; n15656_not
g88143 not n55085 ; n55085_not
g88144 not n43493 ; n43493_not
g88145 not n42890 ; n42890_not
g88146 not n44924 ; n44924_not
g88147 not n55490 ; n55490_not
g88148 not n43484 ; n43484_not
g88149 not n42881 ; n42881_not
g88150 not n55094 ; n55094_not
g88151 not n43475 ; n43475_not
g88152 not n55481 ; n55481_not
g88153 not n44915 ; n44915_not
g88154 not n43466 ; n43466_not
g88155 not n55472 ; n55472_not
g88156 not n15098 ; n15098_not
g88157 not n43457 ; n43457_not
g88158 not n55463 ; n55463_not
g88159 not n43448 ; n43448_not
g88160 not n15809 ; n15809_not
g88161 not n15827 ; n15827_not
g88162 not n15836 ; n15836_not
g88163 not n44870 ; n44870_not
g88164 not n55382 ; n55382_not
g88165 not n15854 ; n15854_not
g88166 not n15845 ; n15845_not
g88167 not n15872 ; n15872_not
g88168 not n55373 ; n55373_not
g88169 not n15881 ; n15881_not
g88170 not n15890 ; n15890_not
g88171 not n43295 ; n43295_not
g88172 not n43385 ; n43385_not
g88173 not n15674 ; n15674_not
g88174 not n55409 ; n55409_not
g88175 not n43376 ; n43376_not
g88176 not n15692 ; n15692_not
g88177 not n43367 ; n43367_not
g88178 not n15719 ; n15719_not
g88179 not n43358 ; n43358_not
g88180 not n55139 ; n55139_not
g88181 not n15764 ; n15764_not
g88182 not n43349 ; n43349_not
g88183 not n55148 ; n55148_not
g88184 not n55391 ; n55391_not
g88185 not n56534 ; n56534_not
g88186 not n44456 ; n44456_not
g88187 not n56525 ; n56525_not
g88188 not n56516 ; n56516_not
g88189 not n56507 ; n56507_not
g88190 not n44438 ; n44438_not
g88191 not n56480 ; n56480_not
g88192 not n56471 ; n56471_not
g88193 not n44429 ; n44429_not
g88194 not n56462 ; n56462_not
g88195 not n56453 ; n56453_not
g88196 not n55913 ; n55913_not
g88197 not n56444 ; n56444_not
g88198 not n56435 ; n56435_not
g88199 not n55922 ; n55922_not
g88200 not n56633 ; n56633_not
g88201 not n44771 ; n44771_not
g88202 not n56624 ; n56624_not
g88203 not n56615 ; n56615_not
g88204 not n56606 ; n56606_not
g88205 not n44483 ; n44483_not
g88206 not n55841 ; n55841_not
g88207 not n44474 ; n44474_not
g88208 not n44780 ; n44780_not
g88209 not n56570 ; n56570_not
g88210 not n56561 ; n56561_not
g88211 not n56552 ; n56552_not
g88212 not n56543 ; n56543_not
g88213 not n56327 ; n56327_not
g88214 not n56318 ; n56318_not
g88215 not n10499 ; n10499_not
g88216 not n56309 ; n56309_not
g88217 not n10589 ; n10589_not
g88218 not n10598 ; n10598_not
g88219 not n56291 ; n56291_not
g88220 not n10679 ; n10679_not
g88221 not n10688 ; n10688_not
g88222 not n10697 ; n10697_not
g88223 not n56282 ; n56282_not
g88224 not n16277 ; n16277_not
g88225 not n56273 ; n56273_not
g88226 not n10769 ; n10769_not
g88227 not n10778 ; n10778_not
g88228 not n10787 ; n10787_not
g88229 not n10796 ; n10796_not
g88230 not n56426 ; n56426_not
g88231 not n55931 ; n55931_not
g88232 not n56417 ; n56417_not
g88233 not n56408 ; n56408_not
g88234 not n56390 ; n56390_not
g88235 not n44393 ; n44393_not
g88236 not n56381 ; n56381_not
g88237 not n44384 ; n44384_not
g88238 not n56372 ; n56372_not
g88239 not n56363 ; n56363_not
g88240 not n56354 ; n56354_not
g88241 not n56345 ; n56345_not
g88242 not n56336 ; n56336_not
g88243 not n44366 ; n44366_not
g88244 not n57308 ; n57308_not
g88245 not n44528 ; n44528_not
g88246 not n44645 ; n44645_not
g88247 not n57290 ; n57290_not
g88248 not n57281 ; n57281_not
g88249 not n44537 ; n44537_not
g88250 not n44636 ; n44636_not
g88251 not n56840 ; n56840_not
g88252 not n57254 ; n57254_not
g88253 not n44717 ; n44717_not
g88254 not n56831 ; n56831_not
g88255 not n44492 ; n44492_not
g88256 not n44627 ; n44627_not
g88257 not n57236 ; n57236_not
g88258 not n57227 ; n57227_not
g88259 not n57218 ; n57218_not
g88260 not n44618 ; n44618_not
g88261 not n57209 ; n57209_not
g88262 not n56804 ; n56804_not
g88263 not n57470 ; n57470_not
g88264 not n44690 ; n44690_not
g88265 not n57452 ; n57452_not
g88266 not n57443 ; n57443_not
g88267 not n57434 ; n57434_not
g88268 not n44681 ; n44681_not
g88269 not n57425 ; n57425_not
g88270 not n56930 ; n56930_not
g88271 not n56921 ; n56921_not
g88272 not n44672 ; n44672_not
g88273 not n57380 ; n57380_not
g88274 not n57371 ; n57371_not
g88275 not n44708 ; n44708_not
g88276 not n44519 ; n44519_not
g88277 not n44663 ; n44663_not
g88278 not n57362 ; n57362_not
g88279 not n57353 ; n57353_not
g88280 not n44654 ; n44654_not
g88281 not n57326 ; n57326_not
g88282 not n56705 ; n56705_not
g88283 not n57038 ; n57038_not
g88284 not n44744 ; n44744_not
g88285 not n56903 ; n56903_not
g88286 not n44546 ; n44546_not
g88287 not n44753 ; n44753_not
g88288 not n56813 ; n56813_not
g88289 not n44762 ; n44762_not
g88290 not n56750 ; n56750_not
g88291 not n56741 ; n56741_not
g88292 not n56723 ; n56723_not
g88293 not n56660 ; n56660_not
g88294 not n56651 ; n56651_not
g88295 not n56642 ; n56642_not
g88296 not n57182 ; n57182_not
g88297 not n57164 ; n57164_not
g88298 not n44609 ; n44609_not
g88299 not n57155 ; n57155_not
g88300 not n57146 ; n57146_not
g88301 not n57137 ; n57137_not
g88302 not n44726 ; n44726_not
g88303 not n44564 ; n44564_not
g88304 not n57092 ; n57092_not
g88305 not n57083 ; n57083_not
g88306 not n44735 ; n44735_not
g88307 not n57074 ; n57074_not
g88308 not n57065 ; n57065_not
g88309 not n44573 ; n44573_not
g88310 not n56714 ; n56714_not
g88311 not n12956 ; n12956_not
g88312 not n12965 ; n12965_not
g88313 not n12974 ; n12974_not
g88314 not n12983 ; n12983_not
g88315 not n43817 ; n43817_not
g88316 not n12992 ; n12992_not
g88317 not n12587 ; n12587_not
g88318 not n12578 ; n12578_not
g88319 not n12569 ; n12569_not
g88320 not n13298 ; n13298_not
g88321 not n12785 ; n12785_not
g88322 not n12794 ; n12794_not
g88323 not n13379 ; n13379_not
g88324 not n13388 ; n13388_not
g88325 not n13397 ; n13397_not
g88326 not n12839 ; n12839_not
g88327 not n12848 ; n12848_not
g88328 not n12857 ; n12857_not
g88329 not n12659 ; n12659_not
g88330 not n12668 ; n12668_not
g88331 not n12686 ; n12686_not
g88332 not n12749 ; n12749_not
g88333 not n56057 ; n56057_not
g88334 not n12866 ; n12866_not
g88335 not n56048 ; n56048_not
g88336 not n12875 ; n12875_not
g88337 not n12884 ; n12884_not
g88338 not n12893 ; n12893_not
g88339 not n12677 ; n12677_not
g88340 not n12929 ; n12929_not
g88341 not n12938 ; n12938_not
g88342 not n12947 ; n12947_not
g88343 not n13568 ; n13568_not
g88344 not n13577 ; n13577_not
g88345 not n55940 ; n55940_not
g88346 not n13586 ; n13586_not
g88347 not n13595 ; n13595_not
g88348 not n13649 ; n13649_not
g88349 not n13658 ; n13658_not
g88350 not n13667 ; n13667_not
g88351 not n13676 ; n13676_not
g88352 not n13685 ; n13685_not
g88353 not n13694 ; n13694_not
g88354 not n13739 ; n13739_not
g88355 not n43907 ; n43907_not
g88356 not n13469 ; n13469_not
g88357 not n13478 ; n13478_not
g88358 not n43862 ; n43862_not
g88359 not n13487 ; n13487_not
g88360 not n13496 ; n13496_not
g88361 not n13559 ; n13559_not
g88362 not n10868 ; n10868_not
g88363 not n11399 ; n11399_not
g88364 not n11498 ; n11498_not
g88365 not n11588 ; n11588_not
g88366 not n11597 ; n11597_not
g88367 not n56219 ; n56219_not
g88368 not n11669 ; n11669_not
g88369 not n11678 ; n11678_not
g88370 not n11687 ; n11687_not
g88371 not n11696 ; n11696_not
g88372 not n11759 ; n11759_not
g88373 not n11768 ; n11768_not
g88374 not n43727 ; n43727_not
g88375 not n11777 ; n11777_not
g88376 not n11786 ; n11786_not
g88377 not n56264 ; n56264_not
g88378 not n10877 ; n10877_not
g88379 not n44447 ; n44447_not
g88380 not n10895 ; n10895_not
g88381 not n10949 ; n10949_not
g88382 not n10967 ; n10967_not
g88383 not n10985 ; n10985_not
g88384 not n10994 ; n10994_not
g88385 not n56255 ; n56255_not
g88386 not n56246 ; n56246_not
g88387 not n44807 ; n44807_not
g88388 not n56237 ; n56237_not
g88389 not n10958 ; n10958_not
g88390 not n56228 ; n56228_not
g88391 not n56156 ; n56156_not
g88392 not n11993 ; n11993_not
g88393 not n55274 ; n55274_not
g88394 not n56147 ; n56147_not
g88395 not n44825 ; n44825_not
g88396 not n55265 ; n55265_not
g88397 not n56138 ; n56138_not
g88398 not n55256 ; n55256_not
g88399 not n56129 ; n56129_not
g88400 not n56093 ; n56093_not
g88401 not n55229 ; n55229_not
g88402 not n44834 ; n44834_not
g88403 not n43772 ; n43772_not
g88404 not n56075 ; n56075_not
g88405 not n12596 ; n12596_not
g88406 not n11795 ; n11795_not
g88407 not n56192 ; n56192_not
g88408 not n44816 ; n44816_not
g88409 not n56183 ; n56183_not
g88410 not n11849 ; n11849_not
g88411 not n56066 ; n56066_not
g88412 not n11858 ; n11858_not
g88413 not n11867 ; n11867_not
g88414 not n11876 ; n11876_not
g88415 not n11885 ; n11885_not
g88416 not n56174 ; n56174_not
g88417 not n11894 ; n11894_not
g88418 not n55292 ; n55292_not
g88419 not n11939 ; n11939_not
g88420 not n56165 ; n56165_not
g88421 not n11948 ; n11948_not
g88422 not n11957 ; n11957_not
g88423 not n11975 ; n11975_not
g88424 not n11984 ; n11984_not
g88425 not n55283 ; n55283_not
g88426 not n54473 ; n54473_not
g88427 not n54392 ; n54392_not
g88428 not n41981 ; n41981_not
g88429 not n54464 ; n54464_not
g88430 not n18581 ; n18581_not
g88431 not n18608 ; n18608_not
g88432 not n18563 ; n18563_not
g88433 not n18617 ; n18617_not
g88434 not n18554 ; n18554_not
g88435 not n54455 ; n54455_not
g88436 not n18626 ; n18626_not
g88437 not n45329 ; n45329_not
g88438 not n18635 ; n18635_not
g88439 not n18545 ; n18545_not
g88440 not n18644 ; n18644_not
g88441 not n54446 ; n54446_not
g88442 not n18653 ; n18653_not
g88443 not n18662 ; n18662_not
g88444 not n54437 ; n54437_not
g88445 not n18671 ; n18671_not
g88446 not n18419 ; n18419_not
g88447 not n18437 ; n18437_not
g88448 not n18455 ; n18455_not
g88449 not n54527 ; n54527_not
g88450 not n18464 ; n18464_not
g88451 not n18482 ; n18482_not
g88452 not n54518 ; n54518_not
g88453 not n18509 ; n18509_not
g88454 not n54509 ; n54509_not
g88455 not n18527 ; n18527_not
g88456 not n41963 ; n41963_not
g88457 not n54491 ; n54491_not
g88458 not n17870 ; n17870_not
g88459 not n54482 ; n54482_not
g88460 not n41972 ; n41972_not
g88461 not n54329 ; n54329_not
g88462 not n18473 ; n18473_not
g88463 not n54356 ; n54356_not
g88464 not n54338 ; n54338_not
g88465 not n18806 ; n18806_not
g88466 not n18815 ; n18815_not
g88467 not n18824 ; n18824_not
g88468 not n18833 ; n18833_not
g88469 not n41990 ; n41990_not
g88470 not n18842 ; n18842_not
g88471 not n18851 ; n18851_not
g88472 not n18428 ; n18428_not
g88473 not n18860 ; n18860_not
g88474 not n45347 ; n45347_not
g88475 not n54293 ; n54293_not
g88476 not n54275 ; n54275_not
g88477 not n18905 ; n18905_not
g88478 not n54266 ; n54266_not
g88479 not n18914 ; n18914_not
g88480 not n41945 ; n41945_not
g88481 not n18923 ; n18923_not
g88482 not n54428 ; n54428_not
g88483 not n18680 ; n18680_not
g88484 not n54419 ; n54419_not
g88485 not n18518 ; n18518_not
g88486 not n18707 ; n18707_not
g88487 not n18716 ; n18716_not
g88488 not n54365 ; n54365_not
g88489 not n18725 ; n18725_not
g88490 not n18734 ; n18734_not
g88491 not n54374 ; n54374_not
g88492 not n45338 ; n45338_not
g88493 not n18743 ; n18743_not
g88494 not n54383 ; n54383_not
g88495 not n53546 ; n53546_not
g88496 not n18752 ; n18752_not
g88497 not n18761 ; n18761_not
g88498 not n18770 ; n18770_not
g88499 not n17780 ; n17780_not
g88500 not n17375 ; n17375_not
g88501 not n54662 ; n54662_not
g88502 not n17384 ; n17384_not
g88503 not n17393 ; n17393_not
g88504 not n54653 ; n54653_not
g88505 not n54644 ; n54644_not
g88506 not n17753 ; n17753_not
g88507 not n54239 ; n54239_not
g88508 not n17429 ; n17429_not
g88509 not n17744 ; n17744_not
g88510 not n17438 ; n17438_not
g88511 not n54635 ; n54635_not
g88512 not n41873 ; n41873_not
g88513 not n45293 ; n45293_not
g88514 not n17447 ; n17447_not
g88515 not n17735 ; n17735_not
g88516 not n17456 ; n17456_not
g88517 not n17465 ; n17465_not
g88518 not n54626 ; n54626_not
g88519 not n17285 ; n17285_not
g88520 not n17825 ; n17825_not
g88521 not n54185 ; n54185_not
g88522 not n41837 ; n41837_not
g88523 not n54725 ; n54725_not
g88524 not n17294 ; n17294_not
g88525 not n54194 ; n54194_not
g88526 not n54716 ; n54716_not
g88527 not n41846 ; n41846_not
g88528 not n54707 ; n54707_not
g88529 not n17339 ; n17339_not
g88530 not n17348 ; n17348_not
g88531 not n54680 ; n54680_not
g88532 not n17357 ; n17357_not
g88533 not n45284 ; n45284_not
g88534 not n54671 ; n54671_not
g88535 not n17366 ; n17366_not
g88536 not n17663 ; n17663_not
g88537 not n17591 ; n17591_not
g88538 not n17654 ; n17654_not
g88539 not n54563 ; n54563_not
g88540 not n17609 ; n17609_not
g88541 not n17645 ; n17645_not
g88542 not n54284 ; n54284_not
g88543 not n54554 ; n54554_not
g88544 not n41918 ; n41918_not
g88545 not n17627 ; n17627_not
g88546 not n54545 ; n54545_not
g88547 not n18329 ; n18329_not
g88548 not n18347 ; n18347_not
g88549 not n41927 ; n41927_not
g88550 not n18365 ; n18365_not
g88551 not n18374 ; n18374_not
g88552 not n41936 ; n41936_not
g88553 not n54536 ; n54536_not
g88554 not n18392 ; n18392_not
g88555 not n17474 ; n17474_not
g88556 not n17483 ; n17483_not
g88557 not n41882 ; n41882_not
g88558 not n17492 ; n17492_not
g88559 not n54617 ; n54617_not
g88560 not n17708 ; n17708_not
g88561 not n41891 ; n41891_not
g88562 not n54608 ; n54608_not
g88563 not n17519 ; n17519_not
g88564 not n17528 ; n17528_not
g88565 not n17690 ; n17690_not
g88566 not n17537 ; n17537_not
g88567 not n54590 ; n54590_not
g88568 not n17546 ; n17546_not
g88569 not n17555 ; n17555_not
g88570 not n54581 ; n54581_not
g88571 not n17564 ; n17564_not
g88572 not n17573 ; n17573_not
g88573 not n54572 ; n54572_not
g88574 not n17582 ; n17582_not
g88575 not n53456 ; n53456_not
g88576 not n19940 ; n19940_not
g88577 not n41378 ; n41378_not
g88578 not n53465 ; n53465_not
g88579 not n53474 ; n53474_not
g88580 not n41387 ; n41387_not
g88581 not n41396 ; n41396_not
g88582 not n45428 ; n45428_not
g88583 not n53519 ; n53519_not
g88584 not n19913 ; n19913_not
g88585 not n19076 ; n19076_not
g88586 not n19067 ; n19067_not
g88587 not n53375 ; n53375_not
g88588 not n19058 ; n19058_not
g88589 not n53384 ; n53384_not
g88590 not n19751 ; n19751_not
g88591 not n19805 ; n19805_not
g88592 not n19814 ; n19814_not
g88593 not n19832 ; n19832_not
g88594 not n19850 ; n19850_not
g88595 not n53429 ; n53429_not
g88596 not n19904 ; n19904_not
g88597 not n19922 ; n19922_not
g88598 not n45419 ; n45419_not
g88599 not n45446 ; n45446_not
g88600 not n53438 ; n53438_not
g88601 not n20849 ; n20849_not
g88602 not n20858 ; n20858_not
g88603 not n20867 ; n20867_not
g88604 not n20876 ; n20876_not
g88605 not n20885 ; n20885_not
g88606 not n20894 ; n20894_not
g88607 not n20678 ; n20678_not
g88608 not n20939 ; n20939_not
g88609 not n20669 ; n20669_not
g88610 not n20948 ; n20948_not
g88611 not n20957 ; n20957_not
g88612 not n20966 ; n20966_not
g88613 not n20975 ; n20975_not
g88614 not n20984 ; n20984_not
g88615 not n20993 ; n20993_not
g88616 not n41297 ; n41297_not
g88617 not n53393 ; n53393_not
g88618 not n41288 ; n41288_not
g88619 not n20588 ; n20588_not
g88620 not n53366 ; n53366_not
g88621 not n20579 ; n20579_not
g88622 not n53528 ; n53528_not
g88623 not n19823 ; n19823_not
g88624 not n20399 ; n20399_not
g88625 not n45437 ; n45437_not
g88626 not n53483 ; n53483_not
g88627 not n20489 ; n20489_not
g88628 not n20597 ; n20597_not
g88629 not n20687 ; n20687_not
g88630 not n20759 ; n20759_not
g88631 not n19148 ; n19148_not
g88632 not n19157 ; n19157_not
g88633 not n45365 ; n45365_not
g88634 not n41855 ; n41855_not
g88635 not n19175 ; n19175_not
g88636 not n54095 ; n54095_not
g88637 not n19193 ; n19193_not
g88638 not n54086 ; n54086_not
g88639 not n18932 ; n18932_not
g88640 not n54248 ; n54248_not
g88641 not n18383 ; n18383_not
g88642 not n18941 ; n18941_not
g88643 not n18950 ; n18950_not
g88644 not n54176 ; n54176_not
g88645 not n18338 ; n18338_not
g88646 not n45356 ; n45356_not
g88647 not n19049 ; n19049_not
g88648 not n19085 ; n19085_not
g88649 not n54158 ; n54158_not
g88650 not n45185 ; n45185_not
g88651 not n19247 ; n19247_not
g88652 not n19238 ; n19238_not
g88653 not n45383 ; n45383_not
g88654 not n53294 ; n53294_not
g88655 not n19166 ; n19166_not
g88656 not n45167 ; n45167_not
g88657 not n45392 ; n45392_not
g88658 not n53339 ; n53339_not
g88659 not n54077 ; n54077_not
g88660 not n41828 ; n41828_not
g88661 not n19265 ; n19265_not
g88662 not n19283 ; n19283_not
g88663 not n19292 ; n19292_not
g88664 not n45176 ; n45176_not
g88665 not n45374 ; n45374_not
g88666 not n19256 ; n19256_not
g88667 not n42485 ; n42485_not
g88668 not n16673 ; n16673_not
g88669 not n16682 ; n16682_not
g88670 not n42494 ; n42494_not
g88671 not n16691 ; n16691_not
g88672 not n16709 ; n16709_not
g88673 not n16718 ; n16718_not
g88674 not n16394 ; n16394_not
g88675 not n16727 ; n16727_not
g88676 not n16736 ; n16736_not
g88677 not n16385 ; n16385_not
g88678 not n16745 ; n16745_not
g88679 not n16754 ; n16754_not
g88680 not n16088 ; n16088_not
g88681 not n16763 ; n16763_not
g88682 not n16097 ; n16097_not
g88683 not n16475 ; n16475_not
g88684 not n16583 ; n16583_not
g88685 not n16592 ; n16592_not
g88686 not n16619 ; n16619_not
g88687 not n16628 ; n16628_not
g88688 not n16448 ; n16448_not
g88689 not n42476 ; n42476_not
g88690 not n16637 ; n16637_not
g88691 not n16439 ; n16439_not
g88692 not n16646 ; n16646_not
g88693 not n16655 ; n16655_not
g88694 not n16664 ; n16664_not
g88695 not n16196 ; n16196_not
g88696 not n16871 ; n16871_not
g88697 not n42539 ; n42539_not
g88698 not n16880 ; n16880_not
g88699 not n16295 ; n16295_not
g88700 not n16907 ; n16907_not
g88701 not n16916 ; n16916_not
g88702 not n16268 ; n16268_not
g88703 not n16925 ; n16925_not
g88704 not n16259 ; n16259_not
g88705 not n16934 ; n16934_not
g88706 not n16943 ; n16943_not
g88707 not n55157 ; n55157_not
g88708 not n16952 ; n16952_not
g88709 not n16961 ; n16961_not
g88710 not n16772 ; n16772_not
g88711 not n16781 ; n16781_not
g88712 not n16790 ; n16790_not
g88713 not n16358 ; n16358_not
g88714 not n16349 ; n16349_not
g88715 not n16808 ; n16808_not
g88716 not n16817 ; n16817_not
g88717 not n45194 ; n45194_not
g88718 not n16826 ; n16826_not
g88719 not n16835 ; n16835_not
g88720 not n16169 ; n16169_not
g88721 not n16844 ; n16844_not
g88722 not n16178 ; n16178_not
g88723 not n16853 ; n16853_not
g88724 not n16187 ; n16187_not
g88725 not n16862 ; n16862_not
g88726 not n15665 ; n15665_not
g88727 not n55193 ; n55193_not
g88728 not n16484 ; n16484_not
g88729 not n42449 ; n42449_not
g88730 not n16538 ; n16538_not
g88731 not n16547 ; n16547_not
g88732 not n16493 ; n16493_not
g88733 not n16556 ; n16556_not
g88734 not n16565 ; n16565_not
g88735 not n16574 ; n16574_not
g88736 not n45149 ; n45149_not
g88737 not n43079 ; n43079_not
g88738 not n16367 ; n16367_not
g88739 not n16457 ; n16457_not
g88740 not n17762 ; n17762_not
g88741 not n54833 ; n54833_not
g88742 not n17672 ; n17672_not
g88743 not n54851 ; n54851_not
g88744 not n54842 ; n54842_not
g88745 not n17717 ; n17717_not
g88746 not n17852 ; n17852_not
g88747 not n54806 ; n54806_not
g88748 not n54149 ; n54149_not
g88749 not n54770 ; n54770_not
g88750 not n54761 ; n54761_not
g88751 not n17249 ; n17249_not
g88752 not n54752 ; n54752_not
g88753 not n17258 ; n17258_not
g88754 not n17843 ; n17843_not
g88755 not n54743 ; n54743_not
g88756 not n17267 ; n17267_not
g88757 not n17834 ; n17834_not
g88758 not n17276 ; n17276_not
g88759 not n54734 ; n54734_not
g88760 not n42458 ; n42458_not
g88761 not n54824 ; n54824_not
g88762 not n17807 ; n17807_not
g88763 not n45275 ; n45275_not
g88764 not n54815 ; n54815_not
g88765 not n17159 ; n17159_not
g88766 not n17168 ; n17168_not
g88767 not n17186 ; n17186_not
g88768 not n45239 ; n45239_not
g88769 not n55067 ; n55067_not
g88770 not n17177 ; n17177_not
g88771 not n17087 ; n17087_not
g88772 not n42629 ; n42629_not
g88773 not n17078 ; n17078_not
g88774 not n45257 ; n45257_not
g88775 not n42566 ; n42566_not
g88776 not n17069 ; n17069_not
g88777 not n17096 ; n17096_not
g88778 not n42575 ; n42575_not
g88779 not n42584 ; n42584_not
g88780 not n42548 ; n42548_not
g88781 not n54860 ; n54860_not
g88782 not n42665 ; n42665_not
g88783 not n42647 ; n42647_not
g88784 not n42656 ; n42656_not
g88785 not n54905 ; n54905_not
g88786 not n54914 ; n54914_not
g88787 not n54932 ; n54932_not
g88788 not n45266 ; n45266_not
g88789 not n42593 ; n42593_not
g88790 not n37094 ; n37094_not
g88791 not n37229 ; n37229_not
g88792 not n34196 ; n34196_not
g88793 not n46634 ; n46634_not
g88794 not n28463 ; n28463_not
g88795 not n37085 ; n37085_not
g88796 not n34088 ; n34088_not
g88797 not n46823 ; n46823_not
g88798 not n34187 ; n34187_not
g88799 not n37238 ; n37238_not
g88800 not n38651 ; n38651_not
g88801 not n34178 ; n34178_not
g88802 not n34097 ; n34097_not
g88803 not n34169 ; n34169_not
g88804 not n37247 ; n37247_not
g88805 not n48074 ; n48074_not
g88806 not n37076 ; n37076_not
g88807 not n37256 ; n37256_not
g88808 not n34448 ; n34448_not
g88809 not n46814 ; n46814_not
g88810 not n34385 ; n34385_not
g88811 not n46517 ; n46517_not
g88812 not n28445 ; n28445_not
g88813 not n48047 ; n48047_not
g88814 not n38525 ; n38525_not
g88815 not n28454 ; n28454_not
g88816 not n34358 ; n34358_not
g88817 not n34349 ; n34349_not
g88818 not n34295 ; n34295_not
g88819 not n34286 ; n34286_not
g88820 not n34277 ; n34277_not
g88821 not n34268 ; n34268_not
g88822 not n34259 ; n34259_not
g88823 not n37049 ; n37049_not
g88824 not n33656 ; n33656_not
g88825 not n46508 ; n46508_not
g88826 not n33665 ; n33665_not
g88827 not n50198 ; n50198_not
g88828 not n27860 ; n27860_not
g88829 not n37319 ; n37319_not
g88830 not n48029 ; n48029_not
g88831 not n33692 ; n33692_not
g88832 not n28508 ; n28508_not
g88833 not n46841 ; n46841_not
g88834 not n37328 ; n37328_not
g88835 not n50288 ; n50288_not
g88836 not n37337 ; n37337_not
g88837 not n33764 ; n33764_not
g88838 not n28517 ; n28517_not
g88839 not n28472 ; n28472_not
g88840 not n48065 ; n48065_not
g88841 not n37265 ; n37265_not
g88842 not n37274 ; n37274_not
g88843 not n48056 ; n48056_not
g88844 not n37283 ; n37283_not
g88845 not n37292 ; n37292_not
g88846 not n38534 ; n38534_not
g88847 not n27851 ; n27851_not
g88848 not n46832 ; n46832_not
g88849 not n38543 ; n38543_not
g88850 not n28481 ; n28481_not
g88851 not n48038 ; n48038_not
g88852 not n28490 ; n28490_not
g88853 not n33647 ; n33647_not
g88854 not n34646 ; n34646_not
g88855 not n37157 ; n37157_not
g88856 not n28346 ; n28346_not
g88857 not n34439 ; n34439_not
g88858 not n49334 ; n49334_not
g88859 not n51629 ; n51629_not
g88860 not n34637 ; n34637_not
g88861 not n28355 ; n28355_not
g88862 not n28364 ; n28364_not
g88863 not n34628 ; n34628_not
g88864 not n34619 ; n34619_not
g88865 not n28373 ; n28373_not
g88866 not n37166 ; n37166_not
g88867 not n49325 ; n49325_not
g88868 not n37139 ; n37139_not
g88869 not n34682 ; n34682_not
g88870 not n46751 ; n46751_not
g88871 not n34673 ; n34673_not
g88872 not n46553 ; n46553_not
g88873 not n37148 ; n37148_not
g88874 not n27815 ; n27815_not
g88875 not n28319 ; n28319_not
g88876 not n34664 ; n34664_not
g88877 not n49343 ; n49343_not
g88878 not n46760 ; n46760_not
g88879 not n27806 ; n27806_not
g88880 not n34655 ; n34655_not
g88881 not n37184 ; n37184_not
g88882 not n34547 ; n34547_not
g88883 not n46805 ; n46805_not
g88884 not n34538 ; n34538_not
g88885 not n27824 ; n27824_not
g88886 not n28427 ; n28427_not
g88887 not n46526 ; n46526_not
g88888 not n34529 ; n34529_not
g88889 not n50837 ; n50837_not
g88890 not n34493 ; n34493_not
g88891 not n28436 ; n28436_not
g88892 not n37193 ; n37193_not
g88893 not n34475 ; n34475_not
g88894 not n34466 ; n34466_not
g88895 not n28382 ; n28382_not
g88896 not n34592 ; n34592_not
g88897 not n34583 ; n34583_not
g88898 not n37175 ; n37175_not
g88899 not n34574 ; n34574_not
g88900 not n28391 ; n28391_not
g88901 not n34565 ; n34565_not
g88902 not n34484 ; n34484_not
g88903 not n34556 ; n34556_not
g88904 not n50828 ; n50828_not
g88905 not n28328 ; n28328_not
g88906 not n28409 ; n28409_not
g88907 not n28418 ; n28418_not
g88908 not n32918 ; n32918_not
g88909 not n32909 ; n32909_not
g88910 not n50873 ; n50873_not
g88911 not n37409 ; n37409_not
g88912 not n32891 ; n32891_not
g88913 not n27914 ; n27914_not
g88914 not n50369 ; n50369_not
g88915 not n32882 ; n32882_not
g88916 not n46922 ; n46922_not
g88917 not n47903 ; n47903_not
g88918 not n32954 ; n32954_not
g88919 not n37391 ; n37391_not
g88920 not n37481 ; n37481_not
g88921 not n50882 ; n50882_not
g88922 not n37382 ; n37382_not
g88923 not n32873 ; n32873_not
g88924 not n37373 ; n37373_not
g88925 not n37445 ; n37445_not
g88926 not n33188 ; n33188_not
g88927 not n33197 ; n33197_not
g88928 not n28571 ; n28571_not
g88929 not n46913 ; n46913_not
g88930 not n33287 ; n33287_not
g88931 not n37436 ; n37436_not
g88932 not n37454 ; n37454_not
g88933 not n37427 ; n37427_not
g88934 not n33269 ; n33269_not
g88935 not n28580 ; n28580_not
g88936 not n32927 ; n32927_not
g88937 not n46463 ; n46463_not
g88938 not n37463 ; n37463_not
g88939 not n37418 ; n37418_not
g88940 not n32819 ; n32819_not
g88941 not n50387 ; n50387_not
g88942 not n32792 ; n32792_not
g88943 not n37526 ; n37526_not
g88944 not n32783 ; n32783_not
g88945 not n32774 ; n32774_not
g88946 not n32765 ; n32765_not
g88947 not n28625 ; n28625_not
g88948 not n32756 ; n32756_not
g88949 not n28634 ; n28634_not
g88950 not n47831 ; n47831_not
g88951 not n46940 ; n46940_not
g88952 not n32747 ; n32747_not
g88953 not n32864 ; n32864_not
g88954 not n37364 ; n37364_not
g88955 not n32963 ; n32963_not
g88956 not n28607 ; n28607_not
g88957 not n37355 ; n37355_not
g88958 not n32855 ; n32855_not
g88959 not n32972 ; n32972_not
g88960 not n50297 ; n50297_not
g88961 not n37346 ; n37346_not
g88962 not n32846 ; n32846_not
g88963 not n28616 ; n28616_not
g88964 not n37508 ; n37508_not
g88965 not n32837 ; n32837_not
g88966 not n50378 ; n50378_not
g88967 not n46931 ; n46931_not
g88968 not n32828 ; n32828_not
g88969 not n33629 ; n33629_not
g88970 not n33593 ; n33593_not
g88971 not n33584 ; n33584_not
g88972 not n33278 ; n33278_not
g88973 not n33575 ; n33575_not
g88974 not n33566 ; n33566_not
g88975 not n33557 ; n33557_not
g88976 not n33548 ; n33548_not
g88977 not n33539 ; n33539_not
g88978 not n33179 ; n33179_not
g88979 not n33737 ; n33737_not
g88980 not n28526 ; n28526_not
g88981 not n33755 ; n33755_not
g88982 not n46850 ; n46850_not
g88983 not n33719 ; n33719_not
g88984 not n28535 ; n28535_not
g88985 not n28544 ; n28544_not
g88986 not n33674 ; n33674_not
g88987 not n33395 ; n33395_not
g88988 not n33377 ; n33377_not
g88989 not n46904 ; n46904_not
g88990 not n33089 ; n33089_not
g88991 not n28562 ; n28562_not
g88992 not n47921 ; n47921_not
g88993 not n33098 ; n33098_not
g88994 not n33359 ; n33359_not
g88995 not n28256 ; n28256_not
g88996 not n33494 ; n33494_not
g88997 not n33485 ; n33485_not
g88998 not n46481 ; n46481_not
g88999 not n33476 ; n33476_not
g89000 not n38570 ; n38570_not
g89001 not n33467 ; n33467_not
g89002 not n33458 ; n33458_not
g89003 not n33449 ; n33449_not
g89004 not n50864 ; n50864_not
g89005 not n46472 ; n46472_not
g89006 not n33368 ; n33368_not
g89007 not n28553 ; n28553_not
g89008 not n27770 ; n27770_not
g89009 not n35186 ; n35186_not
g89010 not n51845 ; n51845_not
g89011 not n46067 ; n46067_not
g89012 not n34763 ; n34763_not
g89013 not n46058 ; n46058_not
g89014 not n39155 ; n39155_not
g89015 not n27833 ; n27833_not
g89016 not n49415 ; n49415_not
g89017 not n46049 ; n46049_not
g89018 not n35168 ; n35168_not
g89019 not n49424 ; n49424_not
g89020 not n39191 ; n39191_not
g89021 not n27743 ; n27743_not
g89022 not n38714 ; n38714_not
g89023 not n46094 ; n46094_not
g89024 not n27752 ; n27752_not
g89025 not n35285 ; n35285_not
g89026 not n27761 ; n27761_not
g89027 not n36554 ; n36554_not
g89028 not n46085 ; n46085_not
g89029 not n38705 ; n38705_not
g89030 not n46535 ; n46535_not
g89031 not n26915 ; n26915_not
g89032 not n35267 ; n35267_not
g89033 not n35258 ; n35258_not
g89034 not n35195 ; n35195_not
g89035 not n51872 ; n51872_not
g89036 not n51863 ; n51863_not
g89037 not n46076 ; n46076_not
g89038 not n35096 ; n35096_not
g89039 not n38660 ; n38660_not
g89040 not n46580 ; n46580_not
g89041 not n49460 ; n49460_not
g89042 not n35087 ; n35087_not
g89043 not n35078 ; n35078_not
g89044 not n36527 ; n36527_not
g89045 not n35069 ; n35069_not
g89046 not n27923 ; n27923_not
g89047 not n46607 ; n46607_not
g89048 not n49505 ; n49505_not
g89049 not n36518 ; n36518_not
g89050 not n45950 ; n45950_not
g89051 not n49514 ; n49514_not
g89052 not n35159 ; n35159_not
g89053 not n39173 ; n39173_not
g89054 not n39164 ; n39164_not
g89055 not n51827 ; n51827_not
g89056 not n46562 ; n46562_not
g89057 not n39182 ; n39182_not
g89058 not n51818 ; n51818_not
g89059 not n49442 ; n49442_not
g89060 not n34790 ; n34790_not
g89061 not n34808 ; n34808_not
g89062 not n27905 ; n27905_not
g89063 not n46490 ; n46490_not
g89064 not n35339 ; n35339_not
g89065 not n35375 ; n35375_not
g89066 not n46157 ; n46157_not
g89067 not n27635 ; n27635_not
g89068 not n46148 ; n46148_not
g89069 not n35366 ; n35366_not
g89070 not n46139 ; n46139_not
g89071 not n27644 ; n27644_not
g89072 not n49352 ; n49352_not
g89073 not n35357 ; n35357_not
g89074 not n27608 ; n27608_not
g89075 not n46193 ; n46193_not
g89076 not n46184 ; n46184_not
g89077 not n27617 ; n27617_not
g89078 not n35393 ; n35393_not
g89079 not n46175 ; n46175_not
g89080 not n35384 ; n35384_not
g89081 not n46166 ; n46166_not
g89082 not n27626 ; n27626_not
g89083 not n26960 ; n26960_not
g89084 not n51908 ; n51908_not
g89085 not n26951 ; n26951_not
g89086 not n27707 ; n27707_not
g89087 not n39128 ; n39128_not
g89088 not n38732 ; n38732_not
g89089 not n34925 ; n34925_not
g89090 not n27716 ; n27716_not
g89091 not n26942 ; n26942_not
g89092 not n27725 ; n27725_not
g89093 not n27734 ; n27734_not
g89094 not n49370 ; n49370_not
g89095 not n38723 ; n38723_not
g89096 not n47912 ; n47912_not
g89097 not n51890 ; n51890_not
g89098 not n27653 ; n27653_not
g89099 not n35348 ; n35348_not
g89100 not n36572 ; n36572_not
g89101 not n27662 ; n27662_not
g89102 not n27671 ; n27671_not
g89103 not n38750 ; n38750_not
g89104 not n36563 ; n36563_not
g89105 not n27680 ; n27680_not
g89106 not n39119 ; n39119_not
g89107 not n38741 ; n38741_not
g89108 not n51917 ; n51917_not
g89109 not n28157 ; n28157_not
g89110 not n38921 ; n38921_not
g89111 not n38930 ; n38930_not
g89112 not n34844 ; n34844_not
g89113 not n28175 ; n28175_not
g89114 not n34835 ; n34835_not
g89115 not n34817 ; n34817_not
g89116 not n51692 ; n51692_not
g89117 not n46661 ; n46661_not
g89118 not n28076 ; n28076_not
g89119 not n49433 ; n49433_not
g89120 not n34862 ; n34862_not
g89121 not n28049 ; n28049_not
g89122 not n39029 ; n39029_not
g89123 not n38903 ; n38903_not
g89124 not n46670 ; n46670_not
g89125 not n28139 ; n28139_not
g89126 not n38912 ; n38912_not
g89127 not n28148 ; n28148_not
g89128 not n46733 ; n46733_not
g89129 not n51665 ; n51665_not
g89130 not n34727 ; n34727_not
g89131 not n34394 ; n34394_not
g89132 not n34718 ; n34718_not
g89133 not n28283 ; n28283_not
g89134 not n46742 ; n46742_not
g89135 not n34709 ; n34709_not
g89136 not n34691 ; n34691_not
g89137 not n38480 ; n38480_not
g89138 not n28292 ; n28292_not
g89139 not n46706 ; n46706_not
g89140 not n34772 ; n34772_not
g89141 not n28229 ; n28229_not
g89142 not n51683 ; n51683_not
g89143 not n46715 ; n46715_not
g89144 not n34754 ; n34754_not
g89145 not n28247 ; n28247_not
g89146 not n46724 ; n46724_not
g89147 not n34745 ; n34745_not
g89148 not n46571 ; n46571_not
g89149 not n34736 ; n34736_not
g89150 not n28274 ; n28274_not
g89151 not n27950 ; n27950_not
g89152 not n49550 ; n49550_not
g89153 not n45941 ; n45941_not
g89154 not n51755 ; n51755_not
g89155 not n49523 ; n49523_not
g89156 not n46625 ; n46625_not
g89157 not n39092 ; n39092_not
g89158 not n51782 ; n51782_not
g89159 not n39137 ; n39137_not
g89160 not n49532 ; n49532_not
g89161 not n27941 ; n27941_not
g89162 not n51773 ; n51773_not
g89163 not n34853 ; n34853_not
g89164 not n48821 ; n48821_not
g89165 not n34952 ; n34952_not
g89166 not n38831 ; n38831_not
g89167 not n39065 ; n39065_not
g89168 not n38840 ; n38840_not
g89169 not n34943 ; n34943_not
g89170 not n34934 ; n34934_not
g89171 not n51728 ; n51728_not
g89172 not n37058 ; n37058_not
g89173 not n28085 ; n28085_not
g89174 not n39047 ; n39047_not
g89175 not n34880 ; n34880_not
g89176 not n51737 ; n51737_not
g89177 not n46616 ; n46616_not
g89178 not n38804 ; n38804_not
g89179 not n34970 ; n34970_not
g89180 not n38813 ; n38813_not
g89181 not n34961 ; n34961_not
g89182 not n39074 ; n39074_not
g89183 not n38822 ; n38822_not
g89184 not n28058 ; n28058_not
g89185 not n46643 ; n46643_not
g89186 not n29714 ; n29714_not
g89187 not n29705 ; n29705_not
g89188 not n47444 ; n47444_not
g89189 not n37634 ; n37634_not
g89190 not n31676 ; n31676_not
g89191 not n31685 ; n31685_not
g89192 not n29660 ; n29660_not
g89193 not n37940 ; n37940_not
g89194 not n29651 ; n29651_not
g89195 not n50981 ; n50981_not
g89196 not n47291 ; n47291_not
g89197 not n38039 ; n38039_not
g89198 not n31397 ; n31397_not
g89199 not n31784 ; n31784_not
g89200 not n47462 ; n47462_not
g89201 not n31766 ; n31766_not
g89202 not n29732 ; n29732_not
g89203 not n37922 ; n37922_not
g89204 not n31748 ; n31748_not
g89205 not n47453 ; n47453_not
g89206 not n29741 ; n29741_not
g89207 not n31739 ; n31739_not
g89208 not n47282 ; n47282_not
g89209 not n37931 ; n37931_not
g89210 not n47138 ; n47138_not
g89211 not n29723 ; n29723_not
g89212 not n31694 ; n31694_not
g89213 not n31289 ; n31289_not
g89214 not n50918 ; n50918_not
g89215 not n47165 ; n47165_not
g89216 not n31496 ; n31496_not
g89217 not n37913 ; n37913_not
g89218 not n47390 ; n47390_not
g89219 not n31478 ; n31478_not
g89220 not n50909 ; n50909_not
g89221 not n47318 ; n47318_not
g89222 not n37904 ; n37904_not
g89223 not n47381 ; n47381_not
g89224 not n29750 ; n29750_not
g89225 not n47372 ; n47372_not
g89226 not n47435 ; n47435_not
g89227 not n29804 ; n29804_not
g89228 not n31388 ; n31388_not
g89229 not n50963 ; n50963_not
g89230 not n31379 ; n31379_not
g89231 not n47426 ; n47426_not
g89232 not n29813 ; n29813_not
g89233 not n50954 ; n50954_not
g89234 not n31469 ; n31469_not
g89235 not n47417 ; n47417_not
g89236 not n47147 ; n47147_not
g89237 not n50936 ; n50936_not
g89238 not n47408 ; n47408_not
g89239 not n31298 ; n31298_not
g89240 not n29507 ; n29507_not
g89241 not n29516 ; n29516_not
g89242 not n29408 ; n29408_not
g89243 not n47237 ; n47237_not
g89244 not n31793 ; n31793_not
g89245 not n47525 ; n47525_not
g89246 not n47246 ; n47246_not
g89247 not n50585 ; n50585_not
g89248 not n47516 ; n47516_not
g89249 not n47075 ; n47075_not
g89250 not n51098 ; n51098_not
g89251 not n47066 ; n47066_not
g89252 not n47507 ; n47507_not
g89253 not n29390 ; n29390_not
g89254 not n29471 ; n29471_not
g89255 not n37841 ; n37841_not
g89256 not n47228 ; n47228_not
g89257 not n50576 ; n50576_not
g89258 not n47543 ; n47543_not
g89259 not n29453 ; n29453_not
g89260 not n37850 ; n37850_not
g89261 not n29444 ; n29444_not
g89262 not n29435 ; n29435_not
g89263 not n51089 ; n51089_not
g89264 not n29426 ; n29426_not
g89265 not n29417 ; n29417_not
g89266 not n47534 ; n47534_not
g89267 not n50594 ; n50594_not
g89268 not n47273 ; n47273_not
g89269 not n29633 ; n29633_not
g89270 not n37472 ; n37472_not
g89271 not n29624 ; n29624_not
g89272 not n29615 ; n29615_not
g89273 not n47057 ; n47057_not
g89274 not n29462 ; n29462_not
g89275 not n31757 ; n31757_not
g89276 not n47048 ; n47048_not
g89277 not n47039 ; n47039_not
g89278 not n47480 ; n47480_not
g89279 not n29642 ; n29642_not
g89280 not n47471 ; n47471_not
g89281 not n30497 ; n30497_not
g89282 not n30956 ; n30956_not
g89283 not n38075 ; n38075_not
g89284 not n37742 ; n37742_not
g89285 not n30488 ; n30488_not
g89286 not n30659 ; n30659_not
g89287 not n30839 ; n30839_not
g89288 not n30668 ; n30668_not
g89289 not n30677 ; n30677_not
g89290 not n37733 ; n37733_not
g89291 not n30848 ; n30848_not
g89292 not n30686 ; n30686_not
g89293 not n50693 ; n50693_not
g89294 not n30857 ; n30857_not
g89295 not n30695 ; n30695_not
g89296 not n30938 ; n30938_not
g89297 not n30776 ; n30776_not
g89298 not n30983 ; n30983_not
g89299 not n30785 ; n30785_not
g89300 not n37760 ; n37760_not
g89301 not n50738 ; n50738_not
g89302 not n30569 ; n30569_not
g89303 not n30578 ; n30578_not
g89304 not n50684 ; n50684_not
g89305 not n30974 ; n30974_not
g89306 not n38066 ; n38066_not
g89307 not n30587 ; n30587_not
g89308 not n30794 ; n30794_not
g89309 not n30596 ; n30596_not
g89310 not n37751 ; n37751_not
g89311 not n37706 ; n37706_not
g89312 not n30884 ; n30884_not
g89313 not n30893 ; n30893_not
g89314 not n30866 ; n30866_not
g89315 not n37661 ; n37661_not
g89316 not n30875 ; n30875_not
g89317 not n37670 ; n37670_not
g89318 not n30758 ; n30758_not
g89319 not n30767 ; n30767_not
g89320 not n37724 ; n37724_not
g89321 not n50729 ; n50729_not
g89322 not n47255 ; n47255_not
g89323 not n37652 ; n37652_not
g89324 not n38138 ; n38138_not
g89325 not n30929 ; n30929_not
g89326 not n38129 ; n38129_not
g89327 not n37715 ; n37715_not
g89328 not n38093 ; n38093_not
g89329 not n31199 ; n31199_not
g89330 not n47345 ; n47345_not
g89331 not n29930 ; n29930_not
g89332 not n37832 ; n37832_not
g89333 not n50846 ; n50846_not
g89334 not n30947 ; n30947_not
g89335 not n38084 ; n38084_not
g89336 not n29840 ; n29840_not
g89337 not n37823 ; n37823_not
g89338 not n50819 ; n50819_not
g89339 not n50891 ; n50891_not
g89340 not n47327 ; n47327_not
g89341 not n47363 ; n47363_not
g89342 not n29903 ; n29903_not
g89343 not n47336 ; n47336_not
g89344 not n47183 ; n47183_not
g89345 not n47354 ; n47354_not
g89346 not n50639 ; n50639_not
g89347 not n29912 ; n29912_not
g89348 not n47192 ; n47192_not
g89349 not n50666 ; n50666_not
g89350 not n38048 ; n38048_not
g89351 not n50765 ; n50765_not
g89352 not n50756 ; n50756_not
g89353 not n50747 ; n50747_not
g89354 not n50675 ; n50675_not
g89355 not n30299 ; n30299_not
g89356 not n30992 ; n30992_not
g89357 not n30389 ; n30389_not
g89358 not n30398 ; n30398_not
g89359 not n29831 ; n29831_not
g89360 not n50648 ; n50648_not
g89361 not n29822 ; n29822_not
g89362 not n37814 ; n37814_not
g89363 not n50792 ; n50792_not
g89364 not n50783 ; n50783_not
g89365 not n37805 ; n37805_not
g89366 not n50657 ; n50657_not
g89367 not n50774 ; n50774_not
g89368 not n29921 ; n29921_not
g89369 not n28733 ; n28733_not
g89370 not n50927 ; n50927_not
g89371 not n28742 ; n28742_not
g89372 not n47723 ; n47723_not
g89373 not n32684 ; n32684_not
g89374 not n32675 ; n32675_not
g89375 not n32657 ; n32657_not
g89376 not n32639 ; n32639_not
g89377 not n50477 ; n50477_not
g89378 not n47714 ; n47714_not
g89379 not n28751 ; n28751_not
g89380 not n32594 ; n32594_not
g89381 not n28760 ; n28760_not
g89382 not n28724 ; n28724_not
g89383 not n50459 ; n50459_not
g89384 not n37607 ; n37607_not
g89385 not n47732 ; n47732_not
g89386 not n32738 ; n32738_not
g89387 not n28184 ; n28184_not
g89388 not n46418 ; n46418_not
g89389 not n32693 ; n32693_not
g89390 not n50468 ; n50468_not
g89391 not n28823 ; n28823_not
g89392 not n28832 ; n28832_not
g89393 not n50495 ; n50495_not
g89394 not n47156 ; n47156_not
g89395 not n32369 ; n32369_not
g89396 not n32378 ; n32378_not
g89397 not n32396 ; n32396_not
g89398 not n38624 ; n38624_not
g89399 not n28841 ; n28841_not
g89400 not n32387 ; n32387_not
g89401 not n38615 ; n38615_not
g89402 not n28850 ; n28850_not
g89403 not n32279 ; n32279_not
g89404 not n47705 ; n47705_not
g89405 not n32567 ; n32567_not
g89406 not n32288 ; n32288_not
g89407 not n32558 ; n32558_not
g89408 not n32549 ; n32549_not
g89409 not n38642 ; n38642_not
g89410 not n50486 ; n50486_not
g89411 not n28805 ; n28805_not
g89412 not n32495 ; n32495_not
g89413 not n28814 ; n28814_not
g89414 not n32486 ; n32486_not
g89415 not n32477 ; n32477_not
g89416 not n32468 ; n32468_not
g89417 not n32459 ; n32459_not
g89418 not n28661 ; n28661_not
g89419 not n28670 ; n28670_not
g89420 not n32936 ; n32936_not
g89421 not n37616 ; n37616_not
g89422 not n37544 ; n37544_not
g89423 not n32729 ; n32729_not
g89424 not n28643 ; n28643_not
g89425 not n37553 ; n37553_not
g89426 not n47813 ; n47813_not
g89427 not n37571 ; n37571_not
g89428 not n28652 ; n28652_not
g89429 not n50396 ; n50396_not
g89430 not n32981 ; n32981_not
g89431 not n47750 ; n47750_not
g89432 not n32648 ; n32648_not
g89433 not n28715 ; n28715_not
g89434 not n47741 ; n47741_not
g89435 not n38633 ; n38633_not
g89436 not n37625 ; n37625_not
g89437 not n28706 ; n28706_not
g89438 not n46436 ; n46436_not
g89439 not n46427 ; n46427_not
g89440 not n46391 ; n46391_not
g89441 not n29354 ; n29354_not
g89442 not n29309 ; n29309_not
g89443 not n29291 ; n29291_not
g89444 not n29282 ; n29282_not
g89445 not n50567 ; n50567_not
g89446 not n29372 ; n29372_not
g89447 not n29381 ; n29381_not
g89448 not n46382 ; n46382_not
g89449 not n29273 ; n29273_not
g89450 not n29264 ; n29264_not
g89451 not n29255 ; n29255_not
g89452 not n29318 ; n29318_not
g89453 not n29246 ; n29246_not
g89454 not n29327 ; n29327_not
g89455 not n38507 ; n38507_not
g89456 not n29336 ; n29336_not
g89457 not n47570 ; n47570_not
g89458 not n29345 ; n29345_not
g89459 not n47552 ; n47552_not
g89460 not n38462 ; n38462_not
g89461 not n47561 ; n47561_not
g89462 not n29363 ; n29363_not
g89463 not n37517 ; n37517_not
g89464 not n47642 ; n47642_not
g89465 not n32099 ; n32099_not
g89466 not n28940 ; n28940_not
g89467 not n47633 ; n47633_not
g89468 not n47624 ; n47624_not
g89469 not n29048 ; n29048_not
g89470 not n29057 ; n29057_not
g89471 not n29066 ; n29066_not
g89472 not n29075 ; n29075_not
g89473 not n47615 ; n47615_not
g89474 not n29084 ; n29084_not
g89475 not n32297 ; n32297_not
g89476 not n47660 ; n47660_not
g89477 not n31982 ; n31982_not
g89478 not n50972 ; n50972_not
g89479 not n37562 ; n37562_not
g89480 not n47651 ; n47651_not
g89481 not n31991 ; n31991_not
g89482 not n32198 ; n32198_not
g89483 not n28904 ; n28904_not
g89484 not n32189 ; n32189_not
g89485 not n29183 ; n29183_not
g89486 not n50558 ; n50558_not
g89487 not n29192 ; n29192_not
g89488 not n29174 ; n29174_not
g89489 not n31973 ; n31973_not
g89490 not n29165 ; n29165_not
g89491 not n29237 ; n29237_not
g89492 not n29129 ; n29129_not
g89493 not n47606 ; n47606_not
g89494 not n50549 ; n50549_not
g89495 not n29138 ; n29138_not
g89496 not n38552 ; n38552_not
g89497 not n35753 ; n35753_not
g89498 not n46229 ; n46229_not
g89499 not n26861 ; n26861_not
g89500 not n36446 ; n36446_not
g89501 not n26870 ; n26870_not
g89502 not n48461 ; n48461_not
g89503 not n48335 ; n48335_not
g89504 not n36437 ; n36437_not
g89505 not n48470 ; n48470_not
g89506 not n39380 ; n39380_not
g89507 not n26834 ; n26834_not
g89508 not n48452 ; n48452_not
g89509 not n49190 ; n49190_not
g89510 not n26843 ; n26843_not
g89511 not n51746 ; n51746_not
g89512 not n36464 ; n36464_not
g89513 not n48317 ; n48317_not
g89514 not n36536 ; n36536_not
g89515 not n26852 ; n26852_not
g89516 not n36455 ; n36455_not
g89517 not n48326 ; n48326_not
g89518 not n26906 ; n26906_not
g89519 not n48344 ; n48344_not
g89520 not n46256 ; n46256_not
g89521 not n36392 ; n36392_not
g89522 not n48353 ; n48353_not
g89523 not n36383 ; n36383_not
g89524 not n48362 ; n48362_not
g89525 not n36428 ; n36428_not
g89526 not n49208 ; n49208_not
g89527 not n36419 ; n36419_not
g89528 not n46238 ; n46238_not
g89529 not n35762 ; n35762_not
g89530 not n48650 ; n48650_not
g89531 not n46247 ; n46247_not
g89532 not n48263 ; n48263_not
g89533 not n26780 ; n26780_not
g89534 not n39308 ; n39308_not
g89535 not n48425 ; n48425_not
g89536 not n49163 ; n49163_not
g89537 not n39317 ; n39317_not
g89538 not n48434 ; n48434_not
g89539 not n39326 ; n39326_not
g89540 not n39272 ; n39272_not
g89541 not n35717 ; n35717_not
g89542 not n36482 ; n36482_not
g89543 not n48254 ; n48254_not
g89544 not n39281 ; n39281_not
g89545 not n49145 ; n49145_not
g89546 not n48416 ; n48416_not
g89547 not n26771 ; n26771_not
g89548 not n39290 ; n39290_not
g89549 not n35726 ; n35726_not
g89550 not n36491 ; n36491_not
g89551 not n49154 ; n49154_not
g89552 not n39362 ; n39362_not
g89553 not n48281 ; n48281_not
g89554 not n26825 ; n26825_not
g89555 not n39623 ; n39623_not
g89556 not n39371 ; n39371_not
g89557 not n48290 ; n48290_not
g89558 not n48308 ; n48308_not
g89559 not n36473 ; n36473_not
g89560 not n49172 ; n49172_not
g89561 not n48272 ; n48272_not
g89562 not n39335 ; n39335_not
g89563 not n39641 ; n39641_not
g89564 not n39344 ; n39344_not
g89565 not n26807 ; n26807_not
g89566 not n48443 ; n48443_not
g89567 not n39353 ; n39353_not
g89568 not n26816 ; n26816_not
g89569 not n49181 ; n49181_not
g89570 not n35537 ; n35537_not
g89571 not n48506 ; n48506_not
g89572 not n36680 ; n36680_not
g89573 not n48560 ; n48560_not
g89574 not n27077 ; n27077_not
g89575 not n35546 ; n35546_not
g89576 not n48515 ; n48515_not
g89577 not n27086 ; n27086_not
g89578 not n46319 ; n46319_not
g89579 not n49244 ; n49244_not
g89580 not n48524 ; n48524_not
g89581 not n35645 ; n35645_not
g89582 not n36257 ; n36257_not
g89583 not n36653 ; n36653_not
g89584 not n35672 ; n35672_not
g89585 not n36248 ; n36248_not
g89586 not n36239 ; n36239_not
g89587 not n35663 ; n35663_not
g89588 not n35519 ; n35519_not
g89589 not n35528 ; n35528_not
g89590 not n36671 ; n36671_not
g89591 not n27059 ; n27059_not
g89592 not n35609 ; n35609_not
g89593 not n27167 ; n27167_not
g89594 not n36644 ; n36644_not
g89595 not n49253 ; n49253_not
g89596 not n27176 ; n27176_not
g89597 not n46346 ; n46346_not
g89598 not n35591 ; n35591_not
g89599 not n27194 ; n27194_not
g89600 not n46355 ; n46355_not
g89601 not n35555 ; n35555_not
g89602 not n36662 ; n36662_not
g89603 not n35564 ; n35564_not
g89604 not n48542 ; n48542_not
g89605 not n35573 ; n35573_not
g89606 not n46328 ; n46328_not
g89607 not n27149 ; n27149_not
g89608 not n35582 ; n35582_not
g89609 not n35627 ; n35627_not
g89610 not n46337 ; n46337_not
g89611 not n48533 ; n48533_not
g89612 not n35618 ; n35618_not
g89613 not n48623 ; n48623_not
g89614 not n48407 ; n48407_not
g89615 not n36356 ; n36356_not
g89616 not n36347 ; n36347_not
g89617 not n35735 ; n35735_not
g89618 not n36581 ; n36581_not
g89619 not n46265 ; n46265_not
g89620 not n49217 ; n49217_not
g89621 not n26924 ; n26924_not
g89622 not n45734 ; n45734_not
g89623 not n48371 ; n48371_not
g89624 not n36374 ; n36374_not
g89625 not n48632 ; n48632_not
g89626 not n39551 ; n39551_not
g89627 not n48380 ; n48380_not
g89628 not n46274 ; n46274_not
g89629 not n36365 ; n36365_not
g89630 not n36284 ; n36284_not
g89631 not n35474 ; n35474_not
g89632 not n48605 ; n48605_not
g89633 not n46292 ; n46292_not
g89634 not n36275 ; n36275_not
g89635 not n35483 ; n35483_not
g89636 not n36266 ; n36266_not
g89637 not n51791 ; n51791_not
g89638 not n35492 ; n35492_not
g89639 not n49235 ; n49235_not
g89640 not n36338 ; n36338_not
g89641 not n36608 ; n36608_not
g89642 not n46283 ; n46283_not
g89643 not n36329 ; n36329_not
g89644 not n35429 ; n35429_not
g89645 not n35708 ; n35708_not
g89646 not n35438 ; n35438_not
g89647 not n39524 ; n39524_not
g89648 not n35447 ; n35447_not
g89649 not n35456 ; n35456_not
g89650 not n49226 ; n49226_not
g89651 not n36626 ; n36626_not
g89652 not n35465 ; n35465_not
g89653 not n36293 ; n36293_not
g89654 not n35690 ; n35690_not
g89655 not n48227 ; n48227_not
g89656 not n36068 ; n36068_not
g89657 not n36059 ; n36059_not
g89658 not n26546 ; n26546_not
g89659 not n48155 ; n48155_not
g89660 not n48236 ; n48236_not
g89661 not n48713 ; n48713_not
g89662 not n48245 ; n48245_not
g89663 not n48164 ; n48164_not
g89664 not n48191 ; n48191_not
g89665 not n48146 ; n48146_not
g89666 not n36086 ; n36086_not
g89667 not n26528 ; n26528_not
g89668 not n48209 ; n48209_not
g89669 not n48731 ; n48731_not
g89670 not n48218 ; n48218_not
g89671 not n26537 ; n26537_not
g89672 not n48722 ; n48722_not
g89673 not n26573 ; n26573_not
g89674 not n48182 ; n48182_not
g89675 not n48740 ; n48740_not
g89676 not n49037 ; n49037_not
g89677 not n26582 ; n26582_not
g89678 not n49046 ; n49046_not
g89679 not n26555 ; n26555_not
g89680 not n35636 ; n35636_not
g89681 not n26564 ; n26564_not
g89682 not n49019 ; n49019_not
g89683 not n48173 ; n48173_not
g89684 not n49028 ; n49028_not
g89685 not n26483 ; n26483_not
g89686 not n48083 ; n48083_not
g89687 not n48092 ; n48092_not
g89688 not n48830 ; n48830_not
g89689 not n36194 ; n36194_not
g89690 not n26492 ; n26492_not
g89691 not n39632 ; n39632_not
g89692 not n36167 ; n36167_not
g89693 not n48119 ; n48119_not
g89694 not n48803 ; n48803_not
g89695 not n45905 ; n45905_not
g89696 not n26474 ; n26474_not
g89697 not n48128 ; n48128_not
g89698 not n45914 ; n45914_not
g89699 not n26285 ; n26285_not
g89700 not n36149 ; n36149_not
g89701 not n48902 ; n48902_not
g89702 not n48911 ; n48911_not
g89703 not n48137 ; n48137_not
g89704 not n26519 ; n26519_not
g89705 not n48920 ; n48920_not
g89706 not n36158 ; n36158_not
g89707 not n36176 ; n36176_not
g89708 not n48641 ; n48641_not
g89709 not n26717 ; n26717_not
g89710 not n49109 ; n49109_not
g89711 not n26726 ; n26726_not
g89712 not n39713 ; n39713_not
g89713 not n39209 ; n39209_not
g89714 not n26690 ; n26690_not
g89715 not n49091 ; n49091_not
g89716 not n39722 ; n39722_not
g89717 not n36077 ; n36077_not
g89718 not n26708 ; n26708_not
g89719 not n39245 ; n39245_not
g89720 not n26753 ; n26753_not
g89721 not n39254 ; n39254_not
g89722 not n49136 ; n49136_not
g89723 not n39263 ; n39263_not
g89724 not n26762 ; n26762_not
g89725 not n26735 ; n26735_not
g89726 not n39218 ; n39218_not
g89727 not n39704 ; n39704_not
g89728 not n49118 ; n49118_not
g89729 not n39227 ; n39227_not
g89730 not n26744 ; n26744_not
g89731 not n49127 ; n49127_not
g89732 not n39236 ; n39236_not
g89733 not n26618 ; n26618_not
g89734 not n26627 ; n26627_not
g89735 not n49064 ; n49064_not
g89736 not n26636 ; n26636_not
g89737 not n26591 ; n26591_not
g89738 not n49055 ; n49055_not
g89739 not n26609 ; n26609_not
g89740 not n45824 ; n45824_not
g89741 not n49082 ; n49082_not
g89742 not n26672 ; n26672_not
g89743 not n26195 ; n26195_not
g89744 not n26681 ; n26681_not
g89745 not n26645 ; n26645_not
g89746 not n49073 ; n49073_not
g89747 not n26654 ; n26654_not
g89748 not n35681 ; n35681_not
g89749 not n26663 ; n26663_not
g89750 not n27563 ; n27563_not
g89751 not n27284 ; n27284_not
g89752 not n27428 ; n27428_not
g89753 not n27545 ; n27545_not
g89754 not n27374 ; n27374_not
g89755 not n49307 ; n49307_not
g89756 not n27437 ; n27437_not
g89757 not n49262 ; n49262_not
g89758 not n27473 ; n27473_not
g89759 not n39083 ; n39083_not
g89760 not n27527 ; n27527_not
g89761 not n35276 ; n35276_not
g89762 not n27392 ; n27392_not
g89763 not n27491 ; n27491_not
g89764 not n27329 ; n27329_not
g89765 not n51836 ; n51836_not
g89766 not n27419 ; n27419_not
g89767 not n27572 ; n27572_not
g89768 not n27383 ; n27383_not
g89769 not n27347 ; n27347_not
g89770 not n27239 ; n27239_not
g89771 not n27536 ; n27536_not
g89772 not n27248 ; n27248_not
g89773 not n48551 ; n48551_not
g89774 not n27338 ; n27338_not
g89775 not n27257 ; n27257_not
g89776 not n27581 ; n27581_not
g89777 not n27518 ; n27518_not
g89778 not n27509 ; n27509_not
g89779 not n27356 ; n27356_not
g89780 not n49280 ; n49280_not
g89781 not n27365 ; n27365_not
g89782 not n27482 ; n27482_not
g89783 not n36617 ; n36617_not
g89784 not n46445 ; n46445_not
g89785 not n51881 ; n51881_not
g89786 not n27554 ; n27554_not
g89787 not n27455 ; n27455_not
g89788 not n27275 ; n27275_not
g89789 not n27095 ; n27095_not
g89790 not n49271 ; n49271_not
g89791 not n39038 ; n39038_not
g89792 not n47822 ; n47822_not
g89793 not n27185 ; n27185_not
g89794 not n27590 ; n27590_not
g89795 not n27464 ; n27464_not
g89796 not n27293 ; n27293_not
g89797 not n27266 ; n27266_not
g89798 not n27446 ; n27446_not
g89799 not n55743 ; n55743_not
g89800 not n16683 ; n16683_not
g89801 not n16638 ; n16638_not
g89802 not n56454 ; n56454_not
g89803 not n56472 ; n56472_not
g89804 not n16692 ; n16692_not
g89805 not n49065 ; n49065_not
g89806 not n35268 ; n35268_not
g89807 not n13965 ; n13965_not
g89808 not n16593 ; n16593_not
g89809 not n55590 ; n55590_not
g89810 not n55608 ; n55608_not
g89811 not n55734 ; n55734_not
g89812 not n37833 ; n37833_not
g89813 not n31794 ; n31794_not
g89814 not n56445 ; n56445_not
g89815 not n55491 ; n55491_not
g89816 not n47913 ; n47913_not
g89817 not n42576 ; n42576_not
g89818 not n37824 ; n37824_not
g89819 not n37509 ; n37509_not
g89820 not n55635 ; n55635_not
g89821 not n55617 ; n55617_not
g89822 not n37518 ; n37518_not
g89823 not n16629 ; n16629_not
g89824 not n42585 ; n42585_not
g89825 not n16656 ; n16656_not
g89826 not n13974 ; n13974_not
g89827 not n16665 ; n16665_not
g89828 not n31929 ; n31929_not
g89829 not n35673 ; n35673_not
g89830 not n55077 ; n55077_not
g89831 not n16575 ; n16575_not
g89832 not n55482 ; n55482_not
g89833 not n55626 ; n55626_not
g89834 not n56481 ; n56481_not
g89835 not n31938 ; n31938_not
g89836 not n16566 ; n16566_not
g89837 not n35277 ; n35277_not
g89838 not n17169 ; n17169_not
g89839 not n16557 ; n16557_not
g89840 not n56490 ; n56490_not
g89841 not n16647 ; n16647_not
g89842 not n42594 ; n42594_not
g89843 not n35925 ; n35925_not
g89844 not n56463 ; n56463_not
g89845 not n16584 ; n16584_not
g89846 not n17178 ; n17178_not
g89847 not n43854 ; n43854_not
g89848 not n16548 ; n16548_not
g89849 not n44439 ; n44439_not
g89850 not n16674 ; n16674_not
g89851 not n56571 ; n56571_not
g89852 not n17079 ; n17079_not
g89853 not n49047 ; n49047_not
g89854 not n55851 ; n55851_not
g89855 not n17376 ; n17376_not
g89856 not n47247 ; n47247_not
g89857 not n31848 ; n31848_not
g89858 not n17367 ; n17367_not
g89859 not n17088 ; n17088_not
g89860 not n44781 ; n44781_not
g89861 not n55707 ; n55707_not
g89862 not n31749 ; n31749_not
g89863 not n17358 ; n17358_not
g89864 not n17097 ; n17097_not
g89865 not n56562 ; n56562_not
g89866 not n17349 ; n17349_not
g89867 not n56553 ; n56553_not
g89868 not n44466 ; n44466_not
g89869 not n55716 ; n55716_not
g89870 not n31857 ; n31857_not
g89871 not n48723 ; n48723_not
g89872 not n56544 ; n56544_not
g89873 not n45249 ; n45249_not
g89874 not n44394 ; n44394_not
g89875 not n44484 ; n44484_not
g89876 not n55833 ; n55833_not
g89877 not n43881 ; n43881_not
g89878 not n42657 ; n42657_not
g89879 not n31767 ; n31767_not
g89880 not n49290 ; n49290_not
g89881 not n55509 ; n55509_not
g89882 not n37482 ; n37482_not
g89883 not n31758 ; n31758_not
g89884 not n42666 ; n42666_not
g89885 not n50586 ; n50586_not
g89886 not n55725 ; n55725_not
g89887 not n55842 ; n55842_not
g89888 not n56580 ; n56580_not
g89889 not n17394 ; n17394_not
g89890 not n36870 ; n36870_not
g89891 not n31839 ; n31839_not
g89892 not n48732 ; n48732_not
g89893 not n47256 ; n47256_not
g89894 not n45258 ; n45258_not
g89895 not n17385 ; n17385_not
g89896 not n55662 ; n55662_not
g89897 not n43863 ; n43863_not
g89898 not n49056 ; n49056_not
g89899 not n35295 ; n35295_not
g89900 not n44961 ; n44961_not
g89901 not n31893 ; n31893_not
g89902 not n37842 ; n37842_not
g89903 not n55059 ; n55059_not
g89904 not n44457 ; n44457_not
g89905 not n56517 ; n56517_not
g89906 not n49407 ; n49407_not
g89907 not n12939 ; n12939_not
g89908 not n55653 ; n55653_not
g89909 not n50568 ; n50568_not
g89910 not n13947 ; n13947_not
g89911 not n44448 ; n44448_not
g89912 not n17196 ; n17196_not
g89913 not n56508 ; n56508_not
g89914 not n55644 ; n55644_not
g89915 not n35934 ; n35934_not
g89916 not n17187 ; n17187_not
g89917 not n13929 ; n13929_not
g89918 not n47238 ; n47238_not
g89919 not n31866 ; n31866_not
g89920 not n17295 ; n17295_not
g89921 not n55680 ; n55680_not
g89922 not n49380 ; n49380_not
g89923 not n37860 ; n37860_not
g89924 not n17286 ; n17286_not
g89925 not n35943 ; n35943_not
g89926 not n12948 ; n12948_not
g89927 not n56535 ; n56535_not
g89928 not n17277 ; n17277_not
g89929 not n31875 ; n31875_not
g89930 not n17268 ; n17268_not
g89931 not n50577 ; n50577_not
g89932 not n55671 ; n55671_not
g89933 not n17259 ; n17259_not
g89934 not n37851 ; n37851_not
g89935 not n12786 ; n12786_not
g89936 not n31884 ; n31884_not
g89937 not n56526 ; n56526_not
g89938 not n55464 ; n55464_not
g89939 not n16854 ; n16854_not
g89940 not n35169 ; n35169_not
g89941 not n16197 ; n16197_not
g89942 not n37761 ; n37761_not
g89943 not n16845 ; n16845_not
g89944 not n12885 ; n12885_not
g89945 not n48642 ; n48642_not
g89946 not n56319 ; n56319_not
g89947 not n55455 ; n55455_not
g89948 not n16188 ; n16188_not
g89949 not n55185 ; n55185_not
g89950 not n16836 ; n16836_not
g89951 not n34773 ; n34773_not
g89952 not n37554 ; n37554_not
g89953 not n55248 ; n55248_not
g89954 not n16179 ; n16179_not
g89955 not n44358 ; n44358_not
g89956 not n16827 ; n16827_not
g89957 not n37752 ; n37752_not
g89958 not n43818 ; n43818_not
g89959 not n49281 ; n49281_not
g89960 not n13857 ; n13857_not
g89961 not n16818 ; n16818_not
g89962 not n36780 ; n36780_not
g89963 not n31947 ; n31947_not
g89964 not n16908 ; n16908_not
g89965 not n49092 ; n49092_not
g89966 not n47193 ; n47193_not
g89967 not n35691 ; n35691_not
g89968 not n55167 ; n55167_not
g89969 not n54933 ; n54933_not
g89970 not n12894 ; n12894_not
g89971 not n16890 ; n16890_not
g89972 not n16881 ; n16881_not
g89973 not n56337 ; n56337_not
g89974 not n55473 ; n55473_not
g89975 not n13875 ; n13875_not
g89976 not n56328 ; n56328_not
g89977 not n16872 ; n16872_not
g89978 not n37770 ; n37770_not
g89979 not n13866 ; n13866_not
g89980 not n16863 ; n16863_not
g89981 not n49425 ; n49425_not
g89982 not n43809 ; n43809_not
g89983 not n47157 ; n47157_not
g89984 not n16098 ; n16098_not
g89985 not n49434 ; n49434_not
g89986 not n16746 ; n16746_not
g89987 not n37572 ; n37572_not
g89988 not n54915 ; n54915_not
g89989 not n32379 ; n32379_not
g89990 not n56292 ; n56292_not
g89991 not n16089 ; n16089_not
g89992 not n37725 ; n37725_not
g89993 not n48633 ; n48633_not
g89994 not n16737 ; n16737_not
g89995 not n42495 ; n42495_not
g89996 not n49119 ; n49119_not
g89997 not n16728 ; n16728_not
g89998 not n55428 ; n55428_not
g89999 not n50496 ; n50496_not
g90000 not n16395 ; n16395_not
g90001 not n54924 ; n54924_not
g90002 not n16719 ; n16719_not
g90003 not n35871 ; n35871_not
g90004 not n47832 ; n47832_not
g90005 not n14199 ; n14199_not
g90006 not n37716 ; n37716_not
g90007 not n47148 ; n47148_not
g90008 not n32199 ; n32199_not
g90009 not n55446 ; n55446_not
g90010 not n36069 ; n36069_not
g90011 not n16809 ; n16809_not
g90012 not n35880 ; n35880_not
g90013 not n55194 ; n55194_not
g90014 not n31974 ; n31974_not
g90015 not n37743 ; n37743_not
g90016 not n45186 ; n45186_not
g90017 not n16791 ; n16791_not
g90018 not n36906 ; n36906_not
g90019 not n16359 ; n16359_not
g90020 not n16782 ; n16782_not
g90021 not n44349 ; n44349_not
g90022 not n16368 ; n16368_not
g90023 not n10599 ; n10599_not
g90024 not n16773 ; n16773_not
g90025 not n47166 ; n47166_not
g90026 not n16764 ; n16764_not
g90027 not n37563 ; n37563_not
g90028 not n45177 ; n45177_not
g90029 not n32289 ; n32289_not
g90030 not n37734 ; n37734_not
g90031 not n55437 ; n55437_not
g90032 not n16755 ; n16755_not
g90033 not n12876 ; n12876_not
g90034 not n13983 ; n13983_not
g90035 not n56418 ; n56418_not
g90036 not n55932 ; n55932_not
g90037 not n55554 ; n55554_not
g90038 not n37527 ; n37527_not
g90039 not n56409 ; n56409_not
g90040 not n31956 ; n31956_not
g90041 not n55941 ; n55941_not
g90042 not n55752 ; n55752_not
g90043 not n55545 ; n55545_not
g90044 not n55536 ; n55536_not
g90045 not n37806 ; n37806_not
g90046 not n35187 ; n35187_not
g90047 not n36078 ; n36078_not
g90048 not n37815 ; n37815_not
g90049 not n55581 ; n55581_not
g90050 not n56436 ; n56436_not
g90051 not n44880 ; n44880_not
g90052 not n55923 ; n55923_not
g90053 not n49074 ; n49074_not
g90054 not n55095 ; n55095_not
g90055 not n55572 ; n55572_not
g90056 not n36087 ; n36087_not
g90057 not n56427 ; n56427_not
g90058 not n35916 ; n35916_not
g90059 not n35178 ; n35178_not
g90060 not n55563 ; n55563_not
g90061 not n43836 ; n43836_not
g90062 not n35682 ; n35682_not
g90063 not n56364 ; n56364_not
g90064 not n55770 ; n55770_not
g90065 not n16278 ; n16278_not
g90066 not n42549 ; n42549_not
g90067 not n16935 ; n16935_not
g90068 not n31983 ; n31983_not
g90069 not n56355 ; n56355_not
g90070 not n44970 ; n44970_not
g90071 not n16926 ; n16926_not
g90072 not n31965 ; n31965_not
g90073 not n48651 ; n48651_not
g90074 not n44376 ; n44376_not
g90075 not n34764 ; n34764_not
g90076 not n16917 ; n16917_not
g90077 not n56346 ; n56346_not
g90078 not n56391 ; n56391_not
g90079 not n13992 ; n13992_not
g90080 not n31677 ; n31677_not
g90081 not n49083 ; n49083_not
g90082 not n55761 ; n55761_not
g90083 not n47922 ; n47922_not
g90084 not n55527 ; n55527_not
g90085 not n55815 ; n55815_not
g90086 not n44790 ; n44790_not
g90087 not n35907 ; n35907_not
g90088 not n56382 ; n56382_not
g90089 not n16971 ; n16971_not
g90090 not n55518 ; n55518_not
g90091 not n50559 ; n50559_not
g90092 not n36609 ; n36609_not
g90093 not n55149 ; n55149_not
g90094 not n56373 ; n56373_not
g90095 not n38058 ; n38058_not
g90096 not n57246 ; n57246_not
g90097 not n17835 ; n17835_not
g90098 not n54816 ; n54816_not
g90099 not n36159 ; n36159_not
g90100 not n55905 ; n55905_not
g90101 not n30993 ; n30993_not
g90102 not n50667 ; n50667_not
g90103 not n49344 ; n49344_not
g90104 not n42396 ; n42396_not
g90105 not n44718 ; n44718_not
g90106 not n30984 ; n30984_not
g90107 not n44538 ; n44538_not
g90108 not n45276 ; n45276_not
g90109 not n30777 ; n30777_not
g90110 not n42387 ; n42387_not
g90111 not n36807 ; n36807_not
g90112 not n44628 ; n44628_not
g90113 not n57228 ; n57228_not
g90114 not n17817 ; n17817_not
g90115 not n36843 ; n36843_not
g90116 not n42378 ; n42378_not
g90117 not n47328 ; n47328_not
g90118 not n54393 ; n54393_not
g90119 not n44646 ; n44646_not
g90120 not n17880 ; n17880_not
g90121 not n17871 ; n17871_not
g90122 not n44934 ; n44934_not
g90123 not n57291 ; n57291_not
g90124 not n43971 ; n43971_not
g90125 not n57282 ; n57282_not
g90126 not n54807 ; n54807_not
g90127 not n36582 ; n36582_not
g90128 not n57273 ; n57273_not
g90129 not n17862 ; n17862_not
g90130 not n56850 ; n56850_not
g90131 not n44637 ; n44637_not
g90132 not n50676 ; n50676_not
g90133 not n56841 ; n56841_not
g90134 not n17844 ; n17844_not
g90135 not n43935 ; n43935_not
g90136 not n36168 ; n36168_not
g90137 not n57174 ; n57174_not
g90138 not n17772 ; n17772_not
g90139 not n48912 ; n48912_not
g90140 not n57156 ; n57156_not
g90141 not n43917 ; n43917_not
g90142 not n42468 ; n42468_not
g90143 not n30849 ; n30849_not
g90144 not n57147 ; n57147_not
g90145 not n30939 ; n30939_not
g90146 not n54834 ; n54834_not
g90147 not n30858 ; n30858_not
g90148 not n48921 ; n48921_not
g90149 not n17754 ; n17754_not
g90150 not n30867 ; n30867_not
g90151 not n17745 ; n17745_not
g90152 not n57138 ; n57138_not
g90153 not n57129 ; n57129_not
g90154 not n46653 ; n46653_not
g90155 not n36096 ; n36096_not
g90156 not n30876 ; n30876_not
g90157 not n30885 ; n30885_not
g90158 not n50658 ; n50658_not
g90159 not n42369 ; n42369_not
g90160 not n30786 ; n30786_not
g90161 not n17790 ; n17790_not
g90162 not n13749 ; n13749_not
g90163 not n44547 ; n44547_not
g90164 not n54825 ; n54825_not
g90165 not n57219 ; n57219_not
g90166 not n43926 ; n43926_not
g90167 not n30795 ; n30795_not
g90168 not n50649 ; n50649_not
g90169 not n44907 ; n44907_not
g90170 not n30957 ; n30957_not
g90171 not n47337 ; n47337_not
g90172 not n30948 ; n30948_not
g90173 not n44619 ; n44619_not
g90174 not n36573 ; n36573_not
g90175 not n48903 ; n48903_not
g90176 not n56814 ; n56814_not
g90177 not n56805 ; n56805_not
g90178 not n30768 ; n30768_not
g90179 not n47283 ; n47283_not
g90180 not n41838 ; n41838_not
g90181 not n54726 ; n54726_not
g90182 not n44682 ; n44682_not
g90183 not n57426 ; n57426_not
g90184 not n47292 ; n47292_not
g90185 not n17961 ; n17961_not
g90186 not n54186 ; n54186_not
g90187 not n36825 ; n36825_not
g90188 not n57417 ; n57417_not
g90189 not n43953 ; n43953_not
g90190 not n36177 ; n36177_not
g90191 not n54735 ; n54735_not
g90192 not n17952 ; n17952_not
g90193 not n56940 ; n56940_not
g90194 not n56931 ; n56931_not
g90195 not n44925 ; n44925_not
g90196 not n57390 ; n57390_not
g90197 not n50694 ; n50694_not
g90198 not n44673 ; n44673_not
g90199 not n43962 ; n43962_not
g90200 not n54681 ; n54681_not
g90201 not n30696 ; n30696_not
g90202 not n57462 ; n57462_not
g90203 not n41847 ; n41847_not
g90204 not n54690 ; n54690_not
g90205 not n17808 ; n17808_not
g90206 not n44691 ; n44691_not
g90207 not n48804 ; n48804_not
g90208 not n54708 ; n54708_not
g90209 not n54195 ; n54195_not
g90210 not n30894 ; n30894_not
g90211 not n57444 ; n57444_not
g90212 not n48066 ; n48066_not
g90213 not n30687 ; n30687_not
g90214 not n54717 ; n54717_not
g90215 not n57435 ; n57435_not
g90216 not n17970 ; n17970_not
g90217 not n57354 ; n57354_not
g90218 not n54762 ; n54762_not
g90219 not n17916 ; n17916_not
g90220 not n17853 ; n17853_not
g90221 not n56904 ; n56904_not
g90222 not n44655 ; n44655_not
g90223 not n57345 ; n57345_not
g90224 not n17907 ; n17907_not
g90225 not n48831 ; n48831_not
g90226 not n30966 ; n30966_not
g90227 not n54771 ; n54771_not
g90228 not n50685 ; n50685_not
g90229 not n48840 ; n48840_not
g90230 not n49317 ; n49317_not
g90231 not n57318 ; n57318_not
g90232 not n54780 ; n54780_not
g90233 not n54159 ; n54159_not
g90234 not n36186 ; n36186_not
g90235 not n44529 ; n44529_not
g90236 not n17943 ; n17943_not
g90237 not n44916 ; n44916_not
g90238 not n57372 ; n57372_not
g90239 not n54744 ; n54744_not
g90240 not n35286 ; n35286_not
g90241 not n36816 ; n36816_not
g90242 not n38085 ; n38085_not
g90243 not n35763 ; n35763_not
g90244 not n44664 ; n44664_not
g90245 not n44709 ; n44709_not
g90246 not n17934 ; n17934_not
g90247 not n43944 ; n43944_not
g90248 not n57363 ; n57363_not
g90249 not n49335 ; n49335_not
g90250 not n36834 ; n36834_not
g90251 not n54753 ; n54753_not
g90252 not n44493 ; n44493_not
g90253 not n38076 ; n38076_not
g90254 not n17925 ; n17925_not
g90255 not n36564 ; n36564_not
g90256 not n35637 ; n35637_not
g90257 not n17556 ; n17556_not
g90258 not n31668 ; n31668_not
g90259 not n56733 ; n56733_not
g90260 not n45267 ; n45267_not
g90261 not n37932 ; n37932_not
g90262 not n35646 ; n35646_not
g90263 not n54906 ; n54906_not
g90264 not n56715 ; n56715_not
g90265 not n31659 ; n31659_not
g90266 not n55950 ; n55950_not
g90267 not n17547 ; n17547_not
g90268 not n55860 ; n55860_not
g90269 not n31596 ; n31596_not
g90270 not n31587 ; n31587_not
g90271 not n17538 ; n17538_not
g90272 not n56706 ; n56706_not
g90273 not n31578 ; n31578_not
g90274 not n35970 ; n35970_not
g90275 not n42099 ; n42099_not
g90276 not n17529 ; n17529_not
g90277 not n44367 ; n44367_not
g90278 not n17592 ; n17592_not
g90279 not n34935 ; n34935_not
g90280 not n48750 ; n48750_not
g90281 not n44754 ; n44754_not
g90282 not n17583 ; n17583_not
g90283 not n12975 ; n12975_not
g90284 not n37941 ; n37941_not
g90285 not n56823 ; n56823_not
g90286 not n56760 ; n56760_not
g90287 not n54096 ; n54096_not
g90288 not n17574 ; n17574_not
g90289 not n31686 ; n31686_not
g90290 not n44763 ; n44763_not
g90291 not n17565 ; n17565_not
g90292 not n56751 ; n56751_not
g90293 not n35961 ; n35961_not
g90294 not n17475 ; n17475_not
g90295 not n13884 ; n13884_not
g90296 not n44772 ; n44772_not
g90297 not n54960 ; n54960_not
g90298 not n17466 ; n17466_not
g90299 not n56616 ; n56616_not
g90300 not n12957 ; n12957_not
g90301 not n37905 ; n37905_not
g90302 not n17457 ; n17457_not
g90303 not n50595 ; n50595_not
g90304 not n42639 ; n42639_not
g90305 not n17448 ; n17448_not
g90306 not n17439 ; n17439_not
g90307 not n56607 ; n56607_not
g90308 not n49038 ; n49038_not
g90309 not n37473 ; n37473_not
g90310 not n35952 ; n35952_not
g90311 not n37923 ; n37923_not
g90312 not n31569 ; n31569_not
g90313 not n56661 ; n56661_not
g90314 not n56652 ; n56652_not
g90315 not n31776 ; n31776_not
g90316 not n43872 ; n43872_not
g90317 not n55806 ; n55806_not
g90318 not n56643 ; n56643_not
g90319 not n37464 ; n37464_not
g90320 not n47904 ; n47904_not
g90321 not n56634 ; n56634_not
g90322 not n17493 ; n17493_not
g90323 not n44952 ; n44952_not
g90324 not n37914 ; n37914_not
g90325 not n12966 ; n12966_not
g90326 not n31785 ; n31785_not
g90327 not n49029 ; n49029_not
g90328 not n54942 ; n54942_not
g90329 not n56625 ; n56625_not
g90330 not n17484 ; n17484_not
g90331 not n42279 ; n42279_not
g90332 not n44736 ; n44736_not
g90333 not n57075 ; n57075_not
g90334 not n17709 ; n17709_not
g90335 not n57066 ; n57066_not
g90336 not n44574 ; n44574_not
g90337 not n54843 ; n54843_not
g90338 not n13794 ; n13794_not
g90339 not n43908 ; n43908_not
g90340 not n31398 ; n31398_not
g90341 not n56724 ; n56724_not
g90342 not n31389 ; n31389_not
g90343 not n17682 ; n17682_not
g90344 not n57057 ; n57057_not
g90345 not n54852 ; n54852_not
g90346 not n44727 ; n44727_not
g90347 not n43980 ; n43980_not
g90348 not n46644 ; n46644_not
g90349 not n42486 ; n42486_not
g90350 not n36852 ; n36852_not
g90351 not n42297 ; n42297_not
g90352 not n48741 ; n48741_not
g90353 not n17727 ; n17727_not
g90354 not n44943 ; n44943_not
g90355 not n48930 ; n48930_not
g90356 not n13767 ; n13767_not
g90357 not n42288 ; n42288_not
g90358 not n12993 ; n12993_not
g90359 not n57084 ; n57084_not
g90360 not n13776 ; n13776_not
g90361 not n37950 ; n37950_not
g90362 not n31479 ; n31479_not
g90363 not n42198 ; n42198_not
g90364 not n17637 ; n17637_not
g90365 not n13839 ; n13839_not
g90366 not n36861 ; n36861_not
g90367 not n17628 ; n17628_not
g90368 not n42189 ; n42189_not
g90369 not n44556 ; n44556_not
g90370 not n49362 ; n49362_not
g90371 not n56913 ; n56913_not
g90372 not n35628 ; n35628_not
g90373 not n42558 ; n42558_not
g90374 not n16962 ; n16962_not
g90375 not n54870 ; n54870_not
g90376 not n31488 ; n31488_not
g90377 not n31299 ; n31299_not
g90378 not n17664 ; n17664_not
g90379 not n44745 ; n44745_not
g90380 not n17655 ; n17655_not
g90381 not n12984 ; n12984_not
g90382 not n54861 ; n54861_not
g90383 not n48039 ; n48039_not
g90384 not n49920 ; n49920_not
g90385 not n49740 ; n49740_not
g90386 not n15729 ; n15729_not
g90387 not n48048 ; n48048_not
g90388 not n37059 ; n37059_not
g90389 not n14793 ; n14793_not
g90390 not n12399 ; n12399_not
g90391 not n43368 ; n43368_not
g90392 not n47346 ; n47346_not
g90393 not n55257 ; n55257_not
g90394 not n54555 ; n54555_not
g90395 not n36636 ; n36636_not
g90396 not n43377 ; n43377_not
g90397 not n15684 ; n15684_not
g90398 not n34098 ; n34098_not
g90399 not n55266 ; n55266_not
g90400 not n48057 ; n48057_not
g90401 not n15666 ; n15666_not
g90402 not n44178 ; n44178_not
g90403 not n33918 ; n33918_not
g90404 not n15774 ; n15774_not
g90405 not n49227 ; n49227_not
g90406 not n49821 ; n49821_not
g90407 not n33927 ; n33927_not
g90408 not n14784 ; n14784_not
g90409 not n33936 ; n33936_not
g90410 not n49830 ; n49830_not
g90411 not n33945 ; n33945_not
g90412 not n33954 ; n33954_not
g90413 not n49470 ; n49470_not
g90414 not n33963 ; n33963_not
g90415 not n45087 ; n45087_not
g90416 not n15756 ; n15756_not
g90417 not n33972 ; n33972_not
g90418 not n33981 ; n33981_not
g90419 not n49902 ; n49902_not
g90420 not n43638 ; n43638_not
g90421 not n15747 ; n15747_not
g90422 not n33990 ; n33990_not
g90423 not n49911 ; n49911_not
g90424 not n44187 ; n44187_not
g90425 not n43359 ; n43359_not
g90426 not n14982 ; n14982_not
g90427 not n15594 ; n15594_not
g90428 not n49236 ; n49236_not
g90429 not n54573 ; n54573_not
g90430 not n55284 ; n55284_not
g90431 not n34368 ; n34368_not
g90432 not n14847 ; n14847_not
g90433 not n55293 ; n55293_not
g90434 not n15585 ; n15585_not
g90435 not n34377 ; n34377_not
g90436 not n15576 ; n15576_not
g90437 not n34908 ; n34908_not
g90438 not n43197 ; n43197_not
g90439 not n54582 ; n54582_not
g90440 not n15567 ; n15567_not
g90441 not n34386 ; n34386_not
g90442 not n34395 ; n34395_not
g90443 not n49308 ; n49308_not
g90444 not n15558 ; n15558_not
g90445 not n12498 ; n12498_not
g90446 not n43773 ; n43773_not
g90447 not n43386 ; n43386_not
g90448 not n15657 ; n15657_not
g90449 not n43764 ; n43764_not
g90450 not n43629 ; n43629_not
g90451 not n36744 ; n36744_not
g90452 not n12489 ; n12489_not
g90453 not n37086 ; n37086_not
g90454 not n14829 ; n14829_not
g90455 not n55275 ; n55275_not
g90456 not n43395 ; n43395_not
g90457 not n14838 ; n14838_not
g90458 not n15639 ; n15639_not
g90459 not n56085 ; n56085_not
g90460 not n44169 ; n44169_not
g90461 not n44835 ; n44835_not
g90462 not n54564 ; n54564_not
g90463 not n37095 ; n37095_not
g90464 not n33684 ; n33684_not
g90465 not n49605 ; n49605_not
g90466 not n11967 ; n11967_not
g90467 not n14748 ; n14748_not
g90468 not n34890 ; n34890_not
g90469 not n50298 ; n50298_not
g90470 not n33729 ; n33729_not
g90471 not n49614 ; n49614_not
g90472 not n43296 ; n43296_not
g90473 not n45096 ; n45096_not
g90474 not n49722 ; n49722_not
g90475 not n14757 ; n14757_not
g90476 not n11985 ; n11985_not
g90477 not n33738 ; n33738_not
g90478 not n33747 ; n33747_not
g90479 not n54519 ; n54519_not
g90480 not n56157 ; n56157_not
g90481 not n35727 ; n35727_not
g90482 not n33756 ; n33756_not
g90483 not n49623 ; n49623_not
g90484 not n49704 ; n49704_not
g90485 not n14487 ; n14487_not
g90486 not n33558 ; n33558_not
g90487 not n43269 ; n43269_not
g90488 not n33288 ; n33288_not
g90489 not n33567 ; n33567_not
g90490 not n33279 ; n33279_not
g90491 not n36591 ; n36591_not
g90492 not n33576 ; n33576_not
g90493 not n49713 ; n49713_not
g90494 not n56166 ; n56166_not
g90495 not n35745 ; n35745_not
g90496 not n33585 ; n33585_not
g90497 not n34953 ; n34953_not
g90498 not n33594 ; n33594_not
g90499 not n47814 ; n47814_not
g90500 not n33639 ; n33639_not
g90501 not n14739 ; n14739_not
g90502 not n48615 ; n48615_not
g90503 not n33657 ; n33657_not
g90504 not n43287 ; n43287_not
g90505 not n56076 ; n56076_not
g90506 not n49218 ; n49218_not
g90507 not n33666 ; n33666_not
g90508 not n43656 ; n43656_not
g90509 not n15846 ; n15846_not
g90510 not n14775 ; n14775_not
g90511 not n15837 ; n15837_not
g90512 not n33855 ; n33855_not
g90513 not n49731 ; n49731_not
g90514 not n56139 ; n56139_not
g90515 not n34944 ; n34944_not
g90516 not n33864 ; n33864_not
g90517 not n15819 ; n15819_not
g90518 not n33675 ; n33675_not
g90519 not n33873 ; n33873_not
g90520 not n33882 ; n33882_not
g90521 not n44196 ; n44196_not
g90522 not n54537 ; n54537_not
g90523 not n33891 ; n33891_not
g90524 not n49803 ; n49803_not
g90525 not n36618 ; n36618_not
g90526 not n15792 ; n15792_not
g90527 not n49812 ; n49812_not
g90528 not n33909 ; n33909_not
g90529 not n54546 ; n54546_not
g90530 not n35718 ; n35718_not
g90531 not n56148 ; n56148_not
g90532 not n33765 ; n33765_not
g90533 not n14766 ; n14766_not
g90534 not n49632 ; n49632_not
g90535 not n33774 ; n33774_not
g90536 not n55158 ; n55158_not
g90537 not n54528 ; n54528_not
g90538 not n49641 ; n49641_not
g90539 not n33783 ; n33783_not
g90540 not n49650 ; n49650_not
g90541 not n33792 ; n33792_not
g90542 not n33819 ; n33819_not
g90543 not n15855 ; n15855_not
g90544 not n43647 ; n43647_not
g90545 not n44826 ; n44826_not
g90546 not n33828 ; n33828_not
g90547 not n33837 ; n33837_not
g90548 not n33846 ; n33846_not
g90549 not n14919 ; n14919_not
g90550 not n15198 ; n15198_not
g90551 not n34719 ; n34719_not
g90552 not n14928 ; n14928_not
g90553 not n48561 ; n48561_not
g90554 not n34728 ; n34728_not
g90555 not n14586 ; n14586_not
g90556 not n15189 ; n15189_not
g90557 not n34854 ; n34854_not
g90558 not n36717 ; n36717_not
g90559 not n55365 ; n55365_not
g90560 not n54672 ; n54672_not
g90561 not n44097 ; n44097_not
g90562 not n34737 ; n34737_not
g90563 not n14937 ; n14937_not
g90564 not n43584 ; n43584_not
g90565 not n15099 ; n15099_not
g90566 not n34746 ; n34746_not
g90567 not n44862 ; n44862_not
g90568 not n44079 ; n44079_not
g90569 not n55347 ; n55347_not
g90570 not n48534 ; n48534_not
g90571 not n12687 ; n12687_not
g90572 not n43494 ; n43494_not
g90573 not n34674 ; n34674_not
g90574 not n49353 ; n49353_not
g90575 not n36654 ; n36654_not
g90576 not n15297 ; n15297_not
g90577 not n54654 ; n54654_not
g90578 not n12678 ; n12678_not
g90579 not n34683 ; n34683_not
g90580 not n55356 ; n55356_not
g90581 not n15288 ; n15288_not
g90582 not n49263 ; n49263_not
g90583 not n15279 ; n15279_not
g90584 not n34692 ; n34692_not
g90585 not n12669 ; n12669_not
g90586 not n54663 ; n54663_not
g90587 not n36735 ; n36735_not
g90588 not n36708 ; n36708_not
g90589 not n47805 ; n47805_not
g90590 not n55383 ; n55383_not
g90591 not n43557 ; n43557_not
g90592 not n34809 ; n34809_not
g90593 not n35196 ; n35196_not
g90594 not n36753 ; n36753_not
g90595 not n55392 ; n55392_not
g90596 not n43566 ; n43566_not
g90597 not n36762 ; n36762_not
g90598 not n34827 ; n34827_not
g90599 not n14964 ; n14964_not
g90600 not n36771 ; n36771_not
g90601 not n12588 ; n12588_not
g90602 not n43575 ; n43575_not
g90603 not n12597 ; n12597_not
g90604 not n14955 ; n14955_not
g90605 not n12579 ; n12579_not
g90606 not n34845 ; n34845_not
g90607 not n55068 ; n55068_not
g90608 not n43539 ; n43539_not
g90609 not n55374 ; n55374_not
g90610 not n49254 ; n49254_not
g90611 not n36726 ; n36726_not
g90612 not n14946 ; n14946_not
g90613 not n43548 ; n43548_not
g90614 not n48552 ; n48552_not
g90615 not n34782 ; n34782_not
g90616 not n44088 ; n44088_not
g90617 not n12696 ; n12696_not
g90618 not n34548 ; n34548_not
g90619 not n56067 ; n56067_not
g90620 not n15477 ; n15477_not
g90621 not n34485 ; n34485_not
g90622 not n12759 ; n12759_not
g90623 not n15468 ; n15468_not
g90624 not n35655 ; n35655_not
g90625 not n12768 ; n12768_not
g90626 not n34557 ; n34557_not
g90627 not n15459 ; n15459_not
g90628 not n54609 ; n54609_not
g90629 not n43449 ; n43449_not
g90630 not n49443 ; n49443_not
g90631 not n14397 ; n14397_not
g90632 not n34566 ; n34566_not
g90633 not n44844 ; n44844_not
g90634 not n14883 ; n14883_not
g90635 not n34476 ; n34476_not
g90636 not n36663 ; n36663_not
g90637 not n34575 ; n34575_not
g90638 not n12777 ; n12777_not
g90639 not n34458 ; n34458_not
g90640 not n14856 ; n14856_not
g90641 not n15549 ; n15549_not
g90642 not n54591 ; n54591_not
g90643 not n14865 ; n14865_not
g90644 not n43782 ; n43782_not
g90645 not n15495 ; n15495_not
g90646 not n14874 ; n14874_not
g90647 not n15486 ; n15486_not
g90648 not n34539 ; n34539_not
g90649 not n34494 ; n34494_not
g90650 not n55329 ; n55329_not
g90651 not n34638 ; n34638_not
g90652 not n43476 ; n43476_not
g90653 not n15378 ; n15378_not
g90654 not n36690 ; n36690_not
g90655 not n55338 ; n55338_not
g90656 not n15369 ; n15369_not
g90657 not n54636 ; n54636_not
g90658 not n49245 ; n49245_not
g90659 not n44853 ; n44853_not
g90660 not n34647 ; n34647_not
g90661 not n48543 ; n48543_not
g90662 not n43485 ; n43485_not
g90663 not n34656 ; n34656_not
g90664 not n43593 ; n43593_not
g90665 not n34665 ; n34665_not
g90666 not n54645 ; n54645_not
g90667 not n34584 ; n34584_not
g90668 not n43458 ; n43458_not
g90669 not n45069 ; n45069_not
g90670 not n54618 ; n54618_not
g90671 not n48570 ; n48570_not
g90672 not n34872 ; n34872_not
g90673 not n34593 ; n34593_not
g90674 not n56058 ; n56058_not
g90675 not n37068 ; n37068_not
g90676 not n43827 ; n43827_not
g90677 not n15396 ; n15396_not
g90678 not n43467 ; n43467_not
g90679 not n14892 ; n14892_not
g90680 not n54627 ; n54627_not
g90681 not n36672 ; n36672_not
g90682 not n34449 ; n34449_not
g90683 not n15387 ; n15387_not
g90684 not n34629 ; n34629_not
g90685 not n15891 ; n15891_not
g90686 not n37617 ; n37617_not
g90687 not n16485 ; n16485_not
g90688 not n35736 ; n35736_not
g90689 not n37626 ; n37626_not
g90690 not n44808 ; n44808_not
g90691 not n15909 ; n15909_not
g90692 not n49164 ; n49164_not
g90693 not n35808 ; n35808_not
g90694 not n15918 ; n15918_not
g90695 not n44295 ; n44295_not
g90696 not n36519 ; n36519_not
g90697 not n15927 ; n15927_not
g90698 not n15936 ; n15936_not
g90699 not n32595 ; n32595_not
g90700 not n16467 ; n16467_not
g90701 not n56238 ; n56238_not
g90702 not n15945 ; n15945_not
g90703 not n16494 ; n16494_not
g90704 not n32658 ; n32658_not
g90705 not n49155 ; n49155_not
g90706 not n32649 ; n32649_not
g90707 not n15873 ; n15873_not
g90708 not n47823 ; n47823_not
g90709 not n56256 ; n56256_not
g90710 not n15882 ; n15882_not
g90711 not n10995 ; n10995_not
g90712 not n56247 ; n56247_not
g90713 not n36942 ; n36942_not
g90714 not n35817 ; n35817_not
g90715 not n32946 ; n32946_not
g90716 not n37608 ; n37608_not
g90717 not n32892 ; n32892_not
g90718 not n32883 ; n32883_not
g90719 not n14469 ; n14469_not
g90720 not n16377 ; n16377_not
g90721 not n32874 ; n32874_not
g90722 not n36951 ; n36951_not
g90723 not n32865 ; n32865_not
g90724 not n44286 ; n44286_not
g90725 not n49524 ; n49524_not
g90726 not n12795 ; n12795_not
g90727 not n32856 ; n32856_not
g90728 not n55419 ; n55419_not
g90729 not n32964 ; n32964_not
g90730 not n15954 ; n15954_not
g90731 not n32586 ; n32586_not
g90732 not n15963 ; n15963_not
g90733 not n54429 ; n54429_not
g90734 not n10968 ; n10968_not
g90735 not n16449 ; n16449_not
g90736 not n15972 ; n15972_not
g90737 not n32919 ; n32919_not
g90738 not n15981 ; n15981_not
g90739 not n32928 ; n32928_not
g90740 not n10959 ; n10959_not
g90741 not n15990 ; n15990_not
g90742 not n48606 ; n48606_not
g90743 not n49515 ; n49515_not
g90744 not n54438 ; n54438_not
g90745 not n49173 ; n49173_not
g90746 not n36537 ; n36537_not
g90747 not n55239 ; n55239_not
g90748 not n32577 ; n32577_not
g90749 not n35097 ; n35097_not
g90750 not n43791 ; n43791_not
g90751 not n50478 ; n50478_not
g90752 not n12858 ; n12858_not
g90753 not n45159 ; n45159_not
g90754 not n10779 ; n10779_not
g90755 not n49137 ; n49137_not
g90756 not n35853 ; n35853_not
g90757 not n16458 ; n16458_not
g90758 not n10788 ; n10788_not
g90759 not n32667 ; n32667_not
g90760 not n36915 ; n36915_not
g90761 not n10689 ; n10689_not
g90762 not n48705 ; n48705_not
g90763 not n49128 ; n49128_not
g90764 not n12867 ; n12867_not
g90765 not n37707 ; n37707_not
g90766 not n50487 ; n50487_not
g90767 not n10698 ; n10698_not
g90768 not n56283 ; n56283_not
g90769 not n54375 ; n54375_not
g90770 not n32298 ; n32298_not
g90771 not n56274 ; n56274_not
g90772 not n35862 ; n35862_not
g90773 not n49452 ; n49452_not
g90774 not n13785 ; n13785_not
g90775 not n32685 ; n32685_not
g90776 not n14298 ; n14298_not
g90777 not n49146 ; n49146_not
g90778 not n10887 ; n10887_not
g90779 not n36528 ; n36528_not
g90780 not n37662 ; n37662_not
g90781 not n42459 ; n42459_not
g90782 not n35088 ; n35088_not
g90783 not n34818 ; n34818_not
g90784 not n35835 ; n35835_not
g90785 not n14379 ; n14379_not
g90786 not n43692 ; n43692_not
g90787 not n36933 ; n36933_not
g90788 not n35079 ; n35079_not
g90789 not n10977 ; n10977_not
g90790 not n35826 ; n35826_not
g90791 not n37680 ; n37680_not
g90792 not n12849 ; n12849_not
g90793 not n10797 ; n10797_not
g90794 not n36924 ; n36924_not
g90795 not n50469 ; n50469_not
g90796 not n32694 ; n32694_not
g90797 not n35844 ; n35844_not
g90798 not n56265 ; n56265_not
g90799 not n32388 ; n32388_not
g90800 not n43683 ; n43683_not
g90801 not n37671 ; n37671_not
g90802 not n14289 ; n14289_not
g90803 not n32937 ; n32937_not
g90804 not n49209 ; n49209_not
g90805 not n34980 ; n34980_not
g90806 not n14649 ; n14649_not
g90807 not n14658 ; n14658_not
g90808 not n33297 ; n33297_not
g90809 not n33198 ; n33198_not
g90810 not n15765 ; n15765_not
g90811 not n33189 ; n33189_not
g90812 not n56193 ; n56193_not
g90813 not n14667 ; n14667_not
g90814 not n37491 ; n37491_not
g90815 not n54465 ; n54465_not
g90816 not n44259 ; n44259_not
g90817 not n36960 ; n36960_not
g90818 not n49533 ; n49533_not
g90819 not n43179 ; n43179_not
g90820 not n43719 ; n43719_not
g90821 not n36546 ; n36546_not
g90822 not n14595 ; n14595_not
g90823 not n35772 ; n35772_not
g90824 not n33369 ; n33369_not
g90825 not n54492 ; n54492_not
g90826 not n43737 ; n43737_not
g90827 not n14694 ; n14694_not
g90828 not n33459 ; n33459_not
g90829 not n56175 ; n56175_not
g90830 not n33468 ; n33468_not
g90831 not n33477 ; n33477_not
g90832 not n33486 ; n33486_not
g90833 not n33495 ; n33495_not
g90834 not n14496 ; n14496_not
g90835 not n34962 ; n34962_not
g90836 not n43665 ; n43665_not
g90837 not n33549 ; n33549_not
g90838 not n54474 ; n54474_not
g90839 not n37446 ; n37446_not
g90840 not n33099 ; n33099_not
g90841 not n43728 ; n43728_not
g90842 not n14676 ; n14676_not
g90843 not n54483 ; n54483_not
g90844 not n56184 ; n56184_not
g90845 not n33387 ; n33387_not
g90846 not n34971 ; n34971_not
g90847 not n14685 ; n14685_not
g90848 not n33396 ; n33396_not
g90849 not n49272 ; n49272_not
g90850 not n47931 ; n47931_not
g90851 not n33378 ; n33378_not
g90852 not n44817 ; n44817_not
g90853 not n32775 ; n32775_not
g90854 not n32766 ; n32766_not
g90855 not n32757 ; n32757_not
g90856 not n32748 ; n32748_not
g90857 not n32739 ; n32739_not
g90858 not n49182 ; n49182_not
g90859 not n10878 ; n10878_not
g90860 not n43746 ; n43746_not
g90861 not n44277 ; n44277_not
g90862 not n32847 ; n32847_not
g90863 not n56229 ; n56229_not
g90864 not n47094 ; n47094_not
g90865 not n16287 ; n16287_not
g90866 not n32973 ; n32973_not
g90867 not n32838 ; n32838_not
g90868 not n54447 ; n54447_not
g90869 not n32829 ; n32829_not
g90870 not n16269 ; n16269_not
g90871 not n35790 ; n35790_not
g90872 not n37581 ; n37581_not
g90873 not n32991 ; n32991_not
g90874 not n50397 ; n50397_not
g90875 not n44871 ; n44871_not
g90876 not n32793 ; n32793_not
g90877 not n32784 ; n32784_not
g90878 not n49542 ; n49542_not
g90879 not n43089 ; n43089_not
g90880 not n50379 ; n50379_not
g90881 not n44268 ; n44268_not
g90882 not n49191 ; n49191_not
g90883 not n32982 ; n32982_not
g90884 not n34863 ; n34863_not
g90885 not n35781 ; n35781_not
g90886 not n14568 ; n14568_not
g90887 not n48660 ; n48660_not
g90888 not n49560 ; n49560_not
g90889 not n36627 ; n36627_not
g90890 not n37536 ; n37536_not
g90891 not n15675 ; n15675_not
g90892 not n11598 ; n11598_not
g90893 not n14559 ; n14559_not
g90894 not n50388 ; n50388_not
g90895 not n54456 ; n54456_not
g90896 not n47841 ; n47841_not
g90897 not n22983 ; n22983_not
g90898 not n22479 ; n22479_not
g90899 not n39075 ; n39075_not
g90900 not n52728 ; n52728_not
g90901 not n22398 ; n22398_not
g90902 not n22389 ; n22389_not
g90903 not n46635 ; n46635_not
g90904 not n27339 ; n27339_not
g90905 not n27348 ; n27348_not
g90906 not n39084 ; n39084_not
g90907 not n27357 ; n27357_not
g90908 not n27366 ; n27366_not
g90909 not n22992 ; n22992_not
g90910 not n27375 ; n27375_not
g90911 not n40992 ; n40992_not
g90912 not n51738 ; n51738_not
g90913 not n46617 ; n46617_not
g90914 not n22893 ; n22893_not
g90915 not n52476 ; n52476_not
g90916 not n38823 ; n38823_not
g90917 not n22596 ; n22596_not
g90918 not n27276 ; n27276_not
g90919 not n22587 ; n22587_not
g90920 not n22578 ; n22578_not
g90921 not n22929 ; n22929_not
g90922 not n22569 ; n22569_not
g90923 not n22938 ; n22938_not
g90924 not n38814 ; n38814_not
g90925 not n22956 ; n22956_not
g90926 not n27285 ; n27285_not
g90927 not n27294 ; n27294_not
g90928 not n22497 ; n22497_not
g90929 not n22974 ; n22974_not
g90930 not n22488 ; n22488_not
g90931 not n38805 ; n38805_not
g90932 not n51765 ; n51765_not
g90933 not n38742 ; n38742_not
g90934 not n40974 ; n40974_not
g90935 not n27465 ; n27465_not
g90936 not n38733 ; n38733_not
g90937 not n45483 ; n45483_not
g90938 not n27951 ; n27951_not
g90939 not n27474 ; n27474_not
g90940 not n38724 ; n38724_not
g90941 not n40965 ; n40965_not
g90942 not n40776 ; n40776_not
g90943 not n40398 ; n40398_not
g90944 not n52287 ; n52287_not
g90945 not n38715 ; n38715_not
g90946 not n27483 ; n27483_not
g90947 not n40956 ; n40956_not
g90948 not n40785 ; n40785_not
g90949 not n27384 ; n27384_not
g90950 not n27393 ; n27393_not
g90951 not n45474 ; n45474_not
g90952 not n38760 ; n38760_not
g90953 not n51747 ; n51747_not
g90954 not n27429 ; n27429_not
g90955 not n27438 ; n27438_not
g90956 not n40983 ; n40983_not
g90957 not n38751 ; n38751_not
g90958 not n40767 ; n40767_not
g90959 not n52296 ; n52296_not
g90960 not n22947 ; n22947_not
g90961 not n27447 ; n27447_not
g90962 not n27456 ; n27456_not
g90963 not n27960 ; n27960_not
g90964 not n38931 ; n38931_not
g90965 not n38922 ; n38922_not
g90966 not n22659 ; n22659_not
g90967 not n28167 ; n28167_not
g90968 not n22668 ; n22668_not
g90969 not n38913 ; n38913_not
g90970 not n22677 ; n22677_not
g90971 not n22686 ; n22686_not
g90972 not n38904 ; n38904_not
g90973 not n52377 ; n52377_not
g90974 not n28149 ; n28149_not
g90975 not n22695 ; n22695_not
g90976 not n52458 ; n52458_not
g90977 not n22749 ; n22749_not
g90978 not n28059 ; n28059_not
g90979 not n22758 ; n22758_not
g90980 not n28086 ; n28086_not
g90981 not n22767 ; n22767_not
g90982 not n27915 ; n27915_not
g90983 not n46581 ; n46581_not
g90984 not n52395 ; n52395_not
g90985 not n38940 ; n38940_not
g90986 not n51693 ; n51693_not
g90987 not n28194 ; n28194_not
g90988 not n52386 ; n52386_not
g90989 not n27249 ; n27249_not
g90990 not n22839 ; n22839_not
g90991 not n38841 ; n38841_not
g90992 not n22848 ; n22848_not
g90993 not n39057 ; n39057_not
g90994 not n40479 ; n40479_not
g90995 not n52467 ; n52467_not
g90996 not n22866 ; n22866_not
g90997 not n27258 ; n27258_not
g90998 not n38832 ; n38832_not
g90999 not n28068 ; n28068_not
g91000 not n27267 ; n27267_not
g91001 not n22884 ; n22884_not
g91002 not n39039 ; n39039_not
g91003 not n22776 ; n22776_not
g91004 not n52368 ; n52368_not
g91005 not n28095 ; n28095_not
g91006 not n22785 ; n22785_not
g91007 not n40497 ; n40497_not
g91008 not n46608 ; n46608_not
g91009 not n38850 ; n38850_not
g91010 not n52359 ; n52359_not
g91011 not n40488 ; n40488_not
g91012 not n45465 ; n45465_not
g91013 not n39129 ; n39129_not
g91014 not n23883 ; n23883_not
g91015 not n27726 ; n27726_not
g91016 not n27717 ; n27717_not
g91017 not n46518 ; n46518_not
g91018 not n23874 ; n23874_not
g91019 not n27708 ; n27708_not
g91020 not n23919 ; n23919_not
g91021 not n40299 ; n40299_not
g91022 not n26952 ; n26952_not
g91023 not n23928 ; n23928_not
g91024 not n52548 ; n52548_not
g91025 not n27690 ; n27690_not
g91026 not n51918 ; n51918_not
g91027 not n23937 ; n23937_not
g91028 not n26961 ; n26961_not
g91029 not n23946 ; n23946_not
g91030 not n23793 ; n23793_not
g91031 not n51873 ; n51873_not
g91032 not n40866 ; n40866_not
g91033 not n23829 ; n23829_not
g91034 not n23838 ; n23838_not
g91035 not n27762 ; n27762_not
g91036 not n40857 ; n40857_not
g91037 not n51882 ; n51882_not
g91038 not n26925 ; n26925_not
g91039 not n27753 ; n27753_not
g91040 not n23856 ; n23856_not
g91041 not n39138 ; n39138_not
g91042 not n46527 ; n46527_not
g91043 not n27744 ; n27744_not
g91044 not n27735 ; n27735_not
g91045 not n52566 ; n52566_not
g91046 not n27645 ; n27645_not
g91047 not n51945 ; n51945_not
g91048 not n23991 ; n23991_not
g91049 not n52179 ; n52179_not
g91050 not n40389 ; n40389_not
g91051 not n27636 ; n27636_not
g91052 not n51954 ; n51954_not
g91053 not n27681 ; n27681_not
g91054 not n26970 ; n26970_not
g91055 not n23955 ; n23955_not
g91056 not n51927 ; n51927_not
g91057 not n27672 ; n27672_not
g91058 not n23964 ; n23964_not
g91059 not n52197 ; n52197_not
g91060 not n23847 ; n23847_not
g91061 not n27663 ; n27663_not
g91062 not n23973 ; n23973_not
g91063 not n52557 ; n52557_not
g91064 not n51936 ; n51936_not
g91065 not n52188 ; n52188_not
g91066 not n45519 ; n45519_not
g91067 not n27654 ; n27654_not
g91068 not n40794 ; n40794_not
g91069 not n23982 ; n23982_not
g91070 not n27537 ; n27537_not
g91071 not n38670 ; n38670_not
g91072 not n40929 ; n40929_not
g91073 not n46590 ; n46590_not
g91074 not n27546 ; n27546_not
g91075 not n38661 ; n38661_not
g91076 not n27906 ; n27906_not
g91077 not n38652 ; n38652_not
g91078 not n51792 ; n51792_not
g91079 not n27555 ; n27555_not
g91080 not n27564 ; n27564_not
g91081 not n27573 ; n27573_not
g91082 not n27582 ; n27582_not
g91083 not n46572 ; n46572_not
g91084 not n27591 ; n27591_not
g91085 not n27609 ; n27609_not
g91086 not n27618 ; n27618_not
g91087 not n27870 ; n27870_not
g91088 not n38706 ; n38706_not
g91089 not n52278 ; n52278_not
g91090 not n27492 ; n27492_not
g91091 not n40947 ; n40947_not
g91092 not n45492 ; n45492_not
g91093 not n27933 ; n27933_not
g91094 not n27519 ; n27519_not
g91095 not n51783 ; n51783_not
g91096 not n40938 ; n40938_not
g91097 not n39147 ; n39147_not
g91098 not n52269 ; n52269_not
g91099 not n27528 ; n27528_not
g91100 not n22857 ; n22857_not
g91101 not n51837 ; n51837_not
g91102 not n23739 ; n23739_not
g91103 not n27825 ; n27825_not
g91104 not n40884 ; n40884_not
g91105 not n27816 ; n27816_not
g91106 not n46545 ; n46545_not
g91107 not n23748 ; n23748_not
g91108 not n23766 ; n23766_not
g91109 not n40875 ; n40875_not
g91110 not n23784 ; n23784_not
g91111 not n51855 ; n51855_not
g91112 not n39165 ; n39165_not
g91113 not n27627 ; n27627_not
g91114 not n27861 ; n27861_not
g91115 not n46563 ; n46563_not
g91116 not n23649 ; n23649_not
g91117 not n23658 ; n23658_not
g91118 not n39183 ; n39183_not
g91119 not n23676 ; n23676_not
g91120 not n39192 ; n39192_not
g91121 not n51828 ; n51828_not
g91122 not n23694 ; n23694_not
g91123 not n27843 ; n27843_not
g91124 not n40893 ; n40893_not
g91125 not n20778 ; n20778_not
g91126 not n52917 ; n52917_not
g91127 not n20859 ; n20859_not
g91128 not n51576 ; n51576_not
g91129 not n20868 ; n20868_not
g91130 not n38544 ; n38544_not
g91131 not n52926 ; n52926_not
g91132 not n20877 ; n20877_not
g91133 not n20886 ; n20886_not
g91134 not n52935 ; n52935_not
g91135 not n28491 ; n28491_not
g91136 not n20895 ; n20895_not
g91137 not n20787 ; n20787_not
g91138 not n28518 ; n28518_not
g91139 not n52890 ; n52890_not
g91140 not n53448 ; n53448_not
g91141 not n45447 ; n45447_not
g91142 not n28509 ; n28509_not
g91143 not n52908 ; n52908_not
g91144 not n38553 ; n38553_not
g91145 not n52962 ; n52962_not
g91146 not n50847 ; n50847_not
g91147 not n20967 ; n20967_not
g91148 not n51594 ; n51594_not
g91149 not n20976 ; n20976_not
g91150 not n52971 ; n52971_not
g91151 not n38535 ; n38535_not
g91152 not n20985 ; n20985_not
g91153 not n41298 ; n41298_not
g91154 not n52980 ; n52980_not
g91155 not n28473 ; n28473_not
g91156 not n20994 ; n20994_not
g91157 not n52944 ; n52944_not
g91158 not n20688 ; n20688_not
g91159 not n20679 ; n20679_not
g91160 not n51585 ; n51585_not
g91161 not n52953 ; n52953_not
g91162 not n28482 ; n28482_not
g91163 not n20949 ; n20949_not
g91164 not n20958 ; n20958_not
g91165 not n52764 ; n52764_not
g91166 not n28554 ; n28554_not
g91167 not n52773 ; n52773_not
g91168 not n52782 ; n52782_not
g91169 not n19833 ; n19833_not
g91170 not n46473 ; n46473_not
g91171 not n52791 ; n52791_not
g91172 not n19824 ; n19824_not
g91173 not n52809 ; n52809_not
g91174 not n53493 ; n53493_not
g91175 not n19815 ; n19815_not
g91176 not n52818 ; n52818_not
g91177 not n19905 ; n19905_not
g91178 not n53529 ; n53529_not
g91179 not n52755 ; n52755_not
g91180 not n53556 ; n53556_not
g91181 not n52746 ; n52746_not
g91182 not n38580 ; n38580_not
g91183 not n53547 ; n53547_not
g91184 not n51549 ; n51549_not
g91185 not n28563 ; n28563_not
g91186 not n52737 ; n52737_not
g91187 not n19860 ; n19860_not
g91188 not n52872 ; n52872_not
g91189 not n41397 ; n41397_not
g91190 not n28545 ; n28545_not
g91191 not n41388 ; n41388_not
g91192 not n20589 ; n20589_not
g91193 not n28536 ; n28536_not
g91194 not n51567 ; n51567_not
g91195 not n52881 ; n52881_not
g91196 not n20697 ; n20697_not
g91197 not n28527 ; n28527_not
g91198 not n20769 ; n20769_not
g91199 not n51558 ; n51558_not
g91200 not n52827 ; n52827_not
g91201 not n45438 ; n45438_not
g91202 not n46482 ; n46482_not
g91203 not n52836 ; n52836_not
g91204 not n53475 ; n53475_not
g91205 not n52845 ; n52845_not
g91206 not n52854 ; n52854_not
g91207 not n53466 ; n53466_not
g91208 not n46491 ; n46491_not
g91209 not n52863 ; n52863_not
g91210 not n19770 ; n19770_not
g91211 not n19752 ; n19752_not
g91212 not n28365 ; n28365_not
g91213 not n21795 ; n21795_not
g91214 not n53187 ; n53187_not
g91215 not n53196 ; n53196_not
g91216 not n28347 ; n28347_not
g91217 not n21849 ; n21849_not
g91218 not n28338 ; n28338_not
g91219 not n21858 ; n21858_not
g91220 not n21867 ; n21867_not
g91221 not n38490 ; n38490_not
g91222 not n21876 ; n21876_not
g91223 not n53268 ; n53268_not
g91224 not n21885 ; n21885_not
g91225 not n21894 ; n21894_not
g91226 not n53295 ; n53295_not
g91227 not n53169 ; n53169_not
g91228 not n28383 ; n28383_not
g91229 not n38508 ; n38508_not
g91230 not n21759 ; n21759_not
g91231 not n21399 ; n21399_not
g91232 not n21768 ; n21768_not
g91233 not n41199 ; n41199_not
g91234 not n53178 ; n53178_not
g91235 not n28374 ; n28374_not
g91236 not n21777 ; n21777_not
g91237 not n53286 ; n53286_not
g91238 not n21786 ; n21786_not
g91239 not n40578 ; n40578_not
g91240 not n28275 ; n28275_not
g91241 not n40569 ; n40569_not
g91242 not n28266 ; n28266_not
g91243 not n51675 ; n51675_not
g91244 not n38463 ; n38463_not
g91245 not n45456 ; n45456_not
g91246 not n40686 ; n40686_not
g91247 not n28239 ; n28239_not
g91248 not n40695 ; n40695_not
g91249 not n21939 ; n21939_not
g91250 not n40596 ; n40596_not
g91251 not n21948 ; n21948_not
g91252 not n51648 ; n51648_not
g91253 not n28293 ; n28293_not
g91254 not n21957 ; n21957_not
g91255 not n21966 ; n21966_not
g91256 not n51657 ; n51657_not
g91257 not n40587 ; n40587_not
g91258 not n21975 ; n21975_not
g91259 not n28284 ; n28284_not
g91260 not n21984 ; n21984_not
g91261 not n21993 ; n21993_not
g91262 not n40677 ; n40677_not
g91263 not n53358 ; n53358_not
g91264 not n28455 ; n28455_not
g91265 not n28446 ; n28446_not
g91266 not n53385 ; n53385_not
g91267 not n53376 ; n53376_not
g91268 not n50838 ; n50838_not
g91269 not n20598 ; n20598_not
g91270 not n28464 ; n28464_not
g91271 not n28437 ; n28437_not
g91272 not n53088 ; n53088_not
g91273 not n53097 ; n53097_not
g91274 not n28428 ; n28428_not
g91275 not n21579 ; n21579_not
g91276 not n21588 ; n21588_not
g91277 not n21498 ; n21498_not
g91278 not n28419 ; n28419_not
g91279 not n21597 ; n21597_not
g91280 not n21489 ; n21489_not
g91281 not n21669 ; n21669_not
g91282 not n21678 ; n21678_not
g91283 not n21687 ; n21687_not
g91284 not n46536 ; n46536_not
g91285 not n21696 ; n21696_not
g91286 not n28392 ; n28392_not
g91287 not n53079 ; n53079_not
g91288 not n27834 ; n27834_not
g91289 not n26187 ; n26187_not
g91290 not n25863 ; n25863_not
g91291 not n26682 ; n26682_not
g91292 not n39750 ; n39750_not
g91293 not n25854 ; n25854_not
g91294 not n45816 ; n45816_not
g91295 not n45663 ; n45663_not
g91296 not n26673 ; n26673_not
g91297 not n52485 ; n52485_not
g91298 not n26196 ; n26196_not
g91299 not n25845 ; n25845_not
g91300 not n26664 ; n26664_not
g91301 not n25089 ; n25089_not
g91302 not n25836 ; n25836_not
g91303 not n26655 ; n26655_not
g91304 not n25098 ; n25098_not
g91305 not n25827 ; n25827_not
g91306 not n26727 ; n26727_not
g91307 not n45636 ; n45636_not
g91308 not n39714 ; n39714_not
g91309 not n26718 ; n26718_not
g91310 not n24972 ; n24972_not
g91311 not n24981 ; n24981_not
g91312 not n25890 ; n25890_not
g91313 not n39723 ; n39723_not
g91314 not n26709 ; n26709_not
g91315 not n45645 ; n45645_not
g91316 not n24990 ; n24990_not
g91317 not n39732 ; n39732_not
g91318 not n25881 ; n25881_not
g91319 not n25359 ; n25359_not
g91320 not n45654 ; n45654_not
g91321 not n25872 ; n25872_not
g91322 not n26691 ; n26691_not
g91323 not n25197 ; n25197_not
g91324 not n25773 ; n25773_not
g91325 not n26592 ; n26592_not
g91326 not n39813 ; n39813_not
g91327 not n26079 ; n26079_not
g91328 not n25764 ; n25764_not
g91329 not n26583 ; n26583_not
g91330 not n26097 ; n26097_not
g91331 not n25980 ; n25980_not
g91332 not n25971 ; n25971_not
g91333 not n25962 ; n25962_not
g91334 not n25953 ; n25953_not
g91335 not n25944 ; n25944_not
g91336 not n45825 ; n45825_not
g91337 not n45690 ; n45690_not
g91338 not n26646 ; n26646_not
g91339 not n25296 ; n25296_not
g91340 not n45834 ; n45834_not
g91341 not n25818 ; n25818_not
g91342 not n45708 ; n45708_not
g91343 not n26637 ; n26637_not
g91344 not n25809 ; n25809_not
g91345 not n26628 ; n26628_not
g91346 not n26619 ; n26619_not
g91347 not n25791 ; n25791_not
g91348 not n25269 ; n25269_not
g91349 not n25179 ; n25179_not
g91350 not n25782 ; n25782_not
g91351 not n39804 ; n39804_not
g91352 not n25188 ; n25188_not
g91353 not n24783 ; n24783_not
g91354 not n39624 ; n39624_not
g91355 not n26817 ; n26817_not
g91356 not n25476 ; n25476_not
g91357 not n24792 ; n24792_not
g91358 not n39633 ; n39633_not
g91359 not n26808 ; n26808_not
g91360 not n24819 ; n24819_not
g91361 not n26790 ; n26790_not
g91362 not n24828 ; n24828_not
g91363 not n39651 ; n39651_not
g91364 not n45771 ; n45771_not
g91365 not n24837 ; n24837_not
g91366 not n26781 ; n26781_not
g91367 not n25449 ; n25449_not
g91368 not n26853 ; n26853_not
g91369 not n24738 ; n24738_not
g91370 not n39606 ; n39606_not
g91371 not n52593 ; n52593_not
g91372 not n24747 ; n24747_not
g91373 not n26844 ; n26844_not
g91374 not n26835 ; n26835_not
g91375 not n24756 ; n24756_not
g91376 not n25494 ; n25494_not
g91377 not n45591 ; n45591_not
g91378 not n24765 ; n24765_not
g91379 not n26826 ; n26826_not
g91380 not n25485 ; n25485_not
g91381 not n24774 ; n24774_not
g91382 not n52575 ; n52575_not
g91383 not n24909 ; n24909_not
g91384 not n45618 ; n45618_not
g91385 not n24918 ; n24918_not
g91386 not n26754 ; n26754_not
g91387 not n24927 ; n24927_not
g91388 not n25926 ; n25926_not
g91389 not n25395 ; n25395_not
g91390 not n24936 ; n24936_not
g91391 not n26745 ; n26745_not
g91392 not n45627 ; n45627_not
g91393 not n24945 ; n24945_not
g91394 not n25917 ; n25917_not
g91395 not n26736 ; n26736_not
g91396 not n25386 ; n25386_not
g91397 not n24954 ; n24954_not
g91398 not n25908 ; n25908_not
g91399 not n24963 ; n24963_not
g91400 not n24846 ; n24846_not
g91401 not n24855 ; n24855_not
g91402 not n26772 ; n26772_not
g91403 not n24864 ; n24864_not
g91404 not n39741 ; n39741_not
g91405 not n45609 ; n45609_not
g91406 not n24873 ; n24873_not
g91407 not n45780 ; n45780_not
g91408 not n24882 ; n24882_not
g91409 not n24891 ; n24891_not
g91410 not n26763 ; n26763_not
g91411 not n25935 ; n25935_not
g91412 not n25584 ; n25584_not
g91413 not n25575 ; n25575_not
g91414 not n25692 ; n25692_not
g91415 not n25566 ; n25566_not
g91416 not n26349 ; n26349_not
g91417 not n25557 ; n25557_not
g91418 not n25548 ; n25548_not
g91419 not n26286 ; n26286_not
g91420 not n26367 ; n26367_not
g91421 not n45915 ; n45915_not
g91422 not n25683 ; n25683_not
g91423 not n25674 ; n25674_not
g91424 not n26277 ; n26277_not
g91425 not n25665 ; n25665_not
g91426 not n25656 ; n25656_not
g91427 not n25647 ; n25647_not
g91428 not n25638 ; n25638_not
g91429 not n25629 ; n25629_not
g91430 not n45906 ; n45906_not
g91431 not n25593 ; n25593_not
g91432 not n39642 ; n39642_not
g91433 not n39930 ; n39930_not
g91434 not n39903 ; n39903_not
g91435 not n26475 ; n26475_not
g91436 not n26439 ; n26439_not
g91437 not n26448 ; n26448_not
g91438 not n39921 ; n39921_not
g91439 not n26457 ; n26457_not
g91440 not n26466 ; n26466_not
g91441 not n39912 ; n39912_not
g91442 not n26295 ; n26295_not
g91443 not n45924 ; n45924_not
g91444 not n26385 ; n26385_not
g91445 not n45843 ; n45843_not
g91446 not n26493 ; n26493_not
g91447 not n26394 ; n26394_not
g91448 not n51666 ; n51666_not
g91449 not n45861 ; n45861_not
g91450 not n26484 ; n26484_not
g91451 not n45870 ; n45870_not
g91452 not n25746 ; n25746_not
g91453 not n39831 ; n39831_not
g91454 not n39534 ; n39534_not
g91455 not n26565 ; n26565_not
g91456 not n25737 ; n25737_not
g91457 not n26556 ; n26556_not
g91458 not n39822 ; n39822_not
g91459 not n25755 ; n25755_not
g91460 not n26574 ; n26574_not
g91461 not n26169 ; n26169_not
g91462 not n45735 ; n45735_not
g91463 not n25719 ; n25719_not
g91464 not n25728 ; n25728_not
g91465 not n26259 ; n26259_not
g91466 not n26538 ; n26538_not
g91467 not n45753 ; n45753_not
g91468 not n26529 ; n26529_not
g91469 not n39543 ; n39543_not
g91470 not n39840 ; n39840_not
g91471 not n39552 ; n39552_not
g91472 not n45726 ; n45726_not
g91473 not n26547 ; n26547_not
g91474 not n24369 ; n24369_not
g91475 not n46392 ; n46392_not
g91476 not n24378 ; n24378_not
g91477 not n24387 ; n24387_not
g91478 not n52647 ; n52647_not
g91479 not n46383 ; n46383_not
g91480 not n24468 ; n24468_not
g91481 not n27177 ; n27177_not
g91482 not n52656 ; n52656_not
g91483 not n24486 ; n24486_not
g91484 not n24495 ; n24495_not
g91485 not n24288 ; n24288_not
g91486 not n23667 ; n23667_not
g91487 not n24297 ; n24297_not
g91488 not n27096 ; n27096_not
g91489 not n52638 ; n52638_not
g91490 not n51846 ; n51846_not
g91491 not n39048 ; n39048_not
g91492 not n24675 ; n24675_not
g91493 not n24693 ; n24693_not
g91494 not n23892 ; n23892_not
g91495 not n51990 ; n51990_not
g91496 not n51981 ; n51981_not
g91497 not n27186 ; n27186_not
g91498 not n24729 ; n24729_not
g91499 not n24684 ; n24684_not
g91500 not n24558 ; n24558_not
g91501 not n46365 ; n46365_not
g91502 not n46374 ; n46374_not
g91503 not n24576 ; n24576_not
g91504 not n24585 ; n24585_not
g91505 not n27195 ; n27195_not
g91506 not n24648 ; n24648_not
g91507 not n24666 ; n24666_not
g91508 not n24099 ; n24099_not
g91509 not n39093 ; n39093_not
g91510 not n23757 ; n23757_not
g91511 not n51891 ; n51891_not
g91512 not n51963 ; n51963_not
g91513 not n40749 ; n40749_not
g91514 not n51972 ; n51972_not
g91515 not n46437 ; n46437_not
g91516 not n46428 ; n46428_not
g91517 not n40659 ; n40659_not
g91518 not n27087 ; n27087_not
g91519 not n24279 ; n24279_not
g91520 not n46455 ; n46455_not
g91521 not n24189 ; n24189_not
g91522 not n52098 ; n52098_not
g91523 not n45528 ; n45528_not
g91524 not n24198 ; n24198_not
g91525 not n52089 ; n52089_not
g91526 not n45564 ; n45564_not
g91527 not n39525 ; n39525_not
g91528 not n52665 ; n52665_not
g91529 not n24459 ; n24459_not
g91530 not n26862 ; n26862_not
g91531 not n24549 ; n24549_not
g91532 not n52692 ; n52692_not
g91533 not n52683 ; n52683_not
g91534 not n45744 ; n45744_not
g91535 not n25458 ; n25458_not
g91536 not n45582 ; n45582_not
g91537 not n51756 ; n51756_not
g91538 not n26880 ; n26880_not
g91539 not n26871 ; n26871_not
g91540 not n25278 ; n25278_not
g91541 not n45573 ; n45573_not
g91542 not n25368 ; n25368_not
g91543 not n26934 ; n26934_not
g91544 not n39561 ; n39561_not
g91545 not n24639 ; n24639_not
g91546 not n45537 ; n45537_not
g91547 not n27159 ; n27159_not
g91548 not n52719 ; n52719_not
g91549 not n45555 ; n45555_not
g91550 not n45546 ; n45546_not
g91551 not n27069 ; n27069_not
g91552 not n24594 ; n24594_not
g91553 not n41928 ; n41928_not
g91554 not n29418 ; n29418_not
g91555 not n18942 ; n18942_not
g91556 not n18375 ; n18375_not
g91557 not n29364 ; n29364_not
g91558 not n18951 ; n18951_not
g91559 not n29382 ; n29382_not
g91560 not n18960 ; n18960_not
g91561 not n51189 ; n51189_not
g91562 not n38472 ; n38472_not
g91563 not n29373 ; n29373_not
g91564 not n51198 ; n51198_not
g91565 not n29454 ; n29454_not
g91566 not n54276 ; n54276_not
g91567 not n41955 ; n41955_not
g91568 not n29445 ; n29445_not
g91569 not n18906 ; n18906_not
g91570 not n38445 ; n38445_not
g91571 not n29436 ; n29436_not
g91572 not n18915 ; n18915_not
g91573 not n18393 ; n18393_not
g91574 not n29355 ; n29355_not
g91575 not n18924 ; n18924_not
g91576 not n18384 ; n18384_not
g91577 not n54258 ; n54258_not
g91578 not n41937 ; n41937_not
g91579 not n38454 ; n38454_not
g91580 not n18933 ; n18933_not
g91581 not n29427 ; n29427_not
g91582 not n29238 ; n29238_not
g91583 not n19095 ; n19095_not
g91584 not n38517 ; n38517_not
g91585 not n29265 ; n29265_not
g91586 not n29274 ; n29274_not
g91587 not n41865 ; n41865_not
g91588 not n29229 ; n29229_not
g91589 not n19158 ; n19158_not
g91590 not n29247 ; n29247_not
g91591 not n19167 ; n19167_not
g91592 not n29157 ; n29157_not
g91593 not n29166 ; n29166_not
g91594 not n45366 ; n45366_not
g91595 not n18348 ; n18348_not
g91596 not n18339 ; n18339_not
g91597 not n41892 ; n41892_not
g91598 not n45357 ; n45357_not
g91599 not n29337 ; n29337_not
g91600 not n41883 ; n41883_not
g91601 not n19068 ; n19068_not
g91602 not n19077 ; n19077_not
g91603 not n54168 ; n54168_not
g91604 not n29472 ; n29472_not
g91605 not n29571 ; n29571_not
g91606 not n18780 ; n18780_not
g91607 not n29463 ; n29463_not
g91608 not n18465 ; n18465_not
g91609 not n29562 ; n29562_not
g91610 not n38391 ; n38391_not
g91611 not n54348 ; n54348_not
g91612 not n51099 ; n51099_not
g91613 not n29553 ; n29553_not
g91614 not n29544 ; n29544_not
g91615 not n29535 ; n29535_not
g91616 not n18807 ; n18807_not
g91617 not n29634 ; n29634_not
g91618 not n18753 ; n18753_not
g91619 not n29625 ; n29625_not
g91620 not n18483 ; n18483_not
g91621 not n38373 ; n38373_not
g91622 not n45339 ; n45339_not
g91623 not n18762 ; n18762_not
g91624 not n18474 ; n18474_not
g91625 not n29607 ; n29607_not
g91626 not n54366 ; n54366_not
g91627 not n18771 ; n18771_not
g91628 not n38382 ; n38382_not
g91629 not n29580 ; n29580_not
g91630 not n41982 ; n41982_not
g91631 not n18852 ; n18852_not
g91632 not n45195 ; n45195_not
g91633 not n29481 ; n29481_not
g91634 not n41973 ; n41973_not
g91635 not n18861 ; n18861_not
g91636 not n38427 ; n38427_not
g91637 not n45348 ; n45348_not
g91638 not n18870 ; n18870_not
g91639 not n47085 ; n47085_not
g91640 not n54285 ; n54285_not
g91641 not n38436 ; n38436_not
g91642 not n18816 ; n18816_not
g91643 not n29526 ; n29526_not
g91644 not n29508 ; n29508_not
g91645 not n18825 ; n18825_not
g91646 not n38409 ; n38409_not
g91647 not n18834 ; n18834_not
g91648 not n29409 ; n29409_not
g91649 not n18438 ; n18438_not
g91650 not n18843 ; n18843_not
g91651 not n18429 ; n18429_not
g91652 not n38418 ; n38418_not
g91653 not n51396 ; n51396_not
g91654 not n19437 ; n19437_not
g91655 not n18744 ; n18744_not
g91656 not n28833 ; n28833_not
g91657 not n19446 ; n19446_not
g91658 not n38625 ; n38625_not
g91659 not n41748 ; n41748_not
g91660 not n19455 ; n19455_not
g91661 not n28824 ; n28824_not
g91662 not n19464 ; n19464_not
g91663 not n38634 ; n38634_not
g91664 not n19383 ; n19383_not
g91665 not n51378 ; n51378_not
g91666 not n18690 ; n18690_not
g91667 not n19248 ; n19248_not
g91668 not n28860 ; n28860_not
g91669 not n19392 ; n19392_not
g91670 not n41766 ; n41766_not
g91671 not n28851 ; n28851_not
g91672 not n51387 ; n51387_not
g91673 not n18708 ; n18708_not
g91674 not n18717 ; n18717_not
g91675 not n19419 ; n19419_not
g91676 not n18726 ; n18726_not
g91677 not n41757 ; n41757_not
g91678 not n28842 ; n28842_not
g91679 not n19428 ; n19428_not
g91680 not n18735 ; n18735_not
g91681 not n19509 ; n19509_not
g91682 not n50928 ; n50928_not
g91683 not n19518 ; n19518_not
g91684 not n53952 ; n53952_not
g91685 not n19176 ; n19176_not
g91686 not n19527 ; n19527_not
g91687 not n28752 ; n28752_not
g91688 not n19536 ; n19536_not
g91689 not n53943 ; n53943_not
g91690 not n28743 ; n28743_not
g91691 not n19545 ; n19545_not
g91692 not n28176 ; n28176_not
g91693 not n41739 ; n41739_not
g91694 not n28815 ; n28815_not
g91695 not n19473 ; n19473_not
g91696 not n28806 ; n28806_not
g91697 not n45384 ; n45384_not
g91698 not n19482 ; n19482_not
g91699 not n50937 ; n50937_not
g91700 not n19491 ; n19491_not
g91701 not n53970 ; n53970_not
g91702 not n28770 ; n28770_not
g91703 not n53961 ; n53961_not
g91704 not n28761 ; n28761_not
g91705 not n29067 ; n29067_not
g91706 not n29085 ; n29085_not
g91707 not n19257 ; n19257_not
g91708 not n54069 ; n54069_not
g91709 not n29076 ; n29076_not
g91710 not n19275 ; n19275_not
g91711 not n51279 ; n51279_not
g91712 not n51288 ; n51288_not
g91713 not n51297 ; n51297_not
g91714 not n19293 ; n19293_not
g91715 not n18609 ; n18609_not
g91716 not n19185 ; n19185_not
g91717 not n29184 ; n29184_not
g91718 not n29175 ; n29175_not
g91719 not n29148 ; n29148_not
g91720 not n54078 ; n54078_not
g91721 not n38562 ; n38562_not
g91722 not n18645 ; n18645_not
g91723 not n50982 ; n50982_not
g91724 not n19347 ; n19347_not
g91725 not n41784 ; n41784_not
g91726 not n18654 ; n18654_not
g91727 not n38607 ; n38607_not
g91728 not n19356 ; n19356_not
g91729 not n18663 ; n18663_not
g91730 not n50973 ; n50973_not
g91731 not n19266 ; n19266_not
g91732 not n19365 ; n19365_not
g91733 not n18672 ; n18672_not
g91734 not n41775 ; n41775_not
g91735 not n51369 ; n51369_not
g91736 not n19374 ; n19374_not
g91737 not n18681 ; n18681_not
g91738 not n50964 ; n50964_not
g91739 not n28950 ; n28950_not
g91740 not n28941 ; n28941_not
g91741 not n53259 ; n53259_not
g91742 not n18618 ; n18618_not
g91743 not n18627 ; n18627_not
g91744 not n28905 ; n28905_not
g91745 not n41793 ; n41793_not
g91746 not n28914 ; n28914_not
g91747 not n19329 ; n19329_not
g91748 not n18636 ; n18636_not
g91749 not n19338 ; n19338_not
g91750 not n45375 ; n45375_not
g91751 not n18249 ; n18249_not
g91752 not n38193 ; n38193_not
g91753 not n18258 ; n18258_not
g91754 not n50748 ; n50748_not
g91755 not n18267 ; n18267_not
g91756 not n50757 ; n50757_not
g91757 not n29913 ; n29913_not
g91758 not n18276 ; n18276_not
g91759 not n50766 ; n50766_not
g91760 not n29922 ; n29922_not
g91761 not n18195 ; n18195_not
g91762 not n30588 ; n30588_not
g91763 not n30579 ; n30579_not
g91764 not n38175 ; n38175_not
g91765 not n30498 ; n30498_not
g91766 not n38184 ; n38184_not
g91767 not n30399 ; n30399_not
g91768 not n17673 ; n17673_not
g91769 not n50739 ; n50739_not
g91770 not n29940 ; n29940_not
g91771 not n50793 ; n50793_not
g91772 not n54294 ; n54294_not
g91773 not n50784 ; n50784_not
g91774 not n50856 ; n50856_not
g91775 not n38238 ; n38238_not
g91776 not n50775 ; n50775_not
g91777 not n18285 ; n18285_not
g91778 not n29931 ; n29931_not
g91779 not n38094 ; n38094_not
g91780 not n18294 ; n18294_not
g91781 not n18357 ; n18357_not
g91782 not n38229 ; n38229_not
g91783 not n18069 ; n18069_not
g91784 not n37653 ; n37653_not
g91785 not n17763 ; n17763_not
g91786 not n18078 ; n18078_not
g91787 not n18087 ; n18087_not
g91788 not n18096 ; n18096_not
g91789 not n41856 ; n41856_not
g91790 not n47265 ; n47265_not
g91791 not n45285 ; n45285_not
g91792 not n17718 ; n17718_not
g91793 not n30669 ; n30669_not
g91794 not n18159 ; n18159_not
g91795 not n54249 ; n54249_not
g91796 not n18168 ; n18168_not
g91797 not n18177 ; n18177_not
g91798 not n38166 ; n38166_not
g91799 not n18186 ; n18186_not
g91800 not n30597 ; n30597_not
g91801 not n38148 ; n38148_not
g91802 not n45294 ; n45294_not
g91803 not n38157 ; n38157_not
g91804 not n29706 ; n29706_not
g91805 not n29751 ; n29751_not
g91806 not n29715 ; n29715_not
g91807 not n38328 ; n38328_not
g91808 not n29742 ; n29742_not
g91809 not n29724 ; n29724_not
g91810 not n29733 ; n29733_not
g91811 not n50991 ; n50991_not
g91812 not n54339 ; n54339_not
g91813 not n29652 ; n29652_not
g91814 not n29661 ; n29661_not
g91815 not n29670 ; n29670_not
g91816 not n18555 ; n18555_not
g91817 not n38319 ; n38319_not
g91818 not n41991 ; n41991_not
g91819 not n38355 ; n38355_not
g91820 not n29643 ; n29643_not
g91821 not n38364 ; n38364_not
g91822 not n18528 ; n18528_not
g91823 not n38337 ; n38337_not
g91824 not n18519 ; n18519_not
g91825 not n38346 ; n38346_not
g91826 not n38265 ; n38265_not
g91827 not n38274 ; n38274_not
g91828 not n18492 ; n18492_not
g91829 not n47175 ; n47175_not
g91830 not n29760 ; n29760_not
g91831 not n38247 ; n38247_not
g91832 not n50874 ; n50874_not
g91833 not n41946 ; n41946_not
g91834 not n38256 ; n38256_not
g91835 not n18447 ; n18447_not
g91836 not n29904 ; n29904_not
g91837 not n50883 ; n50883_not
g91838 not n18573 ; n18573_not
g91839 not n29814 ; n29814_not
g91840 not n29805 ; n29805_not
g91841 not n18564 ; n18564_not
g91842 not n18537 ; n18537_not
g91843 not n38283 ; n38283_not
g91844 not n50919 ; n50919_not
g91845 not n38049 ; n38049_not
g91846 not n38292 ; n38292_not
g91847 not n50946 ; n50946_not
g91848 not n53664 ; n53664_not
g91849 not n53844 ; n53844_not
g91850 not n19086 ; n19086_not
g91851 not n53853 ; n53853_not
g91852 not n53655 ; n53655_not
g91853 not n19680 ; n19680_not
g91854 not n53862 ; n53862_not
g91855 not n41649 ; n41649_not
g91856 not n19671 ; n19671_not
g91857 not n28707 ; n28707_not
g91858 not n53871 ; n53871_not
g91859 not n53682 ; n53682_not
g91860 not n53826 ; n53826_not
g91861 not n19743 ; n19743_not
g91862 not n19734 ; n19734_not
g91863 not n19950 ; n19950_not
g91864 not n51468 ; n51468_not
g91865 not n19725 ; n19725_not
g91866 not n53835 ; n53835_not
g91867 not n19716 ; n19716_not
g91868 not n53673 ; n53673_not
g91869 not n28617 ; n28617_not
g91870 not n19707 ; n19707_not
g91871 not n27924 ; n27924_not
g91872 not n19626 ; n19626_not
g91873 not n19617 ; n19617_not
g91874 not n41496 ; n41496_not
g91875 not n53628 ; n53628_not
g91876 not n41676 ; n41676_not
g91877 not n19608 ; n19608_not
g91878 not n53619 ; n53619_not
g91879 not n28590 ; n28590_not
g91880 not n53907 ; n53907_not
g91881 not n53646 ; n53646_not
g91882 not n19662 ; n19662_not
g91883 not n53880 ; n53880_not
g91884 not n53484 ; n53484_not
g91885 not n41658 ; n41658_not
g91886 not n28608 ; n28608_not
g91887 not n19653 ; n19653_not
g91888 not n53637 ; n53637_not
g91889 not n19644 ; n19644_not
g91890 not n53349 ; n53349_not
g91891 not n28716 ; n28716_not
g91892 not n19635 ; n19635_not
g91893 not n41667 ; n41667_not
g91894 not n51459 ; n51459_not
g91895 not n41586 ; n41586_not
g91896 not n19554 ; n19554_not
g91897 not n53439 ; n53439_not
g91898 not n53763 ; n53763_not
g91899 not n41559 ; n41559_not
g91900 not n50892 ; n50892_not
g91901 not n51495 ; n51495_not
g91902 not n53718 ; n53718_not
g91903 not n53772 ; n53772_not
g91904 not n41595 ; n41595_not
g91905 not n19590 ; n19590_not
g91906 not n53745 ; n53745_not
g91907 not n19581 ; n19581_not
g91908 not n28653 ; n28653_not
g91909 not n41577 ; n41577_not
g91910 not n41568 ; n41568_not
g91911 not n19842 ; n19842_not
g91912 not n53736 ; n53736_not
g91913 not n19572 ; n19572_not
g91914 not n53754 ; n53754_not
g91915 not n19563 ; n19563_not
g91916 not n53727 ; n53727_not
g91917 not n28662 ; n28662_not
g91918 not n19932 ; n19932_not
g91919 not n28635 ; n28635_not
g91920 not n53394 ; n53394_not
g91921 not n53808 ; n53808_not
g91922 not n51477 ; n51477_not
g91923 not n53691 ; n53691_not
g91924 not n53817 ; n53817_not
g91925 not n28626 ; n28626_not
g91926 not n19761 ; n19761_not
g91927 not n28671 ; n28671_not
g91928 not n28644 ; n28644_not
g91929 not n53781 ; n53781_not
g91930 not n19914 ; n19914_not
g91931 not n53709 ; n53709_not
g91932 not n51486 ; n51486_not
g91933 not n28680 ; n28680_not
g91934 not n53790 ; n53790_not
g91935 not n46446 ; n46446_not
g91936 not n41694 ; n41694_not
g91937 not n28581 ; n28581_not
g91938 not n53592 ; n53592_not
g91939 not n28734 ; n28734_not
g91940 not n53583 ; n53583_not
g91941 not n38643 ; n38643_not
g91942 not n41478 ; n41478_not
g91943 not n28572 ; n28572_not
g91944 not n53925 ; n53925_not
g91945 not n45429 ; n45429_not
g91946 not n41469 ; n41469_not
g91947 not n53574 ; n53574_not
g91948 not n41685 ; n41685_not
g91949 not n19923 ; n19923_not
g91950 not n28725 ; n28725_not
g91951 not n41487 ; n41487_not
g91952 not n53934 ; n53934_not
g91953 not n53916 ; n53916_not
g91954 not n45393 ; n45393_not
g91955 not n53565 ; n53565_not
g91956 not n28248 ; n28248_not
g91957 not n51928 ; n51928_not
g91958 not n57337 ; n57337_not
g91959 not n52198 ; n52198_not
g91960 not n54394 ; n54394_not
g91961 not n46843 ; n46843_not
g91962 not n48643 ; n48643_not
g91963 not n52558 ; n52558_not
g91964 not n48607 ; n48607_not
g91965 not n51919 ; n51919_not
g91966 not n47392 ; n47392_not
g91967 not n46924 ; n46924_not
g91968 not n44962 ; n44962_not
g91969 not n45826 ; n45826_not
g91970 not n57346 ; n57346_not
g91971 not n46636 ; n46636_not
g91972 not n56851 ; n56851_not
g91973 not n53692 ; n53692_not
g91974 not n54466 ; n54466_not
g91975 not n56257 ; n56257_not
g91976 not n48814 ; n48814_not
g91977 not n47356 ; n47356_not
g91978 not n50848 ; n50848_not
g91979 not n47824 ; n47824_not
g91980 not n45934 ; n45934_not
g91981 not n47158 ; n47158_not
g91982 not n46195 ; n46195_not
g91983 not n47257 ; n47257_not
g91984 not n47743 ; n47743_not
g91985 not n49156 ; n49156_not
g91986 not n56248 ; n56248_not
g91987 not n54556 ; n54556_not
g91988 not n44791 ; n44791_not
g91989 not n50938 ; n50938_not
g91990 not n57355 ; n57355_not
g91991 not n56905 ; n56905_not
g91992 not n49174 ; n49174_not
g91993 not n56329 ; n56329_not
g91994 not n49093 ; n49093_not
g91995 not n46942 ; n46942_not
g91996 not n46753 ; n46753_not
g91997 not n44881 ; n44881_not
g91998 not n50956 ; n50956_not
g91999 not n53575 ; n53575_not
g92000 not n54493 ; n54493_not
g92001 not n45853 ; n45853_not
g92002 not n44872 ; n44872_not
g92003 not n53539 ; n53539_not
g92004 not n46456 ; n46456_not
g92005 not n52189 ; n52189_not
g92006 not n56239 ; n56239_not
g92007 not n44827 ; n44827_not
g92008 not n44494 ; n44494_not
g92009 not n49165 ; n49165_not
g92010 not n57265 ; n57265_not
g92011 not n44809 ; n44809_not
g92012 not n47770 ; n47770_not
g92013 not n52567 ; n52567_not
g92014 not n50929 ; n50929_not
g92015 not n53674 ; n53674_not
g92016 not n56284 ; n56284_not
g92017 not n44980 ; n44980_not
g92018 not n49129 ; n49129_not
g92019 not n45790 ; n45790_not
g92020 not n56275 ; n56275_not
g92021 not n47752 ; n47752_not
g92022 not n47374 ; n47374_not
g92023 not n44674 ; n44674_not
g92024 not n57274 ; n57274_not
g92025 not n52279 ; n52279_not
g92026 not n51577 ; n51577_not
g92027 not n53683 ; n53683_not
g92028 not n47185 ; n47185_not
g92029 not n50884 ; n50884_not
g92030 not n56293 ; n56293_not
g92031 not n46906 ; n46906_not
g92032 not n47365 ; n47365_not
g92033 not n50857 ; n50857_not
g92034 not n54547 ; n54547_not
g92035 not n46933 ; n46933_not
g92036 not n50893 ; n50893_not
g92037 not n55195 ; n55195_not
g92038 not n57283 ; n57283_not
g92039 not n46159 ; n46159_not
g92040 not n47833 ; n47833_not
g92041 not n56860 ; n56860_not
g92042 not n47761 ; n47761_not
g92043 not n45781 ; n45781_not
g92044 not n46744 ; n46744_not
g92045 not n47167 ; n47167_not
g92046 not n49147 ; n49147_not
g92047 not n48850 ; n48850_not
g92048 not n54295 ; n54295_not
g92049 not n48616 ; n48616_not
g92050 not n52288 ; n52288_not
g92051 not n48841 ; n48841_not
g92052 not n46186 ; n46186_not
g92053 not n53584 ; n53584_not
g92054 not n47383 ; n47383_not
g92055 not n46168 ; n46168_not
g92056 not n45835 ; n45835_not
g92057 not n49138 ; n49138_not
g92058 not n44971 ; n44971_not
g92059 not n46951 ; n46951_not
g92060 not n56266 ; n56266_not
g92061 not n57292 ; n57292_not
g92062 not n46177 ; n46177_not
g92063 not n45925 ; n45925_not
g92064 not n46960 ; n46960_not
g92065 not n56167 ; n56167_not
g92066 not n46276 ; n46276_not
g92067 not n57427 ; n57427_not
g92068 not n51595 ; n51595_not
g92069 not n44773 ; n44773_not
g92070 not n52657 ; n52657_not
g92071 not n48625 ; n48625_not
g92072 not n44890 ; n44890_not
g92073 not n53728 ; n53728_not
g92074 not n56950 ; n56950_not
g92075 not n48067 ; n48067_not
g92076 not n48058 ; n48058_not
g92077 not n53557 ; n53557_not
g92078 not n53395 ; n53395_not
g92079 not n57436 ; n57436_not
g92080 not n47275 ; n47275_not
g92081 not n48805 ; n48805_not
g92082 not n57418 ; n57418_not
g92083 not n48049 ; n48049_not
g92084 not n45736 ; n45736_not
g92085 not n47806 ; n47806_not
g92086 not n44935 ; n44935_not
g92087 not n46267 ; n46267_not
g92088 not n47446 ; n47446_not
g92089 not n56176 ; n56176_not
g92090 not n51766 ; n51766_not
g92091 not n52648 ; n52648_not
g92092 not n56068 ; n56068_not
g92093 not n46780 ; n46780_not
g92094 not n46654 ; n46654_not
g92095 not n51991 ; n51991_not
g92096 not n56086 ; n56086_not
g92097 not n47455 ; n47455_not
g92098 not n52675 ; n52675_not
g92099 not n46285 ; n46285_not
g92100 not n46915 ; n46915_not
g92101 not n54079 ; n54079_not
g92102 not n44692 ; n44692_not
g92103 not n51982 ; n51982_not
g92104 not n48076 ; n48076_not
g92105 not n51658 ; n51658_not
g92106 not n57481 ; n57481_not
g92107 not n45196 ; n45196_not
g92108 not n57490 ; n57490_not
g92109 not n51973 ; n51973_not
g92110 not n53386 ; n53386_not
g92111 not n44926 ; n44926_not
g92112 not n49633 ; n49633_not
g92113 not n49219 ; n49219_not
g92114 not n56158 ; n56158_not
g92115 not n53737 ; n53737_not
g92116 not n56077 ; n56077_not
g92117 not n54349 ; n54349_not
g92118 not n46825 ; n46825_not
g92119 not n56149 ; n56149_not
g92120 not n53566 ; n53566_not
g92121 not n57454 ; n57454_not
g92122 not n46771 ; n46771_not
g92123 not n54574 ; n54574_not
g92124 not n47293 ; n47293_not
g92125 not n54565 ; n54565_not
g92126 not n46834 ; n46834_not
g92127 not n48823 ; n48823_not
g92128 not n57382 ; n57382_not
g92129 not n45871 ; n45871_not
g92130 not n44854 ; n44854_not
g92131 not n49192 ; n49192_not
g92132 not n44818 ; n44818_not
g92133 not n47419 ; n47419_not
g92134 not n44953 ; n44953_not
g92135 not n53449 ; n53449_not
g92136 not n45916 ; n45916_not
g92137 not n51586 ; n51586_not
g92138 not n57364 ; n57364_not
g92139 not n54484 ; n54484_not
g92140 not n46447 ; n46447_not
g92141 not n47428 ; n47428_not
g92142 not n56914 ; n56914_not
g92143 not n48670 ; n48670_not
g92144 not n47914 ; n47914_not
g92145 not n49183 ; n49183_not
g92146 not n52585 ; n52585_not
g92147 not n54196 ; n54196_not
g92148 not n48652 ; n48652_not
g92149 not n56194 ; n56194_not
g92150 not n45745 ; n45745_not
g92151 not n44845 ; n44845_not
g92152 not n51757 ; n51757_not
g92153 not n56185 ; n56185_not
g92154 not n46249 ; n46249_not
g92155 not n56941 ; n56941_not
g92156 not n46258 ; n46258_not
g92157 not n44683 ; n44683_not
g92158 not n47608 ; n47608_not
g92159 not n51748 ; n51748_not
g92160 not n46762 ; n46762_not
g92161 not n44944 ; n44944_not
g92162 not n57409 ; n57409_not
g92163 not n45754 ; n45754_not
g92164 not n47437 ; n47437_not
g92165 not n52099 ; n52099_not
g92166 not n50974 ; n50974_not
g92167 not n53719 ; n53719_not
g92168 not n50983 ; n50983_not
g92169 not n45880 ; n45880_not
g92170 not n57139 ; n57139_not
g92171 not n47707 ; n47707_not
g92172 not n56671 ; n56671_not
g92173 not n56680 ; n56680_not
g92174 not n56662 ; n56662_not
g92175 not n56653 ; n56653_not
g92176 not n56770 ; n56770_not
g92177 not n46690 ; n46690_not
g92178 not n56644 ; n56644_not
g92179 not n49930 ; n49930_not
g92180 not n49912 ; n49912_not
g92181 not n55807 ; n55807_not
g92182 not n49921 ; n49921_not
g92183 not n56761 ; n56761_not
g92184 not n47464 ; n47464_not
g92185 not n53476 ; n53476_not
g92186 not n56743 ; n56743_not
g92187 not n44467 ; n44467_not
g92188 not n44782 ; n44782_not
g92189 not n53629 ; n53629_not
g92190 not n56725 ; n56725_not
g92191 not n56716 ; n56716_not
g92192 not n44458 ; n44458_not
g92193 not n46870 ; n46870_not
g92194 not n44863 ; n44863_not
g92195 not n56608 ; n56608_not
g92196 not n47725 ; n47725_not
g92197 not n44665 ; n44665_not
g92198 not n46672 ; n46672_not
g92199 not n49039 ; n49039_not
g92200 not n57166 ; n57166_not
g92201 not n45097 ; n45097_not
g92202 not n53638 ; n53638_not
g92203 not n46861 ; n46861_not
g92204 not n49903 ; n49903_not
g92205 not n56590 ; n56590_not
g92206 not n56635 ; n56635_not
g92207 not n48742 ; n48742_not
g92208 not n57148 ; n57148_not
g92209 not n46717 ; n46717_not
g92210 not n55816 ; n55816_not
g92211 not n53485 ; n53485_not
g92212 not n56626 ; n56626_not
g92213 not n48913 ; n48913_not
g92214 not n45718 ; n45718_not
g92215 not n47716 ; n47716_not
g92216 not n55168 ; n55168_not
g92217 not n56617 ; n56617_not
g92218 not n46681 ; n46681_not
g92219 not n47851 ; n47851_not
g92220 not n46852 ; n46852_not
g92221 not n57058 ; n57058_not
g92222 not n47518 ; n47518_not
g92223 not n46708 ; n46708_not
g92224 not n57049 ; n57049_not
g92225 not n47635 ; n47635_not
g92226 not n47626 ; n47626_not
g92227 not n46816 ; n46816_not
g92228 not n47644 ; n47644_not
g92229 not n47653 ; n47653_not
g92230 not n47545 ; n47545_not
g92231 not n47662 ; n47662_not
g92232 not n49606 ; n49606_not
g92233 not n45763 ; n45763_not
g92234 not n48931 ; n48931_not
g92235 not n47248 ; n47248_not
g92236 not n56734 ; n56734_not
g92237 not n57094 ; n57094_not
g92238 not n48733 ; n48733_not
g92239 not n57076 ; n57076_not
g92240 not n48940 ; n48940_not
g92241 not n47527 ; n47527_not
g92242 not n48760 ; n48760_not
g92243 not n57067 ; n57067_not
g92244 not n44656 ; n44656_not
g92245 not n47536 ; n47536_not
g92246 not n46483 ; n46483_not
g92247 not n53494 ; n53494_not
g92248 not n48922 ; n48922_not
g92249 not n56833 ; n56833_not
g92250 not n47491 ; n47491_not
g92251 not n44638 ; n44638_not
g92252 not n54259 ; n54259_not
g92253 not n47482 ; n47482_not
g92254 not n56815 ; n56815_not
g92255 not n48706 ; n48706_not
g92256 not n56806 ; n56806_not
g92257 not n47473 ; n47473_not
g92258 not n47671 ; n47671_not
g92259 not n54169 ; n54169_not
g92260 not n51676 ; n51676_not
g92261 not n47554 ; n47554_not
g92262 not n45970 ; n45970_not
g92263 not n47509 ; n47509_not
g92264 not n56923 ; n56923_not
g92265 not n47680 ; n47680_not
g92266 not n46807 ; n46807_not
g92267 not n47581 ; n47581_not
g92268 not n56419 ; n56419_not
g92269 not n49075 ; n49075_not
g92270 not n47590 ; n47590_not
g92271 not n55933 ; n55933_not
g92272 not n49615 ; n49615_not
g92273 not n53656 ; n53656_not
g92274 not n51667 ; n51667_not
g92275 not n52468 ; n52468_not
g92276 not n45673 ; n45673_not
g92277 not n45943 ; n45943_not
g92278 not n55942 ; n55942_not
g92279 not n52477 ; n52477_not
g92280 not n52369 ; n52369_not
g92281 not n54475 ; n54475_not
g92282 not n48661 ; n48661_not
g92283 not n56446 ; n56446_not
g92284 not n46096 ; n46096_not
g92285 not n56824 ; n56824_not
g92286 not n48715 ; n48715_not
g92287 not n56437 ; n56437_not
g92288 not n45691 ; n45691_not
g92289 not n44836 ; n44836_not
g92290 not n56428 ; n56428_not
g92291 not n47338 ; n47338_not
g92292 not n45682 ; n45682_not
g92293 not n44449 ; n44449_not
g92294 not n52495 ; n52495_not
g92295 not n49624 ; n49624_not
g92296 not n56356 ; n56356_not
g92297 not n56347 ; n56347_not
g92298 not n52297 ; n52297_not
g92299 not n47923 ; n47923_not
g92300 not n46735 ; n46735_not
g92301 not n56338 ; n56338_not
g92302 not n44629 ; n44629_not
g92303 not n56392 ; n56392_not
g92304 not n55951 ; n55951_not
g92305 not n44647 ; n44647_not
g92306 not n57238 ; n57238_not
g92307 not n46726 ; n46726_not
g92308 not n50866 ; n50866_not
g92309 not n54538 ; n54538_not
g92310 not n56383 ; n56383_not
g92311 not n53665 ; n53665_not
g92312 not n56374 ; n56374_not
g92313 not n49084 ; n49084_not
g92314 not n47347 ; n47347_not
g92315 not n47617 ; n47617_not
g92316 not n56365 ; n56365_not
g92317 not n48751 ; n48751_not
g92318 not n55861 ; n55861_not
g92319 not n57193 ; n57193_not
g92320 not n56545 ; n56545_not
g92321 not n49048 ; n49048_not
g92322 not n48904 ; n48904_not
g92323 not n45952 ; n45952_not
g92324 not n56536 ; n56536_not
g92325 not n47941 ; n47941_not
g92326 not n54286 ; n54286_not
g92327 not n56527 ; n56527_not
g92328 not n53458 ; n53458_not
g92329 not n56581 ; n56581_not
g92330 not n45961 ; n45961_not
g92331 not n55843 ; n55843_not
g92332 not n51559 ; n51559_not
g92333 not n47734 ; n47734_not
g92334 not n56572 ; n56572_not
g92335 not n46492 ; n46492_not
g92336 not n46663 ; n46663_not
g92337 not n56563 ; n56563_not
g92338 not n55852 ; n55852_not
g92339 not n56554 ; n56554_not
g92340 not n51568 ; n51568_not
g92341 not n52387 ; n52387_not
g92342 not n56482 ; n56482_not
g92343 not n47572 ; n47572_not
g92344 not n56473 ; n56473_not
g92345 not n45808 ; n45808_not
g92346 not n52378 ; n52378_not
g92347 not n55906 ; n55906_not
g92348 not n49066 ; n49066_not
g92349 not n46087 ; n46087_not
g92350 not n56464 ; n56464_not
g92351 not n56455 ; n56455_not
g92352 not n50839 ; n50839_not
g92353 not n55159 ; n55159_not
g92354 not n53647 ; n53647_not
g92355 not n53593 ; n53593_not
g92356 not n56518 ; n56518_not
g92357 not n54529 ; n54529_not
g92358 not n46069 ; n46069_not
g92359 not n52396 ; n52396_not
g92360 not n56509 ; n56509_not
g92361 not n49057 ; n49057_not
g92362 not n47563 ; n47563_not
g92363 not n45844 ; n45844_not
g92364 not n56491 ; n56491_not
g92365 not n46078 ; n46078_not
g92366 not n54691 ; n54691_not
g92367 not n55069 ; n55069_not
g92368 not n54916 ; n54916_not
g92369 not n47932 ; n47932_not
g92370 not n49444 ; n49444_not
g92371 not n50992 ; n50992_not
g92372 not n49570 ; n49570_not
g92373 not n54907 ; n54907_not
g92374 not n51793 ; n51793_not
g92375 not n46573 ; n46573_not
g92376 not n48292 ; n48292_not
g92377 not n55177 ; n55177_not
g92378 not n46555 ; n46555_not
g92379 not n51289 ; n51289_not
g92380 not n54934 ; n54934_not
g92381 not n51298 ; n51298_not
g92382 not n54943 ; n54943_not
g92383 not n49435 ; n49435_not
g92384 not n47176 ; n47176_not
g92385 not n48256 ; n48256_not
g92386 not n54709 ; n54709_not
g92387 not n49525 ; n49525_not
g92388 not n49534 ; n49534_not
g92389 not n48247 ; n48247_not
g92390 not n45187 ; n45187_not
g92391 not n54457 ; n54457_not
g92392 not n53269 ; n53269_not
g92393 not n49462 ; n49462_not
g92394 not n46582 ; n46582_not
g92395 not n48283 ; n48283_not
g92396 not n44755 ; n44755_not
g92397 not n51685 ; n51685_not
g92398 not n49480 ; n49480_not
g92399 not n48274 ; n48274_not
g92400 not n49750 ; n49750_not
g92401 not n49507 ; n49507_not
g92402 not n48265 ; n48265_not
g92403 not n48346 ; n48346_not
g92404 not n49354 ; n49354_not
g92405 not n53881 ; n53881_not
g92406 not n44359 ; n44359_not
g92407 not n49372 ; n49372_not
g92408 not n54673 ; n54673_not
g92409 not n51892 ; n51892_not
g92410 not n48337 ; n48337_not
g92411 not n54583 ; n54583_not
g92412 not n54664 ; n54664_not
g92413 not n55870 ; n55870_not
g92414 not n48355 ; n48355_not
g92415 not n53359 ; n53359_not
g92416 not n53872 ; n53872_not
g92417 not n55825 ; n55825_not
g92418 not n51865 ; n51865_not
g92419 not n44728 ; n44728_not
g92420 not n48319 ; n48319_not
g92421 not n53890 ; n53890_not
g92422 not n51847 ; n51847_not
g92423 not n54682 ; n54682_not
g92424 not n55078 ; n55078_not
g92425 not n51838 ; n51838_not
g92426 not n49417 ; n49417_not
g92427 not n49390 ; n49390_not
g92428 not n49363 ; n49363_not
g92429 not n54088 ; n54088_not
g92430 not n51883 ; n51883_not
g92431 not n48328 ; n48328_not
g92432 not n46528 ; n46528_not
g92433 not n46537 ; n46537_not
g92434 not n44764 ; n44764_not
g92435 not n49723 ; n49723_not
g92436 not n50947 ; n50947_not
g92437 not n44737 ; n44737_not
g92438 not n53980 ; n53980_not
g92439 not n48166 ; n48166_not
g92440 not n53296 ; n53296_not
g92441 not n54376 ; n54376_not
g92442 not n49732 ; n49732_not
g92443 not n53971 ; n53971_not
g92444 not n54790 ; n54790_not
g92445 not n46618 ; n46618_not
g92446 not n49741 ; n49741_not
g92447 not n54817 ; n54817_not
g92448 not n48139 ; n48139_not
g92449 not n48184 ; n48184_not
g92450 not n49705 ; n49705_not
g92451 not n54736 ; n54736_not
g92452 not n53926 ; n53926_not
g92453 not n54808 ; n54808_not
g92454 not n48175 ; n48175_not
g92455 not n49822 ; n49822_not
g92456 not n49714 ; n49714_not
g92457 not n45169 ; n45169_not
g92458 not n53944 ; n53944_not
g92459 not n54763 ; n54763_not
g92460 not n49804 ; n49804_not
g92461 not n54754 ; n54754_not
g92462 not n48148 ; n48148_not
g92463 not n44746 ; n44746_not
g92464 not n53962 ; n53962_not
g92465 not n54745 ; n54745_not
g92466 not n54781 ; n54781_not
g92467 not n48157 ; n48157_not
g92468 not n53953 ; n53953_not
g92469 not n49813 ; n49813_not
g92470 not n53935 ; n53935_not
g92471 not n54772 ; n54772_not
g92472 not n49453 ; n49453_not
g92473 not n54718 ; n54718_not
g92474 not n54439 ; n54439_not
g92475 not n48229 ; n48229_not
g92476 not n51379 ; n51379_not
g92477 not n49543 ; n49543_not
g92478 not n44719 ; n44719_not
g92479 not n49552 ; n49552_not
g92480 not n51775 ; n51775_not
g92481 not n54448 ; n54448_not
g92482 not n48238 ; n48238_not
g92483 not n54880 ; n54880_not
g92484 not n53908 ; n53908_not
g92485 not n49651 ; n49651_not
g92486 not n54727 ; n54727_not
g92487 not n51397 ; n51397_not
g92488 not n46591 ; n46591_not
g92489 not n54835 ; n54835_not
g92490 not n49660 ; n49660_not
g92491 not n49831 ; n49831_not
g92492 not n48193 ; n48193_not
g92493 not n53917 ; n53917_not
g92494 not n54826 ; n54826_not
g92495 not n52486 ; n52486_not
g92496 not n54970 ; n54970_not
g92497 not n54871 ; n54871_not
g92498 not n54862 ; n54862_not
g92499 not n51388 ; n51388_not
g92500 not n49408 ; n49408_not
g92501 not n49642 ; n49642_not
g92502 not n54853 ; n54853_not
g92503 not n49840 ; n49840_not
g92504 not n54844 ; n54844_not
g92505 not n46627 ; n46627_not
g92506 not n46339 ; n46339_not
g92507 not n53773 ; n53773_not
g92508 not n47059 ; n47059_not
g92509 not n54358 ; n54358_not
g92510 not n48526 ; n48526_not
g92511 not n49255 ; n49255_not
g92512 not n46348 ; n46348_not
g92513 not n47068 ; n47068_not
g92514 not n51955 ; n51955_not
g92515 not n47266 ; n47266_not
g92516 not n51964 ; n51964_not
g92517 not n52693 ; n52693_not
g92518 not n48535 ; n48535_not
g92519 not n49246 ; n49246_not
g92520 not n48094 ; n48094_not
g92521 not n54592 ; n54592_not
g92522 not n48508 ; n48508_not
g92523 not n51478 ; n51478_not
g92524 not n46375 ; n46375_not
g92525 not n47095 ; n47095_not
g92526 not n49309 ; n49309_not
g92527 not n46357 ; n46357_not
g92528 not n53809 ; n53809_not
g92529 not n49273 ; n49273_not
g92530 not n53782 ; n53782_not
g92531 not n51487 ; n51487_not
g92532 not n48553 ; n48553_not
g92533 not n47077 ; n47077_not
g92534 not n48517 ; n48517_not
g92535 not n49264 ; n49264_not
g92536 not n52666 ; n52666_not
g92537 not n46366 ; n46366_not
g92538 not n53791 ; n53791_not
g92539 not n46294 ; n46294_not
g92540 not n44917 ; n44917_not
g92541 not n53368 ; n53368_not
g92542 not n49237 ; n49237_not
g92543 not n49228 ; n49228_not
g92544 not n54925 ; n54925_not
g92545 not n56095 ; n56095_not
g92546 not n51946 ; n51946_not
g92547 not n53746 ; n53746_not
g92548 not n51937 ; n51937_not
g92549 not n48571 ; n48571_not
g92550 not n45709 ; n45709_not
g92551 not n48562 ; n48562_not
g92552 not n47086 ; n47086_not
g92553 not n53764 ; n53764_not
g92554 not n54385 ; n54385_not
g92555 not n51496 ; n51496_not
g92556 not n44908 ; n44908_not
g92557 not n54952 ; n54952_not
g92558 not n45079 ; n45079_not
g92559 not n53755 ; n53755_not
g92560 not n48085 ; n48085_not
g92561 not n48580 ; n48580_not
g92562 not n48418 ; n48418_not
g92563 not n53845 ; n53845_not
g92564 not n49327 ; n49327_not
g92565 not n54637 ; n54637_not
g92566 not n48409 ; n48409_not
g92567 not n44377 ; n44377_not
g92568 not n54178 ; n54178_not
g92569 not n55087 ; n55087_not
g92570 not n54655 ; n54655_not
g92571 not n48427 ; n48427_not
g92572 not n53278 ; n53278_not
g92573 not n54646 ; n54646_not
g92574 not n46465 ; n46465_not
g92575 not n51199 ; n51199_not
g92576 not n48373 ; n48373_not
g92577 not n53863 ; n53863_not
g92578 not n49345 ; n49345_not
g92579 not n48364 ; n48364_not
g92580 not n46393 ; n46393_not
g92581 not n55915 ; n55915_not
g92582 not n54628 ; n54628_not
g92583 not n44368 ; n44368_not
g92584 not n53854 ; n53854_not
g92585 not n54619 ; n54619_not
g92586 not n48391 ; n48391_not
g92587 not n52576 ; n52576_not
g92588 not n48382 ; n48382_not
g92589 not n53818 ; n53818_not
g92590 not n48481 ; n48481_not
g92591 not n48472 ; n48472_not
g92592 not n48490 ; n48490_not
g92593 not n49318 ; n49318_not
g92594 not n51469 ; n51469_not
g92595 not n48445 ; n48445_not
g92596 not n46546 ; n46546_not
g92597 not n49282 ; n49282_not
g92598 not n53836 ; n53836_not
g92599 not n48436 ; n48436_not
g92600 not n53827 ; n53827_not
g92601 not n48463 ; n48463_not
g92602 not n47842 ; n47842_not
g92603 not n54268 ; n54268_not
g92604 not n46438 ; n46438_not
g92605 not n48454 ; n48454_not
g92606 not n55960 ; n55960_not
g92607 not n51856 ; n51856_not
g92608 not n15298 ; n15298_not
g92609 not n15289 ; n15289_not
g92610 not n15199 ; n15199_not
g92611 not n18637 ; n18637_not
g92612 not n14596 ; n14596_not
g92613 not n18628 ; n18628_not
g92614 not n35692 ; n35692_not
g92615 not n35683 ; n35683_not
g92616 not n28186 ; n28186_not
g92617 not n39940 ; n39940_not
g92618 not n19285 ; n19285_not
g92619 not n28195 ; n28195_not
g92620 not n23686 ; n23686_not
g92621 not n39931 ; n39931_not
g92622 not n27925 ; n27925_not
g92623 not n18619 ; n18619_not
g92624 not n23596 ; n23596_not
g92625 not n23659 ; n23659_not
g92626 not n23668 ; n23668_not
g92627 not n35638 ; n35638_not
g92628 not n35647 ; n35647_not
g92629 not n39904 ; n39904_not
g92630 not n39913 ; n39913_not
g92631 not n35665 ; n35665_not
g92632 not n39922 ; n39922_not
g92633 not n23758 ; n23758_not
g92634 not n35773 ; n35773_not
g92635 not n18655 ; n18655_not
g92636 not n19267 ; n19267_not
g92637 not n15397 ; n15397_not
g92638 not n18664 ; n18664_not
g92639 not n38473 ; n38473_not
g92640 not n23776 ; n23776_not
g92641 not n18673 ; n18673_not
g92642 not n35782 ; n35782_not
g92643 not n19258 ; n19258_not
g92644 not n15469 ; n15469_not
g92645 not n18682 ; n18682_not
g92646 not n15478 ; n15478_not
g92647 not n28159 ; n28159_not
g92648 not n35728 ; n35728_not
g92649 not n28069 ; n28069_not
g92650 not n35737 ; n35737_not
g92651 not n37573 ; n37573_not
g92652 not n37582 ; n37582_not
g92653 not n23749 ; n23749_not
g92654 not n28096 ; n28096_not
g92655 not n35755 ; n35755_not
g92656 not n18646 ; n18646_not
g92657 not n28078 ; n28078_not
g92658 not n15379 ; n15379_not
g92659 not n15388 ; n15388_not
g92660 not n35449 ; n35449_not
g92661 not n27835 ; n27835_not
g92662 not n35458 ; n35458_not
g92663 not n19348 ; n19348_not
g92664 not n19276 ; n19276_not
g92665 not n35467 ; n35467_not
g92666 not n14974 ; n14974_not
g92667 not n14992 ; n14992_not
g92668 not n19339 ; n19339_not
g92669 not n23488 ; n23488_not
g92670 not n35476 ; n35476_not
g92671 not n35485 ; n35485_not
g92672 not n28285 ; n28285_not
g92673 not n39805 ; n39805_not
g92674 not n35296 ; n35296_not
g92675 not n39760 ; n39760_not
g92676 not n35287 ; n35287_not
g92677 not n39751 ; n39751_not
g92678 not n39733 ; n39733_not
g92679 not n14983 ; n14983_not
g92680 not n22867 ; n22867_not
g92681 not n39742 ; n39742_not
g92682 not n27826 ; n27826_not
g92683 not n35278 ; n35278_not
g92684 not n22849 ; n22849_not
g92685 not n39850 ; n39850_not
g92686 not n35539 ; n35539_not
g92687 not n35548 ; n35548_not
g92688 not n23569 ; n23569_not
g92689 not n35557 ; n35557_not
g92690 not n35566 ; n35566_not
g92691 not n23578 ; n23578_not
g92692 not n35575 ; n35575_not
g92693 not n35197 ; n35197_not
g92694 not n35584 ; n35584_not
g92695 not n23587 ; n23587_not
g92696 not n27916 ; n27916_not
g92697 not n35593 ; n35593_not
g92698 not n37564 ; n37564_not
g92699 not n22858 ; n22858_not
g92700 not n39814 ; n39814_not
g92701 not n28276 ; n28276_not
g92702 not n35494 ; n35494_not
g92703 not n39823 ; n39823_not
g92704 not n23497 ; n23497_not
g92705 not n39832 ; n39832_not
g92706 not n39841 ; n39841_not
g92707 not n28267 ; n28267_not
g92708 not n28258 ; n28258_not
g92709 not n35890 ; n35890_not
g92710 not n18871 ; n18871_not
g92711 not n15829 ; n15829_not
g92712 not n18862 ; n18862_not
g92713 not n39724 ; n39724_not
g92714 not n27853 ; n27853_not
g92715 not n18853 ; n18853_not
g92716 not n15784 ; n15784_not
g92717 not n35881 ; n35881_not
g92718 not n18844 ; n18844_not
g92719 not n18835 ; n18835_not
g92720 not n18808 ; n18808_not
g92721 not n18817 ; n18817_not
g92722 not n35863 ; n35863_not
g92723 not n19177 ; n19177_not
g92724 not n18826 ; n18826_not
g92725 not n15739 ; n15739_not
g92726 not n15757 ; n15757_not
g92727 not n15766 ; n15766_not
g92728 not n35872 ; n35872_not
g92729 not n19168 ; n19168_not
g92730 not n27880 ; n27880_not
g92731 not n23866 ; n23866_not
g92732 not n27871 ; n27871_not
g92733 not n23884 ; n23884_not
g92734 not n18943 ; n18943_not
g92735 not n18952 ; n18952_not
g92736 not n23893 ; n23893_not
g92737 not n18961 ; n18961_not
g92738 not n35917 ; n35917_not
g92739 not n27790 ; n27790_not
g92740 not n35926 ; n35926_not
g92741 not n27772 ; n27772_not
g92742 not n27781 ; n27781_not
g92743 not n35935 ; n35935_not
g92744 not n18970 ; n18970_not
g92745 not n18880 ; n18880_not
g92746 not n18907 ; n18907_not
g92747 not n18916 ; n18916_not
g92748 not n15847 ; n15847_not
g92749 not n18925 ; n18925_not
g92750 not n18934 ; n18934_not
g92751 not n27808 ; n27808_not
g92752 not n35908 ; n35908_not
g92753 not n15559 ; n15559_not
g92754 not n15568 ; n15568_not
g92755 not n18727 ; n18727_not
g92756 not n35746 ; n35746_not
g92757 not n39544 ; n39544_not
g92758 not n15577 ; n15577_not
g92759 not n18736 ; n18736_not
g92760 not n18745 ; n18745_not
g92761 not n35809 ; n35809_not
g92762 not n15586 ; n15586_not
g92763 not n18754 ; n18754_not
g92764 not n15487 ; n15487_not
g92765 not n18691 ; n18691_not
g92766 not n27970 ; n27970_not
g92767 not n15496 ; n15496_not
g92768 not n38464 ; n38464_not
g92769 not n35791 ; n35791_not
g92770 not n18709 ; n18709_not
g92771 not n27961 ; n27961_not
g92772 not n18718 ; n18718_not
g92773 not n15649 ; n15649_not
g92774 not n18781 ; n18781_not
g92775 not n35845 ; n35845_not
g92776 not n39562 ; n39562_not
g92777 not n23839 ; n23839_not
g92778 not n15667 ; n15667_not
g92779 not n15676 ; n15676_not
g92780 not n18790 ; n18790_not
g92781 not n19195 ; n19195_not
g92782 not n23848 ; n23848_not
g92783 not n35854 ; n35854_not
g92784 not n15694 ; n15694_not
g92785 not n35818 ; n35818_not
g92786 not n27943 ; n27943_not
g92787 not n15595 ; n15595_not
g92788 not n18763 ; n18763_not
g92789 not n35827 ; n35827_not
g92790 not n39553 ; n39553_not
g92791 not n18772 ; n18772_not
g92792 not n35836 ; n35836_not
g92793 not n23794 ; n23794_not
g92794 not n28618 ; n28618_not
g92795 not n27934 ; n27934_not
g92796 not n14668 ; n14668_not
g92797 not n40993 ; n40993_not
g92798 not n34819 ; n34819_not
g92799 not n28627 ; n28627_not
g92800 not n34918 ; n34918_not
g92801 not n14659 ; n14659_not
g92802 not n34828 ; n34828_not
g92803 not n28636 ; n28636_not
g92804 not n19186 ; n19186_not
g92805 not n28645 ; n28645_not
g92806 not n22993 ; n22993_not
g92807 not n22966 ; n22966_not
g92808 not n13957 ; n13957_not
g92809 not n14569 ; n14569_not
g92810 not n28672 ; n28672_not
g92811 not n19519 ; n19519_not
g92812 not n40687 ; n40687_not
g92813 not n28663 ; n28663_not
g92814 not n28654 ; n28654_not
g92815 not n40696 ; n40696_not
g92816 not n22984 ; n22984_not
g92817 not n40948 ; n40948_not
g92818 not n38518 ; n38518_not
g92819 not n40786 ; n40786_not
g92820 not n28546 ; n28546_not
g92821 not n40939 ; n40939_not
g92822 not n40795 ; n40795_not
g92823 not n35089 ; n35089_not
g92824 not n28537 ; n28537_not
g92825 not n23299 ; n23299_not
g92826 not n14695 ; n14695_not
g92827 not n19483 ; n19483_not
g92828 not n35098 ; n35098_not
g92829 not n28528 ; n28528_not
g92830 not n28609 ; n28609_not
g92831 not n28591 ; n28591_not
g92832 not n40984 ; n40984_not
g92833 not n28582 ; n28582_not
g92834 not n40975 ; n40975_not
g92835 not n14677 ; n14677_not
g92836 not n28573 ; n28573_not
g92837 not n19492 ; n19492_not
g92838 not n28564 ; n28564_not
g92839 not n14686 ; n14686_not
g92840 not n40966 ; n40966_not
g92841 not n40777 ; n40777_not
g92842 not n28555 ; n28555_not
g92843 not n40957 ; n40957_not
g92844 not n28780 ; n28780_not
g92845 not n41596 ; n41596_not
g92846 not n19564 ; n19564_not
g92847 not n41587 ; n41587_not
g92848 not n13795 ; n13795_not
g92849 not n28771 ; n28771_not
g92850 not n41578 ; n41578_not
g92851 not n13786 ; n13786_not
g92852 not n41569 ; n41569_not
g92853 not n28762 ; n28762_not
g92854 not n28168 ; n28168_not
g92855 not n19555 ; n19555_not
g92856 not n13777 ; n13777_not
g92857 not n28753 ; n28753_not
g92858 not n28744 ; n28744_not
g92859 not n14299 ; n14299_not
g92860 not n41686 ; n41686_not
g92861 not n19582 ; n19582_not
g92862 not n28834 ; n28834_not
g92863 not n34864 ; n34864_not
g92864 not n41677 ; n41677_not
g92865 not n28825 ; n28825_not
g92866 not n41668 ; n41668_not
g92867 not n19573 ; n19573_not
g92868 not n41659 ; n41659_not
g92869 not n28816 ; n28816_not
g92870 not n28807 ; n28807_not
g92871 not n38545 ; n38545_not
g92872 not n37528 ; n37528_not
g92873 not n22939 ; n22939_not
g92874 not n19537 ; n19537_not
g92875 not n14497 ; n14497_not
g92876 not n22948 ; n22948_not
g92877 not n28690 ; n28690_not
g92878 not n41398 ; n41398_not
g92879 not n19528 ; n19528_not
g92880 not n28681 ; n28681_not
g92881 not n37537 ; n37537_not
g92882 not n22876 ; n22876_not
g92883 not n28735 ; n28735_not
g92884 not n41497 ; n41497_not
g92885 not n28726 ; n28726_not
g92886 not n41488 ; n41488_not
g92887 not n22894 ; n22894_not
g92888 not n41479 ; n41479_not
g92889 not n14389 ; n14389_not
g92890 not n34855 ; n34855_not
g92891 not n14479 ; n14479_not
g92892 not n19546 ; n19546_not
g92893 not n28717 ; n28717_not
g92894 not n40867 ; n40867_not
g92895 not n28708 ; n28708_not
g92896 not n19384 ; n19384_not
g92897 not n40399 ; n40399_not
g92898 not n28429 ; n28429_not
g92899 not n19393 ; n19393_not
g92900 not n28438 ; n28438_not
g92901 not n14893 ; n14893_not
g92902 not n34927 ; n34927_not
g92903 not n28447 ; n28447_not
g92904 not n14884 ; n14884_not
g92905 not n28456 ; n28456_not
g92906 not n34945 ; n34945_not
g92907 not n14875 ; n14875_not
g92908 not n27844 ; n27844_not
g92909 not n28465 ; n28465_not
g92910 not n14839 ; n14839_not
g92911 not n34981 ; n34981_not
g92912 not n14848 ; n14848_not
g92913 not n28483 ; n28483_not
g92914 not n34972 ; n34972_not
g92915 not n14857 ; n14857_not
g92916 not n28474 ; n28474_not
g92917 not n34963 ; n34963_not
g92918 not n14866 ; n14866_not
g92919 not n23398 ; n23398_not
g92920 not n34954 ; n34954_not
g92921 not n14947 ; n14947_not
g92922 not n35377 ; n35377_not
g92923 not n28366 ; n28366_not
g92924 not n28357 ; n28357_not
g92925 not n35386 ; n35386_not
g92926 not n19366 ; n19366_not
g92927 not n14956 ; n14956_not
g92928 not n28348 ; n28348_not
g92929 not n14965 ; n14965_not
g92930 not n35395 ; n35395_not
g92931 not n19357 ; n19357_not
g92932 not n28339 ; n28339_not
g92933 not n23479 ; n23479_not
g92934 not n28393 ; n28393_not
g92935 not n19375 ; n19375_not
g92936 not n28384 ; n28384_not
g92937 not n35359 ; n35359_not
g92938 not n28375 ; n28375_not
g92939 not n35368 ; n35368_not
g92940 not n14929 ; n14929_not
g92941 not n14938 ; n14938_not
g92942 not n14758 ; n14758_not
g92943 not n19465 ; n19465_not
g92944 not n34783 ; n34783_not
g92945 not n40759 ; n40759_not
g92946 not n40489 ; n40489_not
g92947 not n40498 ; n40498_not
g92948 not n34774 ; n34774_not
g92949 not n40894 ; n40894_not
g92950 not n40885 ; n40885_not
g92951 not n28519 ; n28519_not
g92952 not n40876 ; n40876_not
g92953 not n19474 ; n19474_not
g92954 not n14749 ; n14749_not
g92955 not n22957 ; n22957_not
g92956 not n38509 ; n38509_not
g92957 not n14785 ; n14785_not
g92958 not n19438 ; n19438_not
g92959 not n14794 ; n14794_not
g92960 not n23389 ; n23389_not
g92961 not n19429 ; n19429_not
g92962 not n34990 ; n34990_not
g92963 not n40669 ; n40669_not
g92964 not n40579 ; n40579_not
g92965 not n40588 ; n40588_not
g92966 not n40597 ; n40597_not
g92967 not n19456 ; n19456_not
g92968 not n14767 ; n14767_not
g92969 not n28492 ; n28492_not
g92970 not n14776 ; n14776_not
g92971 not n19447 ; n19447_not
g92972 not n24964 ; n24964_not
g92973 not n37096 ; n37096_not
g92974 not n17683 ; n17683_not
g92975 not n24973 ; n24973_not
g92976 not n24982 ; n24982_not
g92977 not n39661 ; n39661_not
g92978 not n17674 ; n17674_not
g92979 not n16972 ; n16972_not
g92980 not n36835 ; n36835_not
g92981 not n24991 ; n24991_not
g92982 not n25369 ; n25369_not
g92983 not n39391 ; n39391_not
g92984 not n36583 ; n36583_not
g92985 not n39049 ; n39049_not
g92986 not n17665 ; n17665_not
g92987 not n36826 ; n36826_not
g92988 not n36718 ; n36718_not
g92989 not n25099 ; n25099_not
g92990 not n37168 ; n37168_not
g92991 not n36709 ; n36709_not
g92992 not n37159 ; n37159_not
g92993 not n18277 ; n18277_not
g92994 not n36808 ; n36808_not
g92995 not n36691 ; n36691_not
g92996 not n18268 ; n18268_not
g92997 not n39058 ; n39058_not
g92998 not n39382 ; n39382_not
g92999 not n36817 ; n36817_not
g93000 not n24586 ; n24586_not
g93001 not n36682 ; n36682_not
g93002 not n36592 ; n36592_not
g93003 not n18259 ; n18259_not
g93004 not n17647 ; n17647_not
g93005 not n36853 ; n36853_not
g93006 not n18187 ; n18187_not
g93007 not n24874 ; n24874_not
g93008 not n39616 ; n39616_not
g93009 not n39418 ; n39418_not
g93010 not n24865 ; n24865_not
g93011 not n24856 ; n24856_not
g93012 not n18178 ; n18178_not
g93013 not n36862 ; n36862_not
g93014 not n18169 ; n18169_not
g93015 not n24847 ; n24847_not
g93016 not n17719 ; n17719_not
g93017 not n25459 ; n25459_not
g93018 not n17728 ; n17728_not
g93019 not n24955 ; n24955_not
g93020 not n16963 ; n16963_not
g93021 not n36844 ; n36844_not
g93022 not n25396 ; n25396_not
g93023 not n24946 ; n24946_not
g93024 not n39643 ; n39643_not
g93025 not n36574 ; n36574_not
g93026 not n39634 ; n39634_not
g93027 not n39409 ; n39409_not
g93028 not n24937 ; n24937_not
g93029 not n18196 ; n18196_not
g93030 not n24928 ; n24928_not
g93031 not n16954 ; n16954_not
g93032 not n24919 ; n24919_not
g93033 not n24892 ; n24892_not
g93034 not n37078 ; n37078_not
g93035 not n24883 ; n24883_not
g93036 not n36736 ; n36736_not
g93037 not n36637 ; n36637_not
g93038 not n18385 ; n18385_not
g93039 not n36745 ; n36745_not
g93040 not n37249 ; n37249_not
g93041 not n36790 ; n36790_not
g93042 not n36628 ; n36628_not
g93043 not n39337 ; n39337_not
g93044 not n24649 ; n24649_not
g93045 not n26368 ; n26368_not
g93046 not n26359 ; n26359_not
g93047 not n36754 ; n36754_not
g93048 not n36781 ; n36781_not
g93049 not n18367 ; n18367_not
g93050 not n26296 ; n26296_not
g93051 not n37276 ; n37276_not
g93052 not n37069 ; n37069_not
g93053 not n18457 ; n18457_not
g93054 not n37267 ; n37267_not
g93055 not n18439 ; n18439_not
g93056 not n39319 ; n39319_not
g93057 not n36727 ; n36727_not
g93058 not n37258 ; n37258_not
g93059 not n39085 ; n39085_not
g93060 not n18394 ; n18394_not
g93061 not n39328 ; n39328_not
g93062 not n39355 ; n39355_not
g93063 not n25279 ; n25279_not
g93064 not n39706 ; n39706_not
g93065 not n39364 ; n39364_not
g93066 not n37195 ; n37195_not
g93067 not n18295 ; n18295_not
g93068 not n37186 ; n37186_not
g93069 not n18286 ; n18286_not
g93070 not n24595 ; n24595_not
g93071 not n37177 ; n37177_not
g93072 not n39373 ; n39373_not
g93073 not n26287 ; n26287_not
g93074 not n36772 ; n36772_not
g93075 not n26269 ; n26269_not
g93076 not n36763 ; n36763_not
g93077 not n39346 ; n39346_not
g93078 not n36619 ; n36619_not
g93079 not n26197 ; n26197_not
g93080 not n26179 ; n26179_not
g93081 not n18349 ; n18349_not
g93082 not n26089 ; n26089_not
g93083 not n25198 ; n25198_not
g93084 not n25189 ; n25189_not
g93085 not n17638 ; n17638_not
g93086 not n17953 ; n17953_not
g93087 not n17944 ; n17944_not
g93088 not n36961 ; n36961_not
g93089 not n17935 ; n17935_not
g93090 not n17908 ; n17908_not
g93091 not n17773 ; n17773_not
g93092 not n39517 ; n39517_not
g93093 not n24829 ; n24829_not
g93094 not n17917 ; n17917_not
g93095 not n24838 ; n24838_not
g93096 not n36952 ; n36952_not
g93097 not n17845 ; n17845_not
g93098 not n39508 ; n39508_not
g93099 not n17926 ; n17926_not
g93100 not n39463 ; n39463_not
g93101 not n17980 ; n17980_not
g93102 not n36970 ; n36970_not
g93103 not n17809 ; n17809_not
g93104 not n25288 ; n25288_not
g93105 not n39472 ; n39472_not
g93106 not n39490 ; n39490_not
g93107 not n24469 ; n24469_not
g93108 not n17962 ; n17962_not
g93109 not n17971 ; n17971_not
g93110 not n25378 ; n25378_not
g93111 not n39481 ; n39481_not
g93112 not n17818 ; n17818_not
g93113 not n24766 ; n24766_not
g93114 not n17782 ; n17782_not
g93115 not n18097 ; n18097_not
g93116 not n36547 ; n36547_not
g93117 not n39571 ; n39571_not
g93118 not n36907 ; n36907_not
g93119 not n24757 ; n24757_not
g93120 not n18088 ; n18088_not
g93121 not n17827 ; n17827_not
g93122 not n36538 ; n36538_not
g93123 not n39445 ; n39445_not
g93124 not n36916 ; n36916_not
g93125 not n24748 ; n24748_not
g93126 not n24739 ; n24739_not
g93127 not n17854 ; n17854_not
g93128 not n36871 ; n36871_not
g93129 not n17692 ; n17692_not
g93130 not n39427 ; n39427_not
g93131 not n24559 ; n24559_not
g93132 not n17737 ; n17737_not
g93133 not n24793 ; n24793_not
g93134 not n36880 ; n36880_not
g93135 not n25486 ; n25486_not
g93136 not n24784 ; n24784_not
g93137 not n17755 ; n17755_not
g93138 not n17764 ; n17764_not
g93139 not n24775 ; n24775_not
g93140 not n39436 ; n39436_not
g93141 not n25495 ; n25495_not
g93142 not n36934 ; n36934_not
g93143 not n17863 ; n17863_not
g93144 not n24496 ; n24496_not
g93145 not n39526 ; n39526_not
g93146 not n36943 ; n36943_not
g93147 not n25468 ; n25468_not
g93148 not n17188 ; n17188_not
g93149 not n36925 ; n36925_not
g93150 not n18079 ; n18079_not
g93151 not n39454 ; n39454_not
g93152 not n36529 ; n36529_not
g93153 not n17890 ; n17890_not
g93154 not n23677 ; n23677_not
g93155 not n37483 ; n37483_not
g93156 not n26962 ; n26962_not
g93157 not n26971 ; n26971_not
g93158 not n36196 ; n36196_not
g93159 not n16369 ; n16369_not
g93160 not n16378 ; n16378_not
g93161 not n18448 ; n18448_not
g93162 not n36178 ; n36178_not
g93163 not n27079 ; n27079_not
g93164 not n27196 ; n27196_not
g93165 not n27187 ; n27187_not
g93166 not n37546 ; n37546_not
g93167 not n16468 ; n16468_not
g93168 not n16459 ; n16459_not
g93169 not n27169 ; n27169_not
g93170 not n23767 ; n23767_not
g93171 not n39139 ; n39139_not
g93172 not n27097 ; n27097_not
g93173 not n36169 ; n36169_not
g93174 not n37519 ; n37519_not
g93175 not n26917 ; n26917_not
g93176 not n26908 ; n26908_not
g93177 not n16279 ; n16279_not
g93178 not n39166 ; n39166_not
g93179 not n36295 ; n36295_not
g93180 not n39175 ; n39175_not
g93181 not n16945 ; n16945_not
g93182 not n18484 ; n18484_not
g93183 not n37456 ; n37456_not
g93184 not n37447 ; n37447_not
g93185 not n39184 ; n39184_not
g93186 not n26944 ; n26944_not
g93187 not n36187 ; n36187_not
g93188 not n39157 ; n39157_not
g93189 not n18475 ; n18475_not
g93190 not n36259 ; n36259_not
g93191 not n36268 ; n36268_not
g93192 not n38644 ; n38644_not
g93193 not n36277 ; n36277_not
g93194 not n26926 ; n26926_not
g93195 not n16288 ; n16288_not
g93196 not n37474 ; n37474_not
g93197 not n36286 ; n36286_not
g93198 not n15775 ; n15775_not
g93199 not n37645 ; n37645_not
g93200 not n35971 ; n35971_not
g93201 not n35980 ; n35980_not
g93202 not n18358 ; n18358_not
g93203 not n37627 ; n37627_not
g93204 not n37618 ; n37618_not
g93205 not n26980 ; n26980_not
g93206 not n35944 ; n35944_not
g93207 not n19087 ; n19087_not
g93208 not n19078 ; n19078_not
g93209 not n35953 ; n35953_not
g93210 not n23857 ; n23857_not
g93211 not n26935 ; n26935_not
g93212 not n37609 ; n37609_not
g93213 not n35656 ; n35656_not
g93214 not n35962 ; n35962_not
g93215 not n16477 ; n16477_not
g93216 not n36079 ; n36079_not
g93217 not n37591 ; n37591_not
g93218 not n16495 ; n16495_not
g93219 not n36088 ; n36088_not
g93220 not n39094 ; n39094_not
g93221 not n15685 ; n15685_not
g93222 not n37636 ; n37636_not
g93223 not n16297 ; n16297_not
g93224 not n16387 ; n16387_not
g93225 not n39607 ; n39607_not
g93226 not n39067 ; n39067_not
g93227 not n18574 ; n18574_not
g93228 not n39283 ; n39283_not
g93229 not n36358 ; n36358_not
g93230 not n36349 ; n36349_not
g93231 not n37375 ; n37375_not
g93232 not n18565 ; n18565_not
g93233 not n17179 ; n17179_not
g93234 not n37393 ; n37393_not
g93235 not n24694 ; n24694_not
g93236 not n36394 ; n36394_not
g93237 not n36385 ; n36385_not
g93238 not n18583 ; n18583_not
g93239 not n24685 ; n24685_not
g93240 not n36376 ; n36376_not
g93241 not n39274 ; n39274_not
g93242 not n36367 ; n36367_not
g93243 not n24676 ; n24676_not
g93244 not n37384 ; n37384_not
g93245 not n18529 ; n18529_not
g93246 not n17098 ; n17098_not
g93247 not n37294 ; n37294_not
g93248 not n17089 ; n17089_not
g93249 not n37285 ; n37285_not
g93250 not n36646 ; n36646_not
g93251 not n37366 ; n37366_not
g93252 not n37357 ; n37357_not
g93253 not n36664 ; n36664_not
g93254 not n39292 ; n39292_not
g93255 not n36673 ; n36673_not
g93256 not n18547 ; n18547_not
g93257 not n37348 ; n37348_not
g93258 not n37339 ; n37339_not
g93259 not n24478 ; n24478_not
g93260 not n24568 ; n24568_not
g93261 not n36097 ; n36097_not
g93262 not n39148 ; n39148_not
g93263 not n18538 ; n18538_not
g93264 not n36439 ; n36439_not
g93265 not n36448 ; n36448_not
g93266 not n36457 ; n36457_not
g93267 not n18493 ; n18493_not
g93268 not n39193 ; n39193_not
g93269 not n37438 ; n37438_not
g93270 not n16981 ; n16981_not
g93271 not n24397 ; n24397_not
g93272 not n37429 ; n37429_not
g93273 not n39652 ; n39652_not
g93274 not n36475 ; n36475_not
g93275 not n36466 ; n36466_not
g93276 not n39256 ; n39256_not
g93277 not n18592 ; n18592_not
g93278 not n36556 ; n36556_not
g93279 not n39265 ; n39265_not
g93280 not n39229 ; n39229_not
g93281 not n36484 ; n36484_not
g93282 not n36493 ; n36493_not
g93283 not n24658 ; n24658_not
g93284 not n39238 ; n39238_not
g93285 not n39247 ; n39247_not
g93286 not n20779 ; n20779_not
g93287 not n19915 ; n19915_not
g93288 not n43891 ; n43891_not
g93289 not n30895 ; n30895_not
g93290 not n33973 ; n33973_not
g93291 not n30886 ; n30886_not
g93292 not n30877 ; n30877_not
g93293 not n38635 ; n38635_not
g93294 not n43909 ; n43909_not
g93295 not n43927 ; n43927_not
g93296 not n30868 ; n30868_not
g93297 not n43945 ; n43945_not
g93298 not n38617 ; n38617_not
g93299 not n37780 ; n37780_not
g93300 not n19924 ; n19924_not
g93301 not n33955 ; n33955_not
g93302 not n43936 ; n43936_not
g93303 not n30958 ; n30958_not
g93304 not n30949 ; n30949_not
g93305 not n30859 ; n30859_not
g93306 not n33964 ; n33964_not
g93307 not n37843 ; n37843_not
g93308 not n30769 ; n30769_not
g93309 not n33991 ; n33991_not
g93310 not n37852 ; n37852_not
g93311 not n43846 ; n43846_not
g93312 not n20689 ; n20689_not
g93313 not n43828 ; n43828_not
g93314 not n43819 ; n43819_not
g93315 not n20698 ; n20698_not
g93316 not n37807 ; n37807_not
g93317 not n37816 ; n37816_not
g93318 not n37825 ; n37825_not
g93319 not n43873 ; n43873_not
g93320 not n37834 ; n37834_not
g93321 not n43864 ; n43864_not
g93322 not n30697 ; n30697_not
g93323 not n38095 ; n38095_not
g93324 not n37717 ; n37717_not
g93325 not n30778 ; n30778_not
g93326 not n30787 ; n30787_not
g93327 not n33874 ; n33874_not
g93328 not n37726 ; n37726_not
g93329 not n19942 ; n19942_not
g93330 not n20788 ; n20788_not
g93331 not n43981 ; n43981_not
g93332 not n38086 ; n38086_not
g93333 not n38572 ; n38572_not
g93334 not n30994 ; n30994_not
g93335 not n33667 ; n33667_not
g93336 not n19960 ; n19960_not
g93337 not n38554 ; n38554_not
g93338 not n33847 ; n33847_not
g93339 not n33685 ; n33685_not
g93340 not n33856 ; n33856_not
g93341 not n37708 ; n37708_not
g93342 not n43990 ; n43990_not
g93343 not n33676 ; n33676_not
g93344 not n20797 ; n20797_not
g93345 not n33865 ; n33865_not
g93346 not n37762 ; n37762_not
g93347 not n30976 ; n30976_not
g93348 not n30796 ; n30796_not
g93349 not n38068 ; n38068_not
g93350 not n38590 ; n38590_not
g93351 not n33919 ; n33919_not
g93352 not n43954 ; n43954_not
g93353 not n33928 ; n33928_not
g93354 not n33937 ; n33937_not
g93355 not n37771 ; n37771_not
g93356 not n33946 ; n33946_not
g93357 not n37735 ; n37735_not
g93358 not n33883 ; n33883_not
g93359 not n43972 ; n43972_not
g93360 not n43882 ; n43882_not
g93361 not n37744 ; n37744_not
g93362 not n37753 ; n37753_not
g93363 not n43963 ; n43963_not
g93364 not n33892 ; n33892_not
g93365 not n43585 ; n43585_not
g93366 not n29752 ; n29752_not
g93367 not n10879 ; n10879_not
g93368 not n37915 ; n37915_not
g93369 not n43576 ; n43576_not
g93370 not n10897 ; n10897_not
g93371 not n29860 ; n29860_not
g93372 not n43567 ; n43567_not
g93373 not n34459 ; n34459_not
g93374 not n43558 ; n43558_not
g93375 not n43549 ; n43549_not
g93376 not n10969 ; n10969_not
g93377 not n34549 ; n34549_not
g93378 not n20599 ; n20599_not
g93379 not n43639 ; n43639_not
g93380 not n34486 ; n34486_not
g93381 not n29905 ; n29905_not
g93382 not n34558 ; n34558_not
g93383 not n34567 ; n34567_not
g93384 not n37906 ; n37906_not
g93385 not n34576 ; n34576_not
g93386 not n34585 ; n34585_not
g93387 not n43594 ; n43594_not
g93388 not n34594 ; n34594_not
g93389 not n43468 ; n43468_not
g93390 not n43459 ; n43459_not
g93391 not n34657 ; n34657_not
g93392 not n10888 ; n10888_not
g93393 not n11689 ; n11689_not
g93394 not n11698 ; n11698_not
g93395 not n11779 ; n11779_not
g93396 not n19825 ; n19825_not
g93397 not n29824 ; n29824_not
g93398 not n11788 ; n11788_not
g93399 not n43396 ; n43396_not
g93400 not n10987 ; n10987_not
g93401 not n29851 ; n29851_not
g93402 not n37924 ; n37924_not
g93403 not n29761 ; n29761_not
g93404 not n29842 ; n29842_not
g93405 not n34639 ; n34639_not
g93406 not n29770 ; n29770_not
g93407 not n43495 ; n43495_not
g93408 not n19834 ; n19834_not
g93409 not n34648 ; n34648_not
g93410 not n43486 ; n43486_not
g93411 not n29833 ; n29833_not
g93412 not n43477 ; n43477_not
g93413 not n10978 ; n10978_not
g93414 not n29932 ; n29932_not
g93415 not n43783 ; n43783_not
g93416 not n29941 ; n29941_not
g93417 not n43774 ; n43774_not
g93418 not n33757 ; n33757_not
g93419 not n19870 ; n19870_not
g93420 not n29950 ; n29950_not
g93421 not n34189 ; n34189_not
g93422 not n34198 ; n34198_not
g93423 not n43756 ; n43756_not
g93424 not n34279 ; n34279_not
g93425 not n37861 ; n37861_not
g93426 not n30598 ; n30598_not
g93427 not n30589 ; n30589_not
g93428 not n37870 ; n37870_not
g93429 not n29923 ; n29923_not
g93430 not n34288 ; n34288_not
g93431 not n34468 ; n34468_not
g93432 not n34495 ; n34495_not
g93433 not n43666 ; n43666_not
g93434 not n43657 ; n43657_not
g93435 not n19852 ; n19852_not
g93436 not n43648 ; n43648_not
g93437 not n34297 ; n34297_not
g93438 not n43738 ; n43738_not
g93439 not n43729 ; n43729_not
g93440 not n34369 ; n34369_not
g93441 not n34378 ; n34378_not
g93442 not n43693 ; n43693_not
g93443 not n34396 ; n34396_not
g93444 not n38248 ; n38248_not
g93445 not n32983 ; n32983_not
g93446 not n32974 ; n32974_not
g93447 not n19618 ; n19618_not
g93448 not n38257 ; n38257_not
g93449 not n38392 ; n38392_not
g93450 not n32956 ; n32956_not
g93451 not n38266 ; n38266_not
g93452 not n44539 ; n44539_not
g93453 not n31885 ; n31885_not
g93454 not n31876 ; n31876_not
g93455 not n31867 ; n31867_not
g93456 not n19933 ; n19933_not
g93457 not n31858 ; n31858_not
g93458 not n38275 ; n38275_not
g93459 not n38059 ; n38059_not
g93460 not n31849 ; n31849_not
g93461 not n38383 ; n38383_not
g93462 not n32578 ; n32578_not
g93463 not n19609 ; n19609_not
g93464 not n44548 ; n44548_not
g93465 not n32929 ; n32929_not
g93466 not n32938 ; n32938_not
g93467 not n44476 ; n44476_not
g93468 not n31957 ; n31957_not
g93469 not n31669 ; n31669_not
g93470 not n19636 ; n19636_not
g93471 not n31678 ; n31678_not
g93472 not n31948 ; n31948_not
g93473 not n31939 ; n31939_not
g93474 not n38419 ; n38419_not
g93475 not n31894 ; n31894_not
g93476 not n37942 ; n37942_not
g93477 not n19843 ; n19843_not
g93478 not n31993 ; n31993_not
g93479 not n31975 ; n31975_not
g93480 not n19627 ; n19627_not
g93481 not n38239 ; n38239_not
g93482 not n31984 ; n31984_not
g93483 not n31687 ; n31687_not
g93484 not n31966 ; n31966_not
g93485 not n37933 ; n37933_not
g93486 not n32992 ; n32992_not
g93487 not n32695 ; n32695_not
g93488 not n32497 ; n32497_not
g93489 not n38329 ; n38329_not
g93490 not n32488 ; n32488_not
g93491 not n32479 ; n32479_not
g93492 not n38338 ; n38338_not
g93493 not n32668 ; n32668_not
g93494 not n38293 ; n38293_not
g93495 not n32569 ; n32569_not
g93496 not n32659 ; n32659_not
g93497 not n32677 ; n32677_not
g93498 not n32587 ; n32587_not
g93499 not n32398 ; n32398_not
g93500 not n32299 ; n32299_not
g93501 not n44593 ; n44593_not
g93502 not n38365 ; n38365_not
g93503 not n44575 ; n44575_not
g93504 not n38284 ; n38284_not
g93505 not n44584 ; n44584_not
g93506 not n19591 ; n19591_not
g93507 not n38374 ; n38374_not
g93508 not n38347 ; n38347_not
g93509 not n32389 ; n32389_not
g93510 not n38356 ; n38356_not
g93511 not n44557 ; n44557_not
g93512 not n37654 ; n37654_not
g93513 not n37663 ; n37663_not
g93514 not n33766 ; n33766_not
g93515 not n19726 ; n19726_not
g93516 not n33775 ; n33775_not
g93517 not n44098 ; n44098_not
g93518 not n44089 ; n44089_not
g93519 not n19780 ; n19780_not
g93520 not n33784 ; n33784_not
g93521 not n31759 ; n31759_not
g93522 not n38176 ; n38176_not
g93523 not n37690 ; n37690_not
g93524 not n38167 ; n38167_not
g93525 not n37681 ; n37681_not
g93526 not n38482 ; n38482_not
g93527 not n43792 ; n43792_not
g93528 not n38158 ; n38158_not
g93529 not n31696 ; n31696_not
g93530 not n33694 ; n33694_not
g93531 not n37672 ; n37672_not
g93532 not n19717 ; n19717_not
g93533 not n33388 ; n33388_not
g93534 not n38149 ; n38149_not
g93535 not n19744 ; n19744_not
g93536 not n30967 ; n30967_not
g93537 not n33829 ; n33829_not
g93538 not n38527 ; n38527_not
g93539 not n33838 ; n33838_not
g93540 not n19762 ; n19762_not
g93541 not n31597 ; n31597_not
g93542 not n19735 ; n19735_not
g93543 not n31588 ; n31588_not
g93544 not n43837 ; n43837_not
g93545 not n31579 ; n31579_not
g93546 not n31489 ; n31489_not
g93547 not n33793 ; n33793_not
g93548 not n19753 ; n19753_not
g93549 not n31498 ; n31498_not
g93550 not n31399 ; n31399_not
g93551 not n19654 ; n19654_not
g93552 not n38437 ; n38437_not
g93553 not n44296 ; n44296_not
g93554 not n37960 ; n37960_not
g93555 not n44287 ; n44287_not
g93556 not n19663 ; n19663_not
g93557 not n44386 ; n44386_not
g93558 not n32947 ; n32947_not
g93559 not n19645 ; n19645_not
g93560 not n33289 ; n33289_not
g93561 not n33379 ; n33379_not
g93562 not n38428 ; n38428_not
g93563 not n38194 ; n38194_not
g93564 not n31777 ; n31777_not
g93565 not n31786 ; n31786_not
g93566 not n44197 ; n44197_not
g93567 not n33649 ; n33649_not
g93568 not n19681 ; n19681_not
g93569 not n44188 ; n44188_not
g93570 not n44179 ; n44179_not
g93571 not n38185 ; n38185_not
g93572 not n19690 ; n19690_not
g93573 not n19708 ; n19708_not
g93574 not n31768 ; n31768_not
g93575 not n44278 ; n44278_not
g93576 not n44269 ; n44269_not
g93577 not n38446 ; n38446_not
g93578 not n33298 ; n33298_not
g93579 not n43747 ; n43747_not
g93580 not n19672 ; n19672_not
g93581 not n13678 ; n13678_not
g93582 not n41893 ; n41893_not
g93583 not n29572 ; n29572_not
g93584 not n37492 ; n37492_not
g93585 not n13948 ; n13948_not
g93586 not n42289 ; n42289_not
g93587 not n12688 ; n12688_not
g93588 not n29077 ; n29077_not
g93589 not n42919 ; n42919_not
g93590 not n29383 ; n29383_not
g93591 not n42298 ; n42298_not
g93592 not n12679 ; n12679_not
g93593 not n29275 ; n29275_not
g93594 not n42928 ; n42928_not
g93595 not n13966 ; n13966_not
g93596 not n29374 ; n29374_not
g93597 not n42694 ; n42694_not
g93598 not n13687 ; n13687_not
g93599 not n29473 ; n29473_not
g93600 not n42739 ; n42739_not
g93601 not n29563 ; n29563_not
g93602 not n12778 ; n12778_not
g93603 not n13669 ; n13669_not
g93604 not n29095 ; n29095_not
g93605 not n12769 ; n12769_not
g93606 not n41992 ; n41992_not
g93607 not n13894 ; n13894_not
g93608 not n42595 ; n42595_not
g93609 not n13489 ; n13489_not
g93610 not n34882 ; n34882_not
g93611 not n13498 ; n13498_not
g93612 not n13399 ; n13399_not
g93613 not n13939 ; n13939_not
g93614 not n29086 ; n29086_not
g93615 not n29482 ; n29482_not
g93616 not n42496 ; n42496_not
g93617 not n29392 ; n29392_not
g93618 not n41965 ; n41965_not
g93619 not n29248 ; n29248_not
g93620 not n42955 ; n42955_not
g93621 not n13759 ; n13759_not
g93622 not n42667 ; n42667_not
g93623 not n29329 ; n29329_not
g93624 not n42649 ; n42649_not
g93625 not n11986 ; n11986_not
g93626 not n42469 ; n42469_not
g93627 not n42658 ; n42658_not
g93628 not n41947 ; n41947_not
g93629 not n41938 ; n41938_not
g93630 not n28942 ; n28942_not
g93631 not n34909 ; n34909_not
g93632 not n42964 ; n42964_not
g93633 not n29617 ; n29617_not
g93634 not n13579 ; n13579_not
g93635 not n42937 ; n42937_not
g93636 not n29365 ; n29365_not
g93637 not n42685 ; n42685_not
g93638 not n13588 ; n13588_not
g93639 not n41983 ; n41983_not
g93640 not n29347 ; n29347_not
g93641 not n29338 ; n29338_not
g93642 not n12598 ; n12598_not
g93643 not n29068 ; n29068_not
g93644 not n13975 ; n13975_not
g93645 not n29581 ; n29581_not
g93646 not n42946 ; n42946_not
g93647 not n42676 ; n42676_not
g93648 not n29059 ; n29059_not
g93649 not n12589 ; n12589_not
g93650 not n13597 ; n13597_not
g93651 not n42199 ; n42199_not
g93652 not n42829 ; n42829_not
g93653 not n29437 ; n29437_not
g93654 not n42838 ; n42838_not
g93655 not n29464 ; n29464_not
g93656 not n29428 ; n29428_not
g93657 not n42847 ; n42847_not
g93658 not n42775 ; n42775_not
g93659 not n41956 ; n41956_not
g93660 not n42856 ; n42856_not
g93661 not n29419 ; n29419_not
g93662 not n29176 ; n29176_not
g93663 not n29509 ; n29509_not
g93664 not n29455 ; n29455_not
g93665 not n42793 ; n42793_not
g93666 not n29446 ; n29446_not
g93667 not n42784 ; n42784_not
g93668 not n29194 ; n29194_not
g93669 not n42559 ; n42559_not
g93670 not n29491 ; n29491_not
g93671 not n34837 ; n34837_not
g93672 not n29185 ; n29185_not
g93673 not n29545 ; n29545_not
g93674 not n13867 ; n13867_not
g93675 not n42748 ; n42748_not
g93676 not n29149 ; n29149_not
g93677 not n42883 ; n42883_not
g93678 not n12499 ; n12499_not
g93679 not n29554 ; n29554_not
g93680 not n34792 ; n34792_not
g93681 not n42586 ; n42586_not
g93682 not n42892 ; n42892_not
g93683 not n13876 ; n13876_not
g93684 not n19096 ; n19096_not
g93685 not n29518 ; n29518_not
g93686 not n42865 ; n42865_not
g93687 not n29527 ; n29527_not
g93688 not n13849 ; n13849_not
g93689 not n42766 ; n42766_not
g93690 not n42874 ; n42874_not
g93691 not n29158 ; n29158_not
g93692 not n29536 ; n29536_not
g93693 not n42757 ; n42757_not
g93694 not n12697 ; n12697_not
g93695 not n42379 ; n42379_not
g93696 not n42397 ; n42397_not
g93697 not n29608 ; n29608_not
g93698 not n42388 ; n42388_not
g93699 not n43279 ; n43279_not
g93700 not n13696 ; n13696_not
g93701 not n41848 ; n41848_not
g93702 not n41776 ; n41776_not
g93703 not n34738 ; n34738_not
g93704 not n21499 ; n21499_not
g93705 not n29644 ; n29644_not
g93706 not n28861 ; n28861_not
g93707 not n41767 ; n41767_not
g93708 not n41794 ; n41794_not
g93709 not n29284 ; n29284_not
g93710 not n11959 ; n11959_not
g93711 not n22795 ; n22795_not
g93712 not n34747 ; n34747_not
g93713 not n29806 ; n29806_not
g93714 not n29257 ; n29257_not
g93715 not n43297 ; n43297_not
g93716 not n41785 ; n41785_not
g93717 not n11968 ; n11968_not
g93718 not n28870 ; n28870_not
g93719 not n34684 ; n34684_not
g93720 not n43288 ; n43288_not
g93721 not n41866 ; n41866_not
g93722 not n13885 ; n13885_not
g93723 not n11878 ; n11878_not
g93724 not n34693 ; n34693_not
g93725 not n11887 ; n11887_not
g93726 not n11896 ; n11896_not
g93727 not n43189 ; n43189_not
g93728 not n11995 ; n11995_not
g93729 not n34729 ; n34729_not
g93730 not n34873 ; n34873_not
g93731 not n29734 ; n29734_not
g93732 not n41758 ; n41758_not
g93733 not n41749 ; n41749_not
g93734 not n43099 ; n43099_not
g93735 not n28852 ; n28852_not
g93736 not n11797 ; n11797_not
g93737 not n11869 ; n11869_not
g93738 not n28951 ; n28951_not
g93739 not n43378 ; n43378_not
g93740 not n13993 ; n13993_not
g93741 not n29293 ; n29293_not
g93742 not n42568 ; n42568_not
g93743 not n43369 ; n43369_not
g93744 not n41875 ; n41875_not
g93745 not n13984 ; n13984_not
g93746 not n29815 ; n29815_not
g93747 not n34666 ; n34666_not
g93748 not n43387 ; n43387_not
g93749 not n29635 ; n29635_not
g93750 not n29239 ; n29239_not
g93751 not n42973 ; n42973_not
g93752 not n34675 ; n34675_not
g93753 not n41695 ; n41695_not
g93754 not n42991 ; n42991_not
g93755 not n42478 ; n42478_not
g93756 not n37951 ; n37951_not
g93757 not n41857 ; n41857_not
g93758 not n19807 ; n19807_not
g93759 not n38608 ; n38608_not
g93760 not n28843 ; n28843_not
g93761 not n38563 ; n38563_not
g93762 not n42982 ; n42982_not
g93763 not n28915 ; n28915_not
g93764 not n36692 ; n36692_not
g93765 not n36809 ; n36809_not
g93766 not n22589 ; n22589_not
g93767 not n46826 ; n46826_not
g93768 not n52757 ; n52757_not
g93769 not n53495 ; n53495_not
g93770 not n53198 ; n53198_not
g93771 not n36683 ; n36683_not
g93772 not n46817 ; n46817_not
g93773 not n36782 ; n36782_not
g93774 not n47348 ; n47348_not
g93775 not n19691 ; n19691_not
g93776 not n37196 ; n37196_not
g93777 not n48086 ; n48086_not
g93778 not n52739 ; n52739_not
g93779 not n38195 ; n38195_not
g93780 not n36755 ; n36755_not
g93781 not n47375 ; n47375_not
g93782 not n48095 ; n48095_not
g93783 not n22499 ; n22499_not
g93784 not n19718 ; n19718_not
g93785 not n19709 ; n19709_not
g93786 not n36764 ; n36764_not
g93787 not n22949 ; n22949_not
g93788 not n20798 ; n20798_not
g93789 not n47366 ; n47366_not
g93790 not n21698 ; n21698_not
g93791 not n53486 ; n53486_not
g93792 not n36773 ; n36773_not
g93793 not n38186 ; n38186_not
g93794 not n52748 ; n52748_not
g93795 not n19808 ; n19808_not
g93796 not n21599 ; n21599_not
g93797 not n21689 ; n21689_not
g93798 not n22967 ; n22967_not
g93799 not n38159 ; n38159_not
g93800 not n47519 ; n47519_not
g93801 not n36719 ; n36719_not
g93802 not n48077 ; n48077_not
g93803 not n47393 ; n47393_not
g93804 not n37169 ; n37169_not
g93805 not n24596 ; n24596_not
g93806 not n47357 ; n47357_not
g93807 not n19682 ; n19682_not
g93808 not n36728 ; n36728_not
g93809 not n19727 ; n19727_not
g93810 not n47636 ; n47636_not
g93811 not n47627 ; n47627_not
g93812 not n38096 ; n38096_not
g93813 not n37178 ; n37178_not
g93814 not n46934 ; n46934_not
g93815 not n38168 ; n38168_not
g93816 not n36737 ; n36737_not
g93817 not n22958 ; n22958_not
g93818 not n36791 ; n36791_not
g93819 not n47186 ; n47186_not
g93820 not n37187 ; n37187_not
g93821 not n38177 ; n38177_not
g93822 not n21779 ; n21779_not
g93823 not n47384 ; n47384_not
g93824 not n36746 ; n36746_not
g93825 not n47177 ; n47177_not
g93826 not n36917 ; n36917_not
g93827 not n47591 ; n47591_not
g93828 not n47465 ; n47465_not
g93829 not n52685 ; n52685_not
g93830 not n22778 ; n22778_not
g93831 not n19619 ; n19619_not
g93832 not n22787 ; n22787_not
g93833 not n51965 ; n51965_not
g93834 not n38276 ; n38276_not
g93835 not n47168 ; n47168_not
g93836 not n36926 ; n36926_not
g93837 not n47555 ; n47555_not
g93838 not n51974 ; n51974_not
g93839 not n22598 ; n22598_not
g93840 not n46862 ; n46862_not
g93841 not n38069 ; n38069_not
g93842 not n38258 ; n38258_not
g93843 not n47546 ; n47546_not
g93844 not n36890 ; n36890_not
g93845 not n51929 ; n51929_not
g93846 not n48176 ; n48176_not
g93847 not n47456 ; n47456_not
g93848 not n38267 ; n38267_not
g93849 not n51938 ; n51938_not
g93850 not n36908 ; n36908_not
g93851 not n19844 ; n19844_not
g93852 not n51947 ; n51947_not
g93853 not n46853 ; n46853_not
g93854 not n51956 ; n51956_not
g93855 not n19628 ; n19628_not
g93856 not n22769 ; n22769_not
g93857 not n19853 ; n19853_not
g93858 not n48185 ; n48185_not
g93859 not n52667 ; n52667_not
g93860 not n22868 ; n22868_not
g93861 not n22697 ; n22697_not
g93862 not n19880 ; n19880_not
g93863 not n47483 ; n47483_not
g93864 not n37529 ; n37529_not
g93865 not n46880 ; n46880_not
g93866 not n47564 ; n47564_not
g93867 not n36944 ; n36944_not
g93868 not n47573 ; n47573_not
g93869 not n46871 ; n46871_not
g93870 not n19565 ; n19565_not
g93871 not n22859 ; n22859_not
g93872 not n53549 ; n53549_not
g93873 not n36953 ; n36953_not
g93874 not n24398 ; n24398_not
g93875 not n52658 ; n52658_not
g93876 not n19556 ; n19556_not
g93877 not n19592 ; n19592_not
g93878 not n48194 ; n48194_not
g93879 not n22796 ; n22796_not
g93880 not n47474 ; n47474_not
g93881 not n22886 ; n22886_not
g93882 not n36935 ; n36935_not
g93883 not n38285 ; n38285_not
g93884 not n47582 ; n47582_not
g93885 not n22679 ; n22679_not
g93886 not n22688 ; n22688_not
g93887 not n51983 ; n51983_not
g93888 not n19583 ; n19583_not
g93889 not n24479 ; n24479_not
g93890 not n51992 ; n51992_not
g93891 not n19574 ; n19574_not
g93892 not n52496 ; n52496_not
g93893 not n47528 ; n47528_not
g93894 not n46835 ; n46835_not
g93895 not n37088 ; n37088_not
g93896 not n19655 ; n19655_not
g93897 not n22994 ; n22994_not
g93898 not n53189 ; n53189_not
g93899 not n37493 ; n37493_not
g93900 not n37538 ; n37538_not
g93901 not n46916 ; n46916_not
g93902 not n48149 ; n48149_not
g93903 not n47609 ; n47609_not
g93904 not n37547 ; n37547_not
g93905 not n19673 ; n19673_not
g93906 not n46925 ; n46925_not
g93907 not n47618 ; n47618_not
g93908 not n19664 ; n19664_not
g93909 not n24569 ; n24569_not
g93910 not n48158 ; n48158_not
g93911 not n36854 ; n36854_not
g93912 not n47438 ; n47438_not
g93913 not n22976 ; n22976_not
g93914 not n52478 ; n52478_not
g93915 not n36863 ; n36863_not
g93916 not n47195 ; n47195_not
g93917 not n36872 ; n36872_not
g93918 not n38249 ; n38249_not
g93919 not n19637 ; n19637_not
g93920 not n36881 ; n36881_not
g93921 not n48167 ; n48167_not
g93922 not n47447 ; n47447_not
g93923 not n36818 ; n36818_not
g93924 not n47429 ; n47429_not
g93925 not n52487 ; n52487_not
g93926 not n36827 ; n36827_not
g93927 not n19835 ; n19835_not
g93928 not n47537 ; n47537_not
g93929 not n46844 ; n46844_not
g93930 not n19646 ; n19646_not
g93931 not n36836 ; n36836_not
g93932 not n46907 ; n46907_not
g93933 not n36845 ; n36845_not
g93934 not n23894 ; n23894_not
g93935 not n52964 ; n52964_not
g93936 not n37457 ; n37457_not
g93937 not n52577 ; n52577_not
g93938 not n23678 ; n23678_not
g93939 not n47096 ; n47096_not
g93940 not n23669 ; n23669_not
g93941 not n52955 ; n52955_not
g93942 not n52586 ; n52586_not
g93943 not n20987 ; n20987_not
g93944 not n52991 ; n52991_not
g93945 not n23984 ; n23984_not
g93946 not n20978 ; n20978_not
g93947 not n20969 ; n20969_not
g93948 not n47771 ; n47771_not
g93949 not n47078 ; n47078_not
g93950 not n47087 ; n47087_not
g93951 not n46664 ; n46664_not
g93952 not n52982 ; n52982_not
g93953 not n23993 ; n23993_not
g93954 not n52568 ; n52568_not
g93955 not n47780 ; n47780_not
g93956 not n52973 ; n52973_not
g93957 not n23768 ; n23768_not
g93958 not n47834 ; n47834_not
g93959 not n53288 ; n53288_not
g93960 not n46655 ; n46655_not
g93961 not n23759 ; n23759_not
g93962 not n23579 ; n23579_not
g93963 not n47843 ; n47843_not
g93964 not n52919 ; n52919_not
g93965 not n37583 ; n37583_not
g93966 not n46754 ; n46754_not
g93967 not n37574 ; n37574_not
g93968 not n52946 ; n52946_not
g93969 not n47807 ; n47807_not
g93970 not n52937 ; n52937_not
g93971 not n47816 ; n47816_not
g93972 not n37556 ; n37556_not
g93973 not n46763 ; n46763_not
g93974 not n23777 ; n23777_not
g93975 not n47681 ; n47681_not
g93976 not n23588 ; n23588_not
g93977 not n52928 ; n52928_not
g93978 not n20897 ; n20897_not
g93979 not n47717 ; n47717_not
g93980 not n46727 ; n46727_not
g93981 not n20888 ; n20888_not
g93982 not n20879 ; n20879_not
g93983 not n47726 ; n47726_not
g93984 not n23867 ; n23867_not
g93985 not n53378 ; n53378_not
g93986 not n23939 ; n23939_not
g93987 not n37952 ; n37952_not
g93988 not n47708 ; n47708_not
g93989 not n23849 ; n23849_not
g93990 not n23858 ; n23858_not
g93991 not n46709 ; n46709_not
g93992 not n37592 ; n37592_not
g93993 not n37970 ; n37970_not
g93994 not n20996 ; n20996_not
g93995 not n46718 ; n46718_not
g93996 not n37961 ; n37961_not
g93997 not n23786 ; n23786_not
g93998 not n23876 ; n23876_not
g93999 not n46691 ; n46691_not
g94000 not n47690 ; n47690_not
g94001 not n47753 ; n47753_not
g94002 not n23975 ; n23975_not
g94003 not n46673 ; n46673_not
g94004 not n37637 ; n37637_not
g94005 not n46745 ; n46745_not
g94006 not n37448 ; n37448_not
g94007 not n53396 ; n53396_not
g94008 not n37619 ; n37619_not
g94009 not n47762 ; n47762_not
g94010 not n47069 ; n47069_not
g94011 not n47735 ; n47735_not
g94012 not n46682 ; n46682_not
g94013 not n23948 ; n23948_not
g94014 not n46736 ; n46736_not
g94015 not n23957 ; n23957_not
g94016 not n23696 ; n23696_not
g94017 not n47744 ; n47744_not
g94018 not n37646 ; n37646_not
g94019 not n23966 ; n23966_not
g94020 not n52676 ; n52676_not
g94021 not n21977 ; n21977_not
g94022 not n47492 ; n47492_not
g94023 not n47258 ; n47258_not
g94024 not n23399 ; n23399_not
g94025 not n24686 ; n24686_not
g94026 not n52784 ; n52784_not
g94027 not n20699 ; n20699_not
g94028 not n37385 ; n37385_not
g94029 not n46952 ; n46952_not
g94030 not n47285 ; n47285_not
g94031 not n21968 ; n21968_not
g94032 not n37376 ; n37376_not
g94033 not n47645 ; n47645_not
g94034 not n19763 ; n19763_not
g94035 not n21959 ; n21959_not
g94036 not n36962 ; n36962_not
g94037 not n38078 ; n38078_not
g94038 not n24668 ; n24668_not
g94039 not n46790 ; n46790_not
g94040 not n46961 ; n46961_not
g94041 not n21995 ; n21995_not
g94042 not n21986 ; n21986_not
g94043 not n47654 ; n47654_not
g94044 not n22877 ; n22877_not
g94045 not n24695 ; n24695_not
g94046 not n37394 ; n37394_not
g94047 not n52793 ; n52793_not
g94048 not n21869 ; n21869_not
g94049 not n37286 ; n37286_not
g94050 not n21797 ; n21797_not
g94051 not n53099 ; n53099_not
g94052 not n37277 ; n37277_not
g94053 not n19745 ; n19745_not
g94054 not n37484 ; n37484_not
g94055 not n37268 ; n37268_not
g94056 not n19736 ; n19736_not
g94057 not n48059 ; n48059_not
g94058 not n37259 ; n37259_not
g94059 not n37079 ; n37079_not
g94060 not n19790 ; n19790_not
g94061 not n46943 ; n46943_not
g94062 not n21788 ; n21788_not
g94063 not n21896 ; n21896_not
g94064 not n37367 ; n37367_not
g94065 not n37358 ; n37358_not
g94066 not n52775 ; n52775_not
g94067 not n37349 ; n37349_not
g94068 not n21887 ; n21887_not
g94069 not n47267 ; n47267_not
g94070 not n46808 ; n46808_not
g94071 not n21878 ; n21878_not
g94072 not n52766 ; n52766_not
g94073 not n24659 ; n24659_not
g94074 not n37295 ; n37295_not
g94075 not n53468 ; n53468_not
g94076 not n52865 ; n52865_not
g94077 not n23498 ; n23498_not
g94078 not n24299 ; n24299_not
g94079 not n52856 ; n52856_not
g94080 not n46772 ; n46772_not
g94081 not n47276 ; n47276_not
g94082 not n47906 ; n47906_not
g94083 not n52847 ; n52847_not
g94084 not n47672 ; n47672_not
g94085 not n47861 ; n47861_not
g94086 not n52892 ; n52892_not
g94087 not n52883 ; n52883_not
g94088 not n23687 ; n23687_not
g94089 not n52874 ; n52874_not
g94090 not n47924 ; n47924_not
g94091 not n47933 ; n47933_not
g94092 not n24389 ; n24389_not
g94093 not n52829 ; n52829_not
g94094 not n36980 ; n36980_not
g94095 not n24488 ; n24488_not
g94096 not n24578 ; n24578_not
g94097 not n47951 ; n47951_not
g94098 not n46970 ; n46970_not
g94099 not n47663 ; n47663_not
g94100 not n37466 ; n37466_not
g94101 not n23489 ; n23489_not
g94102 not n52838 ; n52838_not
g94103 not n46781 ; n46781_not
g94104 not n49463 ; n49463_not
g94105 not n34919 ; n34919_not
g94106 not n49571 ; n49571_not
g94107 not n29267 ; n29267_not
g94108 not n34937 ; n34937_not
g94109 not n29249 ; n29249_not
g94110 not n34928 ; n34928_not
g94111 not n29186 ; n29186_not
g94112 not n29159 ; n29159_not
g94113 not n34874 ; n34874_not
g94114 not n29375 ; n29375_not
g94115 not n29393 ; n29393_not
g94116 not n49445 ; n49445_not
g94117 not n34892 ; n34892_not
g94118 not n29357 ; n29357_not
g94119 not n29339 ; n29339_not
g94120 not n29258 ; n29258_not
g94121 not n29294 ; n29294_not
g94122 not n49454 ; n49454_not
g94123 not n29285 ; n29285_not
g94124 not n29195 ; n29195_not
g94125 not n28970 ; n28970_not
g94126 not n51299 ; n51299_not
g94127 not n28952 ; n28952_not
g94128 not n50993 ; n50993_not
g94129 not n49508 ; n49508_not
g94130 not n34883 ; n34883_not
g94131 not n28943 ; n28943_not
g94132 not n28934 ; n28934_not
g94133 not n50984 ; n50984_not
g94134 not n28097 ; n28097_not
g94135 not n29168 ; n29168_not
g94136 not n29078 ; n29078_not
g94137 not n29087 ; n29087_not
g94138 not n49490 ; n49490_not
g94139 not n29096 ; n29096_not
g94140 not n29069 ; n29069_not
g94141 not n29735 ; n29735_not
g94142 not n29726 ; n29726_not
g94143 not n29717 ; n29717_not
g94144 not n49373 ; n49373_not
g94145 not n29708 ; n29708_not
g94146 not n34379 ; n34379_not
g94147 not n29609 ; n29609_not
g94148 not n29618 ; n29618_not
g94149 not n29690 ; n29690_not
g94150 not n29681 ; n29681_not
g94151 not n34757 ; n34757_not
g94152 not n34766 ; n34766_not
g94153 not n29672 ; n29672_not
g94154 not n29663 ; n29663_not
g94155 not n50399 ; n50399_not
g94156 not n50588 ; n50588_not
g94157 not n34298 ; n34298_not
g94158 not n50966 ; n50966_not
g94159 not n50579 ; n50579_not
g94160 not n29807 ; n29807_not
g94161 not n49355 ; n49355_not
g94162 not n29645 ; n29645_not
g94163 not n29771 ; n29771_not
g94164 not n29762 ; n29762_not
g94165 not n50498 ; n50498_not
g94166 not n50489 ; n50489_not
g94167 not n29744 ; n29744_not
g94168 not n49364 ; n49364_not
g94169 not n29537 ; n29537_not
g94170 not n49409 ; n49409_not
g94171 not n29528 ; n29528_not
g94172 not n29519 ; n29519_not
g94173 not n49418 ; n49418_not
g94174 not n34829 ; n34829_not
g94175 not n34847 ; n34847_not
g94176 not n29483 ; n29483_not
g94177 not n29474 ; n29474_not
g94178 not n29465 ; n29465_not
g94179 not n34865 ; n34865_not
g94180 not n29348 ; n29348_not
g94181 not n29654 ; n29654_not
g94182 not n29627 ; n29627_not
g94183 not n49580 ; n49580_not
g94184 not n29582 ; n29582_not
g94185 not n34775 ; n34775_not
g94186 not n29573 ; n29573_not
g94187 not n34784 ; n34784_not
g94188 not n29564 ; n29564_not
g94189 not n29555 ; n29555_not
g94190 not n29492 ; n29492_not
g94191 not n29546 ; n29546_not
g94192 not n51578 ; n51578_not
g94193 not n49427 ; n49427_not
g94194 not n50849 ; n50849_not
g94195 not n51587 ; n51587_not
g94196 not n28475 ; n28475_not
g94197 not n35189 ; n35189_not
g94198 not n35198 ; n35198_not
g94199 not n35288 ; n35288_not
g94200 not n35297 ; n35297_not
g94201 not n27854 ; n27854_not
g94202 not n49472 ; n49472_not
g94203 not n27890 ; n27890_not
g94204 not n50867 ; n50867_not
g94205 not n28529 ; n28529_not
g94206 not n50858 ; n50858_not
g94207 not n27881 ; n27881_not
g94208 not n51569 ; n51569_not
g94209 not n28493 ; n28493_not
g94210 not n34793 ; n34793_not
g94211 not n35396 ; n35396_not
g94212 not n27773 ; n27773_not
g94213 not n27809 ; n27809_not
g94214 not n49319 ; n49319_not
g94215 not n27836 ; n27836_not
g94216 not n35459 ; n35459_not
g94217 not n28295 ; n28295_not
g94218 not n35468 ; n35468_not
g94219 not n49292 ; n49292_not
g94220 not n27845 ; n27845_not
g94221 not n35477 ; n35477_not
g94222 not n35486 ; n35486_not
g94223 not n28277 ; n28277_not
g94224 not n48815 ; n48815_not
g94225 not n48536 ; n48536_not
g94226 not n35495 ; n35495_not
g94227 not n28268 ; n28268_not
g94228 not n51596 ; n51596_not
g94229 not n28457 ; n28457_not
g94230 not n49382 ; n49382_not
g94231 not n28439 ; n28439_not
g94232 not n28385 ; n28385_not
g94233 not n28367 ; n28367_not
g94234 not n35369 ; n35369_not
g94235 not n27791 ; n27791_not
g94236 not n35378 ; n35378_not
g94237 not n35387 ; n35387_not
g94238 not n49337 ; n49337_not
g94239 not n28349 ; n28349_not
g94240 not n28781 ; n28781_not
g94241 not n49544 ; n49544_not
g94242 not n50939 ; n50939_not
g94243 not n28763 ; n28763_not
g94244 not n49553 ; n49553_not
g94245 not n28745 ; n28745_not
g94246 not n28727 ; n28727_not
g94247 not n48824 ; n48824_not
g94248 not n28709 ; n28709_not
g94249 not n28871 ; n28871_not
g94250 not n28853 ; n28853_not
g94251 not n51389 ; n51389_not
g94252 not n28835 ; n28835_not
g94253 not n49535 ; n49535_not
g94254 not n50957 ; n50957_not
g94255 not n51398 ; n51398_not
g94256 not n28817 ; n28817_not
g94257 not n50948 ; n50948_not
g94258 not n50894 ; n50894_not
g94259 not n34838 ; n34838_not
g94260 not n28637 ; n28637_not
g94261 not n49517 ; n49517_not
g94262 not n27944 ; n27944_not
g94263 not n28619 ; n28619_not
g94264 not n28583 ; n28583_not
g94265 not n28565 ; n28565_not
g94266 not n28547 ; n28547_not
g94267 not n27980 ; n27980_not
g94268 not n48833 ; n48833_not
g94269 not n28691 ; n28691_not
g94270 not n49562 ; n49562_not
g94271 not n27971 ; n27971_not
g94272 not n51479 ; n51479_not
g94273 not n28673 ; n28673_not
g94274 not n51488 ; n51488_not
g94275 not n28655 ; n28655_not
g94276 not n51497 ; n51497_not
g94277 not n33479 ; n33479_not
g94278 not n49841 ; n49841_not
g94279 not n33488 ; n33488_not
g94280 not n31769 ; n31769_not
g94281 not n33497 ; n33497_not
g94282 not n31787 ; n31787_not
g94283 not n31778 ; n31778_not
g94284 not n50597 ; n50597_not
g94285 not n33299 ; n33299_not
g94286 not n33569 ; n33569_not
g94287 not n33578 ; n33578_not
g94288 not n33587 ; n33587_not
g94289 not n33596 ; n33596_not
g94290 not n49850 ; n49850_not
g94291 not n31796 ; n31796_not
g94292 not n49814 ; n49814_not
g94293 not n31688 ; n31688_not
g94294 not n49634 ; n49634_not
g94295 not n32984 ; n32984_not
g94296 not n31697 ; n31697_not
g94297 not n49823 ; n49823_not
g94298 not n49625 ; n49625_not
g94299 not n32957 ; n32957_not
g94300 not n32948 ; n32948_not
g94301 not n32939 ; n32939_not
g94302 not n49616 ; n49616_not
g94303 not n33389 ; n33389_not
g94304 not n33398 ; n33398_not
g94305 not n49832 ; n49832_not
g94306 not n31598 ; n31598_not
g94307 not n31589 ; n31589_not
g94308 not n49607 ; n49607_not
g94309 not n33767 ; n33767_not
g94310 not n49643 ; n49643_not
g94311 not n31679 ; n31679_not
g94312 not n33776 ; n33776_not
g94313 not n49652 ; n49652_not
g94314 not n33785 ; n33785_not
g94315 not n49661 ; n49661_not
g94316 not n49670 ; n49670_not
g94317 not n31499 ; n31499_not
g94318 not n33659 ; n33659_not
g94319 not n33677 ; n33677_not
g94320 not n33686 ; n33686_not
g94321 not n32768 ; n32768_not
g94322 not n49706 ; n49706_not
g94323 not n49751 ; n49751_not
g94324 not n32399 ; n32399_not
g94325 not n32777 ; n32777_not
g94326 not n32786 ; n32786_not
g94327 not n31985 ; n31985_not
g94328 not n32795 ; n32795_not
g94329 not n31994 ; n31994_not
g94330 not n49760 ; n49760_not
g94331 not n32489 ; n32489_not
g94332 not n31967 ; n31967_not
g94333 not n32498 ; n32498_not
g94334 not n31958 ; n31958_not
g94335 not n31949 ; n31949_not
g94336 not n32849 ; n32849_not
g94337 not n32858 ; n32858_not
g94338 not n32867 ; n32867_not
g94339 not n31895 ; n31895_not
g94340 not n49733 ; n49733_not
g94341 not n32579 ; n32579_not
g94342 not n32597 ; n32597_not
g94343 not n32669 ; n32669_not
g94344 not n49724 ; n49724_not
g94345 not n32687 ; n32687_not
g94346 not n32588 ; n32588_not
g94347 not n32696 ; n32696_not
g94348 not n49715 ; n49715_not
g94349 not n49742 ; n49742_not
g94350 not n32678 ; n32678_not
g94351 not n32759 ; n32759_not
g94352 not n31886 ; n31886_not
g94353 not n32966 ; n32966_not
g94354 not n32993 ; n32993_not
g94355 not n49805 ; n49805_not
g94356 not n31976 ; n31976_not
g94357 not n32876 ; n32876_not
g94358 not n31877 ; n31877_not
g94359 not n32885 ; n32885_not
g94360 not n31868 ; n31868_not
g94361 not n32894 ; n32894_not
g94362 not n31859 ; n31859_not
g94363 not n29960 ; n29960_not
g94364 not n34199 ; n34199_not
g94365 not n29942 ; n29942_not
g94366 not n29933 ; n29933_not
g94367 not n50795 ; n50795_not
g94368 not n50786 ; n50786_not
g94369 not n34289 ; n34289_not
g94370 not n50777 ; n50777_not
g94371 not n50768 ; n50768_not
g94372 not n50759 ; n50759_not
g94373 not n33992 ; n33992_not
g94374 not n34388 ; n34388_not
g94375 not n49931 ; n49931_not
g94376 not n30869 ; n30869_not
g94377 not n49940 ; n49940_not
g94378 not n33983 ; n33983_not
g94379 not n30797 ; n30797_not
g94380 not n30788 ; n30788_not
g94381 not n30779 ; n30779_not
g94382 not n30698 ; n30698_not
g94383 not n30689 ; n30689_not
g94384 not n29906 ; n29906_not
g94385 not n29951 ; n29951_not
g94386 not n50687 ; n50687_not
g94387 not n50678 ; n50678_not
g94388 not n29861 ; n29861_not
g94389 not n50669 ; n50669_not
g94390 not n29852 ; n29852_not
g94391 not n29843 ; n29843_not
g94392 not n29834 ; n29834_not
g94393 not n29825 ; n29825_not
g94394 not n29780 ; n29780_not
g94395 not n29816 ; n29816_not
g94396 not n34478 ; n34478_not
g94397 not n34496 ; n34496_not
g94398 not n50876 ; n50876_not
g94399 not n29915 ; n29915_not
g94400 not n34469 ; n34469_not
g94401 not n50696 ; n50696_not
g94402 not n49328 ; n49328_not
g94403 not n29870 ; n29870_not
g94404 not n33866 ; n33866_not
g94405 not n49922 ; n49922_not
g94406 not n33875 ; n33875_not
g94407 not n30995 ; n30995_not
g94408 not n30986 ; n30986_not
g94409 not n33884 ; n33884_not
g94410 not n33893 ; n33893_not
g94411 not n33794 ; n33794_not
g94412 not n30959 ; n30959_not
g94413 not n49904 ; n49904_not
g94414 not n30968 ; n30968_not
g94415 not n30977 ; n30977_not
g94416 not n33695 ; n33695_not
g94417 not n33839 ; n33839_not
g94418 not n49913 ; n49913_not
g94419 not n33848 ; n33848_not
g94420 not n33857 ; n33857_not
g94421 not n33965 ; n33965_not
g94422 not n30878 ; n30878_not
g94423 not n33974 ; n33974_not
g94424 not n30887 ; n30887_not
g94425 not n30896 ; n30896_not
g94426 not n33929 ; n33929_not
g94427 not n33938 ; n33938_not
g94428 not n33947 ; n33947_not
g94429 not n33956 ; n33956_not
g94430 not n26378 ; n26378_not
g94431 not n26495 ; n26495_not
g94432 not n48572 ; n48572_not
g94433 not n26297 ; n26297_not
g94434 not n26486 ; n26486_not
g94435 not n48563 ; n48563_not
g94436 not n26477 ; n26477_not
g94437 not n26468 ; n26468_not
g94438 not n36674 ; n36674_not
g94439 not n26459 ; n26459_not
g94440 not n26576 ; n26576_not
g94441 not n48608 ; n48608_not
g94442 not n36629 ; n36629_not
g94443 not n36638 ; n36638_not
g94444 not n51677 ; n51677_not
g94445 not n36656 ; n36656_not
g94446 not n26567 ; n26567_not
g94447 not n26558 ; n26558_not
g94448 not n48590 ; n48590_not
g94449 not n26549 ; n26549_not
g94450 not n51668 ; n51668_not
g94451 not n48518 ; n48518_not
g94452 not n52388 ; n52388_not
g94453 not n36287 ; n36287_not
g94454 not n26369 ; n26369_not
g94455 not n48509 ; n48509_not
g94456 not n36296 ; n36296_not
g94457 not n52397 ; n52397_not
g94458 not n26279 ; n26279_not
g94459 not n48491 ; n48491_not
g94460 not n48545 ; n48545_not
g94461 not n52379 ; n52379_not
g94462 not n26396 ; n26396_not
g94463 not n26387 ; n26387_not
g94464 not n36269 ; n36269_not
g94465 not n36647 ; n36647_not
g94466 not n36278 ; n36278_not
g94467 not n26774 ; n26774_not
g94468 not n48725 ; n48725_not
g94469 not n26765 ; n26765_not
g94470 not n26756 ; n26756_not
g94471 not n36089 ; n36089_not
g94472 not n26747 ; n26747_not
g94473 not n26738 ; n26738_not
g94474 not n36449 ; n36449_not
g94475 not n48707 ; n48707_not
g94476 not n36458 ; n36458_not
g94477 not n36467 ; n36467_not
g94478 not n36476 ; n36476_not
g94479 not n36485 ; n36485_not
g94480 not n26729 ; n26729_not
g94481 not n26837 ; n26837_not
g94482 not n48752 ; n48752_not
g94483 not n36359 ; n36359_not
g94484 not n36368 ; n36368_not
g94485 not n26828 ; n26828_not
g94486 not n48743 ; n48743_not
g94487 not n26819 ; n26819_not
g94488 not n36377 ; n36377_not
g94489 not n36386 ; n36386_not
g94490 not n26792 ; n26792_not
g94491 not n36395 ; n36395_not
g94492 not n26783 ; n26783_not
g94493 not n36098 ; n36098_not
g94494 not n52298 ; n52298_not
g94495 not n48653 ; n48653_not
g94496 not n26648 ; n26648_not
g94497 not n36566 ; n36566_not
g94498 not n26639 ; n26639_not
g94499 not n48635 ; n48635_not
g94500 not n36584 ; n36584_not
g94501 not n26594 ; n26594_not
g94502 not n51686 ; n51686_not
g94503 not n26585 ; n26585_not
g94504 not n36593 ; n36593_not
g94505 not n48617 ; n48617_not
g94506 not n36494 ; n36494_not
g94507 not n26693 ; n26693_not
g94508 not n26684 ; n26684_not
g94509 not n26675 ; n26675_not
g94510 not n48680 ; n48680_not
g94511 not n52289 ; n52289_not
g94512 not n26666 ; n26666_not
g94513 not n26657 ; n26657_not
g94514 not n48662 ; n48662_not
g94515 not n36539 ; n36539_not
g94516 not n36548 ; n36548_not
g94517 not n48329 ; n48329_not
g94518 not n36557 ; n36557_not
g94519 not n25586 ; n25586_not
g94520 not n25577 ; n25577_not
g94521 not n25496 ; n25496_not
g94522 not n52595 ; n52595_not
g94523 not n25568 ; n25568_not
g94524 not n48365 ; n48365_not
g94525 not n25685 ; n25685_not
g94526 not n52199 ; n52199_not
g94527 not n25676 ; n25676_not
g94528 not n48356 ; n48356_not
g94529 not n25667 ; n25667_not
g94530 not n25658 ; n25658_not
g94531 not n48347 ; n48347_not
g94532 not n25649 ; n25649_not
g94533 not n48338 ; n48338_not
g94534 not n25469 ; n25469_not
g94535 not n25595 ; n25595_not
g94536 not n48257 ; n48257_not
g94537 not n48248 ; n48248_not
g94538 not n48239 ; n48239_not
g94539 not n36971 ; n36971_not
g94540 not n25388 ; n25388_not
g94541 not n25298 ; n25298_not
g94542 not n25559 ; n25559_not
g94543 not n48293 ; n48293_not
g94544 not n48284 ; n48284_not
g94545 not n47942 ; n47942_not
g94546 not n48275 ; n48275_not
g94547 not n48266 ; n48266_not
g94548 not n25478 ; n25478_not
g94549 not n25289 ; n25289_not
g94550 not n25946 ; n25946_not
g94551 not n48455 ; n48455_not
g94552 not n25937 ; n25937_not
g94553 not n25928 ; n25928_not
g94554 not n48446 ; n48446_not
g94555 not n25919 ; n25919_not
g94556 not n47852 ; n47852_not
g94557 not n25892 ; n25892_not
g94558 not n25883 ; n25883_not
g94559 not n48437 ; n48437_not
g94560 not n25874 ; n25874_not
g94561 not n26189 ; n26189_not
g94562 not n26099 ; n26099_not
g94563 not n48482 ; n48482_not
g94564 not n25991 ; n25991_not
g94565 not n25982 ; n25982_not
g94566 not n48473 ; n48473_not
g94567 not n25973 ; n25973_not
g94568 not n48464 ; n48464_not
g94569 not n25964 ; n25964_not
g94570 not n25955 ; n25955_not
g94571 not n25793 ; n25793_not
g94572 not n25379 ; n25379_not
g94573 not n25784 ; n25784_not
g94574 not n48392 ; n48392_not
g94575 not n25775 ; n25775_not
g94576 not n25766 ; n25766_not
g94577 not n48383 ; n48383_not
g94578 not n25757 ; n25757_not
g94579 not n25748 ; n25748_not
g94580 not n48374 ; n48374_not
g94581 not n25739 ; n25739_not
g94582 not n25694 ; n25694_not
g94583 not n48428 ; n48428_not
g94584 not n25865 ; n25865_not
g94585 not n48419 ; n48419_not
g94586 not n25856 ; n25856_not
g94587 not n25847 ; n25847_not
g94588 not n25838 ; n25838_not
g94589 not n25829 ; n25829_not
g94590 not n27638 ; n27638_not
g94591 not n35882 ; n35882_not
g94592 not n27647 ; n27647_not
g94593 not n27656 ; n27656_not
g94594 not n35693 ; n35693_not
g94595 not n27665 ; n27665_not
g94596 not n35891 ; n35891_not
g94597 not n27674 ; n27674_not
g94598 not n27683 ; n27683_not
g94599 not n27692 ; n27692_not
g94600 not n27818 ; n27818_not
g94601 not n27719 ; n27719_not
g94602 not n27728 ; n27728_not
g94603 not n27737 ; n27737_not
g94604 not n27539 ; n27539_not
g94605 not n27548 ; n27548_not
g94606 not n27908 ; n27908_not
g94607 not n27557 ; n27557_not
g94608 not n35855 ; n35855_not
g94609 not n48626 ; n48626_not
g94610 not n27566 ; n27566_not
g94611 not n27575 ; n27575_not
g94612 not n35864 ; n35864_not
g94613 not n27584 ; n27584_not
g94614 not n27593 ; n27593_not
g94615 not n35873 ; n35873_not
g94616 not n27629 ; n27629_not
g94617 not n27863 ; n27863_not
g94618 not n35666 ; n35666_not
g94619 not n27764 ; n27764_not
g94620 not n35945 ; n35945_not
g94621 not n26909 ; n26909_not
g94622 not n27755 ; n27755_not
g94623 not n26927 ; n26927_not
g94624 not n27746 ; n27746_not
g94625 not n35657 ; n35657_not
g94626 not n35954 ; n35954_not
g94627 not n26936 ; n26936_not
g94628 not n51893 ; n51893_not
g94629 not n35963 ; n35963_not
g94630 not n26945 ; n26945_not
g94631 not n35648 ; n35648_not
g94632 not n35909 ; n35909_not
g94633 not n51848 ; n51848_not
g94634 not n35918 ; n35918_not
g94635 not n51857 ; n51857_not
g94636 not n35927 ; n35927_not
g94637 not n27782 ; n27782_not
g94638 not n35936 ; n35936_not
g94639 not n51875 ; n51875_not
g94640 not n48671 ; n48671_not
g94641 not n35675 ; n35675_not
g94642 not n28196 ; n28196_not
g94643 not n28187 ; n28187_not
g94644 not n28178 ; n28178_not
g94645 not n28079 ; n28079_not
g94646 not n35738 ; n35738_not
g94647 not n35747 ; n35747_not
g94648 not n48581 ; n48581_not
g94649 not n35765 ; n35765_not
g94650 not n27269 ; n27269_not
g94651 not n28259 ; n28259_not
g94652 not n35549 ; n35549_not
g94653 not n35558 ; n35558_not
g94654 not n35567 ; n35567_not
g94655 not n35576 ; n35576_not
g94656 not n35585 ; n35585_not
g94657 not n27926 ; n27926_not
g94658 not n35594 ; n35594_not
g94659 not n27935 ; n27935_not
g94660 not n51695 ; n51695_not
g94661 not n27458 ; n27458_not
g94662 not n51767 ; n51767_not
g94663 not n27467 ; n27467_not
g94664 not n27953 ; n27953_not
g94665 not n27476 ; n27476_not
g94666 not n27485 ; n27485_not
g94667 not n35819 ; n35819_not
g94668 not n27494 ; n27494_not
g94669 not n35828 ; n35828_not
g94670 not n35837 ; n35837_not
g94671 not n51785 ; n51785_not
g94672 not n35846 ; n35846_not
g94673 not n27278 ; n27278_not
g94674 not n27287 ; n27287_not
g94675 not n35774 ; n35774_not
g94676 not n27296 ; n27296_not
g94677 not n27359 ; n27359_not
g94678 not n27368 ; n27368_not
g94679 not n27377 ; n27377_not
g94680 not n27386 ; n27386_not
g94681 not n35756 ; n35756_not
g94682 not n35783 ; n35783_not
g94683 not n27395 ; n27395_not
g94684 not n27449 ; n27449_not
g94685 not n51758 ; n51758_not
g94686 not n35792 ; n35792_not
g94687 not n36188 ; n36188_not
g94688 not n26981 ; n26981_not
g94689 not n26972 ; n26972_not
g94690 not n27089 ; n27089_not
g94691 not n36179 ; n36179_not
g94692 not n26891 ; n26891_not
g94693 not n26882 ; n26882_not
g94694 not n48770 ; n48770_not
g94695 not n26873 ; n26873_not
g94696 not n26864 ; n26864_not
g94697 not n26855 ; n26855_not
g94698 not n26846 ; n26846_not
g94699 not n36197 ; n36197_not
g94700 not n26954 ; n26954_not
g94701 not n51776 ; n51776_not
g94702 not n26918 ; n26918_not
g94703 not n48716 ; n48716_not
g94704 not n51866 ; n51866_not
g94705 not n35972 ; n35972_not
g94706 not n35981 ; n35981_not
g94707 not n35990 ; n35990_not
g94708 not n26990 ; n26990_not
g94709 not n27197 ; n27197_not
g94710 not n27179 ; n27179_not
g94711 not n48761 ; n48761_not
g94712 not n14579 ; n14579_not
g94713 not n17738 ; n17738_not
g94714 not n40697 ; n40697_not
g94715 not n39428 ; n39428_not
g94716 not n46376 ; n46376_not
g94717 not n45458 ; n45458_not
g94718 not n17729 ; n17729_not
g94719 not n46367 ; n46367_not
g94720 not n39419 ; n39419_not
g94721 not n46385 ; n46385_not
g94722 not n18179 ; n18179_not
g94723 not n18188 ; n18188_not
g94724 not n55709 ; n55709_not
g94725 not n14588 ; n14588_not
g94726 not n40994 ; n40994_not
g94727 not n18197 ; n18197_not
g94728 not n17693 ; n17693_not
g94729 not n45449 ; n45449_not
g94730 not n40985 ; n40985_not
g94731 not n55718 ; n55718_not
g94732 not n17684 ; n17684_not
g94733 not n40976 ; n40976_not
g94734 not n40967 ; n40967_not
g94735 not n45674 ; n45674_not
g94736 not n45935 ; n45935_not
g94737 not n39455 ; n39455_not
g94738 not n46358 ; n46358_not
g94739 not n55673 ; n55673_not
g94740 not n45476 ; n45476_not
g94741 not n14669 ; n14669_not
g94742 not n55682 ; n55682_not
g94743 not n39446 ; n39446_not
g94744 not n18089 ; n18089_not
g94745 not n54980 ; n54980_not
g94746 not n45467 ; n45467_not
g94747 not n55691 ; n55691_not
g94748 not n18098 ; n18098_not
g94749 not n39437 ; n39437_not
g94750 not n39068 ; n39068_not
g94751 not n13679 ; n13679_not
g94752 not n54953 ; n54953_not
g94753 not n18296 ; n18296_not
g94754 not n55745 ; n55745_not
g94755 not n13787 ; n13787_not
g94756 not n41579 ; n41579_not
g94757 not n39356 ; n39356_not
g94758 not n41588 ; n41588_not
g94759 not n41597 ; n41597_not
g94760 not n54944 ; n54944_not
g94761 not n55754 ; n55754_not
g94762 not n39347 ; n39347_not
g94763 not n13796 ; n13796_not
g94764 not n13598 ; n13598_not
g94765 not n18359 ; n18359_not
g94766 not n13589 ; n13589_not
g94767 not n46448 ; n46448_not
g94768 not n39338 ; n39338_not
g94769 not n55763 ; n55763_not
g94770 not n41669 ; n41669_not
g94771 not n18377 ; n18377_not
g94772 not n41678 ; n41678_not
g94773 not n54935 ; n54935_not
g94774 not n46457 ; n46457_not
g94775 not n39329 ; n39329_not
g94776 not n55772 ; n55772_not
g94777 not n54269 ; n54269_not
g94778 not n17675 ; n17675_not
g94779 not n40958 ; n40958_not
g94780 not n39392 ; n39392_not
g94781 not n40949 ; n40949_not
g94782 not n40895 ; n40895_not
g94783 not n40886 ; n40886_not
g94784 not n40877 ; n40877_not
g94785 not n39383 ; n39383_not
g94786 not n18269 ; n18269_not
g94787 not n40859 ; n40859_not
g94788 not n18278 ; n18278_not
g94789 not n55727 ; n55727_not
g94790 not n17648 ; n17648_not
g94791 not n14489 ; n14489_not
g94792 not n14399 ; n14399_not
g94793 not n39374 ; n39374_not
g94794 not n13697 ; n13697_not
g94795 not n39059 ; n39059_not
g94796 not n41489 ; n41489_not
g94797 not n18287 ; n18287_not
g94798 not n41498 ; n41498_not
g94799 not n17639 ; n17639_not
g94800 not n55736 ; n55736_not
g94801 not n13688 ; n13688_not
g94802 not n39365 ; n39365_not
g94803 not n39527 ; n39527_not
g94804 not n46286 ; n46286_not
g94805 not n17855 ; n17855_not
g94806 not n17909 ; n17909_not
g94807 not n55619 ; n55619_not
g94808 not n17918 ; n17918_not
g94809 not n46295 ; n46295_not
g94810 not n45548 ; n45548_not
g94811 not n14795 ; n14795_not
g94812 not n39509 ; n39509_not
g94813 not n14786 ; n14786_not
g94814 not n45719 ; n45719_not
g94815 not n55628 ; n55628_not
g94816 not n17927 ; n17927_not
g94817 not n14777 ; n14777_not
g94818 not n17936 ; n17936_not
g94819 not n45539 ; n45539_not
g94820 not n54179 ; n54179_not
g94821 not n55592 ; n55592_not
g94822 not n45575 ; n45575_not
g94823 not n17189 ; n17189_not
g94824 not n39554 ; n39554_not
g94825 not n17873 ; n17873_not
g94826 not n46268 ; n46268_not
g94827 not n14885 ; n14885_not
g94828 not n14876 ; n14876_not
g94829 not n17864 ; n17864_not
g94830 not n45566 ; n45566_not
g94831 not n17891 ; n17891_not
g94832 not n14867 ; n14867_not
g94833 not n46277 ; n46277_not
g94834 not n14858 ; n14858_not
g94835 not n14849 ; n14849_not
g94836 not n39536 ; n39536_not
g94837 not n45557 ; n45557_not
g94838 not n55646 ; n55646_not
g94839 not n39473 ; n39473_not
g94840 not n55655 ; n55655_not
g94841 not n14696 ; n14696_not
g94842 not n40796 ; n40796_not
g94843 not n17783 ; n17783_not
g94844 not n14687 ; n14687_not
g94845 not n55664 ; n55664_not
g94846 not n39464 ; n39464_not
g94847 not n45494 ; n45494_not
g94848 not n40787 ; n40787_not
g94849 not n17774 ; n17774_not
g94850 not n46349 ; n46349_not
g94851 not n45485 ; n45485_not
g94852 not n14678 ; n14678_not
g94853 not n17765 ; n17765_not
g94854 not n14768 ; n14768_not
g94855 not n14759 ; n14759_not
g94856 not n17945 ; n17945_not
g94857 not n55637 ; n55637_not
g94858 not n40679 ; n40679_not
g94859 not n17954 ; n17954_not
g94860 not n39491 ; n39491_not
g94861 not n40769 ; n40769_not
g94862 not n17828 ; n17828_not
g94863 not n17963 ; n17963_not
g94864 not n17819 ; n17819_not
g94865 not n17972 ; n17972_not
g94866 not n39482 ; n39482_not
g94867 not n17981 ; n17981_not
g94868 not n17990 ; n17990_not
g94869 not n12896 ; n12896_not
g94870 not n39149 ; n39149_not
g94871 not n42848 ; n42848_not
g94872 not n42857 ; n42857_not
g94873 not n45197 ; n45197_not
g94874 not n12887 ; n12887_not
g94875 not n42866 ; n42866_not
g94876 not n12878 ; n12878_not
g94877 not n12689 ; n12689_not
g94878 not n42875 ; n42875_not
g94879 not n12869 ; n12869_not
g94880 not n12698 ; n12698_not
g94881 not n42884 ; n42884_not
g94882 not n12797 ; n12797_not
g94883 not n12788 ; n12788_not
g94884 not n42893 ; n42893_not
g94885 not n45179 ; n45179_not
g94886 not n12779 ; n12779_not
g94887 not n42299 ; n42299_not
g94888 not n54296 ; n54296_not
g94889 not n42929 ; n42929_not
g94890 not n12599 ; n12599_not
g94891 not n42938 ; n42938_not
g94892 not n42479 ; n42479_not
g94893 not n42947 ; n42947_not
g94894 not n55943 ; n55943_not
g94895 not n38645 ; n38645_not
g94896 not n55952 ; n55952_not
g94897 not n13499 ; n13499_not
g94898 not n55970 ; n55970_not
g94899 not n42596 ; n42596_not
g94900 not n54368 ; n54368_not
g94901 not n42749 ; n42749_not
g94902 not n42758 ; n42758_not
g94903 not n46583 ; n46583_not
g94904 not n42767 ; n42767_not
g94905 not n42776 ; n42776_not
g94906 not n12995 ; n12995_not
g94907 not n42569 ; n42569_not
g94908 not n42785 ; n42785_not
g94909 not n46592 ; n46592_not
g94910 not n12986 ; n12986_not
g94911 not n42794 ; n42794_not
g94912 not n12977 ; n12977_not
g94913 not n12968 ; n12968_not
g94914 not n12959 ; n12959_not
g94915 not n18458 ; n18458_not
g94916 not n42839 ; n42839_not
g94917 not n18449 ; n18449_not
g94918 not n56087 ; n56087_not
g94919 not n46628 ; n46628_not
g94920 not n43199 ; n43199_not
g94921 not n56078 ; n56078_not
g94922 not n18368 ; n18368_not
g94923 not n11969 ; n11969_not
g94924 not n11987 ; n11987_not
g94925 not n45953 ; n45953_not
g94926 not n56159 ; n56159_not
g94927 not n42659 ; n42659_not
g94928 not n56168 ; n56168_not
g94929 not n11897 ; n11897_not
g94930 not n11888 ; n11888_not
g94931 not n11879 ; n11879_not
g94932 not n45962 ; n45962_not
g94933 not n45089 ; n45089_not
g94934 not n54188 ; n54188_not
g94935 not n56177 ; n56177_not
g94936 not n56186 ; n56186_not
g94937 not n11798 ; n11798_not
g94938 not n19088 ; n19088_not
g94939 not n11789 ; n11789_not
g94940 not n45971 ; n45971_not
g94941 not n39095 ; n39095_not
g94942 not n42956 ; n42956_not
g94943 not n42965 ; n42965_not
g94944 not n42974 ; n42974_not
g94945 not n11996 ; n11996_not
g94946 not n54278 ; n54278_not
g94947 not n18395 ; n18395_not
g94948 not n42983 ; n42983_not
g94949 not n42992 ; n42992_not
g94950 not n45944 ; n45944_not
g94951 not n39077 ; n39077_not
g94952 not n42389 ; n42389_not
g94953 not n42398 ; n42398_not
g94954 not n56096 ; n56096_not
g94955 not n11699 ; n11699_not
g94956 not n41858 ; n41858_not
g94957 not n41867 ; n41867_not
g94958 not n18539 ; n18539_not
g94959 not n13994 ; n13994_not
g94960 not n55817 ; n55817_not
g94961 not n45359 ; n45359_not
g94962 not n39293 ; n39293_not
g94963 not n41885 ; n41885_not
g94964 not n46493 ; n46493_not
g94965 not n13985 ; n13985_not
g94966 not n18557 ; n18557_not
g94967 not n41948 ; n41948_not
g94968 not n41957 ; n41957_not
g94969 not n39284 ; n39284_not
g94970 not n18575 ; n18575_not
g94971 not n13976 ; n13976_not
g94972 not n41975 ; n41975_not
g94973 not n13967 ; n13967_not
g94974 not n41993 ; n41993_not
g94975 not n55835 ; n55835_not
g94976 not n39275 ; n39275_not
g94977 not n13886 ; n13886_not
g94978 not n13877 ; n13877_not
g94979 not n55853 ; n55853_not
g94980 not n39266 ; n39266_not
g94981 not n45395 ; n45395_not
g94982 not n41687 ; n41687_not
g94983 not n41696 ; n41696_not
g94984 not n55781 ; n55781_not
g94985 not n18467 ; n18467_not
g94986 not n45386 ; n45386_not
g94987 not n41759 ; n41759_not
g94988 not n46475 ; n46475_not
g94989 not n41768 ; n41768_not
g94990 not n41777 ; n41777_not
g94991 not n18485 ; n18485_not
g94992 not n18494 ; n18494_not
g94993 not n55790 ; n55790_not
g94994 not n45377 ; n45377_not
g94995 not n41786 ; n41786_not
g94996 not n41795 ; n41795_not
g94997 not n13895 ; n13895_not
g94998 not n45368 ; n45368_not
g94999 not n55808 ; n55808_not
g95000 not n54359 ; n54359_not
g95001 not n39158 ; n39158_not
g95002 not n42488 ; n42488_not
g95003 not n45269 ; n45269_not
g95004 not n42578 ; n42578_not
g95005 not n39194 ; n39194_not
g95006 not n55925 ; n55925_not
g95007 not n39185 ; n39185_not
g95008 not n54386 ; n54386_not
g95009 not n46565 ; n46565_not
g95010 not n42668 ; n42668_not
g95011 not n42677 ; n42677_not
g95012 not n42686 ; n42686_not
g95013 not n42695 ; n42695_not
g95014 not n18593 ; n18593_not
g95015 not n55862 ; n55862_not
g95016 not n13859 ; n13859_not
g95017 not n41966 ; n41966_not
g95018 not n39257 ; n39257_not
g95019 not n39248 ; n39248_not
g95020 not n39239 ; n39239_not
g95021 not n18548 ; n18548_not
g95022 not n55880 ; n55880_not
g95023 not n13769 ; n13769_not
g95024 not n45296 ; n45296_not
g95025 not n41876 ; n41876_not
g95026 not n46538 ; n46538_not
g95027 not n55907 ; n55907_not
g95028 not n45287 ; n45287_not
g95029 not n46547 ; n46547_not
g95030 not n45278 ; n45278_not
g95031 not n45854 ; n45854_not
g95032 not n55295 ; n55295_not
g95033 not n45863 ; n45863_not
g95034 not n39725 ; n39725_not
g95035 not n16667 ; n16667_not
g95036 not n16199 ; n16199_not
g95037 not n15677 ; n15677_not
g95038 not n16658 ; n16658_not
g95039 not n16649 ; n16649_not
g95040 not n39941 ; n39941_not
g95041 not n16595 ; n16595_not
g95042 not n45845 ; n45845_not
g95043 not n15686 ; n15686_not
g95044 not n15695 ; n15695_not
g95045 not n16586 ; n16586_not
g95046 not n15767 ; n15767_not
g95047 not n55079 ; n55079_not
g95048 not n16766 ; n16766_not
g95049 not n16757 ; n16757_not
g95050 not n16469 ; n16469_not
g95051 not n45881 ; n45881_not
g95052 not n55277 ; n55277_not
g95053 not n39608 ; n39608_not
g95054 not n16748 ; n16748_not
g95055 not n39815 ; n39815_not
g95056 not n55286 ; n55286_not
g95057 not n55097 ; n55097_not
g95058 not n39923 ; n39923_not
g95059 not n16739 ; n16739_not
g95060 not n16694 ; n16694_not
g95061 not n16397 ; n16397_not
g95062 not n17099 ; n17099_not
g95063 not n16379 ; n16379_not
g95064 not n16685 ; n16685_not
g95065 not n39806 ; n39806_not
g95066 not n39932 ; n39932_not
g95067 not n16676 ; n16676_not
g95068 not n16289 ; n16289_not
g95069 not n15956 ; n15956_not
g95070 not n55349 ; n55349_not
g95071 not n39770 ; n39770_not
g95072 not n45818 ; n45818_not
g95073 not n15947 ; n15947_not
g95074 not n46097 ; n46097_not
g95075 not n15938 ; n15938_not
g95076 not n15929 ; n15929_not
g95077 not n55358 ; n55358_not
g95078 not n17369 ; n17369_not
g95079 not n39761 ; n39761_not
g95080 not n17378 ; n17378_not
g95081 not n17387 ; n17387_not
g95082 not n15893 ; n15893_not
g95083 not n17396 ; n17396_not
g95084 not n55367 ; n55367_not
g95085 not n16577 ; n16577_not
g95086 not n16568 ; n16568_not
g95087 not n16559 ; n16559_not
g95088 not n15992 ; n15992_not
g95089 not n45836 ; n45836_not
g95090 not n17198 ; n17198_not
g95091 not n15983 ; n15983_not
g95092 not n46079 ; n46079_not
g95093 not n39950 ; n39950_not
g95094 not n15776 ; n15776_not
g95095 not n15974 ; n15974_not
g95096 not n55178 ; n55178_not
g95097 not n15785 ; n15785_not
g95098 not n17279 ; n17279_not
g95099 not n17288 ; n17288_not
g95100 not n46088 ; n46088_not
g95101 not n15965 ; n15965_not
g95102 not n17297 ; n17297_not
g95103 not n55169 ; n55169_not
g95104 not n16883 ; n16883_not
g95105 not n16892 ; n16892_not
g95106 not n16298 ; n16298_not
g95107 not n16919 ; n16919_not
g95108 not n16928 ; n16928_not
g95109 not n45926 ; n45926_not
g95110 not n16937 ; n16937_not
g95111 not n45980 ; n45980_not
g95112 not n39644 ; n39644_not
g95113 not n45890 ; n45890_not
g95114 not n16946 ; n16946_not
g95115 not n16955 ; n16955_not
g95116 not n16829 ; n16829_not
g95117 not n16793 ; n16793_not
g95118 not n16838 ; n16838_not
g95119 not n16784 ; n16784_not
g95120 not n55187 ; n55187_not
g95121 not n16775 ; n16775_not
g95122 not n16847 ; n16847_not
g95123 not n16856 ; n16856_not
g95124 not n16865 ; n16865_not
g95125 not n16388 ; n16388_not
g95126 not n39860 ; n39860_not
g95127 not n16874 ; n16874_not
g95128 not n39842 ; n39842_not
g95129 not n39617 ; n39617_not
g95130 not n55259 ; n55259_not
g95131 not n39653 ; n39653_not
g95132 not n15857 ; n15857_not
g95133 not n55268 ; n55268_not
g95134 not n39833 ; n39833_not
g95135 not n39662 ; n39662_not
g95136 not n39914 ; n39914_not
g95137 not n16487 ; n16487_not
g95138 not n39824 ; n39824_not
g95139 not n16478 ; n16478_not
g95140 not n16964 ; n16964_not
g95141 not n16973 ; n16973_not
g95142 not n45908 ; n45908_not
g95143 not n39905 ; n39905_not
g95144 not n39851 ; n39851_not
g95145 not n16991 ; n16991_not
g95146 not n17594 ; n17594_not
g95147 not n45647 ; n45647_not
g95148 not n55538 ; n55538_not
g95149 not n14894 ; n14894_not
g95150 not n39626 ; n39626_not
g95151 not n45638 ; n45638_not
g95152 not n17657 ; n17657_not
g95153 not n45764 ; n45764_not
g95154 not n16982 ; n16982_not
g95155 not n17567 ; n17567_not
g95156 not n39671 ; n39671_not
g95157 not n17576 ; n17576_not
g95158 not n46187 ; n46187_not
g95159 not n45665 ; n45665_not
g95160 not n17585 ; n17585_not
g95161 not n45656 ; n45656_not
g95162 not n55529 ; n55529_not
g95163 not n46196 ; n46196_not
g95164 not n14957 ; n14957_not
g95165 not n55574 ; n55574_not
g95166 not n45746 ; n45746_not
g95167 not n14948 ; n14948_not
g95168 not n45593 ; n45593_not
g95169 not n14939 ; n14939_not
g95170 not n17792 ; n17792_not
g95171 not n45584 ; n45584_not
g95172 not n55583 ; n55583_not
g95173 not n17837 ; n17837_not
g95174 not n39563 ; n39563_not
g95175 not n46259 ; n46259_not
g95176 not n45629 ; n45629_not
g95177 not n55547 ; n55547_not
g95178 not n45755 ; n45755_not
g95179 not n14966 ; n14966_not
g95180 not n55556 ; n55556_not
g95181 not n39752 ; n39752_not
g95182 not n39743 ; n39743_not
g95183 not n17747 ; n17747_not
g95184 not n39734 ; n39734_not
g95185 not n55565 ; n55565_not
g95186 not n39581 ; n39581_not
g95187 not n39572 ; n39572_not
g95188 not n17459 ; n17459_not
g95189 not n17468 ; n17468_not
g95190 not n15749 ; n15749_not
g95191 not n54962 ; n54962_not
g95192 not n17477 ; n17477_not
g95193 not n45809 ; n45809_not
g95194 not n17486 ; n17486_not
g95195 not n15659 ; n15659_not
g95196 not n15884 ; n15884_not
g95197 not n15875 ; n15875_not
g95198 not n55376 ; n55376_not
g95199 not n45791 ; n45791_not
g95200 not n39707 ; n39707_not
g95201 not n15866 ; n15866_not
g95202 not n15848 ; n15848_not
g95203 not n15839 ; n15839_not
g95204 not n55385 ; n55385_not
g95205 not n15794 ; n15794_not
g95206 not n55394 ; n55394_not
g95207 not n45773 ; n45773_not
g95208 not n55448 ; n55448_not
g95209 not n15488 ; n15488_not
g95210 not n15479 ; n15479_not
g95211 not n55457 ; n55457_not
g95212 not n55466 ; n55466_not
g95213 not n15398 ; n15398_not
g95214 not n55475 ; n55475_not
g95215 not n15389 ; n15389_not
g95216 not n46169 ; n46169_not
g95217 not n55484 ; n55484_not
g95218 not n54089 ; n54089_not
g95219 not n17549 ; n17549_not
g95220 not n55493 ; n55493_not
g95221 not n45683 ; n45683_not
g95222 not n55088 ; n55088_not
g95223 not n15299 ; n15299_not
g95224 not n17558 ; n17558_not
g95225 not n46178 ; n46178_not
g95226 not n15596 ; n15596_not
g95227 not n17495 ; n17495_not
g95228 not n39716 ; n39716_not
g95229 not n14993 ; n14993_not
g95230 not n15587 ; n15587_not
g95231 not n15578 ; n15578_not
g95232 not n45728 ; n45728_not
g95233 not n15569 ; n15569_not
g95234 not n54926 ; n54926_not
g95235 not n55439 ; n55439_not
g95236 not n15497 ; n15497_not
g95237 not n46466 ; n46466_not
g95238 not n43847 ; n43847_not
g95239 not n56447 ; n56447_not
g95240 not n38753 ; n38753_not
g95241 not n56438 ; n56438_not
g95242 not n43838 ; n43838_not
g95243 not n56816 ; n56816_not
g95244 not n56429 ; n56429_not
g95245 not n56825 ; n56825_not
g95246 not n43829 ; n43829_not
g95247 not n53792 ; n53792_not
g95248 not n56393 ; n56393_not
g95249 not n56843 ; n56843_not
g95250 not n44099 ; n44099_not
g95251 not n56384 ; n56384_not
g95252 not n38744 ; n38744_not
g95253 not n43991 ; n43991_not
g95254 not n53819 ; n53819_not
g95255 not n56555 ; n56555_not
g95256 not n56753 ; n56753_not
g95257 not n38771 ; n38771_not
g95258 not n56546 ; n56546_not
g95259 not n19772 ; n19772_not
g95260 not n56537 ; n56537_not
g95261 not n56528 ; n56528_not
g95262 not n56519 ; n56519_not
g95263 not n56771 ; n56771_not
g95264 not n56780 ; n56780_not
g95265 not n56492 ; n56492_not
g95266 not n38762 ; n38762_not
g95267 not n56483 ; n56483_not
g95268 not n56474 ; n56474_not
g95269 not n56465 ; n56465_not
g95270 not n56456 ; n56456_not
g95271 not n38717 ; n38717_not
g95272 not n56906 ; n56906_not
g95273 not n56267 ; n56267_not
g95274 not n56915 ; n56915_not
g95275 not n38708 ; n38708_not
g95276 not n56258 ; n56258_not
g95277 not n38609 ; n38609_not
g95278 not n53765 ; n53765_not
g95279 not n38618 ; n38618_not
g95280 not n56249 ; n56249_not
g95281 not n53756 ; n53756_not
g95282 not n44189 ; n44189_not
g95283 not n38690 ; n38690_not
g95284 not n56375 ; n56375_not
g95285 not n53783 ; n53783_not
g95286 not n56366 ; n56366_not
g95287 not n56357 ; n56357_not
g95288 not n43793 ; n43793_not
g95289 not n38735 ; n38735_not
g95290 not n56861 ; n56861_not
g95291 not n56348 ; n56348_not
g95292 not n56870 ; n56870_not
g95293 not n56339 ; n56339_not
g95294 not n53774 ; n53774_not
g95295 not n38726 ; n38726_not
g95296 not n19817 ; n19817_not
g95297 not n43784 ; n43784_not
g95298 not n56294 ; n56294_not
g95299 not n56285 ; n56285_not
g95300 not n56276 ; n56276_not
g95301 not n56582 ; n56582_not
g95302 not n38834 ; n38834_not
g95303 not n53936 ; n53936_not
g95304 not n56591 ; n56591_not
g95305 not n43874 ; n43874_not
g95306 not n38825 ; n38825_not
g95307 not n53927 ; n53927_not
g95308 not n56609 ; n56609_not
g95309 not n43883 ; n43883_not
g95310 not n55826 ; n55826_not
g95311 not n38816 ; n38816_not
g95312 not n56618 ; n56618_not
g95313 not n53918 ; n53918_not
g95314 not n56627 ; n56627_not
g95315 not n56636 ; n56636_not
g95316 not n38807 ; n38807_not
g95317 not n38555 ; n38555_not
g95318 not n53909 ; n53909_not
g95319 not n56645 ; n56645_not
g95320 not n43919 ; n43919_not
g95321 not n19187 ; n19187_not
g95322 not n55871 ; n55871_not
g95323 not n38870 ; n38870_not
g95324 not n38519 ; n38519_not
g95325 not n53963 ; n53963_not
g95326 not n53954 ; n53954_not
g95327 not n38861 ; n38861_not
g95328 not n38528 ; n38528_not
g95329 not n19178 ; n19178_not
g95330 not n38852 ; n38852_not
g95331 not n56564 ; n56564_not
g95332 not n53945 ; n53945_not
g95333 not n38843 ; n38843_not
g95334 not n56573 ; n56573_not
g95335 not n43856 ; n43856_not
g95336 not n56708 ; n56708_not
g95337 not n53855 ; n53855_not
g95338 not n53369 ; n53369_not
g95339 not n43973 ; n43973_not
g95340 not n44387 ; n44387_not
g95341 not n53846 ; n53846_not
g95342 not n56726 ; n56726_not
g95343 not n53837 ; n53837_not
g95344 not n43982 ; n43982_not
g95345 not n56735 ; n56735_not
g95346 not n38780 ; n38780_not
g95347 not n38573 ; n38573_not
g95348 not n53828 ; n53828_not
g95349 not n43928 ; n43928_not
g95350 not n56654 ; n56654_not
g95351 not n53891 ; n53891_not
g95352 not n56663 ; n56663_not
g95353 not n44369 ; n44369_not
g95354 not n43937 ; n43937_not
g95355 not n53882 ; n53882_not
g95356 not n19097 ; n19097_not
g95357 not n43946 ; n43946_not
g95358 not n56690 ; n56690_not
g95359 not n53873 ; n53873_not
g95360 not n43892 ; n43892_not
g95361 not n43955 ; n43955_not
g95362 not n38564 ; n38564_not
g95363 not n53864 ; n53864_not
g95364 not n44378 ; n44378_not
g95365 not n43964 ; n43964_not
g95366 not n57275 ; n57275_not
g95367 not n38474 ; n38474_not
g95368 not n19349 ; n19349_not
g95369 not n44567 ; n44567_not
g95370 not n57284 ; n57284_not
g95371 not n53639 ; n53639_not
g95372 not n44558 ; n44558_not
g95373 not n44585 ; n44585_not
g95374 not n19358 ; n19358_not
g95375 not n19367 ; n19367_not
g95376 not n38447 ; n38447_not
g95377 not n19376 ; n19376_not
g95378 not n44594 ; n44594_not
g95379 not n19385 ; n19385_not
g95380 not n19394 ; n19394_not
g95381 not n57257 ; n57257_not
g95382 not n53666 ; n53666_not
g95383 not n19970 ; n19970_not
g95384 not n44468 ; n44468_not
g95385 not n57266 ; n57266_not
g95386 not n53657 ; n53657_not
g95387 not n44549 ; n44549_not
g95388 not n38492 ; n38492_not
g95389 not n44477 ; n44477_not
g95390 not n53648 ; n53648_not
g95391 not n57428 ; n57428_not
g95392 not n53585 ; n53585_not
g95393 not n38384 ; n38384_not
g95394 not n19934 ; n19934_not
g95395 not n56951 ; n56951_not
g95396 not n19475 ; n19475_not
g95397 not n57446 ; n57446_not
g95398 not n19484 ; n19484_not
g95399 not n56960 ; n56960_not
g95400 not n38375 ; n38375_not
g95401 not n53576 ; n53576_not
g95402 not n19925 ; n19925_not
g95403 not n19493 ; n19493_not
g95404 not n57473 ; n57473_not
g95405 not n38366 ; n38366_not
g95406 not n57482 ; n57482_not
g95407 not n38357 ; n38357_not
g95408 not n38348 ; n38348_not
g95409 not n53567 ; n53567_not
g95410 not n38339 ; n38339_not
g95411 not n19529 ; n19529_not
g95412 not n57491 ; n57491_not
g95413 not n19538 ; n19538_not
g95414 not n53558 ; n53558_not
g95415 not n19547 ; n19547_not
g95416 not n38294 ; n38294_not
g95417 not n38438 ; n38438_not
g95418 not n38429 ; n38429_not
g95419 not n57329 ; n57329_not
g95420 not n57338 ; n57338_not
g95421 not n57347 ; n57347_not
g95422 not n19439 ; n19439_not
g95423 not n57356 ; n57356_not
g95424 not n19448 ; n19448_not
g95425 not n57374 ; n57374_not
g95426 not n53594 ; n53594_not
g95427 not n56924 ; n56924_not
g95428 not n38393 ; n38393_not
g95429 not n19457 ; n19457_not
g95430 not n19943 ; n19943_not
g95431 not n57419 ; n57419_not
g95432 not n19466 ; n19466_not
g95433 not n44279 ; n44279_not
g95434 not n44288 ; n44288_not
g95435 not n53729 ; n53729_not
g95436 not n44297 ; n44297_not
g95437 not n38672 ; n38672_not
g95438 not n43694 ; n43694_not
g95439 not n38663 ; n38663_not
g95440 not n43685 ; n43685_not
g95441 not n43757 ; n43757_not
g95442 not n44198 ; n44198_not
g95443 not n56933 ; n56933_not
g95444 not n53747 ; n53747_not
g95445 not n43748 ; n43748_not
g95446 not n19862 ; n19862_not
g95447 not n56195 ; n56195_not
g95448 not n43739 ; n43739_not
g95449 not n38681 ; n38681_not
g95450 not n53738 ; n53738_not
g95451 not n38582 ; n38582_not
g95452 not n44459 ; n44459_not
g95453 not n53459 ; n53459_not
g95454 not n57158 ; n57158_not
g95455 not n44486 ; n44486_not
g95456 not n53684 ; n53684_not
g95457 not n19952 ; n19952_not
g95458 not n53675 ; n53675_not
g95459 not n57185 ; n57185_not
g95460 not n57194 ; n57194_not
g95461 not n38537 ; n38537_not
g95462 not n56834 ; n56834_not
g95463 not n19907 ; n19907_not
g95464 not n57059 ; n57059_not
g95465 not n57068 ; n57068_not
g95466 not n38654 ; n38654_not
g95467 not n57086 ; n57086_not
g95468 not n38627 ; n38627_not
g95469 not n56744 ; n56744_not
g95470 not n44396 ; n44396_not
g95471 not n53693 ; n53693_not
g95472 not n53981 ; n53981_not
g95473 not n38942 ; n38942_not
g95474 not n10997 ; n10997_not
g95475 not n38915 ; n38915_not
g95476 not n19268 ; n19268_not
g95477 not n10979 ; n10979_not
g95478 not n19196 ; n19196_not
g95479 not n43676 ; n43676_not
g95480 not n55961 ; n55961_not
g95481 not n19295 ; n19295_not
g95482 not n10988 ; n10988_not
g95483 not n38483 ; n38483_not
g95484 not n53990 ; n53990_not
g95485 not n38960 ; n38960_not
g95486 not n10889 ; n10889_not
g95487 not n53279 ; n53279_not
g95488 not n43766 ; n43766_not
g95489 not n10799 ; n10799_not
g95490 not n38951 ; n38951_not
g95491 not n38906 ; n38906_not
g95492 not n19277 ; n19277_not
g95493 not n54098 ; n54098_not
g95494 not n55916 ; n55916_not
g95495 not n46556 ; n46556_not
g95496 not n10898 ; n10898_not
g95497 not n19286 ; n19286_not
g95498 not n38924 ; n38924_not
g95499 not n53972 ; n53972_not
g95500 not n38933 ; n38933_not
g95501 not n39582 ; n39582_not
g95502 not n51867 ; n51867_not
g95503 not n32994 ; n32994_not
g95504 not n35748 ; n35748_not
g95505 not n55359 ; n55359_not
g95506 not n48816 ; n48816_not
g95507 not n44478 ; n44478_not
g95508 not n27783 ; n27783_not
g95509 not n29619 ; n29619_not
g95510 not n49419 ; n49419_not
g95511 not n15894 ; n15894_not
g95512 not n56781 ; n56781_not
g95513 not n42966 ; n42966_not
g95514 not n27774 ; n27774_not
g95515 not n35676 ; n35676_not
g95516 not n49068 ; n49068_not
g95517 not n29637 ; n29637_not
g95518 not n51858 ; n51858_not
g95519 not n31689 ; n31689_not
g95520 not n29871 ; n29871_not
g95521 not n28089 ; n28089_not
g95522 not n56754 ; n56754_not
g95523 not n35757 ; n35757_not
g95524 not n31698 ; n31698_not
g95525 not n44199 ; n44199_not
g95526 not n42939 ; n42939_not
g95527 not n49095 ; n49095_not
g95528 not n29880 ; n29880_not
g95529 not n15867 ; n15867_not
g95530 not n27828 ; n27828_not
g95531 not n55377 ; n55377_not
g95532 not n44784 ; n44784_not
g95533 not n29592 ; n29592_not
g95534 not n49086 ; n49086_not
g95535 not n11988 ; n11988_not
g95536 not n42957 ; n42957_not
g95537 not n55368 ; n55368_not
g95538 not n55089 ; n55089_not
g95539 not n49077 ; n49077_not
g95540 not n15885 ; n15885_not
g95541 not n45675 ; n45675_not
g95542 not n55485 ; n55485_not
g95543 not n44469 ; n44469_not
g95544 not n43596 ; n43596_not
g95545 not n15876 ; n15876_not
g95546 not n34749 ; n34749_not
g95547 not n39573 ; n39573_not
g95548 not n42948 ; n42948_not
g95549 not n34839 ; n34839_not
g95550 not n51885 ; n51885_not
g95551 not n31797 ; n31797_not
g95552 not n43992 ; n43992_not
g95553 not n27747 ; n27747_not
g95554 not n48672 ; n48672_not
g95555 not n43587 ; n43587_not
g95556 not n15966 ; n15966_not
g95557 not n29655 ; n29655_not
g95558 not n26892 ; n26892_not
g95559 not n31995 ; n31995_not
g95560 not n35658 ; n35658_not
g95561 not n45828 ; n45828_not
g95562 not n57195 ; n57195_not
g95563 not n44766 ; n44766_not
g95564 not n27396 ; n27396_not
g95565 not n14589 ; n14589_not
g95566 not n43983 ; n43983_not
g95567 not n27738 ; n27738_not
g95568 not n12978 ; n12978_not
g95569 not n11997 ; n11997_not
g95570 not n26883 ; n26883_not
g95571 not n48681 ; n48681_not
g95572 not n26937 ; n26937_not
g95573 not n15975 ; n15975_not
g95574 not n27729 ; n27729_not
g95575 not n56826 ; n56826_not
g95576 not n34767 ; n34767_not
g95577 not n32976 ; n32976_not
g95578 not n56790 ; n56790_not
g95579 not n44775 ; n44775_not
g95580 not n12969 ; n12969_not
g95581 not n48663 ; n48663_not
g95582 not n33588 ; n33588_not
g95583 not n35667 ; n35667_not
g95584 not n31977 ; n31977_not
g95585 not n49059 ; n49059_not
g95586 not n45684 ; n45684_not
g95587 not n55494 ; n55494_not
g95588 not n56943 ; n56943_not
g95589 not n15939 ; n15939_not
g95590 not n29529 ; n29529_not
g95591 not n33597 ; n33597_not
g95592 not n57186 ; n57186_not
g95593 not n27378 ; n27378_not
g95594 not n48573 ; n48573_not
g95595 not n15786 ; n15786_not
g95596 not n27756 ; n27756_not
g95597 not n31986 ; n31986_not
g95598 not n15957 ; n15957_not
g95599 not n34596 ; n34596_not
g95600 not n43749 ; n43749_not
g95601 not n27288 ; n27288_not
g95602 not n27765 ; n27765_not
g95603 not n57177 ; n57177_not
g95604 not n44496 ; n44496_not
g95605 not n15795 ; n15795_not
g95606 not n42975 ; n42975_not
g95607 not n15948 ; n15948_not
g95608 not n51777 ; n51777_not
g95609 not n34686 ; n34686_not
g95610 not n49158 ; n49158_not
g95611 not n56682 ; n56682_not
g95612 not n55962 ; n55962_not
g95613 not n45738 ; n45738_not
g95614 not n42876 ; n42876_not
g95615 not n56961 ; n56961_not
g95616 not n56691 ; n56691_not
g95617 not n55458 ; n55458_not
g95618 not n31779 ; n31779_not
g95619 not n49194 ; n49194_not
g95620 not n45189 ; n45189_not
g95621 not n50886 ; n50886_not
g95622 not n48618 ; n48618_not
g95623 not n55971 ; n55971_not
g95624 not n55467 ; n55467_not
g95625 not n29493 ; n29493_not
g95626 not n43677 ; n43677_not
g95627 not n15669 ; n15669_not
g95628 not n27918 ; n27918_not
g95629 not n33399 ; n33399_not
g95630 not n12699 ; n12699_not
g95631 not n49842 ; n49842_not
g95632 not n49149 ; n49149_not
g95633 not n56709 ; n56709_not
g95634 not n14985 ; n14985_not
g95635 not n34695 ; n34695_not
g95636 not n27936 ; n27936_not
g95637 not n43659 ; n43659_not
g95638 not n42849 ; n42849_not
g95639 not n33489 ; n33489_not
g95640 not n55449 ; n55449_not
g95641 not n42858 ; n42858_not
g95642 not n49185 ; n49185_not
g95643 not n39528 ; n39528_not
g95644 not n44289 ; n44289_not
g95645 not n27963 ; n27963_not
g95646 not n56970 ; n56970_not
g95647 not n51399 ; n51399_not
g95648 not n49176 ; n49176_not
g95649 not n39537 ; n39537_not
g95650 not n34677 ; n34677_not
g95651 not n34668 ; n34668_not
g95652 not n27945 ; n27945_not
g95653 not n44298 ; n44298_not
g95654 not n42867 ; n42867_not
g95655 not n14994 ; n14994_not
g95656 not n27990 ; n27990_not
g95657 not n49167 ; n49167_not
g95658 not n12879 ; n12879_not
g95659 not n51768 ; n51768_not
g95660 not n49833 ; n49833_not
g95661 not n27981 ; n27981_not
g95662 not n12888 ; n12888_not
g95663 not n50589 ; n50589_not
g95664 not n29907 ; n29907_not
g95665 not n33498 ; n33498_not
g95666 not n34479 ; n34479_not
g95667 not n44379 ; n44379_not
g95668 not n48582 ; n48582_not
g95669 not n44388 ; n44388_not
g95670 not n32958 ; n32958_not
g95671 not n43668 ; n43668_not
g95672 not n27873 ; n27873_not
g95673 not n48636 ; n48636_not
g95674 not n56736 ; n56736_not
g95675 not n55395 ; n55395_not
g95676 not n15777 ; n15777_not
g95677 not n12897 ; n12897_not
g95678 not n34587 ; n34587_not
g95679 not n49860 ; n49860_not
g95680 not n42489 ; n42489_not
g95681 not n33579 ; n33579_not
g95682 not n29745 ; n29745_not
g95683 not n56745 ; n56745_not
g95684 not n55386 ; n55386_not
g95685 not n55098 ; n55098_not
g95686 not n27846 ; n27846_not
g95687 not n45783 ; n45783_not
g95688 not n34578 ; n34578_not
g95689 not n45693 ; n45693_not
g95690 not n32967 ; n32967_not
g95691 not n27855 ; n27855_not
g95692 not n42885 ; n42885_not
g95693 not n34794 ; n34794_not
g95694 not n12798 ; n12798_not
g95695 not n49824 ; n49824_not
g95696 not n48591 ; n48591_not
g95697 not n12789 ; n12789_not
g95698 not n34659 ; n34659_not
g95699 not n15687 ; n15687_not
g95700 not n45756 ; n45756_not
g95701 not n51795 ; n51795_not
g95702 not n57078 ; n57078_not
g95703 not n55953 ; n55953_not
g95704 not n39564 ; n39564_not
g95705 not n50598 ; n50598_not
g95706 not n32949 ; n32949_not
g95707 not n34785 ; n34785_not
g95708 not n42894 ; n42894_not
g95709 not n15759 ; n15759_not
g95710 not n44793 ; n44793_not
g95711 not n48627 ; n48627_not
g95712 not n29484 ; n29484_not
g95713 not n45765 ; n45765_not
g95714 not n27891 ; n27891_not
g95715 not n34569 ; n34569_not
g95716 not n29736 ; n29736_not
g95717 not n15696 ; n15696_not
g95718 not n49851 ; n49851_not
g95719 not n55476 ; n55476_not
g95720 not n10989 ; n10989_not
g95721 not n43497 ; n43497_not
g95722 not n26388 ; n26388_not
g95723 not n48906 ; n48906_not
g95724 not n26397 ; n26397_not
g95725 not n32769 ; n32769_not
g95726 not n16578 ; n16578_not
g95727 not n57366 ; n57366_not
g95728 not n11979 ; n11979_not
g95729 not n10998 ; n10998_not
g95730 not n29781 ; n29781_not
g95731 not n49932 ; n49932_not
g95732 not n32778 ; n32778_not
g95733 not n27279 ; n27279_not
g95734 not n57348 ; n57348_not
g95735 not n49338 ; n49338_not
g95736 not n50994 ; n50994_not
g95737 not n29772 ; n29772_not
g95738 not n29790 ; n29790_not
g95739 not n32679 ; n32679_not
g95740 not n44649 ; n44649_not
g95741 not n45918 ; n45918_not
g95742 not n57393 ; n57393_not
g95743 not n56925 ; n56925_not
g95744 not n42669 ; n42669_not
g95745 not n27189 ; n27189_not
g95746 not n39627 ; n39627_not
g95747 not n16596 ; n16596_not
g95748 not n50499 ; n50499_not
g95749 not n16587 ; n16587_not
g95750 not n56916 ; n56916_not
g95751 not n48753 ; n48753_not
g95752 not n39618 ; n39618_not
g95753 not n26379 ; n26379_not
g95754 not n56880 ; n56880_not
g95755 not n48924 ; n48924_not
g95756 not n32796 ; n32796_not
g95757 not n56871 ; n56871_not
g95758 not n44595 ; n44595_not
g95759 not n44487 ; n44487_not
g95760 not n27387 ; n27387_not
g95761 not n26559 ; n26559_not
g95762 not n29754 ; n29754_not
g95763 not n26568 ; n26568_not
g95764 not n48933 ; n48933_not
g95765 not n32499 ; n32499_not
g95766 not n26577 ; n26577_not
g95767 not n49923 ; n49923_not
g95768 not n11898 ; n11898_not
g95769 not n57339 ; n57339_not
g95770 not n16479 ; n16479_not
g95771 not n16569 ; n16569_not
g95772 not n32787 ; n32787_not
g95773 not n27297 ; n27297_not
g95774 not n48915 ; n48915_not
g95775 not n26469 ; n26469_not
g95776 not n26478 ; n26478_not
g95777 not n36099 ; n36099_not
g95778 not n29844 ; n29844_not
g95779 not n26487 ; n26487_not
g95780 not n26496 ; n26496_not
g95781 not n16488 ; n16488_not
g95782 not n27369 ; n27369_not
g95783 not n29817 ; n29817_not
g95784 not n43389 ; n43389_not
g95785 not n32589 ; n32589_not
g95786 not n16758 ; n16758_not
g95787 not n29826 ; n29826_not
g95788 not n48852 ; n48852_not
g95789 not n50958 ; n50958_not
g95790 not n57474 ; n57474_not
g95791 not n16749 ; n16749_not
g95792 not n45936 ; n45936_not
g95793 not n48861 ; n48861_not
g95794 not n57465 ; n57465_not
g95795 not n49950 ; n49950_not
g95796 not n57492 ; n57492_not
g95797 not n51786 ; n51786_not
g95798 not n16794 ; n16794_not
g95799 not n55197 ; n55197_not
g95800 not n43398 ; n43398_not
g95801 not n48834 ; n48834_not
g95802 not n26982 ; n26982_not
g95803 not n16785 ; n16785_not
g95804 not n50949 ; n50949_not
g95805 not n26991 ; n26991_not
g95806 not n34299 ; n34299_not
g95807 not n44694 ; n44694_not
g95808 not n16776 ; n16776_not
g95809 not n36189 ; n36189_not
g95810 not n48843 ; n48843_not
g95811 not n57483 ; n57483_not
g95812 not n16767 ; n16767_not
g95813 not n44667 ; n44667_not
g95814 not n43488 ; n43488_not
g95815 not n45927 ; n45927_not
g95816 not n48762 ; n48762_not
g95817 not n43299 ; n43299_not
g95818 not n50976 ; n50976_not
g95819 not n49941 ; n49941_not
g95820 not n16668 ; n16668_not
g95821 not n54387 ; n54387_not
g95822 not n44658 ; n44658_not
g95823 not n56934 ; n56934_not
g95824 not n29835 ; n29835_not
g95825 not n16659 ; n16659_not
g95826 not n45099 ; n45099_not
g95827 not n32688 ; n32688_not
g95828 not n44685 ; n44685_not
g95829 not n16389 ; n16389_not
g95830 not n16398 ; n16398_not
g95831 not n10899 ; n10899_not
g95832 not n16695 ; n16695_not
g95833 not n48870 ; n48870_not
g95834 not n16686 ; n16686_not
g95835 not n43479 ; n43479_not
g95836 not n27099 ; n27099_not
g95837 not n44676 ; n44676_not
g95838 not n48771 ; n48771_not
g95839 not n16677 ; n16677_not
g95840 not n57438 ; n57438_not
g95841 not n27648 ; n27648_not
g95842 not n56097 ; n56097_not
g95843 not n27657 ; n27657_not
g95844 not n45855 ; n45855_not
g95845 not n43938 ; n43938_not
g95846 not n29682 ; n29682_not
g95847 not n43947 ; n43947_not
g95848 not n43569 ; n43569_not
g95849 not n43956 ; n43956_not
g95850 not n57267 ; n57267_not
g95851 not n27666 ; n27666_not
g95852 not n45846 ; n45846_not
g95853 not n26757 ; n26757_not
g95854 not n26766 ; n26766_not
g95855 not n44559 ; n44559_not
g95856 not n43929 ; n43929_not
g95857 not n32598 ; n32598_not
g95858 not n42993 ; n42993_not
g95859 not n29691 ; n29691_not
g95860 not n26775 ; n26775_not
g95861 not n49329 ; n49329_not
g95862 not n55296 ; n55296_not
g95863 not n26784 ; n26784_not
g95864 not n32895 ; n32895_not
g95865 not n27639 ; n27639_not
g95866 not n44748 ; n44748_not
g95867 not n49374 ; n49374_not
g95868 not n26793 ; n26793_not
g95869 not n15993 ; n15993_not
g95870 not n42984 ; n42984_not
g95871 not n29862 ; n29862_not
g95872 not n43578 ; n43578_not
g95873 not n43965 ; n43965_not
g95874 not n26856 ; n26856_not
g95875 not n26946 ; n26946_not
g95876 not n26865 ; n26865_not
g95877 not n56844 ; n56844_not
g95878 not n55179 ; n55179_not
g95879 not n26874 ; n26874_not
g95880 not n57249 ; n57249_not
g95881 not n29664 ; n29664_not
g95882 not n15984 ; n15984_not
g95883 not n43974 ; n43974_not
g95884 not n56835 ; n56835_not
g95885 not n27675 ; n27675_not
g95886 not n26829 ; n26829_not
g95887 not n27684 ; n27684_not
g95888 not n55188 ; n55188_not
g95889 not n34758 ; n34758_not
g95890 not n29628 ; n29628_not
g95891 not n49383 ; n49383_not
g95892 not n26838 ; n26838_not
g95893 not n44757 ; n44757_not
g95894 not n56088 ; n56088_not
g95895 not n57258 ; n57258_not
g95896 not n27693 ; n27693_not
g95897 not n26847 ; n26847_not
g95898 not n26955 ; n26955_not
g95899 not n29673 ; n29673_not
g95900 not n16497 ; n16497_not
g95901 not n27477 ; n27477_not
g95902 not n27486 ; n27486_not
g95903 not n32859 ; n32859_not
g95904 not n27495 ; n27495_not
g95905 not n26649 ; n26649_not
g95906 not n26658 ; n26658_not
g95907 not n48951 ; n48951_not
g95908 not n26667 ; n26667_not
g95909 not n44739 ; n44739_not
g95910 not n49914 ; n49914_not
g95911 not n26676 ; n26676_not
g95912 not n48726 ; n48726_not
g95913 not n26586 ; n26586_not
g95914 not n44577 ; n44577_not
g95915 not n26595 ; n26595_not
g95916 not n45891 ; n45891_not
g95917 not n11889 ; n11889_not
g95918 not n27459 ; n27459_not
g95919 not n55269 ; n55269_not
g95920 not n49365 ; n49365_not
g95921 not n11799 ; n11799_not
g95922 not n57294 ; n57294_not
g95923 not n44586 ; n44586_not
g95924 not n27468 ; n27468_not
g95925 not n48942 ; n48942_not
g95926 not n27576 ; n27576_not
g95927 not n44568 ; n44568_not
g95928 not n51876 ; n51876_not
g95929 not n27585 ; n27585_not
g95930 not n29709 ; n29709_not
g95931 not n26739 ; n26739_not
g95932 not n45873 ; n45873_not
g95933 not n27594 ; n27594_not
g95934 not n26748 ; n26748_not
g95935 not n49905 ; n49905_not
g95936 not n32886 ; n32886_not
g95937 not n16299 ; n16299_not
g95938 not n48708 ; n48708_not
g95939 not n26685 ; n26685_not
g95940 not n32868 ; n32868_not
g95941 not n26694 ; n26694_not
g95942 not n34389 ; n34389_not
g95943 not n27549 ; n27549_not
g95944 not n29853 ; n29853_not
g95945 not n48960 ; n48960_not
g95946 not n39609 ; n39609_not
g95947 not n55278 ; n55278_not
g95948 not n27558 ; n27558_not
g95949 not n32877 ; n32877_not
g95950 not n48717 ; n48717_not
g95951 not n29718 ; n29718_not
g95952 not n57276 ; n57276_not
g95953 not n27567 ; n27567_not
g95954 not n55287 ; n55287_not
g95955 not n33939 ; n33939_not
g95956 not n44928 ; n44928_not
g95957 not n45459 ; n45459_not
g95958 not n27954 ; n27954_not
g95959 not n33858 ; n33858_not
g95960 not n49527 ; n49527_not
g95961 not n50688 ; n50688_not
g95962 not n14598 ; n14598_not
g95963 not n33948 ; n33948_not
g95964 not n43893 ; n43893_not
g95965 not n13797 ; n13797_not
g95966 not n28665 ; n28665_not
g95967 not n51498 ; n51498_not
g95968 not n55872 ; n55872_not
g95969 not n49509 ; n49509_not
g95970 not n49815 ; n49815_not
g95971 not n33795 ; n33795_not
g95972 not n55692 ; n55692_not
g95973 not n29196 ; n29196_not
g95974 not n33849 ; n33849_not
g95975 not n28647 ; n28647_not
g95976 not n29187 ; n29187_not
g95977 not n34947 ; n34947_not
g95978 not n49716 ; n49716_not
g95979 not n56673 ; n56673_not
g95980 not n49545 ; n49545_not
g95981 not n13599 ; n13599_not
g95982 not n55719 ; n55719_not
g95983 not n41958 ; n41958_not
g95984 not n50796 ; n50796_not
g95985 not n34893 ; n34893_not
g95986 not n13968 ; n13968_not
g95987 not n49554 ; n49554_not
g95988 not n29178 ; n29178_not
g95989 not n13977 ; n13977_not
g95990 not n50679 ; n50679_not
g95991 not n13986 ; n13986_not
g95992 not n13995 ; n13995_not
g95993 not n33876 ; n33876_not
g95994 not n55791 ; n55791_not
g95995 not n51489 ; n51489_not
g95996 not n33867 ; n33867_not
g95997 not n50697 ; n50697_not
g95998 not n44937 ; n44937_not
g95999 not n34848 ; n34848_not
g96000 not n33957 ; n33957_not
g96001 not n28683 ; n28683_not
g96002 not n41877 ; n41877_not
g96003 not n49464 ; n49464_not
g96004 not n45495 ; n45495_not
g96005 not n28539 ; n28539_not
g96006 not n56718 ; n56718_not
g96007 not n33777 ; n33777_not
g96008 not n13698 ; n13698_not
g96009 not n50769 ; n50769_not
g96010 not n55665 ; n55665_not
g96011 not n49473 ; n49473_not
g96012 not n45297 ; n45297_not
g96013 not n41886 ; n41886_not
g96014 not n28557 ; n28557_not
g96015 not n45486 ; n45486_not
g96016 not n30996 ; n30996_not
g96017 not n55647 ; n55647_not
g96018 not n41868 ; n41868_not
g96019 not n29961 ; n29961_not
g96020 not n50778 ; n50778_not
g96021 not n43776 ; n43776_not
g96022 not n49761 ; n49761_not
g96023 not n55656 ; n55656_not
g96024 not n49455 ; n49455_not
g96025 not n49770 ; n49770_not
g96026 not n50859 ; n50859_not
g96027 not n34938 ; n34938_not
g96028 not n33759 ; n33759_not
g96029 not n40797 ; n40797_not
g96030 not n49734 ; n49734_not
g96031 not n29169 ; n29169_not
g96032 not n28593 ; n28593_not
g96033 not n45477 ; n45477_not
g96034 not n33894 ; n33894_not
g96035 not n33786 ; n33786_not
g96036 not n44919 ; n44919_not
g96037 not n43884 ; n43884_not
g96038 not n28629 ; n28629_not
g96039 not n49806 ; n49806_not
g96040 not n55683 ; n55683_not
g96041 not n29952 ; n29952_not
g96042 not n30969 ; n30969_not
g96043 not n45468 ; n45468_not
g96044 not n33885 ; n33885_not
g96045 not n50868 ; n50868_not
g96046 not n55890 ; n55890_not
g96047 not n49482 ; n49482_not
g96048 not n13689 ; n13689_not
g96049 not n28575 ; n28575_not
g96050 not n30978 ; n30978_not
g96051 not n49725 ; n49725_not
g96052 not n29970 ; n29970_not
g96053 not n54990 ; n54990_not
g96054 not n50877 ; n50877_not
g96055 not n13779 ; n13779_not
g96056 not n55674 ; n55674_not
g96057 not n28962 ; n28962_not
g96058 not n49626 ; n49626_not
g96059 not n28863 ; n28863_not
g96060 not n50967 ; n50967_not
g96061 not n49680 ; n49680_not
g96062 not n34983 ; n34983_not
g96063 not n45378 ; n45378_not
g96064 not n33975 ; n33975_not
g96065 not n43794 ; n43794_not
g96066 not n55863 ; n55863_not
g96067 not n49635 ; n49635_not
g96068 not n28980 ; n28980_not
g96069 not n41985 ; n41985_not
g96070 not n29916 ; n29916_not
g96071 not n34992 ; n34992_not
g96072 not n44982 ; n44982_not
g96073 not n28971 ; n28971_not
g96074 not n41967 ; n41967_not
g96075 not n49617 ; n49617_not
g96076 not n28845 ; n28845_not
g96077 not n44973 ; n44973_not
g96078 not n45387 ; n45387_not
g96079 not n13887 ; n13887_not
g96080 not n28944 ; n28944_not
g96081 not n49662 ; n49662_not
g96082 not n28953 ; n28953_not
g96083 not n55818 ; n55818_not
g96084 not n41895 ; n41895_not
g96085 not n49671 ; n49671_not
g96086 not n28881 ; n28881_not
g96087 not n49644 ; n49644_not
g96088 not n34875 ; n34875_not
g96089 not n45369 ; n45369_not
g96090 not n28908 ; n28908_not
g96091 not n49518 ; n49518_not
g96092 not n28917 ; n28917_not
g96093 not n55827 ; n55827_not
g96094 not n34974 ; n34974_not
g96095 not n49653 ; n49653_not
g96096 not n13896 ; n13896_not
g96097 not n34965 ; n34965_not
g96098 not n28935 ; n28935_not
g96099 not n33966 ; n33966_not
g96100 not n49563 ; n49563_not
g96101 not n41976 ; n41976_not
g96102 not n28737 ; n28737_not
g96103 not n49572 ; n49572_not
g96104 not n50787 ; n50787_not
g96105 not n55737 ; n55737_not
g96106 not n13869 ; n13869_not
g96107 not n28755 ; n28755_not
g96108 not n49581 ; n49581_not
g96109 not n29088 ; n29088_not
g96110 not n34884 ; n34884_not
g96111 not n54963 ; n54963_not
g96112 not n49707 ; n49707_not
g96113 not n40869 ; n40869_not
g96114 not n55728 ; n55728_not
g96115 not n14499 ; n14499_not
g96116 not n28719 ; n28719_not
g96117 not n34956 ; n34956_not
g96118 not n44946 ; n44946_not
g96119 not n29943 ; n29943_not
g96120 not n54954 ; n54954_not
g96121 not n28809 ; n28809_not
g96122 not n55764 ; n55764_not
g96123 not n44964 ; n44964_not
g96124 not n28827 ; n28827_not
g96125 not n43848 ; n43848_not
g96126 not n45396 ; n45396_not
g96127 not n49608 ; n49608_not
g96128 not n43839 ; n43839_not
g96129 not n55773 ; n55773_not
g96130 not n55746 ; n55746_not
g96131 not n55845 ; n55845_not
g96132 not n28773 ; n28773_not
g96133 not n55881 ; n55881_not
g96134 not n44955 ; n44955_not
g96135 not n49590 ; n49590_not
g96136 not n55836 ; n55836_not
g96137 not n54945 ; n54945_not
g96138 not n28791 ; n28791_not
g96139 not n55755 ; n55755_not
g96140 not n43866 ; n43866_not
g96141 not n29385 ; n29385_not
g96142 not n35487 ; n35487_not
g96143 not n49293 ; n49293_not
g96144 not n51579 ; n51579_not
g96145 not n28287 ; n28287_not
g96146 not n44847 ; n44847_not
g96147 not n55548 ; n55548_not
g96148 not n51588 ; n51588_not
g96149 not n29394 ; n29394_not
g96150 not n35478 ; n35478_not
g96151 not n33696 ; n33696_not
g96152 not n34398 ; n34398_not
g96153 not n45639 ; n45639_not
g96154 not n55980 ; n55980_not
g96155 not n35496 ; n35496_not
g96156 not n31599 ; n31599_not
g96157 not n49284 ; n49284_not
g96158 not n28269 ; n28269_not
g96159 not n16956 ; n16956_not
g96160 not n48537 ; n48537_not
g96161 not n33687 ; n33687_not
g96162 not n14976 ; n14976_not
g96163 not n49257 ; n49257_not
g96164 not n29376 ; n29376_not
g96165 not n35298 ; n35298_not
g96166 not n49248 ; n49248_not
g96167 not n55566 ; n55566_not
g96168 not n35397 ; n35397_not
g96169 not n49239 ; n49239_not
g96170 not n42696 ; n42696_not
g96171 not n56853 ; n56853_not
g96172 not n42687 ; n42687_not
g96173 not n35469 ; n35469_not
g96174 not n51597 ; n51597_not
g96175 not n55557 ; n55557_not
g96176 not n49275 ; n49275_not
g96177 not n39726 ; n39726_not
g96178 not n49266 ; n49266_not
g96179 not n27819 ; n27819_not
g96180 not n43686 ; n43686_not
g96181 not n45666 ; n45666_not
g96182 not n33669 ; n33669_not
g96183 not n29466 ; n29466_not
g96184 not n45657 ; n45657_not
g96185 not n43758 ; n43758_not
g96186 not n28179 ; n28179_not
g96187 not n42795 ; n42795_not
g96188 not n35685 ; n35685_not
g96189 not n34488 ; n34488_not
g96190 not n49428 ; n49428_not
g96191 not n12987 ; n12987_not
g96192 not n28188 ; n28188_not
g96193 not n44829 ; n44829_not
g96194 not n34857 ; n34857_not
g96195 not n42786 ; n42786_not
g96196 not n28197 ; n28197_not
g96197 not n45648 ; n45648_not
g96198 not n27909 ; n27909_not
g96199 not n35568 ; n35568_not
g96200 not n29439 ; n29439_not
g96201 not n29349 ; n29349_not
g96202 not n35559 ; n35559_not
g96203 not n44838 ; n44838_not
g96204 not n55539 ; n55539_not
g96205 not n29358 ; n29358_not
g96206 not n42759 ; n42759_not
g96207 not n51678 ; n51678_not
g96208 not n48546 ; n48546_not
g96209 not n35595 ; n35595_not
g96210 not n12996 ; n12996_not
g96211 not n42777 ; n42777_not
g96212 not n43767 ; n43767_not
g96213 not n51687 ; n51687_not
g96214 not n35586 ; n35586_not
g96215 not n42768 ; n42768_not
g96216 not n29457 ; n29457_not
g96217 not n29448 ; n29448_not
g96218 not n35577 ; n35577_not
g96219 not n42579 ; n42579_not
g96220 not n44883 ; n44883_not
g96221 not n55908 ; n55908_not
g96222 not n56763 ; n56763_not
g96223 not n55629 ; n55629_not
g96224 not n45279 ; n45279_not
g96225 not n29277 ; n29277_not
g96226 not n55917 ; n55917_not
g96227 not n43857 ; n43857_not
g96228 not n28485 ; n28485_not
g96229 not n29268 ; n29268_not
g96230 not n29286 ; n29286_not
g96231 not n49752 ; n49752_not
g96232 not n45549 ; n45549_not
g96233 not n49437 ; n49437_not
g96234 not n44991 ; n44991_not
g96235 not n49743 ; n49743_not
g96236 not n45288 ; n45288_not
g96237 not n29259 ; n29259_not
g96238 not n30987 ; n30987_not
g96239 not n44397 ; n44397_not
g96240 not n40599 ; n40599_not
g96241 not n44892 ; n44892_not
g96242 not n27864 ; n27864_not
g96243 not n40689 ; n40689_not
g96244 not n55638 ; n55638_not
g96245 not n40779 ; n40779_not
g96246 not n28377 ; n28377_not
g96247 not n55584 ; n55584_not
g96248 not n55935 ; n55935_not
g96249 not n28395 ; n28395_not
g96250 not n29925 ; n29925_not
g96251 not n44865 ; n44865_not
g96252 not n45576 ; n45576_not
g96253 not n35388 ; n35388_not
g96254 not n55926 ; n55926_not
g96255 not n55575 ; n55575_not
g96256 not n29367 ; n29367_not
g96257 not n45594 ; n45594_not
g96258 not n28359 ; n28359_not
g96259 not n35379 ; n35379_not
g96260 not n44856 ; n44856_not
g96261 not n49347 ; n49347_not
g96262 not n45585 ; n45585_not
g96263 not n42678 ; n42678_not
g96264 not n28467 ; n28467_not
g96265 not n29295 ; n29295_not
g96266 not n56808 ; n56808_not
g96267 not n49392 ; n49392_not
g96268 not n28296 ; n28296_not
g96269 not n44874 ; n44874_not
g96270 not n45558 ; n45558_not
g96271 not n42498 ; n42498_not
g96272 not n55593 ; n55593_not
g96273 not n28449 ; n28449_not
g96274 not n42588 ; n42588_not
g96275 not n45567 ; n45567_not
g96276 not n18783 ; n18783_not
g96277 not n47682 ; n47682_not
g96278 not n53586 ; n53586_not
g96279 not n45990 ; n45990_not
g96280 not n52875 ; n52875_not
g96281 not n18468 ; n18468_not
g96282 not n47673 ; n47673_not
g96283 not n53577 ; n53577_not
g96284 not n23679 ; n23679_not
g96285 not n18774 ; n18774_not
g96286 not n47664 ; n47664_not
g96287 not n52866 ; n52866_not
g96288 not n53568 ; n53568_not
g96289 not n47655 ; n47655_not
g96290 not n53559 ; n53559_not
g96291 not n18765 ; n18765_not
g96292 not n47646 ; n47646_not
g96293 not n52857 ; n52857_not
g96294 not n39159 ; n39159_not
g96295 not n47637 ; n47637_not
g96296 not n46575 ; n46575_not
g96297 not n39168 ; n39168_not
g96298 not n37476 ; n37476_not
g96299 not n47628 ; n47628_not
g96300 not n47736 ; n47736_not
g96301 not n47844 ; n47844_not
g96302 not n18828 ; n18828_not
g96303 not n45963 ; n45963_not
g96304 not n18819 ; n18819_not
g96305 not n47727 ; n47727_not
g96306 not n37494 ; n37494_not
g96307 not n47853 ; n47853_not
g96308 not n45972 ; n45972_not
g96309 not n47718 ; n47718_not
g96310 not n18792 ; n18792_not
g96311 not n45981 ; n45981_not
g96312 not n47709 ; n47709_not
g96313 not n46593 ; n46593_not
g96314 not n18459 ; n18459_not
g96315 not n52893 ; n52893_not
g96316 not n53595 ; n53595_not
g96317 not n23697 ; n23697_not
g96318 not n52884 ; n52884_not
g96319 not n47691 ; n47691_not
g96320 not n47871 ; n47871_not
g96321 not n23688 ; n23688_not
g96322 not n47565 ; n47565_not
g96323 not n24498 ; n24498_not
g96324 not n18675 ; n18675_not
g96325 not n47943 ; n47943_not
g96326 not n47556 ; n47556_not
g96327 not n24588 ; n24588_not
g96328 not n18666 ; n18666_not
g96329 not n47547 ; n47547_not
g96330 not n18657 ; n18657_not
g96331 not n46089 ; n46089_not
g96332 not n18648 ; n18648_not
g96333 not n47538 ; n47538_not
g96334 not n47529 ; n47529_not
g96335 not n47961 ; n47961_not
g96336 not n18639 ; n18639_not
g96337 not n36990 ; n36990_not
g96338 not n46098 ; n46098_not
g96339 not n18549 ; n18549_not
g96340 not n18558 ; n18558_not
g96341 not n54459 ; n54459_not
g96342 not n39249 ; n39249_not
g96343 not n24678 ; n24678_not
g96344 not n54468 ; n54468_not
g96345 not n18756 ; n18756_not
g96346 not n52848 ; n52848_not
g96347 not n18747 ; n18747_not
g96348 not n47619 ; n47619_not
g96349 not n37458 ; n37458_not
g96350 not n47916 ; n47916_not
g96351 not n18738 ; n18738_not
g96352 not n52839 ; n52839_not
g96353 not n46557 ; n46557_not
g96354 not n54396 ; n54396_not
g96355 not n39195 ; n39195_not
g96356 not n18729 ; n18729_not
g96357 not n18495 ; n18495_not
g96358 not n47592 ; n47592_not
g96359 not n54369 ; n54369_not
g96360 not n46548 ; n46548_not
g96361 not n24399 ; n24399_not
g96362 not n47583 ; n47583_not
g96363 not n36981 ; n36981_not
g96364 not n18693 ; n18693_not
g96365 not n47574 ; n47574_not
g96366 not n47934 ; n47934_not
g96367 not n18684 ; n18684_not
g96368 not n37638 ; n37638_not
g96369 not n53829 ; n53829_not
g96370 not n23976 ; n23976_not
g96371 not n18963 ; n18963_not
g96372 not n18954 ; n18954_not
g96373 not n18369 ; n18369_not
g96374 not n47349 ; n47349_not
g96375 not n47079 ; n47079_not
g96376 not n37629 ; n37629_not
g96377 not n52992 ; n52992_not
g96378 not n18945 ; n18945_not
g96379 not n18378 ; n18378_not
g96380 not n23985 ; n23985_not
g96381 not n53793 ; n53793_not
g96382 not n18936 ; n18936_not
g96383 not n46647 ; n46647_not
g96384 not n53784 ; n53784_not
g96385 not n52983 ; n52983_not
g96386 not n53775 ; n53775_not
g96387 not n46629 ; n46629_not
g96388 not n23994 ; n23994_not
g96389 not n45945 ; n45945_not
g96390 not n39069 ; n39069_not
g96391 not n52974 ; n52974_not
g96392 not n47097 ; n47097_not
g96393 not n18927 ; n18927_not
g96394 not n23868 ; n23868_not
g96395 not n37674 ; n37674_not
g96396 not n53946 ; n53946_not
g96397 not n53937 ; n53937_not
g96398 not n53928 ; n53928_not
g96399 not n23859 ; n23859_not
g96400 not n37665 ; n37665_not
g96401 not n53919 ; n53919_not
g96402 not n23949 ; n23949_not
g96403 not n53892 ; n53892_not
g96404 not n37656 ; n37656_not
g96405 not n18990 ; n18990_not
g96406 not n23958 ; n23958_not
g96407 not n53883 ; n53883_not
g96408 not n53874 ; n53874_not
g96409 not n54198 ; n54198_not
g96410 not n53865 ; n53865_not
g96411 not n37647 ; n37647_not
g96412 not n53856 ; n53856_not
g96413 not n23967 ; n23967_not
g96414 not n18981 ; n18981_not
g96415 not n53847 ; n53847_not
g96416 not n18972 ; n18972_not
g96417 not n53838 ; n53838_not
g96418 not n23778 ; n23778_not
g96419 not n47781 ; n47781_not
g96420 not n53685 ; n53685_not
g96421 not n37548 ; n37548_not
g96422 not n53676 ; n53676_not
g96423 not n47772 ; n47772_not
g96424 not n47826 ; n47826_not
g96425 not n37539 ; n37539_not
g96426 not n52929 ; n52929_not
g96427 not n18864 ; n18864_not
g96428 not n47763 ; n47763_not
g96429 not n53667 ; n53667_not
g96430 not n23769 ; n23769_not
g96431 not n47754 ; n47754_not
g96432 not n18855 ; n18855_not
g96433 not n53658 ; n53658_not
g96434 not n45954 ; n45954_not
g96435 not n18846 ; n18846_not
g96436 not n47745 ; n47745_not
g96437 not n53649 ; n53649_not
g96438 not n18837 ; n18837_not
g96439 not n37593 ; n37593_not
g96440 not n53766 ; n53766_not
g96441 not n52965 ; n52965_not
g96442 not n53757 ; n53757_not
g96443 not n46638 ; n46638_not
g96444 not n52578 ; n52578_not
g96445 not n39087 ; n39087_not
g96446 not n18918 ; n18918_not
g96447 not n53748 ; n53748_not
g96448 not n52956 ; n52956_not
g96449 not n37584 ; n37584_not
g96450 not n18909 ; n18909_not
g96451 not n53739 ; n53739_not
g96452 not n18891 ; n18891_not
g96453 not n52947 ; n52947_not
g96454 not n18882 ; n18882_not
g96455 not n37566 ; n37566_not
g96456 not n54288 ; n54288_not
g96457 not n47808 ; n47808_not
g96458 not n52587 ; n52587_not
g96459 not n23787 ; n23787_not
g96460 not n52938 ; n52938_not
g96461 not n18873 ; n18873_not
g96462 not n47790 ; n47790_not
g96463 not n53694 ; n53694_not
g96464 not n52596 ; n52596_not
g96465 not n54594 ; n54594_not
g96466 not n36756 ; n36756_not
g96467 not n46395 ; n46395_not
g96468 not n36765 ; n36765_not
g96469 not n18198 ; n18198_not
g96470 not n36774 ; n36774_not
g96471 not n17694 ; n17694_not
g96472 not n36783 ; n36783_not
g96473 not n24939 ; n24939_not
g96474 not n24948 ; n24948_not
g96475 not n18189 ; n18189_not
g96476 not n47439 ; n47439_not
g96477 not n36792 ; n36792_not
g96478 not n46359 ; n46359_not
g96479 not n36819 ; n36819_not
g96480 not n46377 ; n46377_not
g96481 not n47448 ; n47448_not
g96482 not n36828 ; n36828_not
g96483 not n39429 ; n39429_not
g96484 not n36837 ; n36837_not
g96485 not n17739 ; n17739_not
g96486 not n48159 ; n48159_not
g96487 not n17748 ; n17748_not
g96488 not n54639 ; n54639_not
g96489 not n36846 ; n36846_not
g96490 not n18099 ; n18099_not
g96491 not n24957 ; n24957_not
g96492 not n36855 ; n36855_not
g96493 not n47457 ; n47457_not
g96494 not n24876 ; n24876_not
g96495 not n46278 ; n46278_not
g96496 not n37188 ; n37188_not
g96497 not n18288 ; n18288_not
g96498 not n54558 ; n54558_not
g96499 not n37179 ; n37179_not
g96500 not n46287 ; n46287_not
g96501 not n39375 ; n39375_not
g96502 not n46296 ; n46296_not
g96503 not n18279 ; n18279_not
g96504 not n24885 ; n24885_not
g96505 not n24894 ; n24894_not
g96506 not n17649 ; n17649_not
g96507 not n36684 ; n36684_not
g96508 not n39384 ; n39384_not
g96509 not n54279 ; n54279_not
g96510 not n54567 ; n54567_not
g96511 not n36693 ; n36693_not
g96512 not n17658 ; n17658_not
g96513 not n24579 ; n24579_not
g96514 not n39393 ; n39393_not
g96515 not n54576 ; n54576_not
g96516 not n36729 ; n36729_not
g96517 not n36738 ; n36738_not
g96518 not n54585 ; n54585_not
g96519 not n36747 ; n36747_not
g96520 not n17685 ; n17685_not
g96521 not n37098 ; n37098_not
g96522 not n54666 ; n54666_not
g96523 not n52677 ; n52677_not
g96524 not n24489 ; n24489_not
g96525 not n47493 ; n47493_not
g96526 not n52668 ; n52668_not
g96527 not n36927 ; n36927_not
g96528 not n39465 ; n39465_not
g96529 not n17784 ; n17784_not
g96530 not n36936 ; n36936_not
g96531 not n54675 ; n54675_not
g96532 not n17793 ; n17793_not
g96533 not n54684 ; n54684_not
g96534 not n36945 ; n36945_not
g96535 not n39474 ; n39474_not
g96536 not n54693 ; n54693_not
g96537 not n36954 ; n36954_not
g96538 not n17991 ; n17991_not
g96539 not n17982 ; n17982_not
g96540 not n36963 ; n36963_not
g96541 not n39483 ; n39483_not
g96542 not n39438 ; n39438_not
g96543 not n36864 ; n36864_not
g96544 not n46368 ; n46368_not
g96545 not n48168 ; n48168_not
g96546 not n36873 ; n36873_not
g96547 not n24966 ; n24966_not
g96548 not n47466 ; n47466_not
g96549 not n24975 ; n24975_not
g96550 not n36882 ; n36882_not
g96551 not n24984 ; n24984_not
g96552 not n48177 ; n48177_not
g96553 not n36891 ; n36891_not
g96554 not n39447 ; n39447_not
g96555 not n52695 ; n52695_not
g96556 not n24993 ; n24993_not
g96557 not n47475 ; n47475_not
g96558 not n54648 ; n54648_not
g96559 not n48186 ; n48186_not
g96560 not n39456 ; n39456_not
g96561 not n36909 ; n36909_not
g96562 not n54657 ; n54657_not
g96563 not n47484 ; n47484_not
g96564 not n17775 ; n17775_not
g96565 not n36918 ; n36918_not
g96566 not n48195 ; n48195_not
g96567 not n17892 ; n17892_not
g96568 not n37368 ; n37368_not
g96569 not n17919 ; n17919_not
g96570 not n24669 ; n24669_not
g96571 not n37359 ; n37359_not
g96572 not n54495 ; n54495_not
g96573 not n52776 ; n52776_not
g96574 not n39294 ; n39294_not
g96575 not n17928 ; n17928_not
g96576 not n52686 ; n52686_not
g96577 not n24759 ; n24759_not
g96578 not n17937 ; n17937_not
g96579 not n17946 ; n17946_not
g96580 not n24768 ; n24768_not
g96581 not n17955 ; n17955_not
g96582 not n46179 ; n46179_not
g96583 not n46485 ; n46485_not
g96584 not n47394 ; n47394_not
g96585 not n17964 ; n17964_not
g96586 not n17973 ; n17973_not
g96587 not n52767 ; n52767_not
g96588 not n47385 ; n47385_not
g96589 not n46188 ; n46188_not
g96590 not n37395 ; n37395_not
g96591 not n39258 ; n39258_not
g96592 not n18594 ; n18594_not
g96593 not n52794 ; n52794_not
g96594 not n39267 ; n39267_not
g96595 not n24696 ; n24696_not
g96596 not n39276 ; n39276_not
g96597 not n52785 ; n52785_not
g96598 not n54477 ; n54477_not
g96599 not n37386 ; n37386_not
g96600 not n18576 ; n18576_not
g96601 not n39285 ; n39285_not
g96602 not n37377 ; n37377_not
g96603 not n54486 ; n54486_not
g96604 not n18567 ; n18567_not
g96605 not n48078 ; n48078_not
g96606 not n37089 ; n37089_not
g96607 not n47376 ; n47376_not
g96608 not n39339 ; n39339_not
g96609 not n24795 ; n24795_not
g96610 not n39078 ; n39078_not
g96611 not n48087 ; n48087_not
g96612 not n52749 ; n52749_not
g96613 not n39348 ; n39348_not
g96614 not n18297 ; n18297_not
g96615 not n39357 ; n39357_not
g96616 not n24849 ; n24849_not
g96617 not n48096 ; n48096_not
g96618 not n54549 ; n54549_not
g96619 not n24858 ; n24858_not
g96620 not n46269 ; n46269_not
g96621 not n24867 ; n24867_not
g96622 not n37197 ; n37197_not
g96623 not n39366 ; n39366_not
g96624 not n24777 ; n24777_not
g96625 not n37296 ; n37296_not
g96626 not n47367 ; n47367_not
g96627 not n37287 ; n37287_not
g96628 not n47358 ; n47358_not
g96629 not n46197 ; n46197_not
g96630 not n18477 ; n18477_not
g96631 not n46656 ; n46656_not
g96632 not n24786 ; n24786_not
g96633 not n37278 ; n37278_not
g96634 not n37269 ; n37269_not
g96635 not n46467 ; n46467_not
g96636 not n48069 ; n48069_not
g96637 not n52758 ; n52758_not
g96638 not n46458 ; n46458_not
g96639 not n18387 ; n18387_not
g96640 not n20979 ; n20979_not
g96641 not n38628 ; n38628_not
g96642 not n20988 ; n20988_not
g96643 not n46683 ; n46683_not
g96644 not n19575 ; n19575_not
g96645 not n20997 ; n20997_not
g96646 not n53388 ; n53388_not
g96647 not n38682 ; n38682_not
g96648 not n19584 ; n19584_not
g96649 not n46692 ; n46692_not
g96650 not n19593 ; n19593_not
g96651 not n19854 ; n19854_not
g96652 not n19845 ; n19845_not
g96653 not n38619 ; n38619_not
g96654 not n38691 ; n38691_not
g96655 not n37980 ; n37980_not
g96656 not n19629 ; n19629_not
g96657 not n19638 ; n19638_not
g96658 not n19827 ; n19827_not
g96659 not n37971 ; n37971_not
g96660 not n38637 ; n38637_not
g96661 not n19476 ; n19476_not
g96662 not n20889 ; n20889_not
g96663 not n19917 ; n19917_not
g96664 not n46674 ; n46674_not
g96665 not n20898 ; n20898_not
g96666 not n38655 ; n38655_not
g96667 not n19485 ; n19485_not
g96668 not n46665 ; n46665_not
g96669 not n19494 ; n19494_not
g96670 not n38664 ; n38664_not
g96671 not n19890 ; n19890_not
g96672 not n19539 ; n19539_not
g96673 not n19548 ; n19548_not
g96674 not n38673 ; n38673_not
g96675 not n19557 ; n19557_not
g96676 not n19872 ; n19872_not
g96677 not n19566 ; n19566_not
g96678 not n38745 ; n38745_not
g96679 not n21699 ; n21699_not
g96680 not n37935 ; n37935_not
g96681 not n46764 ; n46764_not
g96682 not n47286 ; n47286_not
g96683 not n53298 ; n53298_not
g96684 not n37926 ; n37926_not
g96685 not n46773 ; n46773_not
g96686 not n47277 ; n47277_not
g96687 not n21789 ; n21789_not
g96688 not n37917 ; n37917_not
g96689 not n37467 ; n37467_not
g96690 not n38754 ; n38754_not
g96691 not n21798 ; n21798_not
g96692 not n19719 ; n19719_not
g96693 not n46782 ; n46782_not
g96694 not n37908 ; n37908_not
g96695 not n19782 ; n19782_not
g96696 not n21879 ; n21879_not
g96697 not n38583 ; n38583_not
g96698 not n21888 ; n21888_not
g96699 not n46719 ; n46719_not
g96700 not n38709 ; n38709_not
g96701 not n19647 ; n19647_not
g96702 not n38718 ; n38718_not
g96703 not n19656 ; n19656_not
g96704 not n46728 ; n46728_not
g96705 not n38727 ; n38727_not
g96706 not n19665 ; n19665_not
g96707 not n46737 ; n46737_not
g96708 not n19674 ; n19674_not
g96709 not n19809 ; n19809_not
g96710 not n37953 ; n37953_not
g96711 not n20799 ; n20799_not
g96712 not n38736 ; n38736_not
g96713 not n46746 ; n46746_not
g96714 not n19683 ; n19683_not
g96715 not n19692 ; n19692_not
g96716 not n37944 ; n37944_not
g96717 not n46755 ; n46755_not
g96718 not n19953 ; n19953_not
g96719 not n46917 ; n46917_not
g96720 not n46908 ; n46908_not
g96721 not n38079 ; n38079_not
g96722 not n47088 ; n47088_not
g96723 not n46890 ; n46890_not
g96724 not n53496 ; n53496_not
g96725 not n19980 ; n19980_not
g96726 not n46881 ; n46881_not
g96727 not n46872 ; n46872_not
g96728 not n19818 ; n19818_not
g96729 not n46863 ; n46863_not
g96730 not n38457 ; n38457_not
g96731 not n46854 ; n46854_not
g96732 not n38466 ; n38466_not
g96733 not n46845 ; n46845_not
g96734 not n19908 ; n19908_not
g96735 not n46980 ; n46980_not
g96736 not n46971 ; n46971_not
g96737 not n19863 ; n19863_not
g96738 not n46962 ; n46962_not
g96739 not n46953 ; n46953_not
g96740 not n19935 ; n19935_not
g96741 not n46944 ; n46944_not
g96742 not n47178 ; n47178_not
g96743 not n46935 ; n46935_not
g96744 not n47187 ; n47187_not
g96745 not n46926 ; n46926_not
g96746 not n19944 ; n19944_not
g96747 not n19395 ; n19395_not
g96748 not n38529 ; n38529_not
g96749 not n53469 ; n53469_not
g96750 not n38547 ; n38547_not
g96751 not n19962 ; n19962_not
g96752 not n47295 ; n47295_not
g96753 not n38565 ; n38565_not
g96754 not n38088 ; n38088_not
g96755 not n38574 ; n38574_not
g96756 not n19449 ; n19449_not
g96757 not n38592 ; n38592_not
g96758 not n19458 ; n19458_not
g96759 not n19467 ; n19467_not
g96760 not n46836 ; n46836_not
g96761 not n46386 ; n46386_not
g96762 not n53478 ; n53478_not
g96763 not n46827 ; n46827_not
g96764 not n38475 ; n38475_not
g96765 not n38484 ; n38484_not
g96766 not n46818 ; n46818_not
g96767 not n46809 ; n46809_not
g96768 not n19359 ; n19359_not
g96769 not n19368 ; n19368_not
g96770 not n46791 ; n46791_not
g96771 not n19377 ; n19377_not
g96772 not n47268 ; n47268_not
g96773 not n19386 ; n19386_not
g96774 not n19773 ; n19773_not
g96775 not n22959 ; n22959_not
g96776 not n53991 ; n53991_not
g96777 not n53289 ; n53289_not
g96778 not n37755 ; n37755_not
g96779 not n22599 ; n22599_not
g96780 not n37557 ; n37557_not
g96781 not n22887 ; n22887_not
g96782 not n37746 ; n37746_not
g96783 not n22878 ; n22878_not
g96784 not n38907 ; n38907_not
g96785 not n22869 ; n22869_not
g96786 not n22689 ; n22689_not
g96787 not n38862 ; n38862_not
g96788 not n22986 ; n22986_not
g96789 not n53955 ; n53955_not
g96790 not n52488 ; n52488_not
g96791 not n37782 ; n37782_not
g96792 not n38871 ; n38871_not
g96793 not n19188 ; n19188_not
g96794 not n47196 ; n47196_not
g96795 not n53964 ; n53964_not
g96796 not n53973 ; n53973_not
g96797 not n22977 ; n22977_not
g96798 not n22968 ; n22968_not
g96799 not n37773 ; n37773_not
g96800 not n38880 ; n38880_not
g96801 not n53982 ; n53982_not
g96802 not n52497 ; n52497_not
g96803 not n19197 ; n19197_not
g96804 not n37764 ; n37764_not
g96805 not n38952 ; n38952_not
g96806 not n46566 ; n46566_not
g96807 not n38961 ; n38961_not
g96808 not n23796 ; n23796_not
g96809 not n37692 ; n37692_not
g96810 not n23886 ; n23886_not
g96811 not n37683 ; n37683_not
g96812 not n23877 ; n23877_not
g96813 not n19098 ; n19098_not
g96814 not n38916 ; n38916_not
g96815 not n38493 ; n38493_not
g96816 not n37737 ; n37737_not
g96817 not n22698 ; n22698_not
g96818 not n19278 ; n19278_not
g96819 not n38925 ; n38925_not
g96820 not n23499 ; n23499_not
g96821 not n19287 ; n19287_not
g96822 not n22779 ; n22779_not
g96823 not n37728 ; n37728_not
g96824 not n22797 ; n22797_not
g96825 not n19296 ; n19296_not
g96826 not n22788 ; n22788_not
g96827 not n38934 ; n38934_not
g96828 not n23589 ; n23589_not
g96829 not n23598 ; n23598_not
g96830 not n37719 ; n37719_not
g96831 not n38943 ; n38943_not
g96832 not n37872 ; n37872_not
g96833 not n53199 ; n53199_not
g96834 not n37863 ; n37863_not
g96835 not n21897 ; n21897_not
g96836 not n38763 ; n38763_not
g96837 not n19728 ; n19728_not
g96838 not n19737 ; n19737_not
g96839 not n21969 ; n21969_not
g96840 not n21978 ; n21978_not
g96841 not n21987 ; n21987_not
g96842 not n38772 ; n38772_not
g96843 not n21996 ; n21996_not
g96844 not n19746 ; n19746_not
g96845 not n37890 ; n37890_not
g96846 not n46476 ; n46476_not
g96847 not n38781 ; n38781_not
g96848 not n37881 ; n37881_not
g96849 not n53379 ; n53379_not
g96850 not n38808 ; n38808_not
g96851 not n37809 ; n37809_not
g96852 not n38817 ; n38817_not
g96853 not n38826 ; n38826_not
g96854 not n38835 ; n38835_not
g96855 not n22896 ; n22896_not
g96856 not n38538 ; n38538_not
g96857 not n38844 ; n38844_not
g96858 not n37791 ; n37791_not
g96859 not n38853 ; n38853_not
g96860 not n37854 ; n37854_not
g96861 not n38790 ; n38790_not
g96862 not n37845 ; n37845_not
g96863 not n37836 ; n37836_not
g96864 not n37827 ; n37827_not
g96865 not n37818 ; n37818_not
g96866 not n17478 ; n17478_not
g96867 not n26289 ; n26289_not
g96868 not n36675 ; n36675_not
g96869 not n17469 ; n17469_not
g96870 not n47817 ; n47817_not
g96871 not n54972 ; n54972_not
g96872 not n39708 ; n39708_not
g96873 not n36297 ; n36297_not
g96874 not n16848 ; n16848_not
g96875 not n25974 ; n25974_not
g96876 not n17496 ; n17496_not
g96877 not n48474 ; n48474_not
g96878 not n25983 ; n25983_not
g96879 not n25992 ; n25992_not
g96880 not n48483 ; n48483_not
g96881 not n16839 ; n16839_not
g96882 not n17487 ; n17487_not
g96883 not n26199 ; n26199_not
g96884 not n39717 ; n39717_not
g96885 not n48492 ; n48492_not
g96886 not n48528 ; n48528_not
g96887 not n17388 ; n17388_not
g96888 not n17379 ; n17379_not
g96889 not n48555 ; n48555_not
g96890 not n48519 ; n48519_not
g96891 not n36639 ; n36639_not
g96892 not n36288 ; n36288_not
g96893 not n45819 ; n45819_not
g96894 not n36279 ; n36279_not
g96895 not n36648 ; n36648_not
g96896 not n36657 ; n36657_not
g96897 not n17397 ; n17397_not
g96898 not n25794 ; n25794_not
g96899 not n36396 ; n36396_not
g96900 not n54099 ; n54099_not
g96901 not n54891 ; n54891_not
g96902 not n39663 ; n39663_not
g96903 not n16929 ; n16929_not
g96904 not n17577 ; n17577_not
g96905 not n25839 ; n25839_not
g96906 not n36387 ; n36387_not
g96907 not n16974 ; n16974_not
g96908 not n17568 ; n17568_not
g96909 not n25848 ; n25848_not
g96910 not n36378 ; n36378_not
g96911 not n25857 ; n25857_not
g96912 not n17559 ; n17559_not
g96913 not n16983 ; n16983_not
g96914 not n48375 ; n48375_not
g96915 not n54873 ; n54873_not
g96916 not n25749 ; n25749_not
g96917 not n17595 ; n17595_not
g96918 not n25758 ; n25758_not
g96919 not n48384 ; n48384_not
g96920 not n45774 ; n45774_not
g96921 not n16947 ; n16947_not
g96922 not n25767 ; n25767_not
g96923 not n39654 ; n39654_not
g96924 not n25389 ; n25389_not
g96925 not n25776 ; n25776_not
g96926 not n16938 ; n16938_not
g96927 not n54882 ; n54882_not
g96928 not n48393 ; n48393_not
g96929 not n25785 ; n25785_not
g96930 not n17586 ; n17586_not
g96931 not n48447 ; n48447_not
g96932 not n16875 ; n16875_not
g96933 not n25929 ; n25929_not
g96934 not n25299 ; n25299_not
g96935 not n16866 ; n16866_not
g96936 not n25938 ; n25938_not
g96937 not n48456 ; n48456_not
g96938 not n54927 ; n54927_not
g96939 not n25947 ; n25947_not
g96940 not n16857 ; n16857_not
g96941 not n25956 ; n25956_not
g96942 not n26919 ; n26919_not
g96943 not n48465 ; n48465_not
g96944 not n25965 ; n25965_not
g96945 not n25866 ; n25866_not
g96946 not n47862 ; n47862_not
g96947 not n36594 ; n36594_not
g96948 not n48429 ; n48429_not
g96949 not n36369 ; n36369_not
g96950 not n16992 ; n16992_not
g96951 not n39681 ; n39681_not
g96952 not n25875 ; n25875_not
g96953 not n54909 ; n54909_not
g96954 not n16893 ; n16893_not
g96955 not n48438 ; n48438_not
g96956 not n25884 ; n25884_not
g96957 not n16884 ; n16884_not
g96958 not n25893 ; n25893_not
g96959 not n54918 ; n54918_not
g96960 not n48735 ; n48735_not
g96961 not n36495 ; n36495_not
g96962 not n48690 ; n48690_not
g96963 not n48807 ; n48807_not
g96964 not n36198 ; n36198_not
g96965 not n26964 ; n26964_not
g96966 not n35766 ; n35766_not
g96967 not n45909 ; n45909_not
g96968 not n48780 ; n48780_not
g96969 not n17199 ; n17199_not
g96970 not n17298 ; n17298_not
g96971 not n17289 ; n17289_not
g96972 not n36666 ; n36666_not
g96973 not n36459 ; n36459_not
g96974 not n39672 ; n39672_not
g96975 not n36468 ; n36468_not
g96976 not n36477 ; n36477_not
g96977 not n36486 ; n36486_not
g96978 not n45864 ; n45864_not
g96979 not n48645 ; n48645_not
g96980 not n36576 ; n36576_not
g96981 not n51696 ; n51696_not
g96982 not n36558 ; n36558_not
g96983 not n36549 ; n36549_not
g96984 not n25587 ; n25587_not
g96985 not n25578 ; n25578_not
g96986 not n54828 ; n54828_not
g96987 not n25569 ; n25569_not
g96988 not n17865 ; n17865_not
g96989 not n48294 ; n48294_not
g96990 not n17847 ; n17847_not
g96991 not n17829 ; n17829_not
g96992 not n54819 ; n54819_not
g96993 not n54846 ; n54846_not
g96994 not n47907 ; n47907_not
g96995 not n36567 ; n36567_not
g96996 not n48348 ; n48348_not
g96997 not n25659 ; n25659_not
g96998 not n54855 ; n54855_not
g96999 not n25668 ; n25668_not
g97000 not n17757 ; n17757_not
g97001 not n54837 ; n54837_not
g97002 not n39591 ; n39591_not
g97003 not n25596 ; n25596_not
g97004 not n25479 ; n25479_not
g97005 not n48339 ; n48339_not
g97006 not n48258 ; n48258_not
g97007 not n54765 ; n54765_not
g97008 not n54756 ; n54756_not
g97009 not n48249 ; n48249_not
g97010 not n54747 ; n54747_not
g97011 not n17838 ; n17838_not
g97012 not n36972 ; n36972_not
g97013 not n25398 ; n25398_not
g97014 not n54189 ; n54189_not
g97015 not n54729 ; n54729_not
g97016 not n39492 ; n39492_not
g97017 not n54738 ; n54738_not
g97018 not n39546 ; n39546_not
g97019 not n48276 ; n48276_not
g97020 not n54783 ; n54783_not
g97021 not n54792 ; n54792_not
g97022 not n48285 ; n48285_not
g97023 not n17874 ; n17874_not
g97024 not n39519 ; n39519_not
g97025 not n54774 ; n54774_not
g97026 not n47952 ; n47952_not
g97027 not n48267 ; n48267_not
g97028 not n25488 ; n25488_not
g97029 not n45729 ; n45729_not
g97030 not n25677 ; n25677_not
g97031 not n25686 ; n25686_not
g97032 not n48357 ; n48357_not
g97033 not n17667 ; n17667_not
g97034 not n48366 ; n48366_not
g97035 not n39636 ; n39636_not
g97036 not n25695 ; n25695_not
g97037 not n54864 ; n54864_not
g97038 not n51868 ; n51868_not
g97039 not n23995 ; n23995_not
g97040 not n51697 ; n51697_not
g97041 not n56476 ; n56476_not
g97042 not n14599 ; n14599_not
g97043 not n51994 ; n51994_not
g97044 not n28657 ; n28657_not
g97045 not n55837 ; n55837_not
g97046 not n56467 ; n56467_not
g97047 not n16696 ; n16696_not
g97048 not n13699 ; n13699_not
g97049 not n26749 ; n26749_not
g97050 not n56458 ; n56458_not
g97051 not n28468 ; n28468_not
g97052 not n18649 ; n18649_not
g97053 not n56818 ; n56818_not
g97054 not n14788 ; n14788_not
g97055 not n28648 ; n28648_not
g97056 not n51985 ; n51985_not
g97057 not n55288 ; n55288_not
g97058 not n20998 ; n20998_not
g97059 not n16399 ; n16399_not
g97060 not n56449 ; n56449_not
g97061 not n53389 ; n53389_not
g97062 not n21997 ; n21997_not
g97063 not n30997 ; n30997_not
g97064 not n26785 ; n26785_not
g97065 not n24949 ; n24949_not
g97066 not n54973 ; n54973_not
g97067 not n56755 ; n56755_not
g97068 not n56548 ; n56548_not
g97069 not n26776 ; n26776_not
g97070 not n56539 ; n56539_not
g97071 not n16687 ; n16687_not
g97072 not n14896 ; n14896_not
g97073 not n51886 ; n51886_not
g97074 not n51967 ; n51967_not
g97075 not n19774 ; n19774_not
g97076 not n14869 ; n14869_not
g97077 not n56773 ; n56773_not
g97078 not n26767 ; n26767_not
g97079 not n24598 ; n24598_not
g97080 not n18658 ; n18658_not
g97081 not n51877 ; n51877_not
g97082 not n56494 ; n56494_not
g97083 not n26758 ; n26758_not
g97084 not n30979 ; n30979_not
g97085 not n51976 ; n51976_not
g97086 not n56485 ; n56485_not
g97087 not n54784 ; n54784_not
g97088 not n27487 ; n27487_not
g97089 not n56791 ; n56791_not
g97090 not n16768 ; n16768_not
g97091 not n55684 ; n55684_not
g97092 not n26668 ; n26668_not
g97093 not n20899 ; n20899_not
g97094 not n24958 ; n24958_not
g97095 not n25696 ; n25696_not
g97096 not n26659 ; n26659_not
g97097 not n16777 ; n16777_not
g97098 not n20989 ; n20989_not
g97099 not n56881 ; n56881_not
g97100 not n56890 ; n56890_not
g97101 not n31699 ; n31699_not
g97102 not n24967 ; n24967_not
g97103 not n16849 ; n16849_not
g97104 not n16795 ; n16795_not
g97105 not n16786 ; n16786_not
g97106 not n56269 ; n56269_not
g97107 not n24976 ; n24976_not
g97108 not n14887 ; n14887_not
g97109 not n56908 ; n56908_not
g97110 not n16489 ; n16489_not
g97111 not n56278 ; n56278_not
g97112 not n56287 ; n56287_not
g97113 not n19819 ; n19819_not
g97114 not n29098 ; n29098_not
g97115 not n56296 ; n56296_not
g97116 not n55279 ; n55279_not
g97117 not n52786 ; n52786_not
g97118 not n19792 ; n19792_not
g97119 not n16759 ; n16759_not
g97120 not n55693 ; n55693_not
g97121 not n56836 ; n56836_not
g97122 not n54775 ; n54775_not
g97123 not n56395 ; n56395_not
g97124 not n25768 ; n25768_not
g97125 not n55099 ; n55099_not
g97126 not n14797 ; n14797_not
g97127 not n56845 ; n56845_not
g97128 not n56386 ; n56386_not
g97129 not n26677 ; n26677_not
g97130 not n56863 ; n56863_not
g97131 not n23986 ; n23986_not
g97132 not n26686 ; n26686_not
g97133 not n17749 ; n17749_not
g97134 not n13897 ; n13897_not
g97135 not n56359 ; n56359_not
g97136 not n27919 ; n27919_not
g97137 not n56368 ; n56368_not
g97138 not n26695 ; n26695_not
g97139 not n28639 ; n28639_not
g97140 not n56377 ; n56377_not
g97141 not n27667 ; n27667_not
g97142 not n28477 ; n28477_not
g97143 not n27739 ; n27739_not
g97144 not n18685 ; n18685_not
g97145 not n28684 ; n28684_not
g97146 not n16579 ; n16579_not
g97147 not n15994 ; n15994_not
g97148 not n17659 ; n17659_not
g97149 not n21988 ; n21988_not
g97150 not n56674 ; n56674_not
g97151 not n26866 ; n26866_not
g97152 not n16588 ; n16588_not
g97153 not n21979 ; n21979_not
g97154 not n26956 ; n26956_not
g97155 not n26857 ; n26857_not
g97156 not n56683 ; n56683_not
g97157 not n17668 ; n17668_not
g97158 not n52678 ; n52678_not
g97159 not n26965 ; n26965_not
g97160 not n18676 ; n18676_not
g97161 not n56665 ; n56665_not
g97162 not n17587 ; n17587_not
g97163 not n54577 ; n54577_not
g97164 not n54883 ; n54883_not
g97165 not n26848 ; n26848_not
g97166 not n21898 ; n21898_not
g97167 not n29188 ; n29188_not
g97168 not n55594 ; n55594_not
g97169 not n56656 ; n56656_not
g97170 not n16597 ; n16597_not
g97171 not n56647 ; n56647_not
g97172 not n52597 ; n52597_not
g97173 not n17839 ; n17839_not
g97174 not n30898 ; n30898_not
g97175 not n24886 ; n24886_not
g97176 not n26893 ; n26893_not
g97177 not n51895 ; n51895_not
g97178 not n22789 ; n22789_not
g97179 not n15976 ; n15976_not
g97180 not n56629 ; n56629_not
g97181 not n24895 ; n24895_not
g97182 not n56638 ; n56638_not
g97183 not n27946 ; n27946_not
g97184 not n17857 ; n17857_not
g97185 not n50689 ; n50689_not
g97186 not n25786 ; n25786_not
g97187 not n22798 ; n22798_not
g97188 not n54568 ; n54568_not
g97189 not n15985 ; n15985_not
g97190 not n26884 ; n26884_not
g97191 not n28396 ; n28396_not
g97192 not n28693 ; n28693_not
g97193 not n26947 ; n26947_not
g97194 not n50698 ; n50698_not
g97195 not n26875 ; n26875_not
g97196 not n24589 ; n24589_not
g97197 not n55792 ; n55792_not
g97198 not n55297 ; n55297_not
g97199 not n21799 ; n21799_not
g97200 not n28666 ; n28666_not
g97201 not n51949 ; n51949_not
g97202 not n27685 ; n27685_not
g97203 not n54793 ; n54793_not
g97204 not n56584 ; n56584_not
g97205 not n16678 ; n16678_not
g97206 not n21889 ; n21889_not
g97207 not n54478 ; n54478_not
g97208 not n26992 ; n26992_not
g97209 not n56575 ; n56575_not
g97210 not n14779 ; n14779_not
g97211 not n26794 ; n26794_not
g97212 not n56566 ; n56566_not
g97213 not n25498 ; n25498_not
g97214 not n56746 ; n56746_not
g97215 not n30988 ; n30988_not
g97216 not n19765 ; n19765_not
g97217 not n51958 ; n51958_not
g97218 not n56557 ; n56557_not
g97219 not n54586 ; n54586_not
g97220 not n26839 ; n26839_not
g97221 not n51688 ; n51688_not
g97222 not n55189 ; n55189_not
g97223 not n15697 ; n15697_not
g97224 not n55828 ; n55828_not
g97225 not n27964 ; n27964_not
g97226 not n25777 ; n25777_not
g97227 not n54964 ; n54964_not
g97228 not n54595 ; n54595_not
g97229 not n17875 ; n17875_not
g97230 not n16669 ; n16669_not
g97231 not n29269 ; n29269_not
g97232 not n18667 ; n18667_not
g97233 not n27469 ; n27469_not
g97234 not n55198 ; n55198_not
g97235 not n56728 ; n56728_not
g97236 not n14878 ; n14878_not
g97237 not n28675 ; n28675_not
g97238 not n17695 ; n17695_not
g97239 not n28459 ; n28459_not
g97240 not n56593 ; n56593_not
g97241 not n54739 ; n54739_not
g97242 not n55657 ; n55657_not
g97243 not n14698 ; n14698_not
g97244 not n19990 ; n19990_not
g97245 not n54676 ; n54676_not
g97246 not n27649 ; n27649_not
g97247 not n24688 ; n24688_not
g97248 not n29089 ; n29089_not
g97249 not n19297 ; n19297_not
g97250 not n53488 ; n53488_not
g97251 not n55648 ; n55648_not
g97252 not n57286 ; n57286_not
g97253 not n54874 ; n54874_not
g97254 not n24697 ; n24697_not
g97255 not n54469 ; n54469_not
g97256 not n54685 ; n54685_not
g97257 not n31996 ; n31996_not
g97258 not n17794 ; n17794_not
g97259 not n26497 ; n26497_not
g97260 not n25399 ; n25399_not
g97261 not n54667 ; n54667_not
g97262 not n14689 ; n14689_not
g97263 not n17785 ; n17785_not
g97264 not n26569 ; n26569_not
g97265 not n50788 ; n50788_not
g97266 not n19972 ; n19972_not
g97267 not n26578 ; n26578_not
g97268 not n26596 ; n26596_not
g97269 not n56854 ; n56854_not
g97270 not n28495 ; n28495_not
g97271 not n53479 ; n53479_not
g97272 not n57268 ; n57268_not
g97273 not n27586 ; n27586_not
g97274 not n26587 ; n26587_not
g97275 not n18595 ; n18595_not
g97276 not n19783 ; n19783_not
g97277 not n26929 ; n26929_not
g97278 not n57259 ; n57259_not
g97279 not n56935 ; n56935_not
g97280 not n56944 ; n56944_not
g97281 not n13879 ; n13879_not
g97282 not n51787 ; n51787_not
g97283 not n19855 ; n19855_not
g97284 not n54199 ; n54199_not
g97285 not n57457 ; n57457_not
g97286 not n56971 ; n56971_not
g97287 not n17596 ; n17596_not
g97288 not n19864 ; n19864_not
g97289 not n57466 ; n57466_not
g97290 not n51778 ; n51778_not
g97291 not n55855 ; n55855_not
g97292 not n57475 ; n57475_not
g97293 not n56980 ; n56980_not
g97294 not n19918 ; n19918_not
g97295 not n16957 ; n16957_not
g97296 not n19873 ; n19873_not
g97297 not n19909 ; n19909_not
g97298 not n57484 ; n57484_not
g97299 not n26974 ; n26974_not
g97300 not n55639 ; n55639_not
g97301 not n19828 ; n19828_not
g97302 not n19963 ; n19963_not
g97303 not n19954 ; n19954_not
g97304 not n27874 ; n27874_not
g97305 not n52795 ; n52795_not
g97306 not n57394 ; n57394_not
g97307 not n54694 ; n54694_not
g97308 not n56926 ; n56926_not
g97309 not n19945 ; n19945_not
g97310 not n57385 ; n57385_not
g97311 not n51796 ; n51796_not
g97312 not n50797 ; n50797_not
g97313 not n57358 ; n57358_not
g97314 not n54766 ; n54766_not
g97315 not n56179 ; n56179_not
g97316 not n54865 ; n54865_not
g97317 not n31789 ; n31789_not
g97318 not n23968 ; n23968_not
g97319 not n53398 ; n53398_not
g97320 not n27559 ; n27559_not
g97321 not n28585 ; n28585_not
g97322 not n16876 ; n16876_not
g97323 not n13789 ; n13789_not
g97324 not n16885 ; n16885_not
g97325 not n54757 ; n54757_not
g97326 not n28576 ; n28576_not
g97327 not n19882 ; n19882_not
g97328 not n24994 ; n24994_not
g97329 not n16993 ; n16993_not
g97330 not n26488 ; n26488_not
g97331 not n54649 ; n54649_not
g97332 not n16894 ; n16894_not
g97333 not n26479 ; n26479_not
g97334 not n56719 ; n56719_not
g97335 not n27568 ; n27568_not
g97336 not n17758 ; n17758_not
g97337 not n23977 ; n23977_not
g97338 not n19837 ; n19837_not
g97339 not n50887 ; n50887_not
g97340 not n16858 ; n16858_not
g97341 not n55882 ; n55882_not
g97342 not n28594 ; n28594_not
g97343 not n55675 ; n55675_not
g97344 not n50878 ; n50878_not
g97345 not n18577 ; n18577_not
g97346 not n56188 ; n56188_not
g97347 not n16867 ; n16867_not
g97348 not n56953 ; n56953_not
g97349 not n24985 ; n24985_not
g97350 not n56197 ; n56197_not
g97351 not n16498 ; n16498_not
g97352 not n31798 ; n31798_not
g97353 not n23959 ; n23959_not
g97354 not n27199 ; n27199_not
g97355 not n55873 ; n55873_not
g97356 not n24499 ; n24499_not
g97357 not n54748 ; n54748_not
g97358 not n57169 ; n57169_not
g97359 not n27595 ; n27595_not
g97360 not n31969 ; n31969_not
g97361 not n28549 ; n28549_not
g97362 not n31978 ; n31978_not
g97363 not n18559 ; n18559_not
g97364 not n16948 ; n16948_not
g97365 not n57178 ; n57178_not
g97366 not n29179 ; n29179_not
g97367 not n28486 ; n28486_not
g97368 not n57187 ; n57187_not
g97369 not a[10] ; a[10]_not
g97370 not n28288 ; n28288_not
g97371 not n57196 ; n57196_not
g97372 not n56809 ; n56809_not
g97373 not n25759 ; n25759_not
g97374 not n16984 ; n16984_not
g97375 not n27577 ; n27577_not
g97376 not n52687 ; n52687_not
g97377 not n17848 ; n17848_not
g97378 not n16939 ; n16939_not
g97379 not n50869 ; n50869_not
g97380 not n28567 ; n28567_not
g97381 not n18568 ; n18568_not
g97382 not n28558 ; n28558_not
g97383 not n31879 ; n31879_not
g97384 not n16966 ; n16966_not
g97385 not n26398 ; n26398_not
g97386 not n54658 ; n54658_not
g97387 not n50779 ; n50779_not
g97388 not n55666 ; n55666_not
g97389 not n56764 ; n56764_not
g97390 not n26389 ; n26389_not
g97391 not n19927 ; n19927_not
g97392 not n31897 ; n31897_not
g97393 not n57097 ; n57097_not
g97394 not n31888 ; n31888_not
g97395 not n29674 ; n29674_not
g97396 not n28945 ; n28945_not
g97397 not n18919 ; n18919_not
g97398 not n17497 ; n17497_not
g97399 not n14995 ; n14995_not
g97400 not n17569 ; n17569_not
g97401 not n18388 ; n18388_not
g97402 not n29683 ; n29683_not
g97403 not n52966 ; n52966_not
g97404 not n27694 ; n27694_not
g97405 not n15589 ; n15589_not
g97406 not n14977 ; n14977_not
g97407 not n27496 ; n27496_not
g97408 not n29692 ; n29692_not
g97409 not n54937 ; n54937_not
g97410 not n28864 ; n28864_not
g97411 not n25975 ; n25975_not
g97412 not n56098 ; n56098_not
g97413 not n52975 ; n52975_not
g97414 not n24778 ; n24778_not
g97415 not n18928 ; n18928_not
g97416 not n29593 ; n29593_not
g97417 not n25984 ; n25984_not
g97418 not n50599 ; n50599_not
g97419 not n55558 ; n55558_not
g97420 not n52984 ; n52984_not
g97421 not n29719 ; n29719_not
g97422 not n25993 ; n25993_not
g97423 not n18487 ; n18487_not
g97424 not n27955 ; n27955_not
g97425 not n29566 ; n29566_not
g97426 not n29557 ; n29557_not
g97427 not n29629 ; n29629_not
g97428 not n29548 ; n29548_not
g97429 not n27478 ; n27478_not
g97430 not n29539 ; n29539_not
g97431 not n52849 ; n52849_not
g97432 not n18883 ; n18883_not
g97433 not n52948 ; n52948_not
g97434 not n28873 ; n28873_not
g97435 not n29647 ; n29647_not
g97436 not n23797 ; n23797_not
g97437 not n18892 ; n18892_not
g97438 not n29656 ; n29656_not
g97439 not n11998 ; n11998_not
g97440 not n25966 ; n25966_not
g97441 not n29638 ; n29638_not
g97442 not n29278 ; n29278_not
g97443 not n29665 ; n29665_not
g97444 not n52957 ; n52957_not
g97445 not n54928 ; n54928_not
g97446 not n50968 ; n50968_not
g97447 not n54838 ; n54838_not
g97448 not n17479 ; n17479_not
g97449 not n15499 ; n15499_not
g97450 not n50986 ; n50986_not
g97451 not n29791 ; n29791_not
g97452 not n28846 ; n28846_not
g97453 not n18982 ; n18982_not
g97454 not n55783 ; n55783_not
g97455 not n29782 ; n29782_not
g97456 not n29359 ; n29359_not
g97457 not n11899 ; n11899_not
g97458 not n27748 ; n27748_not
g97459 not n29809 ; n29809_not
g97460 not n28189 ; n28189_not
g97461 not n18991 ; n18991_not
g97462 not n18469 ; n18469_not
g97463 not n50959 ; n50959_not
g97464 not n26299 ; n26299_not
g97465 not n52399 ; n52399_not
g97466 not n15598 ; n15598_not
g97467 not n18379 ; n18379_not
g97468 not n14986 ; n14986_not
g97469 not n18937 ; n18937_not
g97470 not n27928 ; n27928_not
g97471 not n18946 ; n18946_not
g97472 not n29746 ; n29746_not
g97473 not n55945 ; n55945_not
g97474 not n52498 ; n52498_not
g97475 not n18973 ; n18973_not
g97476 not n25678 ; n25678_not
g97477 not n28855 ; n28855_not
g97478 not n15679 ; n15679_not
g97479 not n27829 ; n27829_not
g97480 not n27289 ; n27289_not
g97481 not n18964 ; n18964_not
g97482 not n52993 ; n52993_not
g97483 not n25597 ; n25597_not
g97484 not n17488 ; n17488_not
g97485 not n29764 ; n29764_not
g97486 not n18955 ; n18955_not
g97487 not n54487 ; n54487_not
g97488 not n28936 ; n28936_not
g97489 not n12988 ; n12988_not
g97490 not n52885 ; n52885_not
g97491 not n18784 ; n18784_not
g97492 not n25876 ; n25876_not
g97493 not n23698 ; n23698_not
g97494 not n12979 ; n12979_not
g97495 not n52894 ; n52894_not
g97496 not n29395 ; n29395_not
g97497 not n17677 ; n17677_not
g97498 not n12898 ; n12898_not
g97499 not n18793 ; n18793_not
g97500 not n55477 ; n55477_not
g97501 not n25885 ; n25885_not
g97502 not n18478 ; n18478_not
g97503 not n27298 ; n27298_not
g97504 not n29494 ; n29494_not
g97505 not n24769 ; n24769_not
g97506 not n55963 ; n55963_not
g97507 not n25894 ; n25894_not
g97508 not n55468 ; n55468_not
g97509 not n27388 ; n27388_not
g97510 not n55990 ; n55990_not
g97511 not n29368 ; n29368_not
g97512 not n54856 ; n54856_not
g97513 not n28279 ; n28279_not
g97514 not n52867 ; n52867_not
g97515 not n14959 ; n14959_not
g97516 not n18775 ; n18775_not
g97517 not n54496 ; n54496_not
g97518 not n25867 ; n25867_not
g97519 not n55495 ; n55495_not
g97520 not n29449 ; n29449_not
g97521 not n29476 ; n29476_not
g97522 not n27856 ; n27856_not
g97523 not n29467 ; n29467_not
g97524 not n28099 ; n28099_not
g97525 not n55486 ; n55486_not
g97526 not n23689 ; n23689_not
g97527 not n52876 ; n52876_not
g97528 not n55972 ; n55972_not
g97529 not n12997 ; n12997_not
g97530 not n27658 ; n27658_not
g97531 not n25858 ; n25858_not
g97532 not n18766 ; n18766_not
g97533 not n25669 ; n25669_not
g97534 not n25939 ; n25939_not
g97535 not n25849 ; n25849_not
g97536 not n18865 ; n18865_not
g97537 not n52777 ; n52777_not
g97538 not n54847 ; n54847_not
g97539 not n25948 ; n25948_not
g97540 not n23779 ; n23779_not
g97541 not n18757 ; n18757_not
g97542 not n29575 ; n29575_not
g97543 not n54298 ; n54298_not
g97544 not n28891 ; n28891_not
g97545 not n28882 ; n28882_not
g97546 not n29584 ; n29584_not
g97547 not n18874 ; n18874_not
g97548 not n52939 ; n52939_not
g97549 not n25957 ; n25957_not
g97550 not n23788 ; n23788_not
g97551 not n50977 ; n50977_not
g97552 not n52588 ; n52588_not
g97553 not n27379 ; n27379_not
g97554 not n12889 ; n12889_not
g97555 not n52858 ; n52858_not
g97556 not n18829 ; n18829_not
g97557 not n18838 ; n18838_not
g97558 not n28918 ; n28918_not
g97559 not n28954 ; n28954_not
g97560 not n55549 ; n55549_not
g97561 not n55459 ; n55459_not
g97562 not n18847 ; n18847_not
g97563 not n52768 ; n52768_not
g97564 not n27973 ; n27973_not
g97565 not n28909 ; n28909_not
g97566 not n14968 ; n14968_not
g97567 not n27991 ; n27991_not
g97568 not n12799 ; n12799_not
g97569 not n18856 ; n18856_not
g97570 not n27397 ; n27397_not
g97571 not n27676 ; n27676_not
g97572 not n25687 ; n25687_not
g97573 not n29962 ; n29962_not
g97574 not n17389 ; n17389_not
g97575 not n27766 ; n27766_not
g97576 not n55576 ; n55576_not
g97577 not n54289 ; n54289_not
g97578 not n54397 ; n54397_not
g97579 not n28981 ; n28981_not
g97580 not n29980 ; n29980_not
g97581 not n28765 ; n28765_not
g97582 not n55747 ; n55747_not
g97583 not n29953 ; n29953_not
g97584 not n19198 ; n19198_not
g97585 not n15895 ; n15895_not
g97586 not n28369 ; n28369_not
g97587 not n28756 ; n28756_not
g97588 not n27784 ; n27784_not
g97589 not n53299 ; n53299_not
g97590 not n55918 ; n55918_not
g97591 not n55891 ; n55891_not
g97592 not n22969 ; n22969_not
g97593 not n24859 ; n24859_not
g97594 not n27757 ; n27757_not
g97595 not n22888 ; n22888_not
g97596 not n22897 ; n22897_not
g97597 not n17398 ; n17398_not
g97598 not n28783 ; n28783_not
g97599 not n29863 ; n29863_not
g97600 not n29935 ; n29935_not
g97601 not n29854 ; n29854_not
g97602 not n29845 ; n29845_not
g97603 not n28774 ; n28774_not
g97604 not n55369 ; n55369_not
g97605 not n27793 ; n27793_not
g97606 not n29836 ; n29836_not
g97607 not n15886 ; n15886_not
g97608 not n29827 ; n29827_not
g97609 not n54829 ; n54829_not
g97610 not n15958 ; n15958_not
g97611 not n17299 ; n17299_not
g97612 not n15787 ; n15787_not
g97613 not n24877 ; n24877_not
g97614 not n28378 ; n28378_not
g97615 not n28729 ; n28729_not
g97616 not n28387 ; n28387_not
g97617 not n15967 ; n15967_not
g97618 not n22879 ; n22879_not
g97619 not n55585 ; n55585_not
g97620 not n55846 ; n55846_not
g97621 not n54559 ; n54559_not
g97622 not n55729 ; n55729_not
g97623 not n22699 ; n22699_not
g97624 not n30889 ; n30889_not
g97625 not n29926 ; n29926_not
g97626 not n24868 ; n24868_not
g97627 not n24679 ; n24679_not
g97628 not n29917 ; n29917_not
g97629 not n22978 ; n22978_not
g97630 not n22987 ; n22987_not
g97631 not n15796 ; n15796_not
g97632 not n27775 ; n27775_not
g97633 not n28747 ; n28747_not
g97634 not n54955 ; n54955_not
g97635 not n25795 ; n25795_not
g97636 not n30799 ; n30799_not
g97637 not n18694 ; n18694_not
g97638 not n28738 ; n28738_not
g97639 not n22996 ; n22996_not
g97640 not n55738 ; n55738_not
g97641 not n15949 ; n15949_not
g97642 not n28828 ; n28828_not
g97643 not n54982 ; n54982_not
g97644 not n29755 ; n29755_not
g97645 not n55387 ; n55387_not
g97646 not n29872 ; n29872_not
g97647 not n29881 ; n29881_not
g97648 not n54379 ; n54379_not
g97649 not n23869 ; n23869_not
g97650 not n52759 ; n52759_not
g97651 not n24787 ; n24787_not
g97652 not n27883 ; n27883_not
g97653 not n15769 ; n15769_not
g97654 not n25489 ; n25489_not
g97655 not n18748 ; n18748_not
g97656 not n10999 ; n10999_not
g97657 not n18397 ; n18397_not
g97658 not n23878 ; n23878_not
g97659 not n28837 ; n28837_not
g97660 not n27865 ; n27865_not
g97661 not n55396 ; n55396_not
g97662 not n23887 ; n23887_not
g97663 not n55774 ; n55774_not
g97664 not n19288 ; n19288_not
g97665 not n17767 ; n17767_not
g97666 not n55378 ; n55378_not
g97667 not n55927 ; n55927_not
g97668 not n55756 ; n55756_not
g97669 not n28792 ; n28792_not
g97670 not n55936 ; n55936_not
g97671 not n15868 ; n15868_not
g97672 not n29890 ; n29890_not
g97673 not n18739 ; n18739_not
g97674 not n24796 ; n24796_not
g97675 not n54892 ; n54892_not
g97676 not n25579 ; n25579_not
g97677 not n15877 ; n15877_not
g97678 not n52696 ; n52696_not
g97679 not n55981 ; n55981_not
g97680 not n50896 ; n50896_not
g97681 not n17578 ; n17578_not
g97682 not n55765 ; n55765_not
g97683 not n25588 ; n25588_not
g97684 not n55567 ; n55567_not
g97685 not n28819 ; n28819_not
g97686 not n27838 ; n27838_not
g97687 not n35947 ; n35947_not
g97688 not n38692 ; n38692_not
g97689 not n48916 ; n48916_not
g97690 not n35938 ; n35938_not
g97691 not n35929 ; n35929_not
g97692 not n35893 ; n35893_not
g97693 not n37747 ; n37747_not
g97694 not n47647 ; n47647_not
g97695 not n34777 ; n34777_not
g97696 not n41968 ; n41968_not
g97697 not n35884 ; n35884_not
g97698 not n48907 ; n48907_not
g97699 not n37558 ; n37558_not
g97700 not n39385 ; n39385_not
g97701 not n39178 ; n39178_not
g97702 not n41977 ; n41977_not
g97703 not n35875 ; n35875_not
g97704 not n39790 ; n39790_not
g97705 not n47656 ; n47656_not
g97706 not n37765 ; n37765_not
g97707 not n48736 ; n48736_not
g97708 not n37549 ; n37549_not
g97709 not n48934 ; n48934_not
g97710 not n41878 ; n41878_not
g97711 not n47629 ; n47629_not
g97712 not n38683 ; n38683_not
g97713 not n35965 ; n35965_not
g97714 not n45829 ; n45829_not
g97715 not n41887 ; n41887_not
g97716 not n41896 ; n41896_not
g97717 not n34795 ; n34795_not
g97718 not n39772 ; n39772_not
g97719 not n35956 ; n35956_not
g97720 not n48925 ; n48925_not
g97721 not n37756 ; n37756_not
g97722 not n47638 ; n47638_not
g97723 not n39781 ; n39781_not
g97724 not n47674 ; n47674_not
g97725 not n48880 ; n48880_not
g97726 not n34768 ; n34768_not
g97727 not n49384 ; n49384_not
g97728 not n39808 ; n39808_not
g97729 not n35848 ; n35848_not
g97730 not n35839 ; n35839_not
g97731 not n45388 ; n45388_not
g97732 not n38746 ; n38746_not
g97733 not n41995 ; n41995_not
g97734 not n47683 ; n47683_not
g97735 not n48871 ; n48871_not
g97736 not n44389 ; n44389_not
g97737 not n38584 ; n38584_not
g97738 not n39817 ; n39817_not
g97739 not n49159 ; n49159_not
g97740 not n41599 ; n41599_not
g97741 not n38719 ; n38719_not
g97742 not n38728 ; n38728_not
g97743 not n37738 ; n37738_not
g97744 not n37567 ; n37567_not
g97745 not n41986 ; n41986_not
g97746 not n35866 ; n35866_not
g97747 not n47665 ; n47665_not
g97748 not n39682 ; n39682_not
g97749 not n45397 ; n45397_not
g97750 not n34759 ; n34759_not
g97751 not n38737 ; n38737_not
g97752 not n39376 ; n39376_not
g97753 not n49393 ; n49393_not
g97754 not n39673 ; n39673_not
g97755 not n35857 ; n35857_not
g97756 not n37729 ; n37729_not
g97757 not n38593 ; n38593_not
g97758 not n48763 ; n48763_not
g97759 not n45469 ; n45469_not
g97760 not n47566 ; n47566_not
g97761 not n38278 ; n38278_not
g97762 not n34885 ; n34885_not
g97763 not n44938 ; n44938_not
g97764 not n39718 ; n39718_not
g97765 not n38269 ; n38269_not
g97766 not n47575 ; n47575_not
g97767 not n38575 ; n38575_not
g97768 not n39736 ; n39736_not
g97769 not n44587 ; n44587_not
g97770 not n47584 ; n47584_not
g97771 not n38197 ; n38197_not
g97772 not n37792 ; n37792_not
g97773 not n43894 ; n43894_not
g97774 not n38188 ; n38188_not
g97775 not n38179 ; n38179_not
g97776 not n38629 ; n38629_not
g97777 not n38368 ; n38368_not
g97778 not n47539 ; n47539_not
g97779 not n37846 ; n37846_not
g97780 not n35992 ; n35992_not
g97781 not n38359 ; n38359_not
g97782 not n38539 ; n38539_not
g97783 not n42787 ; n42787_not
g97784 not n38557 ; n38557_not
g97785 not n37837 ; n37837_not
g97786 not n47548 ; n47548_not
g97787 not n42778 ; n42778_not
g97788 not n42769 ; n42769_not
g97789 not n37828 ; n37828_not
g97790 not n38296 ; n38296_not
g97791 not n42589 ; n42589_not
g97792 not n38287 ; n38287_not
g97793 not n34894 ; n34894_not
g97794 not n47557 ; n47557_not
g97795 not n37819 ; n37819_not
g97796 not n42679 ; n42679_not
g97797 not n49078 ; n49078_not
g97798 not n39754 ; n39754_not
g97799 not n37783 ; n37783_not
g97800 not n42598 ; n42598_not
g97801 not n35983 ; n35983_not
g97802 not n48952 ; n48952_not
g97803 not n34849 ; n34849_not
g97804 not n49087 ; n49087_not
g97805 not n39763 ; n39763_not
g97806 not n49096 ; n49096_not
g97807 not n48727 ; n48727_not
g97808 not n38674 ; n38674_not
g97809 not n48943 ; n48943_not
g97810 not n47188 ; n47188_not
g97811 not n39394 ; n39394_not
g97812 not n35974 ; n35974_not
g97813 not n37774 ; n37774_not
g97814 not n47593 ; n47593_not
g97815 not n38647 ; n38647_not
g97816 not n47197 ; n47197_not
g97817 not n48970 ; n48970_not
g97818 not n38656 ; n38656_not
g97819 not n38638 ; n38638_not
g97820 not n49438 ; n49438_not
g97821 not n42697 ; n42697_not
g97822 not n38665 ; n38665_not
g97823 not n34867 ; n34867_not
g97824 not n44929 ; n44929_not
g97825 not n49069 ; n49069_not
g97826 not n39709 ; n39709_not
g97827 not n48718 ; n48718_not
g97828 not n49429 ; n49429_not
g97829 not n39745 ; n39745_not
g97830 not n48961 ; n48961_not
g97831 not n42688 ; n42688_not
g97832 not n47764 ; n47764_not
g97833 not n38791 ; n38791_not
g97834 not n47773 ; n47773_not
g97835 not n37594 ; n37594_not
g97836 not n47098 ; n47098_not
g97837 not n48745 ; n48745_not
g97838 not n44857 ; n44857_not
g97839 not n49249 ; n49249_not
g97840 not n39295 ; n39295_not
g97841 not n48169 ; n48169_not
g97842 not n47782 ; n47782_not
g97843 not n48178 ; n48178_not
g97844 not n46495 ; n46495_not
g97845 not n34597 ; n34597_not
g97846 not n39862 ; n39862_not
g97847 not n49258 ; n49258_not
g97848 not n48088 ; n48088_not
g97849 not n37657 ; n37657_not
g97850 not n41698 ; n41698_not
g97851 not n48097 ; n48097_not
g97852 not n41689 ; n41689_not
g97853 not n39853 ; n39853_not
g97854 not n44875 ; n44875_not
g97855 not n43849 ; n43849_not
g97856 not n34669 ; n34669_not
g97857 not n43399 ; n43399_not
g97858 not n49348 ; n49348_not
g97859 not n47737 ; n47737_not
g97860 not n37648 ; n37648_not
g97861 not n47746 ; n47746_not
g97862 not n37639 ; n37639_not
g97863 not n48772 ; n48772_not
g97864 not n49339 ; n49339_not
g97865 not n47755 ; n47755_not
g97866 not n44866 ; n44866_not
g97867 not n49294 ; n49294_not
g97868 not n38818 ; n38818_not
g97869 not n34498 ; n34498_not
g97870 not n47809 ; n47809_not
g97871 not n38548 ; n38548_not
g97872 not n45298 ; n45298_not
g97873 not n43498 ; n43498_not
g97874 not n38827 ; n38827_not
g97875 not n33994 ; n33994_not
g97876 not n40897 ; n40897_not
g97877 not n38836 ; n38836_not
g97878 not n40969 ; n40969_not
g97879 not n40978 ; n40978_not
g97880 not n47818 ; n47818_not
g97881 not n48259 ; n48259_not
g97882 not n39277 ; n39277_not
g97883 not n47791 ; n47791_not
g97884 not n48187 ; n48187_not
g97885 not n34588 ; n34588_not
g97886 not n40879 ; n40879_not
g97887 not n48196 ; n48196_not
g97888 not n39286 ; n39286_not
g97889 not n49267 ; n49267_not
g97890 not n34579 ; n34579_not
g97891 not n38809 ; n38809_not
g97892 not n40888 ; n40888_not
g97893 not n43489 ; n43489_not
g97894 not n37576 ; n37576_not
g97895 not n49276 ; n49276_not
g97896 not n44848 ; n44848_not
g97897 not n34489 ; n34489_not
g97898 not n49285 ; n49285_not
g97899 not n49177 ; n49177_not
g97900 not n46468 ; n46468_not
g97901 not n39664 ; n39664_not
g97902 not n38773 ; n38773_not
g97903 not n39826 ; n39826_not
g97904 not n34399 ; n34399_not
g97905 not n49186 ; n49186_not
g97906 not n48844 ; n48844_not
g97907 not n41779 ; n41779_not
g97908 not n35776 ; n35776_not
g97909 not n37693 ; n37693_not
g97910 not n41788 ; n41788_not
g97911 not n49195 ; n49195_not
g97912 not n45865 ; n45865_not
g97913 not n43867 ; n43867_not
g97914 not n34696 ; n34696_not
g97915 not n45856 ; n45856_not
g97916 not n39367 ; n39367_not
g97917 not n48862 ; n48862_not
g97918 not n45379 ; n45379_not
g97919 not n38755 ; n38755_not
g97920 not n49168 ; n49168_not
g97921 not n35794 ; n35794_not
g97922 not n49375 ; n49375_not
g97923 not n39358 ; n39358_not
g97924 not n48781 ; n48781_not
g97925 not n38764 ; n38764_not
g97926 not n47692 ; n47692_not
g97927 not n48853 ; n48853_not
g97928 not n44893 ; n44893_not
g97929 not n35785 ; n35785_not
g97930 not n38782 ; n38782_not
g97931 not n34687 ; n34687_not
g97932 not n39844 ; n39844_not
g97933 not n36199 ; n36199_not
g97934 not n48808 ; n48808_not
g97935 not n43858 ; n43858_not
g97936 not n47728 ; n47728_not
g97937 not n46486 ; n46486_not
g97938 not n37666 ; n37666_not
g97939 not n48079 ; n48079_not
g97940 not n34678 ; n34678_not
g97941 not n46477 ; n46477_not
g97942 not n48790 ; n48790_not
g97943 not n37684 ; n37684_not
g97944 not n39349 ; n39349_not
g97945 not n39835 ; n39835_not
g97946 not n47719 ; n47719_not
g97947 not n39079 ; n39079_not
g97948 not n41797 ; n41797_not
g97949 not n44884 ; n44884_not
g97950 not n45874 ; n45874_not
g97951 not n39088 ; n39088_not
g97952 not n44398 ; n44398_not
g97953 not n37675 ; n37675_not
g97954 not n42859 ; n42859_not
g97955 not n43678 ; n43678_not
g97956 not n39457 ; n39457_not
g97957 not n42868 ; n42868_not
g97958 not n39475 ; n39475_not
g97959 not n42877 ; n42877_not
g97960 not n45586 ; n45586_not
g97961 not n39448 ; n39448_not
g97962 not n42886 ; n42886_not
g97963 not n39574 ; n39574_not
g97964 not n35695 ; n35695_not
g97965 not n39439 ; n39439_not
g97966 not n48556 ; n48556_not
g97967 not n34858 ; n34858_not
g97968 not n48835 ; n48835_not
g97969 not n43669 ; n43669_not
g97970 not n45595 ; n45595_not
g97971 not n38089 ; n38089_not
g97972 not n45658 ; n45658_not
g97973 not n37954 ; n37954_not
g97974 not n47296 ; n47296_not
g97975 not n39466 ; n39466_not
g97976 not n43687 ; n43687_not
g97977 not n49555 ; n49555_not
g97978 not n35668 ; n35668_not
g97979 not n35677 ; n35677_not
g97980 not n43759 ; n43759_not
g97981 not n37936 ; n37936_not
g97982 not n42985 ; n42985_not
g97983 not n37927 ; n37927_not
g97984 not n48592 ; n48592_not
g97985 not n34993 ; n34993_not
g97986 not n43768 ; n43768_not
g97987 not n37459 ; n37459_not
g97988 not n47449 ; n47449_not
g97989 not n42994 ; n42994_not
g97990 not n44992 ; n44992_not
g97991 not n47287 ; n47287_not
g97992 not n42895 ; n42895_not
g97993 not n45667 ; n45667_not
g97994 not n45577 ; n45577_not
g97995 not n43696 ; n43696_not
g97996 not n42949 ; n42949_not
g97997 not n42958 ; n42958_not
g97998 not n39583 ; n39583_not
g97999 not n42967 ; n42967_not
g98000 not n35758 ; n35758_not
g98001 not n35767 ; n35767_not
g98002 not n48583 ; n48583_not
g98003 not n45568 ; n45568_not
g98004 not n42976 ; n42976_not
g98005 not n47359 ; n47359_not
g98006 not n49492 ; n49492_not
g98007 not n38098 ; n38098_not
g98008 not n34939 ; n34939_not
g98009 not n47278 ; n47278_not
g98010 not n49357 ; n49357_not
g98011 not n39484 ; n39484_not
g98012 not n34948 ; n34948_not
g98013 not n47368 ; n47368_not
g98014 not n34957 ; n34957_not
g98015 not n49519 ; n49519_not
g98016 not n34966 ; n34966_not
g98017 not n34975 ; n34975_not
g98018 not n49447 ; n49447_not
g98019 not n39538 ; n39538_not
g98020 not n49465 ; n49465_not
g98021 not n49474 ; n49474_not
g98022 not n43579 ; n43579_not
g98023 not n39493 ; n39493_not
g98024 not n43588 ; n43588_not
g98025 not n45739 ; n45739_not
g98026 not n47395 ; n47395_not
g98027 not n37963 ; n37963_not
g98028 not n42796 ; n42796_not
g98029 not n48547 ; n48547_not
g98030 not n49564 ; n49564_not
g98031 not n43597 ; n43597_not
g98032 not n34984 ; n34984_not
g98033 not n37990 ; n37990_not
g98034 not n47377 ; n47377_not
g98035 not n37981 ; n37981_not
g98036 not n49537 ; n49537_not
g98037 not n45649 ; n45649_not
g98038 not n39556 ; n39556_not
g98039 not n47386 ; n47386_not
g98040 not n44965 ; n44965_not
g98041 not n38458 ; n38458_not
g98042 not n46378 ; n46378_not
g98043 not n45784 ; n45784_not
g98044 not n38467 ; n38467_not
g98045 not n39268 ; n39268_not
g98046 not n39259 ; n39259_not
g98047 not n48673 ; n48673_not
g98048 not n37873 ; n37873_not
g98049 not n39691 ; n39691_not
g98050 not n46369 ; n46369_not
g98051 not n44974 ; n44974_not
g98052 not n45775 ; n45775_not
g98053 not n47494 ; n47494_not
g98054 not n37882 ; n37882_not
g98055 not n38449 ; n38449_not
g98056 not n45487 ; n45487_not
g98057 not n39187 ; n39187_not
g98058 not n46387 ; n46387_not
g98059 not n37864 ; n37864_not
g98060 not n38395 ; n38395_not
g98061 not n38386 ; n38386_not
g98062 not n45478 ; n45478_not
g98063 not n44947 ; n44947_not
g98064 not n37855 ; n37855_not
g98065 not n38377 ; n38377_not
g98066 not n46396 ; n46396_not
g98067 not n43876 ; n43876_not
g98068 not n48682 ; n48682_not
g98069 not n45496 ; n45496_not
g98070 not n44956 ; n44956_not
g98071 not n48691 ; n48691_not
g98072 not n38485 ; n38485_not
g98073 not n38494 ; n38494_not
g98074 not n49483 ; n49483_not
g98075 not n45199 ; n45199_not
g98076 not n39628 ; n39628_not
g98077 not n43786 ; n43786_not
g98078 not n45766 ; n45766_not
g98079 not n37468 ; n37468_not
g98080 not n45685 ; n45685_not
g98081 not n47467 ; n47467_not
g98082 not n45559 ; n45559_not
g98083 not n37918 ; n37918_not
g98084 not n47458 ; n47458_not
g98085 not n37909 ; n37909_not
g98086 not n49528 ; n49528_not
g98087 not n45694 ; n45694_not
g98088 not n39619 ; n39619_not
g98089 not n37891 ; n37891_not
g98090 not n47089 ; n47089_not
g98091 not n35686 ; n35686_not
g98092 not n42499 ; n42499_not
g98093 not n47485 ; n47485_not
g98094 not n39646 ; n39646_not
g98095 not n44983 ; n44983_not
g98096 not n48628 ; n48628_not
g98097 not n37477 ; n37477_not
g98098 not n47476 ; n47476_not
g98099 not n48637 ; n48637_not
g98100 not n48646 ; n48646_not
g98101 not n48286 ; n48286_not
g98102 not n48277 ; n48277_not
g98103 not n32986 ; n32986_not
g98104 not n44794 ; n44794_not
g98105 not n38935 ; n38935_not
g98106 not n36676 ; n36676_not
g98107 not n47944 ; n47944_not
g98108 not n48268 ; n48268_not
g98109 not n36649 ; n36649_not
g98110 not n32968 ; n32968_not
g98111 not n44659 ; n44659_not
g98112 not n32959 ; n32959_not
g98113 not n40699 ; n40699_not
g98114 not n40789 ; n40789_not
g98115 not n39916 ; n39916_not
g98116 not n38926 ; n38926_not
g98117 not n45793 ; n45793_not
g98118 not n46567 ; n46567_not
g98119 not n33985 ; n33985_not
g98120 not n47908 ; n47908_not
g98121 not n47827 ; n47827_not
g98122 not n38962 ; n38962_not
g98123 not n38953 ; n38953_not
g98124 not n48493 ; n48493_not
g98125 not n44497 ; n44497_not
g98126 not n38944 ; n38944_not
g98127 not n46558 ; n46558_not
g98128 not n48295 ; n48295_not
g98129 not n32887 ; n32887_not
g98130 not n48484 ; n48484_not
g98131 not n39907 ; n39907_not
g98132 not n36667 ; n36667_not
g98133 not n48475 ; n48475_not
g98134 not n44668 ; n44668_not
g98135 not n37486 ; n37486_not
g98136 not n32599 ; n32599_not
g98137 not n48466 ; n48466_not
g98138 not n32878 ; n32878_not
g98139 not n32869 ; n32869_not
g98140 not n44677 ; n44677_not
g98141 not n48457 ; n48457_not
g98142 not n46639 ; n46639_not
g98143 not n36658 ; n36658_not
g98144 not n38917 ; n38917_not
g98145 not n45289 ; n45289_not
g98146 not n46648 ; n46648_not
g98147 not n38908 ; n38908_not
g98148 not n47953 ; n47953_not
g98149 not n47881 ; n47881_not
g98150 not n32896 ; n32896_not
g98151 not n47962 ; n47962_not
g98152 not n48565 ; n48565_not
g98153 not n47971 ; n47971_not
g98154 not n33697 ; n33697_not
g98155 not n45838 ; n45838_not
g98156 not n33499 ; n33499_not
g98157 not n36991 ; n36991_not
g98158 not n33679 ; n33679_not
g98159 not n39952 ; n39952_not
g98160 not n48448 ; n48448_not
g98161 not n48376 ; n48376_not
g98162 not n36577 ; n36577_not
g98163 not n44767 ; n44767_not
g98164 not n39934 ; n39934_not
g98165 not n44596 ; n44596_not
g98166 not n39169 ; n39169_not
g98167 not n33589 ; n33589_not
g98168 not n44749 ; n44749_not
g98169 not n44569 ; n44569_not
g98170 not n47872 ; n47872_not
g98171 not n47863 ; n47863_not
g98172 not n44758 ; n44758_not
g98173 not n48394 ; n48394_not
g98174 not n44479 ; n44479_not
g98175 not n39943 ; n39943_not
g98176 not n33769 ; n33769_not
g98177 not n47854 ; n47854_not
g98178 not n46585 ; n46585_not
g98179 not n48439 ; n48439_not
g98180 not n48385 ; n48385_not
g98181 not n48349 ; n48349_not
g98182 not n44488 ; n44488_not
g98183 not n46576 ; n46576_not
g98184 not n37099 ; n37099_not
g98185 not n36559 ; n36559_not
g98186 not n44785 ; n44785_not
g98187 not n39925 ; n39925_not
g98188 not n45883 ; n45883_not
g98189 not n39970 ; n39970_not
g98190 not n47917 ; n47917_not
g98191 not n32977 ; n32977_not
g98192 not n33598 ; n33598_not
g98193 not n45676 ; n45676_not
g98194 not n44776 ; n44776_not
g98195 not n48367 ; n48367_not
g98196 not n39592 ; n39592_not
g98197 not n36568 ; n36568_not
g98198 not n48358 ; n48358_not
g98199 not n39961 ; n39961_not
g98200 not n47926 ; n47926_not
g98201 not n32788 ; n32788_not
g98202 not n45919 ; n45919_not
g98203 not n44839 ; n44839_not
g98204 not n43777 ; n43777_not
g98205 not n38881 ; n38881_not
g98206 not n36586 ; n36586_not
g98207 not n32779 ; n32779_not
g98208 not n32689 ; n32689_not
g98209 not n40996 ; n40996_not
g98210 not n32797 ; n32797_not
g98211 not n38863 ; n38863_not
g98212 not n45748 ; n45748_not
g98213 not n45928 ; n45928_not
g98214 not n38872 ; n38872_not
g98215 not n39097 ; n39097_not
g98216 not n48655 ; n48655_not
g98217 not n39880 ; n39880_not
g98218 not n44686 ; n44686_not
g98219 not n44695 ; n44695_not
g98220 not n39637 ; n39637_not
g98221 not n47836 ; n47836_not
g98222 not n39871 ; n39871_not
g98223 not n32698 ; n32698_not
g98224 not n40987 ; n40987_not
g98225 not n39547 ; n39547_not
g98226 not n38890 ; n38890_not
g98227 not n36973 ; n36973_not
g98228 not n38845 ; n38845_not
g98229 not n38854 ; n38854_not
g98230 not n17885 ; n17885_not
g98231 not n35768 ; n35768_not
g98232 not b[10] ; b[10]_not
g98233 not n15977 ; n15977_not
g98234 not n24689 ; n24689_not
g98235 not n51797 ; n51797_not
g98236 not n25688 ; n25688_not
g98237 not n25796 ; n25796_not
g98238 not n39548 ; n39548_not
g98239 not n37298 ; n37298_not
g98240 not n45668 ; n45668_not
g98241 not n47873 ; n47873_not
g98242 not n49097 ; n49097_not
g98243 not n39953 ; n39953_not
g98244 not n35867 ; n35867_not
g98245 not n45677 ; n45677_not
g98246 not n27893 ; n27893_not
g98247 not n24779 ; n24779_not
g98248 not n39638 ; n39638_not
g98249 not n25697 ; n25697_not
g98250 not n35858 ; n35858_not
g98251 not n37487 ; n37487_not
g98252 not n37469 ; n37469_not
g98253 not n37289 ; n37289_not
g98254 not n34985 ; n34985_not
g98255 not n27776 ; n27776_not
g98256 not n39962 ; n39962_not
g98257 not n27938 ; n27938_not
g98258 not n14699 ; n14699_not
g98259 not n49394 ; n49394_not
g98260 not n15959 ; n15959_not
g98261 not n45569 ; n45569_not
g98262 not n55496 ; n55496_not
g98263 not n34976 ; n34976_not
g98264 not n36866 ; n36866_not
g98265 not n34967 ; n34967_not
g98266 not n54785 ; n54785_not
g98267 not n51599 ; n51599_not
g98268 not n45848 ; n45848_not
g98269 not n34994 ; n34994_not
g98270 not n16958 ; n16958_not
g98271 not n35849 ; n35849_not
g98272 not n28478 ; n28478_not
g98273 not n51788 ; n51788_not
g98274 not n15968 ; n15968_not
g98275 not n54866 ; n54866_not
g98276 not n24788 ; n24788_not
g98277 not n39629 ; n39629_not
g98278 not n25679 ; n25679_not
g98279 not n36569 ; n36569_not
g98280 not n36857 ; n36857_not
g98281 not n15599 ; n15599_not
g98282 not n52967 ; n52967_not
g98283 not n45758 ; n45758_not
g98284 not n47882 ; n47882_not
g98285 not n48656 ; n48656_not
g98286 not n36839 ; n36839_not
g98287 not n35894 ; n35894_not
g98288 not n52769 ; n52769_not
g98289 not n17894 ; n17894_not
g98290 not n15986 ; n15986_not
g98291 not n45776 ; n45776_not
g98292 not n25778 ; n25778_not
g98293 not n49079 ; n49079_not
g98294 not n34778 ; n34778_not
g98295 not n21989 ; n21989_not
g98296 not n55298 ; n55298_not
g98297 not n39593 ; n39593_not
g98298 not n54884 ; n54884_not
g98299 not n15689 ; n15689_not
g98300 not n15995 ; n15995_not
g98301 not n25769 ; n25769_not
g98302 not n48647 ; n48647_not
g98303 not n54776 ; n54776_not
g98304 not n39539 ; n39539_not
g98305 not n49439 ; n49439_not
g98306 not n37892 ; n37892_not
g98307 not n45389 ; n45389_not
g98308 not n21998 ; n21998_not
g98309 not n28496 ; n28496_not
g98310 not n55289 ; n55289_not
g98311 not n35687 ; n35687_not
g98312 not n37379 ; n37379_not
g98313 not n52949 ; n52949_not
g98314 not n54893 ; n54893_not
g98315 not n39656 ; n39656_not
g98316 not n35876 ; n35876_not
g98317 not n46199 ; n46199_not
g98318 not n27785 ; n27785_not
g98319 not n52958 ; n52958_not
g98320 not n27866 ; n27866_not
g98321 not n37883 ; n37883_not
g98322 not n27875 ; n27875_not
g98323 not n49088 ; n49088_not
g98324 not n16967 ; n16967_not
g98325 not n21899 ; n21899_not
g98326 not n54875 ; n54875_not
g98327 not n45659 ; n45659_not
g98328 not n37478 ; n37478_not
g98329 not n36578 ; n36578_not
g98330 not n35678 ; n35678_not
g98331 not n27848 ; n27848_not
g98332 not n35696 ; n35696_not
g98333 not n48638 ; n48638_not
g98334 not n35885 ; n35885_not
g98335 not n52778 ; n52778_not
g98336 not n36848 ; n36848_not
g98337 not n25787 ; n25787_not
g98338 not n45398 ; n45398_not
g98339 not n37388 ; n37388_not
g98340 not n34769 ; n34769_not
g98341 not n52688 ; n52688_not
g98342 not n39566 ; n39566_not
g98343 not n45479 ; n45479_not
g98344 not n35579 ; n35579_not
g98345 not n24986 ; n24986_not
g98346 not n35588 ; n35588_not
g98347 not n56189 ; n56189_not
g98348 not n35399 ; n35399_not
g98349 not n36983 ; n36983_not
g98350 not n48557 ; n48557_not
g98351 not n37955 ; n37955_not
g98352 not n35597 ; n35597_not
g98353 not n49259 ; n49259_not
g98354 not n47297 ; n47297_not
g98355 not n14978 ; n14978_not
g98356 not n36947 ; n36947_not
g98357 not n55379 ; n55379_not
g98358 not n47954 ; n47954_not
g98359 not n27929 ; n27929_not
g98360 not n14969 ; n14969_not
g98361 not n34958 ; n34958_not
g98362 not n15869 ; n15869_not
g98363 not n15779 ; n15779_not
g98364 not n36929 ; n36929_not
g98365 not n17795 ; n17795_not
g98366 not n35489 ; n35489_not
g98367 not n27794 ; n27794_not
g98368 not n27965 ; n27965_not
g98369 not n49349 ; n49349_not
g98370 not n35498 ; n35498_not
g98371 not n54794 ; n54794_not
g98372 not n36938 ; n36938_not
g98373 not n28199 ; n28199_not
g98374 not n52697 ; n52697_not
g98375 not n51698 ; n51698_not
g98376 not n48566 ; n48566_not
g98377 not n45587 ; n45587_not
g98378 not n27956 ; n27956_not
g98379 not n14879 ; n14879_not
g98380 not n37946 ; n37946_not
g98381 not n24959 ; n24959_not
g98382 not n36965 ; n36965_not
g98383 not n14897 ; n14897_not
g98384 not n47972 ; n47972_not
g98385 not n37973 ; n37973_not
g98386 not n55388 ; n55388_not
g98387 not n49286 ; n49286_not
g98388 not n24968 ; n24968_not
g98389 not n48539 ; n48539_not
g98390 not n47963 ; n47963_not
g98391 not n49295 ; n49295_not
g98392 not n36974 ; n36974_not
g98393 not n17867 ; n17867_not
g98394 not n17876 ; n17876_not
g98395 not n45488 ; n45488_not
g98396 not n36956 ; n36956_not
g98397 not n45785 ; n45785_not
g98398 not n14888 ; n14888_not
g98399 not n49268 ; n49268_not
g98400 not n48548 ; n48548_not
g98401 not n49277 ; n49277_not
g98402 not n45596 ; n45596_not
g98403 not n45497 ; n45497_not
g98404 not n28298 ; n28298_not
g98405 not n27839 ; n27839_not
g98406 not n15797 ; n15797_not
g98407 not n24977 ; n24977_not
g98408 not n17849 ; n17849_not
g98409 not n25598 ; n25598_not
g98410 not n52976 ; n52976_not
g98411 not n49169 ; n49169_not
g98412 not n39971 ; n39971_not
g98413 not n45578 ; n45578_not
g98414 not n27983 ; n27983_not
g98415 not n34949 ; n34949_not
g98416 not n36884 ; n36884_not
g98417 not n49178 ; n49178_not
g98418 not n17687 ; n17687_not
g98419 not n37928 ; n37928_not
g98420 not n48593 ; n48593_not
g98421 not n54848 ; n54848_not
g98422 not n55478 ; n55478_not
g98423 not n25589 ; n25589_not
g98424 not n24797 ; n24797_not
g98425 not n55487 ; n55487_not
g98426 not n37919 ; n37919_not
g98427 not n54857 ; n54857_not
g98428 not n35795 ; n35795_not
g98429 not n49385 ; n49385_not
g98430 not n36875 ; n36875_not
g98431 not n17669 ; n17669_not
g98432 not n39584 ; n39584_not
g98433 not n14987 ; n14987_not
g98434 not n47909 ; n47909_not
g98435 not n56198 ; n56198_not
g98436 not n45686 ; n45686_not
g98437 not n35786 ; n35786_not
g98438 not n49196 ; n49196_not
g98439 not n55469 ; n55469_not
g98440 not n47927 ; n47927_not
g98441 not n15887 ; n15887_not
g98442 not n24878 ; n24878_not
g98443 not n17759 ; n17759_not
g98444 not n14798 ; n14798_not
g98445 not n28388 ; n28388_not
g98446 not n47288 ; n47288_not
g98447 not n24599 ; n24599_not
g98448 not n52598 ; n52598_not
g98449 not n52994 ; n52994_not
g98450 not n17777 ; n17777_not
g98451 not n45749 ; n45749_not
g98452 not n24887 ; n24887_not
g98453 not n55397 ; n55397_not
g98454 not n15878 ; n15878_not
g98455 not n24896 ; n24896_not
g98456 not n49187 ; n49187_not
g98457 not n49367 ; n49367_not
g98458 not n45695 ; n45695_not
g98459 not n52985 ; n52985_not
g98460 not n37937 ; n37937_not
g98461 not n15896 ; n15896_not
g98462 not n36893 ; n36893_not
g98463 not n35777 ; n35777_not
g98464 not n37991 ; n37991_not
g98465 not n39980 ; n39980_not
g98466 not n24995 ; n24995_not
g98467 not n47918 ; n47918_not
g98468 not n54839 ; n54839_not
g98469 not n25499 ; n25499_not
g98470 not n37199 ; n37199_not
g98471 not n24869 ; n24869_not
g98472 not n39557 ; n39557_not
g98473 not n14789 ; n14789_not
g98474 not n23888 ; n23888_not
g98475 not n47864 ; n47864_not
g98476 not n26984 ; n26984_not
g98477 not n37685 ; n37685_not
g98478 not n23879 ; n23879_not
g98479 not n45866 ; n45866_not
g98480 not n55775 ; n55775_not
g98481 not n48791 ; n48791_not
g98482 not n55766 ; n55766_not
g98483 not n39890 ; n39890_not
g98484 not n37694 ; n37694_not
g98485 not n55667 ; n55667_not
g98486 not n39827 ; n39827_not
g98487 not n23798 ; n23798_not
g98488 not n55757 ; n55757_not
g98489 not n23789 ; n23789_not
g98490 not n48782 ; n48782_not
g98491 not n48575 ; n48575_not
g98492 not n13997 ; n13997_not
g98493 not n52877 ; n52877_not
g98494 not n55748 ; n55748_not
g98495 not n55658 ; n55658_not
g98496 not n39845 ; n39845_not
g98497 not n48809 ; n48809_not
g98498 not n45929 ; n45929_not
g98499 not n36596 ; n36596_not
g98500 not n41789 ; n41789_not
g98501 not n48818 ; n48818_not
g98502 not n54389 ; n54389_not
g98503 not n37676 ; n37676_not
g98504 not n55676 ; n55676_not
g98505 not n26957 ; n26957_not
g98506 not n23699 ; n23699_not
g98507 not n40988 ; n40988_not
g98508 not n41798 ; n41798_not
g98509 not n26966 ; n26966_not
g98510 not n36659 ; n36659_not
g98511 not n39836 ; n39836_not
g98512 not n48827 ; n48827_not
g98513 not n40979 ; n40979_not
g98514 not n23897 ; n23897_not
g98515 not n36668 ; n36668_not
g98516 not n52886 ; n52886_not
g98517 not n13889 ; n13889_not
g98518 not n36695 ; n36695_not
g98519 not n16499 ; n16499_not
g98520 not n40799 ; n40799_not
g98521 not n41996 ; n41996_not
g98522 not n41987 ; n41987_not
g98523 not n55847 ; n55847_not
g98524 not n55694 ; n55694_not
g98525 not n52859 ; n52859_not
g98526 not n39917 ; n39917_not
g98527 not n55685 ; n55685_not
g98528 not n39791 ; n39791_not
g98529 not n37739 ; n37739_not
g98530 not n45893 ; n45893_not
g98531 not n36749 ; n36749_not
g98532 not n41978 ; n41978_not
g98533 not n36758 ; n36758_not
g98534 not n55865 ; n55865_not
g98535 not n39908 ; n39908_not
g98536 not n39818 ; n39818_not
g98537 not n13988 ; n13988_not
g98538 not n41888 ; n41888_not
g98539 not n41897 ; n41897_not
g98540 not n40898 ; n40898_not
g98541 not n55739 ; n55739_not
g98542 not n48773 ; n48773_not
g98543 not n13979 ; n13979_not
g98544 not n52868 ; n52868_not
g98545 not n36686 ; n36686_not
g98546 not n55649 ; n55649_not
g98547 not n40889 ; n40889_not
g98548 not n37577 ; n37577_not
g98549 not n39809 ; n39809_not
g98550 not n55838 ; n55838_not
g98551 not n47891 ; n47891_not
g98552 not n37568 ; n37568_not
g98553 not n39674 ; n39674_not
g98554 not n37586 ; n37586_not
g98555 not n48728 ; n48728_not
g98556 not n35939 ; n35939_not
g98557 not n39863 ; n39863_not
g98558 not n55199 ; n55199_not
g98559 not n48737 ; n48737_not
g98560 not n36389 ; n36389_not
g98561 not n39872 ; n39872_not
g98562 not n45974 ; n45974_not
g98563 not n39647 ; n39647_not
g98564 not n47846 ; n47846_not
g98565 not n48665 ; n48665_not
g98566 not n54974 ; n54974_not
g98567 not n45983 ; n45983_not
g98568 not n36497 ; n36497_not
g98569 not n54965 ; n54965_not
g98570 not n48692 ; n48692_not
g98571 not n45956 ; n45956_not
g98572 not n47819 ; n47819_not
g98573 not n36488 ; n36488_not
g98574 not n47828 ; n47828_not
g98575 not n36479 ; n36479_not
g98576 not n35993 ; n35993_not
g98577 not n48683 ; n48683_not
g98578 not n37559 ; n37559_not
g98579 not n35984 ; n35984_not
g98580 not n35975 ; n35975_not
g98581 not n45965 ; n45965_not
g98582 not n35966 ; n35966_not
g98583 not n35957 ; n35957_not
g98584 not n35948 ; n35948_not
g98585 not n36398 ; n36398_not
g98586 not n45884 ; n45884_not
g98587 not n36299 ; n36299_not
g98588 not n23969 ; n23969_not
g98589 not n37649 ; n37649_not
g98590 not n39854 ; n39854_not
g98591 not n54938 ; n54938_not
g98592 not n45938 ; n45938_not
g98593 not n39881 ; n39881_not
g98594 not n54983 ; n54983_not
g98595 not n54929 ; n54929_not
g98596 not n37658 ; n37658_not
g98597 not n41699 ; n41699_not
g98598 not n16994 ; n16994_not
g98599 not n52895 ; n52895_not
g98600 not n26939 ; n26939_not
g98601 not n40997 ; n40997_not
g98602 not n45875 ; n45875_not
g98603 not n37667 ; n37667_not
g98604 not n23996 ; n23996_not
g98605 not n48755 ; n48755_not
g98606 not n16949 ; n16949_not
g98607 not n23987 ; n23987_not
g98608 not n45992 ; n45992_not
g98609 not n23978 ; n23978_not
g98610 not n45947 ; n45947_not
g98611 not n16976 ; n16976_not
g98612 not n37496 ; n37496_not
g98613 not n37838 ; n37838_not
g98614 not n25949 ; n25949_not
g98615 not n37847 ; n37847_not
g98616 not n55586 ; n55586_not
g98617 not n39728 ; n39728_not
g98618 not n36794 ; n36794_not
g98619 not n54947 ; n54947_not
g98620 not n26975 ; n26975_not
g98621 not n39188 ; n39188_not
g98622 not n37856 ; n37856_not
g98623 not n39719 ; n39719_not
g98624 not n39197 ; n39197_not
g98625 not n55982 ; n55982_not
g98626 not n25976 ; n25976_not
g98627 not n47936 ; n47936_not
g98628 not n47837 ; n47837_not
g98629 not n51959 ; n51959_not
g98630 not n51887 ; n51887_not
g98631 not n12899 ; n12899_not
g98632 not n25967 ; n25967_not
g98633 not n12989 ; n12989_not
g98634 not n12998 ; n12998_not
g98635 not n22799 ; n22799_not
g98636 not n51896 ; n51896_not
g98637 not n36785 ; n36785_not
g98638 not n37829 ; n37829_not
g98639 not n25958 ; n25958_not
g98640 not n25859 ; n25859_not
g98641 not n52796 ; n52796_not
g98642 not n39683 ; n39683_not
g98643 not n37874 ; n37874_not
g98644 not n55559 ; n55559_not
g98645 not n51878 ; n51878_not
g98646 not n39944 ; n39944_not
g98647 not n36587 ; n36587_not
g98648 not n52787 ; n52787_not
g98649 not n39935 ; n39935_not
g98650 not n25895 ; n25895_not
g98651 not n25886 ; n25886_not
g98652 not n55577 ; n55577_not
g98653 not n37865 ; n37865_not
g98654 not n37397 ; n37397_not
g98655 not n25877 ; n25877_not
g98656 not n47981 ; n47981_not
g98657 not n25868 ; n25868_not
g98658 not n55568 ; n55568_not
g98659 not n45794 ; n45794_not
g98660 not n55892 ; n55892_not
g98661 not n36767 ; n36767_not
g98662 not a[20] ; a[20]_not
g98663 not n37766 ; n37766_not
g98664 not n55595 ; n55595_not
g98665 not n22979 ; n22979_not
g98666 not n39764 ; n39764_not
g98667 not n37775 ; n37775_not
g98668 not n22988 ; n22988_not
g98669 not n45299 ; n45299_not
g98670 not n45839 ; n45839_not
g98671 not n22889 ; n22889_not
g98672 not n37748 ; n37748_not
g98673 not n13799 ; n13799_not
g98674 not n48746 ; n48746_not
g98675 not n22898 ; n22898_not
g98676 not n39782 ; n39782_not
g98677 not n39692 ; n39692_not
g98678 not n55883 ; n55883_not
g98679 not n39773 ; n39773_not
g98680 not n37757 ; n37757_not
g98681 not n47198 ; n47198_not
g98682 not n51986 ; n51986_not
g98683 not n25994 ; n25994_not
g98684 not n39737 ; n39737_not
g98685 not n37793 ; n37793_not
g98686 not n25985 ; n25985_not
g98687 not n51977 ; n51977_not
g98688 not n36776 ; n36776_not
g98689 not n51968 ; n51968_not
g98690 not n55973 ; n55973_not
g98691 not n42599 ; n42599_not
g98692 not n22997 ; n22997_not
g98693 not n39755 ; n39755_not
g98694 not n54992 ; n54992_not
g98695 not n55928 ; n55928_not
g98696 not n55937 ; n55937_not
g98697 not n39746 ; n39746_not
g98698 not n39926 ; n39926_not
g98699 not n44597 ; n44597_not
g98700 not n37784 ; n37784_not
g98701 not n51995 ; n51995_not
g98702 not n55955 ; n55955_not
g98703 not n46694 ; n46694_not
g98704 not n29459 ; n29459_not
g98705 not n34598 ; n34598_not
g98706 not n49808 ; n49808_not
g98707 not n29468 ; n29468_not
g98708 not n34859 ; n34859_not
g98709 not n56684 ; n56684_not
g98710 not n38549 ; n38549_not
g98711 not n56666 ; n56666_not
g98712 not n43976 ; n43976_not
g98713 not n46991 ; n46991_not
g98714 not n53579 ; n53579_not
g98715 not n49817 ; n49817_not
g98716 not n43499 ; n43499_not
g98717 not n18776 ; n18776_not
g98718 not n29486 ; n29486_not
g98719 not n43949 ; n43949_not
g98720 not n19379 ; n19379_not
g98721 not n43688 ; n43688_not
g98722 not n39179 ; n39179_not
g98723 not n49790 ; n49790_not
g98724 not n34877 ; n34877_not
g98725 not n53975 ; n53975_not
g98726 not n38639 ; n38639_not
g98727 not n19919 ; n19919_not
g98728 not n29738 ; n29738_not
g98729 not n56846 ; n56846_not
g98730 not n50888 ; n50888_not
g98731 not n53984 ; n53984_not
g98732 not n53588 ; n53588_not
g98733 not n56396 ; n56396_not
g98734 not n53993 ; n53993_not
g98735 not n19577 ; n19577_not
g98736 not n54596 ; n54596_not
g98737 not n44849 ; n44849_not
g98738 not n34589 ; n34589_not
g98739 not n19892 ; n19892_not
g98740 not n46397 ; n46397_not
g98741 not n44759 ; n44759_not
g98742 not n43967 ; n43967_not
g98743 not n43958 ; n43958_not
g98744 not n49844 ; n49844_not
g98745 not n46775 ; n46775_not
g98746 not n56648 ; n56648_not
g98747 not n38495 ; n38495_not
g98748 not n46586 ; n46586_not
g98749 not n38990 ; n38990_not
g98750 not n46973 ; n46973_not
g98751 not n30989 ; n30989_not
g98752 not n56855 ; n56855_not
g98753 not n29549 ; n29549_not
g98754 not n54578 ; n54578_not
g98755 not n56459 ; n56459_not
g98756 not n49853 ; n49853_not
g98757 not n38189 ; n38189_not
g98758 not n29558 ; n29558_not
g98759 not n19847 ; n19847_not
g98760 not n33869 ; n33869_not
g98761 not n46964 ; n46964_not
g98762 not n56639 ; n56639_not
g98763 not n18758 ; n18758_not
g98764 not n34787 ; n34787_not
g98765 not n46577 ; n46577_not
g98766 not n56675 ; n56675_not
g98767 not n49826 ; n49826_not
g98768 not n46847 ; n46847_not
g98769 not n29909 ; n29909_not
g98770 not n54587 ; n54587_not
g98771 not n19874 ; n19874_not
g98772 not n18767 ; n18767_not
g98773 not n34679 ; n34679_not
g98774 not n19586 ; n19586_not
g98775 not n49835 ; n49835_not
g98776 not n29747 ; n29747_not
g98777 not n56657 ; n56657_not
g98778 not n34688 ; n34688_not
g98779 not n46982 ; n46982_not
g98780 not n56693 ; n56693_not
g98781 not n19865 ; n19865_not
g98782 not n34697 ; n34697_not
g98783 not n17678 ; n17678_not
g98784 not n56819 ; n56819_not
g98785 not n43985 ; n43985_not
g98786 not n29927 ; n29927_not
g98787 not n46388 ; n46388_not
g98788 not n29198 ; n29198_not
g98789 not n19982 ; n19982_not
g98790 not n18686 ; n18686_not
g98791 not n49475 ; n49475_not
g98792 not n19559 ; n19559_not
g98793 not n18794 ; n18794_not
g98794 not n49727 ; n49727_not
g98795 not n46595 ; n46595_not
g98796 not n44948 ; n44948_not
g98797 not n46838 ; n46838_not
g98798 not n34895 ; n34895_not
g98799 not n29918 ; n29918_not
g98800 not n49736 ; n49736_not
g98801 not n19388 ; n19388_not
g98802 not n53939 ; n53939_not
g98803 not n33689 ; n33689_not
g98804 not n49745 ; n49745_not
g98805 not n53669 ; n53669_not
g98806 not n46676 ; n46676_not
g98807 not n19568 ; n19568_not
g98808 not n49754 ; n49754_not
g98809 not n29279 ; n29279_not
g98810 not n56891 ; n56891_not
g98811 not n56594 ; n56594_not
g98812 not n38459 ; n38459_not
g98813 not n48971 ; n48971_not
g98814 not n38477 ; n38477_not
g98815 not n49493 ; n49493_not
g98816 not n29099 ; n29099_not
g98817 not n33599 ; n33599_not
g98818 not n48980 ; n48980_not
g98819 not n49484 ; n49484_not
g98820 not n31799 ; n31799_not
g98821 not n49709 ; n49709_not
g98822 not n49565 ; n49565_not
g98823 not n48836 ; n48836_not
g98824 not n33986 ; n33986_not
g98825 not n43886 ; n43886_not
g98826 not n49718 ; n49718_not
g98827 not n34499 ; n34499_not
g98828 not n53687 ; n53687_not
g98829 not n53957 ; n53957_not
g98830 not n18569 ; n18569_not
g98831 not n29369 ; n29369_not
g98832 not n29288 ; n29288_not
g98833 not n57278 ; n57278_not
g98834 not n56378 ; n56378_not
g98835 not n49448 ; n49448_not
g98836 not n29378 ; n29378_not
g98837 not n50879 ; n50879_not
g98838 not n49781 ; n49781_not
g98839 not n54488 ; n54488_not
g98840 not n18785 ; n18785_not
g98841 not n53966 ; n53966_not
g98842 not n19937 ; n19937_not
g98843 not n38585 ; n38585_not
g98844 not n38594 ; n38594_not
g98845 not n56387 ; n56387_not
g98846 not n53696 ; n53696_not
g98847 not n56873 ; n56873_not
g98848 not n46685 ; n46685_not
g98849 not n33797 ; n33797_not
g98850 not n19964 ; n19964_not
g98851 not n19955 ; n19955_not
g98852 not n49763 ; n49763_not
g98853 not n53678 ; n53678_not
g98854 not n29297 ; n29297_not
g98855 not n33896 ; n33896_not
g98856 not n56864 ; n56864_not
g98857 not n33779 ; n33779_not
g98858 not n44939 ; n44939_not
g98859 not n56369 ; n56369_not
g98860 not n33788 ; n33788_not
g98861 not n53948 ; n53948_not
g98862 not n49772 ; n49772_not
g98863 not n53597 ; n53597_not
g98864 not n38567 ; n38567_not
g98865 not n46478 ; n46478_not
g98866 not n18389 ; n18389_not
g98867 not n56783 ; n56783_not
g98868 not n56558 ; n56558_not
g98869 not n50996 ; n50996_not
g98870 not n44399 ; n44399_not
g98871 not n39089 ; n39089_not
g98872 not n46568 ; n46568_not
g98873 not n54299 ; n54299_not
g98874 not n29648 ; n29648_not
g98875 not n46487 ; n46487_not
g98876 not n49358 ; n49358_not
g98877 not n49943 ; n49943_not
g98878 not n19694 ; n19694_not
g98879 not n29792 ; n29792_not
g98880 not n56567 ; n56567_not
g98881 not n46883 ; n46883_not
g98882 not n29765 ; n29765_not
g98883 not n38468 ; n38468_not
g98884 not n53849 ; n53849_not
g98885 not n39098 ; n39098_not
g98886 not n43859 ; n43859_not
g98887 not n50978 ; n50978_not
g98888 not n29729 ; n29729_not
g98889 not n33977 ; n33977_not
g98890 not n19766 ; n19766_not
g98891 not n18299 ; n18299_not
g98892 not n17948 ; n17948_not
g98893 not n56756 ; n56756_not
g98894 not n29756 ; n29756_not
g98895 not a[11] ; a[11]_not
g98896 not n38279 ; n38279_not
g98897 not n44786 ; n44786_not
g98898 not n56765 ; n56765_not
g98899 not n46766 ; n46766_not
g98900 not n19757 ; n19757_not
g98901 not n19748 ; n19748_not
g98902 not n44885 ; n44885_not
g98903 not n19739 ; n19739_not
g98904 not n49934 ; n49934_not
g98905 not n29774 ; n29774_not
g98906 not n33995 ; n33995_not
g98907 not n44858 ; n44858_not
g98908 not n46892 ; n46892_not
g98909 not n46748 ; n46748_not
g98910 not n57089 ; n57089_not
g98911 not n19667 ; n19667_not
g98912 not n38297 ; n38297_not
g98913 not n17993 ; n17993_not
g98914 not n44867 ; n44867_not
g98915 not n56828 ; n56828_not
g98916 not n17966 ; n17966_not
g98917 not n49970 ; n49970_not
g98918 not n44795 ; n44795_not
g98919 not n19298 ; n19298_not
g98920 not n17975 ; n17975_not
g98921 not n53876 ; n53876_not
g98922 not n53885 ; n53885_not
g98923 not n19658 ; n19658_not
g98924 not n17984 ; n17984_not
g98925 not n46757 ; n46757_not
g98926 not n46496 ; n46496_not
g98927 not n19649 ; n19649_not
g98928 not n46865 ; n46865_not
g98929 not n19685 ; n19685_not
g98930 not n54398 ; n54398_not
g98931 not n18479 ; n18479_not
g98932 not n17957 ; n17957_not
g98933 not n50969 ; n50969_not
g98934 not n56576 ; n56576_not
g98935 not n46739 ; n46739_not
g98936 not n49952 ; n49952_not
g98937 not n53858 ; n53858_not
g98938 not n53894 ; n53894_not
g98939 not n19676 ; n19676_not
g98940 not n44876 ; n44876_not
g98941 not n57098 ; n57098_not
g98942 not n38288 ; n38288_not
g98943 not n18497 ; n18497_not
g98944 not n49961 ; n49961_not
g98945 not n56729 ; n56729_not
g98946 not n56585 ; n56585_not
g98947 not n46874 ; n46874_not
g98948 not n29819 ; n29819_not
g98949 not n53867 ; n53867_not
g98950 not n33968 ; n33968_not
g98951 not n33959 ; n33959_not
g98952 not n18749 ; n18749_not
g98953 not n19595 ; n19595_not
g98954 not n56486 ; n56486_not
g98955 not n46946 ; n46946_not
g98956 not n46937 ; n46937_not
g98957 not n29594 ; n29594_not
g98958 not n57179 ; n57179_not
g98959 not n43877 ; n43877_not
g98960 not n44498 ; n44498_not
g98961 not n54497 ; n54497_not
g98962 not n53777 ; n53777_not
g98963 not n44489 ; n44489_not
g98964 not n33887 ; n33887_not
g98965 not n38972 ; n38972_not
g98966 not n18488 ; n18488_not
g98967 not n49880 ; n49880_not
g98968 not n56495 ; n56495_not
g98969 not n56468 ; n56468_not
g98970 not n49862 ; n49862_not
g98971 not n29567 ; n29567_not
g98972 not n44768 ; n44768_not
g98973 not n38648 ; n38648_not
g98974 not n53759 ; n53759_not
g98975 not n33878 ; n33878_not
g98976 not n18695 ; n18695_not
g98977 not n38198 ; n38198_not
g98978 not n29576 ; n29576_not
g98979 not n57188 ; n57188_not
g98980 not n46955 ; n46955_not
g98981 not n29477 ; n29477_not
g98982 not n56477 ; n56477_not
g98983 not n19829 ; n19829_not
g98984 not n43994 ; n43994_not
g98985 not n29585 ; n29585_not
g98986 not n38558 ; n38558_not
g98987 not n54569 ; n54569_not
g98988 not n49871 ; n49871_not
g98989 not n53768 ; n53768_not
g98990 not n46856 ; n46856_not
g98991 not n49907 ; n49907_not
g98992 not n44894 ; n44894_not
g98993 not n19775 ; n19775_not
g98994 not n49916 ; n49916_not
g98995 not n56774 ; n56774_not
g98996 not n49925 ; n49925_not
g98997 not n56549 ; n56549_not
g98998 not n53786 ; n53786_not
g98999 not n29639 ; n29639_not
g99000 not n46928 ; n46928_not
g99001 not n43868 ; n43868_not
g99002 not n38981 ; n38981_not
g99003 not n56738 ; n56738_not
g99004 not n53795 ; n53795_not
g99005 not n44777 ; n44777_not
g99006 not n46919 ; n46919_not
g99007 not n53399 ; n53399_not
g99008 not n17939 ; n17939_not
g99009 not n19784 ; n19784_not
g99010 not n48854 ; n48854_not
g99011 not n32879 ; n32879_not
g99012 not n48845 ; n48845_not
g99013 not n56945 ; n56945_not
g99014 not n56954 ; n56954_not
g99015 not n27974 ; n27974_not
g99016 not n38099 ; n38099_not
g99017 not n28694 ; n28694_not
g99018 not n32888 ; n32888_not
g99019 not n53498 ; n53498_not
g99020 not n19793 ; n19793_not
g99021 not n44678 ; n44678_not
g99022 not n48881 ; n48881_not
g99023 not n18866 ; n18866_not
g99024 not n48872 ; n48872_not
g99025 not n48863 ; n48863_not
g99026 not n49547 ; n49547_not
g99027 not n57449 ; n57449_not
g99028 not n28676 ; n28676_not
g99029 not n29963 ; n29963_not
g99030 not n44669 ; n44669_not
g99031 not n49592 ; n49592_not
g99032 not n19487 ; n19487_not
g99033 not n28766 ; n28766_not
g99034 not n32897 ; n32897_not
g99035 not n56936 ; n56936_not
g99036 not n32969 ; n32969_not
g99037 not n32978 ; n32978_not
g99038 not n28784 ; n28784_not
g99039 not n18938 ; n18938_not
g99040 not n54695 ; n54695_not
g99041 not n56981 ; n56981_not
g99042 not n43679 ; n43679_not
g99043 not n49574 ; n49574_not
g99044 not n18929 ; n18929_not
g99045 not n19838 ; n19838_not
g99046 not n29972 ; n29972_not
g99047 not n49583 ; n49583_not
g99048 not n28748 ; n28748_not
g99049 not n18668 ; n18668_not
g99050 not n55946 ; n55946_not
g99051 not n46649 ; n46649_not
g99052 not n38387 ; n38387_not
g99053 not n28568 ; n28568_not
g99054 not n54758 ; n54758_not
g99055 not n46298 ; n46298_not
g99056 not n18893 ; n18893_not
g99057 not n56279 ; n56279_not
g99058 not n48962 ; n48962_not
g99059 not n28586 ; n28586_not
g99060 not n57476 ; n57476_not
g99061 not n44687 ; n44687_not
g99062 not n49457 ; n49457_not
g99063 not n32699 ; n32699_not
g99064 not n18875 ; n18875_not
g99065 not n27884 ; n27884_not
g99066 not n19469 ; n19469_not
g99067 not n56963 ; n56963_not
g99068 not n56990 ; n56990_not
g99069 not n17858 ; n17858_not
g99070 not n46289 ; n46289_not
g99071 not n54767 ; n54767_not
g99072 not n57494 ; n57494_not
g99073 not n44696 ; n44696_not
g99074 not n18884 ; n18884_not
g99075 not n29990 ; n29990_not
g99076 not n48917 ; n48917_not
g99077 not n48908 ; n48908_not
g99078 not n18659 ; n18659_not
g99079 not n43598 ; n43598_not
g99080 not n50897 ; n50897_not
g99081 not n46793 ; n46793_not
g99082 not n49529 ; n49529_not
g99083 not n32798 ; n32798_not
g99084 not n28658 ; n28658_not
g99085 not n18398 ; n18398_not
g99086 not n48890 ; n48890_not
g99087 not n29981 ; n29981_not
g99088 not n57458 ; n57458_not
g99089 not n43589 ; n43589_not
g99090 not n48953 ; n48953_not
g99091 not n56288 ; n56288_not
g99092 not n54749 ; n54749_not
g99093 not n57467 ; n57467_not
g99094 not n56297 ; n56297_not
g99095 not n31979 ; n31979_not
g99096 not n48944 ; n48944_not
g99097 not n19478 ; n19478_not
g99098 not n55991 ; n55991_not
g99099 not n48935 ; n48935_not
g99100 not n48926 ; n48926_not
g99101 not n32789 ; n32789_not
g99102 not n28946 ; n28946_not
g99103 not n18983 ; n18983_not
g99104 not n57377 ; n57377_not
g99105 not n49673 ; n49673_not
g99106 not n43796 ; n43796_not
g99107 not n28955 ; n28955_not
g99108 not n43697 ; n43697_not
g99109 not n44975 ; n44975_not
g99110 not n19973 ; n19973_not
g99111 not n43778 ; n43778_not
g99112 not n28892 ; n28892_not
g99113 not n38369 ; n38369_not
g99114 not n31898 ; n31898_not
g99115 not n50987 ; n50987_not
g99116 not n49655 ; n49655_not
g99117 not n38396 ; n38396_not
g99118 not n17768 ; n17768_not
g99119 not n28919 ; n28919_not
g99120 not n29945 ; n29945_not
g99121 not n31889 ; n31889_not
g99122 not n46784 ; n46784_not
g99123 not n28937 ; n28937_not
g99124 not n49664 ; n49664_not
g99125 not n18992 ; n18992_not
g99126 not n43787 ; n43787_not
g99127 not n19397 ; n19397_not
g99128 not n28991 ; n28991_not
g99129 not n28973 ; n28973_not
g99130 not n53489 ; n53489_not
g99131 not n54479 ; n54479_not
g99132 not n46829 ; n46829_not
g99133 not n44957 ; n44957_not
g99134 not n49691 ; n49691_not
g99135 not n46667 ; n46667_not
g99136 not n56909 ; n56909_not
g99137 not n49682 ; n49682_not
g99138 not n55856 ; n55856_not
g99139 not n37964 ; n37964_not
g99140 not n28964 ; n28964_not
g99141 not n44966 ; n44966_not
g99142 not n28982 ; n28982_not
g99143 not n31988 ; n31988_not
g99144 not n49538 ; n49538_not
g99145 not n49619 ; n49619_not
g99146 not n28838 ; n28838_not
g99147 not n43769 ; n43769_not
g99148 not n18956 ; n18956_not
g99149 not n49628 ; n49628_not
g99150 not n54677 ; n54677_not
g99151 not n56918 ; n56918_not
g99152 not n28856 ; n28856_not
g99153 not n18857 ; n18857_not
g99154 not n38378 ; n38378_not
g99155 not n18947 ; n18947_not
g99156 not n19883 ; n19883_not
g99157 not n32996 ; n32996_not
g99158 not n54686 ; n54686_not
g99159 not n34868 ; n34868_not
g99160 not n44993 ; n44993_not
g99161 not n54668 ; n54668_not
g99162 not n29936 ; n29936_not
g99163 not n46658 ; n46658_not
g99164 not n28874 ; n28874_not
g99165 not n44984 ; n44984_not
g99166 not n19928 ; n19928_not
g99167 not n19496 ; n19496_not
g99168 not n49646 ; n49646_not
g99169 not n18677 ; n18677_not
g99170 not n54659 ; n54659_not
g99171 not n57395 ; n57395_not
g99172 not n18848 ; n18848_not
g99173 not n49637 ; n49637_not
g99174 not n18974 ; n18974_not
g99175 not n18839 ; n18839_not
g99176 not n18965 ; n18965_not
g99177 not n57386 ; n57386_not
g99178 not n32987 ; n32987_not
g99179 not n18588 ; n18588_not
g99180 not n46785 ; n46785_not
g99181 not n17958 ; n17958_not
g99182 not n46776 ; n46776_not
g99183 not n46758 ; n46758_not
g99184 not b[11] ; b[11]_not
g99185 not n17976 ; n17976_not
g99186 not n53589 ; n53589_not
g99187 not n53598 ; n53598_not
g99188 not n47874 ; n47874_not
g99189 not n38892 ; n38892_not
g99190 not n18696 ; n18696_not
g99191 not n38919 ; n38919_not
g99192 not n46794 ; n46794_not
g99193 not n18669 ; n18669_not
g99194 not n47883 ; n47883_not
g99195 not n18678 ; n18678_not
g99196 not n38928 ; n38928_not
g99197 not n17994 ; n17994_not
g99198 not b[20] ; b[20]_not
g99199 not n17985 ; n17985_not
g99200 not n19398 ; n19398_not
g99201 not n17967 ; n17967_not
g99202 not n18687 ; n18687_not
g99203 not n37488 ; n37488_not
g99204 not n53994 ; n53994_not
g99205 not n19389 ; n19389_not
g99206 not n39909 ; n39909_not
g99207 not n46767 ; n46767_not
g99208 not n17949 ; n17949_not
g99209 not n39891 ; n39891_not
g99210 not n16599 ; n16599_not
g99211 not n38685 ; n38685_not
g99212 not n18975 ; n18975_not
g99213 not n38874 ; n38874_not
g99214 not n39972 ; n39972_not
g99215 not n46659 ; n46659_not
g99216 not n48099 ; n48099_not
g99217 not n38694 ; n38694_not
g99218 not n18966 ; n18966_not
g99219 not n38865 ; n38865_not
g99220 not n39981 ; n39981_not
g99221 not n18957 ; n18957_not
g99222 not n24879 ; n24879_not
g99223 not n18849 ; n18849_not
g99224 not n38739 ; n38739_not
g99225 not n38748 ; n38748_not
g99226 not n18948 ; n18948_not
g99227 not a[12] ; a[12]_not
g99228 not n39954 ; n39954_not
g99229 not n38676 ; n38676_not
g99230 not n18993 ; n18993_not
g99231 not n24789 ; n24789_not
g99232 not n46668 ; n46668_not
g99233 not n39963 ; n39963_not
g99234 not n18984 ; n18984_not
g99235 not n24798 ; n24798_not
g99236 not n38883 ; n38883_not
g99237 not n52698 ; n52698_not
g99238 not n18399 ; n18399_not
g99239 not n24987 ; n24987_not
g99240 not n18867 ; n18867_not
g99241 not n18894 ; n18894_not
g99242 not n24996 ; n24996_not
g99243 not n38775 ; n38775_not
g99244 not n45768 ; n45768_not
g99245 not n38766 ; n38766_not
g99246 not n18885 ; n18885_not
g99247 not n15699 ; n15699_not
g99248 not n39567 ; n39567_not
g99249 not n48189 ; n48189_not
g99250 not n18876 ; n18876_not
g99251 not n39099 ; n39099_not
g99252 not n24888 ; n24888_not
g99253 not n38856 ; n38856_not
g99254 not n24897 ; n24897_not
g99255 not n45795 ; n45795_not
g99256 not n18939 ; n18939_not
g99257 not n38847 ; n38847_not
g99258 not n45786 ; n45786_not
g99259 not n18858 ; n18858_not
g99260 not n38838 ; n38838_not
g99261 not n38829 ; n38829_not
g99262 not n39990 ; n39990_not
g99263 not n38793 ; n38793_not
g99264 not n38757 ; n38757_not
g99265 not n24969 ; n24969_not
g99266 not n15789 ; n15789_not
g99267 not n24978 ; n24978_not
g99268 not n38784 ; n38784_not
g99269 not n38973 ; n38973_not
g99270 not n36975 ; n36975_not
g99271 not n47919 ; n47919_not
g99272 not n18759 ; n18759_not
g99273 not n38982 ; n38982_not
g99274 not n18768 ; n18768_not
g99275 not n47928 ; n47928_not
g99276 not n36984 ; n36984_not
g99277 not n18777 ; n18777_not
g99278 not n46578 ; n46578_not
g99279 not n45876 ; n45876_not
g99280 not n18786 ; n18786_not
g99281 not n47946 ; n47946_not
g99282 not n18795 ; n18795_not
g99283 not n38964 ; n38964_not
g99284 not n38658 ; n38658_not
g99285 not n38955 ; n38955_not
g99286 not n47964 ; n47964_not
g99287 not n39936 ; n39936_not
g99288 not n37479 ; n37479_not
g99289 not n39198 ; n39198_not
g99290 not n54399 ; n54399_not
g99291 not n18498 ; n18498_not
g99292 not n38937 ; n38937_not
g99293 not n18597 ; n18597_not
g99294 not n39918 ; n39918_not
g99295 not n46749 ; n46749_not
g99296 not n38946 ; n38946_not
g99297 not n38478 ; n38478_not
g99298 not n38469 ; n38469_not
g99299 not n45885 ; n45885_not
g99300 not n18489 ; n18489_not
g99301 not n39927 ; n39927_not
g99302 not n39945 ; n39945_not
g99303 not n46686 ; n46686_not
g99304 not n47991 ; n47991_not
g99305 not n46596 ; n46596_not
g99306 not n37389 ; n37389_not
g99307 not n46677 ; n46677_not
g99308 not n39594 ; n39594_not
g99309 not n37299 ; n37299_not
g99310 not n47973 ; n47973_not
g99311 not n38667 ; n38667_not
g99312 not n37398 ; n37398_not
g99313 not n46587 ; n46587_not
g99314 not n46695 ; n46695_not
g99315 not n23889 ; n23889_not
g99316 not n24699 ; n24699_not
g99317 not n45858 ; n45858_not
g99318 not n47487 ; n47487_not
g99319 not n16968 ; n16968_not
g99320 not n17886 ; n17886_not
g99321 not n19974 ; n19974_not
g99322 not n37974 ; n37974_not
g99323 not n37965 ; n37965_not
g99324 not n53499 ; n53499_not
g99325 not n47496 ; n47496_not
g99326 not n19983 ; n19983_not
g99327 not n39288 ; n39288_not
g99328 not n37884 ; n37884_not
g99329 not n53796 ; n53796_not
g99330 not n39666 ; n39666_not
g99331 not n37875 ; n37875_not
g99332 not n54894 ; n54894_not
g99333 not n16977 ; n16977_not
g99334 not n39279 ; n39279_not
g99335 not n53787 ; n53787_not
g99336 not n39459 ; n39459_not
g99337 not n16959 ; n16959_not
g99338 not n17778 ; n17778_not
g99339 not n54867 ; n54867_not
g99340 not n19929 ; n19929_not
g99341 not n47469 ; n47469_not
g99342 not n17598 ; n17598_not
g99343 not n17769 ; n17769_not
g99344 not n19938 ; n19938_not
g99345 not n39639 ; n39639_not
g99346 not n39648 ; n39648_not
g99347 not n54876 ; n54876_not
g99348 not n17589 ; n17589_not
g99349 not n47478 ; n47478_not
g99350 not n39297 ; n39297_not
g99351 not n37893 ; n37893_not
g99352 not n54885 ; n54885_not
g99353 not n19965 ; n19965_not
g99354 not n53679 ; n53679_not
g99355 not n38559 ; n38559_not
g99356 not n53769 ; n53769_not
g99357 not n38298 ; n38298_not
g99358 not n19947 ; n19947_not
g99359 not n47559 ; n47559_not
g99360 not n38289 ; n38289_not
g99361 not n53688 ; n53688_not
g99362 not n47568 ; n47568_not
g99363 not n54957 ; n54957_not
g99364 not n47577 ; n47577_not
g99365 not n38577 ; n38577_not
g99366 not n37794 ; n37794_not
g99367 not n47586 ; n47586_not
g99368 not n53697 ; n53697_not
g99369 not n22899 ; n22899_not
g99370 not n38595 ; n38595_not
g99371 not n38199 ; n38199_not
g99372 not n47595 ; n47595_not
g99373 not n54858 ; n54858_not
g99374 not n39684 ; n39684_not
g99375 not n39693 ; n39693_not
g99376 not n19992 ; n19992_not
g99377 not n38487 ; n38487_not
g99378 not n37866 ; n37866_not
g99379 not n17499 ; n17499_not
g99380 not n53778 ; n53778_not
g99381 not n38397 ; n38397_not
g99382 not n37497 ; n37497_not
g99383 not n54939 ; n54939_not
g99384 not n37857 ; n37857_not
g99385 not n38388 ; n38388_not
g99386 not n38379 ; n38379_not
g99387 not n37848 ; n37848_not
g99388 not n37839 ; n37839_not
g99389 not n46398 ; n46398_not
g99390 not n39729 ; n39729_not
g99391 not n37695 ; n37695_not
g99392 not n39549 ; n39549_not
g99393 not n37686 ; n37686_not
g99394 not n39486 ; n39486_not
g99395 not n37677 ; n37677_not
g99396 not n53958 ; n53958_not
g99397 not n37668 ; n37668_not
g99398 not n37659 ; n37659_not
g99399 not n17877 ; n17877_not
g99400 not n54795 ; n54795_not
g99401 not n39495 ; n39495_not
g99402 not n47379 ; n47379_not
g99403 not n19785 ; n19785_not
g99404 not n53967 ; n53967_not
g99405 not n37983 ; n37983_not
g99406 not n19794 ; n19794_not
g99407 not n47388 ; n47388_not
g99408 not n39558 ; n39558_not
g99409 not n39477 ; n39477_not
g99410 not n53895 ; n53895_not
g99411 not n17859 ; n17859_not
g99412 not n47397 ; n47397_not
g99413 not n54768 ; n54768_not
g99414 not n17895 ; n17895_not
g99415 not n54777 ; n54777_not
g99416 not n37785 ; n37785_not
g99417 not n37776 ; n37776_not
g99418 not n54759 ; n54759_not
g99419 not n37767 ; n37767_not
g99420 not n37758 ; n37758_not
g99421 not n46299 ; n46299_not
g99422 not n37749 ; n37749_not
g99423 not n47298 ; n47298_not
g99424 not n53949 ; n53949_not
g99425 not n54786 ; n54786_not
g99426 not n17868 ; n17868_not
g99427 not n45696 ; n45696_not
g99428 not n19875 ; n19875_not
g99429 not n37938 ; n37938_not
g99430 not n54687 ; n54687_not
g99431 not n17697 ; n17697_not
g99432 not n39396 ; n39396_not
g99433 not n37929 ; n37929_not
g99434 not n19884 ; n19884_not
g99435 not n45759 ; n45759_not
g99436 not n54849 ; n54849_not
g99437 not n17679 ; n17679_not
g99438 not n19893 ; n19893_not
g99439 not n39387 ; n39387_not
g99440 not n54678 ; n54678_not
g99441 not n39378 ; n39378_not
g99442 not n39468 ; n39468_not
g99443 not n39369 ; n39369_not
g99444 not n54669 ; n54669_not
g99445 not n53976 ; n53976_not
g99446 not n53886 ; n53886_not
g99447 not n53877 ; n53877_not
g99448 not n19839 ; n19839_not
g99449 not n53985 ; n53985_not
g99450 not n19848 ; n19848_not
g99451 not n17787 ; n17787_not
g99452 not n39576 ; n39576_not
g99453 not n53868 ; n53868_not
g99454 not n54696 ; n54696_not
g99455 not n53859 ; n53859_not
g99456 not n47775 ; n47775_not
g99457 not n46866 ; n46866_not
g99458 not n37596 ; n37596_not
g99459 not n45984 ; n45984_not
g99460 not n46857 ; n46857_not
g99461 not n47784 ; n47784_not
g99462 not n45894 ; n45894_not
g99463 not n45975 ; n45975_not
g99464 not n54498 ; n54498_not
g99465 not n46497 ; n46497_not
g99466 not n46488 ; n46488_not
g99467 not n16896 ; n16896_not
g99468 not n19596 ; n19596_not
g99469 not n47793 ; n47793_not
g99470 not n16887 ; n16887_not
g99471 not n39864 ; n39864_not
g99472 not n46848 ; n46848_not
g99473 not n19587 ; n19587_not
g99474 not n39846 ; n39846_not
g99475 not n46884 ; n46884_not
g99476 not n54588 ; n54588_not
g99477 not n19686 ; n19686_not
g99478 not n19677 ; n19677_not
g99479 not n54579 ; n54579_not
g99480 not n47739 ; n47739_not
g99481 not n46875 ; n46875_not
g99482 not n47748 ; n47748_not
g99483 not n39855 ; n39855_not
g99484 not n16986 ; n16986_not
g99485 not n19668 ; n19668_not
g99486 not n47757 ; n47757_not
g99487 not n47766 ; n47766_not
g99488 not n38568 ; n38568_not
g99489 not n19659 ; n19659_not
g99490 not n45993 ; n45993_not
g99491 not n16797 ; n16797_not
g99492 not n47838 ; n47838_not
g99493 not n16788 ; n16788_not
g99494 not n39873 ; n39873_not
g99495 not n16779 ; n16779_not
g99496 not n19488 ; n19488_not
g99497 not n45948 ; n45948_not
g99498 not n45939 ; n45939_not
g99499 not n47856 ; n47856_not
g99500 not n19479 ; n19479_not
g99501 not n39882 ; n39882_not
g99502 not n16698 ; n16698_not
g99503 not n16689 ; n16689_not
g99504 not n23799 ; n23799_not
g99505 not n16878 ; n16878_not
g99506 not n54489 ; n54489_not
g99507 not n37578 ; n37578_not
g99508 not n19578 ; n19578_not
g99509 not n37569 ; n37569_not
g99510 not n19767 ; n19767_not
g99511 not n45966 ; n45966_not
g99512 not n16869 ; n16869_not
g99513 not n19569 ; n19569_not
g99514 not n46839 ; n46839_not
g99515 not n45957 ; n45957_not
g99516 not n18579 ; n18579_not
g99517 not n47829 ; n47829_not
g99518 not n19497 ; n19497_not
g99519 not n39765 ; n39765_not
g99520 not n46983 ; n46983_not
g99521 not n46974 ; n46974_not
g99522 not n19857 ; n19857_not
g99523 not n39774 ; n39774_not
g99524 not n46965 ; n46965_not
g99525 not n39783 ; n39783_not
g99526 not n47649 ; n47649_not
g99527 not n46956 ; n46956_not
g99528 not n39738 ; n39738_not
g99529 not n38649 ; n38649_not
g99530 not n54597 ; n54597_not
g99531 not n22989 ; n22989_not
g99532 not n17688 ; n17688_not
g99533 not n22998 ; n22998_not
g99534 not n54975 ; n54975_not
g99535 not n54984 ; n54984_not
g99536 not n39747 ; n39747_not
g99537 not n46992 ; n46992_not
g99538 not n39756 ; n39756_not
g99539 not n47694 ; n47694_not
g99540 not n39819 ; n39819_not
g99541 not n37587 ; n37587_not
g99542 not n39828 ; n39828_not
g99543 not n19758 ; n19758_not
g99544 not n46893 ; n46893_not
g99545 not n39837 ; n39837_not
g99546 not n39657 ; n39657_not
g99547 not n19695 ; n19695_not
g99548 not n47658 ; n47658_not
g99549 not n46947 ; n46947_not
g99550 not n46938 ; n46938_not
g99551 not n39792 ; n39792_not
g99552 not n47667 ; n47667_not
g99553 not n45849 ; n45849_not
g99554 not n47676 ; n47676_not
g99555 not n46929 ; n46929_not
g99556 not n47685 ; n47685_not
g99557 not n49593 ; n49593_not
g99558 not n28758 ; n28758_not
g99559 not n49584 ; n49584_not
g99560 not n55947 ; n55947_not
g99561 not n49575 ; n49575_not
g99562 not n27984 ; n27984_not
g99563 not n55956 ; n55956_not
g99564 not n44994 ; n44994_not
g99565 not n49557 ; n49557_not
g99566 not n28686 ; n28686_not
g99567 not n44985 ; n44985_not
g99568 not n49539 ; n49539_not
g99569 not n44976 ; n44976_not
g99570 not n50898 ; n50898_not
g99571 not n43599 ; n43599_not
g99572 not n28668 ; n28668_not
g99573 not n49638 ; n49638_not
g99574 not n28866 ; n28866_not
g99575 not n43779 ; n43779_not
g99576 not n55893 ; n55893_not
g99577 not n34869 ; n34869_not
g99578 not n49629 ; n49629_not
g99579 not n28848 ; n28848_not
g99580 not n43698 ; n43698_not
g99581 not n28794 ; n28794_not
g99582 not n49548 ; n49548_not
g99583 not n43689 ; n43689_not
g99584 not n55938 ; n55938_not
g99585 not n28776 ; n28776_not
g99586 not n49449 ; n49449_not
g99587 not n34788 ; n34788_not
g99588 not n34779 ; n34779_not
g99589 not n28488 ; n28488_not
g99590 not n49395 ; n49395_not
g99591 not n49377 ; n49377_not
g99592 not n28398 ; n28398_not
g99593 not n49359 ; n49359_not
g99594 not n44895 ; n44895_not
g99595 not n44886 ; n44886_not
g99596 not n27786 ; n27786_not
g99597 not n44877 ; n44877_not
g99598 not n27795 ; n27795_not
g99599 not n28299 ; n28299_not
g99600 not n55983 ; n55983_not
g99601 not n50889 ; n50889_not
g99602 not n55992 ; n55992_not
g99603 not n28596 ; n28596_not
g99604 not n44967 ; n44967_not
g99605 not n49494 ; n49494_not
g99606 not n49485 ; n49485_not
g99607 not n28578 ; n28578_not
g99608 not n44958 ; n44958_not
g99609 not n44949 ; n44949_not
g99610 not n27894 ; n27894_not
g99611 not n49467 ; n49467_not
g99612 not n29379 ; n29379_not
g99613 not n49773 ; n49773_not
g99614 not n29298 ; n29298_not
g99615 not n49764 ; n49764_not
g99616 not n49458 ; n49458_not
g99617 not n29289 ; n29289_not
g99618 not n49755 ; n49755_not
g99619 not n49746 ; n49746_not
g99620 not n49737 ; n49737_not
g99621 not n43896 ; n43896_not
g99622 not n49728 ; n49728_not
g99623 not n29199 ; n29199_not
g99624 not n49719 ; n49719_not
g99625 not n29478 ; n29478_not
g99626 not n49809 ; n49809_not
g99627 not n29388 ; n29388_not
g99628 not n56676 ; n56676_not
g99629 not n49791 ; n49791_not
g99630 not n29397 ; n29397_not
g99631 not n55794 ; n55794_not
g99632 not n34887 ; n34887_not
g99633 not n49782 ; n49782_not
g99634 not n28956 ; n28956_not
g99635 not n55866 ; n55866_not
g99636 not n49674 ; n49674_not
g99637 not n50997 ; n50997_not
g99638 not n28947 ; n28947_not
g99639 not n50988 ; n50988_not
g99640 not n49665 ; n49665_not
g99641 not n49656 ; n49656_not
g99642 not n34878 ; n34878_not
g99643 not n50979 ; n50979_not
g99644 not n43788 ; n43788_not
g99645 not n49647 ; n49647_not
g99646 not a[30] ; a[30]_not
g99647 not n28884 ; n28884_not
g99648 not n43878 ; n43878_not
g99649 not n49692 ; n49692_not
g99650 not n43869 ; n43869_not
g99651 not n28992 ; n28992_not
g99652 not n28983 ; n28983_not
g99653 not n55848 ; n55848_not
g99654 not n49683 ; n49683_not
g99655 not n28974 ; n28974_not
g99656 not n28965 ; n28965_not
g99657 not n55857 ; n55857_not
g99658 not n48693 ; n48693_not
g99659 not n27669 ; n27669_not
g99660 not n35769 ; n35769_not
g99661 not n42798 ; n42798_not
g99662 not n42789 ; n42789_not
g99663 not n26976 ; n26976_not
g99664 not n51897 ; n51897_not
g99665 not n26985 ; n26985_not
g99666 not a[21] ; a[21]_not
g99667 not n35589 ; n35589_not
g99668 not n51888 ; n51888_not
g99669 not n51969 ; n51969_not
g99670 not n35598 ; n35598_not
g99671 not n27777 ; n27777_not
g99672 not n27768 ; n27768_not
g99673 not n27759 ; n27759_not
g99674 not n44697 ; n44697_not
g99675 not n42879 ; n42879_not
g99676 not n44688 ; n44688_not
g99677 not n27696 ; n27696_not
g99678 not n44679 ; n44679_not
g99679 not n27687 ; n27687_not
g99680 not n27678 ; n27678_not
g99681 not n26967 ; n26967_not
g99682 not n27489 ; n27489_not
g99683 not n35985 ; n35985_not
g99684 not n35976 ; n35976_not
g99685 not n35967 ; n35967_not
g99686 not n27399 ; n27399_not
g99687 not n48738 ; n48738_not
g99688 not n41898 ; n41898_not
g99689 not n35958 ; n35958_not
g99690 not n35949 ; n35949_not
g99691 not n55875 ; n55875_not
g99692 not n35895 ; n35895_not
g99693 not n48747 ; n48747_not
g99694 not n44589 ; n44589_not
g99695 not n27597 ; n27597_not
g99696 not n51978 ; n51978_not
g99697 not n55965 ; n55965_not
g99698 not n27588 ; n27588_not
g99699 not n51987 ; n51987_not
g99700 not n42699 ; n42699_not
g99701 not n27579 ; n27579_not
g99702 not n51996 ; n51996_not
g99703 not n35994 ; n35994_not
g99704 not n27498 ; n27498_not
g99705 not n41799 ; n41799_not
g99706 not n42888 ; n42888_not
g99707 not n35697 ; n35697_not
g99708 not n48576 ; n48576_not
g99709 not n42897 ; n42897_not
g99710 not n42969 ; n42969_not
g99711 not n42978 ; n42978_not
g99712 not n42987 ; n42987_not
g99713 not n27993 ; n27993_not
g99714 not n27975 ; n27975_not
g99715 not n27966 ; n27966_not
g99716 not n42996 ; n42996_not
g99717 not n44796 ; n44796_not
g99718 not n27948 ; n27948_not
g99719 not n27849 ; n27849_not
g99720 not n44868 ; n44868_not
g99721 not n44859 ; n44859_not
g99722 not n49296 ; n49296_not
g99723 not n35499 ; n35499_not
g99724 not n27876 ; n27876_not
g99725 not n27885 ; n27885_not
g99726 not n27939 ; n27939_not
g99727 not n48558 ; n48558_not
g99728 not n48567 ; n48567_not
g99729 not n35688 ; n35688_not
g99730 not n44769 ; n44769_not
g99731 not n48648 ; n48648_not
g99732 not n48657 ; n48657_not
g99733 not n48666 ; n48666_not
g99734 not n44787 ; n44787_not
g99735 not n44778 ; n44778_not
g99736 not n51798 ; n51798_not
g99737 not n27858 ; n27858_not
g99738 not n33987 ; n33987_not
g99739 not n56577 ; n56577_not
g99740 not n57099 ; n57099_not
g99741 not n56586 ; n56586_not
g99742 not n56739 ; n56739_not
g99743 not n56595 ; n56595_not
g99744 not n44499 ; n44499_not
g99745 not n56487 ; n56487_not
g99746 not n33888 ; n33888_not
g99747 not n56496 ; n56496_not
g99748 not n33897 ; n33897_not
g99749 not n56784 ; n56784_not
g99750 not n56775 ; n56775_not
g99751 not n33969 ; n33969_not
g99752 not n56766 ; n56766_not
g99753 not n33978 ; n33978_not
g99754 not n56559 ; n56559_not
g99755 not n33996 ; n33996_not
g99756 not n56568 ; n56568_not
g99757 not n56199 ; n56199_not
g99758 not n29982 ; n29982_not
g99759 not n56946 ; n56946_not
g99760 not n29973 ; n29973_not
g99761 not n56928 ; n56928_not
g99762 not n33789 ; n33789_not
g99763 not n29955 ; n29955_not
g99764 not n33798 ; n33798_not
g99765 not n29829 ; n29829_not
g99766 not n29838 ; n29838_not
g99767 not n29847 ; n29847_not
g99768 not n29856 ; n29856_not
g99769 not n29937 ; n29937_not
g99770 not n56289 ; n56289_not
g99771 not n56649 ; n56649_not
g99772 not n56658 ; n56658_not
g99773 not n56667 ; n56667_not
g99774 not n56694 ; n56694_not
g99775 not n56685 ; n56685_not
g99776 not n29928 ; n29928_not
g99777 not n56991 ; n56991_not
g99778 not n29946 ; n29946_not
g99779 not n56973 ; n56973_not
g99780 not n50799 ; n50799_not
g99781 not n29991 ; n29991_not
g99782 not n56955 ; n56955_not
g99783 not n43995 ; n43995_not
g99784 not n32979 ; n32979_not
g99785 not n32988 ; n32988_not
g99786 not n31998 ; n31998_not
g99787 not n57396 ; n57396_not
g99788 not n43986 ; n43986_not
g99789 not n32997 ; n32997_not
g99790 not n43977 ; n43977_not
g99791 not n57387 ; n57387_not
g99792 not n31899 ; n31899_not
g99793 not n57378 ; n57378_not
g99794 not n56919 ; n56919_not
g99795 not n43968 ; n43968_not
g99796 not n57486 ; n57486_not
g99797 not n57468 ; n57468_not
g99798 not n31989 ; n31989_not
g99799 not n57459 ; n57459_not
g99800 not n56964 ; n56964_not
g99801 not n56388 ; n56388_not
g99802 not n56397 ; n56397_not
g99803 not n56829 ; n56829_not
g99804 not n30999 ; n30999_not
g99805 not n56469 ; n56469_not
g99806 not n57198 ; n57198_not
g99807 not n56478 ; n56478_not
g99808 not n33879 ; n33879_not
g99809 not n57369 ; n57369_not
g99810 not n43959 ; n43959_not
g99811 not n56298 ; n56298_not
g99812 not n56874 ; n56874_not
g99813 not n57297 ; n57297_not
g99814 not n56865 ; n56865_not
g99815 not n33699 ; n33699_not
g99816 not n56856 ; n56856_not
g99817 not n56379 ; n56379_not
g99818 not n56748 ; n56748_not
g99819 not n29568 ; n29568_not
g99820 not n29676 ; n29676_not
g99821 not n29559 ; n29559_not
g99822 not n29667 ; n29667_not
g99823 not n49890 ; n49890_not
g99824 not n29658 ; n29658_not
g99825 not n29649 ; n29649_not
g99826 not n49881 ; n49881_not
g99827 not n29766 ; n29766_not
g99828 not n34689 ; n34689_not
g99829 not n29694 ; n29694_not
g99830 not n29757 ; n29757_not
g99831 not n34698 ; n34698_not
g99832 not n49926 ; n49926_not
g99833 not n29739 ; n29739_not
g99834 not n49368 ; n49368_not
g99835 not n49917 ; n49917_not
g99836 not n49908 ; n49908_not
g99837 not n29586 ; n29586_not
g99838 not n29577 ; n29577_not
g99839 not n29685 ; n29685_not
g99840 not n43887 ; n43887_not
g99841 not n49854 ; n49854_not
g99842 not n34797 ; n34797_not
g99843 not n49845 ; n49845_not
g99844 not n49836 ; n49836_not
g99845 not n29496 ; n29496_not
g99846 not n49827 ; n49827_not
g99847 not n49818 ; n49818_not
g99848 not n34599 ; n34599_not
g99849 not n29595 ; n29595_not
g99850 not n49872 ; n49872_not
g99851 not n49863 ; n49863_not
g99852 not n29487 ; n29487_not
g99853 not n43797 ; n43797_not
g99854 not n29883 ; n29883_not
g99855 not n29874 ; n29874_not
g99856 not n29865 ; n29865_not
g99857 not n56883 ; n56883_not
g99858 not n29892 ; n29892_not
g99859 not n56793 ; n56793_not
g99860 not n29793 ; n29793_not
g99861 not n49944 ; n49944_not
g99862 not n29784 ; n29784_not
g99863 not n49935 ; n49935_not
g99864 not n49980 ; n49980_not
g99865 not n56838 ; n56838_not
g99866 not n29775 ; n29775_not
g99867 not n49971 ; n49971_not
g99868 not n49962 ; n49962_not
g99869 not n49953 ; n49953_not
g99870 not n26679 ; n26679_not
g99871 not n48279 ; n48279_not
g99872 not n26688 ; n26688_not
g99873 not n40998 ; n40998_not
g99874 not n26697 ; n26697_not
g99875 not n40989 ; n40989_not
g99876 not n36489 ; n36489_not
g99877 not n40899 ; n40899_not
g99878 not n26769 ; n26769_not
g99879 not n36399 ; n36399_not
g99880 not n26778 ; n26778_not
g99881 not n48198 ; n48198_not
g99882 not n48468 ; n48468_not
g99883 not n48459 ; n48459_not
g99884 not n48585 ; n48585_not
g99885 not n36669 ; n36669_not
g99886 not n54993 ; n54993_not
g99887 not n48396 ; n48396_not
g99888 not n48387 ; n48387_not
g99889 not n26589 ; n26589_not
g99890 not n48378 ; n48378_not
g99891 not n26598 ; n26598_not
g99892 not n36588 ; n36588_not
g99893 not n48369 ; n48369_not
g99894 not n36579 ; n36579_not
g99895 not n48297 ; n48297_not
g99896 not n13998 ; n13998_not
g99897 not n48675 ; n48675_not
g99898 not n13989 ; n13989_not
g99899 not n48288 ; n48288_not
g99900 not n35859 ; n35859_not
g99901 not n26895 ; n26895_not
g99902 not n48783 ; n48783_not
g99903 not n48792 ; n48792_not
g99904 not n55785 ; n55785_not
g99905 not n35796 ; n35796_not
g99906 not n26949 ; n26949_not
g99907 not n48819 ; n48819_not
g99908 not n35778 ; n35778_not
g99909 not n35787 ; n35787_not
g99910 not n48828 ; n48828_not
g99911 not n26787 ; n26787_not
g99912 not n26796 ; n26796_not
g99913 not n26859 ; n26859_not
g99914 not n35886 ; n35886_not
g99915 not n54948 ; n54948_not
g99916 not n48765 ; n48765_not
g99917 not n26868 ; n26868_not
g99918 not n35877 ; n35877_not
g99919 not n26877 ; n26877_not
g99920 not n35868 ; n35868_not
g99921 not n26886 ; n26886_not
g99922 not n36939 ; n36939_not
g99923 not n47937 ; n47937_not
g99924 not n14799 ; n14799_not
g99925 not n36894 ; n36894_not
g99926 not n36885 ; n36885_not
g99927 not n36876 ; n36876_not
g99928 not n36867 ; n36867_not
g99929 not n36858 ; n36858_not
g99930 not n45678 ; n45678_not
g99931 not n36849 ; n36849_not
g99932 not n47892 ; n47892_not
g99933 not n14988 ; n14988_not
g99934 not n36993 ; n36993_not
g99935 not n47982 ; n47982_not
g99936 not n14898 ; n14898_not
g99937 not n36957 ; n36957_not
g99938 not n36948 ; n36948_not
g99939 not n14889 ; n14889_not
g99940 not n36777 ; n36777_not
g99941 not n48477 ; n48477_not
g99942 not n48486 ; n48486_not
g99943 not n36768 ; n36768_not
g99944 not n48495 ; n48495_not
g99945 not n36759 ; n36759_not
g99946 not n36696 ; n36696_not
g99947 not n36687 ; n36687_not
g99948 not n36678 ; n36678_not
g99949 not n26499 ; n26499_not
g99950 not n14997 ; n14997_not
g99951 not n14979 ; n14979_not
g99952 not n36597 ; n36597_not
g99953 not n36795 ; n36795_not
g99954 not n47847 ; n47847_not
g99955 not n36786 ; n36786_not
g99956 not n26994 ; n26994_not
g99957 not n41988 ; n41988_not
g99958 not n13899 ; n13899_not
g99959 not n48756 ; n48756_not
g99960 not n41997 ; n41997_not
g99961 not b[21] ; b[21]_not
g99962 not n47677 ; n47677_not
g99963 not n15979 ; n15979_not
g99964 not n39397 ; n39397_not
g99965 not b[12] ; b[12]_not
g99966 not n49963 ; n49963_not
g99967 not n19669 ; n19669_not
g99968 not n29794 ; n29794_not
g99969 not n55588 ; n55588_not
g99970 not n46876 ; n46876_not
g99971 not n46867 ; n46867_not
g99972 not n25987 ; n25987_not
g99973 not n29767 ; n29767_not
g99974 not n53698 ; n53698_not
g99975 not n29677 ; n29677_not
g99976 not n17995 ; n17995_not
g99977 not n55597 ; n55597_not
g99978 not n25996 ; n25996_not
g99979 not b[30] ; b[30]_not
g99980 not n49972 ; n49972_not
g99981 not n36796 ; n36796_not
g99982 not n48478 ; n48478_not
g99983 not n48199 ; n48199_not
g99984 not n29668 ; n29668_not
g99985 not n35977 ; n35977_not
g99986 not n36994 ; n36994_not
g99987 not n18499 ; n18499_not
g99988 not n29776 ; n29776_not
g99989 not n49945 ; n49945_not
g99990 not n15988 ; n15988_not
g99991 not n38569 ; n38569_not
g99992 not n19696 ; n19696_not
g99993 not n50989 ; n50989_not
g99994 not n48469 ; n48469_not
g99995 not n38785 ; n38785_not
g99996 not n47938 ; n47938_not
g99997 not n36778 ; n36778_not
g99998 not n49936 ; n49936_not
g99999 not n56785 ; n56785_not
g100000 not n46894 ; n46894_not
g100001 not n47929 ; n47929_not
g100002 not n50998 ; n50998_not
g100003 not n38794 ; n38794_not
g100004 not n25978 ; n25978_not
g100005 not n56776 ; n56776_not
g100006 not n48766 ; n48766_not
g100007 not n38767 ; n38767_not
g100008 not n47956 ; n47956_not
g100009 not n36985 ; n36985_not
g100010 not n49954 ; n49954_not
g100011 not n29659 ; n29659_not
g100012 not n19678 ; n19678_not
g100013 not n29785 ; n29785_not
g100014 not n47839 ; n47839_not
g100015 not n36787 ; n36787_not
g100016 not n22999 ; n22999_not
g100017 not n19687 ; n19687_not
g100018 not n25969 ; n25969_not
g100019 not n38776 ; n38776_not
g100020 not n46885 ; n46885_not
g100021 not n15997 ; n15997_not
g100022 not n39739 ; n39739_not
g100023 not n43789 ; n43789_not
g100024 not n46498 ; n46498_not
g100025 not n56875 ; n56875_not
g100026 not n17896 ; n17896_not
g100027 not n56866 ; n56866_not
g100028 not n29893 ; n29893_not
g100029 not n48946 ; n48946_not
g100030 not n52798 ; n52798_not
g100031 not n19579 ; n19579_not
g100032 not n29884 ; n29884_not
g100033 not n41998 ; n41998_not
g100034 not n50899 ; n50899_not
g100035 not n19588 ; n19588_not
g100036 not n29875 ; n29875_not
g100037 not n45598 ; n45598_not
g100038 not n46849 ; n46849_not
g100039 not n48883 ; n48883_not
g100040 not n33889 ; n33889_not
g100041 not n25798 ; n25798_not
g100042 not n38848 ; n38848_not
g100043 not n33898 ; n33898_not
g100044 not n55579 ; n55579_not
g100045 not n52789 ; n52789_not
g100046 not n38839 ; n38839_not
g100047 not n33979 ; n33979_not
g100048 not n14989 ; n14989_not
g100049 not n56893 ; n56893_not
g100050 not n33997 ; n33997_not
g100051 not n17878 ; n17878_not
g100052 not n36589 ; n36589_not
g100053 not n17869 ; n17869_not
g100054 not n38749 ; n38749_not
g100055 not n47983 ; n47983_not
g100056 not n29848 ; n29848_not
g100057 not n46858 ; n46858_not
g100058 not n47848 ; n47848_not
g100059 not n49981 ; n49981_not
g100060 not n29686 ; n29686_not
g100061 not n17968 ; n17968_not
g100062 not n45868 ; n45868_not
g100063 not n17977 ; n17977_not
g100064 not n39298 ; n39298_not
g100065 not n53689 ; n53689_not
g100066 not n25897 ; n25897_not
g100067 not n27499 ; n27499_not
g100068 not n45589 ; n45589_not
g100069 not n29839 ; n29839_not
g100070 not n17986 ; n17986_not
g100071 not n47857 ; n47857_not
g100072 not n43798 ; n43798_not
g100073 not n25879 ; n25879_not
g100074 not n19597 ; n19597_not
g100075 not n39289 ; n39289_not
g100076 not n29866 ; n29866_not
g100077 not n38758 ; n38758_not
g100078 not n47974 ; n47974_not
g100079 not n36598 ; n36598_not
g100080 not n49990 ; n49990_not
g100081 not n56848 ; n56848_not
g100082 not n25888 ; n25888_not
g100083 not n29857 ; n29857_not
g100084 not n17959 ; n17959_not
g100085 not n29695 ; n29695_not
g100086 not n49837 ; n49837_not
g100087 not n29398 ; n29398_not
g100088 not n46984 ; n46984_not
g100089 not n52879 ; n52879_not
g100090 not n43888 ; n43888_not
g100091 not n56686 ; n56686_not
g100092 not n49828 ; n49828_not
g100093 not n48964 ; n48964_not
g100094 not n29488 ; n29488_not
g100095 not n49819 ; n49819_not
g100096 not n48577 ; n48577_not
g100097 not n29479 ; n29479_not
g100098 not n38668 ; n38668_not
g100099 not n46993 ; n46993_not
g100100 not n29389 ; n29389_not
g100101 not n19885 ; n19885_not
g100102 not n55669 ; n55669_not
g100103 not n43897 ; n43897_not
g100104 not n39379 ; n39379_not
g100105 not n49855 ; n49855_not
g100106 not n38857 ; n38857_not
g100107 not n36679 ; n36679_not
g100108 not n19849 ; n19849_not
g100109 not n38686 ; n38686_not
g100110 not n45499 ; n45499_not
g100111 not n29497 ; n29497_not
g100112 not n46975 ; n46975_not
g100113 not n49846 ; n49846_not
g100114 not n54994 ; n54994_not
g100115 not n56695 ; n56695_not
g100116 not n48568 ; n48568_not
g100117 not n38677 ; n38677_not
g100118 not n19867 ; n19867_not
g100119 not n48595 ; n48595_not
g100120 not n53779 ; n53779_not
g100121 not n55678 ; n55678_not
g100122 not n29299 ; n29299_not
g100123 not n38587 ; n38587_not
g100124 not n38875 ; n38875_not
g100125 not n49783 ; n49783_not
g100126 not n54985 ; n54985_not
g100127 not n19939 ; n19939_not
g100128 not n17698 ; n17698_not
g100129 not n55786 ; n55786_not
g100130 not n49774 ; n49774_not
g100131 not n34897 ; n34897_not
g100132 not n38866 ; n38866_not
g100133 not n19894 ; n19894_not
g100134 not n55948 ; n55948_not
g100135 not n56677 ; n56677_not
g100136 not n44599 ; n44599_not
g100137 not n38659 ; n38659_not
g100138 not n52888 ; n52888_not
g100139 not n17689 ; n17689_not
g100140 not n55957 ; n55957_not
g100141 not n55498 ; n55498_not
g100142 not n49792 ; n49792_not
g100143 not n47866 ; n47866_not
g100144 not n34879 ; n34879_not
g100145 not n49378 ; n49378_not
g100146 not n15898 ; n15898_not
g100147 not n48487 ; n48487_not
g100148 not n15889 ; n15889_not
g100149 not n25789 ; n25789_not
g100150 not n25699 ; n25699_not
g100151 not n17599 ; n17599_not
g100152 not n48496 ; n48496_not
g100153 not n49891 ; n49891_not
g100154 not n45886 ; n45886_not
g100155 not n48955 ; n48955_not
g100156 not n36769 ; n36769_not
g100157 not n56758 ; n56758_not
g100158 not a[13] ; a[13]_not
g100159 not n29749 ; n29749_not
g100160 not n49927 ; n49927_not
g100161 not n19768 ; n19768_not
g100162 not n38578 ; n38578_not
g100163 not n49918 ; n49918_not
g100164 not n49369 ; n49369_not
g100165 not n19777 ; n19777_not
g100166 not n49909 ; n49909_not
g100167 not n39388 ; n39388_not
g100168 not n29596 ; n29596_not
g100169 not n46948 ; n46948_not
g100170 not n49873 ; n49873_not
g100171 not n29587 ; n29587_not
g100172 not n43879 ; n43879_not
g100173 not n37399 ; n37399_not
g100174 not n29578 ; n29578_not
g100175 not n46957 ; n46957_not
g100176 not n38695 ; n38695_not
g100177 not n29569 ; n29569_not
g100178 not n47884 ; n47884_not
g100179 not n49864 ; n49864_not
g100180 not n36688 ; n36688_not
g100181 not n35995 ; n35995_not
g100182 not n34789 ; n34789_not
g100183 not n46966 ; n46966_not
g100184 not n19795 ; n19795_not
g100185 not n49882 ; n49882_not
g100186 not n35986 ; n35986_not
g100187 not n47893 ; n47893_not
g100188 not n45895 ; n45895_not
g100189 not n36697 ; n36697_not
g100190 not n46939 ; n46939_not
g100191 not n36958 ; n36958_not
g100192 not n18589 ; n18589_not
g100193 not n39577 ; n39577_not
g100194 not n36949 ; n36949_not
g100195 not n46597 ; n46597_not
g100196 not n57298 ; n57298_not
g100197 not n57289 ; n57289_not
g100198 not n53869 ; n53869_not
g100199 not n43978 ; n43978_not
g100200 not n53878 ; n53878_not
g100201 not n53887 ; n53887_not
g100202 not n48919 ; n48919_not
g100203 not n46669 ; n46669_not
g100204 not n53896 ; n53896_not
g100205 not n15799 ; n15799_not
g100206 not n43969 ; n43969_not
g100207 not n56884 ; n56884_not
g100208 not n53995 ; n53995_not
g100209 not n46588 ; n46588_not
g100210 not n55687 ; n55687_not
g100211 not n56839 ; n56839_not
g100212 not n45796 ; n45796_not
g100213 not n48289 ; n48289_not
g100214 not n46696 ; n46696_not
g100215 not n47668 ; n47668_not
g100216 not n43987 ; n43987_not
g100217 not n46678 ; n46678_not
g100218 not n53959 ; n53959_not
g100219 not n47947 ; n47947_not
g100220 not n53968 ; n53968_not
g100221 not n53599 ; n53599_not
g100222 not n53977 ; n53977_not
g100223 not n53986 ; n53986_not
g100224 not n46687 ; n46687_not
g100225 not n35878 ; n35878_not
g100226 not n31999 ; n31999_not
g100227 not n39469 ; n39469_not
g100228 not n56965 ; n56965_not
g100229 not n55858 ; n55858_not
g100230 not n56956 ; n56956_not
g100231 not n48748 ; n48748_not
g100232 not n53788 ; n53788_not
g100233 not n55399 ; n55399_not
g100234 not n47992 ; n47992_not
g100235 not n47659 ; n47659_not
g100236 not n39478 ; n39478_not
g100237 not n39559 ; n39559_not
g100238 not n57478 ; n57478_not
g100239 not n39487 ; n39487_not
g100240 not n56974 ; n56974_not
g100241 not n35887 ; n35887_not
g100242 not n32998 ; n32998_not
g100243 not n43996 ; n43996_not
g100244 not n56929 ; n56929_not
g100245 not n55867 ; n55867_not
g100246 not n32989 ; n32989_not
g100247 not n57388 ; n57388_not
g100248 not n35896 ; n35896_not
g100249 not n45778 ; n45778_not
g100250 not n57379 ; n57379_not
g100251 not n32899 ; n32899_not
g100252 not n53797 ; n53797_not
g100253 not n39496 ; n39496_not
g100254 not n39568 ; n39568_not
g100255 not n14998 ; n14998_not
g100256 not n35869 ; n35869_not
g100257 not n43699 ; n43699_not
g100258 not n48379 ; n48379_not
g100259 not n46795 ; n46795_not
g100260 not n29947 ; n29947_not
g100261 not n19399 ; n19399_not
g100262 not n48937 ; n48937_not
g100263 not n46786 ; n46786_not
g100264 not n38893 ; n38893_not
g100265 not n29938 ; n29938_not
g100266 not n56983 ; n56983_not
g100267 not n48388 ; n48388_not
g100268 not n33799 ; n33799_not
g100269 not n35968 ; n35968_not
g100270 not n48757 ; n48757_not
g100271 not n19498 ; n19498_not
g100272 not n48397 ; n48397_not
g100273 not n29956 ; n29956_not
g100274 not n38884 ; n38884_not
g100275 not n29983 ; n29983_not
g100276 not n29974 ; n29974_not
g100277 not n18598 ; n18598_not
g100278 not n56938 ; n56938_not
g100279 not n29965 ; n29965_not
g100280 not n19489 ; n19489_not
g100281 not n33988 ; n33988_not
g100282 not n36877 ; n36877_not
g100283 not n38965 ; n38965_not
g100284 not n39694 ; n39694_not
g100285 not n45688 ; n45688_not
g100286 not n55489 ; n55489_not
g100287 not n56749 ; n56749_not
g100288 not n38956 ; n38956_not
g100289 not n36868 ; n36868_not
g100290 not n38992 ; n38992_not
g100291 not n48298 ; n48298_not
g100292 not n38974 ; n38974_not
g100293 not n55885 ; n55885_not
g100294 not n36895 ; n36895_not
g100295 not n56794 ; n56794_not
g100296 not n38983 ; n38983_not
g100297 not n48928 ; n48928_not
g100298 not n36886 ; n36886_not
g100299 not n45679 ; n45679_not
g100300 not n46768 ; n46768_not
g100301 not n48892 ; n48892_not
g100302 not n55696 ; n55696_not
g100303 not n46777 ; n46777_not
g100304 not a[40] ; a[40]_not
g100305 not n38947 ; n38947_not
g100306 not n38479 ; n38479_not
g100307 not n36859 ; n36859_not
g100308 not n38938 ; n38938_not
g100309 not n35959 ; n35959_not
g100310 not n38488 ; n38488_not
g100311 not n46759 ; n46759_not
g100312 not n38929 ; n38929_not
g100313 not n28678 ; n28678_not
g100314 not n26779 ; n26779_not
g100315 not n55768 ; n55768_not
g100316 not n28669 ; n28669_not
g100317 not n26896 ; n26896_not
g100318 not n35797 ; n35797_not
g100319 not n26788 ; n26788_not
g100320 not n37579 ; n37579_not
g100321 not n28696 ; n28696_not
g100322 not n55993 ; n55993_not
g100323 not n39649 ; n39649_not
g100324 not n28687 ; n28687_not
g100325 not n55759 ; n55759_not
g100326 not n49549 ; n49549_not
g100327 not n16879 ; n16879_not
g100328 not n55966 ; n55966_not
g100329 not n42997 ; n42997_not
g100330 not n28597 ; n28597_not
g100331 not n37498 ; n37498_not
g100332 not n49495 ; n49495_not
g100333 not n48991 ; n48991_not
g100334 not n26797 ; n26797_not
g100335 not n27976 ; n27976_not
g100336 not n37588 ; n37588_not
g100337 not n54958 ; n54958_not
g100338 not n42988 ; n42988_not
g100339 not n35788 ; n35788_not
g100340 not n16888 ; n16888_not
g100341 not n27958 ; n27958_not
g100342 not n26995 ; n26995_not
g100343 not n48775 ; n48775_not
g100344 not n47749 ; n47749_not
g100345 not n13999 ; n13999_not
g100346 not n28786 ; n28786_not
g100347 not n48793 ; n48793_not
g100348 not n28777 ; n28777_not
g100349 not n27895 ; n27895_not
g100350 not n19858 ; n19858_not
g100351 not n35599 ; n35599_not
g100352 not n48856 ; n48856_not
g100353 not n39199 ; n39199_not
g100354 not n42979 ; n42979_not
g100355 not n28795 ; n28795_not
g100356 not n27886 ; n27886_not
g100357 not n45967 ; n45967_not
g100358 not n49576 ; n49576_not
g100359 not n27994 ; n27994_not
g100360 not n55777 ; n55777_not
g100361 not n49567 ; n49567_not
g100362 not n47569 ; n47569_not
g100363 not n49594 ; n49594_not
g100364 not n47578 ; n47578_not
g100365 not n16996 ; n16996_not
g100366 not n28768 ; n28768_not
g100367 not n42799 ; n42799_not
g100368 not n28759 ; n28759_not
g100369 not n49585 ; n49585_not
g100370 not n49558 ; n49558_not
g100371 not n45769 ; n45769_not
g100372 not n23998 ; n23998_not
g100373 not n45985 ; n45985_not
g100374 not n17797 ; n17797_not
g100375 not n27796 ; n27796_not
g100376 not n47767 ; n47767_not
g100377 not n51898 ; n51898_not
g100378 not n52978 ; n52978_not
g100379 not n37993 ; n37993_not
g100380 not n52996 ; n52996_not
g100381 not n27985 ; n27985_not
g100382 not n17779 ; n17779_not
g100383 not n16969 ; n16969_not
g100384 not n27778 ; n27778_not
g100385 not n26878 ; n26878_not
g100386 not n48847 ; n48847_not
g100387 not n37948 ; n37948_not
g100388 not n49288 ; n49288_not
g100389 not n37957 ; n37957_not
g100390 not n35779 ; n35779_not
g100391 not n37966 ; n37966_not
g100392 not n49279 ; n49279_not
g100393 not n26869 ; n26869_not
g100394 not n23989 ; n23989_not
g100395 not n26977 ; n26977_not
g100396 not n52987 ; n52987_not
g100397 not n47389 ; n47389_not
g100398 not n47776 ; n47776_not
g100399 not n49297 ; n49297_not
g100400 not n27859 ; n27859_not
g100401 not n27949 ; n27949_not
g100402 not n45994 ; n45994_not
g100403 not n37975 ; n37975_not
g100404 not n39667 ; n39667_not
g100405 not n47398 ; n47398_not
g100406 not n49477 ; n49477_not
g100407 not n42898 ; n42898_not
g100408 not n42889 ; n42889_not
g100409 not n16978 ; n16978_not
g100410 not n49459 ; n49459_not
g100411 not n45976 ; n45976_not
g100412 not n47785 ; n47785_not
g100413 not n49198 ; n49198_not
g100414 not n28588 ; n28588_not
g100415 not n52897 ; n52897_not
g100416 not n28579 ; n28579_not
g100417 not n16897 ; n16897_not
g100418 not n26887 ; n26887_not
g100419 not n49189 ; n49189_not
g100420 not n52969 ; n52969_not
g100421 not n54949 ; n54949_not
g100422 not n49387 ; n49387_not
g100423 not n35698 ; n35698_not
g100424 not n47758 ; n47758_not
g100425 not n28399 ; n28399_not
g100426 not n34798 ; n34798_not
g100427 not n48586 ; n48586_not
g100428 not n28498 ; n28498_not
g100429 not n28489 ; n28489_not
g100430 not n26986 ; n26986_not
g100431 not n39586 ; n39586_not
g100432 not n48829 ; n48829_not
g100433 not n28975 ; n28975_not
g100434 not n23899 ; n23899_not
g100435 not n19984 ; n19984_not
g100436 not n49684 ; n49684_not
g100437 not n19993 ; n19993_not
g100438 not n45949 ; n45949_not
g100439 not n28984 ; n28984_not
g100440 not n27688 ; n27688_not
g100441 not n37597 ; n37597_not
g100442 not n48667 ; n48667_not
g100443 not n39658 ; n39658_not
g100444 not n28993 ; n28993_not
g100445 not n45859 ; n45859_not
g100446 not n28948 ; n28948_not
g100447 not n49675 ; n49675_not
g100448 not n16789 ; n16789_not
g100449 not n55795 ; n55795_not
g100450 not n37984 ; n37984_not
g100451 not n28939 ; n28939_not
g100452 not a[31] ; a[31]_not
g100453 not n28966 ; n28966_not
g100454 not n48838 ; n48838_not
g100455 not n48658 ; n48658_not
g100456 not n19975 ; n19975_not
g100457 not n54967 ; n54967_not
g100458 not n47497 ; n47497_not
g100459 not n49747 ; n49747_not
g100460 not n37489 ; n37489_not
g100461 not n49468 ; n49468_not
g100462 not n49738 ; n49738_not
g100463 not n49729 ; n49729_not
g100464 not n16699 ; n16699_not
g100465 not n27697 ; n27697_not
g100466 not n49765 ; n49765_not
g100467 not n48874 ; n48874_not
g100468 not n19957 ; n19957_not
g100469 not n38299 ; n38299_not
g100470 not n49756 ; n49756_not
g100471 not n34888 ; n34888_not
g100472 not n48676 ; n48676_not
g100473 not n39676 ; n39676_not
g100474 not n48973 ; n48973_not
g100475 not n49693 ; n49693_not
g100476 not n16987 ; n16987_not
g100477 not n47596 ; n47596_not
g100478 not n38389 ; n38389_not
g100479 not n38398 ; n38398_not
g100480 not n47686 ; n47686_not
g100481 not n26599 ; n26599_not
g100482 not n38497 ; n38497_not
g100483 not n27589 ; n27589_not
g100484 not n28867 ; n28867_not
g100485 not n49639 ; n49639_not
g100486 not n28876 ; n28876_not
g100487 not n27679 ; n27679_not
g100488 not n55975 ; n55975_not
g100489 not n49099 ; n49099_not
g100490 not n34978 ; n34978_not
g100491 not n26959 ; n26959_not
g100492 not n27598 ; n27598_not
g100493 not n55876 ; n55876_not
g100494 not n47587 ; n47587_not
g100495 not a[22] ; a[22]_not
g100496 not n28894 ; n28894_not
g100497 not n48685 ; n48685_not
g100498 not n28885 ; n28885_not
g100499 not n26689 ; n26689_not
g100500 not n27868 ; n27868_not
g100501 not n34996 ; n34996_not
g100502 not n45958 ; n45958_not
g100503 not n28849 ; n28849_not
g100504 not n34987 ; n34987_not
g100505 not n36499 ; n36499_not
g100506 not n26698 ; n26698_not
g100507 not n17788 ; n17788_not
g100508 not n47479 ; n47479_not
g100509 not n28858 ; n28858_not
g100510 not n47695 ; n47695_not
g100511 not n48982 ; n48982_not
g100512 not n48865 ; n48865_not
g100513 not n49657 ; n49657_not
g100514 not n16798 ; n16798_not
g100515 not n49666 ; n49666_not
g100516 not n19948 ; n19948_not
g100517 not n34969 ; n34969_not
g100518 not n47488 ; n47488_not
g100519 not n49648 ; n49648_not
g100520 not b[13] ; b[13]_not
g100521 not n56795 ; n56795_not
g100522 not n39686 ; n39686_not
g100523 not n55787 ; n55787_not
g100524 not n44798 ; n44798_not
g100525 not n39974 ; n39974_not
g100526 not b[31] ; b[31]_not
g100527 not n39794 ; n39794_not
g100528 not n57497 ; n57497_not
g100529 not n39857 ; n39857_not
g100530 not n55868 ; n55868_not
g100531 not n45698 ; n45698_not
g100532 not n38678 ; n38678_not
g100533 not n38768 ; n38768_not
g100534 not n16997 ; n16997_not
g100535 not n39992 ; n39992_not
g100536 not n39776 ; n39776_not
g100537 not n39479 ; n39479_not
g100538 not n54878 ; n54878_not
g100539 not n16988 ; n16988_not
g100540 not n57299 ; n57299_not
g100541 not n39569 ; n39569_not
g100542 not n56975 ; n56975_not
g100543 not n14999 ; n14999_not
g100544 not n17789 ; n17789_not
g100545 not n45977 ; n45977_not
g100546 not n38759 ; n38759_not
g100547 not n15899 ; n15899_not
g100548 not n38687 ; n38687_not
g100549 not n54698 ; n54698_not
g100550 not n39848 ; n39848_not
g100551 not b[40] ; b[40]_not
g100552 not b[22] ; b[22]_not
g100553 not n39983 ; n39983_not
g100554 not n18869 ; n18869_not
g100555 not n45869 ; n45869_not
g100556 not n39785 ; n39785_not
g100557 not n45959 ; n45959_not
g100558 not n39839 ; n39839_not
g100559 not n39488 ; n39488_not
g100560 not n44699 ; n44699_not
g100561 not n46598 ; n46598_not
g100562 not n56786 ; n56786_not
g100563 not n56939 ; n56939_not
g100564 not n56984 ; n56984_not
g100565 not n18788 ; n18788_not
g100566 not n45779 ; n45779_not
g100567 not n39389 ; n39389_not
g100568 not n38669 ; n38669_not
g100569 not n38696 ; n38696_not
g100570 not n39578 ; n39578_not
g100571 not n42998 ; n42998_not
g100572 not n55796 ; n55796_not
g100573 not n45968 ; n45968_not
g100574 not n54599 ; n54599_not
g100575 not n54896 ; n54896_not
g100576 not n39596 ; n39596_not
g100577 not n39668 ; n39668_not
g100578 not n18797 ; n18797_not
g100579 not n54887 ; n54887_not
g100580 not n45788 ; n45788_not
g100581 not n39398 ; n39398_not
g100582 not n44789 ; n44789_not
g100583 not a[14] ; a[14]_not
g100584 not n45986 ; n45986_not
g100585 not n56876 ; n56876_not
g100586 not n39659 ; n39659_not
g100587 not n55877 ; n55877_not
g100588 not n17699 ; n17699_not
g100589 not n18779 ; n18779_not
g100590 not n42989 ; n42989_not
g100591 not n16979 ; n16979_not
g100592 not n39497 ; n39497_not
g100593 not n39299 ; n39299_not
g100594 not n42899 ; n42899_not
g100595 not n56885 ; n56885_not
g100596 not n39965 ; n39965_not
g100597 not n56894 ; n56894_not
g100598 not n56849 ; n56849_not
g100599 not n54689 ; n54689_not
g100600 not n55769 ; n55769_not
g100601 not n55778 ; n55778_not
g100602 not n45995 ; n45995_not
g100603 not n57398 ; n57398_not
g100604 not n56966 ; n56966_not
g100605 not n54869 ; n54869_not
g100606 not a[50] ; a[50]_not
g100607 not n16799 ; n16799_not
g100608 not n55598 ; n55598_not
g100609 not n55886 ; n55886_not
g100610 not n44888 ; n44888_not
g100611 not n56498 ; n56498_not
g100612 not n38939 ; n38939_not
g100613 not n56768 ; n56768_not
g100614 not n44987 ; n44987_not
g100615 not n54995 ; n54995_not
g100616 not n39677 ; n39677_not
g100617 not n55967 ; n55967_not
g100618 not n44978 ; n44978_not
g100619 not n38849 ; n38849_not
g100620 not n39749 ; n39749_not
g100621 not n44897 ; n44897_not
g100622 not n45689 ; n45689_not
g100623 not n54968 ; n54968_not
g100624 not n44996 ; n44996_not
g100625 not n39758 ; n39758_not
g100626 not n54797 ; n54797_not
g100627 not n55589 ; n55589_not
g100628 not n39866 ; n39866_not
g100629 not n54959 ; n54959_not
g100630 not n38777 ; n38777_not
g100631 not n56489 ; n56489_not
g100632 not n38795 ; n38795_not
g100633 not n17798 ; n17798_not
g100634 not n38948 ; n38948_not
g100635 not n45878 ; n45878_not
g100636 not n39929 ; n39929_not
g100637 not n44879 ; n44879_not
g100638 not n38786 ; n38786_not
g100639 not n38894 ; n38894_not
g100640 not n56678 ; n56678_not
g100641 not n15998 ; n15998_not
g100642 not n43889 ; n43889_not
g100643 not n38876 ; n38876_not
g100644 not n15989 ; n15989_not
g100645 not n39893 ; n39893_not
g100646 not n43898 ; n43898_not
g100647 not n39884 ; n39884_not
g100648 not n38885 ; n38885_not
g100649 not n55958 ; n55958_not
g100650 not n56669 ; n56669_not
g100651 not n55679 ; n55679_not
g100652 not n55688 ; n55688_not
g100653 not n55697 ; n55697_not
g100654 not n38867 ; n38867_not
g100655 not n44969 ; n44969_not
g100656 not n43799 ; n43799_not
g100657 not n45896 ; n45896_not
g100658 not n38858 ; n38858_not
g100659 not a[32] ; a[32]_not
g100660 not n56597 ; n56597_not
g100661 not n56588 ; n56588_not
g100662 not n39875 ; n39875_not
g100663 not n56579 ; n56579_not
g100664 not n56696 ; n56696_not
g100665 not n54977 ; n54977_not
g100666 not n56993 ; n56993_not
g100667 not n54788 ; n54788_not
g100668 not n39938 ; n39938_not
g100669 not n18689 ; n18689_not
g100670 not n54779 ; n54779_not
g100671 not n39947 ; n39947_not
g100672 not n55499 ; n55499_not
g100673 not a[23] ; a[23]_not
g100674 not n39587 ; n39587_not
g100675 not n39956 ; n39956_not
g100676 not n56759 ; n56759_not
g100677 not a[41] ; a[41]_not
g100678 not n18698 ; n18698_not
g100679 not n55895 ; n55895_not
g100680 not n56858 ; n56858_not
g100681 not n45599 ; n45599_not
g100682 not n55976 ; n55976_not
g100683 not n56399 ; n56399_not
g100684 not n38957 ; n38957_not
g100685 not n55985 ; n55985_not
g100686 not n38966 ; n38966_not
g100687 not n38984 ; n38984_not
g100688 not n39767 ; n39767_not
g100689 not n16898 ; n16898_not
g100690 not n56948 ; n56948_not
g100691 not n38993 ; n38993_not
g100692 not n16889 ; n16889_not
g100693 not n29885 ; n29885_not
g100694 not n47858 ; n47858_not
g100695 not n37679 ; n37679_not
g100696 not n19994 ; n19994_not
g100697 not n29894 ; n29894_not
g100698 not n37688 ; n37688_not
g100699 not n28769 ; n28769_not
g100700 not n19985 ; n19985_not
g100701 not n48956 ; n48956_not
g100702 not n37589 ; n37589_not
g100703 not n34898 ; n34898_not
g100704 not n52799 ; n52799_not
g100705 not n37949 ; n37949_not
g100706 not n37697 ; n37697_not
g100707 not n28778 ; n28778_not
g100708 not n47696 ; n47696_not
g100709 not n51989 ; n51989_not
g100710 not n29867 ; n29867_not
g100711 not n47768 ; n47768_not
g100712 not n47759 ; n47759_not
g100713 not n38597 ; n38597_not
g100714 not n38579 ; n38579_not
g100715 not n52997 ; n52997_not
g100716 not n19949 ; n19949_not
g100717 not n19967 ; n19967_not
g100718 not n48965 ; n48965_not
g100719 not n29876 ; n29876_not
g100720 not n51998 ; n51998_not
g100721 not n38489 ; n38489_not
g100722 not n49559 ; n49559_not
g100723 not n47867 ; n47867_not
g100724 not n49469 ; n49469_not
g100725 not n37598 ; n37598_not
g100726 not n49568 ; n49568_not
g100727 not n47669 ; n47669_not
g100728 not n48929 ; n48929_not
g100729 not n34889 ; n34889_not
g100730 not n28796 ; n28796_not
g100731 not n25979 ; n25979_not
g100732 not n19895 ; n19895_not
g100733 not n25988 ; n25988_not
g100734 not n25997 ; n25997_not
g100735 not n46994 ; n46994_not
g100736 not n29993 ; n29993_not
g100737 not n46985 ; n46985_not
g100738 not n46976 ; n46976_not
g100739 not n48947 ; n48947_not
g100740 not n37976 ; n37976_not
g100741 not n49478 ; n49478_not
g100742 not n47687 ; n47687_not
g100743 not n19958 ; n19958_not
g100744 not n36599 ; n36599_not
g100745 not n28787 ; n28787_not
g100746 not n47678 ; n47678_not
g100747 not n25889 ; n25889_not
g100748 not n37985 ; n37985_not
g100749 not n37994 ; n37994_not
g100750 not n25898 ; n25898_not
g100751 not n48938 ; n48938_not
g100752 not n47849 ; n47849_not
g100753 not n29957 ; n29957_not
g100754 not n48992 ; n48992_not
g100755 not n47894 ; n47894_not
g100756 not n46895 ; n46895_not
g100757 not n19769 ; n19769_not
g100758 not n52988 ; n52988_not
g100759 not n37499 ; n37499_not
g100760 not n52979 ; n52979_not
g100761 not n19787 ; n19787_not
g100762 not n38588 ; n38588_not
g100763 not n29966 ; n29966_not
g100764 not n29498 ; n29498_not
g100765 not n46868 ; n46868_not
g100766 not n29858 ; n29858_not
g100767 not n32999 ; n32999_not
g100768 not n52889 ; n52889_not
g100769 not n29849 ; n29849_not
g100770 not n46877 ; n46877_not
g100771 not n52898 ; n52898_not
g100772 not n29948 ; n29948_not
g100773 not n29489 ; n29489_not
g100774 not n46886 ; n46886_not
g100775 not n26987 ; n26987_not
g100776 not n23999 ; n23999_not
g100777 not n19877 ; n19877_not
g100778 not n48974 ; n48974_not
g100779 not n47777 ; n47777_not
g100780 not n28697 ; n28697_not
g100781 not n25799 ; n25799_not
g100782 not n29984 ; n29984_not
g100783 not n26996 ; n26996_not
g100784 not n28679 ; n28679_not
g100785 not n46949 ; n46949_not
g100786 not n48983 ; n48983_not
g100787 not n46958 ; n46958_not
g100788 not n47786 ; n47786_not
g100789 not n28688 ; n28688_not
g100790 not n46967 ; n46967_not
g100791 not n19859 ; n19859_not
g100792 not n27599 ; n27599_not
g100793 not n37868 ; n37868_not
g100794 not n28886 ; n28886_not
g100795 not n47399 ; n47399_not
g100796 not n48398 ; n48398_not
g100797 not n33989 ; n33989_not
g100798 not n48785 ; n48785_not
g100799 not n37958 ; n37958_not
g100800 not n48389 ; n48389_not
g100801 not n47579 ; n47579_not
g100802 not n48479 ; n48479_not
g100803 not n26969 ; n26969_not
g100804 not n37877 ; n37877_not
g100805 not n37886 ; n37886_not
g100806 not n48578 ; n48578_not
g100807 not n48587 ; n48587_not
g100808 not n33998 ; n33998_not
g100809 not n37859 ; n37859_not
g100810 not n37895 ; n37895_not
g100811 not n34979 ; n34979_not
g100812 not n47498 ; n47498_not
g100813 not n48677 ; n48677_not
g100814 not n47489 ; n47489_not
g100815 not n28958 ; n28958_not
g100816 not n26699 ; n26699_not
g100817 not n26798 ; n26798_not
g100818 not n48695 ; n48695_not
g100819 not n26789 ; n26789_not
g100820 not n28976 ; n28976_not
g100821 not n26897 ; n26897_not
g100822 not n28895 ; n28895_not
g100823 not n26888 ; n26888_not
g100824 not n26879 ; n26879_not
g100825 not n48668 ; n48668_not
g100826 not n48767 ; n48767_not
g100827 not n48299 ; n48299_not
g100828 not n50999 ; n50999_not
g100829 not n48758 ; n48758_not
g100830 not n46859 ; n46859_not
g100831 not n48875 ; n48875_not
g100832 not n28859 ; n28859_not
g100833 not n48866 ; n48866_not
g100834 not n28985 ; n28985_not
g100835 not n48776 ; n48776_not
g100836 not n46796 ; n46796_not
g100837 not n46787 ; n46787_not
g100838 not n46778 ; n46778_not
g100839 not n19778 ; n19778_not
g100840 not n46769 ; n46769_not
g100841 not n34997 ; n34997_not
g100842 not n19868 ; n19868_not
g100843 not n48893 ; n48893_not
g100844 not n37769 ; n37769_not
g100845 not n37778 ; n37778_not
g100846 not n48884 ; n48884_not
g100847 not n34988 ; n34988_not
g100848 not n48839 ; n48839_not
g100849 not n48497 ; n48497_not
g100850 not n37787 ; n37787_not
g100851 not n47597 ; n47597_not
g100852 not n37796 ; n37796_not
g100853 not n47588 ; n47588_not
g100854 not n48488 ; n48488_not
g100855 not n28877 ; n28877_not
g100856 not n48857 ; n48857_not
g100857 not n28868 ; n28868_not
g100858 not n36689 ; n36689_not
g100859 not n46697 ; n46697_not
g100860 not n48848 ; n48848_not
g100861 not n46688 ; n46688_not
g100862 not n46679 ; n46679_not
g100863 not n36968 ; n36968_not
g100864 not n47993 ; n47993_not
g100865 not n24899 ; n24899_not
g100866 not n49388 ; n49388_not
g100867 not n18968 ; n18968_not
g100868 not n29687 ; n29687_not
g100869 not n49379 ; n49379_not
g100870 not n18977 ; n18977_not
g100871 not n47984 ; n47984_not
g100872 not n47957 ; n47957_not
g100873 not n29696 ; n29696_not
g100874 not n18896 ; n18896_not
g100875 not n49298 ; n49298_not
g100876 not n24998 ; n24998_not
g100877 not n18959 ; n18959_not
g100878 not n18995 ; n18995_not
g100879 not n36995 ; n36995_not
g100880 not n47966 ; n47966_not
g100881 not n18986 ; n18986_not
g100882 not n29795 ; n29795_not
g100883 not n28589 ; n28589_not
g100884 not n47939 ; n47939_not
g100885 not n36986 ; n36986_not
g100886 not n47948 ; n47948_not
g100887 not n27896 ; n27896_not
g100888 not n49487 ; n49487_not
g100889 not n29669 ; n29669_not
g100890 not n27878 ; n27878_not
g100891 not n27779 ; n27779_not
g100892 not n28499 ; n28499_not
g100893 not n49199 ; n49199_not
g100894 not n29678 ; n29678_not
g100895 not n29759 ; n29759_not
g100896 not n27995 ; n27995_not
g100897 not n29777 ; n29777_not
g100898 not n38975 ; n38975_not
g100899 not n49397 ; n49397_not
g100900 not n48596 ; n48596_not
g100901 not n27986 ; n27986_not
g100902 not n29786 ; n29786_not
g100903 not n27959 ; n27959_not
g100904 not n27968 ; n27968_not
g100905 not n18878 ; n18878_not
g100906 not n36977 ; n36977_not
g100907 not n18887 ; n18887_not
g100908 not n27869 ; n27869_not
g100909 not n24989 ; n24989_not
g100910 not n38498 ; n38498_not
g100911 not n34799 ; n34799_not
g100912 not n47876 ; n47876_not
g100913 not n27689 ; n27689_not
g100914 not n27788 ; n27788_not
g100915 not n27698 ; n27698_not
g100916 not n48686 ; n48686_not
g100917 not n28598 ; n28598_not
g100918 not n29597 ; n29597_not
g100919 not n29688 ; n29688_not
g100920 not b[14] ; b[14]_not
g100921 not n54798 ; n54798_not
g100922 not n28977 ; n28977_not
g100923 not n39759 ; n39759_not
g100924 not n37896 ; n37896_not
g100925 not b[50] ; b[50]_not
g100926 not n24999 ; n24999_not
g100927 not b[32] ; b[32]_not
g100928 not n49857 ; n49857_not
g100929 not b[41] ; b[41]_not
g100930 not b[23] ; b[23]_not
g100931 not n49929 ; n49929_not
g100932 not n44979 ; n44979_not
g100933 not n48687 ; n48687_not
g100934 not n39975 ; n39975_not
g100935 not n54789 ; n54789_not
g100936 not n54879 ; n54879_not
g100937 not n49866 ; n49866_not
g100938 not n54987 ; n54987_not
g100939 not n36699 ; n36699_not
g100940 not n29697 ; n29697_not
g100941 not n56589 ; n56589_not
g100942 not n29787 ; n29787_not
g100943 not n25899 ; n25899_not
g100944 not n49695 ; n49695_not
g100945 not a[42] ; a[42]_not
g100946 not n49668 ; n49668_not
g100947 not n28995 ; n28995_not
g100948 not n36879 ; n36879_not
g100949 not n39966 ; n39966_not
g100950 not n44799 ; n44799_not
g100951 not n49677 ; n49677_not
g100952 not n36798 ; n36798_not
g100953 not n28959 ; n28959_not
g100954 not n49938 ; n49938_not
g100955 not n39993 ; n39993_not
g100956 not n48588 ; n48588_not
g100957 not n16989 ; n16989_not
g100958 not n45789 ; n45789_not
g100959 not n39678 ; n39678_not
g100960 not n45798 ; n45798_not
g100961 not n36897 ; n36897_not
g100962 not n16998 ; n16998_not
g100963 not n29769 ; n29769_not
g100964 not n37869 ; n37869_not
g100965 not n55698 ; n55698_not
g100966 not n39696 ; n39696_not
g100967 not n49686 ; n49686_not
g100968 not n49947 ; n49947_not
g100969 not n49893 ; n49893_not
g100970 not n39984 ; n39984_not
g100971 not n43998 ; n43998_not
g100972 not n48597 ; n48597_not
g100973 not n37878 ; n37878_not
g100974 not n55689 ; n55689_not
g100975 not n54969 ; n54969_not
g100976 not n56796 ; n56796_not
g100977 not n37887 ; n37887_not
g100978 not n39579 ; n39579_not
g100979 not n36789 ; n36789_not
g100980 not n37788 ; n37788_not
g100981 not n49956 ; n49956_not
g100982 not n48678 ; n48678_not
g100983 not n54888 ; n54888_not
g100984 not n56778 ; n56778_not
g100985 not n49875 ; n49875_not
g100986 not n28986 ; n28986_not
g100987 not n54978 ; n54978_not
g100988 not n56769 ; n56769_not
g100989 not n39669 ; n39669_not
g100990 not n37797 ; n37797_not
g100991 not n36888 ; n36888_not
g100992 not n29679 ; n29679_not
g100993 not n54897 ; n54897_not
g100994 not n47994 ; n47994_not
g100995 not n49884 ; n49884_not
g100996 not n15999 ; n15999_not
g100997 not n36969 ; n36969_not
g100998 not n39858 ; n39858_not
g100999 not n29598 ; n29598_not
g101000 not a[15] ; a[15]_not
g101001 not n29589 ; n29589_not
g101002 not n44988 ; n44988_not
g101003 not n47877 ; n47877_not
g101004 not n56868 ; n56868_not
g101005 not n49398 ; n49398_not
g101006 not n56976 ; n56976_not
g101007 not n45888 ; n45888_not
g101008 not n49992 ; n49992_not
g101009 not n16899 ; n16899_not
g101010 not n44997 ; n44997_not
g101011 not n47796 ; n47796_not
g101012 not n49767 ; n49767_not
g101013 not n55779 ; n55779_not
g101014 not n45879 ; n45879_not
g101015 not a[33] ; a[33]_not
g101016 not n47976 ; n47976_not
g101017 not n39939 ; n39939_not
g101018 not n49749 ; n49749_not
g101019 not n49983 ; n49983_not
g101020 not n39849 ; n39849_not
g101021 not n34899 ; n34899_not
g101022 not n47868 ; n47868_not
g101023 not n36996 ; n36996_not
g101024 not n49758 ; n49758_not
g101025 not n49389 ; n49389_not
g101026 not n54699 ; n54699_not
g101027 not n43899 ; n43899_not
g101028 not n47958 ; n47958_not
g101029 not n56985 ; n56985_not
g101030 not n47949 ; n47949_not
g101031 not n37599 ; n37599_not
g101032 not n39876 ; n39876_not
g101033 not n29958 ; n29958_not
g101034 not n49794 ; n49794_not
g101035 not n56679 ; n56679_not
g101036 not n39894 ; n39894_not
g101037 not n49848 ; n49848_not
g101038 not n29499 ; n29499_not
g101039 not n39885 ; n39885_not
g101040 not n47859 ; n47859_not
g101041 not n49839 ; n49839_not
g101042 not n56688 ; n56688_not
g101043 not n29994 ; n29994_not
g101044 not n49299 ; n49299_not
g101045 not n56958 ; n56958_not
g101046 not n39867 ; n39867_not
g101047 not n55797 ; n55797_not
g101048 not n49776 ; n49776_not
g101049 not n56886 ; n56886_not
g101050 not n29976 ; n29976_not
g101051 not n47886 ; n47886_not
g101052 not n49785 ; n49785_not
g101053 not n29967 ; n29967_not
g101054 not n56895 ; n56895_not
g101055 not n39948 ; n39948_not
g101056 not n49965 ; n49965_not
g101057 not n39777 ; n39777_not
g101058 not n49488 ; n49488_not
g101059 not n25989 ; n25989_not
g101060 not n25998 ; n25998_not
g101061 not n49479 ; n49479_not
g101062 not n39786 ; n39786_not
g101063 not n39597 ; n39597_not
g101064 not n37779 ; n37779_not
g101065 not n44889 ; n44889_not
g101066 not n39588 ; n39588_not
g101067 not n39957 ; n39957_not
g101068 not n56598 ; n56598_not
g101069 not n39768 ; n39768_not
g101070 not n44898 ; n44898_not
g101071 not n29985 ; n29985_not
g101072 not n37698 ; n37698_not
g101073 not n47967 ; n47967_not
g101074 not n37689 ; n37689_not
g101075 not n51999 ; n51999_not
g101076 not n36978 ; n36978_not
g101077 not n39687 ; n39687_not
g101078 not n49974 ; n49974_not
g101079 not n39795 ; n39795_not
g101080 not n43989 ; n43989_not
g101081 not n19689 ; n19689_not
g101082 not n38589 ; n38589_not
g101083 not n19698 ; n19698_not
g101084 not n26997 ; n26997_not
g101085 not n19797 ; n19797_not
g101086 not n55968 ; n55968_not
g101087 not n52989 ; n52989_not
g101088 not n53799 ; n53799_not
g101089 not n52998 ; n52998_not
g101090 not n19779 ; n19779_not
g101091 not n55995 ; n55995_not
g101092 not n38769 ; n38769_not
g101093 not n55977 ; n55977_not
g101094 not n48975 ; n48975_not
g101095 not n19869 ; n19869_not
g101096 not n38679 ; n38679_not
g101097 not n19599 ; n19599_not
g101098 not n28689 ; n28689_not
g101099 not n38688 ; n38688_not
g101100 not n38697 ; n38697_not
g101101 not n48984 ; n48984_not
g101102 not n38598 ; n38598_not
g101103 not n18969 ; n18969_not
g101104 not n35988 ; n35988_not
g101105 not n48696 ; n48696_not
g101106 not n38787 ; n38787_not
g101107 not n53889 ; n53889_not
g101108 not n35979 ; n35979_not
g101109 not n53898 ; n53898_not
g101110 not n55986 ; n55986_not
g101111 not n48993 ; n48993_not
g101112 not n35997 ; n35997_not
g101113 not n38778 ; n38778_not
g101114 not n18996 ; n18996_not
g101115 not n18987 ; n18987_not
g101116 not n18978 ; n18978_not
g101117 not n37986 ; n37986_not
g101118 not n48939 ; n48939_not
g101119 not n19959 ; n19959_not
g101120 not n19968 ; n19968_not
g101121 not n28779 ; n28779_not
g101122 not n48948 ; n48948_not
g101123 not n49596 ; n49596_not
g101124 not n37959 ; n37959_not
g101125 not n28797 ; n28797_not
g101126 not n49578 ; n49578_not
g101127 not n55887 ; n55887_not
g101128 not n37995 ; n37995_not
g101129 not n55599 ; n55599_not
g101130 not n28788 ; n28788_not
g101131 not n19977 ; n19977_not
g101132 not n48966 ; n48966_not
g101133 not n52899 ; n52899_not
g101134 not n28698 ; n28698_not
g101135 not n19887 ; n19887_not
g101136 not n19995 ; n19995_not
g101137 not n48957 ; n48957_not
g101138 not n49587 ; n49587_not
g101139 not a[60] ; a[60]_not
g101140 not n49569 ; n49569_not
g101141 not n38499 ; n38499_not
g101142 not n38976 ; n38976_not
g101143 not n38967 ; n38967_not
g101144 not n27996 ; n27996_not
g101145 not n38985 ; n38985_not
g101146 not n57489 ; n57489_not
g101147 not n38958 ; n38958_not
g101148 not n38994 ; n38994_not
g101149 not n27969 ; n27969_not
g101150 not n38949 ; n38949_not
g101151 not n27879 ; n27879_not
g101152 not n27978 ; n27978_not
g101153 not n18699 ; n18699_not
g101154 not a[24] ; a[24]_not
g101155 not n38859 ; n38859_not
g101156 not n38796 ; n38796_not
g101157 not n27789 ; n27789_not
g101158 not n18897 ; n18897_not
g101159 not n18888 ; n18888_not
g101160 not n18879 ; n18879_not
g101161 not n18789 ; n18789_not
g101162 not n56994 ; n56994_not
g101163 not n18798 ; n18798_not
g101164 not n57498 ; n57498_not
g101165 not n38895 ; n38895_not
g101166 not n38886 ; n38886_not
g101167 not n38877 ; n38877_not
g101168 not n38868 ; n38868_not
g101169 not n56949 ; n56949_not
g101170 not n27798 ; n27798_not
g101171 not n49497 ; n49497_not
g101172 not n27699 ; n27699_not
g101173 not n28599 ; n28599_not
g101174 not n35799 ; n35799_not
g101175 not n53979 ; n53979_not
g101176 not n35898 ; n35898_not
g101177 not n35889 ; n35889_not
g101178 not n53988 ; n53988_not
g101179 not n27888 ; n27888_not
g101180 not n53997 ; n53997_not
g101181 not n17799 ; n17799_not
g101182 not n28887 ; n28887_not
g101183 not n55878 ; n55878_not
g101184 not n48876 ; n48876_not
g101185 not n48768 ; n48768_not
g101186 not n55896 ; n55896_not
g101187 not n48867 ; n48867_not
g101188 not n19788 ; n19788_not
g101189 not n37968 ; n37968_not
g101190 not n48858 ; n48858_not
g101191 not n34989 ; n34989_not
g101192 not n17979 ; n17979_not
g101193 not n56859 ; n56859_not
g101194 not n49659 ; n49659_not
g101195 not n26889 ; n26889_not
g101196 not n48885 ; n48885_not
g101197 not n28896 ; n28896_not
g101198 not n48777 ; n48777_not
g101199 not n26898 ; n26898_not
g101200 not n55788 ; n55788_not
g101201 not n17898 ; n17898_not
g101202 not n26799 ; n26799_not
g101203 not n26979 ; n26979_not
g101204 not n28878 ; n28878_not
g101205 not n17889 ; n17889_not
g101206 not n28869 ; n28869_not
g101207 not n48795 ; n48795_not
g101208 not n48849 ; n48849_not
g101209 not n48786 ; n48786_not
g101210 not n56499 ; n56499_not
g101211 not n19878 ; n19878_not
g101212 not n34998 ; n34998_not
g101213 not n17997 ; n17997_not
g101214 not n45699 ; n45699_not
g101215 not a[51] ; a[51]_not
g101216 not n17988 ; n17988_not
g101217 not n48894 ; n48894_not
g101218 not n43999 ; n43999_not
g101219 not n29599 ; n29599_not
g101220 not n39976 ; n39976_not
g101221 not b[15] ; b[15]_not
g101222 not n48949 ; n48949_not
g101223 not b[33] ; b[33]_not
g101224 not n49669 ; n49669_not
g101225 not n54898 ; n54898_not
g101226 not b[24] ; b[24]_not
g101227 not n28969 ; n28969_not
g101228 not n28897 ; n28897_not
g101229 not n49399 ; n49399_not
g101230 not n35899 ; n35899_not
g101231 not n34999 ; n34999_not
g101232 not n27799 ; n27799_not
g101233 not n48598 ; n48598_not
g101234 not n28879 ; n28879_not
g101235 not n48688 ; n48688_not
g101236 not n27988 ; n27988_not
g101237 not b[42] ; b[42]_not
g101238 not n36898 ; n36898_not
g101239 not n49867 ; n49867_not
g101240 not b[60] ; b[60]_not
g101241 not n48697 ; n48697_not
g101242 not n54889 ; n54889_not
g101243 not n55789 ; n55789_not
g101244 not n49687 ; n49687_not
g101245 not n49885 ; n49885_not
g101246 not n27979 ; n27979_not
g101247 not n49894 ; n49894_not
g101248 not n48985 ; n48985_not
g101249 not n54979 ; n54979_not
g101250 not n48778 ; n48778_not
g101251 not n47968 ; n47968_not
g101252 not n28888 ; n28888_not
g101253 not n36979 ; n36979_not
g101254 not n28978 ; n28978_not
g101255 not n48994 ; n48994_not
g101256 not n27889 ; n27889_not
g101257 not n54988 ; n54988_not
g101258 not n49489 ; n49489_not
g101259 not n39985 ; n39985_not
g101260 not n49678 ; n49678_not
g101261 not n48958 ; n48958_not
g101262 not n36988 ; n36988_not
g101263 not n49876 ; n49876_not
g101264 not n47959 ; n47959_not
g101265 not n48787 ; n48787_not
g101266 not a[25] ; a[25]_not
g101267 not b[51] ; b[51]_not
g101268 not n48976 ; n48976_not
g101269 not n39994 ; n39994_not
g101270 not n44899 ; n44899_not
g101271 not n47977 ; n47977_not
g101272 not n48967 ; n48967_not
g101273 not n27898 ; n27898_not
g101274 not n39796 ; n39796_not
g101275 not n39787 ; n39787_not
g101276 not n39778 ; n39778_not
g101277 not n48895 ; n48895_not
g101278 not n39769 ; n39769_not
g101279 not n47869 ; n47869_not
g101280 not n49579 ; n49579_not
g101281 not n39967 ; n39967_not
g101282 not n39859 ; n39859_not
g101283 not n44989 ; n44989_not
g101284 not n44998 ; n44998_not
g101285 not n49696 ; n49696_not
g101286 not n47797 ; n47797_not
g101287 not n48886 ; n48886_not
g101288 not n49759 ; n49759_not
g101289 not n55897 ; n55897_not
g101290 not n28699 ; n28699_not
g101291 not n39895 ; n39895_not
g101292 not n28789 ; n28789_not
g101293 not n39886 ; n39886_not
g101294 not n39868 ; n39868_not
g101295 not n55888 ; n55888_not
g101296 not n39877 ; n39877_not
g101297 not n28798 ; n28798_not
g101298 not n56599 ; n56599_not
g101299 not n49588 ; n49588_not
g101300 not n48499 ; n48499_not
g101301 not n39958 ; n39958_not
g101302 not n39949 ; n39949_not
g101303 not n49597 ; n49597_not
g101304 not n36799 ; n36799_not
g101305 not n28996 ; n28996_not
g101306 not n26989 ; n26989_not
g101307 not n35989 ; n35989_not
g101308 not n55987 ; n55987_not
g101309 not n35998 ; n35998_not
g101310 not n49795 ; n49795_not
g101311 not n36889 ; n36889_not
g101312 not n28987 ; n28987_not
g101313 not n48796 ; n48796_not
g101314 not n49858 ; n49858_not
g101315 not n49849 ; n49849_not
g101316 not n55798 ; n55798_not
g101317 not n56698 ; n56698_not
g101318 not n55996 ; n55996_not
g101319 not n49498 ; n49498_not
g101320 not n48868 ; n48868_not
g101321 not n49768 ; n49768_not
g101322 not n55978 ; n55978_not
g101323 not n48859 ; n48859_not
g101324 not n54799 ; n54799_not
g101325 not n47887 ; n47887_not
g101326 not n48877 ; n48877_not
g101327 not n47878 ; n47878_not
g101328 not n49786 ; n49786_not
g101329 not a[34] ; a[34]_not
g101330 not n49777 ; n49777_not
g101331 not n19978 ; n19978_not
g101332 not n54997 ; n54997_not
g101333 not n37969 ; n37969_not
g101334 not n29986 ; n29986_not
g101335 not n56995 ; n56995_not
g101336 not n49984 ; n49984_not
g101337 not n38977 ; n38977_not
g101338 not n39697 ; n39697_not
g101339 not n29977 ; n29977_not
g101340 not n29995 ; n29995_not
g101341 not n37996 ; n37996_not
g101342 not n37897 ; n37897_not
g101343 not n37888 ; n37888_not
g101344 not n37879 ; n37879_not
g101345 not n49957 ; n49957_not
g101346 not n49975 ; n49975_not
g101347 not n19969 ; n19969_not
g101348 not n49966 ; n49966_not
g101349 not n47599 ; n47599_not
g101350 not n19897 ; n19897_not
g101351 not n47689 ; n47689_not
g101352 not n29968 ; n29968_not
g101353 not n47698 ; n47698_not
g101354 not n46996 ; n46996_not
g101355 not n56689 ; n56689_not
g101356 not n18799 ; n18799_not
g101357 not n19879 ; n19879_not
g101358 not n56986 ; n56986_not
g101359 not n46969 ; n46969_not
g101360 not n16999 ; n16999_not
g101361 not n46978 ; n46978_not
g101362 not n46987 ; n46987_not
g101363 not n56896 ; n56896_not
g101364 not n49993 ; n49993_not
g101365 not n39688 ; n39688_not
g101366 not n38599 ; n38599_not
g101367 not n39679 ; n39679_not
g101368 not n19987 ; n19987_not
g101369 not n46699 ; n46699_not
g101370 not n37699 ; n37699_not
g101371 not n39499 ; n39499_not
g101372 not n39589 ; n39589_not
g101373 not n46789 ; n46789_not
g101374 not n38995 ; n38995_not
g101375 not n19699 ; n19699_not
g101376 not n19798 ; n19798_not
g101377 not n39598 ; n39598_not
g101378 not n19789 ; n19789_not
g101379 not n46798 ; n46798_not
g101380 not n17899 ; n17899_not
g101381 not n37789 ; n37789_not
g101382 not n37978 ; n37978_not
g101383 not n37798 ; n37798_not
g101384 not n49939 ; n49939_not
g101385 not n56869 ; n56869_not
g101386 not a[43] ; a[43]_not
g101387 not a[52] ; a[52]_not
g101388 not n45799 ; n45799_not
g101389 not n49948 ; n49948_not
g101390 not n17989 ; n17989_not
g101391 not n46897 ; n46897_not
g101392 not n46888 ; n46888_not
g101393 not n46879 ; n46879_not
g101394 not n19888 ; n19888_not
g101395 not n56779 ; n56779_not
g101396 not n17998 ; n17998_not
g101397 not n29896 ; n29896_not
g101398 not n18979 ; n18979_not
g101399 not n18988 ; n18988_not
g101400 not n29887 ; n29887_not
g101401 not n18997 ; n18997_not
g101402 not n53899 ; n53899_not
g101403 not n29878 ; n29878_not
g101404 not a[16] ; a[16]_not
g101405 not n18898 ; n18898_not
g101406 not n29869 ; n29869_not
g101407 not n47986 ; n47986_not
g101408 not n45988 ; n45988_not
g101409 not n45898 ; n45898_not
g101410 not n47896 ; n47896_not
g101411 not n56878 ; n56878_not
g101412 not n45979 ; n45979_not
g101413 not n29797 ; n29797_not
g101414 not n53989 ; n53989_not
g101415 not n29788 ; n29788_not
g101416 not n56788 ; n56788_not
g101417 not n29779 ; n29779_not
g101418 not n18889 ; n18889_not
g101419 not n57499 ; n57499_not
g101420 not a[61] ; a[61]_not
g101421 not n53998 ; n53998_not
g101422 not n47788 ; n47788_not
g101423 not n56968 ; n56968_not
g101424 not n45997 ; n45997_not
g101425 not n56959 ; n56959_not
g101426 not n47779 ; n47779_not
g101427 not n45889 ; n45889_not
g101428 not b[43] ; b[43]_not
g101429 not b[34] ; b[34]_not
g101430 not b[16] ; b[16]_not
g101431 not n55988 ; n55988_not
g101432 not n19799 ; n19799_not
g101433 not b[25] ; b[25]_not
g101434 not n46997 ; n46997_not
g101435 not n19889 ; n19889_not
g101436 not n49499 ; n49499_not
g101437 not a[62] ; a[62]_not
g101438 not b[52] ; b[52]_not
g101439 not n55997 ; n55997_not
g101440 not n56996 ; n56996_not
g101441 not n49877 ; n49877_not
g101442 not n49787 ; n49787_not
g101443 not n55898 ; n55898_not
g101444 not n49679 ; n49679_not
g101445 not n49778 ; n49778_not
g101446 not n49697 ; n49697_not
g101447 not n48788 ; n48788_not
g101448 not n38888 ; n38888_not
g101449 not n38978 ; n38978_not
g101450 not n46799 ; n46799_not
g101451 not n49895 ; n49895_not
g101452 not n38699 ; n38699_not
g101453 not n49769 ; n49769_not
g101454 not n46988 ; n46988_not
g101455 not n38879 ; n38879_not
g101456 not n49886 ; n49886_not
g101457 not n46979 ; n46979_not
g101458 not n26999 ; n26999_not
g101459 not n49598 ; n49598_not
g101460 not a[26] ; a[26]_not
g101461 not a[53] ; a[53]_not
g101462 not n56879 ; n56879_not
g101463 not n49589 ; n49589_not
g101464 not n46889 ; n46889_not
g101465 not n35999 ; n35999_not
g101466 not n38789 ; n38789_not
g101467 not n19988 ; n19988_not
g101468 not n49688 ; n49688_not
g101469 not n38897 ; n38897_not
g101470 not n19979 ; n19979_not
g101471 not n56969 ; n56969_not
g101472 not n37979 ; n37979_not
g101473 not n48698 ; n48698_not
g101474 not n53999 ; n53999_not
g101475 not n28799 ; n28799_not
g101476 not n49796 ; n49796_not
g101477 not n49868 ; n49868_not
g101478 not n17999 ; n17999_not
g101479 not b[61] ; b[61]_not
g101480 not n49859 ; n49859_not
g101481 not n38798 ; n38798_not
g101482 not n19997 ; n19997_not
g101483 not n19898 ; n19898_not
g101484 not n46898 ; n46898_not
g101485 not n39869 ; n39869_not
g101486 not n29996 ; n29996_not
g101487 not n29969 ; n29969_not
g101488 not n47789 ; n47789_not
g101489 not n47879 ; n47879_not
g101490 not n45899 ; n45899_not
g101491 not n56978 ; n56978_not
g101492 not n45989 ; n45989_not
g101493 not n39797 ; n39797_not
g101494 not n39788 ; n39788_not
g101495 not n27989 ; n27989_not
g101496 not n49994 ; n49994_not
g101497 not n39779 ; n39779_not
g101498 not n45998 ; n45998_not
g101499 not n47897 ; n47897_not
g101500 not n29978 ; n29978_not
g101501 not n29987 ; n29987_not
g101502 not n47888 ; n47888_not
g101503 not n39896 ; n39896_not
g101504 not n39887 ; n39887_not
g101505 not n47798 ; n47798_not
g101506 not n39878 ; n39878_not
g101507 not n49985 ; n49985_not
g101508 not n49976 ; n49976_not
g101509 not n56699 ; n56699_not
g101510 not n47699 ; n47699_not
g101511 not n38987 ; n38987_not
g101512 not n36998 ; n36998_not
g101513 not n47978 ; n47978_not
g101514 not n29699 ; n29699_not
g101515 not n36899 ; n36899_not
g101516 not n47969 ; n47969_not
g101517 not n47996 ; n47996_not
g101518 not n39995 ; n39995_not
g101519 not n39986 ; n39986_not
g101520 not n39977 ; n39977_not
g101521 not n56798 ; n56798_not
g101522 not n39968 ; n39968_not
g101523 not a[35] ; a[35]_not
g101524 not n39959 ; n39959_not
g101525 not a[17] ; a[17]_not
g101526 not n47987 ; n47987_not
g101527 not n27899 ; n27899_not
g101528 not n39599 ; n39599_not
g101529 not n29879 ; n29879_not
g101530 not n36989 ; n36989_not
g101531 not n29888 ; n29888_not
g101532 not n56888 ; n56888_not
g101533 not n56789 ; n56789_not
g101534 not n49949 ; n49949_not
g101535 not n27998 ; n27998_not
g101536 not n48797 ; n48797_not
g101537 not n37988 ; n37988_not
g101538 not n28889 ; n28889_not
g101539 not n54989 ; n54989_not
g101540 not n49967 ; n49967_not
g101541 not n38969 ; n38969_not
g101542 not n28997 ; n28997_not
g101543 not n49958 ; n49958_not
g101544 not n39689 ; n39689_not
g101545 not n39698 ; n39698_not
g101546 not n28979 ; n28979_not
g101547 not a[44] ; a[44]_not
g101548 not n54998 ; n54998_not
g101549 not n28988 ; n28988_not
g101550 not b[17] ; b[17]_not
g101551 not b[53] ; b[53]_not
g101552 not b[44] ; b[44]_not
g101553 not b[62] ; b[62]_not
g101554 not b[26] ; b[26]_not
g101555 not n48996 ; n48996_not
g101556 not b[35] ; b[35]_not
g101557 not n48987 ; n48987_not
g101558 not a[63] ; a[63]_not
g101559 not n48969 ; n48969_not
g101560 not n48978 ; n48978_not
g101561 not n56979 ; n56979_not
g101562 not n49698 ; n49698_not
g101563 not n49968 ; n49968_not
g101564 not n49977 ; n49977_not
g101565 not n56997 ; n56997_not
g101566 not n56988 ; n56988_not
g101567 not n49986 ; n49986_not
g101568 not n49995 ; n49995_not
g101569 not n49779 ; n49779_not
g101570 not a[45] ; a[45]_not
g101571 not n49869 ; n49869_not
g101572 not n49878 ; n49878_not
g101573 not n49887 ; n49887_not
g101574 not n49896 ; n49896_not
g101575 not n49959 ; n49959_not
g101576 not n49689 ; n49689_not
g101577 not a[36] ; a[36]_not
g101578 not n49788 ; n49788_not
g101579 not n49797 ; n49797_not
g101580 not n56898 ; n56898_not
g101581 not n29898 ; n29898_not
g101582 not n29889 ; n29889_not
g101583 not n48888 ; n48888_not
g101584 not n48879 ; n48879_not
g101585 not a[27] ; a[27]_not
g101586 not n55998 ; n55998_not
g101587 not n48897 ; n48897_not
g101588 not n28899 ; n28899_not
g101589 not n56799 ; n56799_not
g101590 not n56889 ; n56889_not
g101591 not a[54] ; a[54]_not
g101592 not n49599 ; n49599_not
g101593 not n46899 ; n46899_not
g101594 not n46989 ; n46989_not
g101595 not n46998 ; n46998_not
g101596 not n47889 ; n47889_not
g101597 not n37998 ; n37998_not
g101598 not n38979 ; n38979_not
g101599 not n38988 ; n38988_not
g101600 not n19899 ; n19899_not
g101601 not n36999 ; n36999_not
g101602 not n47979 ; n47979_not
g101603 not n47988 ; n47988_not
g101604 not n47898 ; n47898_not
g101605 not n37989 ; n37989_not
g101606 not n19989 ; n19989_not
g101607 not n19998 ; n19998_not
g101608 not n39699 ; n39699_not
g101609 not n54999 ; n54999_not
g101610 not n47799 ; n47799_not
g101611 not n37899 ; n37899_not
g101612 not a[18] ; a[18]_not
g101613 not n48798 ; n48798_not
g101614 not n47997 ; n47997_not
g101615 not n27999 ; n27999_not
g101616 not n38799 ; n38799_not
g101617 not n38889 ; n38889_not
g101618 not n38898 ; n38898_not
g101619 not n45999 ; n45999_not
g101620 not n38997 ; n38997_not
g101621 not n18999 ; n18999_not
g101622 not b[18] ; b[18]_not
g101623 not n29998 ; n29998_not
g101624 not b[27] ; b[27]_not
g101625 not b[36] ; b[36]_not
g101626 not n48889 ; n48889_not
g101627 not b[45] ; b[45]_not
g101628 not n48997 ; n48997_not
g101629 not n47989 ; n47989_not
g101630 not b[54] ; b[54]_not
g101631 not n48898 ; n48898_not
g101632 not b[63] ; b[63]_not
g101633 not a[46] ; a[46]_not
g101634 not n47998 ; n47998_not
g101635 not a[19] ; a[19]_not
g101636 not n48979 ; n48979_not
g101637 not n39979 ; n39979_not
g101638 not n39988 ; n39988_not
g101639 not n38989 ; n38989_not
g101640 not n56989 ; n56989_not
g101641 not n39799 ; n39799_not
g101642 not n48988 ; n48988_not
g101643 not n38899 ; n38899_not
g101644 not n56998 ; n56998_not
g101645 not n39997 ; n39997_not
g101646 not a[55] ; a[55]_not
g101647 not n19999 ; n19999_not
g101648 not n56899 ; n56899_not
g101649 not n39889 ; n39889_not
g101650 not n47899 ; n47899_not
g101651 not n37999 ; n37999_not
g101652 not n39898 ; n39898_not
g101653 not a[37] ; a[37]_not
g101654 not n38998 ; n38998_not
g101655 not n29989 ; n29989_not
g101656 not a[28] ; a[28]_not
g101657 not n49997 ; n49997_not
g101658 not n49979 ; n49979_not
g101659 not b[28] ; b[28]_not
g101660 not n49799 ; n49799_not
g101661 not b[55] ; b[55]_not
g101662 not b[37] ; b[37]_not
g101663 not n29999 ; n29999_not
g101664 not b[19] ; b[19]_not
g101665 not n49889 ; n49889_not
g101666 not b[46] ; b[46]_not
g101667 not n47999 ; n47999_not
g101668 not n48998 ; n48998_not
g101669 not n49988 ; n49988_not
g101670 not n39998 ; n39998_not
g101671 not a[38] ; a[38]_not
g101672 not n48989 ; n48989_not
g101673 not n39899 ; n39899_not
g101674 not n56999 ; n56999_not
g101675 not n39989 ; n39989_not
g101676 not n49898 ; n49898_not
g101677 not n48899 ; n48899_not
g101678 not a[56] ; a[56]_not
g101679 not n38999 ; n38999_not
g101680 not a[29] ; a[29]_not
g101681 not a[47] ; a[47]_not
g101682 not b[29] ; b[29]_not
g101683 not b[38] ; b[38]_not
g101684 not b[47] ; b[47]_not
g101685 not a[48] ; a[48]_not
g101686 not b[56] ; b[56]_not
g101687 not a[57] ; a[57]_not
g101688 not n49998 ; n49998_not
g101689 not n49989 ; n49989_not
g101690 not a[39] ; a[39]_not
g101691 not n39999 ; n39999_not
g101692 not n49899 ; n49899_not
g101693 not b[39] ; b[39]_not
g101694 not b[48] ; b[48]_not
g101695 not a[49] ; a[49]_not
g101696 not b[57] ; b[57]_not
g101697 not n49999 ; n49999_not
g101698 not a[58] ; a[58]_not
g101699 not b[49] ; b[49]_not
g101700 not b[58] ; b[58]_not
g101701 not a[59] ; a[59]_not
g101702 not b[59] ; b[59]_not
g101703 not quotient[6] ; quotient[6]_not
g101704 not quotient[9] ; quotient[9]_not
g101705 not quotient[30] ; quotient[30]_not
g101706 not quotient[12] ; quotient[12]_not
g101707 not quotient[21] ; quotient[21]_not
g101708 not quotient[50] ; quotient[50]_not
g101709 not quotient[23] ; quotient[23]_not
g101710 not quotient[32] ; quotient[32]_not
g101711 not quotient[41] ; quotient[41]_not
g101712 not quotient[24] ; quotient[24]_not
g101713 not quotient[51] ; quotient[51]_not
g101714 not quotient[15] ; quotient[15]_not
g101715 not quotient[60] ; quotient[60]_not
g101716 not quotient[33] ; quotient[33]_not
g101717 not quotient[42] ; quotient[42]_not
g101718 not quotient[35] ; quotient[35]_not
g101719 not quotient[26] ; quotient[26]_not
g101720 not quotient[44] ; quotient[44]_not
g101721 not quotient[53] ; quotient[53]_not
g101722 not quotient[36] ; quotient[36]_not
g101723 not quotient[45] ; quotient[45]_not
g101724 not quotient[18] ; quotient[18]_not
g101725 not quotient[27] ; quotient[27]_not
g101726 not quotient[54] ; quotient[54]_not
g101727 not quotient[56] ; quotient[56]_not
g101728 not quotient[29] ; quotient[29]_not
g101729 not quotient[38] ; quotient[38]_not
g101730 not quotient[47] ; quotient[47]_not
g101731 not quotient[39] ; quotient[39]_not
g101732 not quotient[48] ; quotient[48]_not
g101733 not quotient[57] ; quotient[57]_not
o quotient[0]
o quotient[59]
o quotient[62]
o quotient[63]
o remainder[0]
o remainder[1]
o remainder[2]
o remainder[3]
o remainder[4]
o remainder[5]
o remainder[6]
o remainder[7]
o remainder[8]
o remainder[9]
o remainder[10]
o remainder[11]
o remainder[12]
o remainder[13]
o remainder[14]
o remainder[15]
o remainder[16]
o remainder[17]
o remainder[18]
o remainder[19]
o remainder[20]
o remainder[21]
o remainder[22]
o remainder[23]
o remainder[24]
o remainder[25]
o remainder[26]
o remainder[27]
o remainder[28]
o remainder[29]
o remainder[30]
o remainder[31]
o remainder[32]
o remainder[33]
o remainder[34]
o remainder[35]
o remainder[36]
o remainder[37]
o remainder[38]
o remainder[39]
o remainder[40]
o remainder[41]
o remainder[42]
o remainder[43]
o remainder[44]
o remainder[45]
o remainder[46]
o remainder[47]
o remainder[48]
o remainder[49]
o remainder[50]
o remainder[51]
o remainder[52]
o remainder[53]
o remainder[54]
o remainder[55]
o remainder[56]
o remainder[57]
o remainder[58]
o remainder[59]
o remainder[60]
o remainder[61]
o remainder[62]
o remainder[63]
